module tt_um_corey (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire _15494_;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire _15551_;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire _15622_;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire _15631_;
 wire _15632_;
 wire _15633_;
 wire _15634_;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire _15658_;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire _15705_;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire _15714_;
 wire _15715_;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire _15735_;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire _15754_;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire _15759_;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire _15773_;
 wire _15774_;
 wire _15775_;
 wire _15776_;
 wire _15777_;
 wire _15778_;
 wire _15779_;
 wire _15780_;
 wire _15781_;
 wire _15782_;
 wire _15783_;
 wire _15784_;
 wire _15785_;
 wire _15786_;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15803_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15808_;
 wire _15809_;
 wire _15810_;
 wire _15811_;
 wire _15812_;
 wire _15813_;
 wire _15814_;
 wire _15815_;
 wire _15816_;
 wire _15817_;
 wire _15818_;
 wire _15819_;
 wire _15820_;
 wire _15821_;
 wire _15822_;
 wire _15823_;
 wire _15824_;
 wire _15825_;
 wire _15826_;
 wire _15827_;
 wire _15828_;
 wire _15829_;
 wire _15830_;
 wire _15831_;
 wire _15832_;
 wire _15833_;
 wire _15834_;
 wire _15835_;
 wire _15836_;
 wire _15837_;
 wire _15838_;
 wire _15839_;
 wire _15840_;
 wire _15841_;
 wire _15842_;
 wire _15843_;
 wire _15844_;
 wire _15845_;
 wire _15846_;
 wire _15847_;
 wire _15848_;
 wire _15849_;
 wire _15850_;
 wire _15851_;
 wire _15852_;
 wire _15853_;
 wire _15854_;
 wire _15855_;
 wire _15856_;
 wire _15857_;
 wire _15858_;
 wire _15859_;
 wire _15860_;
 wire _15861_;
 wire _15862_;
 wire _15863_;
 wire _15864_;
 wire _15865_;
 wire _15866_;
 wire _15867_;
 wire _15868_;
 wire _15869_;
 wire _15870_;
 wire _15871_;
 wire _15872_;
 wire _15873_;
 wire _15874_;
 wire _15875_;
 wire _15876_;
 wire _15877_;
 wire _15878_;
 wire _15879_;
 wire _15880_;
 wire _15881_;
 wire _15882_;
 wire _15883_;
 wire _15884_;
 wire _15885_;
 wire _15886_;
 wire _15887_;
 wire _15888_;
 wire _15889_;
 wire _15890_;
 wire _15891_;
 wire _15892_;
 wire _15893_;
 wire _15894_;
 wire _15895_;
 wire _15896_;
 wire _15897_;
 wire _15898_;
 wire _15899_;
 wire _15900_;
 wire _15901_;
 wire _15902_;
 wire _15903_;
 wire _15904_;
 wire _15905_;
 wire _15906_;
 wire _15907_;
 wire _15908_;
 wire _15909_;
 wire _15910_;
 wire _15911_;
 wire _15912_;
 wire _15913_;
 wire _15914_;
 wire _15915_;
 wire _15916_;
 wire _15917_;
 wire _15918_;
 wire _15919_;
 wire _15920_;
 wire _15921_;
 wire _15922_;
 wire _15923_;
 wire _15924_;
 wire _15925_;
 wire _15926_;
 wire _15927_;
 wire _15928_;
 wire _15929_;
 wire _15930_;
 wire _15931_;
 wire _15932_;
 wire _15933_;
 wire _15934_;
 wire _15935_;
 wire _15936_;
 wire _15937_;
 wire _15938_;
 wire _15939_;
 wire _15940_;
 wire _15941_;
 wire _15942_;
 wire _15943_;
 wire _15944_;
 wire _15945_;
 wire _15946_;
 wire _15947_;
 wire _15948_;
 wire _15949_;
 wire _15950_;
 wire _15951_;
 wire _15952_;
 wire _15953_;
 wire _15954_;
 wire _15955_;
 wire _15956_;
 wire _15957_;
 wire _15958_;
 wire _15959_;
 wire _15960_;
 wire _15961_;
 wire _15962_;
 wire _15963_;
 wire _15964_;
 wire _15965_;
 wire _15966_;
 wire _15967_;
 wire _15968_;
 wire _15969_;
 wire _15970_;
 wire _15971_;
 wire _15972_;
 wire _15973_;
 wire _15974_;
 wire _15975_;
 wire _15976_;
 wire _15977_;
 wire _15978_;
 wire _15979_;
 wire _15980_;
 wire _15981_;
 wire _15982_;
 wire _15983_;
 wire _15984_;
 wire _15985_;
 wire _15986_;
 wire _15987_;
 wire _15988_;
 wire _15989_;
 wire _15990_;
 wire _15991_;
 wire _15992_;
 wire _15993_;
 wire _15994_;
 wire _15995_;
 wire _15996_;
 wire _15997_;
 wire _15998_;
 wire _15999_;
 wire _16000_;
 wire _16001_;
 wire _16002_;
 wire _16003_;
 wire _16004_;
 wire _16005_;
 wire _16006_;
 wire _16007_;
 wire _16008_;
 wire _16009_;
 wire _16010_;
 wire _16011_;
 wire _16012_;
 wire _16013_;
 wire _16014_;
 wire _16015_;
 wire _16016_;
 wire _16017_;
 wire _16018_;
 wire _16019_;
 wire _16020_;
 wire _16021_;
 wire _16022_;
 wire _16023_;
 wire _16024_;
 wire _16025_;
 wire _16026_;
 wire _16027_;
 wire _16028_;
 wire _16029_;
 wire _16030_;
 wire _16031_;
 wire _16032_;
 wire _16033_;
 wire _16034_;
 wire _16035_;
 wire _16036_;
 wire _16037_;
 wire _16038_;
 wire _16039_;
 wire _16040_;
 wire _16041_;
 wire _16042_;
 wire _16043_;
 wire _16044_;
 wire _16045_;
 wire _16046_;
 wire _16047_;
 wire _16048_;
 wire _16049_;
 wire _16050_;
 wire _16051_;
 wire _16052_;
 wire _16053_;
 wire _16054_;
 wire _16055_;
 wire _16056_;
 wire _16057_;
 wire _16058_;
 wire _16059_;
 wire _16060_;
 wire _16061_;
 wire _16062_;
 wire _16063_;
 wire _16064_;
 wire _16065_;
 wire _16066_;
 wire _16067_;
 wire _16068_;
 wire _16069_;
 wire _16070_;
 wire _16071_;
 wire _16072_;
 wire _16073_;
 wire _16074_;
 wire _16075_;
 wire _16076_;
 wire _16077_;
 wire _16078_;
 wire _16079_;
 wire _16080_;
 wire _16081_;
 wire _16082_;
 wire _16083_;
 wire _16084_;
 wire _16085_;
 wire _16086_;
 wire _16087_;
 wire _16088_;
 wire _16089_;
 wire _16090_;
 wire _16091_;
 wire _16092_;
 wire _16093_;
 wire _16094_;
 wire _16095_;
 wire _16096_;
 wire _16097_;
 wire _16098_;
 wire _16099_;
 wire _16100_;
 wire _16101_;
 wire _16102_;
 wire _16103_;
 wire _16104_;
 wire _16105_;
 wire _16106_;
 wire _16107_;
 wire _16108_;
 wire _16109_;
 wire _16110_;
 wire _16111_;
 wire _16112_;
 wire _16113_;
 wire _16114_;
 wire _16115_;
 wire _16116_;
 wire _16117_;
 wire _16118_;
 wire _16119_;
 wire _16120_;
 wire _16121_;
 wire _16122_;
 wire _16123_;
 wire _16124_;
 wire _16125_;
 wire _16126_;
 wire _16127_;
 wire _16128_;
 wire _16129_;
 wire _16130_;
 wire _16131_;
 wire _16132_;
 wire _16133_;
 wire _16134_;
 wire _16135_;
 wire _16136_;
 wire _16137_;
 wire _16138_;
 wire _16139_;
 wire _16140_;
 wire _16141_;
 wire _16142_;
 wire _16143_;
 wire _16144_;
 wire _16145_;
 wire _16146_;
 wire _16147_;
 wire _16148_;
 wire _16149_;
 wire _16150_;
 wire _16151_;
 wire _16152_;
 wire _16153_;
 wire _16154_;
 wire _16155_;
 wire _16156_;
 wire _16157_;
 wire _16158_;
 wire _16159_;
 wire _16160_;
 wire _16161_;
 wire _16162_;
 wire _16163_;
 wire _16164_;
 wire _16165_;
 wire _16166_;
 wire _16167_;
 wire _16168_;
 wire _16169_;
 wire _16170_;
 wire _16171_;
 wire _16172_;
 wire _16173_;
 wire _16174_;
 wire _16175_;
 wire _16176_;
 wire _16177_;
 wire _16178_;
 wire _16179_;
 wire _16180_;
 wire _16181_;
 wire _16182_;
 wire _16183_;
 wire _16184_;
 wire _16185_;
 wire _16186_;
 wire _16187_;
 wire _16188_;
 wire _16189_;
 wire _16190_;
 wire _16191_;
 wire _16192_;
 wire _16193_;
 wire _16194_;
 wire _16195_;
 wire _16196_;
 wire _16197_;
 wire _16198_;
 wire _16199_;
 wire _16200_;
 wire _16201_;
 wire _16202_;
 wire _16203_;
 wire _16204_;
 wire _16205_;
 wire _16206_;
 wire _16207_;
 wire _16208_;
 wire _16209_;
 wire _16210_;
 wire _16211_;
 wire _16212_;
 wire _16213_;
 wire _16214_;
 wire _16215_;
 wire _16216_;
 wire _16217_;
 wire _16218_;
 wire _16219_;
 wire _16220_;
 wire _16221_;
 wire _16222_;
 wire _16223_;
 wire _16224_;
 wire _16225_;
 wire _16226_;
 wire _16227_;
 wire _16228_;
 wire _16229_;
 wire _16230_;
 wire _16231_;
 wire _16232_;
 wire _16233_;
 wire _16234_;
 wire _16235_;
 wire _16236_;
 wire _16237_;
 wire _16238_;
 wire _16239_;
 wire _16240_;
 wire _16241_;
 wire _16242_;
 wire _16243_;
 wire _16244_;
 wire _16245_;
 wire _16246_;
 wire _16247_;
 wire _16248_;
 wire _16249_;
 wire _16250_;
 wire _16251_;
 wire _16252_;
 wire _16253_;
 wire _16254_;
 wire _16255_;
 wire _16256_;
 wire _16257_;
 wire _16258_;
 wire _16259_;
 wire _16260_;
 wire _16261_;
 wire _16262_;
 wire _16263_;
 wire _16264_;
 wire _16265_;
 wire _16266_;
 wire _16267_;
 wire _16268_;
 wire _16269_;
 wire _16270_;
 wire _16271_;
 wire _16272_;
 wire _16273_;
 wire _16274_;
 wire _16275_;
 wire _16276_;
 wire _16277_;
 wire _16278_;
 wire _16279_;
 wire _16280_;
 wire _16281_;
 wire _16282_;
 wire _16283_;
 wire _16284_;
 wire _16285_;
 wire _16286_;
 wire _16287_;
 wire _16288_;
 wire _16289_;
 wire _16290_;
 wire _16291_;
 wire _16292_;
 wire _16293_;
 wire _16294_;
 wire _16295_;
 wire _16296_;
 wire _16297_;
 wire _16298_;
 wire _16299_;
 wire _16300_;
 wire _16301_;
 wire _16302_;
 wire _16303_;
 wire _16304_;
 wire _16305_;
 wire _16306_;
 wire _16307_;
 wire _16308_;
 wire _16309_;
 wire _16310_;
 wire _16311_;
 wire _16312_;
 wire _16313_;
 wire _16314_;
 wire _16315_;
 wire _16316_;
 wire _16317_;
 wire _16318_;
 wire _16319_;
 wire _16320_;
 wire _16321_;
 wire _16322_;
 wire _16323_;
 wire _16324_;
 wire _16325_;
 wire _16326_;
 wire _16327_;
 wire _16328_;
 wire _16329_;
 wire _16330_;
 wire _16331_;
 wire _16332_;
 wire _16333_;
 wire _16334_;
 wire _16335_;
 wire _16336_;
 wire _16337_;
 wire _16338_;
 wire _16339_;
 wire _16340_;
 wire _16341_;
 wire _16342_;
 wire _16343_;
 wire _16344_;
 wire _16345_;
 wire _16346_;
 wire _16347_;
 wire _16348_;
 wire _16349_;
 wire _16350_;
 wire _16351_;
 wire _16352_;
 wire _16353_;
 wire _16354_;
 wire _16355_;
 wire _16356_;
 wire _16357_;
 wire _16358_;
 wire _16359_;
 wire _16360_;
 wire _16361_;
 wire _16362_;
 wire _16363_;
 wire _16364_;
 wire _16365_;
 wire _16366_;
 wire _16367_;
 wire _16368_;
 wire _16369_;
 wire _16370_;
 wire _16371_;
 wire _16372_;
 wire _16373_;
 wire _16374_;
 wire _16375_;
 wire _16376_;
 wire _16377_;
 wire _16378_;
 wire _16379_;
 wire _16380_;
 wire _16381_;
 wire _16382_;
 wire _16383_;
 wire _16384_;
 wire _16385_;
 wire _16386_;
 wire _16387_;
 wire _16388_;
 wire _16389_;
 wire _16390_;
 wire _16391_;
 wire _16392_;
 wire _16393_;
 wire _16394_;
 wire _16395_;
 wire _16396_;
 wire _16397_;
 wire _16398_;
 wire _16399_;
 wire _16400_;
 wire _16401_;
 wire _16402_;
 wire _16403_;
 wire _16404_;
 wire _16405_;
 wire _16406_;
 wire _16407_;
 wire _16408_;
 wire _16409_;
 wire _16410_;
 wire _16411_;
 wire _16412_;
 wire _16413_;
 wire _16414_;
 wire _16415_;
 wire _16416_;
 wire _16417_;
 wire _16418_;
 wire _16419_;
 wire _16420_;
 wire _16421_;
 wire _16422_;
 wire _16423_;
 wire _16424_;
 wire _16425_;
 wire _16426_;
 wire _16427_;
 wire _16428_;
 wire _16429_;
 wire _16430_;
 wire _16431_;
 wire _16432_;
 wire _16433_;
 wire _16434_;
 wire _16435_;
 wire _16436_;
 wire _16437_;
 wire _16438_;
 wire _16439_;
 wire _16440_;
 wire _16441_;
 wire _16442_;
 wire _16443_;
 wire _16444_;
 wire _16445_;
 wire _16446_;
 wire _16447_;
 wire _16448_;
 wire _16449_;
 wire _16450_;
 wire _16451_;
 wire _16452_;
 wire _16453_;
 wire _16454_;
 wire _16455_;
 wire _16456_;
 wire _16457_;
 wire _16458_;
 wire _16459_;
 wire _16460_;
 wire _16461_;
 wire _16462_;
 wire _16463_;
 wire _16464_;
 wire _16465_;
 wire _16466_;
 wire _16467_;
 wire _16468_;
 wire _16469_;
 wire _16470_;
 wire _16471_;
 wire _16472_;
 wire _16473_;
 wire _16474_;
 wire _16475_;
 wire _16476_;
 wire _16477_;
 wire _16478_;
 wire _16479_;
 wire _16480_;
 wire _16481_;
 wire _16482_;
 wire _16483_;
 wire _16484_;
 wire _16485_;
 wire _16486_;
 wire _16487_;
 wire _16488_;
 wire _16489_;
 wire _16490_;
 wire _16491_;
 wire _16492_;
 wire _16493_;
 wire _16494_;
 wire _16495_;
 wire _16496_;
 wire _16497_;
 wire _16498_;
 wire _16499_;
 wire _16500_;
 wire _16501_;
 wire _16502_;
 wire _16503_;
 wire _16504_;
 wire _16505_;
 wire _16506_;
 wire _16507_;
 wire _16508_;
 wire _16509_;
 wire _16510_;
 wire _16511_;
 wire _16512_;
 wire _16513_;
 wire _16514_;
 wire _16515_;
 wire _16516_;
 wire _16517_;
 wire _16518_;
 wire _16519_;
 wire _16520_;
 wire _16521_;
 wire _16522_;
 wire _16523_;
 wire _16524_;
 wire _16525_;
 wire _16526_;
 wire _16527_;
 wire _16528_;
 wire _16529_;
 wire _16530_;
 wire _16531_;
 wire _16532_;
 wire _16533_;
 wire _16534_;
 wire _16535_;
 wire _16536_;
 wire _16537_;
 wire _16538_;
 wire _16539_;
 wire _16540_;
 wire _16541_;
 wire _16542_;
 wire _16543_;
 wire _16544_;
 wire _16545_;
 wire _16546_;
 wire _16547_;
 wire _16548_;
 wire _16549_;
 wire _16550_;
 wire _16551_;
 wire _16552_;
 wire _16553_;
 wire _16554_;
 wire _16555_;
 wire _16556_;
 wire _16557_;
 wire _16558_;
 wire _16559_;
 wire _16560_;
 wire _16561_;
 wire _16562_;
 wire _16563_;
 wire _16564_;
 wire _16565_;
 wire _16566_;
 wire _16567_;
 wire _16568_;
 wire _16569_;
 wire _16570_;
 wire _16571_;
 wire _16572_;
 wire _16573_;
 wire _16574_;
 wire _16575_;
 wire _16576_;
 wire _16577_;
 wire _16578_;
 wire _16579_;
 wire _16580_;
 wire _16581_;
 wire _16582_;
 wire _16583_;
 wire _16584_;
 wire _16585_;
 wire _16586_;
 wire _16587_;
 wire _16588_;
 wire _16589_;
 wire _16590_;
 wire _16591_;
 wire _16592_;
 wire _16593_;
 wire _16594_;
 wire _16595_;
 wire _16596_;
 wire _16597_;
 wire _16598_;
 wire _16599_;
 wire _16600_;
 wire _16601_;
 wire _16602_;
 wire _16603_;
 wire _16604_;
 wire _16605_;
 wire _16606_;
 wire _16607_;
 wire _16608_;
 wire _16609_;
 wire _16610_;
 wire _16611_;
 wire _16612_;
 wire _16613_;
 wire _16614_;
 wire _16615_;
 wire _16616_;
 wire _16617_;
 wire _16618_;
 wire _16619_;
 wire _16620_;
 wire _16621_;
 wire _16622_;
 wire _16623_;
 wire _16624_;
 wire _16625_;
 wire _16626_;
 wire _16627_;
 wire _16628_;
 wire _16629_;
 wire _16630_;
 wire _16631_;
 wire _16632_;
 wire _16633_;
 wire _16634_;
 wire _16635_;
 wire _16636_;
 wire _16637_;
 wire _16638_;
 wire _16639_;
 wire _16640_;
 wire _16641_;
 wire _16642_;
 wire _16643_;
 wire _16644_;
 wire _16645_;
 wire _16646_;
 wire _16647_;
 wire _16648_;
 wire _16649_;
 wire _16650_;
 wire _16651_;
 wire _16652_;
 wire _16653_;
 wire _16654_;
 wire _16655_;
 wire _16656_;
 wire _16657_;
 wire _16658_;
 wire _16659_;
 wire _16660_;
 wire _16661_;
 wire _16662_;
 wire _16663_;
 wire _16664_;
 wire _16665_;
 wire _16666_;
 wire _16667_;
 wire _16668_;
 wire _16669_;
 wire _16670_;
 wire _16671_;
 wire _16672_;
 wire _16673_;
 wire _16674_;
 wire _16675_;
 wire _16676_;
 wire _16677_;
 wire _16678_;
 wire _16679_;
 wire _16680_;
 wire _16681_;
 wire _16682_;
 wire _16683_;
 wire _16684_;
 wire _16685_;
 wire _16686_;
 wire _16687_;
 wire _16688_;
 wire _16689_;
 wire _16690_;
 wire _16691_;
 wire _16692_;
 wire _16693_;
 wire _16694_;
 wire _16695_;
 wire _16696_;
 wire _16697_;
 wire _16698_;
 wire _16699_;
 wire _16700_;
 wire _16701_;
 wire _16702_;
 wire _16703_;
 wire _16704_;
 wire _16705_;
 wire _16706_;
 wire _16707_;
 wire _16708_;
 wire _16709_;
 wire _16710_;
 wire _16711_;
 wire _16712_;
 wire _16713_;
 wire _16714_;
 wire _16715_;
 wire _16716_;
 wire _16717_;
 wire _16718_;
 wire _16719_;
 wire _16720_;
 wire _16721_;
 wire _16722_;
 wire _16723_;
 wire _16724_;
 wire _16725_;
 wire _16726_;
 wire _16727_;
 wire _16728_;
 wire _16729_;
 wire _16730_;
 wire _16731_;
 wire _16732_;
 wire _16733_;
 wire _16734_;
 wire _16735_;
 wire _16736_;
 wire _16737_;
 wire _16738_;
 wire _16739_;
 wire _16740_;
 wire _16741_;
 wire _16742_;
 wire _16743_;
 wire _16744_;
 wire _16745_;
 wire _16746_;
 wire _16747_;
 wire _16748_;
 wire _16749_;
 wire _16750_;
 wire _16751_;
 wire _16752_;
 wire _16753_;
 wire _16754_;
 wire _16755_;
 wire _16756_;
 wire _16757_;
 wire _16758_;
 wire _16759_;
 wire _16760_;
 wire _16761_;
 wire _16762_;
 wire _16763_;
 wire _16764_;
 wire _16765_;
 wire _16766_;
 wire _16767_;
 wire _16768_;
 wire _16769_;
 wire _16770_;
 wire _16771_;
 wire _16772_;
 wire _16773_;
 wire _16774_;
 wire _16775_;
 wire _16776_;
 wire _16777_;
 wire _16778_;
 wire _16779_;
 wire _16780_;
 wire _16781_;
 wire _16782_;
 wire _16783_;
 wire _16784_;
 wire _16785_;
 wire _16786_;
 wire _16787_;
 wire _16788_;
 wire _16789_;
 wire _16790_;
 wire _16791_;
 wire _16792_;
 wire _16793_;
 wire _16794_;
 wire _16795_;
 wire _16796_;
 wire _16797_;
 wire _16798_;
 wire _16799_;
 wire _16800_;
 wire _16801_;
 wire _16802_;
 wire _16803_;
 wire _16804_;
 wire _16805_;
 wire _16806_;
 wire _16807_;
 wire _16808_;
 wire _16809_;
 wire _16810_;
 wire _16811_;
 wire _16812_;
 wire _16813_;
 wire _16814_;
 wire _16815_;
 wire _16816_;
 wire _16817_;
 wire _16818_;
 wire _16819_;
 wire _16820_;
 wire _16821_;
 wire _16822_;
 wire _16823_;
 wire _16824_;
 wire _16825_;
 wire _16826_;
 wire _16827_;
 wire _16828_;
 wire _16829_;
 wire _16830_;
 wire _16831_;
 wire _16832_;
 wire _16833_;
 wire _16834_;
 wire _16835_;
 wire _16836_;
 wire _16837_;
 wire _16838_;
 wire _16839_;
 wire _16840_;
 wire _16841_;
 wire _16842_;
 wire _16843_;
 wire _16844_;
 wire _16845_;
 wire _16846_;
 wire _16847_;
 wire _16848_;
 wire _16849_;
 wire _16850_;
 wire _16851_;
 wire _16852_;
 wire _16853_;
 wire _16854_;
 wire _16855_;
 wire _16856_;
 wire _16857_;
 wire _16858_;
 wire _16859_;
 wire _16860_;
 wire _16861_;
 wire _16862_;
 wire _16863_;
 wire _16864_;
 wire _16865_;
 wire _16866_;
 wire _16867_;
 wire _16868_;
 wire _16869_;
 wire _16870_;
 wire _16871_;
 wire _16872_;
 wire _16873_;
 wire _16874_;
 wire _16875_;
 wire _16876_;
 wire _16877_;
 wire _16878_;
 wire _16879_;
 wire _16880_;
 wire _16881_;
 wire _16882_;
 wire _16883_;
 wire _16884_;
 wire _16885_;
 wire _16886_;
 wire _16887_;
 wire _16888_;
 wire _16889_;
 wire _16890_;
 wire _16891_;
 wire _16892_;
 wire _16893_;
 wire _16894_;
 wire _16895_;
 wire _16896_;
 wire _16897_;
 wire _16898_;
 wire _16899_;
 wire _16900_;
 wire _16901_;
 wire _16902_;
 wire _16903_;
 wire _16904_;
 wire _16905_;
 wire _16906_;
 wire _16907_;
 wire _16908_;
 wire _16909_;
 wire _16910_;
 wire _16911_;
 wire _16912_;
 wire _16913_;
 wire _16914_;
 wire _16915_;
 wire _16916_;
 wire _16917_;
 wire _16918_;
 wire _16919_;
 wire _16920_;
 wire _16921_;
 wire _16922_;
 wire _16923_;
 wire _16924_;
 wire _16925_;
 wire _16926_;
 wire _16927_;
 wire _16928_;
 wire _16929_;
 wire _16930_;
 wire _16931_;
 wire _16932_;
 wire _16933_;
 wire _16934_;
 wire _16935_;
 wire _16936_;
 wire _16937_;
 wire _16938_;
 wire _16939_;
 wire _16940_;
 wire _16941_;
 wire _16942_;
 wire _16943_;
 wire _16944_;
 wire _16945_;
 wire _16946_;
 wire _16947_;
 wire _16948_;
 wire _16949_;
 wire _16950_;
 wire _16951_;
 wire _16952_;
 wire _16953_;
 wire _16954_;
 wire _16955_;
 wire _16956_;
 wire _16957_;
 wire _16958_;
 wire _16959_;
 wire _16960_;
 wire _16961_;
 wire _16962_;
 wire _16963_;
 wire _16964_;
 wire _16965_;
 wire _16966_;
 wire _16967_;
 wire _16968_;
 wire _16969_;
 wire _16970_;
 wire _16971_;
 wire _16972_;
 wire _16973_;
 wire _16974_;
 wire _16975_;
 wire _16976_;
 wire _16977_;
 wire _16978_;
 wire _16979_;
 wire _16980_;
 wire _16981_;
 wire _16982_;
 wire _16983_;
 wire _16984_;
 wire _16985_;
 wire _16986_;
 wire _16987_;
 wire _16988_;
 wire _16989_;
 wire _16990_;
 wire _16991_;
 wire _16992_;
 wire _16993_;
 wire _16994_;
 wire _16995_;
 wire _16996_;
 wire _16997_;
 wire _16998_;
 wire _16999_;
 wire _17000_;
 wire _17001_;
 wire _17002_;
 wire _17003_;
 wire _17004_;
 wire _17005_;
 wire _17006_;
 wire _17007_;
 wire _17008_;
 wire _17009_;
 wire _17010_;
 wire _17011_;
 wire _17012_;
 wire _17013_;
 wire _17014_;
 wire _17015_;
 wire _17016_;
 wire _17017_;
 wire _17018_;
 wire _17019_;
 wire _17020_;
 wire _17021_;
 wire _17022_;
 wire _17023_;
 wire _17024_;
 wire _17025_;
 wire _17026_;
 wire _17027_;
 wire _17028_;
 wire _17029_;
 wire _17030_;
 wire _17031_;
 wire _17032_;
 wire _17033_;
 wire _17034_;
 wire _17035_;
 wire _17036_;
 wire _17037_;
 wire _17038_;
 wire _17039_;
 wire _17040_;
 wire _17041_;
 wire _17042_;
 wire _17043_;
 wire _17044_;
 wire _17045_;
 wire _17046_;
 wire _17047_;
 wire _17048_;
 wire _17049_;
 wire _17050_;
 wire _17051_;
 wire _17052_;
 wire _17053_;
 wire _17054_;
 wire _17055_;
 wire _17056_;
 wire _17057_;
 wire _17058_;
 wire _17059_;
 wire _17060_;
 wire _17061_;
 wire _17062_;
 wire _17063_;
 wire _17064_;
 wire _17065_;
 wire _17066_;
 wire _17067_;
 wire _17068_;
 wire _17069_;
 wire _17070_;
 wire _17071_;
 wire _17072_;
 wire _17073_;
 wire _17074_;
 wire _17075_;
 wire _17076_;
 wire _17077_;
 wire _17078_;
 wire _17079_;
 wire _17080_;
 wire _17081_;
 wire _17082_;
 wire _17083_;
 wire _17084_;
 wire _17085_;
 wire _17086_;
 wire _17087_;
 wire _17088_;
 wire _17089_;
 wire _17090_;
 wire _17091_;
 wire _17092_;
 wire _17093_;
 wire _17094_;
 wire _17095_;
 wire _17096_;
 wire _17097_;
 wire _17098_;
 wire _17099_;
 wire _17100_;
 wire _17101_;
 wire _17102_;
 wire _17103_;
 wire _17104_;
 wire _17105_;
 wire _17106_;
 wire _17107_;
 wire _17108_;
 wire _17109_;
 wire _17110_;
 wire _17111_;
 wire _17112_;
 wire _17113_;
 wire _17114_;
 wire _17115_;
 wire _17116_;
 wire _17117_;
 wire _17118_;
 wire _17119_;
 wire _17120_;
 wire _17121_;
 wire _17122_;
 wire _17123_;
 wire _17124_;
 wire _17125_;
 wire _17126_;
 wire _17127_;
 wire _17128_;
 wire _17129_;
 wire _17130_;
 wire _17131_;
 wire _17132_;
 wire _17133_;
 wire _17134_;
 wire _17135_;
 wire _17136_;
 wire _17137_;
 wire _17138_;
 wire _17139_;
 wire _17140_;
 wire _17141_;
 wire _17142_;
 wire _17143_;
 wire _17144_;
 wire _17145_;
 wire _17146_;
 wire _17147_;
 wire _17148_;
 wire _17149_;
 wire _17150_;
 wire _17151_;
 wire _17152_;
 wire _17153_;
 wire _17154_;
 wire _17155_;
 wire _17156_;
 wire _17157_;
 wire _17158_;
 wire _17159_;
 wire _17160_;
 wire _17161_;
 wire _17162_;
 wire _17163_;
 wire _17164_;
 wire _17165_;
 wire _17166_;
 wire _17167_;
 wire _17168_;
 wire _17169_;
 wire _17170_;
 wire _17171_;
 wire _17172_;
 wire _17173_;
 wire _17174_;
 wire _17175_;
 wire _17176_;
 wire _17177_;
 wire _17178_;
 wire _17179_;
 wire _17180_;
 wire _17181_;
 wire _17182_;
 wire _17183_;
 wire _17184_;
 wire _17185_;
 wire _17186_;
 wire _17187_;
 wire _17188_;
 wire _17189_;
 wire _17190_;
 wire _17191_;
 wire _17192_;
 wire _17193_;
 wire _17194_;
 wire _17195_;
 wire _17196_;
 wire _17197_;
 wire _17198_;
 wire _17199_;
 wire _17200_;
 wire _17201_;
 wire _17202_;
 wire _17203_;
 wire _17204_;
 wire _17205_;
 wire _17206_;
 wire _17207_;
 wire _17208_;
 wire _17209_;
 wire _17210_;
 wire _17211_;
 wire _17212_;
 wire _17213_;
 wire _17214_;
 wire _17215_;
 wire _17216_;
 wire _17217_;
 wire _17218_;
 wire _17219_;
 wire _17220_;
 wire _17221_;
 wire _17222_;
 wire _17223_;
 wire _17224_;
 wire _17225_;
 wire _17226_;
 wire _17227_;
 wire _17228_;
 wire _17229_;
 wire _17230_;
 wire _17231_;
 wire _17232_;
 wire _17233_;
 wire _17234_;
 wire _17235_;
 wire _17236_;
 wire _17237_;
 wire _17238_;
 wire _17239_;
 wire _17240_;
 wire _17241_;
 wire _17242_;
 wire _17243_;
 wire _17244_;
 wire _17245_;
 wire _17246_;
 wire _17247_;
 wire _17248_;
 wire _17249_;
 wire _17250_;
 wire _17251_;
 wire _17252_;
 wire _17253_;
 wire _17254_;
 wire _17255_;
 wire _17256_;
 wire _17257_;
 wire _17258_;
 wire _17259_;
 wire _17260_;
 wire _17261_;
 wire _17262_;
 wire _17263_;
 wire _17264_;
 wire _17265_;
 wire _17266_;
 wire _17267_;
 wire _17268_;
 wire _17269_;
 wire _17270_;
 wire _17271_;
 wire _17272_;
 wire _17273_;
 wire _17274_;
 wire _17275_;
 wire _17276_;
 wire _17277_;
 wire _17278_;
 wire _17279_;
 wire _17280_;
 wire _17281_;
 wire _17282_;
 wire _17283_;
 wire _17284_;
 wire _17285_;
 wire _17286_;
 wire _17287_;
 wire _17288_;
 wire _17289_;
 wire _17290_;
 wire _17291_;
 wire _17292_;
 wire _17293_;
 wire _17294_;
 wire _17295_;
 wire _17296_;
 wire _17297_;
 wire _17298_;
 wire _17299_;
 wire _17300_;
 wire _17301_;
 wire _17302_;
 wire _17303_;
 wire _17304_;
 wire _17305_;
 wire _17306_;
 wire _17307_;
 wire _17308_;
 wire _17309_;
 wire _17310_;
 wire _17311_;
 wire _17312_;
 wire _17313_;
 wire _17314_;
 wire _17315_;
 wire _17316_;
 wire _17317_;
 wire _17318_;
 wire _17319_;
 wire _17320_;
 wire _17321_;
 wire _17322_;
 wire _17323_;
 wire _17324_;
 wire _17325_;
 wire _17326_;
 wire _17327_;
 wire _17328_;
 wire _17329_;
 wire _17330_;
 wire _17331_;
 wire _17332_;
 wire _17333_;
 wire _17334_;
 wire _17335_;
 wire _17336_;
 wire _17337_;
 wire _17338_;
 wire _17339_;
 wire _17340_;
 wire _17341_;
 wire _17342_;
 wire _17343_;
 wire _17344_;
 wire _17345_;
 wire _17346_;
 wire _17347_;
 wire _17348_;
 wire _17349_;
 wire _17350_;
 wire _17351_;
 wire _17352_;
 wire _17353_;
 wire _17354_;
 wire _17355_;
 wire _17356_;
 wire _17357_;
 wire _17358_;
 wire _17359_;
 wire _17360_;
 wire _17361_;
 wire _17362_;
 wire _17363_;
 wire _17364_;
 wire _17365_;
 wire _17366_;
 wire _17367_;
 wire _17368_;
 wire _17369_;
 wire _17370_;
 wire _17371_;
 wire _17372_;
 wire _17373_;
 wire _17374_;
 wire _17375_;
 wire _17376_;
 wire _17377_;
 wire _17378_;
 wire _17379_;
 wire _17380_;
 wire _17381_;
 wire _17382_;
 wire _17383_;
 wire _17384_;
 wire _17385_;
 wire _17386_;
 wire _17387_;
 wire _17388_;
 wire _17389_;
 wire _17390_;
 wire _17391_;
 wire _17392_;
 wire _17393_;
 wire _17394_;
 wire _17395_;
 wire _17396_;
 wire _17397_;
 wire _17398_;
 wire _17399_;
 wire _17400_;
 wire _17401_;
 wire _17402_;
 wire _17403_;
 wire _17404_;
 wire _17405_;
 wire _17406_;
 wire _17407_;
 wire _17408_;
 wire _17409_;
 wire _17410_;
 wire _17411_;
 wire _17412_;
 wire _17413_;
 wire _17414_;
 wire _17415_;
 wire _17416_;
 wire _17417_;
 wire _17418_;
 wire _17419_;
 wire _17420_;
 wire _17421_;
 wire _17422_;
 wire _17423_;
 wire _17424_;
 wire _17425_;
 wire _17426_;
 wire _17427_;
 wire _17428_;
 wire _17429_;
 wire _17430_;
 wire _17431_;
 wire _17432_;
 wire _17433_;
 wire _17434_;
 wire _17435_;
 wire _17436_;
 wire _17437_;
 wire _17438_;
 wire _17439_;
 wire _17440_;
 wire _17441_;
 wire _17442_;
 wire _17443_;
 wire _17444_;
 wire _17445_;
 wire _17446_;
 wire _17447_;
 wire _17448_;
 wire _17449_;
 wire _17450_;
 wire _17451_;
 wire _17452_;
 wire _17453_;
 wire _17454_;
 wire _17455_;
 wire _17456_;
 wire _17457_;
 wire _17458_;
 wire _17459_;
 wire _17460_;
 wire _17461_;
 wire _17462_;
 wire _17463_;
 wire _17464_;
 wire _17465_;
 wire _17466_;
 wire _17467_;
 wire _17468_;
 wire _17469_;
 wire _17470_;
 wire _17471_;
 wire _17472_;
 wire _17473_;
 wire _17474_;
 wire _17475_;
 wire _17476_;
 wire _17477_;
 wire _17478_;
 wire _17479_;
 wire _17480_;
 wire _17481_;
 wire _17482_;
 wire _17483_;
 wire _17484_;
 wire _17485_;
 wire _17486_;
 wire _17487_;
 wire _17488_;
 wire _17489_;
 wire _17490_;
 wire _17491_;
 wire _17492_;
 wire _17493_;
 wire _17494_;
 wire _17495_;
 wire _17496_;
 wire _17497_;
 wire _17498_;
 wire _17499_;
 wire _17500_;
 wire _17501_;
 wire _17502_;
 wire _17503_;
 wire _17504_;
 wire _17505_;
 wire _17506_;
 wire _17507_;
 wire _17508_;
 wire _17509_;
 wire _17510_;
 wire _17511_;
 wire _17512_;
 wire _17513_;
 wire _17514_;
 wire _17515_;
 wire _17516_;
 wire _17517_;
 wire _17518_;
 wire _17519_;
 wire _17520_;
 wire _17521_;
 wire _17522_;
 wire _17523_;
 wire _17524_;
 wire _17525_;
 wire _17526_;
 wire _17527_;
 wire _17528_;
 wire _17529_;
 wire _17530_;
 wire _17531_;
 wire _17532_;
 wire _17533_;
 wire _17534_;
 wire _17535_;
 wire _17536_;
 wire _17537_;
 wire _17538_;
 wire _17539_;
 wire _17540_;
 wire _17541_;
 wire _17542_;
 wire _17543_;
 wire _17544_;
 wire _17545_;
 wire _17546_;
 wire _17547_;
 wire _17548_;
 wire _17549_;
 wire _17550_;
 wire _17551_;
 wire _17552_;
 wire _17553_;
 wire _17554_;
 wire _17555_;
 wire _17556_;
 wire _17557_;
 wire _17558_;
 wire _17559_;
 wire _17560_;
 wire _17561_;
 wire _17562_;
 wire _17563_;
 wire _17564_;
 wire _17565_;
 wire _17566_;
 wire _17567_;
 wire _17568_;
 wire _17569_;
 wire _17570_;
 wire _17571_;
 wire _17572_;
 wire _17573_;
 wire _17574_;
 wire _17575_;
 wire _17576_;
 wire _17577_;
 wire _17578_;
 wire _17579_;
 wire _17580_;
 wire _17581_;
 wire _17582_;
 wire _17583_;
 wire _17584_;
 wire _17585_;
 wire _17586_;
 wire _17587_;
 wire _17588_;
 wire _17589_;
 wire _17590_;
 wire _17591_;
 wire _17592_;
 wire _17593_;
 wire _17594_;
 wire _17595_;
 wire _17596_;
 wire _17597_;
 wire _17598_;
 wire _17599_;
 wire _17600_;
 wire _17601_;
 wire _17602_;
 wire _17603_;
 wire _17604_;
 wire _17605_;
 wire _17606_;
 wire _17607_;
 wire _17608_;
 wire _17609_;
 wire _17610_;
 wire _17611_;
 wire _17612_;
 wire _17613_;
 wire _17614_;
 wire _17615_;
 wire _17616_;
 wire _17617_;
 wire _17618_;
 wire _17619_;
 wire _17620_;
 wire _17621_;
 wire _17622_;
 wire _17623_;
 wire _17624_;
 wire _17625_;
 wire _17626_;
 wire _17627_;
 wire _17628_;
 wire _17629_;
 wire _17630_;
 wire _17631_;
 wire _17632_;
 wire _17633_;
 wire _17634_;
 wire _17635_;
 wire _17636_;
 wire _17637_;
 wire _17638_;
 wire _17639_;
 wire _17640_;
 wire _17641_;
 wire _17642_;
 wire _17643_;
 wire _17644_;
 wire _17645_;
 wire _17646_;
 wire _17647_;
 wire _17648_;
 wire _17649_;
 wire _17650_;
 wire _17651_;
 wire _17652_;
 wire _17653_;
 wire _17654_;
 wire _17655_;
 wire _17656_;
 wire _17657_;
 wire _17658_;
 wire _17659_;
 wire _17660_;
 wire _17661_;
 wire _17662_;
 wire _17663_;
 wire _17664_;
 wire _17665_;
 wire _17666_;
 wire _17667_;
 wire _17668_;
 wire _17669_;
 wire _17670_;
 wire _17671_;
 wire _17672_;
 wire _17673_;
 wire _17674_;
 wire _17675_;
 wire _17676_;
 wire _17677_;
 wire _17678_;
 wire _17679_;
 wire _17680_;
 wire _17681_;
 wire _17682_;
 wire _17683_;
 wire _17684_;
 wire _17685_;
 wire _17686_;
 wire _17687_;
 wire _17688_;
 wire _17689_;
 wire _17690_;
 wire _17691_;
 wire _17692_;
 wire _17693_;
 wire _17694_;
 wire _17695_;
 wire _17696_;
 wire _17697_;
 wire _17698_;
 wire _17699_;
 wire _17700_;
 wire _17701_;
 wire _17702_;
 wire _17703_;
 wire _17704_;
 wire _17705_;
 wire _17706_;
 wire _17707_;
 wire _17708_;
 wire _17709_;
 wire _17710_;
 wire _17711_;
 wire _17712_;
 wire _17713_;
 wire _17714_;
 wire _17715_;
 wire _17716_;
 wire _17717_;
 wire _17718_;
 wire _17719_;
 wire _17720_;
 wire _17721_;
 wire _17722_;
 wire _17723_;
 wire _17724_;
 wire _17725_;
 wire _17726_;
 wire _17727_;
 wire _17728_;
 wire _17729_;
 wire _17730_;
 wire _17731_;
 wire _17732_;
 wire _17733_;
 wire _17734_;
 wire _17735_;
 wire _17736_;
 wire _17737_;
 wire _17738_;
 wire _17739_;
 wire _17740_;
 wire _17741_;
 wire _17742_;
 wire _17743_;
 wire _17744_;
 wire _17745_;
 wire _17746_;
 wire _17747_;
 wire _17748_;
 wire _17749_;
 wire _17750_;
 wire _17751_;
 wire _17752_;
 wire _17753_;
 wire _17754_;
 wire _17755_;
 wire _17756_;
 wire _17757_;
 wire _17758_;
 wire _17759_;
 wire _17760_;
 wire _17761_;
 wire _17762_;
 wire _17763_;
 wire _17764_;
 wire _17765_;
 wire _17766_;
 wire _17767_;
 wire _17768_;
 wire _17769_;
 wire _17770_;
 wire _17771_;
 wire _17772_;
 wire _17773_;
 wire _17774_;
 wire _17775_;
 wire _17776_;
 wire _17777_;
 wire _17778_;
 wire _17779_;
 wire _17780_;
 wire _17781_;
 wire _17782_;
 wire _17783_;
 wire _17784_;
 wire _17785_;
 wire _17786_;
 wire _17787_;
 wire _17788_;
 wire _17789_;
 wire _17790_;
 wire _17791_;
 wire _17792_;
 wire _17793_;
 wire _17794_;
 wire _17795_;
 wire _17796_;
 wire _17797_;
 wire _17798_;
 wire _17799_;
 wire _17800_;
 wire _17801_;
 wire _17802_;
 wire _17803_;
 wire _17804_;
 wire _17805_;
 wire _17806_;
 wire _17807_;
 wire _17808_;
 wire _17809_;
 wire _17810_;
 wire _17811_;
 wire _17812_;
 wire _17813_;
 wire _17814_;
 wire _17815_;
 wire _17816_;
 wire _17817_;
 wire _17818_;
 wire _17819_;
 wire _17820_;
 wire _17821_;
 wire _17822_;
 wire _17823_;
 wire _17824_;
 wire _17825_;
 wire _17826_;
 wire _17827_;
 wire _17828_;
 wire _17829_;
 wire _17830_;
 wire _17831_;
 wire _17832_;
 wire _17833_;
 wire _17834_;
 wire _17835_;
 wire _17836_;
 wire _17837_;
 wire _17838_;
 wire _17839_;
 wire _17840_;
 wire _17841_;
 wire _17842_;
 wire _17843_;
 wire _17844_;
 wire _17845_;
 wire _17846_;
 wire _17847_;
 wire _17848_;
 wire _17849_;
 wire _17850_;
 wire _17851_;
 wire _17852_;
 wire _17853_;
 wire _17854_;
 wire _17855_;
 wire _17856_;
 wire _17857_;
 wire _17858_;
 wire _17859_;
 wire _17860_;
 wire _17861_;
 wire _17862_;
 wire _17863_;
 wire _17864_;
 wire _17865_;
 wire _17866_;
 wire _17867_;
 wire _17868_;
 wire _17869_;
 wire _17870_;
 wire _17871_;
 wire _17872_;
 wire _17873_;
 wire _17874_;
 wire _17875_;
 wire _17876_;
 wire _17877_;
 wire _17878_;
 wire _17879_;
 wire _17880_;
 wire _17881_;
 wire _17882_;
 wire _17883_;
 wire _17884_;
 wire _17885_;
 wire _17886_;
 wire _17887_;
 wire _17888_;
 wire _17889_;
 wire _17890_;
 wire _17891_;
 wire _17892_;
 wire _17893_;
 wire _17894_;
 wire _17895_;
 wire _17896_;
 wire _17897_;
 wire _17898_;
 wire _17899_;
 wire _17900_;
 wire _17901_;
 wire _17902_;
 wire _17903_;
 wire _17904_;
 wire _17905_;
 wire _17906_;
 wire _17907_;
 wire _17908_;
 wire _17909_;
 wire _17910_;
 wire _17911_;
 wire _17912_;
 wire _17913_;
 wire _17914_;
 wire _17915_;
 wire _17916_;
 wire _17917_;
 wire _17918_;
 wire _17919_;
 wire _17920_;
 wire _17921_;
 wire _17922_;
 wire _17923_;
 wire _17924_;
 wire _17925_;
 wire _17926_;
 wire _17927_;
 wire _17928_;
 wire _17929_;
 wire _17930_;
 wire _17931_;
 wire _17932_;
 wire _17933_;
 wire _17934_;
 wire _17935_;
 wire _17936_;
 wire _17937_;
 wire _17938_;
 wire _17939_;
 wire _17940_;
 wire _17941_;
 wire _17942_;
 wire _17943_;
 wire _17944_;
 wire _17945_;
 wire _17946_;
 wire _17947_;
 wire _17948_;
 wire _17949_;
 wire _17950_;
 wire _17951_;
 wire _17952_;
 wire _17953_;
 wire _17954_;
 wire _17955_;
 wire _17956_;
 wire _17957_;
 wire _17958_;
 wire _17959_;
 wire _17960_;
 wire _17961_;
 wire _17962_;
 wire _17963_;
 wire _17964_;
 wire _17965_;
 wire _17966_;
 wire _17967_;
 wire _17968_;
 wire _17969_;
 wire _17970_;
 wire _17971_;
 wire _17972_;
 wire _17973_;
 wire _17974_;
 wire _17975_;
 wire _17976_;
 wire _17977_;
 wire _17978_;
 wire _17979_;
 wire _17980_;
 wire _17981_;
 wire _17982_;
 wire _17983_;
 wire _17984_;
 wire _17985_;
 wire _17986_;
 wire _17987_;
 wire _17988_;
 wire _17989_;
 wire _17990_;
 wire _17991_;
 wire _17992_;
 wire _17993_;
 wire _17994_;
 wire _17995_;
 wire _17996_;
 wire _17997_;
 wire _17998_;
 wire _17999_;
 wire _18000_;
 wire _18001_;
 wire _18002_;
 wire _18003_;
 wire _18004_;
 wire _18005_;
 wire _18006_;
 wire _18007_;
 wire _18008_;
 wire _18009_;
 wire _18010_;
 wire _18011_;
 wire _18012_;
 wire _18013_;
 wire _18014_;
 wire _18015_;
 wire _18016_;
 wire _18017_;
 wire _18018_;
 wire _18019_;
 wire _18020_;
 wire _18021_;
 wire _18022_;
 wire _18023_;
 wire _18024_;
 wire _18025_;
 wire _18026_;
 wire _18027_;
 wire _18028_;
 wire _18029_;
 wire _18030_;
 wire _18031_;
 wire _18032_;
 wire _18033_;
 wire _18034_;
 wire _18035_;
 wire _18036_;
 wire _18037_;
 wire _18038_;
 wire _18039_;
 wire _18040_;
 wire _18041_;
 wire _18042_;
 wire _18043_;
 wire _18044_;
 wire _18045_;
 wire _18046_;
 wire _18047_;
 wire _18048_;
 wire _18049_;
 wire _18050_;
 wire _18051_;
 wire _18052_;
 wire _18053_;
 wire _18054_;
 wire _18055_;
 wire _18056_;
 wire _18057_;
 wire _18058_;
 wire _18059_;
 wire _18060_;
 wire _18061_;
 wire _18062_;
 wire _18063_;
 wire _18064_;
 wire _18065_;
 wire _18066_;
 wire _18067_;
 wire _18068_;
 wire _18069_;
 wire _18070_;
 wire _18071_;
 wire _18072_;
 wire _18073_;
 wire _18074_;
 wire _18075_;
 wire _18076_;
 wire _18077_;
 wire _18078_;
 wire _18079_;
 wire _18080_;
 wire _18081_;
 wire _18082_;
 wire _18083_;
 wire _18084_;
 wire _18085_;
 wire _18086_;
 wire _18087_;
 wire _18088_;
 wire _18089_;
 wire _18090_;
 wire _18091_;
 wire _18092_;
 wire _18093_;
 wire _18094_;
 wire _18095_;
 wire _18096_;
 wire _18097_;
 wire _18098_;
 wire _18099_;
 wire _18100_;
 wire _18101_;
 wire _18102_;
 wire _18103_;
 wire _18104_;
 wire _18105_;
 wire _18106_;
 wire _18107_;
 wire _18108_;
 wire _18109_;
 wire _18110_;
 wire _18111_;
 wire _18112_;
 wire _18113_;
 wire _18114_;
 wire _18115_;
 wire _18116_;
 wire _18117_;
 wire _18118_;
 wire _18119_;
 wire _18120_;
 wire _18121_;
 wire _18122_;
 wire _18123_;
 wire _18124_;
 wire _18125_;
 wire _18126_;
 wire _18127_;
 wire _18128_;
 wire _18129_;
 wire _18130_;
 wire _18131_;
 wire _18132_;
 wire _18133_;
 wire _18134_;
 wire _18135_;
 wire _18136_;
 wire _18137_;
 wire _18138_;
 wire _18139_;
 wire _18140_;
 wire _18141_;
 wire _18142_;
 wire _18143_;
 wire _18144_;
 wire _18145_;
 wire _18146_;
 wire _18147_;
 wire _18148_;
 wire _18149_;
 wire _18150_;
 wire _18151_;
 wire _18152_;
 wire _18153_;
 wire _18154_;
 wire _18155_;
 wire _18156_;
 wire _18157_;
 wire _18158_;
 wire _18159_;
 wire _18160_;
 wire _18161_;
 wire _18162_;
 wire _18163_;
 wire _18164_;
 wire _18165_;
 wire _18166_;
 wire _18167_;
 wire _18168_;
 wire _18169_;
 wire _18170_;
 wire _18171_;
 wire _18172_;
 wire _18173_;
 wire _18174_;
 wire _18175_;
 wire _18176_;
 wire _18177_;
 wire _18178_;
 wire _18179_;
 wire _18180_;
 wire _18181_;
 wire _18182_;
 wire _18183_;
 wire _18184_;
 wire _18185_;
 wire _18186_;
 wire _18187_;
 wire _18188_;
 wire _18189_;
 wire _18190_;
 wire _18191_;
 wire _18192_;
 wire _18193_;
 wire _18194_;
 wire _18195_;
 wire _18196_;
 wire _18197_;
 wire _18198_;
 wire _18199_;
 wire _18200_;
 wire _18201_;
 wire _18202_;
 wire _18203_;
 wire _18204_;
 wire _18205_;
 wire _18206_;
 wire _18207_;
 wire _18208_;
 wire _18209_;
 wire _18210_;
 wire _18211_;
 wire _18212_;
 wire _18213_;
 wire _18214_;
 wire _18215_;
 wire _18216_;
 wire _18217_;
 wire _18218_;
 wire _18219_;
 wire _18220_;
 wire _18221_;
 wire _18222_;
 wire _18223_;
 wire _18224_;
 wire _18225_;
 wire _18226_;
 wire _18227_;
 wire _18228_;
 wire _18229_;
 wire _18230_;
 wire _18231_;
 wire _18232_;
 wire _18233_;
 wire _18234_;
 wire _18235_;
 wire _18236_;
 wire _18237_;
 wire _18238_;
 wire _18239_;
 wire _18240_;
 wire _18241_;
 wire _18242_;
 wire _18243_;
 wire _18244_;
 wire _18245_;
 wire _18246_;
 wire _18247_;
 wire _18248_;
 wire _18249_;
 wire _18250_;
 wire _18251_;
 wire _18252_;
 wire _18253_;
 wire _18254_;
 wire _18255_;
 wire _18256_;
 wire _18257_;
 wire _18258_;
 wire _18259_;
 wire _18260_;
 wire _18261_;
 wire _18262_;
 wire _18263_;
 wire _18264_;
 wire _18265_;
 wire _18266_;
 wire _18267_;
 wire _18268_;
 wire _18269_;
 wire _18270_;
 wire _18271_;
 wire _18272_;
 wire _18273_;
 wire _18274_;
 wire _18275_;
 wire _18276_;
 wire _18277_;
 wire _18278_;
 wire _18279_;
 wire _18280_;
 wire _18281_;
 wire _18282_;
 wire _18283_;
 wire _18284_;
 wire _18285_;
 wire _18286_;
 wire _18287_;
 wire _18288_;
 wire _18289_;
 wire _18290_;
 wire _18291_;
 wire _18292_;
 wire _18293_;
 wire _18294_;
 wire _18295_;
 wire _18296_;
 wire _18297_;
 wire _18298_;
 wire _18299_;
 wire _18300_;
 wire _18301_;
 wire _18302_;
 wire _18303_;
 wire _18304_;
 wire _18305_;
 wire _18306_;
 wire _18307_;
 wire _18308_;
 wire _18309_;
 wire _18310_;
 wire _18311_;
 wire _18312_;
 wire _18313_;
 wire _18314_;
 wire _18315_;
 wire _18316_;
 wire _18317_;
 wire _18318_;
 wire _18319_;
 wire _18320_;
 wire _18321_;
 wire _18322_;
 wire _18323_;
 wire _18324_;
 wire _18325_;
 wire _18326_;
 wire _18327_;
 wire _18328_;
 wire _18329_;
 wire _18330_;
 wire _18331_;
 wire _18332_;
 wire _18333_;
 wire _18334_;
 wire _18335_;
 wire _18336_;
 wire _18337_;
 wire _18338_;
 wire _18339_;
 wire _18340_;
 wire _18341_;
 wire _18342_;
 wire _18343_;
 wire _18344_;
 wire _18345_;
 wire _18346_;
 wire _18347_;
 wire _18348_;
 wire _18349_;
 wire _18350_;
 wire _18351_;
 wire _18352_;
 wire _18353_;
 wire _18354_;
 wire _18355_;
 wire _18356_;
 wire _18357_;
 wire _18358_;
 wire _18359_;
 wire _18360_;
 wire _18361_;
 wire _18362_;
 wire _18363_;
 wire _18364_;
 wire _18365_;
 wire _18366_;
 wire _18367_;
 wire _18368_;
 wire _18369_;
 wire _18370_;
 wire _18371_;
 wire _18372_;
 wire _18373_;
 wire _18374_;
 wire _18375_;
 wire _18376_;
 wire _18377_;
 wire _18378_;
 wire _18379_;
 wire _18380_;
 wire _18381_;
 wire _18382_;
 wire _18383_;
 wire _18384_;
 wire _18385_;
 wire _18386_;
 wire _18387_;
 wire _18388_;
 wire _18389_;
 wire _18390_;
 wire _18391_;
 wire _18392_;
 wire _18393_;
 wire _18394_;
 wire _18395_;
 wire _18396_;
 wire _18397_;
 wire _18398_;
 wire _18399_;
 wire _18400_;
 wire _18401_;
 wire _18402_;
 wire _18403_;
 wire _18404_;
 wire _18405_;
 wire _18406_;
 wire _18407_;
 wire _18408_;
 wire _18409_;
 wire _18410_;
 wire _18411_;
 wire _18412_;
 wire _18413_;
 wire _18414_;
 wire _18415_;
 wire _18416_;
 wire _18417_;
 wire _18418_;
 wire _18419_;
 wire _18420_;
 wire _18421_;
 wire _18422_;
 wire _18423_;
 wire _18424_;
 wire _18425_;
 wire _18426_;
 wire _18427_;
 wire _18428_;
 wire _18429_;
 wire _18430_;
 wire _18431_;
 wire _18432_;
 wire _18433_;
 wire _18434_;
 wire _18435_;
 wire _18436_;
 wire _18437_;
 wire _18438_;
 wire _18439_;
 wire _18440_;
 wire _18441_;
 wire _18442_;
 wire _18443_;
 wire _18444_;
 wire _18445_;
 wire _18446_;
 wire _18447_;
 wire _18448_;
 wire _18449_;
 wire _18450_;
 wire _18451_;
 wire _18452_;
 wire _18453_;
 wire _18454_;
 wire _18455_;
 wire _18456_;
 wire _18457_;
 wire _18458_;
 wire _18459_;
 wire _18460_;
 wire _18461_;
 wire _18462_;
 wire _18463_;
 wire _18464_;
 wire _18465_;
 wire _18466_;
 wire _18467_;
 wire _18468_;
 wire _18469_;
 wire _18470_;
 wire _18471_;
 wire _18472_;
 wire _18473_;
 wire _18474_;
 wire _18475_;
 wire _18476_;
 wire _18477_;
 wire _18478_;
 wire _18479_;
 wire _18480_;
 wire _18481_;
 wire _18482_;
 wire _18483_;
 wire _18484_;
 wire _18485_;
 wire _18486_;
 wire _18487_;
 wire _18488_;
 wire _18489_;
 wire _18490_;
 wire _18491_;
 wire _18492_;
 wire _18493_;
 wire _18494_;
 wire _18495_;
 wire _18496_;
 wire _18497_;
 wire _18498_;
 wire _18499_;
 wire _18500_;
 wire _18501_;
 wire _18502_;
 wire _18503_;
 wire _18504_;
 wire _18505_;
 wire _18506_;
 wire _18507_;
 wire _18508_;
 wire _18509_;
 wire _18510_;
 wire _18511_;
 wire _18512_;
 wire _18513_;
 wire _18514_;
 wire _18515_;
 wire _18516_;
 wire _18517_;
 wire _18518_;
 wire _18519_;
 wire _18520_;
 wire _18521_;
 wire _18522_;
 wire _18523_;
 wire _18524_;
 wire _18525_;
 wire _18526_;
 wire _18527_;
 wire _18528_;
 wire _18529_;
 wire _18530_;
 wire _18531_;
 wire _18532_;
 wire _18533_;
 wire _18534_;
 wire _18535_;
 wire _18536_;
 wire _18537_;
 wire _18538_;
 wire _18539_;
 wire _18540_;
 wire _18541_;
 wire _18542_;
 wire _18543_;
 wire _18544_;
 wire _18545_;
 wire _18546_;
 wire _18547_;
 wire _18548_;
 wire _18549_;
 wire _18550_;
 wire _18551_;
 wire _18552_;
 wire _18553_;
 wire _18554_;
 wire _18555_;
 wire _18556_;
 wire _18557_;
 wire _18558_;
 wire _18559_;
 wire _18560_;
 wire _18561_;
 wire _18562_;
 wire _18563_;
 wire _18564_;
 wire _18565_;
 wire _18566_;
 wire _18567_;
 wire _18568_;
 wire _18569_;
 wire _18570_;
 wire _18571_;
 wire _18572_;
 wire _18573_;
 wire _18574_;
 wire _18575_;
 wire _18576_;
 wire _18577_;
 wire _18578_;
 wire _18579_;
 wire _18580_;
 wire _18581_;
 wire _18582_;
 wire _18583_;
 wire _18584_;
 wire _18585_;
 wire _18586_;
 wire _18587_;
 wire _18588_;
 wire _18589_;
 wire _18590_;
 wire _18591_;
 wire _18592_;
 wire _18593_;
 wire _18594_;
 wire _18595_;
 wire _18596_;
 wire _18597_;
 wire _18598_;
 wire _18599_;
 wire _18600_;
 wire _18601_;
 wire _18602_;
 wire _18603_;
 wire _18604_;
 wire _18605_;
 wire _18606_;
 wire _18607_;
 wire _18608_;
 wire _18609_;
 wire _18610_;
 wire _18611_;
 wire _18612_;
 wire _18613_;
 wire _18614_;
 wire _18615_;
 wire _18616_;
 wire _18617_;
 wire _18618_;
 wire _18619_;
 wire _18620_;
 wire _18621_;
 wire _18622_;
 wire _18623_;
 wire _18624_;
 wire _18625_;
 wire _18626_;
 wire _18627_;
 wire _18628_;
 wire _18629_;
 wire _18630_;
 wire _18631_;
 wire _18632_;
 wire _18633_;
 wire _18634_;
 wire _18635_;
 wire _18636_;
 wire _18637_;
 wire _18638_;
 wire _18639_;
 wire _18640_;
 wire _18641_;
 wire _18642_;
 wire _18643_;
 wire _18644_;
 wire _18645_;
 wire _18646_;
 wire _18647_;
 wire _18648_;
 wire _18649_;
 wire _18650_;
 wire _18651_;
 wire _18652_;
 wire _18653_;
 wire _18654_;
 wire _18655_;
 wire _18656_;
 wire _18657_;
 wire _18658_;
 wire _18659_;
 wire _18660_;
 wire _18661_;
 wire _18662_;
 wire _18663_;
 wire _18664_;
 wire _18665_;
 wire _18666_;
 wire _18667_;
 wire _18668_;
 wire _18669_;
 wire _18670_;
 wire _18671_;
 wire _18672_;
 wire _18673_;
 wire _18674_;
 wire _18675_;
 wire _18676_;
 wire _18677_;
 wire _18678_;
 wire _18679_;
 wire _18680_;
 wire _18681_;
 wire _18682_;
 wire _18683_;
 wire _18684_;
 wire _18685_;
 wire _18686_;
 wire _18687_;
 wire _18688_;
 wire _18689_;
 wire _18690_;
 wire _18691_;
 wire _18692_;
 wire _18693_;
 wire _18694_;
 wire _18695_;
 wire _18696_;
 wire _18697_;
 wire _18698_;
 wire _18699_;
 wire _18700_;
 wire _18701_;
 wire _18702_;
 wire _18703_;
 wire _18704_;
 wire _18705_;
 wire _18706_;
 wire _18707_;
 wire _18708_;
 wire _18709_;
 wire _18710_;
 wire _18711_;
 wire _18712_;
 wire _18713_;
 wire _18714_;
 wire _18715_;
 wire _18716_;
 wire _18717_;
 wire _18718_;
 wire _18719_;
 wire _18720_;
 wire _18721_;
 wire _18722_;
 wire _18723_;
 wire _18724_;
 wire _18725_;
 wire _18726_;
 wire _18727_;
 wire _18728_;
 wire _18729_;
 wire _18730_;
 wire _18731_;
 wire _18732_;
 wire _18733_;
 wire _18734_;
 wire _18735_;
 wire _18736_;
 wire _18737_;
 wire _18738_;
 wire _18739_;
 wire _18740_;
 wire _18741_;
 wire _18742_;
 wire _18743_;
 wire _18744_;
 wire _18745_;
 wire _18746_;
 wire _18747_;
 wire _18748_;
 wire _18749_;
 wire _18750_;
 wire _18751_;
 wire _18752_;
 wire _18753_;
 wire _18754_;
 wire _18755_;
 wire _18756_;
 wire _18757_;
 wire _18758_;
 wire _18759_;
 wire _18760_;
 wire _18761_;
 wire _18762_;
 wire _18763_;
 wire _18764_;
 wire _18765_;
 wire _18766_;
 wire _18767_;
 wire _18768_;
 wire _18769_;
 wire _18770_;
 wire _18771_;
 wire _18772_;
 wire _18773_;
 wire _18774_;
 wire _18775_;
 wire _18776_;
 wire _18777_;
 wire _18778_;
 wire _18779_;
 wire _18780_;
 wire _18781_;
 wire _18782_;
 wire _18783_;
 wire _18784_;
 wire _18785_;
 wire _18786_;
 wire _18787_;
 wire _18788_;
 wire _18789_;
 wire _18790_;
 wire _18791_;
 wire _18792_;
 wire _18793_;
 wire _18794_;
 wire _18795_;
 wire _18796_;
 wire _18797_;
 wire _18798_;
 wire _18799_;
 wire _18800_;
 wire _18801_;
 wire _18802_;
 wire _18803_;
 wire _18804_;
 wire _18805_;
 wire _18806_;
 wire _18807_;
 wire _18808_;
 wire _18809_;
 wire _18810_;
 wire _18811_;
 wire _18812_;
 wire _18813_;
 wire _18814_;
 wire _18815_;
 wire _18816_;
 wire _18817_;
 wire _18818_;
 wire _18819_;
 wire _18820_;
 wire _18821_;
 wire _18822_;
 wire _18823_;
 wire _18824_;
 wire _18825_;
 wire _18826_;
 wire _18827_;
 wire _18828_;
 wire _18829_;
 wire _18830_;
 wire _18831_;
 wire _18832_;
 wire _18833_;
 wire _18834_;
 wire _18835_;
 wire _18836_;
 wire _18837_;
 wire _18838_;
 wire _18839_;
 wire _18840_;
 wire _18841_;
 wire _18842_;
 wire _18843_;
 wire _18844_;
 wire _18845_;
 wire _18846_;
 wire _18847_;
 wire _18848_;
 wire _18849_;
 wire _18850_;
 wire _18851_;
 wire _18852_;
 wire _18853_;
 wire _18854_;
 wire _18855_;
 wire _18856_;
 wire _18857_;
 wire _18858_;
 wire _18859_;
 wire _18860_;
 wire _18861_;
 wire _18862_;
 wire _18863_;
 wire _18864_;
 wire _18865_;
 wire _18866_;
 wire _18867_;
 wire _18868_;
 wire _18869_;
 wire _18870_;
 wire _18871_;
 wire _18872_;
 wire _18873_;
 wire _18874_;
 wire _18875_;
 wire _18876_;
 wire _18877_;
 wire _18878_;
 wire _18879_;
 wire _18880_;
 wire _18881_;
 wire _18882_;
 wire _18883_;
 wire _18884_;
 wire _18885_;
 wire _18886_;
 wire _18887_;
 wire _18888_;
 wire _18889_;
 wire _18890_;
 wire _18891_;
 wire _18892_;
 wire _18893_;
 wire _18894_;
 wire _18895_;
 wire _18896_;
 wire _18897_;
 wire _18898_;
 wire _18899_;
 wire _18900_;
 wire _18901_;
 wire _18902_;
 wire _18903_;
 wire _18904_;
 wire _18905_;
 wire _18906_;
 wire _18907_;
 wire _18908_;
 wire _18909_;
 wire _18910_;
 wire _18911_;
 wire _18912_;
 wire _18913_;
 wire _18914_;
 wire _18915_;
 wire _18916_;
 wire _18917_;
 wire _18918_;
 wire _18919_;
 wire _18920_;
 wire _18921_;
 wire _18922_;
 wire _18923_;
 wire _18924_;
 wire _18925_;
 wire _18926_;
 wire _18927_;
 wire _18928_;
 wire _18929_;
 wire _18930_;
 wire _18931_;
 wire _18932_;
 wire _18933_;
 wire _18934_;
 wire _18935_;
 wire _18936_;
 wire _18937_;
 wire _18938_;
 wire _18939_;
 wire _18940_;
 wire _18941_;
 wire _18942_;
 wire _18943_;
 wire _18944_;
 wire _18945_;
 wire _18946_;
 wire _18947_;
 wire _18948_;
 wire _18949_;
 wire _18950_;
 wire _18951_;
 wire _18952_;
 wire _18953_;
 wire _18954_;
 wire _18955_;
 wire _18956_;
 wire _18957_;
 wire _18958_;
 wire _18959_;
 wire _18960_;
 wire _18961_;
 wire _18962_;
 wire _18963_;
 wire _18964_;
 wire _18965_;
 wire _18966_;
 wire _18967_;
 wire _18968_;
 wire _18969_;
 wire _18970_;
 wire _18971_;
 wire _18972_;
 wire _18973_;
 wire _18974_;
 wire _18975_;
 wire _18976_;
 wire _18977_;
 wire _18978_;
 wire _18979_;
 wire _18980_;
 wire _18981_;
 wire _18982_;
 wire _18983_;
 wire _18984_;
 wire _18985_;
 wire _18986_;
 wire _18987_;
 wire _18988_;
 wire _18989_;
 wire _18990_;
 wire _18991_;
 wire _18992_;
 wire _18993_;
 wire _18994_;
 wire _18995_;
 wire _18996_;
 wire _18997_;
 wire _18998_;
 wire _18999_;
 wire _19000_;
 wire _19001_;
 wire _19002_;
 wire _19003_;
 wire _19004_;
 wire _19005_;
 wire _19006_;
 wire _19007_;
 wire _19008_;
 wire _19009_;
 wire _19010_;
 wire _19011_;
 wire _19012_;
 wire _19013_;
 wire _19014_;
 wire _19015_;
 wire _19016_;
 wire _19017_;
 wire _19018_;
 wire _19019_;
 wire _19020_;
 wire _19021_;
 wire _19022_;
 wire _19023_;
 wire _19024_;
 wire _19025_;
 wire _19026_;
 wire _19027_;
 wire _19028_;
 wire _19029_;
 wire _19030_;
 wire _19031_;
 wire _19032_;
 wire _19033_;
 wire _19034_;
 wire _19035_;
 wire _19036_;
 wire _19037_;
 wire _19038_;
 wire _19039_;
 wire _19040_;
 wire _19041_;
 wire _19042_;
 wire _19043_;
 wire _19044_;
 wire _19045_;
 wire _19046_;
 wire _19047_;
 wire _19048_;
 wire _19049_;
 wire _19050_;
 wire _19051_;
 wire _19052_;
 wire _19053_;
 wire _19054_;
 wire _19055_;
 wire _19056_;
 wire _19057_;
 wire _19058_;
 wire _19059_;
 wire _19060_;
 wire _19061_;
 wire _19062_;
 wire _19063_;
 wire _19064_;
 wire _19065_;
 wire _19066_;
 wire _19067_;
 wire _19068_;
 wire _19069_;
 wire _19070_;
 wire _19071_;
 wire _19072_;
 wire _19073_;
 wire _19074_;
 wire _19075_;
 wire _19076_;
 wire _19077_;
 wire _19078_;
 wire _19079_;
 wire _19080_;
 wire _19081_;
 wire _19082_;
 wire _19083_;
 wire _19084_;
 wire _19085_;
 wire _19086_;
 wire _19087_;
 wire _19088_;
 wire _19089_;
 wire _19090_;
 wire _19091_;
 wire _19092_;
 wire _19093_;
 wire _19094_;
 wire _19095_;
 wire _19096_;
 wire _19097_;
 wire _19098_;
 wire _19099_;
 wire _19100_;
 wire _19101_;
 wire _19102_;
 wire _19103_;
 wire _19104_;
 wire _19105_;
 wire _19106_;
 wire _19107_;
 wire _19108_;
 wire _19109_;
 wire _19110_;
 wire _19111_;
 wire _19112_;
 wire _19113_;
 wire _19114_;
 wire _19115_;
 wire _19116_;
 wire _19117_;
 wire _19118_;
 wire _19119_;
 wire _19120_;
 wire _19121_;
 wire _19122_;
 wire _19123_;
 wire _19124_;
 wire _19125_;
 wire _19126_;
 wire _19127_;
 wire _19128_;
 wire _19129_;
 wire _19130_;
 wire _19131_;
 wire _19132_;
 wire _19133_;
 wire _19134_;
 wire _19135_;
 wire _19136_;
 wire _19137_;
 wire _19138_;
 wire _19139_;
 wire _19140_;
 wire _19141_;
 wire _19142_;
 wire _19143_;
 wire _19144_;
 wire _19145_;
 wire _19146_;
 wire _19147_;
 wire _19148_;
 wire _19149_;
 wire _19150_;
 wire _19151_;
 wire _19152_;
 wire _19153_;
 wire _19154_;
 wire _19155_;
 wire _19156_;
 wire _19157_;
 wire _19158_;
 wire _19159_;
 wire _19160_;
 wire _19161_;
 wire _19162_;
 wire _19163_;
 wire _19164_;
 wire _19165_;
 wire _19166_;
 wire _19167_;
 wire _19168_;
 wire _19169_;
 wire _19170_;
 wire _19171_;
 wire _19172_;
 wire _19173_;
 wire _19174_;
 wire _19175_;
 wire _19176_;
 wire _19177_;
 wire _19178_;
 wire _19179_;
 wire _19180_;
 wire _19181_;
 wire _19182_;
 wire _19183_;
 wire _19184_;
 wire _19185_;
 wire _19186_;
 wire _19187_;
 wire _19188_;
 wire _19189_;
 wire _19190_;
 wire _19191_;
 wire _19192_;
 wire _19193_;
 wire _19194_;
 wire _19195_;
 wire _19196_;
 wire _19197_;
 wire _19198_;
 wire _19199_;
 wire _19200_;
 wire _19201_;
 wire _19202_;
 wire _19203_;
 wire _19204_;
 wire _19205_;
 wire _19206_;
 wire _19207_;
 wire _19208_;
 wire _19209_;
 wire _19210_;
 wire _19211_;
 wire _19212_;
 wire _19213_;
 wire _19214_;
 wire _19215_;
 wire _19216_;
 wire _19217_;
 wire _19218_;
 wire _19219_;
 wire _19220_;
 wire _19221_;
 wire _19222_;
 wire _19223_;
 wire _19224_;
 wire _19225_;
 wire _19226_;
 wire _19227_;
 wire _19228_;
 wire _19229_;
 wire _19230_;
 wire _19231_;
 wire _19232_;
 wire _19233_;
 wire _19234_;
 wire _19235_;
 wire _19236_;
 wire _19237_;
 wire _19238_;
 wire _19239_;
 wire _19240_;
 wire _19241_;
 wire _19242_;
 wire _19243_;
 wire _19244_;
 wire _19245_;
 wire _19246_;
 wire _19247_;
 wire _19248_;
 wire _19249_;
 wire _19250_;
 wire _19251_;
 wire _19252_;
 wire _19253_;
 wire _19254_;
 wire _19255_;
 wire _19256_;
 wire _19257_;
 wire _19258_;
 wire _19259_;
 wire _19260_;
 wire _19261_;
 wire _19262_;
 wire _19263_;
 wire _19264_;
 wire _19265_;
 wire _19266_;
 wire _19267_;
 wire _19268_;
 wire _19269_;
 wire _19270_;
 wire _19271_;
 wire _19272_;
 wire _19273_;
 wire _19274_;
 wire _19275_;
 wire _19276_;
 wire _19277_;
 wire _19278_;
 wire _19279_;
 wire _19280_;
 wire _19281_;
 wire _19282_;
 wire _19283_;
 wire _19284_;
 wire _19285_;
 wire _19286_;
 wire _19287_;
 wire _19288_;
 wire _19289_;
 wire _19290_;
 wire _19291_;
 wire _19292_;
 wire _19293_;
 wire _19294_;
 wire _19295_;
 wire _19296_;
 wire _19297_;
 wire _19298_;
 wire _19299_;
 wire _19300_;
 wire _19301_;
 wire _19302_;
 wire _19303_;
 wire _19304_;
 wire _19305_;
 wire _19306_;
 wire _19307_;
 wire _19308_;
 wire _19309_;
 wire _19310_;
 wire _19311_;
 wire _19312_;
 wire _19313_;
 wire _19314_;
 wire _19315_;
 wire _19316_;
 wire _19317_;
 wire _19318_;
 wire _19319_;
 wire _19320_;
 wire _19321_;
 wire _19322_;
 wire _19323_;
 wire _19324_;
 wire _19325_;
 wire _19326_;
 wire _19327_;
 wire _19328_;
 wire _19329_;
 wire _19330_;
 wire _19331_;
 wire _19332_;
 wire _19333_;
 wire _19334_;
 wire _19335_;
 wire _19336_;
 wire _19337_;
 wire _19338_;
 wire _19339_;
 wire _19340_;
 wire _19341_;
 wire _19342_;
 wire _19343_;
 wire _19344_;
 wire _19345_;
 wire _19346_;
 wire _19347_;
 wire _19348_;
 wire _19349_;
 wire _19350_;
 wire _19351_;
 wire _19352_;
 wire _19353_;
 wire _19354_;
 wire _19355_;
 wire _19356_;
 wire _19357_;
 wire _19358_;
 wire _19359_;
 wire _19360_;
 wire _19361_;
 wire _19362_;
 wire _19363_;
 wire _19364_;
 wire _19365_;
 wire _19366_;
 wire _19367_;
 wire _19368_;
 wire _19369_;
 wire _19370_;
 wire _19371_;
 wire _19372_;
 wire _19373_;
 wire _19374_;
 wire _19375_;
 wire _19376_;
 wire _19377_;
 wire _19378_;
 wire _19379_;
 wire _19380_;
 wire _19381_;
 wire _19382_;
 wire _19383_;
 wire _19384_;
 wire _19385_;
 wire _19386_;
 wire _19387_;
 wire _19388_;
 wire _19389_;
 wire _19390_;
 wire _19391_;
 wire _19392_;
 wire _19393_;
 wire _19394_;
 wire _19395_;
 wire _19396_;
 wire _19397_;
 wire _19398_;
 wire _19399_;
 wire _19400_;
 wire _19401_;
 wire _19402_;
 wire _19403_;
 wire _19404_;
 wire _19405_;
 wire _19406_;
 wire _19407_;
 wire _19408_;
 wire _19409_;
 wire _19410_;
 wire _19411_;
 wire _19412_;
 wire _19413_;
 wire _19414_;
 wire _19415_;
 wire _19416_;
 wire _19417_;
 wire _19418_;
 wire _19419_;
 wire _19420_;
 wire _19421_;
 wire _19422_;
 wire _19423_;
 wire _19424_;
 wire _19425_;
 wire _19426_;
 wire _19427_;
 wire _19428_;
 wire _19429_;
 wire _19430_;
 wire _19431_;
 wire _19432_;
 wire _19433_;
 wire _19434_;
 wire _19435_;
 wire _19436_;
 wire _19437_;
 wire _19438_;
 wire _19439_;
 wire _19440_;
 wire _19441_;
 wire _19442_;
 wire _19443_;
 wire _19444_;
 wire _19445_;
 wire _19446_;
 wire _19447_;
 wire _19448_;
 wire _19449_;
 wire _19450_;
 wire _19451_;
 wire _19452_;
 wire _19453_;
 wire _19454_;
 wire _19455_;
 wire _19456_;
 wire _19457_;
 wire _19458_;
 wire _19459_;
 wire _19460_;
 wire _19461_;
 wire _19462_;
 wire _19463_;
 wire _19464_;
 wire _19465_;
 wire _19466_;
 wire _19467_;
 wire _19468_;
 wire _19469_;
 wire _19470_;
 wire _19471_;
 wire _19472_;
 wire _19473_;
 wire _19474_;
 wire _19475_;
 wire _19476_;
 wire _19477_;
 wire _19478_;
 wire _19479_;
 wire _19480_;
 wire _19481_;
 wire _19482_;
 wire _19483_;
 wire _19484_;
 wire _19485_;
 wire _19486_;
 wire _19487_;
 wire _19488_;
 wire _19489_;
 wire _19490_;
 wire _19491_;
 wire _19492_;
 wire _19493_;
 wire _19494_;
 wire _19495_;
 wire _19496_;
 wire _19497_;
 wire _19498_;
 wire _19499_;
 wire _19500_;
 wire _19501_;
 wire _19502_;
 wire _19503_;
 wire _19504_;
 wire _19505_;
 wire _19506_;
 wire _19507_;
 wire _19508_;
 wire _19509_;
 wire _19510_;
 wire _19511_;
 wire _19512_;
 wire _19513_;
 wire _19514_;
 wire _19515_;
 wire _19516_;
 wire _19517_;
 wire _19518_;
 wire _19519_;
 wire _19520_;
 wire _19521_;
 wire _19522_;
 wire _19523_;
 wire _19524_;
 wire _19525_;
 wire _19526_;
 wire _19527_;
 wire _19528_;
 wire _19529_;
 wire _19530_;
 wire _19531_;
 wire _19532_;
 wire _19533_;
 wire _19534_;
 wire _19535_;
 wire _19536_;
 wire _19537_;
 wire _19538_;
 wire _19539_;
 wire _19540_;
 wire _19541_;
 wire _19542_;
 wire _19543_;
 wire _19544_;
 wire _19545_;
 wire _19546_;
 wire _19547_;
 wire _19548_;
 wire _19549_;
 wire _19550_;
 wire _19551_;
 wire _19552_;
 wire _19553_;
 wire _19554_;
 wire _19555_;
 wire _19556_;
 wire _19557_;
 wire _19558_;
 wire _19559_;
 wire _19560_;
 wire _19561_;
 wire _19562_;
 wire _19563_;
 wire _19564_;
 wire _19565_;
 wire _19566_;
 wire _19567_;
 wire _19568_;
 wire _19569_;
 wire _19570_;
 wire _19571_;
 wire _19572_;
 wire _19573_;
 wire _19574_;
 wire _19575_;
 wire _19576_;
 wire _19577_;
 wire _19578_;
 wire _19579_;
 wire _19580_;
 wire _19581_;
 wire _19582_;
 wire _19583_;
 wire _19584_;
 wire _19585_;
 wire _19586_;
 wire _19587_;
 wire _19588_;
 wire _19589_;
 wire _19590_;
 wire _19591_;
 wire _19592_;
 wire _19593_;
 wire _19594_;
 wire _19595_;
 wire _19596_;
 wire _19597_;
 wire _19598_;
 wire _19599_;
 wire _19600_;
 wire _19601_;
 wire _19602_;
 wire _19603_;
 wire _19604_;
 wire _19605_;
 wire _19606_;
 wire _19607_;
 wire _19608_;
 wire _19609_;
 wire _19610_;
 wire _19611_;
 wire _19612_;
 wire _19613_;
 wire _19614_;
 wire _19615_;
 wire _19616_;
 wire _19617_;
 wire _19618_;
 wire _19619_;
 wire _19620_;
 wire _19621_;
 wire _19622_;
 wire _19623_;
 wire _19624_;
 wire _19625_;
 wire _19626_;
 wire _19627_;
 wire _19628_;
 wire _19629_;
 wire _19630_;
 wire _19631_;
 wire _19632_;
 wire _19633_;
 wire _19634_;
 wire _19635_;
 wire _19636_;
 wire _19637_;
 wire _19638_;
 wire _19639_;
 wire _19640_;
 wire _19641_;
 wire _19642_;
 wire _19643_;
 wire _19644_;
 wire _19645_;
 wire _19646_;
 wire _19647_;
 wire _19648_;
 wire _19649_;
 wire _19650_;
 wire _19651_;
 wire _19652_;
 wire _19653_;
 wire _19654_;
 wire _19655_;
 wire _19656_;
 wire _19657_;
 wire _19658_;
 wire _19659_;
 wire _19660_;
 wire _19661_;
 wire _19662_;
 wire _19663_;
 wire _19664_;
 wire _19665_;
 wire _19666_;
 wire _19667_;
 wire _19668_;
 wire _19669_;
 wire _19670_;
 wire _19671_;
 wire _19672_;
 wire _19673_;
 wire _19674_;
 wire _19675_;
 wire _19676_;
 wire _19677_;
 wire _19678_;
 wire _19679_;
 wire _19680_;
 wire _19681_;
 wire _19682_;
 wire _19683_;
 wire _19684_;
 wire _19685_;
 wire _19686_;
 wire _19687_;
 wire _19688_;
 wire _19689_;
 wire _19690_;
 wire _19691_;
 wire _19692_;
 wire _19693_;
 wire _19694_;
 wire _19695_;
 wire _19696_;
 wire _19697_;
 wire _19698_;
 wire _19699_;
 wire _19700_;
 wire _19701_;
 wire _19702_;
 wire _19703_;
 wire _19704_;
 wire _19705_;
 wire _19706_;
 wire _19707_;
 wire _19708_;
 wire _19709_;
 wire _19710_;
 wire _19711_;
 wire _19712_;
 wire _19713_;
 wire _19714_;
 wire _19715_;
 wire _19716_;
 wire _19717_;
 wire _19718_;
 wire _19719_;
 wire _19720_;
 wire _19721_;
 wire _19722_;
 wire _19723_;
 wire _19724_;
 wire _19725_;
 wire _19726_;
 wire _19727_;
 wire _19728_;
 wire _19729_;
 wire _19730_;
 wire _19731_;
 wire _19732_;
 wire _19733_;
 wire _19734_;
 wire _19735_;
 wire _19736_;
 wire _19737_;
 wire _19738_;
 wire _19739_;
 wire _19740_;
 wire _19741_;
 wire _19742_;
 wire _19743_;
 wire _19744_;
 wire _19745_;
 wire _19746_;
 wire _19747_;
 wire _19748_;
 wire _19749_;
 wire _19750_;
 wire _19751_;
 wire _19752_;
 wire _19753_;
 wire _19754_;
 wire _19755_;
 wire _19756_;
 wire _19757_;
 wire _19758_;
 wire _19759_;
 wire _19760_;
 wire _19761_;
 wire _19762_;
 wire _19763_;
 wire _19764_;
 wire _19765_;
 wire _19766_;
 wire _19767_;
 wire _19768_;
 wire _19769_;
 wire _19770_;
 wire _19771_;
 wire _19772_;
 wire _19773_;
 wire _19774_;
 wire _19775_;
 wire _19776_;
 wire _19777_;
 wire _19778_;
 wire _19779_;
 wire _19780_;
 wire _19781_;
 wire _19782_;
 wire _19783_;
 wire _19784_;
 wire _19785_;
 wire _19786_;
 wire _19787_;
 wire _19788_;
 wire _19789_;
 wire _19790_;
 wire _19791_;
 wire _19792_;
 wire _19793_;
 wire _19794_;
 wire _19795_;
 wire _19796_;
 wire _19797_;
 wire _19798_;
 wire _19799_;
 wire _19800_;
 wire _19801_;
 wire _19802_;
 wire _19803_;
 wire _19804_;
 wire _19805_;
 wire _19806_;
 wire _19807_;
 wire _19808_;
 wire _19809_;
 wire _19810_;
 wire _19811_;
 wire _19812_;
 wire _19813_;
 wire _19814_;
 wire _19815_;
 wire _19816_;
 wire _19817_;
 wire _19818_;
 wire _19819_;
 wire _19820_;
 wire _19821_;
 wire _19822_;
 wire _19823_;
 wire _19824_;
 wire _19825_;
 wire _19826_;
 wire _19827_;
 wire _19828_;
 wire _19829_;
 wire _19830_;
 wire _19831_;
 wire _19832_;
 wire _19833_;
 wire _19834_;
 wire _19835_;
 wire _19836_;
 wire _19837_;
 wire _19838_;
 wire _19839_;
 wire _19840_;
 wire _19841_;
 wire _19842_;
 wire _19843_;
 wire _19844_;
 wire _19845_;
 wire _19846_;
 wire _19847_;
 wire _19848_;
 wire _19849_;
 wire _19850_;
 wire _19851_;
 wire _19852_;
 wire _19853_;
 wire _19854_;
 wire _19855_;
 wire _19856_;
 wire _19857_;
 wire _19858_;
 wire _19859_;
 wire _19860_;
 wire _19861_;
 wire _19862_;
 wire _19863_;
 wire _19864_;
 wire _19865_;
 wire _19866_;
 wire _19867_;
 wire _19868_;
 wire _19869_;
 wire _19870_;
 wire _19871_;
 wire _19872_;
 wire _19873_;
 wire _19874_;
 wire _19875_;
 wire _19876_;
 wire _19877_;
 wire _19878_;
 wire _19879_;
 wire _19880_;
 wire _19881_;
 wire _19882_;
 wire _19883_;
 wire _19884_;
 wire _19885_;
 wire _19886_;
 wire _19887_;
 wire _19888_;
 wire _19889_;
 wire _19890_;
 wire _19891_;
 wire _19892_;
 wire _19893_;
 wire _19894_;
 wire _19895_;
 wire _19896_;
 wire _19897_;
 wire _19898_;
 wire _19899_;
 wire _19900_;
 wire _19901_;
 wire _19902_;
 wire _19903_;
 wire _19904_;
 wire _19905_;
 wire _19906_;
 wire _19907_;
 wire _19908_;
 wire _19909_;
 wire _19910_;
 wire _19911_;
 wire _19912_;
 wire _19913_;
 wire _19914_;
 wire _19915_;
 wire _19916_;
 wire _19917_;
 wire _19918_;
 wire _19919_;
 wire _19920_;
 wire _19921_;
 wire _19922_;
 wire _19923_;
 wire _19924_;
 wire _19925_;
 wire _19926_;
 wire _19927_;
 wire _19928_;
 wire _19929_;
 wire _19930_;
 wire _19931_;
 wire _19932_;
 wire _19933_;
 wire _19934_;
 wire _19935_;
 wire _19936_;
 wire _19937_;
 wire _19938_;
 wire _19939_;
 wire _19940_;
 wire _19941_;
 wire _19942_;
 wire _19943_;
 wire _19944_;
 wire _19945_;
 wire _19946_;
 wire _19947_;
 wire _19948_;
 wire _19949_;
 wire _19950_;
 wire _19951_;
 wire _19952_;
 wire _19953_;
 wire _19954_;
 wire _19955_;
 wire _19956_;
 wire _19957_;
 wire _19958_;
 wire _19959_;
 wire _19960_;
 wire _19961_;
 wire _19962_;
 wire _19963_;
 wire _19964_;
 wire _19965_;
 wire _19966_;
 wire _19967_;
 wire _19968_;
 wire _19969_;
 wire _19970_;
 wire _19971_;
 wire _19972_;
 wire _19973_;
 wire _19974_;
 wire _19975_;
 wire _19976_;
 wire _19977_;
 wire _19978_;
 wire _19979_;
 wire _19980_;
 wire _19981_;
 wire _19982_;
 wire _19983_;
 wire _19984_;
 wire _19985_;
 wire _19986_;
 wire _19987_;
 wire _19988_;
 wire _19989_;
 wire _19990_;
 wire _19991_;
 wire _19992_;
 wire _19993_;
 wire _19994_;
 wire _19995_;
 wire _19996_;
 wire _19997_;
 wire _19998_;
 wire _19999_;
 wire _20000_;
 wire _20001_;
 wire _20002_;
 wire _20003_;
 wire _20004_;
 wire _20005_;
 wire _20006_;
 wire _20007_;
 wire _20008_;
 wire _20009_;
 wire _20010_;
 wire _20011_;
 wire _20012_;
 wire _20013_;
 wire _20014_;
 wire _20015_;
 wire _20016_;
 wire _20017_;
 wire _20018_;
 wire _20019_;
 wire _20020_;
 wire _20021_;
 wire _20022_;
 wire _20023_;
 wire _20024_;
 wire _20025_;
 wire _20026_;
 wire _20027_;
 wire _20028_;
 wire _20029_;
 wire _20030_;
 wire _20031_;
 wire _20032_;
 wire _20033_;
 wire _20034_;
 wire _20035_;
 wire _20036_;
 wire _20037_;
 wire _20038_;
 wire _20039_;
 wire _20040_;
 wire _20041_;
 wire _20042_;
 wire _20043_;
 wire _20044_;
 wire _20045_;
 wire _20046_;
 wire _20047_;
 wire _20048_;
 wire _20049_;
 wire _20050_;
 wire _20051_;
 wire _20052_;
 wire _20053_;
 wire _20054_;
 wire _20055_;
 wire _20056_;
 wire _20057_;
 wire _20058_;
 wire _20059_;
 wire _20060_;
 wire _20061_;
 wire _20062_;
 wire _20063_;
 wire _20064_;
 wire _20065_;
 wire _20066_;
 wire _20067_;
 wire _20068_;
 wire _20069_;
 wire _20070_;
 wire _20071_;
 wire _20072_;
 wire _20073_;
 wire _20074_;
 wire _20075_;
 wire _20076_;
 wire _20077_;
 wire _20078_;
 wire _20079_;
 wire _20080_;
 wire _20081_;
 wire _20082_;
 wire _20083_;
 wire _20084_;
 wire _20085_;
 wire _20086_;
 wire _20087_;
 wire _20088_;
 wire _20089_;
 wire _20090_;
 wire _20091_;
 wire _20092_;
 wire _20093_;
 wire _20094_;
 wire _20095_;
 wire _20096_;
 wire _20097_;
 wire _20098_;
 wire _20099_;
 wire _20100_;
 wire _20101_;
 wire _20102_;
 wire _20103_;
 wire _20104_;
 wire _20105_;
 wire _20106_;
 wire _20107_;
 wire _20108_;
 wire _20109_;
 wire _20110_;
 wire _20111_;
 wire _20112_;
 wire _20113_;
 wire _20114_;
 wire _20115_;
 wire _20116_;
 wire _20117_;
 wire _20118_;
 wire _20119_;
 wire _20120_;
 wire _20121_;
 wire _20122_;
 wire _20123_;
 wire _20124_;
 wire _20125_;
 wire _20126_;
 wire _20127_;
 wire _20128_;
 wire _20129_;
 wire _20130_;
 wire _20131_;
 wire _20132_;
 wire _20133_;
 wire _20134_;
 wire _20135_;
 wire _20136_;
 wire _20137_;
 wire _20138_;
 wire _20139_;
 wire _20140_;
 wire _20141_;
 wire _20142_;
 wire _20143_;
 wire _20144_;
 wire _20145_;
 wire _20146_;
 wire _20147_;
 wire _20148_;
 wire _20149_;
 wire _20150_;
 wire _20151_;
 wire _20152_;
 wire _20153_;
 wire _20154_;
 wire _20155_;
 wire _20156_;
 wire _20157_;
 wire _20158_;
 wire _20159_;
 wire _20160_;
 wire _20161_;
 wire _20162_;
 wire _20163_;
 wire _20164_;
 wire _20165_;
 wire _20166_;
 wire _20167_;
 wire _20168_;
 wire _20169_;
 wire _20170_;
 wire _20171_;
 wire _20172_;
 wire _20173_;
 wire _20174_;
 wire _20175_;
 wire _20176_;
 wire _20177_;
 wire _20178_;
 wire _20179_;
 wire _20180_;
 wire _20181_;
 wire _20182_;
 wire _20183_;
 wire _20184_;
 wire _20185_;
 wire _20186_;
 wire _20187_;
 wire _20188_;
 wire _20189_;
 wire _20190_;
 wire _20191_;
 wire _20192_;
 wire _20193_;
 wire _20194_;
 wire _20195_;
 wire _20196_;
 wire _20197_;
 wire _20198_;
 wire _20199_;
 wire _20200_;
 wire _20201_;
 wire _20202_;
 wire _20203_;
 wire _20204_;
 wire _20205_;
 wire _20206_;
 wire _20207_;
 wire _20208_;
 wire _20209_;
 wire _20210_;
 wire _20211_;
 wire _20212_;
 wire _20213_;
 wire _20214_;
 wire _20215_;
 wire _20216_;
 wire _20217_;
 wire _20218_;
 wire _20219_;
 wire _20220_;
 wire _20221_;
 wire _20222_;
 wire _20223_;
 wire _20224_;
 wire _20225_;
 wire _20226_;
 wire _20227_;
 wire _20228_;
 wire _20229_;
 wire _20230_;
 wire _20231_;
 wire _20232_;
 wire _20233_;
 wire _20234_;
 wire _20235_;
 wire _20236_;
 wire _20237_;
 wire _20238_;
 wire _20239_;
 wire _20240_;
 wire _20241_;
 wire _20242_;
 wire _20243_;
 wire _20244_;
 wire _20245_;
 wire _20246_;
 wire _20247_;
 wire _20248_;
 wire _20249_;
 wire _20250_;
 wire _20251_;
 wire _20252_;
 wire _20253_;
 wire _20254_;
 wire _20255_;
 wire _20256_;
 wire _20257_;
 wire _20258_;
 wire _20259_;
 wire _20260_;
 wire _20261_;
 wire _20262_;
 wire _20263_;
 wire _20264_;
 wire _20265_;
 wire _20266_;
 wire _20267_;
 wire _20268_;
 wire _20269_;
 wire _20270_;
 wire _20271_;
 wire _20272_;
 wire _20273_;
 wire _20274_;
 wire _20275_;
 wire _20276_;
 wire _20277_;
 wire _20278_;
 wire _20279_;
 wire _20280_;
 wire _20281_;
 wire _20282_;
 wire _20283_;
 wire _20284_;
 wire _20285_;
 wire _20286_;
 wire _20287_;
 wire _20288_;
 wire _20289_;
 wire _20290_;
 wire _20291_;
 wire _20292_;
 wire _20293_;
 wire _20294_;
 wire _20295_;
 wire _20296_;
 wire _20297_;
 wire _20298_;
 wire _20299_;
 wire _20300_;
 wire _20301_;
 wire _20302_;
 wire _20303_;
 wire _20304_;
 wire _20305_;
 wire _20306_;
 wire _20307_;
 wire _20308_;
 wire _20309_;
 wire _20310_;
 wire _20311_;
 wire _20312_;
 wire _20313_;
 wire _20314_;
 wire _20315_;
 wire _20316_;
 wire _20317_;
 wire _20318_;
 wire _20319_;
 wire _20320_;
 wire _20321_;
 wire _20322_;
 wire _20323_;
 wire _20324_;
 wire _20325_;
 wire _20326_;
 wire _20327_;
 wire _20328_;
 wire _20329_;
 wire _20330_;
 wire _20331_;
 wire _20332_;
 wire _20333_;
 wire _20334_;
 wire _20335_;
 wire _20336_;
 wire _20337_;
 wire _20338_;
 wire _20339_;
 wire _20340_;
 wire _20341_;
 wire _20342_;
 wire _20343_;
 wire _20344_;
 wire _20345_;
 wire _20346_;
 wire _20347_;
 wire _20348_;
 wire _20349_;
 wire _20350_;
 wire _20351_;
 wire _20352_;
 wire _20353_;
 wire _20354_;
 wire _20355_;
 wire _20356_;
 wire _20357_;
 wire _20358_;
 wire _20359_;
 wire _20360_;
 wire _20361_;
 wire _20362_;
 wire _20363_;
 wire _20364_;
 wire _20365_;
 wire _20366_;
 wire _20367_;
 wire _20368_;
 wire _20369_;
 wire _20370_;
 wire _20371_;
 wire _20372_;
 wire _20373_;
 wire _20374_;
 wire _20375_;
 wire _20376_;
 wire _20377_;
 wire _20378_;
 wire _20379_;
 wire _20380_;
 wire _20381_;
 wire _20382_;
 wire _20383_;
 wire _20384_;
 wire _20385_;
 wire _20386_;
 wire _20387_;
 wire _20388_;
 wire _20389_;
 wire _20390_;
 wire _20391_;
 wire _20392_;
 wire _20393_;
 wire _20394_;
 wire _20395_;
 wire _20396_;
 wire _20397_;
 wire _20398_;
 wire _20399_;
 wire _20400_;
 wire _20401_;
 wire _20402_;
 wire _20403_;
 wire _20404_;
 wire _20405_;
 wire _20406_;
 wire _20407_;
 wire _20408_;
 wire _20409_;
 wire _20410_;
 wire _20411_;
 wire _20412_;
 wire _20413_;
 wire _20414_;
 wire _20415_;
 wire _20416_;
 wire _20417_;
 wire _20418_;
 wire _20419_;
 wire _20420_;
 wire _20421_;
 wire _20422_;
 wire _20423_;
 wire _20424_;
 wire _20425_;
 wire _20426_;
 wire _20427_;
 wire _20428_;
 wire _20429_;
 wire _20430_;
 wire _20431_;
 wire _20432_;
 wire _20433_;
 wire _20434_;
 wire _20435_;
 wire _20436_;
 wire _20437_;
 wire _20438_;
 wire _20439_;
 wire _20440_;
 wire _20441_;
 wire _20442_;
 wire _20443_;
 wire _20444_;
 wire _20445_;
 wire _20446_;
 wire _20447_;
 wire _20448_;
 wire _20449_;
 wire _20450_;
 wire _20451_;
 wire _20452_;
 wire _20453_;
 wire _20454_;
 wire _20455_;
 wire _20456_;
 wire _20457_;
 wire _20458_;
 wire _20459_;
 wire _20460_;
 wire _20461_;
 wire _20462_;
 wire _20463_;
 wire _20464_;
 wire _20465_;
 wire _20466_;
 wire _20467_;
 wire _20468_;
 wire _20469_;
 wire _20470_;
 wire _20471_;
 wire _20472_;
 wire _20473_;
 wire _20474_;
 wire _20475_;
 wire _20476_;
 wire _20477_;
 wire _20478_;
 wire _20479_;
 wire _20480_;
 wire _20481_;
 wire _20482_;
 wire _20483_;
 wire _20484_;
 wire _20485_;
 wire _20486_;
 wire _20487_;
 wire _20488_;
 wire _20489_;
 wire _20490_;
 wire _20491_;
 wire _20492_;
 wire _20493_;
 wire _20494_;
 wire _20495_;
 wire _20496_;
 wire _20497_;
 wire _20498_;
 wire _20499_;
 wire _20500_;
 wire _20501_;
 wire _20502_;
 wire _20503_;
 wire _20504_;
 wire _20505_;
 wire _20506_;
 wire _20507_;
 wire _20508_;
 wire _20509_;
 wire _20510_;
 wire _20511_;
 wire _20512_;
 wire _20513_;
 wire _20514_;
 wire _20515_;
 wire _20516_;
 wire _20517_;
 wire _20518_;
 wire _20519_;
 wire _20520_;
 wire _20521_;
 wire _20522_;
 wire _20523_;
 wire _20524_;
 wire _20525_;
 wire _20526_;
 wire _20527_;
 wire _20528_;
 wire _20529_;
 wire _20530_;
 wire _20531_;
 wire _20532_;
 wire _20533_;
 wire _20534_;
 wire _20535_;
 wire _20536_;
 wire _20537_;
 wire _20538_;
 wire _20539_;
 wire _20540_;
 wire _20541_;
 wire _20542_;
 wire _20543_;
 wire _20544_;
 wire _20545_;
 wire _20546_;
 wire _20547_;
 wire _20548_;
 wire _20549_;
 wire _20550_;
 wire _20551_;
 wire _20552_;
 wire _20553_;
 wire _20554_;
 wire _20555_;
 wire _20556_;
 wire _20557_;
 wire _20558_;
 wire _20559_;
 wire _20560_;
 wire _20561_;
 wire _20562_;
 wire _20563_;
 wire _20564_;
 wire _20565_;
 wire _20566_;
 wire _20567_;
 wire _20568_;
 wire _20569_;
 wire _20570_;
 wire _20571_;
 wire _20572_;
 wire _20573_;
 wire _20574_;
 wire _20575_;
 wire _20576_;
 wire _20577_;
 wire _20578_;
 wire _20579_;
 wire _20580_;
 wire _20581_;
 wire _20582_;
 wire _20583_;
 wire _20584_;
 wire _20585_;
 wire _20586_;
 wire _20587_;
 wire _20588_;
 wire _20589_;
 wire _20590_;
 wire _20591_;
 wire _20592_;
 wire _20593_;
 wire _20594_;
 wire _20595_;
 wire _20596_;
 wire _20597_;
 wire _20598_;
 wire _20599_;
 wire _20600_;
 wire _20601_;
 wire _20602_;
 wire _20603_;
 wire _20604_;
 wire _20605_;
 wire _20606_;
 wire _20607_;
 wire _20608_;
 wire _20609_;
 wire _20610_;
 wire _20611_;
 wire _20612_;
 wire _20613_;
 wire _20614_;
 wire _20615_;
 wire _20616_;
 wire _20617_;
 wire _20618_;
 wire _20619_;
 wire _20620_;
 wire _20621_;
 wire _20622_;
 wire _20623_;
 wire _20624_;
 wire _20625_;
 wire _20626_;
 wire _20627_;
 wire _20628_;
 wire _20629_;
 wire _20630_;
 wire _20631_;
 wire _20632_;
 wire _20633_;
 wire _20634_;
 wire _20635_;
 wire _20636_;
 wire _20637_;
 wire _20638_;
 wire _20639_;
 wire _20640_;
 wire _20641_;
 wire _20642_;
 wire _20643_;
 wire _20644_;
 wire _20645_;
 wire _20646_;
 wire _20647_;
 wire _20648_;
 wire _20649_;
 wire _20650_;
 wire _20651_;
 wire _20652_;
 wire _20653_;
 wire _20654_;
 wire _20655_;
 wire _20656_;
 wire _20657_;
 wire _20658_;
 wire _20659_;
 wire _20660_;
 wire _20661_;
 wire _20662_;
 wire _20663_;
 wire _20664_;
 wire _20665_;
 wire _20666_;
 wire _20667_;
 wire _20668_;
 wire _20669_;
 wire _20670_;
 wire _20671_;
 wire _20672_;
 wire _20673_;
 wire _20674_;
 wire _20675_;
 wire _20676_;
 wire _20677_;
 wire _20678_;
 wire _20679_;
 wire _20680_;
 wire _20681_;
 wire _20682_;
 wire _20683_;
 wire _20684_;
 wire _20685_;
 wire _20686_;
 wire _20687_;
 wire _20688_;
 wire _20689_;
 wire _20690_;
 wire _20691_;
 wire _20692_;
 wire _20693_;
 wire _20694_;
 wire _20695_;
 wire _20696_;
 wire _20697_;
 wire _20698_;
 wire _20699_;
 wire _20700_;
 wire _20701_;
 wire _20702_;
 wire _20703_;
 wire _20704_;
 wire _20705_;
 wire _20706_;
 wire _20707_;
 wire _20708_;
 wire _20709_;
 wire _20710_;
 wire _20711_;
 wire _20712_;
 wire _20713_;
 wire _20714_;
 wire _20715_;
 wire _20716_;
 wire _20717_;
 wire _20718_;
 wire _20719_;
 wire _20720_;
 wire _20721_;
 wire _20722_;
 wire _20723_;
 wire _20724_;
 wire _20725_;
 wire _20726_;
 wire _20727_;
 wire _20728_;
 wire _20729_;
 wire _20730_;
 wire _20731_;
 wire _20732_;
 wire _20733_;
 wire _20734_;
 wire _20735_;
 wire _20736_;
 wire _20737_;
 wire _20738_;
 wire _20739_;
 wire _20740_;
 wire _20741_;
 wire _20742_;
 wire _20743_;
 wire _20744_;
 wire _20745_;
 wire _20746_;
 wire _20747_;
 wire _20748_;
 wire _20749_;
 wire _20750_;
 wire _20751_;
 wire _20752_;
 wire _20753_;
 wire _20754_;
 wire _20755_;
 wire _20756_;
 wire _20757_;
 wire _20758_;
 wire _20759_;
 wire _20760_;
 wire _20761_;
 wire _20762_;
 wire _20763_;
 wire _20764_;
 wire _20765_;
 wire _20766_;
 wire _20767_;
 wire _20768_;
 wire _20769_;
 wire _20770_;
 wire _20771_;
 wire _20772_;
 wire _20773_;
 wire _20774_;
 wire _20775_;
 wire _20776_;
 wire _20777_;
 wire _20778_;
 wire _20779_;
 wire _20780_;
 wire _20781_;
 wire _20782_;
 wire _20783_;
 wire _20784_;
 wire _20785_;
 wire _20786_;
 wire _20787_;
 wire _20788_;
 wire _20789_;
 wire _20790_;
 wire _20791_;
 wire _20792_;
 wire _20793_;
 wire _20794_;
 wire _20795_;
 wire _20796_;
 wire _20797_;
 wire _20798_;
 wire _20799_;
 wire _20800_;
 wire _20801_;
 wire _20802_;
 wire _20803_;
 wire _20804_;
 wire _20805_;
 wire _20806_;
 wire _20807_;
 wire _20808_;
 wire _20809_;
 wire _20810_;
 wire _20811_;
 wire _20812_;
 wire _20813_;
 wire _20814_;
 wire _20815_;
 wire _20816_;
 wire _20817_;
 wire _20818_;
 wire _20819_;
 wire _20820_;
 wire _20821_;
 wire _20822_;
 wire _20823_;
 wire _20824_;
 wire _20825_;
 wire _20826_;
 wire _20827_;
 wire _20828_;
 wire _20829_;
 wire _20830_;
 wire _20831_;
 wire _20832_;
 wire _20833_;
 wire _20834_;
 wire _20835_;
 wire _20836_;
 wire _20837_;
 wire _20838_;
 wire _20839_;
 wire _20840_;
 wire _20841_;
 wire _20842_;
 wire _20843_;
 wire _20844_;
 wire _20845_;
 wire _20846_;
 wire _20847_;
 wire _20848_;
 wire _20849_;
 wire _20850_;
 wire _20851_;
 wire _20852_;
 wire _20853_;
 wire _20854_;
 wire _20855_;
 wire _20856_;
 wire _20857_;
 wire _20858_;
 wire _20859_;
 wire _20860_;
 wire _20861_;
 wire _20862_;
 wire _20863_;
 wire _20864_;
 wire _20865_;
 wire _20866_;
 wire _20867_;
 wire _20868_;
 wire _20869_;
 wire _20870_;
 wire _20871_;
 wire _20872_;
 wire _20873_;
 wire _20874_;
 wire _20875_;
 wire _20876_;
 wire _20877_;
 wire _20878_;
 wire _20879_;
 wire _20880_;
 wire _20881_;
 wire _20882_;
 wire _20883_;
 wire _20884_;
 wire _20885_;
 wire _20886_;
 wire _20887_;
 wire _20888_;
 wire _20889_;
 wire _20890_;
 wire _20891_;
 wire _20892_;
 wire _20893_;
 wire _20894_;
 wire _20895_;
 wire _20896_;
 wire _20897_;
 wire _20898_;
 wire _20899_;
 wire _20900_;
 wire _20901_;
 wire _20902_;
 wire _20903_;
 wire _20904_;
 wire _20905_;
 wire _20906_;
 wire _20907_;
 wire _20908_;
 wire _20909_;
 wire _20910_;
 wire _20911_;
 wire _20912_;
 wire _20913_;
 wire _20914_;
 wire _20915_;
 wire _20916_;
 wire _20917_;
 wire _20918_;
 wire _20919_;
 wire _20920_;
 wire _20921_;
 wire _20922_;
 wire _20923_;
 wire _20924_;
 wire _20925_;
 wire _20926_;
 wire _20927_;
 wire _20928_;
 wire _20929_;
 wire _20930_;
 wire _20931_;
 wire _20932_;
 wire _20933_;
 wire _20934_;
 wire _20935_;
 wire _20936_;
 wire _20937_;
 wire _20938_;
 wire _20939_;
 wire _20940_;
 wire _20941_;
 wire _20942_;
 wire _20943_;
 wire _20944_;
 wire _20945_;
 wire _20946_;
 wire _20947_;
 wire _20948_;
 wire _20949_;
 wire _20950_;
 wire _20951_;
 wire _20952_;
 wire _20953_;
 wire _20954_;
 wire _20955_;
 wire _20956_;
 wire _20957_;
 wire _20958_;
 wire _20959_;
 wire _20960_;
 wire _20961_;
 wire _20962_;
 wire _20963_;
 wire _20964_;
 wire _20965_;
 wire _20966_;
 wire _20967_;
 wire _20968_;
 wire _20969_;
 wire _20970_;
 wire _20971_;
 wire _20972_;
 wire _20973_;
 wire _20974_;
 wire _20975_;
 wire _20976_;
 wire _20977_;
 wire _20978_;
 wire _20979_;
 wire _20980_;
 wire _20981_;
 wire _20982_;
 wire _20983_;
 wire _20984_;
 wire _20985_;
 wire _20986_;
 wire _20987_;
 wire _20988_;
 wire _20989_;
 wire _20990_;
 wire _20991_;
 wire _20992_;
 wire _20993_;
 wire _20994_;
 wire _20995_;
 wire _20996_;
 wire _20997_;
 wire _20998_;
 wire _20999_;
 wire _21000_;
 wire _21001_;
 wire _21002_;
 wire _21003_;
 wire _21004_;
 wire _21005_;
 wire _21006_;
 wire _21007_;
 wire _21008_;
 wire _21009_;
 wire _21010_;
 wire _21011_;
 wire _21012_;
 wire _21013_;
 wire _21014_;
 wire _21015_;
 wire _21016_;
 wire _21017_;
 wire _21018_;
 wire _21019_;
 wire _21020_;
 wire _21021_;
 wire _21022_;
 wire _21023_;
 wire _21024_;
 wire _21025_;
 wire _21026_;
 wire _21027_;
 wire _21028_;
 wire _21029_;
 wire _21030_;
 wire _21031_;
 wire _21032_;
 wire _21033_;
 wire _21034_;
 wire _21035_;
 wire _21036_;
 wire _21037_;
 wire _21038_;
 wire _21039_;
 wire _21040_;
 wire _21041_;
 wire _21042_;
 wire _21043_;
 wire _21044_;
 wire _21045_;
 wire _21046_;
 wire _21047_;
 wire _21048_;
 wire _21049_;
 wire _21050_;
 wire _21051_;
 wire _21052_;
 wire _21053_;
 wire _21054_;
 wire _21055_;
 wire _21056_;
 wire _21057_;
 wire _21058_;
 wire _21059_;
 wire _21060_;
 wire _21061_;
 wire _21062_;
 wire _21063_;
 wire _21064_;
 wire _21065_;
 wire _21066_;
 wire _21067_;
 wire _21068_;
 wire _21069_;
 wire _21070_;
 wire _21071_;
 wire _21072_;
 wire _21073_;
 wire _21074_;
 wire _21075_;
 wire _21076_;
 wire _21077_;
 wire _21078_;
 wire _21079_;
 wire _21080_;
 wire _21081_;
 wire _21082_;
 wire _21083_;
 wire _21084_;
 wire _21085_;
 wire _21086_;
 wire _21087_;
 wire _21088_;
 wire _21089_;
 wire _21090_;
 wire _21091_;
 wire _21092_;
 wire _21093_;
 wire _21094_;
 wire _21095_;
 wire _21096_;
 wire _21097_;
 wire _21098_;
 wire _21099_;
 wire _21100_;
 wire _21101_;
 wire _21102_;
 wire _21103_;
 wire _21104_;
 wire _21105_;
 wire _21106_;
 wire _21107_;
 wire _21108_;
 wire _21109_;
 wire _21110_;
 wire _21111_;
 wire _21112_;
 wire _21113_;
 wire _21114_;
 wire _21115_;
 wire _21116_;
 wire _21117_;
 wire _21118_;
 wire _21119_;
 wire _21120_;
 wire _21121_;
 wire _21122_;
 wire _21123_;
 wire _21124_;
 wire _21125_;
 wire _21126_;
 wire _21127_;
 wire _21128_;
 wire _21129_;
 wire _21130_;
 wire _21131_;
 wire _21132_;
 wire _21133_;
 wire _21134_;
 wire _21135_;
 wire _21136_;
 wire _21137_;
 wire _21138_;
 wire _21139_;
 wire _21140_;
 wire _21141_;
 wire _21142_;
 wire _21143_;
 wire _21144_;
 wire _21145_;
 wire _21146_;
 wire _21147_;
 wire _21148_;
 wire _21149_;
 wire _21150_;
 wire _21151_;
 wire _21152_;
 wire _21153_;
 wire _21154_;
 wire _21155_;
 wire _21156_;
 wire _21157_;
 wire _21158_;
 wire _21159_;
 wire _21160_;
 wire _21161_;
 wire _21162_;
 wire _21163_;
 wire _21164_;
 wire _21165_;
 wire _21166_;
 wire _21167_;
 wire _21168_;
 wire _21169_;
 wire _21170_;
 wire _21171_;
 wire _21172_;
 wire _21173_;
 wire _21174_;
 wire _21175_;
 wire _21176_;
 wire _21177_;
 wire _21178_;
 wire _21179_;
 wire _21180_;
 wire _21181_;
 wire _21182_;
 wire _21183_;
 wire _21184_;
 wire _21185_;
 wire _21186_;
 wire _21187_;
 wire _21188_;
 wire _21189_;
 wire _21190_;
 wire _21191_;
 wire _21192_;
 wire _21193_;
 wire _21194_;
 wire _21195_;
 wire _21196_;
 wire _21197_;
 wire _21198_;
 wire _21199_;
 wire _21200_;
 wire _21201_;
 wire _21202_;
 wire _21203_;
 wire _21204_;
 wire _21205_;
 wire _21206_;
 wire _21207_;
 wire _21208_;
 wire _21209_;
 wire _21210_;
 wire _21211_;
 wire _21212_;
 wire _21213_;
 wire _21214_;
 wire _21215_;
 wire _21216_;
 wire _21217_;
 wire _21218_;
 wire _21219_;
 wire _21220_;
 wire _21221_;
 wire _21222_;
 wire _21223_;
 wire _21224_;
 wire _21225_;
 wire _21226_;
 wire _21227_;
 wire _21228_;
 wire _21229_;
 wire _21230_;
 wire _21231_;
 wire _21232_;
 wire _21233_;
 wire _21234_;
 wire _21235_;
 wire _21236_;
 wire _21237_;
 wire _21238_;
 wire _21239_;
 wire _21240_;
 wire _21241_;
 wire _21242_;
 wire _21243_;
 wire _21244_;
 wire _21245_;
 wire _21246_;
 wire _21247_;
 wire _21248_;
 wire _21249_;
 wire _21250_;
 wire _21251_;
 wire _21252_;
 wire _21253_;
 wire _21254_;
 wire _21255_;
 wire _21256_;
 wire _21257_;
 wire _21258_;
 wire _21259_;
 wire _21260_;
 wire _21261_;
 wire _21262_;
 wire _21263_;
 wire _21264_;
 wire _21265_;
 wire _21266_;
 wire _21267_;
 wire _21268_;
 wire _21269_;
 wire _21270_;
 wire _21271_;
 wire _21272_;
 wire _21273_;
 wire _21274_;
 wire _21275_;
 wire _21276_;
 wire _21277_;
 wire _21278_;
 wire _21279_;
 wire _21280_;
 wire _21281_;
 wire _21282_;
 wire _21283_;
 wire _21284_;
 wire _21285_;
 wire _21286_;
 wire _21287_;
 wire _21288_;
 wire _21289_;
 wire _21290_;
 wire _21291_;
 wire _21292_;
 wire _21293_;
 wire _21294_;
 wire _21295_;
 wire _21296_;
 wire _21297_;
 wire _21298_;
 wire _21299_;
 wire _21300_;
 wire _21301_;
 wire _21302_;
 wire _21303_;
 wire _21304_;
 wire _21305_;
 wire _21306_;
 wire _21307_;
 wire _21308_;
 wire _21309_;
 wire _21310_;
 wire _21311_;
 wire _21312_;
 wire _21313_;
 wire _21314_;
 wire _21315_;
 wire _21316_;
 wire _21317_;
 wire _21318_;
 wire _21319_;
 wire _21320_;
 wire _21321_;
 wire _21322_;
 wire _21323_;
 wire _21324_;
 wire _21325_;
 wire _21326_;
 wire _21327_;
 wire _21328_;
 wire _21329_;
 wire _21330_;
 wire _21331_;
 wire _21332_;
 wire _21333_;
 wire _21334_;
 wire _21335_;
 wire _21336_;
 wire _21337_;
 wire _21338_;
 wire _21339_;
 wire _21340_;
 wire _21341_;
 wire _21342_;
 wire _21343_;
 wire _21344_;
 wire _21345_;
 wire _21346_;
 wire _21347_;
 wire _21348_;
 wire _21349_;
 wire _21350_;
 wire _21351_;
 wire _21352_;
 wire _21353_;
 wire _21354_;
 wire _21355_;
 wire _21356_;
 wire _21357_;
 wire _21358_;
 wire _21359_;
 wire _21360_;
 wire _21361_;
 wire _21362_;
 wire _21363_;
 wire _21364_;
 wire _21365_;
 wire _21366_;
 wire _21367_;
 wire _21368_;
 wire _21369_;
 wire _21370_;
 wire _21371_;
 wire _21372_;
 wire _21373_;
 wire _21374_;
 wire _21375_;
 wire _21376_;
 wire _21377_;
 wire _21378_;
 wire _21379_;
 wire _21380_;
 wire _21381_;
 wire _21382_;
 wire _21383_;
 wire _21384_;
 wire _21385_;
 wire _21386_;
 wire _21387_;
 wire _21388_;
 wire _21389_;
 wire _21390_;
 wire _21391_;
 wire _21392_;
 wire _21393_;
 wire _21394_;
 wire _21395_;
 wire _21396_;
 wire _21397_;
 wire _21398_;
 wire _21399_;
 wire _21400_;
 wire _21401_;
 wire _21402_;
 wire _21403_;
 wire _21404_;
 wire _21405_;
 wire _21406_;
 wire _21407_;
 wire _21408_;
 wire _21409_;
 wire _21410_;
 wire _21411_;
 wire _21412_;
 wire _21413_;
 wire _21414_;
 wire _21415_;
 wire _21416_;
 wire _21417_;
 wire _21418_;
 wire _21419_;
 wire _21420_;
 wire _21421_;
 wire _21422_;
 wire _21423_;
 wire _21424_;
 wire _21425_;
 wire _21426_;
 wire _21427_;
 wire _21428_;
 wire _21429_;
 wire _21430_;
 wire _21431_;
 wire _21432_;
 wire _21433_;
 wire _21434_;
 wire _21435_;
 wire _21436_;
 wire _21437_;
 wire _21438_;
 wire _21439_;
 wire _21440_;
 wire _21441_;
 wire _21442_;
 wire _21443_;
 wire _21444_;
 wire _21445_;
 wire _21446_;
 wire _21447_;
 wire _21448_;
 wire _21449_;
 wire _21450_;
 wire _21451_;
 wire _21452_;
 wire _21453_;
 wire _21454_;
 wire _21455_;
 wire _21456_;
 wire _21457_;
 wire _21458_;
 wire _21459_;
 wire _21460_;
 wire _21461_;
 wire _21462_;
 wire _21463_;
 wire _21464_;
 wire _21465_;
 wire _21466_;
 wire _21467_;
 wire _21468_;
 wire _21469_;
 wire _21470_;
 wire _21471_;
 wire _21472_;
 wire _21473_;
 wire _21474_;
 wire _21475_;
 wire _21476_;
 wire _21477_;
 wire _21478_;
 wire _21479_;
 wire _21480_;
 wire _21481_;
 wire _21482_;
 wire _21483_;
 wire _21484_;
 wire _21485_;
 wire _21486_;
 wire _21487_;
 wire _21488_;
 wire _21489_;
 wire _21490_;
 wire _21491_;
 wire _21492_;
 wire _21493_;
 wire _21494_;
 wire _21495_;
 wire _21496_;
 wire _21497_;
 wire _21498_;
 wire _21499_;
 wire _21500_;
 wire _21501_;
 wire _21502_;
 wire _21503_;
 wire _21504_;
 wire _21505_;
 wire _21506_;
 wire _21507_;
 wire _21508_;
 wire _21509_;
 wire _21510_;
 wire _21511_;
 wire _21512_;
 wire _21513_;
 wire _21514_;
 wire _21515_;
 wire _21516_;
 wire _21517_;
 wire _21518_;
 wire _21519_;
 wire _21520_;
 wire _21521_;
 wire _21522_;
 wire _21523_;
 wire _21524_;
 wire _21525_;
 wire _21526_;
 wire _21527_;
 wire _21528_;
 wire _21529_;
 wire _21530_;
 wire _21531_;
 wire _21532_;
 wire _21533_;
 wire _21534_;
 wire _21535_;
 wire _21536_;
 wire _21537_;
 wire _21538_;
 wire _21539_;
 wire _21540_;
 wire _21541_;
 wire _21542_;
 wire _21543_;
 wire _21544_;
 wire _21545_;
 wire _21546_;
 wire _21547_;
 wire _21548_;
 wire _21549_;
 wire _21550_;
 wire _21551_;
 wire _21552_;
 wire _21553_;
 wire _21554_;
 wire _21555_;
 wire _21556_;
 wire _21557_;
 wire _21558_;
 wire _21559_;
 wire _21560_;
 wire _21561_;
 wire _21562_;
 wire _21563_;
 wire _21564_;
 wire _21565_;
 wire _21566_;
 wire _21567_;
 wire _21568_;
 wire _21569_;
 wire _21570_;
 wire _21571_;
 wire _21572_;
 wire _21573_;
 wire _21574_;
 wire _21575_;
 wire _21576_;
 wire _21577_;
 wire _21578_;
 wire _21579_;
 wire _21580_;
 wire _21581_;
 wire _21582_;
 wire _21583_;
 wire _21584_;
 wire _21585_;
 wire _21586_;
 wire _21587_;
 wire _21588_;
 wire _21589_;
 wire _21590_;
 wire _21591_;
 wire _21592_;
 wire _21593_;
 wire _21594_;
 wire _21595_;
 wire _21596_;
 wire _21597_;
 wire _21598_;
 wire _21599_;
 wire _21600_;
 wire _21601_;
 wire _21602_;
 wire _21603_;
 wire _21604_;
 wire _21605_;
 wire _21606_;
 wire _21607_;
 wire _21608_;
 wire _21609_;
 wire _21610_;
 wire _21611_;
 wire _21612_;
 wire _21613_;
 wire _21614_;
 wire _21615_;
 wire _21616_;
 wire _21617_;
 wire _21618_;
 wire _21619_;
 wire _21620_;
 wire _21621_;
 wire _21622_;
 wire _21623_;
 wire _21624_;
 wire _21625_;
 wire _21626_;
 wire _21627_;
 wire _21628_;
 wire _21629_;
 wire _21630_;
 wire _21631_;
 wire _21632_;
 wire _21633_;
 wire _21634_;
 wire _21635_;
 wire _21636_;
 wire _21637_;
 wire _21638_;
 wire _21639_;
 wire _21640_;
 wire _21641_;
 wire _21642_;
 wire _21643_;
 wire _21644_;
 wire _21645_;
 wire _21646_;
 wire _21647_;
 wire _21648_;
 wire _21649_;
 wire _21650_;
 wire _21651_;
 wire _21652_;
 wire _21653_;
 wire _21654_;
 wire _21655_;
 wire _21656_;
 wire _21657_;
 wire _21658_;
 wire _21659_;
 wire _21660_;
 wire _21661_;
 wire _21662_;
 wire _21663_;
 wire _21664_;
 wire _21665_;
 wire _21666_;
 wire _21667_;
 wire _21668_;
 wire _21669_;
 wire _21670_;
 wire _21671_;
 wire _21672_;
 wire _21673_;
 wire _21674_;
 wire _21675_;
 wire _21676_;
 wire _21677_;
 wire _21678_;
 wire _21679_;
 wire _21680_;
 wire _21681_;
 wire _21682_;
 wire _21683_;
 wire _21684_;
 wire _21685_;
 wire _21686_;
 wire _21687_;
 wire _21688_;
 wire _21689_;
 wire _21690_;
 wire _21691_;
 wire _21692_;
 wire _21693_;
 wire _21694_;
 wire _21695_;
 wire _21696_;
 wire _21697_;
 wire _21698_;
 wire _21699_;
 wire _21700_;
 wire _21701_;
 wire _21702_;
 wire _21703_;
 wire _21704_;
 wire _21705_;
 wire _21706_;
 wire _21707_;
 wire _21708_;
 wire _21709_;
 wire _21710_;
 wire _21711_;
 wire _21712_;
 wire _21713_;
 wire _21714_;
 wire _21715_;
 wire _21716_;
 wire _21717_;
 wire _21718_;
 wire _21719_;
 wire _21720_;
 wire _21721_;
 wire _21722_;
 wire _21723_;
 wire _21724_;
 wire _21725_;
 wire _21726_;
 wire _21727_;
 wire _21728_;
 wire _21729_;
 wire _21730_;
 wire _21731_;
 wire _21732_;
 wire _21733_;
 wire _21734_;
 wire _21735_;
 wire _21736_;
 wire _21737_;
 wire _21738_;
 wire _21739_;
 wire _21740_;
 wire _21741_;
 wire _21742_;
 wire _21743_;
 wire _21744_;
 wire _21745_;
 wire _21746_;
 wire _21747_;
 wire _21748_;
 wire _21749_;
 wire _21750_;
 wire _21751_;
 wire _21752_;
 wire _21753_;
 wire _21754_;
 wire _21755_;
 wire _21756_;
 wire _21757_;
 wire _21758_;
 wire _21759_;
 wire _21760_;
 wire _21761_;
 wire _21762_;
 wire _21763_;
 wire _21764_;
 wire _21765_;
 wire _21766_;
 wire _21767_;
 wire _21768_;
 wire _21769_;
 wire _21770_;
 wire _21771_;
 wire _21772_;
 wire _21773_;
 wire _21774_;
 wire _21775_;
 wire _21776_;
 wire _21777_;
 wire _21778_;
 wire _21779_;
 wire _21780_;
 wire _21781_;
 wire _21782_;
 wire _21783_;
 wire _21784_;
 wire _21785_;
 wire _21786_;
 wire _21787_;
 wire _21788_;
 wire _21789_;
 wire _21790_;
 wire _21791_;
 wire _21792_;
 wire _21793_;
 wire _21794_;
 wire _21795_;
 wire _21796_;
 wire _21797_;
 wire _21798_;
 wire _21799_;
 wire _21800_;
 wire _21801_;
 wire _21802_;
 wire _21803_;
 wire _21804_;
 wire _21805_;
 wire _21806_;
 wire _21807_;
 wire _21808_;
 wire _21809_;
 wire _21810_;
 wire _21811_;
 wire _21812_;
 wire _21813_;
 wire _21814_;
 wire _21815_;
 wire _21816_;
 wire _21817_;
 wire _21818_;
 wire _21819_;
 wire _21820_;
 wire _21821_;
 wire _21822_;
 wire _21823_;
 wire _21824_;
 wire _21825_;
 wire _21826_;
 wire _21827_;
 wire _21828_;
 wire _21829_;
 wire _21830_;
 wire _21831_;
 wire _21832_;
 wire _21833_;
 wire _21834_;
 wire _21835_;
 wire _21836_;
 wire _21837_;
 wire _21838_;
 wire _21839_;
 wire _21840_;
 wire _21841_;
 wire _21842_;
 wire _21843_;
 wire _21844_;
 wire _21845_;
 wire _21846_;
 wire _21847_;
 wire _21848_;
 wire _21849_;
 wire _21850_;
 wire _21851_;
 wire _21852_;
 wire _21853_;
 wire _21854_;
 wire _21855_;
 wire _21856_;
 wire _21857_;
 wire _21858_;
 wire _21859_;
 wire _21860_;
 wire _21861_;
 wire _21862_;
 wire _21863_;
 wire _21864_;
 wire _21865_;
 wire _21866_;
 wire _21867_;
 wire _21868_;
 wire _21869_;
 wire _21870_;
 wire _21871_;
 wire _21872_;
 wire _21873_;
 wire _21874_;
 wire _21875_;
 wire _21876_;
 wire _21877_;
 wire _21878_;
 wire _21879_;
 wire _21880_;
 wire _21881_;
 wire _21882_;
 wire _21883_;
 wire _21884_;
 wire _21885_;
 wire _21886_;
 wire _21887_;
 wire _21888_;
 wire _21889_;
 wire _21890_;
 wire _21891_;
 wire _21892_;
 wire _21893_;
 wire _21894_;
 wire _21895_;
 wire _21896_;
 wire _21897_;
 wire _21898_;
 wire _21899_;
 wire _21900_;
 wire _21901_;
 wire _21902_;
 wire _21903_;
 wire _21904_;
 wire _21905_;
 wire _21906_;
 wire _21907_;
 wire _21908_;
 wire _21909_;
 wire _21910_;
 wire _21911_;
 wire _21912_;
 wire _21913_;
 wire _21914_;
 wire _21915_;
 wire _21916_;
 wire _21917_;
 wire _21918_;
 wire _21919_;
 wire _21920_;
 wire _21921_;
 wire _21922_;
 wire _21923_;
 wire _21924_;
 wire _21925_;
 wire _21926_;
 wire _21927_;
 wire _21928_;
 wire _21929_;
 wire _21930_;
 wire _21931_;
 wire _21932_;
 wire _21933_;
 wire _21934_;
 wire _21935_;
 wire _21936_;
 wire _21937_;
 wire _21938_;
 wire _21939_;
 wire _21940_;
 wire _21941_;
 wire _21942_;
 wire _21943_;
 wire _21944_;
 wire _21945_;
 wire _21946_;
 wire _21947_;
 wire _21948_;
 wire _21949_;
 wire _21950_;
 wire _21951_;
 wire _21952_;
 wire _21953_;
 wire _21954_;
 wire _21955_;
 wire _21956_;
 wire _21957_;
 wire _21958_;
 wire _21959_;
 wire _21960_;
 wire _21961_;
 wire _21962_;
 wire _21963_;
 wire _21964_;
 wire _21965_;
 wire _21966_;
 wire _21967_;
 wire _21968_;
 wire _21969_;
 wire _21970_;
 wire _21971_;
 wire _21972_;
 wire _21973_;
 wire _21974_;
 wire _21975_;
 wire _21976_;
 wire _21977_;
 wire _21978_;
 wire _21979_;
 wire _21980_;
 wire _21981_;
 wire _21982_;
 wire _21983_;
 wire _21984_;
 wire _21985_;
 wire _21986_;
 wire _21987_;
 wire _21988_;
 wire _21989_;
 wire _21990_;
 wire _21991_;
 wire _21992_;
 wire _21993_;
 wire _21994_;
 wire _21995_;
 wire _21996_;
 wire _21997_;
 wire _21998_;
 wire _21999_;
 wire _22000_;
 wire _22001_;
 wire _22002_;
 wire _22003_;
 wire _22004_;
 wire _22005_;
 wire _22006_;
 wire _22007_;
 wire _22008_;
 wire _22009_;
 wire _22010_;
 wire _22011_;
 wire _22012_;
 wire _22013_;
 wire _22014_;
 wire _22015_;
 wire _22016_;
 wire _22017_;
 wire _22018_;
 wire _22019_;
 wire _22020_;
 wire _22021_;
 wire _22022_;
 wire _22023_;
 wire _22024_;
 wire _22025_;
 wire _22026_;
 wire _22027_;
 wire _22028_;
 wire _22029_;
 wire _22030_;
 wire _22031_;
 wire _22032_;
 wire _22033_;
 wire _22034_;
 wire _22035_;
 wire _22036_;
 wire _22037_;
 wire _22038_;
 wire _22039_;
 wire _22040_;
 wire _22041_;
 wire _22042_;
 wire _22043_;
 wire _22044_;
 wire _22045_;
 wire _22046_;
 wire _22047_;
 wire _22048_;
 wire _22049_;
 wire _22050_;
 wire _22051_;
 wire _22052_;
 wire _22053_;
 wire _22054_;
 wire _22055_;
 wire _22056_;
 wire _22057_;
 wire _22058_;
 wire _22059_;
 wire _22060_;
 wire _22061_;
 wire _22062_;
 wire _22063_;
 wire _22064_;
 wire _22065_;
 wire _22066_;
 wire _22067_;
 wire _22068_;
 wire _22069_;
 wire _22070_;
 wire _22071_;
 wire _22072_;
 wire _22073_;
 wire _22074_;
 wire _22075_;
 wire _22076_;
 wire _22077_;
 wire _22078_;
 wire _22079_;
 wire _22080_;
 wire _22081_;
 wire _22082_;
 wire _22083_;
 wire _22084_;
 wire _22085_;
 wire _22086_;
 wire _22087_;
 wire _22088_;
 wire _22089_;
 wire _22090_;
 wire _22091_;
 wire _22092_;
 wire _22093_;
 wire _22094_;
 wire _22095_;
 wire _22096_;
 wire _22097_;
 wire _22098_;
 wire _22099_;
 wire _22100_;
 wire _22101_;
 wire _22102_;
 wire _22103_;
 wire _22104_;
 wire _22105_;
 wire _22106_;
 wire _22107_;
 wire _22108_;
 wire _22109_;
 wire _22110_;
 wire _22111_;
 wire _22112_;
 wire _22113_;
 wire _22114_;
 wire _22115_;
 wire _22116_;
 wire _22117_;
 wire _22118_;
 wire _22119_;
 wire _22120_;
 wire _22121_;
 wire _22122_;
 wire _22123_;
 wire _22124_;
 wire _22125_;
 wire _22126_;
 wire _22127_;
 wire _22128_;
 wire _22129_;
 wire _22130_;
 wire _22131_;
 wire _22132_;
 wire _22133_;
 wire _22134_;
 wire _22135_;
 wire _22136_;
 wire _22137_;
 wire _22138_;
 wire _22139_;
 wire _22140_;
 wire _22141_;
 wire _22142_;
 wire _22143_;
 wire _22144_;
 wire _22145_;
 wire _22146_;
 wire _22147_;
 wire _22148_;
 wire _22149_;
 wire _22150_;
 wire _22151_;
 wire _22152_;
 wire _22153_;
 wire _22154_;
 wire _22155_;
 wire _22156_;
 wire _22157_;
 wire _22158_;
 wire _22159_;
 wire _22160_;
 wire _22161_;
 wire _22162_;
 wire _22163_;
 wire _22164_;
 wire _22165_;
 wire _22166_;
 wire _22167_;
 wire _22168_;
 wire _22169_;
 wire _22170_;
 wire _22171_;
 wire _22172_;
 wire _22173_;
 wire _22174_;
 wire _22175_;
 wire _22176_;
 wire _22177_;
 wire _22178_;
 wire _22179_;
 wire _22180_;
 wire _22181_;
 wire _22182_;
 wire _22183_;
 wire _22184_;
 wire _22185_;
 wire _22186_;
 wire _22187_;
 wire _22188_;
 wire _22189_;
 wire _22190_;
 wire _22191_;
 wire _22192_;
 wire _22193_;
 wire _22194_;
 wire _22195_;
 wire _22196_;
 wire _22197_;
 wire _22198_;
 wire _22199_;
 wire _22200_;
 wire _22201_;
 wire _22202_;
 wire _22203_;
 wire _22204_;
 wire _22205_;
 wire _22206_;
 wire _22207_;
 wire _22208_;
 wire _22209_;
 wire _22210_;
 wire _22211_;
 wire _22212_;
 wire _22213_;
 wire _22214_;
 wire _22215_;
 wire _22216_;
 wire _22217_;
 wire _22218_;
 wire _22219_;
 wire _22220_;
 wire _22221_;
 wire _22222_;
 wire _22223_;
 wire _22224_;
 wire _22225_;
 wire _22226_;
 wire _22227_;
 wire _22228_;
 wire _22229_;
 wire _22230_;
 wire _22231_;
 wire _22232_;
 wire _22233_;
 wire _22234_;
 wire _22235_;
 wire _22236_;
 wire _22237_;
 wire _22238_;
 wire _22239_;
 wire _22240_;
 wire _22241_;
 wire _22242_;
 wire _22243_;
 wire _22244_;
 wire _22245_;
 wire _22246_;
 wire _22247_;
 wire _22248_;
 wire _22249_;
 wire _22250_;
 wire _22251_;
 wire _22252_;
 wire _22253_;
 wire _22254_;
 wire _22255_;
 wire _22256_;
 wire _22257_;
 wire _22258_;
 wire _22259_;
 wire _22260_;
 wire _22261_;
 wire _22262_;
 wire _22263_;
 wire _22264_;
 wire _22265_;
 wire _22266_;
 wire _22267_;
 wire _22268_;
 wire _22269_;
 wire _22270_;
 wire _22271_;
 wire _22272_;
 wire _22273_;
 wire _22274_;
 wire _22275_;
 wire _22276_;
 wire _22277_;
 wire _22278_;
 wire _22279_;
 wire _22280_;
 wire _22281_;
 wire _22282_;
 wire _22283_;
 wire _22284_;
 wire _22285_;
 wire _22286_;
 wire _22287_;
 wire _22288_;
 wire _22289_;
 wire _22290_;
 wire _22291_;
 wire _22292_;
 wire _22293_;
 wire _22294_;
 wire _22295_;
 wire _22296_;
 wire _22297_;
 wire _22298_;
 wire _22299_;
 wire _22300_;
 wire _22301_;
 wire _22302_;
 wire _22303_;
 wire _22304_;
 wire _22305_;
 wire _22306_;
 wire _22307_;
 wire _22308_;
 wire _22309_;
 wire _22310_;
 wire _22311_;
 wire _22312_;
 wire _22313_;
 wire _22314_;
 wire _22315_;
 wire _22316_;
 wire _22317_;
 wire _22318_;
 wire _22319_;
 wire _22320_;
 wire _22321_;
 wire _22322_;
 wire _22323_;
 wire _22324_;
 wire _22325_;
 wire _22326_;
 wire _22327_;
 wire _22328_;
 wire _22329_;
 wire _22330_;
 wire _22331_;
 wire _22332_;
 wire _22333_;
 wire _22334_;
 wire _22335_;
 wire _22336_;
 wire _22337_;
 wire _22338_;
 wire _22339_;
 wire _22340_;
 wire _22341_;
 wire _22342_;
 wire _22343_;
 wire _22344_;
 wire _22345_;
 wire _22346_;
 wire _22347_;
 wire _22348_;
 wire _22349_;
 wire _22350_;
 wire _22351_;
 wire _22352_;
 wire _22353_;
 wire _22354_;
 wire _22355_;
 wire _22356_;
 wire _22357_;
 wire _22358_;
 wire _22359_;
 wire _22360_;
 wire _22361_;
 wire _22362_;
 wire _22363_;
 wire _22364_;
 wire _22365_;
 wire _22366_;
 wire _22367_;
 wire _22368_;
 wire _22369_;
 wire _22370_;
 wire _22371_;
 wire _22372_;
 wire _22373_;
 wire _22374_;
 wire _22375_;
 wire _22376_;
 wire _22377_;
 wire _22378_;
 wire _22379_;
 wire _22380_;
 wire _22381_;
 wire _22382_;
 wire _22383_;
 wire _22384_;
 wire _22385_;
 wire _22386_;
 wire _22387_;
 wire _22388_;
 wire _22389_;
 wire _22390_;
 wire _22391_;
 wire _22392_;
 wire _22393_;
 wire _22394_;
 wire _22395_;
 wire _22396_;
 wire _22397_;
 wire _22398_;
 wire _22399_;
 wire _22400_;
 wire _22401_;
 wire _22402_;
 wire _22403_;
 wire _22404_;
 wire _22405_;
 wire _22406_;
 wire _22407_;
 wire _22408_;
 wire _22409_;
 wire _22410_;
 wire _22411_;
 wire _22412_;
 wire _22413_;
 wire _22414_;
 wire _22415_;
 wire _22416_;
 wire _22417_;
 wire _22418_;
 wire _22419_;
 wire _22420_;
 wire _22421_;
 wire _22422_;
 wire _22423_;
 wire _22424_;
 wire _22425_;
 wire _22426_;
 wire _22427_;
 wire _22428_;
 wire _22429_;
 wire _22430_;
 wire _22431_;
 wire _22432_;
 wire _22433_;
 wire _22434_;
 wire _22435_;
 wire _22436_;
 wire _22437_;
 wire _22438_;
 wire _22439_;
 wire _22440_;
 wire _22441_;
 wire _22442_;
 wire _22443_;
 wire _22444_;
 wire _22445_;
 wire _22446_;
 wire _22447_;
 wire _22448_;
 wire _22449_;
 wire _22450_;
 wire _22451_;
 wire _22452_;
 wire _22453_;
 wire _22454_;
 wire _22455_;
 wire _22456_;
 wire _22457_;
 wire _22458_;
 wire _22459_;
 wire _22460_;
 wire _22461_;
 wire _22462_;
 wire _22463_;
 wire _22464_;
 wire _22465_;
 wire _22466_;
 wire _22467_;
 wire _22468_;
 wire _22469_;
 wire _22470_;
 wire _22471_;
 wire _22472_;
 wire _22473_;
 wire _22474_;
 wire _22475_;
 wire _22476_;
 wire _22477_;
 wire _22478_;
 wire _22479_;
 wire _22480_;
 wire _22481_;
 wire _22482_;
 wire _22483_;
 wire _22484_;
 wire _22485_;
 wire _22486_;
 wire _22487_;
 wire _22488_;
 wire _22489_;
 wire _22490_;
 wire _22491_;
 wire _22492_;
 wire _22493_;
 wire _22494_;
 wire _22495_;
 wire _22496_;
 wire _22497_;
 wire _22498_;
 wire _22499_;
 wire _22500_;
 wire _22501_;
 wire _22502_;
 wire _22503_;
 wire _22504_;
 wire _22505_;
 wire _22506_;
 wire _22507_;
 wire _22508_;
 wire _22509_;
 wire _22510_;
 wire _22511_;
 wire _22512_;
 wire _22513_;
 wire _22514_;
 wire _22515_;
 wire _22516_;
 wire _22517_;
 wire _22518_;
 wire _22519_;
 wire _22520_;
 wire _22521_;
 wire _22522_;
 wire _22523_;
 wire _22524_;
 wire _22525_;
 wire _22526_;
 wire _22527_;
 wire _22528_;
 wire _22529_;
 wire _22530_;
 wire _22531_;
 wire _22532_;
 wire _22533_;
 wire _22534_;
 wire _22535_;
 wire _22536_;
 wire _22537_;
 wire _22538_;
 wire _22539_;
 wire _22540_;
 wire _22541_;
 wire _22542_;
 wire _22543_;
 wire _22544_;
 wire _22545_;
 wire _22546_;
 wire _22547_;
 wire _22548_;
 wire _22549_;
 wire _22550_;
 wire _22551_;
 wire _22552_;
 wire _22553_;
 wire _22554_;
 wire _22555_;
 wire _22556_;
 wire _22557_;
 wire _22558_;
 wire _22559_;
 wire _22560_;
 wire _22561_;
 wire _22562_;
 wire _22563_;
 wire _22564_;
 wire _22565_;
 wire _22566_;
 wire _22567_;
 wire _22568_;
 wire _22569_;
 wire _22570_;
 wire _22571_;
 wire _22572_;
 wire _22573_;
 wire _22574_;
 wire _22575_;
 wire _22576_;
 wire _22577_;
 wire _22578_;
 wire _22579_;
 wire _22580_;
 wire _22581_;
 wire _22582_;
 wire _22583_;
 wire _22584_;
 wire _22585_;
 wire _22586_;
 wire _22587_;
 wire _22588_;
 wire _22589_;
 wire _22590_;
 wire _22591_;
 wire _22592_;
 wire _22593_;
 wire _22594_;
 wire _22595_;
 wire _22596_;
 wire _22597_;
 wire _22598_;
 wire _22599_;
 wire _22600_;
 wire _22601_;
 wire _22602_;
 wire _22603_;
 wire _22604_;
 wire _22605_;
 wire _22606_;
 wire _22607_;
 wire _22608_;
 wire _22609_;
 wire _22610_;
 wire _22611_;
 wire _22612_;
 wire _22613_;
 wire _22614_;
 wire _22615_;
 wire _22616_;
 wire _22617_;
 wire _22618_;
 wire _22619_;
 wire _22620_;
 wire _22621_;
 wire _22622_;
 wire _22623_;
 wire _22624_;
 wire _22625_;
 wire _22626_;
 wire _22627_;
 wire _22628_;
 wire _22629_;
 wire _22630_;
 wire _22631_;
 wire _22632_;
 wire _22633_;
 wire _22634_;
 wire _22635_;
 wire _22636_;
 wire _22637_;
 wire _22638_;
 wire _22639_;
 wire _22640_;
 wire _22641_;
 wire _22642_;
 wire _22643_;
 wire _22644_;
 wire _22645_;
 wire _22646_;
 wire _22647_;
 wire _22648_;
 wire _22649_;
 wire _22650_;
 wire _22651_;
 wire _22652_;
 wire _22653_;
 wire _22654_;
 wire _22655_;
 wire _22656_;
 wire _22657_;
 wire _22658_;
 wire _22659_;
 wire _22660_;
 wire _22661_;
 wire _22662_;
 wire _22663_;
 wire _22664_;
 wire _22665_;
 wire _22666_;
 wire _22667_;
 wire _22668_;
 wire _22669_;
 wire _22670_;
 wire _22671_;
 wire _22672_;
 wire _22673_;
 wire _22674_;
 wire _22675_;
 wire _22676_;
 wire _22677_;
 wire _22678_;
 wire _22679_;
 wire _22680_;
 wire _22681_;
 wire _22682_;
 wire _22683_;
 wire _22684_;
 wire _22685_;
 wire _22686_;
 wire _22687_;
 wire _22688_;
 wire _22689_;
 wire _22690_;
 wire _22691_;
 wire _22692_;
 wire _22693_;
 wire _22694_;
 wire _22695_;
 wire _22696_;
 wire _22697_;
 wire _22698_;
 wire _22699_;
 wire _22700_;
 wire _22701_;
 wire _22702_;
 wire _22703_;
 wire _22704_;
 wire _22705_;
 wire _22706_;
 wire _22707_;
 wire _22708_;
 wire _22709_;
 wire _22710_;
 wire _22711_;
 wire _22712_;
 wire _22713_;
 wire _22714_;
 wire _22715_;
 wire _22716_;
 wire _22717_;
 wire _22718_;
 wire _22719_;
 wire _22720_;
 wire _22721_;
 wire _22722_;
 wire _22723_;
 wire _22724_;
 wire _22725_;
 wire _22726_;
 wire _22727_;
 wire _22728_;
 wire _22729_;
 wire _22730_;
 wire _22731_;
 wire _22732_;
 wire _22733_;
 wire _22734_;
 wire _22735_;
 wire _22736_;
 wire _22737_;
 wire _22738_;
 wire _22739_;
 wire _22740_;
 wire _22741_;
 wire _22742_;
 wire _22743_;
 wire _22744_;
 wire _22745_;
 wire _22746_;
 wire _22747_;
 wire _22748_;
 wire _22749_;
 wire _22750_;
 wire _22751_;
 wire _22752_;
 wire _22753_;
 wire _22754_;
 wire _22755_;
 wire _22756_;
 wire _22757_;
 wire _22758_;
 wire _22759_;
 wire _22760_;
 wire _22761_;
 wire _22762_;
 wire _22763_;
 wire _22764_;
 wire _22765_;
 wire _22766_;
 wire _22767_;
 wire _22768_;
 wire _22769_;
 wire _22770_;
 wire _22771_;
 wire _22772_;
 wire _22773_;
 wire _22774_;
 wire _22775_;
 wire _22776_;
 wire _22777_;
 wire _22778_;
 wire _22779_;
 wire _22780_;
 wire _22781_;
 wire _22782_;
 wire _22783_;
 wire _22784_;
 wire _22785_;
 wire _22786_;
 wire _22787_;
 wire _22788_;
 wire _22789_;
 wire _22790_;
 wire _22791_;
 wire _22792_;
 wire _22793_;
 wire _22794_;
 wire _22795_;
 wire _22796_;
 wire _22797_;
 wire _22798_;
 wire _22799_;
 wire _22800_;
 wire _22801_;
 wire _22802_;
 wire _22803_;
 wire _22804_;
 wire _22805_;
 wire _22806_;
 wire _22807_;
 wire _22808_;
 wire _22809_;
 wire _22810_;
 wire _22811_;
 wire _22812_;
 wire _22813_;
 wire _22814_;
 wire _22815_;
 wire _22816_;
 wire _22817_;
 wire _22818_;
 wire _22819_;
 wire _22820_;
 wire _22821_;
 wire _22822_;
 wire _22823_;
 wire _22824_;
 wire _22825_;
 wire _22826_;
 wire _22827_;
 wire _22828_;
 wire _22829_;
 wire _22830_;
 wire _22831_;
 wire _22832_;
 wire _22833_;
 wire _22834_;
 wire _22835_;
 wire _22836_;
 wire _22837_;
 wire _22838_;
 wire _22839_;
 wire _22840_;
 wire _22841_;
 wire _22842_;
 wire _22843_;
 wire _22844_;
 wire _22845_;
 wire _22846_;
 wire _22847_;
 wire _22848_;
 wire _22849_;
 wire _22850_;
 wire _22851_;
 wire _22852_;
 wire _22853_;
 wire _22854_;
 wire _22855_;
 wire _22856_;
 wire _22857_;
 wire _22858_;
 wire _22859_;
 wire _22860_;
 wire _22861_;
 wire _22862_;
 wire _22863_;
 wire _22864_;
 wire _22865_;
 wire _22866_;
 wire _22867_;
 wire _22868_;
 wire _22869_;
 wire _22870_;
 wire _22871_;
 wire _22872_;
 wire _22873_;
 wire _22874_;
 wire _22875_;
 wire _22876_;
 wire _22877_;
 wire _22878_;
 wire _22879_;
 wire _22880_;
 wire _22881_;
 wire _22882_;
 wire _22883_;
 wire _22884_;
 wire _22885_;
 wire _22886_;
 wire _22887_;
 wire _22888_;
 wire _22889_;
 wire _22890_;
 wire _22891_;
 wire _22892_;
 wire _22893_;
 wire _22894_;
 wire _22895_;
 wire _22896_;
 wire _22897_;
 wire _22898_;
 wire _22899_;
 wire _22900_;
 wire _22901_;
 wire _22902_;
 wire _22903_;
 wire _22904_;
 wire _22905_;
 wire _22906_;
 wire _22907_;
 wire _22908_;
 wire _22909_;
 wire _22910_;
 wire _22911_;
 wire _22912_;
 wire _22913_;
 wire _22914_;
 wire _22915_;
 wire _22916_;
 wire _22917_;
 wire _22918_;
 wire _22919_;
 wire _22920_;
 wire _22921_;
 wire _22922_;
 wire _22923_;
 wire _22924_;
 wire _22925_;
 wire _22926_;
 wire _22927_;
 wire _22928_;
 wire _22929_;
 wire _22930_;
 wire _22931_;
 wire _22932_;
 wire _22933_;
 wire _22934_;
 wire _22935_;
 wire _22936_;
 wire _22937_;
 wire _22938_;
 wire _22939_;
 wire _22940_;
 wire _22941_;
 wire _22942_;
 wire _22943_;
 wire _22944_;
 wire _22945_;
 wire _22946_;
 wire _22947_;
 wire _22948_;
 wire _22949_;
 wire _22950_;
 wire _22951_;
 wire _22952_;
 wire _22953_;
 wire _22954_;
 wire _22955_;
 wire _22956_;
 wire _22957_;
 wire _22958_;
 wire _22959_;
 wire _22960_;
 wire _22961_;
 wire _22962_;
 wire _22963_;
 wire _22964_;
 wire _22965_;
 wire _22966_;
 wire _22967_;
 wire _22968_;
 wire _22969_;
 wire _22970_;
 wire _22971_;
 wire _22972_;
 wire _22973_;
 wire _22974_;
 wire _22975_;
 wire _22976_;
 wire _22977_;
 wire _22978_;
 wire _22979_;
 wire _22980_;
 wire _22981_;
 wire _22982_;
 wire _22983_;
 wire _22984_;
 wire _22985_;
 wire _22986_;
 wire _22987_;
 wire _22988_;
 wire _22989_;
 wire _22990_;
 wire _22991_;
 wire _22992_;
 wire _22993_;
 wire _22994_;
 wire _22995_;
 wire _22996_;
 wire _22997_;
 wire _22998_;
 wire _22999_;
 wire _23000_;
 wire _23001_;
 wire _23002_;
 wire _23003_;
 wire _23004_;
 wire _23005_;
 wire _23006_;
 wire _23007_;
 wire _23008_;
 wire _23009_;
 wire _23010_;
 wire _23011_;
 wire _23012_;
 wire _23013_;
 wire _23014_;
 wire _23015_;
 wire _23016_;
 wire _23017_;
 wire _23018_;
 wire _23019_;
 wire _23020_;
 wire _23021_;
 wire _23022_;
 wire _23023_;
 wire _23024_;
 wire _23025_;
 wire _23026_;
 wire _23027_;
 wire _23028_;
 wire _23029_;
 wire _23030_;
 wire _23031_;
 wire _23032_;
 wire _23033_;
 wire _23034_;
 wire _23035_;
 wire _23036_;
 wire _23037_;
 wire _23038_;
 wire _23039_;
 wire _23040_;
 wire _23041_;
 wire _23042_;
 wire _23043_;
 wire _23044_;
 wire _23045_;
 wire _23046_;
 wire _23047_;
 wire _23048_;
 wire _23049_;
 wire _23050_;
 wire _23051_;
 wire _23052_;
 wire _23053_;
 wire _23054_;
 wire _23055_;
 wire _23056_;
 wire _23057_;
 wire _23058_;
 wire _23059_;
 wire _23060_;
 wire _23061_;
 wire _23062_;
 wire _23063_;
 wire _23064_;
 wire _23065_;
 wire _23066_;
 wire _23067_;
 wire _23068_;
 wire _23069_;
 wire _23070_;
 wire _23071_;
 wire _23072_;
 wire _23073_;
 wire _23074_;
 wire _23075_;
 wire _23076_;
 wire _23077_;
 wire _23078_;
 wire _23079_;
 wire _23080_;
 wire _23081_;
 wire _23082_;
 wire _23083_;
 wire _23084_;
 wire _23085_;
 wire _23086_;
 wire _23087_;
 wire _23088_;
 wire _23089_;
 wire _23090_;
 wire _23091_;
 wire _23092_;
 wire _23093_;
 wire _23094_;
 wire _23095_;
 wire _23096_;
 wire _23097_;
 wire _23098_;
 wire _23099_;
 wire _23100_;
 wire _23101_;
 wire _23102_;
 wire _23103_;
 wire _23104_;
 wire _23105_;
 wire _23106_;
 wire _23107_;
 wire _23108_;
 wire _23109_;
 wire _23110_;
 wire _23111_;
 wire _23112_;
 wire _23113_;
 wire _23114_;
 wire _23115_;
 wire _23116_;
 wire _23117_;
 wire _23118_;
 wire _23119_;
 wire _23120_;
 wire _23121_;
 wire _23122_;
 wire _23123_;
 wire _23124_;
 wire _23125_;
 wire _23126_;
 wire _23127_;
 wire _23128_;
 wire _23129_;
 wire _23130_;
 wire _23131_;
 wire _23132_;
 wire _23133_;
 wire _23134_;
 wire _23135_;
 wire _23136_;
 wire _23137_;
 wire _23138_;
 wire _23139_;
 wire _23140_;
 wire _23141_;
 wire _23142_;
 wire _23143_;
 wire _23144_;
 wire _23145_;
 wire _23146_;
 wire _23147_;
 wire _23148_;
 wire _23149_;
 wire _23150_;
 wire _23151_;
 wire _23152_;
 wire _23153_;
 wire _23154_;
 wire _23155_;
 wire _23156_;
 wire _23157_;
 wire _23158_;
 wire _23159_;
 wire _23160_;
 wire _23161_;
 wire _23162_;
 wire _23163_;
 wire _23164_;
 wire _23165_;
 wire _23166_;
 wire _23167_;
 wire _23168_;
 wire _23169_;
 wire _23170_;
 wire _23171_;
 wire _23172_;
 wire _23173_;
 wire _23174_;
 wire _23175_;
 wire _23176_;
 wire _23177_;
 wire _23178_;
 wire _23179_;
 wire _23180_;
 wire _23181_;
 wire _23182_;
 wire _23183_;
 wire _23184_;
 wire _23185_;
 wire _23186_;
 wire _23187_;
 wire _23188_;
 wire _23189_;
 wire _23190_;
 wire _23191_;
 wire _23192_;
 wire _23193_;
 wire _23194_;
 wire _23195_;
 wire _23196_;
 wire _23197_;
 wire _23198_;
 wire _23199_;
 wire _23200_;
 wire _23201_;
 wire _23202_;
 wire _23203_;
 wire _23204_;
 wire _23205_;
 wire _23206_;
 wire _23207_;
 wire _23208_;
 wire _23209_;
 wire _23210_;
 wire _23211_;
 wire _23212_;
 wire _23213_;
 wire _23214_;
 wire _23215_;
 wire _23216_;
 wire _23217_;
 wire _23218_;
 wire _23219_;
 wire _23220_;
 wire _23221_;
 wire _23222_;
 wire _23223_;
 wire _23224_;
 wire _23225_;
 wire _23226_;
 wire _23227_;
 wire _23228_;
 wire _23229_;
 wire _23230_;
 wire _23231_;
 wire _23232_;
 wire _23233_;
 wire _23234_;
 wire _23235_;
 wire _23236_;
 wire _23237_;
 wire _23238_;
 wire _23239_;
 wire _23240_;
 wire _23241_;
 wire _23242_;
 wire _23243_;
 wire _23244_;
 wire _23245_;
 wire _23246_;
 wire _23247_;
 wire _23248_;
 wire _23249_;
 wire _23250_;
 wire _23251_;
 wire _23252_;
 wire _23253_;
 wire _23254_;
 wire _23255_;
 wire _23256_;
 wire _23257_;
 wire _23258_;
 wire _23259_;
 wire _23260_;
 wire _23261_;
 wire _23262_;
 wire _23263_;
 wire _23264_;
 wire _23265_;
 wire _23266_;
 wire _23267_;
 wire _23268_;
 wire _23269_;
 wire _23270_;
 wire _23271_;
 wire _23272_;
 wire _23273_;
 wire _23274_;
 wire _23275_;
 wire _23276_;
 wire _23277_;
 wire _23278_;
 wire _23279_;
 wire _23280_;
 wire _23281_;
 wire _23282_;
 wire _23283_;
 wire _23284_;
 wire _23285_;
 wire _23286_;
 wire _23287_;
 wire _23288_;
 wire _23289_;
 wire _23290_;
 wire _23291_;
 wire _23292_;
 wire _23293_;
 wire _23294_;
 wire _23295_;
 wire _23296_;
 wire _23297_;
 wire _23298_;
 wire _23299_;
 wire _23300_;
 wire _23301_;
 wire _23302_;
 wire _23303_;
 wire _23304_;
 wire _23305_;
 wire _23306_;
 wire _23307_;
 wire _23308_;
 wire _23309_;
 wire _23310_;
 wire _23311_;
 wire _23312_;
 wire _23313_;
 wire _23314_;
 wire _23315_;
 wire _23316_;
 wire _23317_;
 wire _23318_;
 wire _23319_;
 wire _23320_;
 wire _23321_;
 wire _23322_;
 wire _23323_;
 wire _23324_;
 wire _23325_;
 wire _23326_;
 wire _23327_;
 wire _23328_;
 wire _23329_;
 wire _23330_;
 wire _23331_;
 wire _23332_;
 wire _23333_;
 wire _23334_;
 wire _23335_;
 wire _23336_;
 wire _23337_;
 wire _23338_;
 wire _23339_;
 wire _23340_;
 wire _23341_;
 wire _23342_;
 wire _23343_;
 wire _23344_;
 wire _23345_;
 wire _23346_;
 wire _23347_;
 wire _23348_;
 wire _23349_;
 wire _23350_;
 wire _23351_;
 wire _23352_;
 wire _23353_;
 wire _23354_;
 wire _23355_;
 wire _23356_;
 wire _23357_;
 wire _23358_;
 wire _23359_;
 wire _23360_;
 wire _23361_;
 wire _23362_;
 wire _23363_;
 wire _23364_;
 wire _23365_;
 wire _23366_;
 wire _23367_;
 wire _23368_;
 wire _23369_;
 wire _23370_;
 wire _23371_;
 wire _23372_;
 wire _23373_;
 wire _23374_;
 wire _23375_;
 wire _23376_;
 wire _23377_;
 wire _23378_;
 wire _23379_;
 wire _23380_;
 wire _23381_;
 wire _23382_;
 wire _23383_;
 wire _23384_;
 wire _23385_;
 wire _23386_;
 wire _23387_;
 wire _23388_;
 wire _23389_;
 wire _23390_;
 wire _23391_;
 wire _23392_;
 wire _23393_;
 wire _23394_;
 wire _23395_;
 wire _23396_;
 wire _23397_;
 wire _23398_;
 wire _23399_;
 wire _23400_;
 wire _23401_;
 wire _23402_;
 wire _23403_;
 wire _23404_;
 wire _23405_;
 wire _23406_;
 wire _23407_;
 wire _23408_;
 wire _23409_;
 wire _23410_;
 wire _23411_;
 wire _23412_;
 wire _23413_;
 wire _23414_;
 wire _23415_;
 wire _23416_;
 wire _23417_;
 wire _23418_;
 wire _23419_;
 wire _23420_;
 wire _23421_;
 wire _23422_;
 wire _23423_;
 wire _23424_;
 wire _23425_;
 wire _23426_;
 wire _23427_;
 wire _23428_;
 wire _23429_;
 wire _23430_;
 wire _23431_;
 wire _23432_;
 wire _23433_;
 wire _23434_;
 wire _23435_;
 wire _23436_;
 wire _23437_;
 wire _23438_;
 wire _23439_;
 wire _23440_;
 wire _23441_;
 wire _23442_;
 wire _23443_;
 wire _23444_;
 wire _23445_;
 wire _23446_;
 wire _23447_;
 wire _23448_;
 wire _23449_;
 wire _23450_;
 wire _23451_;
 wire _23452_;
 wire _23453_;
 wire _23454_;
 wire _23455_;
 wire _23456_;
 wire _23457_;
 wire _23458_;
 wire _23459_;
 wire _23460_;
 wire _23461_;
 wire _23462_;
 wire _23463_;
 wire _23464_;
 wire _23465_;
 wire _23466_;
 wire _23467_;
 wire _23468_;
 wire _23469_;
 wire _23470_;
 wire _23471_;
 wire _23472_;
 wire _23473_;
 wire _23474_;
 wire _23475_;
 wire _23476_;
 wire _23477_;
 wire _23478_;
 wire _23479_;
 wire _23480_;
 wire _23481_;
 wire _23482_;
 wire _23483_;
 wire _23484_;
 wire _23485_;
 wire _23486_;
 wire _23487_;
 wire _23488_;
 wire _23489_;
 wire _23490_;
 wire _23491_;
 wire _23492_;
 wire _23493_;
 wire _23494_;
 wire _23495_;
 wire _23496_;
 wire _23497_;
 wire _23498_;
 wire _23499_;
 wire _23500_;
 wire _23501_;
 wire _23502_;
 wire _23503_;
 wire _23504_;
 wire _23505_;
 wire _23506_;
 wire _23507_;
 wire _23508_;
 wire _23509_;
 wire _23510_;
 wire _23511_;
 wire _23512_;
 wire _23513_;
 wire _23514_;
 wire _23515_;
 wire _23516_;
 wire _23517_;
 wire _23518_;
 wire _23519_;
 wire _23520_;
 wire _23521_;
 wire _23522_;
 wire _23523_;
 wire _23524_;
 wire _23525_;
 wire _23526_;
 wire _23527_;
 wire _23528_;
 wire _23529_;
 wire _23530_;
 wire _23531_;
 wire _23532_;
 wire _23533_;
 wire _23534_;
 wire _23535_;
 wire _23536_;
 wire _23537_;
 wire _23538_;
 wire _23539_;
 wire _23540_;
 wire _23541_;
 wire _23542_;
 wire _23543_;
 wire _23544_;
 wire _23545_;
 wire _23546_;
 wire _23547_;
 wire _23548_;
 wire _23549_;
 wire _23550_;
 wire _23551_;
 wire _23552_;
 wire _23553_;
 wire _23554_;
 wire _23555_;
 wire _23556_;
 wire _23557_;
 wire _23558_;
 wire _23559_;
 wire _23560_;
 wire _23561_;
 wire _23562_;
 wire _23563_;
 wire _23564_;
 wire _23565_;
 wire _23566_;
 wire _23567_;
 wire _23568_;
 wire _23569_;
 wire _23570_;
 wire _23571_;
 wire _23572_;
 wire _23573_;
 wire _23574_;
 wire _23575_;
 wire _23576_;
 wire _23577_;
 wire _23578_;
 wire _23579_;
 wire _23580_;
 wire _23581_;
 wire _23582_;
 wire _23583_;
 wire _23584_;
 wire _23585_;
 wire _23586_;
 wire _23587_;
 wire _23588_;
 wire _23589_;
 wire _23590_;
 wire _23591_;
 wire _23592_;
 wire _23593_;
 wire _23594_;
 wire _23595_;
 wire _23596_;
 wire _23597_;
 wire _23598_;
 wire _23599_;
 wire _23600_;
 wire _23601_;
 wire _23602_;
 wire _23603_;
 wire _23604_;
 wire _23605_;
 wire _23606_;
 wire _23607_;
 wire _23608_;
 wire _23609_;
 wire _23610_;
 wire _23611_;
 wire _23612_;
 wire _23613_;
 wire _23614_;
 wire _23615_;
 wire _23616_;
 wire _23617_;
 wire _23618_;
 wire _23619_;
 wire _23620_;
 wire _23621_;
 wire _23622_;
 wire _23623_;
 wire _23624_;
 wire _23625_;
 wire _23626_;
 wire _23627_;
 wire _23628_;
 wire _23629_;
 wire _23630_;
 wire _23631_;
 wire _23632_;
 wire _23633_;
 wire _23634_;
 wire _23635_;
 wire _23636_;
 wire _23637_;
 wire _23638_;
 wire _23639_;
 wire _23640_;
 wire _23641_;
 wire _23642_;
 wire _23643_;
 wire _23644_;
 wire _23645_;
 wire _23646_;
 wire _23647_;
 wire _23648_;
 wire _23649_;
 wire _23650_;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire accepting;
 wire \byte_cnt[0] ;
 wire \byte_cnt[1] ;
 wire \byte_cnt[2] ;
 wire \byte_cnt[3] ;
 wire \byte_cnt[4] ;
 wire \byte_cnt[5] ;
 wire \inv_cycles[0] ;
 wire \inv_cycles[1] ;
 wire \inv_cycles[2] ;
 wire \inv_cycles[3] ;
 wire \inv_cycles[4] ;
 wire \inv_cycles[5] ;
 wire \inv_cycles[6] ;
 wire \inv_cycles[7] ;
 wire \inv_cycles[8] ;
 wire \inv_cycles[9] ;
 wire inv_done;
 wire inv_go;
 wire \inv_result[0] ;
 wire \inv_result[100] ;
 wire \inv_result[101] ;
 wire \inv_result[102] ;
 wire \inv_result[103] ;
 wire \inv_result[104] ;
 wire \inv_result[105] ;
 wire \inv_result[106] ;
 wire \inv_result[107] ;
 wire \inv_result[108] ;
 wire \inv_result[109] ;
 wire \inv_result[10] ;
 wire \inv_result[110] ;
 wire \inv_result[111] ;
 wire \inv_result[112] ;
 wire \inv_result[113] ;
 wire \inv_result[114] ;
 wire \inv_result[115] ;
 wire \inv_result[116] ;
 wire \inv_result[117] ;
 wire \inv_result[118] ;
 wire \inv_result[119] ;
 wire \inv_result[11] ;
 wire \inv_result[120] ;
 wire \inv_result[121] ;
 wire \inv_result[122] ;
 wire \inv_result[123] ;
 wire \inv_result[124] ;
 wire \inv_result[125] ;
 wire \inv_result[126] ;
 wire \inv_result[127] ;
 wire \inv_result[128] ;
 wire \inv_result[129] ;
 wire \inv_result[12] ;
 wire \inv_result[130] ;
 wire \inv_result[131] ;
 wire \inv_result[132] ;
 wire \inv_result[133] ;
 wire \inv_result[134] ;
 wire \inv_result[135] ;
 wire \inv_result[136] ;
 wire \inv_result[137] ;
 wire \inv_result[138] ;
 wire \inv_result[139] ;
 wire \inv_result[13] ;
 wire \inv_result[140] ;
 wire \inv_result[141] ;
 wire \inv_result[142] ;
 wire \inv_result[143] ;
 wire \inv_result[144] ;
 wire \inv_result[145] ;
 wire \inv_result[146] ;
 wire \inv_result[147] ;
 wire \inv_result[148] ;
 wire \inv_result[149] ;
 wire \inv_result[14] ;
 wire \inv_result[150] ;
 wire \inv_result[151] ;
 wire \inv_result[152] ;
 wire \inv_result[153] ;
 wire \inv_result[154] ;
 wire \inv_result[155] ;
 wire \inv_result[156] ;
 wire \inv_result[157] ;
 wire \inv_result[158] ;
 wire \inv_result[159] ;
 wire \inv_result[15] ;
 wire \inv_result[160] ;
 wire \inv_result[161] ;
 wire \inv_result[162] ;
 wire \inv_result[163] ;
 wire \inv_result[164] ;
 wire \inv_result[165] ;
 wire \inv_result[166] ;
 wire \inv_result[167] ;
 wire \inv_result[168] ;
 wire \inv_result[169] ;
 wire \inv_result[16] ;
 wire \inv_result[170] ;
 wire \inv_result[171] ;
 wire \inv_result[172] ;
 wire \inv_result[173] ;
 wire \inv_result[174] ;
 wire \inv_result[175] ;
 wire \inv_result[176] ;
 wire \inv_result[177] ;
 wire \inv_result[178] ;
 wire \inv_result[179] ;
 wire \inv_result[17] ;
 wire \inv_result[180] ;
 wire \inv_result[181] ;
 wire \inv_result[182] ;
 wire \inv_result[183] ;
 wire \inv_result[184] ;
 wire \inv_result[185] ;
 wire \inv_result[186] ;
 wire \inv_result[187] ;
 wire \inv_result[188] ;
 wire \inv_result[189] ;
 wire \inv_result[18] ;
 wire \inv_result[190] ;
 wire \inv_result[191] ;
 wire \inv_result[192] ;
 wire \inv_result[193] ;
 wire \inv_result[194] ;
 wire \inv_result[195] ;
 wire \inv_result[196] ;
 wire \inv_result[197] ;
 wire \inv_result[198] ;
 wire \inv_result[199] ;
 wire \inv_result[19] ;
 wire \inv_result[1] ;
 wire \inv_result[200] ;
 wire \inv_result[201] ;
 wire \inv_result[202] ;
 wire \inv_result[203] ;
 wire \inv_result[204] ;
 wire \inv_result[205] ;
 wire \inv_result[206] ;
 wire \inv_result[207] ;
 wire \inv_result[208] ;
 wire \inv_result[209] ;
 wire \inv_result[20] ;
 wire \inv_result[210] ;
 wire \inv_result[211] ;
 wire \inv_result[212] ;
 wire \inv_result[213] ;
 wire \inv_result[214] ;
 wire \inv_result[215] ;
 wire \inv_result[216] ;
 wire \inv_result[217] ;
 wire \inv_result[218] ;
 wire \inv_result[219] ;
 wire \inv_result[21] ;
 wire \inv_result[220] ;
 wire \inv_result[221] ;
 wire \inv_result[222] ;
 wire \inv_result[223] ;
 wire \inv_result[224] ;
 wire \inv_result[225] ;
 wire \inv_result[226] ;
 wire \inv_result[227] ;
 wire \inv_result[228] ;
 wire \inv_result[229] ;
 wire \inv_result[22] ;
 wire \inv_result[230] ;
 wire \inv_result[231] ;
 wire \inv_result[232] ;
 wire \inv_result[233] ;
 wire \inv_result[234] ;
 wire \inv_result[235] ;
 wire \inv_result[236] ;
 wire \inv_result[237] ;
 wire \inv_result[238] ;
 wire \inv_result[239] ;
 wire \inv_result[23] ;
 wire \inv_result[240] ;
 wire \inv_result[241] ;
 wire \inv_result[242] ;
 wire \inv_result[243] ;
 wire \inv_result[244] ;
 wire \inv_result[245] ;
 wire \inv_result[246] ;
 wire \inv_result[247] ;
 wire \inv_result[248] ;
 wire \inv_result[249] ;
 wire \inv_result[24] ;
 wire \inv_result[250] ;
 wire \inv_result[251] ;
 wire \inv_result[252] ;
 wire \inv_result[253] ;
 wire \inv_result[254] ;
 wire \inv_result[255] ;
 wire \inv_result[25] ;
 wire \inv_result[26] ;
 wire \inv_result[27] ;
 wire \inv_result[28] ;
 wire \inv_result[29] ;
 wire \inv_result[2] ;
 wire \inv_result[30] ;
 wire \inv_result[31] ;
 wire \inv_result[32] ;
 wire \inv_result[33] ;
 wire \inv_result[34] ;
 wire \inv_result[35] ;
 wire \inv_result[36] ;
 wire \inv_result[37] ;
 wire \inv_result[38] ;
 wire \inv_result[39] ;
 wire \inv_result[3] ;
 wire \inv_result[40] ;
 wire \inv_result[41] ;
 wire \inv_result[42] ;
 wire \inv_result[43] ;
 wire \inv_result[44] ;
 wire \inv_result[45] ;
 wire \inv_result[46] ;
 wire \inv_result[47] ;
 wire \inv_result[48] ;
 wire \inv_result[49] ;
 wire \inv_result[4] ;
 wire \inv_result[50] ;
 wire \inv_result[51] ;
 wire \inv_result[52] ;
 wire \inv_result[53] ;
 wire \inv_result[54] ;
 wire \inv_result[55] ;
 wire \inv_result[56] ;
 wire \inv_result[57] ;
 wire \inv_result[58] ;
 wire \inv_result[59] ;
 wire \inv_result[5] ;
 wire \inv_result[60] ;
 wire \inv_result[61] ;
 wire \inv_result[62] ;
 wire \inv_result[63] ;
 wire \inv_result[64] ;
 wire \inv_result[65] ;
 wire \inv_result[66] ;
 wire \inv_result[67] ;
 wire \inv_result[68] ;
 wire \inv_result[69] ;
 wire \inv_result[6] ;
 wire \inv_result[70] ;
 wire \inv_result[71] ;
 wire \inv_result[72] ;
 wire \inv_result[73] ;
 wire \inv_result[74] ;
 wire \inv_result[75] ;
 wire \inv_result[76] ;
 wire \inv_result[77] ;
 wire \inv_result[78] ;
 wire \inv_result[79] ;
 wire \inv_result[7] ;
 wire \inv_result[80] ;
 wire \inv_result[81] ;
 wire \inv_result[82] ;
 wire \inv_result[83] ;
 wire \inv_result[84] ;
 wire \inv_result[85] ;
 wire \inv_result[86] ;
 wire \inv_result[87] ;
 wire \inv_result[88] ;
 wire \inv_result[89] ;
 wire \inv_result[8] ;
 wire \inv_result[90] ;
 wire \inv_result[91] ;
 wire \inv_result[92] ;
 wire \inv_result[93] ;
 wire \inv_result[94] ;
 wire \inv_result[95] ;
 wire \inv_result[96] ;
 wire \inv_result[97] ;
 wire \inv_result[98] ;
 wire \inv_result[99] ;
 wire \inv_result[9] ;
 wire next_loaded;
 wire parity_error;
 wire \perf_double[0] ;
 wire \perf_double[1] ;
 wire \perf_double[2] ;
 wire \perf_double[3] ;
 wire \perf_double[4] ;
 wire \perf_double[5] ;
 wire \perf_double[6] ;
 wire \perf_double[7] ;
 wire \perf_double[8] ;
 wire \perf_double[9] ;
 wire \perf_total[0] ;
 wire \perf_total[1] ;
 wire \perf_total[2] ;
 wire \perf_total[3] ;
 wire \perf_total[4] ;
 wire \perf_total[5] ;
 wire \perf_total[6] ;
 wire \perf_total[7] ;
 wire \perf_total[8] ;
 wire \perf_total[9] ;
 wire \perf_triple[0] ;
 wire \perf_triple[1] ;
 wire \perf_triple[2] ;
 wire \perf_triple[3] ;
 wire \perf_triple[4] ;
 wire \perf_triple[5] ;
 wire \perf_triple[6] ;
 wire \perf_triple[7] ;
 wire \perf_triple[8] ;
 wire \perf_triple[9] ;
 wire pipe_pending;
 wire rd_prev;
 wire \shift_reg[0] ;
 wire \shift_reg[100] ;
 wire \shift_reg[101] ;
 wire \shift_reg[102] ;
 wire \shift_reg[103] ;
 wire \shift_reg[104] ;
 wire \shift_reg[105] ;
 wire \shift_reg[106] ;
 wire \shift_reg[107] ;
 wire \shift_reg[108] ;
 wire \shift_reg[109] ;
 wire \shift_reg[10] ;
 wire \shift_reg[110] ;
 wire \shift_reg[111] ;
 wire \shift_reg[112] ;
 wire \shift_reg[113] ;
 wire \shift_reg[114] ;
 wire \shift_reg[115] ;
 wire \shift_reg[116] ;
 wire \shift_reg[117] ;
 wire \shift_reg[118] ;
 wire \shift_reg[119] ;
 wire \shift_reg[11] ;
 wire \shift_reg[120] ;
 wire \shift_reg[121] ;
 wire \shift_reg[122] ;
 wire \shift_reg[123] ;
 wire \shift_reg[124] ;
 wire \shift_reg[125] ;
 wire \shift_reg[126] ;
 wire \shift_reg[127] ;
 wire \shift_reg[128] ;
 wire \shift_reg[129] ;
 wire \shift_reg[12] ;
 wire \shift_reg[130] ;
 wire \shift_reg[131] ;
 wire \shift_reg[132] ;
 wire \shift_reg[133] ;
 wire \shift_reg[134] ;
 wire \shift_reg[135] ;
 wire \shift_reg[136] ;
 wire \shift_reg[137] ;
 wire \shift_reg[138] ;
 wire \shift_reg[139] ;
 wire \shift_reg[13] ;
 wire \shift_reg[140] ;
 wire \shift_reg[141] ;
 wire \shift_reg[142] ;
 wire \shift_reg[143] ;
 wire \shift_reg[144] ;
 wire \shift_reg[145] ;
 wire \shift_reg[146] ;
 wire \shift_reg[147] ;
 wire \shift_reg[148] ;
 wire \shift_reg[149] ;
 wire \shift_reg[14] ;
 wire \shift_reg[150] ;
 wire \shift_reg[151] ;
 wire \shift_reg[152] ;
 wire \shift_reg[153] ;
 wire \shift_reg[154] ;
 wire \shift_reg[155] ;
 wire \shift_reg[156] ;
 wire \shift_reg[157] ;
 wire \shift_reg[158] ;
 wire \shift_reg[159] ;
 wire \shift_reg[15] ;
 wire \shift_reg[160] ;
 wire \shift_reg[161] ;
 wire \shift_reg[162] ;
 wire \shift_reg[163] ;
 wire \shift_reg[164] ;
 wire \shift_reg[165] ;
 wire \shift_reg[166] ;
 wire \shift_reg[167] ;
 wire \shift_reg[168] ;
 wire \shift_reg[169] ;
 wire \shift_reg[16] ;
 wire \shift_reg[170] ;
 wire \shift_reg[171] ;
 wire \shift_reg[172] ;
 wire \shift_reg[173] ;
 wire \shift_reg[174] ;
 wire \shift_reg[175] ;
 wire \shift_reg[176] ;
 wire \shift_reg[177] ;
 wire \shift_reg[178] ;
 wire \shift_reg[179] ;
 wire \shift_reg[17] ;
 wire \shift_reg[180] ;
 wire \shift_reg[181] ;
 wire \shift_reg[182] ;
 wire \shift_reg[183] ;
 wire \shift_reg[184] ;
 wire \shift_reg[185] ;
 wire \shift_reg[186] ;
 wire \shift_reg[187] ;
 wire \shift_reg[188] ;
 wire \shift_reg[189] ;
 wire \shift_reg[18] ;
 wire \shift_reg[190] ;
 wire \shift_reg[191] ;
 wire \shift_reg[192] ;
 wire \shift_reg[193] ;
 wire \shift_reg[194] ;
 wire \shift_reg[195] ;
 wire \shift_reg[196] ;
 wire \shift_reg[197] ;
 wire \shift_reg[198] ;
 wire \shift_reg[199] ;
 wire \shift_reg[19] ;
 wire \shift_reg[1] ;
 wire \shift_reg[200] ;
 wire \shift_reg[201] ;
 wire \shift_reg[202] ;
 wire \shift_reg[203] ;
 wire \shift_reg[204] ;
 wire \shift_reg[205] ;
 wire \shift_reg[206] ;
 wire \shift_reg[207] ;
 wire \shift_reg[208] ;
 wire \shift_reg[209] ;
 wire \shift_reg[20] ;
 wire \shift_reg[210] ;
 wire \shift_reg[211] ;
 wire \shift_reg[212] ;
 wire \shift_reg[213] ;
 wire \shift_reg[214] ;
 wire \shift_reg[215] ;
 wire \shift_reg[216] ;
 wire \shift_reg[217] ;
 wire \shift_reg[218] ;
 wire \shift_reg[219] ;
 wire \shift_reg[21] ;
 wire \shift_reg[220] ;
 wire \shift_reg[221] ;
 wire \shift_reg[222] ;
 wire \shift_reg[223] ;
 wire \shift_reg[224] ;
 wire \shift_reg[225] ;
 wire \shift_reg[226] ;
 wire \shift_reg[227] ;
 wire \shift_reg[228] ;
 wire \shift_reg[229] ;
 wire \shift_reg[22] ;
 wire \shift_reg[230] ;
 wire \shift_reg[231] ;
 wire \shift_reg[232] ;
 wire \shift_reg[233] ;
 wire \shift_reg[234] ;
 wire \shift_reg[235] ;
 wire \shift_reg[236] ;
 wire \shift_reg[237] ;
 wire \shift_reg[238] ;
 wire \shift_reg[239] ;
 wire \shift_reg[23] ;
 wire \shift_reg[240] ;
 wire \shift_reg[241] ;
 wire \shift_reg[242] ;
 wire \shift_reg[243] ;
 wire \shift_reg[244] ;
 wire \shift_reg[245] ;
 wire \shift_reg[246] ;
 wire \shift_reg[247] ;
 wire \shift_reg[248] ;
 wire \shift_reg[249] ;
 wire \shift_reg[24] ;
 wire \shift_reg[250] ;
 wire \shift_reg[251] ;
 wire \shift_reg[252] ;
 wire \shift_reg[253] ;
 wire \shift_reg[254] ;
 wire \shift_reg[255] ;
 wire \shift_reg[256] ;
 wire \shift_reg[257] ;
 wire \shift_reg[258] ;
 wire \shift_reg[259] ;
 wire \shift_reg[25] ;
 wire \shift_reg[260] ;
 wire \shift_reg[261] ;
 wire \shift_reg[262] ;
 wire \shift_reg[263] ;
 wire \shift_reg[264] ;
 wire \shift_reg[265] ;
 wire \shift_reg[266] ;
 wire \shift_reg[267] ;
 wire \shift_reg[268] ;
 wire \shift_reg[269] ;
 wire \shift_reg[26] ;
 wire \shift_reg[270] ;
 wire \shift_reg[271] ;
 wire \shift_reg[27] ;
 wire \shift_reg[28] ;
 wire \shift_reg[29] ;
 wire \shift_reg[2] ;
 wire \shift_reg[30] ;
 wire \shift_reg[31] ;
 wire \shift_reg[32] ;
 wire \shift_reg[33] ;
 wire \shift_reg[34] ;
 wire \shift_reg[35] ;
 wire \shift_reg[36] ;
 wire \shift_reg[37] ;
 wire \shift_reg[38] ;
 wire \shift_reg[39] ;
 wire \shift_reg[3] ;
 wire \shift_reg[40] ;
 wire \shift_reg[41] ;
 wire \shift_reg[42] ;
 wire \shift_reg[43] ;
 wire \shift_reg[44] ;
 wire \shift_reg[45] ;
 wire \shift_reg[46] ;
 wire \shift_reg[47] ;
 wire \shift_reg[48] ;
 wire \shift_reg[49] ;
 wire \shift_reg[4] ;
 wire \shift_reg[50] ;
 wire \shift_reg[51] ;
 wire \shift_reg[52] ;
 wire \shift_reg[53] ;
 wire \shift_reg[54] ;
 wire \shift_reg[55] ;
 wire \shift_reg[56] ;
 wire \shift_reg[57] ;
 wire \shift_reg[58] ;
 wire \shift_reg[59] ;
 wire \shift_reg[5] ;
 wire \shift_reg[60] ;
 wire \shift_reg[61] ;
 wire \shift_reg[62] ;
 wire \shift_reg[63] ;
 wire \shift_reg[64] ;
 wire \shift_reg[65] ;
 wire \shift_reg[66] ;
 wire \shift_reg[67] ;
 wire \shift_reg[68] ;
 wire \shift_reg[69] ;
 wire \shift_reg[6] ;
 wire \shift_reg[70] ;
 wire \shift_reg[71] ;
 wire \shift_reg[72] ;
 wire \shift_reg[73] ;
 wire \shift_reg[74] ;
 wire \shift_reg[75] ;
 wire \shift_reg[76] ;
 wire \shift_reg[77] ;
 wire \shift_reg[78] ;
 wire \shift_reg[79] ;
 wire \shift_reg[7] ;
 wire \shift_reg[80] ;
 wire \shift_reg[81] ;
 wire \shift_reg[82] ;
 wire \shift_reg[83] ;
 wire \shift_reg[84] ;
 wire \shift_reg[85] ;
 wire \shift_reg[86] ;
 wire \shift_reg[87] ;
 wire \shift_reg[88] ;
 wire \shift_reg[89] ;
 wire \shift_reg[8] ;
 wire \shift_reg[90] ;
 wire \shift_reg[91] ;
 wire \shift_reg[92] ;
 wire \shift_reg[93] ;
 wire \shift_reg[94] ;
 wire \shift_reg[95] ;
 wire \shift_reg[96] ;
 wire \shift_reg[97] ;
 wire \shift_reg[98] ;
 wire \shift_reg[99] ;
 wire \shift_reg[9] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \trng_data[0] ;
 wire \trng_data[1] ;
 wire \trng_data[2] ;
 wire \trng_data[3] ;
 wire \trng_data[4] ;
 wire \trng_data[5] ;
 wire \trng_data[6] ;
 wire \trng_data[7] ;
 wire trng_ready;
 wire \u_inv.counter[0] ;
 wire \u_inv.counter[1] ;
 wire \u_inv.counter[2] ;
 wire \u_inv.counter[3] ;
 wire \u_inv.counter[4] ;
 wire \u_inv.counter[5] ;
 wire \u_inv.counter[6] ;
 wire \u_inv.counter[7] ;
 wire \u_inv.counter[8] ;
 wire \u_inv.counter[9] ;
 wire \u_inv.d_next[0] ;
 wire \u_inv.d_next[100] ;
 wire \u_inv.d_next[101] ;
 wire \u_inv.d_next[102] ;
 wire \u_inv.d_next[103] ;
 wire \u_inv.d_next[104] ;
 wire \u_inv.d_next[105] ;
 wire \u_inv.d_next[106] ;
 wire \u_inv.d_next[107] ;
 wire \u_inv.d_next[108] ;
 wire \u_inv.d_next[109] ;
 wire \u_inv.d_next[10] ;
 wire \u_inv.d_next[110] ;
 wire \u_inv.d_next[111] ;
 wire \u_inv.d_next[112] ;
 wire \u_inv.d_next[113] ;
 wire \u_inv.d_next[114] ;
 wire \u_inv.d_next[115] ;
 wire \u_inv.d_next[116] ;
 wire \u_inv.d_next[117] ;
 wire \u_inv.d_next[118] ;
 wire \u_inv.d_next[119] ;
 wire \u_inv.d_next[11] ;
 wire \u_inv.d_next[120] ;
 wire \u_inv.d_next[121] ;
 wire \u_inv.d_next[122] ;
 wire \u_inv.d_next[123] ;
 wire \u_inv.d_next[124] ;
 wire \u_inv.d_next[125] ;
 wire \u_inv.d_next[126] ;
 wire \u_inv.d_next[127] ;
 wire \u_inv.d_next[128] ;
 wire \u_inv.d_next[129] ;
 wire \u_inv.d_next[12] ;
 wire \u_inv.d_next[130] ;
 wire \u_inv.d_next[131] ;
 wire \u_inv.d_next[132] ;
 wire \u_inv.d_next[133] ;
 wire \u_inv.d_next[134] ;
 wire \u_inv.d_next[135] ;
 wire \u_inv.d_next[136] ;
 wire \u_inv.d_next[137] ;
 wire \u_inv.d_next[138] ;
 wire \u_inv.d_next[139] ;
 wire \u_inv.d_next[13] ;
 wire \u_inv.d_next[140] ;
 wire \u_inv.d_next[141] ;
 wire \u_inv.d_next[142] ;
 wire \u_inv.d_next[143] ;
 wire \u_inv.d_next[144] ;
 wire \u_inv.d_next[145] ;
 wire \u_inv.d_next[146] ;
 wire \u_inv.d_next[147] ;
 wire \u_inv.d_next[148] ;
 wire \u_inv.d_next[149] ;
 wire \u_inv.d_next[14] ;
 wire \u_inv.d_next[150] ;
 wire \u_inv.d_next[151] ;
 wire \u_inv.d_next[152] ;
 wire \u_inv.d_next[153] ;
 wire \u_inv.d_next[154] ;
 wire \u_inv.d_next[155] ;
 wire \u_inv.d_next[156] ;
 wire \u_inv.d_next[157] ;
 wire \u_inv.d_next[158] ;
 wire \u_inv.d_next[159] ;
 wire \u_inv.d_next[15] ;
 wire \u_inv.d_next[160] ;
 wire \u_inv.d_next[161] ;
 wire \u_inv.d_next[162] ;
 wire \u_inv.d_next[163] ;
 wire \u_inv.d_next[164] ;
 wire \u_inv.d_next[165] ;
 wire \u_inv.d_next[166] ;
 wire \u_inv.d_next[167] ;
 wire \u_inv.d_next[168] ;
 wire \u_inv.d_next[169] ;
 wire \u_inv.d_next[16] ;
 wire \u_inv.d_next[170] ;
 wire \u_inv.d_next[171] ;
 wire \u_inv.d_next[172] ;
 wire \u_inv.d_next[173] ;
 wire \u_inv.d_next[174] ;
 wire \u_inv.d_next[175] ;
 wire \u_inv.d_next[176] ;
 wire \u_inv.d_next[177] ;
 wire \u_inv.d_next[178] ;
 wire \u_inv.d_next[179] ;
 wire \u_inv.d_next[17] ;
 wire \u_inv.d_next[180] ;
 wire \u_inv.d_next[181] ;
 wire \u_inv.d_next[182] ;
 wire \u_inv.d_next[183] ;
 wire \u_inv.d_next[184] ;
 wire \u_inv.d_next[185] ;
 wire \u_inv.d_next[186] ;
 wire \u_inv.d_next[187] ;
 wire \u_inv.d_next[188] ;
 wire \u_inv.d_next[189] ;
 wire \u_inv.d_next[18] ;
 wire \u_inv.d_next[190] ;
 wire \u_inv.d_next[191] ;
 wire \u_inv.d_next[192] ;
 wire \u_inv.d_next[193] ;
 wire \u_inv.d_next[194] ;
 wire \u_inv.d_next[195] ;
 wire \u_inv.d_next[196] ;
 wire \u_inv.d_next[197] ;
 wire \u_inv.d_next[198] ;
 wire \u_inv.d_next[199] ;
 wire \u_inv.d_next[19] ;
 wire \u_inv.d_next[1] ;
 wire \u_inv.d_next[200] ;
 wire \u_inv.d_next[201] ;
 wire \u_inv.d_next[202] ;
 wire \u_inv.d_next[203] ;
 wire \u_inv.d_next[204] ;
 wire \u_inv.d_next[205] ;
 wire \u_inv.d_next[206] ;
 wire \u_inv.d_next[207] ;
 wire \u_inv.d_next[208] ;
 wire \u_inv.d_next[209] ;
 wire \u_inv.d_next[20] ;
 wire \u_inv.d_next[210] ;
 wire \u_inv.d_next[211] ;
 wire \u_inv.d_next[212] ;
 wire \u_inv.d_next[213] ;
 wire \u_inv.d_next[214] ;
 wire \u_inv.d_next[215] ;
 wire \u_inv.d_next[216] ;
 wire \u_inv.d_next[217] ;
 wire \u_inv.d_next[218] ;
 wire \u_inv.d_next[219] ;
 wire \u_inv.d_next[21] ;
 wire \u_inv.d_next[220] ;
 wire \u_inv.d_next[221] ;
 wire \u_inv.d_next[222] ;
 wire \u_inv.d_next[223] ;
 wire \u_inv.d_next[224] ;
 wire \u_inv.d_next[225] ;
 wire \u_inv.d_next[226] ;
 wire \u_inv.d_next[227] ;
 wire \u_inv.d_next[228] ;
 wire \u_inv.d_next[229] ;
 wire \u_inv.d_next[22] ;
 wire \u_inv.d_next[230] ;
 wire \u_inv.d_next[231] ;
 wire \u_inv.d_next[232] ;
 wire \u_inv.d_next[233] ;
 wire \u_inv.d_next[234] ;
 wire \u_inv.d_next[235] ;
 wire \u_inv.d_next[236] ;
 wire \u_inv.d_next[237] ;
 wire \u_inv.d_next[238] ;
 wire \u_inv.d_next[239] ;
 wire \u_inv.d_next[23] ;
 wire \u_inv.d_next[240] ;
 wire \u_inv.d_next[241] ;
 wire \u_inv.d_next[242] ;
 wire \u_inv.d_next[243] ;
 wire \u_inv.d_next[244] ;
 wire \u_inv.d_next[245] ;
 wire \u_inv.d_next[246] ;
 wire \u_inv.d_next[247] ;
 wire \u_inv.d_next[248] ;
 wire \u_inv.d_next[249] ;
 wire \u_inv.d_next[24] ;
 wire \u_inv.d_next[250] ;
 wire \u_inv.d_next[251] ;
 wire \u_inv.d_next[252] ;
 wire \u_inv.d_next[253] ;
 wire \u_inv.d_next[254] ;
 wire \u_inv.d_next[255] ;
 wire \u_inv.d_next[256] ;
 wire \u_inv.d_next[25] ;
 wire \u_inv.d_next[26] ;
 wire \u_inv.d_next[27] ;
 wire \u_inv.d_next[28] ;
 wire \u_inv.d_next[29] ;
 wire \u_inv.d_next[2] ;
 wire \u_inv.d_next[30] ;
 wire \u_inv.d_next[31] ;
 wire \u_inv.d_next[32] ;
 wire \u_inv.d_next[33] ;
 wire \u_inv.d_next[34] ;
 wire \u_inv.d_next[35] ;
 wire \u_inv.d_next[36] ;
 wire \u_inv.d_next[37] ;
 wire \u_inv.d_next[38] ;
 wire \u_inv.d_next[39] ;
 wire \u_inv.d_next[3] ;
 wire \u_inv.d_next[40] ;
 wire \u_inv.d_next[41] ;
 wire \u_inv.d_next[42] ;
 wire \u_inv.d_next[43] ;
 wire \u_inv.d_next[44] ;
 wire \u_inv.d_next[45] ;
 wire \u_inv.d_next[46] ;
 wire \u_inv.d_next[47] ;
 wire \u_inv.d_next[48] ;
 wire \u_inv.d_next[49] ;
 wire \u_inv.d_next[4] ;
 wire \u_inv.d_next[50] ;
 wire \u_inv.d_next[51] ;
 wire \u_inv.d_next[52] ;
 wire \u_inv.d_next[53] ;
 wire \u_inv.d_next[54] ;
 wire \u_inv.d_next[55] ;
 wire \u_inv.d_next[56] ;
 wire \u_inv.d_next[57] ;
 wire \u_inv.d_next[58] ;
 wire \u_inv.d_next[59] ;
 wire \u_inv.d_next[5] ;
 wire \u_inv.d_next[60] ;
 wire \u_inv.d_next[61] ;
 wire \u_inv.d_next[62] ;
 wire \u_inv.d_next[63] ;
 wire \u_inv.d_next[64] ;
 wire \u_inv.d_next[65] ;
 wire \u_inv.d_next[66] ;
 wire \u_inv.d_next[67] ;
 wire \u_inv.d_next[68] ;
 wire \u_inv.d_next[69] ;
 wire \u_inv.d_next[6] ;
 wire \u_inv.d_next[70] ;
 wire \u_inv.d_next[71] ;
 wire \u_inv.d_next[72] ;
 wire \u_inv.d_next[73] ;
 wire \u_inv.d_next[74] ;
 wire \u_inv.d_next[75] ;
 wire \u_inv.d_next[76] ;
 wire \u_inv.d_next[77] ;
 wire \u_inv.d_next[78] ;
 wire \u_inv.d_next[79] ;
 wire \u_inv.d_next[7] ;
 wire \u_inv.d_next[80] ;
 wire \u_inv.d_next[81] ;
 wire \u_inv.d_next[82] ;
 wire \u_inv.d_next[83] ;
 wire \u_inv.d_next[84] ;
 wire \u_inv.d_next[85] ;
 wire \u_inv.d_next[86] ;
 wire \u_inv.d_next[87] ;
 wire \u_inv.d_next[88] ;
 wire \u_inv.d_next[89] ;
 wire \u_inv.d_next[8] ;
 wire \u_inv.d_next[90] ;
 wire \u_inv.d_next[91] ;
 wire \u_inv.d_next[92] ;
 wire \u_inv.d_next[93] ;
 wire \u_inv.d_next[94] ;
 wire \u_inv.d_next[95] ;
 wire \u_inv.d_next[96] ;
 wire \u_inv.d_next[97] ;
 wire \u_inv.d_next[98] ;
 wire \u_inv.d_next[99] ;
 wire \u_inv.d_next[9] ;
 wire \u_inv.d_reg[0] ;
 wire \u_inv.d_reg[100] ;
 wire \u_inv.d_reg[101] ;
 wire \u_inv.d_reg[102] ;
 wire \u_inv.d_reg[103] ;
 wire \u_inv.d_reg[104] ;
 wire \u_inv.d_reg[105] ;
 wire \u_inv.d_reg[106] ;
 wire \u_inv.d_reg[107] ;
 wire \u_inv.d_reg[108] ;
 wire \u_inv.d_reg[109] ;
 wire \u_inv.d_reg[10] ;
 wire \u_inv.d_reg[110] ;
 wire \u_inv.d_reg[111] ;
 wire \u_inv.d_reg[112] ;
 wire \u_inv.d_reg[113] ;
 wire \u_inv.d_reg[114] ;
 wire \u_inv.d_reg[115] ;
 wire \u_inv.d_reg[116] ;
 wire \u_inv.d_reg[117] ;
 wire \u_inv.d_reg[118] ;
 wire \u_inv.d_reg[119] ;
 wire \u_inv.d_reg[11] ;
 wire \u_inv.d_reg[120] ;
 wire \u_inv.d_reg[121] ;
 wire \u_inv.d_reg[122] ;
 wire \u_inv.d_reg[123] ;
 wire \u_inv.d_reg[124] ;
 wire \u_inv.d_reg[125] ;
 wire \u_inv.d_reg[126] ;
 wire \u_inv.d_reg[127] ;
 wire \u_inv.d_reg[128] ;
 wire \u_inv.d_reg[129] ;
 wire \u_inv.d_reg[12] ;
 wire \u_inv.d_reg[130] ;
 wire \u_inv.d_reg[131] ;
 wire \u_inv.d_reg[132] ;
 wire \u_inv.d_reg[133] ;
 wire \u_inv.d_reg[134] ;
 wire \u_inv.d_reg[135] ;
 wire \u_inv.d_reg[136] ;
 wire \u_inv.d_reg[137] ;
 wire \u_inv.d_reg[138] ;
 wire \u_inv.d_reg[139] ;
 wire \u_inv.d_reg[13] ;
 wire \u_inv.d_reg[140] ;
 wire \u_inv.d_reg[141] ;
 wire \u_inv.d_reg[142] ;
 wire \u_inv.d_reg[143] ;
 wire \u_inv.d_reg[144] ;
 wire \u_inv.d_reg[145] ;
 wire \u_inv.d_reg[146] ;
 wire \u_inv.d_reg[147] ;
 wire \u_inv.d_reg[148] ;
 wire \u_inv.d_reg[149] ;
 wire \u_inv.d_reg[14] ;
 wire \u_inv.d_reg[150] ;
 wire \u_inv.d_reg[151] ;
 wire \u_inv.d_reg[152] ;
 wire \u_inv.d_reg[153] ;
 wire \u_inv.d_reg[154] ;
 wire \u_inv.d_reg[155] ;
 wire \u_inv.d_reg[156] ;
 wire \u_inv.d_reg[157] ;
 wire \u_inv.d_reg[158] ;
 wire \u_inv.d_reg[159] ;
 wire \u_inv.d_reg[15] ;
 wire \u_inv.d_reg[160] ;
 wire \u_inv.d_reg[161] ;
 wire \u_inv.d_reg[162] ;
 wire \u_inv.d_reg[163] ;
 wire \u_inv.d_reg[164] ;
 wire \u_inv.d_reg[165] ;
 wire \u_inv.d_reg[166] ;
 wire \u_inv.d_reg[167] ;
 wire \u_inv.d_reg[168] ;
 wire \u_inv.d_reg[169] ;
 wire \u_inv.d_reg[16] ;
 wire \u_inv.d_reg[170] ;
 wire \u_inv.d_reg[171] ;
 wire \u_inv.d_reg[172] ;
 wire \u_inv.d_reg[173] ;
 wire \u_inv.d_reg[174] ;
 wire \u_inv.d_reg[175] ;
 wire \u_inv.d_reg[176] ;
 wire \u_inv.d_reg[177] ;
 wire \u_inv.d_reg[178] ;
 wire \u_inv.d_reg[179] ;
 wire \u_inv.d_reg[17] ;
 wire \u_inv.d_reg[180] ;
 wire \u_inv.d_reg[181] ;
 wire \u_inv.d_reg[182] ;
 wire \u_inv.d_reg[183] ;
 wire \u_inv.d_reg[184] ;
 wire \u_inv.d_reg[185] ;
 wire \u_inv.d_reg[186] ;
 wire \u_inv.d_reg[187] ;
 wire \u_inv.d_reg[188] ;
 wire \u_inv.d_reg[189] ;
 wire \u_inv.d_reg[18] ;
 wire \u_inv.d_reg[190] ;
 wire \u_inv.d_reg[191] ;
 wire \u_inv.d_reg[192] ;
 wire \u_inv.d_reg[193] ;
 wire \u_inv.d_reg[194] ;
 wire \u_inv.d_reg[195] ;
 wire \u_inv.d_reg[196] ;
 wire \u_inv.d_reg[197] ;
 wire \u_inv.d_reg[198] ;
 wire \u_inv.d_reg[199] ;
 wire \u_inv.d_reg[19] ;
 wire \u_inv.d_reg[1] ;
 wire \u_inv.d_reg[200] ;
 wire \u_inv.d_reg[201] ;
 wire \u_inv.d_reg[202] ;
 wire \u_inv.d_reg[203] ;
 wire \u_inv.d_reg[204] ;
 wire \u_inv.d_reg[205] ;
 wire \u_inv.d_reg[206] ;
 wire \u_inv.d_reg[207] ;
 wire \u_inv.d_reg[208] ;
 wire \u_inv.d_reg[209] ;
 wire \u_inv.d_reg[20] ;
 wire \u_inv.d_reg[210] ;
 wire \u_inv.d_reg[211] ;
 wire \u_inv.d_reg[212] ;
 wire \u_inv.d_reg[213] ;
 wire \u_inv.d_reg[214] ;
 wire \u_inv.d_reg[215] ;
 wire \u_inv.d_reg[216] ;
 wire \u_inv.d_reg[217] ;
 wire \u_inv.d_reg[218] ;
 wire \u_inv.d_reg[219] ;
 wire \u_inv.d_reg[21] ;
 wire \u_inv.d_reg[220] ;
 wire \u_inv.d_reg[221] ;
 wire \u_inv.d_reg[222] ;
 wire \u_inv.d_reg[223] ;
 wire \u_inv.d_reg[224] ;
 wire \u_inv.d_reg[225] ;
 wire \u_inv.d_reg[226] ;
 wire \u_inv.d_reg[227] ;
 wire \u_inv.d_reg[228] ;
 wire \u_inv.d_reg[229] ;
 wire \u_inv.d_reg[22] ;
 wire \u_inv.d_reg[230] ;
 wire \u_inv.d_reg[231] ;
 wire \u_inv.d_reg[232] ;
 wire \u_inv.d_reg[233] ;
 wire \u_inv.d_reg[234] ;
 wire \u_inv.d_reg[235] ;
 wire \u_inv.d_reg[236] ;
 wire \u_inv.d_reg[237] ;
 wire \u_inv.d_reg[238] ;
 wire \u_inv.d_reg[239] ;
 wire \u_inv.d_reg[23] ;
 wire \u_inv.d_reg[240] ;
 wire \u_inv.d_reg[241] ;
 wire \u_inv.d_reg[242] ;
 wire \u_inv.d_reg[243] ;
 wire \u_inv.d_reg[244] ;
 wire \u_inv.d_reg[245] ;
 wire \u_inv.d_reg[246] ;
 wire \u_inv.d_reg[247] ;
 wire \u_inv.d_reg[248] ;
 wire \u_inv.d_reg[249] ;
 wire \u_inv.d_reg[24] ;
 wire \u_inv.d_reg[250] ;
 wire \u_inv.d_reg[251] ;
 wire \u_inv.d_reg[252] ;
 wire \u_inv.d_reg[253] ;
 wire \u_inv.d_reg[254] ;
 wire \u_inv.d_reg[255] ;
 wire \u_inv.d_reg[256] ;
 wire \u_inv.d_reg[25] ;
 wire \u_inv.d_reg[26] ;
 wire \u_inv.d_reg[27] ;
 wire \u_inv.d_reg[28] ;
 wire \u_inv.d_reg[29] ;
 wire \u_inv.d_reg[2] ;
 wire \u_inv.d_reg[30] ;
 wire \u_inv.d_reg[31] ;
 wire \u_inv.d_reg[32] ;
 wire \u_inv.d_reg[33] ;
 wire \u_inv.d_reg[34] ;
 wire \u_inv.d_reg[35] ;
 wire \u_inv.d_reg[36] ;
 wire \u_inv.d_reg[37] ;
 wire \u_inv.d_reg[38] ;
 wire \u_inv.d_reg[39] ;
 wire \u_inv.d_reg[3] ;
 wire \u_inv.d_reg[40] ;
 wire \u_inv.d_reg[41] ;
 wire \u_inv.d_reg[42] ;
 wire \u_inv.d_reg[43] ;
 wire \u_inv.d_reg[44] ;
 wire \u_inv.d_reg[45] ;
 wire \u_inv.d_reg[46] ;
 wire \u_inv.d_reg[47] ;
 wire \u_inv.d_reg[48] ;
 wire \u_inv.d_reg[49] ;
 wire \u_inv.d_reg[4] ;
 wire \u_inv.d_reg[50] ;
 wire \u_inv.d_reg[51] ;
 wire \u_inv.d_reg[52] ;
 wire \u_inv.d_reg[53] ;
 wire \u_inv.d_reg[54] ;
 wire \u_inv.d_reg[55] ;
 wire \u_inv.d_reg[56] ;
 wire \u_inv.d_reg[57] ;
 wire \u_inv.d_reg[58] ;
 wire \u_inv.d_reg[59] ;
 wire \u_inv.d_reg[5] ;
 wire \u_inv.d_reg[60] ;
 wire \u_inv.d_reg[61] ;
 wire \u_inv.d_reg[62] ;
 wire \u_inv.d_reg[63] ;
 wire \u_inv.d_reg[64] ;
 wire \u_inv.d_reg[65] ;
 wire \u_inv.d_reg[66] ;
 wire \u_inv.d_reg[67] ;
 wire \u_inv.d_reg[68] ;
 wire \u_inv.d_reg[69] ;
 wire \u_inv.d_reg[6] ;
 wire \u_inv.d_reg[70] ;
 wire \u_inv.d_reg[71] ;
 wire \u_inv.d_reg[72] ;
 wire \u_inv.d_reg[73] ;
 wire \u_inv.d_reg[74] ;
 wire \u_inv.d_reg[75] ;
 wire \u_inv.d_reg[76] ;
 wire \u_inv.d_reg[77] ;
 wire \u_inv.d_reg[78] ;
 wire \u_inv.d_reg[79] ;
 wire \u_inv.d_reg[7] ;
 wire \u_inv.d_reg[80] ;
 wire \u_inv.d_reg[81] ;
 wire \u_inv.d_reg[82] ;
 wire \u_inv.d_reg[83] ;
 wire \u_inv.d_reg[84] ;
 wire \u_inv.d_reg[85] ;
 wire \u_inv.d_reg[86] ;
 wire \u_inv.d_reg[87] ;
 wire \u_inv.d_reg[88] ;
 wire \u_inv.d_reg[89] ;
 wire \u_inv.d_reg[8] ;
 wire \u_inv.d_reg[90] ;
 wire \u_inv.d_reg[91] ;
 wire \u_inv.d_reg[92] ;
 wire \u_inv.d_reg[93] ;
 wire \u_inv.d_reg[94] ;
 wire \u_inv.d_reg[95] ;
 wire \u_inv.d_reg[96] ;
 wire \u_inv.d_reg[97] ;
 wire \u_inv.d_reg[98] ;
 wire \u_inv.d_reg[99] ;
 wire \u_inv.d_reg[9] ;
 wire \u_inv.delta_double[0] ;
 wire \u_inv.delta_reg[1] ;
 wire \u_inv.delta_reg[2] ;
 wire \u_inv.delta_reg[3] ;
 wire \u_inv.delta_reg[4] ;
 wire \u_inv.delta_reg[5] ;
 wire \u_inv.delta_reg[6] ;
 wire \u_inv.delta_reg[7] ;
 wire \u_inv.delta_reg[8] ;
 wire \u_inv.delta_reg[9] ;
 wire \u_inv.f_next[0] ;
 wire \u_inv.f_next[100] ;
 wire \u_inv.f_next[101] ;
 wire \u_inv.f_next[102] ;
 wire \u_inv.f_next[103] ;
 wire \u_inv.f_next[104] ;
 wire \u_inv.f_next[105] ;
 wire \u_inv.f_next[106] ;
 wire \u_inv.f_next[107] ;
 wire \u_inv.f_next[108] ;
 wire \u_inv.f_next[109] ;
 wire \u_inv.f_next[10] ;
 wire \u_inv.f_next[110] ;
 wire \u_inv.f_next[111] ;
 wire \u_inv.f_next[112] ;
 wire \u_inv.f_next[113] ;
 wire \u_inv.f_next[114] ;
 wire \u_inv.f_next[115] ;
 wire \u_inv.f_next[116] ;
 wire \u_inv.f_next[117] ;
 wire \u_inv.f_next[118] ;
 wire \u_inv.f_next[119] ;
 wire \u_inv.f_next[11] ;
 wire \u_inv.f_next[120] ;
 wire \u_inv.f_next[121] ;
 wire \u_inv.f_next[122] ;
 wire \u_inv.f_next[123] ;
 wire \u_inv.f_next[124] ;
 wire \u_inv.f_next[125] ;
 wire \u_inv.f_next[126] ;
 wire \u_inv.f_next[127] ;
 wire \u_inv.f_next[128] ;
 wire \u_inv.f_next[129] ;
 wire \u_inv.f_next[12] ;
 wire \u_inv.f_next[130] ;
 wire \u_inv.f_next[131] ;
 wire \u_inv.f_next[132] ;
 wire \u_inv.f_next[133] ;
 wire \u_inv.f_next[134] ;
 wire \u_inv.f_next[135] ;
 wire \u_inv.f_next[136] ;
 wire \u_inv.f_next[137] ;
 wire \u_inv.f_next[138] ;
 wire \u_inv.f_next[139] ;
 wire \u_inv.f_next[13] ;
 wire \u_inv.f_next[140] ;
 wire \u_inv.f_next[141] ;
 wire \u_inv.f_next[142] ;
 wire \u_inv.f_next[143] ;
 wire \u_inv.f_next[144] ;
 wire \u_inv.f_next[145] ;
 wire \u_inv.f_next[146] ;
 wire \u_inv.f_next[147] ;
 wire \u_inv.f_next[148] ;
 wire \u_inv.f_next[149] ;
 wire \u_inv.f_next[14] ;
 wire \u_inv.f_next[150] ;
 wire \u_inv.f_next[151] ;
 wire \u_inv.f_next[152] ;
 wire \u_inv.f_next[153] ;
 wire \u_inv.f_next[154] ;
 wire \u_inv.f_next[155] ;
 wire \u_inv.f_next[156] ;
 wire \u_inv.f_next[157] ;
 wire \u_inv.f_next[158] ;
 wire \u_inv.f_next[159] ;
 wire \u_inv.f_next[15] ;
 wire \u_inv.f_next[160] ;
 wire \u_inv.f_next[161] ;
 wire \u_inv.f_next[162] ;
 wire \u_inv.f_next[163] ;
 wire \u_inv.f_next[164] ;
 wire \u_inv.f_next[165] ;
 wire \u_inv.f_next[166] ;
 wire \u_inv.f_next[167] ;
 wire \u_inv.f_next[168] ;
 wire \u_inv.f_next[169] ;
 wire \u_inv.f_next[16] ;
 wire \u_inv.f_next[170] ;
 wire \u_inv.f_next[171] ;
 wire \u_inv.f_next[172] ;
 wire \u_inv.f_next[173] ;
 wire \u_inv.f_next[174] ;
 wire \u_inv.f_next[175] ;
 wire \u_inv.f_next[176] ;
 wire \u_inv.f_next[177] ;
 wire \u_inv.f_next[178] ;
 wire \u_inv.f_next[179] ;
 wire \u_inv.f_next[17] ;
 wire \u_inv.f_next[180] ;
 wire \u_inv.f_next[181] ;
 wire \u_inv.f_next[182] ;
 wire \u_inv.f_next[183] ;
 wire \u_inv.f_next[184] ;
 wire \u_inv.f_next[185] ;
 wire \u_inv.f_next[186] ;
 wire \u_inv.f_next[187] ;
 wire \u_inv.f_next[188] ;
 wire \u_inv.f_next[189] ;
 wire \u_inv.f_next[18] ;
 wire \u_inv.f_next[190] ;
 wire \u_inv.f_next[191] ;
 wire \u_inv.f_next[192] ;
 wire \u_inv.f_next[193] ;
 wire \u_inv.f_next[194] ;
 wire \u_inv.f_next[195] ;
 wire \u_inv.f_next[196] ;
 wire \u_inv.f_next[197] ;
 wire \u_inv.f_next[198] ;
 wire \u_inv.f_next[199] ;
 wire \u_inv.f_next[19] ;
 wire \u_inv.f_next[1] ;
 wire \u_inv.f_next[200] ;
 wire \u_inv.f_next[201] ;
 wire \u_inv.f_next[202] ;
 wire \u_inv.f_next[203] ;
 wire \u_inv.f_next[204] ;
 wire \u_inv.f_next[205] ;
 wire \u_inv.f_next[206] ;
 wire \u_inv.f_next[207] ;
 wire \u_inv.f_next[208] ;
 wire \u_inv.f_next[209] ;
 wire \u_inv.f_next[20] ;
 wire \u_inv.f_next[210] ;
 wire \u_inv.f_next[211] ;
 wire \u_inv.f_next[212] ;
 wire \u_inv.f_next[213] ;
 wire \u_inv.f_next[214] ;
 wire \u_inv.f_next[215] ;
 wire \u_inv.f_next[216] ;
 wire \u_inv.f_next[217] ;
 wire \u_inv.f_next[218] ;
 wire \u_inv.f_next[219] ;
 wire \u_inv.f_next[21] ;
 wire \u_inv.f_next[220] ;
 wire \u_inv.f_next[221] ;
 wire \u_inv.f_next[222] ;
 wire \u_inv.f_next[223] ;
 wire \u_inv.f_next[224] ;
 wire \u_inv.f_next[225] ;
 wire \u_inv.f_next[226] ;
 wire \u_inv.f_next[227] ;
 wire \u_inv.f_next[228] ;
 wire \u_inv.f_next[229] ;
 wire \u_inv.f_next[22] ;
 wire \u_inv.f_next[230] ;
 wire \u_inv.f_next[231] ;
 wire \u_inv.f_next[232] ;
 wire \u_inv.f_next[233] ;
 wire \u_inv.f_next[234] ;
 wire \u_inv.f_next[235] ;
 wire \u_inv.f_next[236] ;
 wire \u_inv.f_next[237] ;
 wire \u_inv.f_next[238] ;
 wire \u_inv.f_next[239] ;
 wire \u_inv.f_next[23] ;
 wire \u_inv.f_next[240] ;
 wire \u_inv.f_next[241] ;
 wire \u_inv.f_next[242] ;
 wire \u_inv.f_next[243] ;
 wire \u_inv.f_next[244] ;
 wire \u_inv.f_next[245] ;
 wire \u_inv.f_next[246] ;
 wire \u_inv.f_next[247] ;
 wire \u_inv.f_next[248] ;
 wire \u_inv.f_next[249] ;
 wire \u_inv.f_next[24] ;
 wire \u_inv.f_next[250] ;
 wire \u_inv.f_next[251] ;
 wire \u_inv.f_next[252] ;
 wire \u_inv.f_next[253] ;
 wire \u_inv.f_next[254] ;
 wire \u_inv.f_next[255] ;
 wire \u_inv.f_next[256] ;
 wire \u_inv.f_next[25] ;
 wire \u_inv.f_next[26] ;
 wire \u_inv.f_next[27] ;
 wire \u_inv.f_next[28] ;
 wire \u_inv.f_next[29] ;
 wire \u_inv.f_next[2] ;
 wire \u_inv.f_next[30] ;
 wire \u_inv.f_next[31] ;
 wire \u_inv.f_next[32] ;
 wire \u_inv.f_next[33] ;
 wire \u_inv.f_next[34] ;
 wire \u_inv.f_next[35] ;
 wire \u_inv.f_next[36] ;
 wire \u_inv.f_next[37] ;
 wire \u_inv.f_next[38] ;
 wire \u_inv.f_next[39] ;
 wire \u_inv.f_next[3] ;
 wire \u_inv.f_next[40] ;
 wire \u_inv.f_next[41] ;
 wire \u_inv.f_next[42] ;
 wire \u_inv.f_next[43] ;
 wire \u_inv.f_next[44] ;
 wire \u_inv.f_next[45] ;
 wire \u_inv.f_next[46] ;
 wire \u_inv.f_next[47] ;
 wire \u_inv.f_next[48] ;
 wire \u_inv.f_next[49] ;
 wire \u_inv.f_next[4] ;
 wire \u_inv.f_next[50] ;
 wire \u_inv.f_next[51] ;
 wire \u_inv.f_next[52] ;
 wire \u_inv.f_next[53] ;
 wire \u_inv.f_next[54] ;
 wire \u_inv.f_next[55] ;
 wire \u_inv.f_next[56] ;
 wire \u_inv.f_next[57] ;
 wire \u_inv.f_next[58] ;
 wire \u_inv.f_next[59] ;
 wire \u_inv.f_next[5] ;
 wire \u_inv.f_next[60] ;
 wire \u_inv.f_next[61] ;
 wire \u_inv.f_next[62] ;
 wire \u_inv.f_next[63] ;
 wire \u_inv.f_next[64] ;
 wire \u_inv.f_next[65] ;
 wire \u_inv.f_next[66] ;
 wire \u_inv.f_next[67] ;
 wire \u_inv.f_next[68] ;
 wire \u_inv.f_next[69] ;
 wire \u_inv.f_next[6] ;
 wire \u_inv.f_next[70] ;
 wire \u_inv.f_next[71] ;
 wire \u_inv.f_next[72] ;
 wire \u_inv.f_next[73] ;
 wire \u_inv.f_next[74] ;
 wire \u_inv.f_next[75] ;
 wire \u_inv.f_next[76] ;
 wire \u_inv.f_next[77] ;
 wire \u_inv.f_next[78] ;
 wire \u_inv.f_next[79] ;
 wire \u_inv.f_next[7] ;
 wire \u_inv.f_next[80] ;
 wire \u_inv.f_next[81] ;
 wire \u_inv.f_next[82] ;
 wire \u_inv.f_next[83] ;
 wire \u_inv.f_next[84] ;
 wire \u_inv.f_next[85] ;
 wire \u_inv.f_next[86] ;
 wire \u_inv.f_next[87] ;
 wire \u_inv.f_next[88] ;
 wire \u_inv.f_next[89] ;
 wire \u_inv.f_next[8] ;
 wire \u_inv.f_next[90] ;
 wire \u_inv.f_next[91] ;
 wire \u_inv.f_next[92] ;
 wire \u_inv.f_next[93] ;
 wire \u_inv.f_next[94] ;
 wire \u_inv.f_next[95] ;
 wire \u_inv.f_next[96] ;
 wire \u_inv.f_next[97] ;
 wire \u_inv.f_next[98] ;
 wire \u_inv.f_next[99] ;
 wire \u_inv.f_next[9] ;
 wire \u_inv.f_reg[0] ;
 wire \u_inv.f_reg[100] ;
 wire \u_inv.f_reg[101] ;
 wire \u_inv.f_reg[102] ;
 wire \u_inv.f_reg[103] ;
 wire \u_inv.f_reg[104] ;
 wire \u_inv.f_reg[105] ;
 wire \u_inv.f_reg[106] ;
 wire \u_inv.f_reg[107] ;
 wire \u_inv.f_reg[108] ;
 wire \u_inv.f_reg[109] ;
 wire \u_inv.f_reg[10] ;
 wire \u_inv.f_reg[110] ;
 wire \u_inv.f_reg[111] ;
 wire \u_inv.f_reg[112] ;
 wire \u_inv.f_reg[113] ;
 wire \u_inv.f_reg[114] ;
 wire \u_inv.f_reg[115] ;
 wire \u_inv.f_reg[116] ;
 wire \u_inv.f_reg[117] ;
 wire \u_inv.f_reg[118] ;
 wire \u_inv.f_reg[119] ;
 wire \u_inv.f_reg[11] ;
 wire \u_inv.f_reg[120] ;
 wire \u_inv.f_reg[121] ;
 wire \u_inv.f_reg[122] ;
 wire \u_inv.f_reg[123] ;
 wire \u_inv.f_reg[124] ;
 wire \u_inv.f_reg[125] ;
 wire \u_inv.f_reg[126] ;
 wire \u_inv.f_reg[127] ;
 wire \u_inv.f_reg[128] ;
 wire \u_inv.f_reg[129] ;
 wire \u_inv.f_reg[12] ;
 wire \u_inv.f_reg[130] ;
 wire \u_inv.f_reg[131] ;
 wire \u_inv.f_reg[132] ;
 wire \u_inv.f_reg[133] ;
 wire \u_inv.f_reg[134] ;
 wire \u_inv.f_reg[135] ;
 wire \u_inv.f_reg[136] ;
 wire \u_inv.f_reg[137] ;
 wire \u_inv.f_reg[138] ;
 wire \u_inv.f_reg[139] ;
 wire \u_inv.f_reg[13] ;
 wire \u_inv.f_reg[140] ;
 wire \u_inv.f_reg[141] ;
 wire \u_inv.f_reg[142] ;
 wire \u_inv.f_reg[143] ;
 wire \u_inv.f_reg[144] ;
 wire \u_inv.f_reg[145] ;
 wire \u_inv.f_reg[146] ;
 wire \u_inv.f_reg[147] ;
 wire \u_inv.f_reg[148] ;
 wire \u_inv.f_reg[149] ;
 wire \u_inv.f_reg[14] ;
 wire \u_inv.f_reg[150] ;
 wire \u_inv.f_reg[151] ;
 wire \u_inv.f_reg[152] ;
 wire \u_inv.f_reg[153] ;
 wire \u_inv.f_reg[154] ;
 wire \u_inv.f_reg[155] ;
 wire \u_inv.f_reg[156] ;
 wire \u_inv.f_reg[157] ;
 wire \u_inv.f_reg[158] ;
 wire \u_inv.f_reg[159] ;
 wire \u_inv.f_reg[15] ;
 wire \u_inv.f_reg[160] ;
 wire \u_inv.f_reg[161] ;
 wire \u_inv.f_reg[162] ;
 wire \u_inv.f_reg[163] ;
 wire \u_inv.f_reg[164] ;
 wire \u_inv.f_reg[165] ;
 wire \u_inv.f_reg[166] ;
 wire \u_inv.f_reg[167] ;
 wire \u_inv.f_reg[168] ;
 wire \u_inv.f_reg[169] ;
 wire \u_inv.f_reg[16] ;
 wire \u_inv.f_reg[170] ;
 wire \u_inv.f_reg[171] ;
 wire \u_inv.f_reg[172] ;
 wire \u_inv.f_reg[173] ;
 wire \u_inv.f_reg[174] ;
 wire \u_inv.f_reg[175] ;
 wire \u_inv.f_reg[176] ;
 wire \u_inv.f_reg[177] ;
 wire \u_inv.f_reg[178] ;
 wire \u_inv.f_reg[179] ;
 wire \u_inv.f_reg[17] ;
 wire \u_inv.f_reg[180] ;
 wire \u_inv.f_reg[181] ;
 wire \u_inv.f_reg[182] ;
 wire \u_inv.f_reg[183] ;
 wire \u_inv.f_reg[184] ;
 wire \u_inv.f_reg[185] ;
 wire \u_inv.f_reg[186] ;
 wire \u_inv.f_reg[187] ;
 wire \u_inv.f_reg[188] ;
 wire \u_inv.f_reg[189] ;
 wire \u_inv.f_reg[18] ;
 wire \u_inv.f_reg[190] ;
 wire \u_inv.f_reg[191] ;
 wire \u_inv.f_reg[192] ;
 wire \u_inv.f_reg[193] ;
 wire \u_inv.f_reg[194] ;
 wire \u_inv.f_reg[195] ;
 wire \u_inv.f_reg[196] ;
 wire \u_inv.f_reg[197] ;
 wire \u_inv.f_reg[198] ;
 wire \u_inv.f_reg[199] ;
 wire \u_inv.f_reg[19] ;
 wire \u_inv.f_reg[1] ;
 wire \u_inv.f_reg[200] ;
 wire \u_inv.f_reg[201] ;
 wire \u_inv.f_reg[202] ;
 wire \u_inv.f_reg[203] ;
 wire \u_inv.f_reg[204] ;
 wire \u_inv.f_reg[205] ;
 wire \u_inv.f_reg[206] ;
 wire \u_inv.f_reg[207] ;
 wire \u_inv.f_reg[208] ;
 wire \u_inv.f_reg[209] ;
 wire \u_inv.f_reg[20] ;
 wire \u_inv.f_reg[210] ;
 wire \u_inv.f_reg[211] ;
 wire \u_inv.f_reg[212] ;
 wire \u_inv.f_reg[213] ;
 wire \u_inv.f_reg[214] ;
 wire \u_inv.f_reg[215] ;
 wire \u_inv.f_reg[216] ;
 wire \u_inv.f_reg[217] ;
 wire \u_inv.f_reg[218] ;
 wire \u_inv.f_reg[219] ;
 wire \u_inv.f_reg[21] ;
 wire \u_inv.f_reg[220] ;
 wire \u_inv.f_reg[221] ;
 wire \u_inv.f_reg[222] ;
 wire \u_inv.f_reg[223] ;
 wire \u_inv.f_reg[224] ;
 wire \u_inv.f_reg[225] ;
 wire \u_inv.f_reg[226] ;
 wire \u_inv.f_reg[227] ;
 wire \u_inv.f_reg[228] ;
 wire \u_inv.f_reg[229] ;
 wire \u_inv.f_reg[22] ;
 wire \u_inv.f_reg[230] ;
 wire \u_inv.f_reg[231] ;
 wire \u_inv.f_reg[232] ;
 wire \u_inv.f_reg[233] ;
 wire \u_inv.f_reg[234] ;
 wire \u_inv.f_reg[235] ;
 wire \u_inv.f_reg[236] ;
 wire \u_inv.f_reg[237] ;
 wire \u_inv.f_reg[238] ;
 wire \u_inv.f_reg[239] ;
 wire \u_inv.f_reg[23] ;
 wire \u_inv.f_reg[240] ;
 wire \u_inv.f_reg[241] ;
 wire \u_inv.f_reg[242] ;
 wire \u_inv.f_reg[243] ;
 wire \u_inv.f_reg[244] ;
 wire \u_inv.f_reg[245] ;
 wire \u_inv.f_reg[246] ;
 wire \u_inv.f_reg[247] ;
 wire \u_inv.f_reg[248] ;
 wire \u_inv.f_reg[249] ;
 wire \u_inv.f_reg[24] ;
 wire \u_inv.f_reg[250] ;
 wire \u_inv.f_reg[251] ;
 wire \u_inv.f_reg[252] ;
 wire \u_inv.f_reg[253] ;
 wire \u_inv.f_reg[254] ;
 wire \u_inv.f_reg[255] ;
 wire \u_inv.f_reg[256] ;
 wire \u_inv.f_reg[25] ;
 wire \u_inv.f_reg[26] ;
 wire \u_inv.f_reg[27] ;
 wire \u_inv.f_reg[28] ;
 wire \u_inv.f_reg[29] ;
 wire \u_inv.f_reg[2] ;
 wire \u_inv.f_reg[30] ;
 wire \u_inv.f_reg[31] ;
 wire \u_inv.f_reg[32] ;
 wire \u_inv.f_reg[33] ;
 wire \u_inv.f_reg[34] ;
 wire \u_inv.f_reg[35] ;
 wire \u_inv.f_reg[36] ;
 wire \u_inv.f_reg[37] ;
 wire \u_inv.f_reg[38] ;
 wire \u_inv.f_reg[39] ;
 wire \u_inv.f_reg[3] ;
 wire \u_inv.f_reg[40] ;
 wire \u_inv.f_reg[41] ;
 wire \u_inv.f_reg[42] ;
 wire \u_inv.f_reg[43] ;
 wire \u_inv.f_reg[44] ;
 wire \u_inv.f_reg[45] ;
 wire \u_inv.f_reg[46] ;
 wire \u_inv.f_reg[47] ;
 wire \u_inv.f_reg[48] ;
 wire \u_inv.f_reg[49] ;
 wire \u_inv.f_reg[4] ;
 wire \u_inv.f_reg[50] ;
 wire \u_inv.f_reg[51] ;
 wire \u_inv.f_reg[52] ;
 wire \u_inv.f_reg[53] ;
 wire \u_inv.f_reg[54] ;
 wire \u_inv.f_reg[55] ;
 wire \u_inv.f_reg[56] ;
 wire \u_inv.f_reg[57] ;
 wire \u_inv.f_reg[58] ;
 wire \u_inv.f_reg[59] ;
 wire \u_inv.f_reg[5] ;
 wire \u_inv.f_reg[60] ;
 wire \u_inv.f_reg[61] ;
 wire \u_inv.f_reg[62] ;
 wire \u_inv.f_reg[63] ;
 wire \u_inv.f_reg[64] ;
 wire \u_inv.f_reg[65] ;
 wire \u_inv.f_reg[66] ;
 wire \u_inv.f_reg[67] ;
 wire \u_inv.f_reg[68] ;
 wire \u_inv.f_reg[69] ;
 wire \u_inv.f_reg[6] ;
 wire \u_inv.f_reg[70] ;
 wire \u_inv.f_reg[71] ;
 wire \u_inv.f_reg[72] ;
 wire \u_inv.f_reg[73] ;
 wire \u_inv.f_reg[74] ;
 wire \u_inv.f_reg[75] ;
 wire \u_inv.f_reg[76] ;
 wire \u_inv.f_reg[77] ;
 wire \u_inv.f_reg[78] ;
 wire \u_inv.f_reg[79] ;
 wire \u_inv.f_reg[7] ;
 wire \u_inv.f_reg[80] ;
 wire \u_inv.f_reg[81] ;
 wire \u_inv.f_reg[82] ;
 wire \u_inv.f_reg[83] ;
 wire \u_inv.f_reg[84] ;
 wire \u_inv.f_reg[85] ;
 wire \u_inv.f_reg[86] ;
 wire \u_inv.f_reg[87] ;
 wire \u_inv.f_reg[88] ;
 wire \u_inv.f_reg[89] ;
 wire \u_inv.f_reg[8] ;
 wire \u_inv.f_reg[90] ;
 wire \u_inv.f_reg[91] ;
 wire \u_inv.f_reg[92] ;
 wire \u_inv.f_reg[93] ;
 wire \u_inv.f_reg[94] ;
 wire \u_inv.f_reg[95] ;
 wire \u_inv.f_reg[96] ;
 wire \u_inv.f_reg[97] ;
 wire \u_inv.f_reg[98] ;
 wire \u_inv.f_reg[99] ;
 wire \u_inv.f_reg[9] ;
 wire \u_inv.input_reg[0] ;
 wire \u_inv.input_reg[100] ;
 wire \u_inv.input_reg[101] ;
 wire \u_inv.input_reg[102] ;
 wire \u_inv.input_reg[103] ;
 wire \u_inv.input_reg[104] ;
 wire \u_inv.input_reg[105] ;
 wire \u_inv.input_reg[106] ;
 wire \u_inv.input_reg[107] ;
 wire \u_inv.input_reg[108] ;
 wire \u_inv.input_reg[109] ;
 wire \u_inv.input_reg[10] ;
 wire \u_inv.input_reg[110] ;
 wire \u_inv.input_reg[111] ;
 wire \u_inv.input_reg[112] ;
 wire \u_inv.input_reg[113] ;
 wire \u_inv.input_reg[114] ;
 wire \u_inv.input_reg[115] ;
 wire \u_inv.input_reg[116] ;
 wire \u_inv.input_reg[117] ;
 wire \u_inv.input_reg[118] ;
 wire \u_inv.input_reg[119] ;
 wire \u_inv.input_reg[11] ;
 wire \u_inv.input_reg[120] ;
 wire \u_inv.input_reg[121] ;
 wire \u_inv.input_reg[122] ;
 wire \u_inv.input_reg[123] ;
 wire \u_inv.input_reg[124] ;
 wire \u_inv.input_reg[125] ;
 wire \u_inv.input_reg[126] ;
 wire \u_inv.input_reg[127] ;
 wire \u_inv.input_reg[128] ;
 wire \u_inv.input_reg[129] ;
 wire \u_inv.input_reg[12] ;
 wire \u_inv.input_reg[130] ;
 wire \u_inv.input_reg[131] ;
 wire \u_inv.input_reg[132] ;
 wire \u_inv.input_reg[133] ;
 wire \u_inv.input_reg[134] ;
 wire \u_inv.input_reg[135] ;
 wire \u_inv.input_reg[136] ;
 wire \u_inv.input_reg[137] ;
 wire \u_inv.input_reg[138] ;
 wire \u_inv.input_reg[139] ;
 wire \u_inv.input_reg[13] ;
 wire \u_inv.input_reg[140] ;
 wire \u_inv.input_reg[141] ;
 wire \u_inv.input_reg[142] ;
 wire \u_inv.input_reg[143] ;
 wire \u_inv.input_reg[144] ;
 wire \u_inv.input_reg[145] ;
 wire \u_inv.input_reg[146] ;
 wire \u_inv.input_reg[147] ;
 wire \u_inv.input_reg[148] ;
 wire \u_inv.input_reg[149] ;
 wire \u_inv.input_reg[14] ;
 wire \u_inv.input_reg[150] ;
 wire \u_inv.input_reg[151] ;
 wire \u_inv.input_reg[152] ;
 wire \u_inv.input_reg[153] ;
 wire \u_inv.input_reg[154] ;
 wire \u_inv.input_reg[155] ;
 wire \u_inv.input_reg[156] ;
 wire \u_inv.input_reg[157] ;
 wire \u_inv.input_reg[158] ;
 wire \u_inv.input_reg[159] ;
 wire \u_inv.input_reg[15] ;
 wire \u_inv.input_reg[160] ;
 wire \u_inv.input_reg[161] ;
 wire \u_inv.input_reg[162] ;
 wire \u_inv.input_reg[163] ;
 wire \u_inv.input_reg[164] ;
 wire \u_inv.input_reg[165] ;
 wire \u_inv.input_reg[166] ;
 wire \u_inv.input_reg[167] ;
 wire \u_inv.input_reg[168] ;
 wire \u_inv.input_reg[169] ;
 wire \u_inv.input_reg[16] ;
 wire \u_inv.input_reg[170] ;
 wire \u_inv.input_reg[171] ;
 wire \u_inv.input_reg[172] ;
 wire \u_inv.input_reg[173] ;
 wire \u_inv.input_reg[174] ;
 wire \u_inv.input_reg[175] ;
 wire \u_inv.input_reg[176] ;
 wire \u_inv.input_reg[177] ;
 wire \u_inv.input_reg[178] ;
 wire \u_inv.input_reg[179] ;
 wire \u_inv.input_reg[17] ;
 wire \u_inv.input_reg[180] ;
 wire \u_inv.input_reg[181] ;
 wire \u_inv.input_reg[182] ;
 wire \u_inv.input_reg[183] ;
 wire \u_inv.input_reg[184] ;
 wire \u_inv.input_reg[185] ;
 wire \u_inv.input_reg[186] ;
 wire \u_inv.input_reg[187] ;
 wire \u_inv.input_reg[188] ;
 wire \u_inv.input_reg[189] ;
 wire \u_inv.input_reg[18] ;
 wire \u_inv.input_reg[190] ;
 wire \u_inv.input_reg[191] ;
 wire \u_inv.input_reg[192] ;
 wire \u_inv.input_reg[193] ;
 wire \u_inv.input_reg[194] ;
 wire \u_inv.input_reg[195] ;
 wire \u_inv.input_reg[196] ;
 wire \u_inv.input_reg[197] ;
 wire \u_inv.input_reg[198] ;
 wire \u_inv.input_reg[199] ;
 wire \u_inv.input_reg[19] ;
 wire \u_inv.input_reg[1] ;
 wire \u_inv.input_reg[200] ;
 wire \u_inv.input_reg[201] ;
 wire \u_inv.input_reg[202] ;
 wire \u_inv.input_reg[203] ;
 wire \u_inv.input_reg[204] ;
 wire \u_inv.input_reg[205] ;
 wire \u_inv.input_reg[206] ;
 wire \u_inv.input_reg[207] ;
 wire \u_inv.input_reg[208] ;
 wire \u_inv.input_reg[209] ;
 wire \u_inv.input_reg[20] ;
 wire \u_inv.input_reg[210] ;
 wire \u_inv.input_reg[211] ;
 wire \u_inv.input_reg[212] ;
 wire \u_inv.input_reg[213] ;
 wire \u_inv.input_reg[214] ;
 wire \u_inv.input_reg[215] ;
 wire \u_inv.input_reg[216] ;
 wire \u_inv.input_reg[217] ;
 wire \u_inv.input_reg[218] ;
 wire \u_inv.input_reg[219] ;
 wire \u_inv.input_reg[21] ;
 wire \u_inv.input_reg[220] ;
 wire \u_inv.input_reg[221] ;
 wire \u_inv.input_reg[222] ;
 wire \u_inv.input_reg[223] ;
 wire \u_inv.input_reg[224] ;
 wire \u_inv.input_reg[225] ;
 wire \u_inv.input_reg[226] ;
 wire \u_inv.input_reg[227] ;
 wire \u_inv.input_reg[228] ;
 wire \u_inv.input_reg[229] ;
 wire \u_inv.input_reg[22] ;
 wire \u_inv.input_reg[230] ;
 wire \u_inv.input_reg[231] ;
 wire \u_inv.input_reg[232] ;
 wire \u_inv.input_reg[233] ;
 wire \u_inv.input_reg[234] ;
 wire \u_inv.input_reg[235] ;
 wire \u_inv.input_reg[236] ;
 wire \u_inv.input_reg[237] ;
 wire \u_inv.input_reg[238] ;
 wire \u_inv.input_reg[239] ;
 wire \u_inv.input_reg[23] ;
 wire \u_inv.input_reg[240] ;
 wire \u_inv.input_reg[241] ;
 wire \u_inv.input_reg[242] ;
 wire \u_inv.input_reg[243] ;
 wire \u_inv.input_reg[244] ;
 wire \u_inv.input_reg[245] ;
 wire \u_inv.input_reg[246] ;
 wire \u_inv.input_reg[247] ;
 wire \u_inv.input_reg[248] ;
 wire \u_inv.input_reg[249] ;
 wire \u_inv.input_reg[24] ;
 wire \u_inv.input_reg[250] ;
 wire \u_inv.input_reg[251] ;
 wire \u_inv.input_reg[252] ;
 wire \u_inv.input_reg[253] ;
 wire \u_inv.input_reg[254] ;
 wire \u_inv.input_reg[255] ;
 wire \u_inv.input_reg[25] ;
 wire \u_inv.input_reg[26] ;
 wire \u_inv.input_reg[27] ;
 wire \u_inv.input_reg[28] ;
 wire \u_inv.input_reg[29] ;
 wire \u_inv.input_reg[2] ;
 wire \u_inv.input_reg[30] ;
 wire \u_inv.input_reg[31] ;
 wire \u_inv.input_reg[32] ;
 wire \u_inv.input_reg[33] ;
 wire \u_inv.input_reg[34] ;
 wire \u_inv.input_reg[35] ;
 wire \u_inv.input_reg[36] ;
 wire \u_inv.input_reg[37] ;
 wire \u_inv.input_reg[38] ;
 wire \u_inv.input_reg[39] ;
 wire \u_inv.input_reg[3] ;
 wire \u_inv.input_reg[40] ;
 wire \u_inv.input_reg[41] ;
 wire \u_inv.input_reg[42] ;
 wire \u_inv.input_reg[43] ;
 wire \u_inv.input_reg[44] ;
 wire \u_inv.input_reg[45] ;
 wire \u_inv.input_reg[46] ;
 wire \u_inv.input_reg[47] ;
 wire \u_inv.input_reg[48] ;
 wire \u_inv.input_reg[49] ;
 wire \u_inv.input_reg[4] ;
 wire \u_inv.input_reg[50] ;
 wire \u_inv.input_reg[51] ;
 wire \u_inv.input_reg[52] ;
 wire \u_inv.input_reg[53] ;
 wire \u_inv.input_reg[54] ;
 wire \u_inv.input_reg[55] ;
 wire \u_inv.input_reg[56] ;
 wire \u_inv.input_reg[57] ;
 wire \u_inv.input_reg[58] ;
 wire \u_inv.input_reg[59] ;
 wire \u_inv.input_reg[5] ;
 wire \u_inv.input_reg[60] ;
 wire \u_inv.input_reg[61] ;
 wire \u_inv.input_reg[62] ;
 wire \u_inv.input_reg[63] ;
 wire \u_inv.input_reg[64] ;
 wire \u_inv.input_reg[65] ;
 wire \u_inv.input_reg[66] ;
 wire \u_inv.input_reg[67] ;
 wire \u_inv.input_reg[68] ;
 wire \u_inv.input_reg[69] ;
 wire \u_inv.input_reg[6] ;
 wire \u_inv.input_reg[70] ;
 wire \u_inv.input_reg[71] ;
 wire \u_inv.input_reg[72] ;
 wire \u_inv.input_reg[73] ;
 wire \u_inv.input_reg[74] ;
 wire \u_inv.input_reg[75] ;
 wire \u_inv.input_reg[76] ;
 wire \u_inv.input_reg[77] ;
 wire \u_inv.input_reg[78] ;
 wire \u_inv.input_reg[79] ;
 wire \u_inv.input_reg[7] ;
 wire \u_inv.input_reg[80] ;
 wire \u_inv.input_reg[81] ;
 wire \u_inv.input_reg[82] ;
 wire \u_inv.input_reg[83] ;
 wire \u_inv.input_reg[84] ;
 wire \u_inv.input_reg[85] ;
 wire \u_inv.input_reg[86] ;
 wire \u_inv.input_reg[87] ;
 wire \u_inv.input_reg[88] ;
 wire \u_inv.input_reg[89] ;
 wire \u_inv.input_reg[8] ;
 wire \u_inv.input_reg[90] ;
 wire \u_inv.input_reg[91] ;
 wire \u_inv.input_reg[92] ;
 wire \u_inv.input_reg[93] ;
 wire \u_inv.input_reg[94] ;
 wire \u_inv.input_reg[95] ;
 wire \u_inv.input_reg[96] ;
 wire \u_inv.input_reg[97] ;
 wire \u_inv.input_reg[98] ;
 wire \u_inv.input_reg[99] ;
 wire \u_inv.input_reg[9] ;
 wire \u_inv.input_valid ;
 wire \u_inv.load_input ;
 wire \u_inv.state[0] ;
 wire \u_inv.state[1] ;
 wire \u_trng.bit_cnt[0] ;
 wire \u_trng.bit_cnt[1] ;
 wire \u_trng.bit_cnt[2] ;
 wire \u_trng.entropy_bit ;
 wire \u_trng.entropy_ff1 ;
 wire \u_trng.entropy_raw ;
 wire \u_trng.have_prev ;
 wire \u_trng.prev_sample ;
 wire \u_trng.u_ro5.and_out ;
 wire \u_trng.u_ro5.c[0] ;
 wire \u_trng.u_ro5.c[1] ;
 wire \u_trng.u_ro5.c[2] ;
 wire \u_trng.u_ro5.c[3] ;
 wire \u_trng.u_ro5.c[4] ;
 wire \u_trng.u_ro7.and_out ;
 wire \u_trng.u_ro7.c[0] ;
 wire \u_trng.u_ro7.c[1] ;
 wire \u_trng.u_ro7.c[2] ;
 wire \u_trng.u_ro7.c[3] ;
 wire \u_trng.u_ro7.c[4] ;
 wire \u_trng.u_ro7.c[5] ;
 wire \u_trng.u_ro7.c[6] ;
 wire \u_trng.u_ro9.and_out ;
 wire \u_trng.u_ro9.c[0] ;
 wire \u_trng.u_ro9.c[1] ;
 wire \u_trng.u_ro9.c[2] ;
 wire \u_trng.u_ro9.c[3] ;
 wire \u_trng.u_ro9.c[4] ;
 wire \u_trng.u_ro9.c[5] ;
 wire \u_trng.u_ro9.c[6] ;
 wire \u_trng.u_ro9.c[7] ;
 wire \u_trng.u_ro9.c[8] ;
 wire net1060;
 wire net1061;
 wire net15;
 wire net16;
 wire net1062;
 wire net1063;
 wire clknet_leaf_0_clk;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire wr_prev;
 wire net5065;
 wire net5066;
 wire net5067;
 wire net5068;
 wire net5069;
 wire net5070;
 wire net5071;
 wire net5072;
 wire net5073;
 wire net5074;
 wire net5075;
 wire net5076;
 wire net5077;
 wire net5078;
 wire net5079;
 wire net5080;
 wire net5081;
 wire net5082;
 wire net5083;
 wire net5084;
 wire net5085;
 wire net5086;
 wire net5087;
 wire net5088;
 wire net5089;
 wire net5090;
 wire net5091;
 wire net5092;
 wire net5093;
 wire net5094;
 wire net5095;
 wire net5096;
 wire net5097;
 wire net5098;
 wire net5099;
 wire net5100;
 wire net5101;
 wire net5102;
 wire net5103;
 wire net5104;
 wire net5105;
 wire net5106;
 wire net5107;
 wire net5108;
 wire net5109;
 wire net5110;
 wire net5111;
 wire net5112;
 wire net5113;
 wire net5114;
 wire net5115;
 wire net5116;
 wire net5117;
 wire net5118;
 wire net5119;
 wire net5120;
 wire net5121;
 wire net5122;
 wire net5123;
 wire net5124;
 wire net5125;
 wire net5126;
 wire net5127;
 wire net5128;
 wire net5129;
 wire net5130;
 wire net5131;
 wire net5132;
 wire net5133;
 wire net5134;
 wire net5135;
 wire net5136;
 wire net5137;
 wire net5138;
 wire net5139;
 wire net5140;
 wire net5141;
 wire net5142;
 wire net5143;
 wire net5144;
 wire net5145;
 wire net5146;
 wire net5147;
 wire net5148;
 wire net5149;
 wire net5150;
 wire net5151;
 wire net5152;
 wire net5153;
 wire net5154;
 wire net5155;
 wire net5156;
 wire net5157;
 wire net5158;
 wire net5159;
 wire net5160;
 wire net5161;
 wire net5162;
 wire net5163;
 wire net5164;
 wire net5165;
 wire net5166;
 wire net5167;
 wire net5168;
 wire net5169;
 wire net5170;
 wire net5171;
 wire net5172;
 wire net5173;
 wire net5174;
 wire net5175;
 wire net5176;
 wire net5177;
 wire net5178;
 wire net5179;
 wire net5180;
 wire net5181;
 wire net5182;
 wire net5183;
 wire net5184;
 wire net5185;
 wire net5186;
 wire net5187;
 wire net5188;
 wire net5189;
 wire net5190;
 wire net5191;
 wire net5192;
 wire net5193;
 wire net5194;
 wire net5195;
 wire net5196;
 wire net5197;
 wire net5198;
 wire net5199;
 wire net5200;
 wire net5201;
 wire net5202;
 wire net5203;
 wire net5204;
 wire net5205;
 wire net5206;
 wire net5207;
 wire net5208;
 wire net5209;
 wire net5210;
 wire net5211;
 wire net5212;
 wire net5213;
 wire net5214;
 wire net5215;
 wire net5216;
 wire net5217;
 wire net5218;
 wire net5219;
 wire net5220;
 wire net5221;
 wire net5222;
 wire net5223;
 wire net5224;
 wire net5225;
 wire net5226;
 wire net5227;
 wire net5228;
 wire net5229;
 wire net5230;
 wire net5231;
 wire net5232;
 wire net5233;
 wire net5234;
 wire net5235;
 wire net5236;
 wire net5237;
 wire net5238;
 wire net5239;
 wire net5240;
 wire net5241;
 wire net5242;
 wire net5243;
 wire net5244;
 wire net5245;
 wire net5246;
 wire net5247;
 wire net5248;
 wire net5249;
 wire net5250;
 wire net5251;
 wire net5252;
 wire net5253;
 wire net5254;
 wire net5255;
 wire net5256;
 wire net5257;
 wire net5258;
 wire net5259;
 wire net5260;
 wire net5261;
 wire net5262;
 wire net5263;
 wire net5264;
 wire net5265;
 wire net5266;
 wire net5267;
 wire net5268;
 wire net5269;
 wire net5270;
 wire net5271;
 wire net5272;
 wire net5273;
 wire net5274;
 wire net5275;
 wire net5276;
 wire net5277;
 wire net5278;
 wire net5279;
 wire net5280;
 wire net5281;
 wire net5282;
 wire net5283;
 wire net5284;
 wire net5285;
 wire net5286;
 wire net5287;
 wire net5288;
 wire net5289;
 wire net5290;
 wire net5291;
 wire net5292;
 wire net5293;
 wire net5294;
 wire net5295;
 wire net5296;
 wire net5297;
 wire net5298;
 wire net5299;
 wire net5300;
 wire net5301;
 wire net5302;
 wire net5303;
 wire net5304;
 wire net5305;
 wire net5306;
 wire net5307;
 wire net5308;
 wire net5309;
 wire net5310;
 wire net5311;
 wire net5312;
 wire net5313;
 wire net5314;
 wire net5315;
 wire net5316;
 wire net5317;
 wire net5318;
 wire net5319;
 wire net5320;
 wire net5321;
 wire net5322;
 wire net5323;
 wire net5324;
 wire net5325;
 wire net5326;
 wire net5327;
 wire net5328;
 wire net5329;
 wire net5330;
 wire net5331;
 wire net5332;
 wire net5333;
 wire net5334;
 wire net5335;
 wire net5336;
 wire net5337;
 wire net5338;
 wire net5339;
 wire net5340;
 wire net5341;
 wire net5342;
 wire net5343;
 wire net5344;
 wire net5345;
 wire net5346;
 wire net5347;
 wire net5348;
 wire net1141;
 wire net5350;
 wire net5351;
 wire net5352;
 wire net5353;
 wire net5354;
 wire net5355;
 wire net5356;
 wire net5357;
 wire net5358;
 wire net5359;
 wire net5360;
 wire net5361;
 wire net5362;
 wire net5363;
 wire net5364;
 wire net5365;
 wire net5366;
 wire net5367;
 wire net5368;
 wire net5369;
 wire net5370;
 wire net5371;
 wire net5372;
 wire net5373;
 wire net5374;
 wire net5375;
 wire net5376;
 wire net5377;
 wire net5378;
 wire net5379;
 wire net5380;
 wire net5381;
 wire net5382;
 wire net5383;
 wire net5384;
 wire net5385;
 wire net5386;
 wire net5387;
 wire net5388;
 wire net5389;
 wire net5390;
 wire net5391;
 wire net5392;
 wire net5393;
 wire net5394;
 wire net5395;
 wire net5396;
 wire net5397;
 wire net5398;
 wire net5399;
 wire net5400;
 wire net5401;
 wire net5402;
 wire net5403;
 wire net5404;
 wire net5405;
 wire net5406;
 wire net5407;
 wire net5408;
 wire net5409;
 wire net5410;
 wire net5411;
 wire net5412;
 wire net5413;
 wire net5414;
 wire net5415;
 wire net5416;
 wire net5417;
 wire net5418;
 wire net5419;
 wire net5420;
 wire net5421;
 wire net5422;
 wire net5423;
 wire net5424;
 wire net5425;
 wire net5426;
 wire net5427;
 wire net5428;
 wire net5429;
 wire net5430;
 wire net5431;
 wire net5432;
 wire net5433;
 wire net5434;
 wire net5435;
 wire net5436;
 wire net5437;
 wire net5438;
 wire net5439;
 wire net5440;
 wire net5441;
 wire net5442;
 wire net5443;
 wire net5444;
 wire net5445;
 wire net5446;
 wire net5447;
 wire net5448;
 wire net5449;
 wire net5450;
 wire net5451;
 wire net5452;
 wire net5453;
 wire net5454;
 wire net5455;
 wire net5456;
 wire net5457;
 wire net5458;
 wire net5459;
 wire net5460;
 wire net5461;
 wire net5462;
 wire net5463;
 wire net5464;
 wire net5465;
 wire net5466;
 wire net5467;
 wire net5468;
 wire net5469;
 wire net5470;
 wire net5471;
 wire net5472;
 wire net5473;
 wire net5474;
 wire net5475;
 wire net5476;
 wire net5477;
 wire net5478;
 wire net5479;
 wire net5480;
 wire net5481;
 wire net5482;
 wire net5483;
 wire net5484;
 wire net5485;
 wire net5486;
 wire net5487;
 wire net5488;
 wire net5489;
 wire net5490;
 wire net5491;
 wire net5492;
 wire net5493;
 wire net5494;
 wire net5495;
 wire net5496;
 wire net5497;
 wire net5498;
 wire net5499;
 wire net5500;
 wire net5501;
 wire net5502;
 wire net5503;
 wire net5504;
 wire net5505;
 wire net5506;
 wire net5507;
 wire net5508;
 wire net5509;
 wire net5510;
 wire net5511;
 wire net5512;
 wire net5513;
 wire net5514;
 wire net5515;
 wire net5516;
 wire net5517;
 wire net5518;
 wire net5519;
 wire net5520;
 wire net5521;
 wire net5522;
 wire net5523;
 wire net5524;
 wire net5525;
 wire net5526;
 wire net5527;
 wire net5528;
 wire net5529;
 wire net5530;
 wire net5531;
 wire net5532;
 wire net5533;
 wire net5534;
 wire net5535;
 wire net5536;
 wire net5537;
 wire net5538;
 wire net5539;
 wire net5540;
 wire net5541;
 wire net5542;
 wire net5543;
 wire net5544;
 wire net5545;
 wire net5546;
 wire net5547;
 wire net5548;
 wire net5549;
 wire net5550;
 wire net5551;
 wire net5552;
 wire net5553;
 wire net5554;
 wire net5555;
 wire net5556;
 wire net5557;
 wire net5558;
 wire net5559;
 wire net5560;
 wire net5561;
 wire net5562;
 wire net5563;
 wire net5564;
 wire net5565;
 wire net5566;
 wire net5567;
 wire net5568;
 wire net5569;
 wire net5570;
 wire net5571;
 wire net5572;
 wire net5573;
 wire net5574;
 wire net5575;
 wire net5576;
 wire net5577;
 wire net5578;
 wire net5579;
 wire net5580;
 wire net5581;
 wire net5582;
 wire net5583;
 wire net5584;
 wire net5585;
 wire net5586;
 wire net5587;
 wire net5588;
 wire net5589;
 wire net5590;
 wire net5591;
 wire net5592;
 wire net5593;
 wire net5594;
 wire net5595;
 wire net5596;
 wire net5597;
 wire net5598;
 wire net5599;
 wire net5600;
 wire net5601;
 wire net5602;
 wire net5603;
 wire net5604;
 wire net5605;
 wire net5606;
 wire net5607;
 wire net5608;
 wire net5609;
 wire net5610;
 wire net5611;
 wire net5612;
 wire net5613;
 wire net5614;
 wire net5615;
 wire net5616;
 wire net5617;
 wire net5618;
 wire net5619;
 wire net5620;
 wire net5621;
 wire net5622;
 wire net5623;
 wire net5624;
 wire net5625;
 wire net5626;
 wire net5627;
 wire net5628;
 wire net5629;
 wire net5630;
 wire net5631;
 wire net5632;
 wire net5633;
 wire net5634;
 wire net5635;
 wire net5636;
 wire net5637;
 wire net5638;
 wire net5639;
 wire net5640;
 wire net5641;
 wire net5642;
 wire net5643;
 wire net5644;
 wire net5645;
 wire net5646;
 wire net5647;
 wire net5648;
 wire net5649;
 wire net5650;
 wire net5651;
 wire net5652;
 wire net5653;
 wire net5654;
 wire net5655;
 wire net5656;
 wire net5657;
 wire net5658;
 wire net5659;
 wire net5660;
 wire net5661;
 wire net5662;
 wire net5663;
 wire net5664;
 wire net5665;
 wire net5666;
 wire net5667;
 wire net5668;
 wire net5669;
 wire net5670;
 wire net5671;
 wire net5672;
 wire net5673;
 wire net5674;
 wire net5675;
 wire net5676;
 wire net5677;
 wire net5678;
 wire net5679;
 wire net5680;
 wire net5681;
 wire net5682;
 wire net5683;
 wire net5684;
 wire net5685;
 wire net5686;
 wire net5687;
 wire net5688;
 wire net5689;
 wire net5690;
 wire net5691;
 wire net5692;
 wire net5693;
 wire net5694;
 wire net5695;
 wire net5696;
 wire net5697;
 wire net5698;
 wire net5699;
 wire net5700;
 wire net5701;
 wire net5702;
 wire net5703;
 wire net5704;
 wire net5705;
 wire net5706;
 wire net5707;
 wire net5708;
 wire net5709;
 wire net5710;
 wire net5711;
 wire net5712;
 wire net5713;
 wire net5714;
 wire net5715;
 wire net5716;
 wire net5717;
 wire net5718;
 wire net5719;
 wire net5720;
 wire net5721;
 wire net5722;
 wire net5723;
 wire net5724;
 wire net5725;
 wire net5726;
 wire net5727;
 wire net5728;
 wire net5729;
 wire net5730;
 wire net5731;
 wire net5732;
 wire net5733;
 wire net5734;
 wire net5735;
 wire net5736;
 wire net5737;
 wire net5738;
 wire net5739;
 wire net5740;
 wire net5741;
 wire net5742;
 wire net5743;
 wire net5744;
 wire net5745;
 wire net5746;
 wire net5747;
 wire net5748;
 wire net5749;
 wire net5750;
 wire net5751;
 wire net5752;
 wire net5753;
 wire net5754;
 wire net5755;
 wire net5756;
 wire net5757;
 wire net5758;
 wire net5759;
 wire net5760;
 wire net5761;
 wire net5762;
 wire net5763;
 wire net5764;
 wire net5765;
 wire net5766;
 wire net5767;
 wire net5768;
 wire net5769;
 wire net5770;
 wire net5771;
 wire net5772;
 wire net5773;
 wire net5774;
 wire net5775;
 wire net5776;
 wire net5777;
 wire net5778;
 wire net5779;
 wire net5780;
 wire net5781;
 wire net5782;
 wire net5783;
 wire net5784;
 wire net5785;
 wire net5786;
 wire net5787;
 wire net5788;
 wire net5789;
 wire net5790;
 wire net5791;
 wire net5792;
 wire net5793;
 wire net5794;
 wire net5795;
 wire net5796;
 wire net5797;
 wire net5798;
 wire net5799;
 wire net5800;
 wire net5801;
 wire net5802;
 wire net5803;
 wire net5804;
 wire net5805;
 wire net5806;
 wire net5807;
 wire net5808;
 wire net5809;
 wire net5810;
 wire net5811;
 wire net5812;
 wire net5813;
 wire net5814;
 wire net5815;
 wire net5816;
 wire net5817;
 wire net5818;
 wire net5819;
 wire net5820;
 wire net5821;
 wire net5822;
 wire net5823;
 wire net5824;
 wire net5825;
 wire net5826;
 wire net5827;
 wire net5828;
 wire net5829;
 wire net5830;
 wire net5831;
 wire net5832;
 wire net5833;
 wire net5834;
 wire net5835;
 wire net5836;
 wire net5837;
 wire net5838;
 wire net5839;
 wire net5840;
 wire net5841;
 wire net5842;
 wire net5843;
 wire net5844;
 wire net5845;
 wire net5846;
 wire net5847;
 wire net5848;
 wire net5849;
 wire net5850;
 wire net5851;
 wire net5852;
 wire net5853;
 wire net5854;
 wire net5855;
 wire net5856;
 wire net5857;
 wire net5858;
 wire net5859;
 wire net5860;
 wire net5861;
 wire net5862;
 wire net5863;
 wire net5864;
 wire net5865;
 wire net5866;
 wire net5867;
 wire net5868;
 wire net5869;
 wire net5870;
 wire net5871;
 wire net5872;
 wire net5873;
 wire net5874;
 wire net5875;
 wire net5876;
 wire net5877;
 wire net5878;
 wire net5879;
 wire net5880;
 wire net5881;
 wire net5882;
 wire net5883;
 wire net5884;
 wire net5885;
 wire net5886;
 wire net5887;
 wire net5888;
 wire net5889;
 wire net5890;
 wire net5891;
 wire net5892;
 wire net5893;
 wire net5894;
 wire net5895;
 wire net5896;
 wire net5897;
 wire net5898;
 wire net5899;
 wire net5900;
 wire net5901;
 wire net5902;
 wire net5903;
 wire net5904;
 wire net5905;
 wire net5906;
 wire net5907;
 wire net5908;
 wire net5909;
 wire net5910;
 wire net5911;
 wire net5912;
 wire net5913;
 wire net5914;
 wire net5915;
 wire net5916;
 wire net5917;
 wire net5918;
 wire net5919;
 wire net5920;
 wire net5921;
 wire net5922;
 wire net5923;
 wire net5924;
 wire net5925;
 wire net5926;
 wire net5927;
 wire net5928;
 wire net5929;
 wire net5930;
 wire net5931;
 wire net5932;
 wire net5933;
 wire net5934;
 wire net5935;
 wire net5936;
 wire net5937;
 wire net5938;
 wire net5939;
 wire net5940;
 wire net5941;
 wire net5942;
 wire net5943;
 wire net5944;
 wire net5945;
 wire net5946;
 wire net5947;
 wire net5948;
 wire net5949;
 wire net5950;
 wire net5951;
 wire net5952;
 wire net5953;
 wire net5954;
 wire net5955;
 wire net5956;
 wire net5957;
 wire net5958;
 wire net5959;
 wire net5960;
 wire net5961;
 wire net5962;
 wire net5963;
 wire net5964;
 wire net5965;
 wire net5966;
 wire net5967;
 wire net5968;
 wire net5969;
 wire net5970;
 wire net5971;
 wire net5972;
 wire net5973;
 wire net5974;
 wire net5975;
 wire net5976;
 wire net5977;
 wire net5978;
 wire net5979;
 wire net5980;
 wire net5981;
 wire net5982;
 wire net5983;
 wire net5984;
 wire net5985;
 wire net5986;
 wire net5987;
 wire net5988;
 wire net5989;
 wire net5990;
 wire net5991;
 wire net5992;
 wire net5993;
 wire net5994;
 wire net5995;
 wire net5996;
 wire net5997;
 wire net5998;
 wire net5999;
 wire net6000;
 wire net6001;
 wire net6002;
 wire net6003;
 wire net6004;
 wire net6005;
 wire net6006;
 wire net6007;
 wire net6008;
 wire net6009;
 wire net6010;
 wire net6011;
 wire net6012;
 wire net6013;
 wire net6014;
 wire net6015;
 wire net6016;
 wire net6017;
 wire net6018;
 wire net6019;
 wire net6020;
 wire net6021;
 wire net6022;
 wire net6023;
 wire net6024;
 wire net6025;
 wire net6026;
 wire net6027;
 wire net6028;
 wire net6029;
 wire net6030;
 wire net6031;
 wire net6032;
 wire net6033;
 wire net6034;
 wire net6035;
 wire net6036;
 wire net6037;
 wire net6038;
 wire net6039;
 wire net6040;
 wire net6041;
 wire net6042;
 wire net6043;
 wire net6044;
 wire net6045;
 wire net6046;
 wire net6047;
 wire net6048;
 wire net6049;
 wire net6050;
 wire net6051;
 wire net6052;
 wire net6053;
 wire net6054;
 wire net6055;
 wire net6056;
 wire net6057;
 wire net6058;
 wire net6059;
 wire net6060;
 wire net6061;
 wire net6062;
 wire net6063;
 wire net6064;
 wire net6065;
 wire net6066;
 wire net6067;
 wire net6068;
 wire net6069;
 wire net6070;
 wire net6071;
 wire net6072;
 wire net6073;
 wire net6074;
 wire net6075;
 wire net6076;
 wire net6077;
 wire net6078;
 wire net6079;
 wire net6080;
 wire net6081;
 wire net6082;
 wire net6083;
 wire net6084;
 wire net6085;
 wire net6086;
 wire net6087;
 wire net6088;
 wire net6089;
 wire net6090;
 wire net6091;
 wire net6092;
 wire net6093;
 wire net6094;
 wire net6095;
 wire net6096;
 wire net6097;
 wire net6098;
 wire net6099;
 wire net6100;
 wire net6101;
 wire net6102;
 wire net6103;
 wire net6104;
 wire net6105;
 wire net6106;
 wire net6107;
 wire net6108;
 wire net6109;
 wire net6110;
 wire net6111;
 wire net6112;
 wire net6113;
 wire net6114;
 wire net6115;
 wire net6116;
 wire net6117;
 wire net6118;
 wire net6119;
 wire net6120;
 wire net6121;
 wire net6122;
 wire net6123;
 wire net6124;
 wire net6125;
 wire net6126;
 wire net6127;
 wire net6128;
 wire net6129;
 wire net6130;
 wire net6131;
 wire net6132;
 wire net6133;
 wire net6134;
 wire net6135;
 wire net6136;
 wire net6137;
 wire net6138;
 wire net6139;
 wire net6140;
 wire net6141;
 wire net6142;
 wire net6143;
 wire net6144;
 wire net6145;
 wire net6146;
 wire net6147;
 wire net6148;
 wire net6149;
 wire net6150;
 wire net6151;
 wire net6152;
 wire net6153;
 wire net6154;
 wire net6155;
 wire net6156;
 wire net6157;
 wire net6158;
 wire net6159;
 wire net6160;
 wire net6161;
 wire net6162;
 wire net6163;
 wire net6164;
 wire net6165;
 wire net6166;
 wire net6167;
 wire net6168;
 wire net6169;
 wire net6170;
 wire net6171;
 wire net6172;
 wire net6173;
 wire net6174;
 wire net6175;
 wire net6176;
 wire net6177;
 wire net6178;
 wire net6179;
 wire net6180;
 wire net6181;
 wire net6182;
 wire net6183;
 wire net6184;
 wire net6185;
 wire net6186;
 wire net6187;
 wire net6188;
 wire net6189;
 wire net6190;
 wire net6191;
 wire net6192;
 wire net6193;
 wire net6194;
 wire net6195;
 wire net6196;
 wire net6197;
 wire net6198;
 wire net6199;
 wire net6200;
 wire net6201;
 wire net6202;
 wire net6203;
 wire net6204;
 wire net6205;
 wire net6206;
 wire net6207;
 wire net6208;
 wire net6209;
 wire net6210;
 wire net6211;
 wire net6212;
 wire net6213;
 wire net6214;
 wire net6215;
 wire net6216;
 wire net6217;
 wire net6218;
 wire net6219;
 wire net6220;
 wire net6221;
 wire net6222;
 wire net6223;
 wire net6224;
 wire net6225;
 wire net6226;
 wire net6227;
 wire net6228;
 wire net6229;
 wire net6230;
 wire net6231;
 wire net6232;
 wire net6233;
 wire net6234;
 wire net6235;
 wire net6236;
 wire net6237;
 wire net6238;
 wire net6239;
 wire net6240;
 wire net6241;
 wire net6242;
 wire net6243;
 wire net6244;
 wire net6245;
 wire net6246;
 wire net6247;
 wire net6248;
 wire net6249;
 wire net6250;
 wire net6251;
 wire net6252;
 wire net6253;
 wire net6254;
 wire net6255;
 wire net6256;
 wire net6257;
 wire net6258;
 wire net6259;
 wire net6260;
 wire net6261;
 wire net6262;
 wire net6263;
 wire net6264;
 wire net6265;
 wire net6266;
 wire net6267;
 wire net6268;
 wire net6269;
 wire net6270;
 wire net6271;
 wire net6272;
 wire net6273;
 wire net6274;
 wire net6275;
 wire net6276;
 wire net6277;
 wire net6278;
 wire net6279;
 wire net6280;
 wire net6281;
 wire net6282;
 wire net6283;
 wire net6284;
 wire net6285;
 wire net6286;
 wire net6287;
 wire net6288;
 wire net6289;
 wire net6290;
 wire net6291;
 wire net6292;
 wire net6293;
 wire net6294;
 wire net6295;
 wire net6296;
 wire net6297;
 wire net6298;
 wire net6299;
 wire net6300;
 wire net6301;
 wire net6302;
 wire net6303;
 wire net6304;
 wire net6305;
 wire net6306;
 wire net6307;
 wire net6308;
 wire net6309;
 wire net6310;
 wire net6311;
 wire net6312;
 wire net6313;
 wire net6314;
 wire net6315;
 wire net6316;
 wire net6317;
 wire net6318;
 wire net6319;
 wire net6320;
 wire net6321;
 wire net6322;
 wire net6323;
 wire net6324;
 wire net6325;
 wire net6326;
 wire net6327;
 wire net6328;
 wire net6329;
 wire net6330;
 wire net6331;
 wire net6332;
 wire net6333;
 wire net6334;
 wire net6335;
 wire net6336;
 wire net6337;
 wire net6338;
 wire net6339;
 wire net6340;
 wire net6341;
 wire net6342;
 wire net6343;
 wire net6344;
 wire net6345;
 wire net6346;
 wire net6347;
 wire net6348;
 wire net6349;
 wire net6350;
 wire net6351;
 wire net6352;
 wire net6353;
 wire net6354;
 wire net6355;
 wire net6356;
 wire net6357;
 wire net6358;
 wire net6359;
 wire net6360;
 wire net6361;
 wire net6362;
 wire net6363;
 wire net6364;
 wire net6365;
 wire net6366;
 wire net6367;
 wire net6368;
 wire net6369;
 wire net6370;
 wire net6371;
 wire net6372;
 wire net6373;
 wire net6374;
 wire net6375;
 wire net6376;
 wire net6377;
 wire net6378;
 wire net6379;
 wire net6380;
 wire net6381;
 wire net6382;
 wire net6383;
 wire net6384;
 wire net6385;
 wire net6386;
 wire net6387;
 wire net6388;
 wire net6389;
 wire net6390;
 wire net6391;
 wire net6392;
 wire net6393;
 wire net6394;
 wire net6395;
 wire net6396;
 wire net6397;
 wire net6398;
 wire net6399;
 wire net6400;
 wire net6401;
 wire net6402;
 wire net6403;
 wire net6404;
 wire net6405;
 wire net6406;
 wire net6407;
 wire net6408;
 wire net6409;
 wire net6410;
 wire net6411;
 wire net6412;
 wire net6413;
 wire net6414;
 wire net6415;
 wire net6416;
 wire net6417;
 wire net6418;
 wire net6419;
 wire net6420;
 wire net6421;
 wire net6422;
 wire net6423;
 wire net6424;
 wire net6425;
 wire net6426;
 wire net6427;
 wire net6428;
 wire net6429;
 wire net6430;
 wire net6431;
 wire net6432;
 wire net6433;
 wire net6434;
 wire net6435;
 wire net6436;
 wire net6437;
 wire net6438;
 wire net6439;
 wire net6440;
 wire net6441;
 wire net6442;
 wire net6443;
 wire net6444;
 wire net6445;
 wire net6446;
 wire net6447;
 wire net6448;
 wire net6449;
 wire net6450;
 wire net6451;
 wire net6452;
 wire net6453;
 wire net6454;
 wire net6455;
 wire net6456;
 wire net6457;
 wire net6458;
 wire net6459;
 wire net6460;
 wire net6461;
 wire net6462;
 wire net6463;
 wire net6464;
 wire net6465;
 wire net6466;
 wire net6467;
 wire net6468;
 wire net6469;
 wire net6470;
 wire net6471;
 wire net6472;
 wire net6473;
 wire net6474;
 wire net6475;
 wire net6476;
 wire net6477;
 wire net6478;
 wire net6479;
 wire net6480;
 wire net6481;
 wire net6482;
 wire net6483;
 wire net6484;
 wire net6485;
 wire net6486;
 wire net6487;
 wire net6488;
 wire net6489;
 wire net6490;
 wire net6491;
 wire net6492;
 wire net6493;
 wire net6494;
 wire net6495;
 wire net6496;
 wire net6497;
 wire net6498;
 wire net6499;
 wire net6500;
 wire net6501;
 wire net6502;
 wire net6503;
 wire net6504;
 wire net6505;
 wire net6506;
 wire net6507;
 wire net6508;
 wire net6509;
 wire net6510;
 wire net6511;
 wire net6512;
 wire net6513;
 wire net6514;
 wire net6515;
 wire net6516;
 wire net6517;
 wire net6518;
 wire net6519;
 wire net6520;
 wire net6521;
 wire net6522;
 wire net6523;
 wire net6524;
 wire net6525;
 wire net6526;
 wire net6527;
 wire net6528;
 wire net6529;
 wire net6530;
 wire net6531;
 wire net6532;
 wire net6533;
 wire net6534;
 wire net6535;
 wire net6536;
 wire net6537;
 wire net6538;
 wire net6539;
 wire net6540;
 wire net6541;
 wire net6542;
 wire net6543;
 wire net6544;
 wire net6545;
 wire net6546;
 wire net6547;
 wire net6548;
 wire net6549;
 wire net6550;
 wire net6551;
 wire net6552;
 wire net6553;
 wire net6554;
 wire net6555;
 wire net6556;
 wire net6557;
 wire net6558;
 wire net6559;
 wire net6560;
 wire net6561;
 wire net6562;
 wire net6563;
 wire net6564;
 wire net6565;
 wire net6566;
 wire net6567;
 wire net6568;
 wire net6569;
 wire net6570;
 wire net6571;
 wire net6572;
 wire net6573;
 wire net6574;
 wire net6575;
 wire net6576;
 wire net6577;
 wire net6578;
 wire net6579;
 wire net6580;
 wire net6581;
 wire net6582;
 wire net6583;
 wire net6584;
 wire net6585;
 wire net6586;
 wire net6587;
 wire net6588;
 wire net6589;
 wire net6590;
 wire net6591;
 wire net6592;
 wire net6593;
 wire net6594;
 wire net6595;
 wire net6596;
 wire net6597;
 wire net6598;
 wire net6599;
 wire net6600;
 wire net6601;
 wire net6602;
 wire net6603;
 wire net6604;
 wire net6605;
 wire net6606;
 wire net6607;
 wire net6608;
 wire net6609;
 wire net6610;
 wire net6611;
 wire net6612;
 wire net6613;
 wire net6614;
 wire net6615;
 wire net6616;
 wire net6617;
 wire net6618;
 wire net6619;
 wire net6620;
 wire net6621;
 wire net6622;
 wire net6623;
 wire net6624;
 wire net6625;
 wire net6626;
 wire net6627;
 wire net6628;
 wire net6629;
 wire net6630;
 wire net6631;
 wire net6632;
 wire net6633;
 wire net6634;
 wire net6635;
 wire net6636;
 wire net6637;
 wire net6638;
 wire net6639;
 wire net6640;
 wire net6641;
 wire net6642;
 wire net6643;
 wire net6644;
 wire net6645;
 wire net6646;
 wire net6647;
 wire net6648;
 wire net6649;
 wire net6650;
 wire net6651;
 wire net6652;
 wire net6653;
 wire net6654;
 wire net6655;
 wire net6656;
 wire net6657;
 wire net6658;
 wire net6659;
 wire net6660;
 wire net6661;
 wire net6662;
 wire net6663;
 wire net6664;
 wire net6665;
 wire net6666;
 wire net6667;
 wire net6668;
 wire net6669;
 wire net6670;
 wire net6671;
 wire net6672;
 wire net6673;
 wire net6674;
 wire net6675;
 wire net6676;
 wire net6677;
 wire net6678;
 wire net6679;
 wire net6680;
 wire net6681;
 wire net6682;
 wire net6683;
 wire net6684;
 wire net6685;
 wire net6686;
 wire net6687;
 wire net6688;
 wire net6689;
 wire net6690;
 wire net6691;
 wire net6692;
 wire net6693;
 wire net6694;
 wire net6695;
 wire net6696;
 wire net6697;
 wire net6698;
 wire net6699;
 wire net6700;
 wire net6701;
 wire net6702;
 wire net6703;
 wire net6704;
 wire net6705;
 wire net6706;
 wire net6707;
 wire net6708;
 wire net6709;
 wire net6710;
 wire net6711;
 wire net6712;
 wire net6713;
 wire net6714;
 wire net6715;
 wire net6716;
 wire net6717;
 wire net6718;
 wire net6719;
 wire net6720;
 wire net6721;
 wire net6722;
 wire net6723;
 wire net6724;
 wire net6725;
 wire net6726;
 wire net6727;
 wire net6728;
 wire net6729;
 wire net6730;
 wire net6731;
 wire net6732;
 wire net6733;
 wire net6734;
 wire net6735;
 wire net6736;
 wire net6737;
 wire net6738;
 wire net6739;
 wire net6740;
 wire net6741;
 wire net6742;
 wire net6743;
 wire net6744;
 wire net6745;
 wire net6746;
 wire net6747;
 wire net6748;
 wire net6749;
 wire net6750;
 wire net6751;
 wire net6752;
 wire net6753;
 wire net6754;
 wire net6755;
 wire net6756;
 wire net6757;
 wire net6758;
 wire net6759;
 wire net6760;
 wire net6761;
 wire net6762;
 wire net6763;
 wire net6764;
 wire net6765;
 wire net6766;
 wire net6767;
 wire net6768;
 wire net6769;
 wire net6770;
 wire net6771;
 wire net6772;
 wire net6773;
 wire net6774;
 wire net6775;
 wire net6776;
 wire net6777;
 wire net6778;
 wire net6779;
 wire net6780;
 wire net6781;
 wire net6782;
 wire net6783;
 wire net6784;
 wire net6785;
 wire net6786;
 wire net6787;
 wire net6788;
 wire net6789;
 wire net6790;
 wire net6791;
 wire net6792;
 wire net6793;
 wire net6794;
 wire net6795;
 wire net6796;
 wire net6797;
 wire net6798;
 wire net6799;
 wire net6800;
 wire net6801;
 wire net6802;
 wire net6803;
 wire net6804;
 wire net6805;
 wire net6806;
 wire net6807;
 wire net6808;
 wire net6809;
 wire net6810;
 wire net6811;
 wire net6812;
 wire net6813;
 wire net6814;
 wire net6815;
 wire net6816;
 wire net6817;
 wire net6818;
 wire net6819;
 wire net6820;
 wire net6821;
 wire net6822;
 wire net6823;
 wire net6824;
 wire net6825;
 wire net6826;
 wire net6827;
 wire net6828;
 wire net6829;
 wire net6830;
 wire net6831;
 wire net6832;
 wire net6833;
 wire net6834;
 wire net6835;
 wire net6836;
 wire net6837;
 wire net6838;
 wire net6839;
 wire net6840;
 wire net6841;
 wire net6842;
 wire net6843;
 wire net6844;
 wire net6845;
 wire net6846;
 wire net6847;
 wire net6848;
 wire net6849;
 wire net6850;
 wire net6851;
 wire net6852;
 wire net6853;
 wire net6854;
 wire net6855;
 wire net6856;
 wire net6857;
 wire net6858;
 wire net6859;
 wire net6860;
 wire net6861;
 wire net6862;
 wire net6863;
 wire net6864;
 wire net6865;
 wire net6866;
 wire net6867;
 wire net6868;
 wire net6869;
 wire net6870;
 wire net6871;
 wire net6872;
 wire net6873;
 wire net6874;
 wire net6875;
 wire net6876;
 wire net6877;
 wire net6878;
 wire net6879;
 wire net6880;
 wire net6881;
 wire net6882;
 wire net6883;
 wire net6884;
 wire net6885;
 wire net6886;
 wire net6887;
 wire net6888;
 wire net6889;
 wire net6890;
 wire net6891;
 wire net6892;
 wire net6893;
 wire net6894;
 wire net6895;
 wire net6896;
 wire net6897;
 wire net6898;
 wire net6899;
 wire net6900;
 wire net6901;
 wire net6902;
 wire net6903;
 wire net6904;
 wire net6905;
 wire net6906;
 wire net6907;
 wire net6908;
 wire net6909;
 wire net6910;
 wire net6911;
 wire net6912;
 wire net6913;
 wire net6914;
 wire net6915;
 wire net6916;
 wire net6917;
 wire net6918;
 wire net6919;
 wire net6920;
 wire net6921;
 wire net6922;
 wire net6923;
 wire net6924;
 wire net6925;
 wire net6926;
 wire net6927;
 wire net6928;
 wire net6929;
 wire net6930;
 wire net6931;
 wire net6932;
 wire net6933;
 wire net6934;
 wire net6935;
 wire net6936;
 wire net6937;
 wire net6938;
 wire net6939;
 wire net6940;
 wire net6941;
 wire net6942;
 wire net6943;
 wire net6944;
 wire net6945;
 wire net6946;
 wire net6947;
 wire net6948;
 wire net6949;
 wire net6950;
 wire net6951;
 wire net6952;
 wire net6953;
 wire net6954;
 wire net6955;
 wire net6956;
 wire net6957;
 wire net6958;
 wire net6959;
 wire net6960;
 wire net6961;
 wire net6962;
 wire net6963;
 wire net6964;
 wire net6965;
 wire net6966;
 wire net6967;
 wire net6968;
 wire net6969;
 wire net6970;
 wire net6971;
 wire net6972;
 wire net6973;
 wire net6974;
 wire net6975;
 wire net6976;
 wire net6977;
 wire net6978;
 wire net6979;
 wire net6980;
 wire net6981;
 wire net6982;
 wire net6983;
 wire net6984;
 wire net6985;
 wire net6986;
 wire net6987;
 wire net6988;
 wire net6989;
 wire net6990;
 wire net6991;
 wire net6992;
 wire net6993;
 wire net6994;
 wire net6995;
 wire net6996;
 wire net6997;
 wire net6998;
 wire net6999;
 wire net7000;
 wire net7001;
 wire net7002;
 wire net7003;
 wire net7004;
 wire net7005;
 wire net7006;
 wire net7007;
 wire net7008;
 wire net7009;
 wire net7010;
 wire net7011;
 wire net7012;
 wire net7013;
 wire net7014;
 wire net7015;
 wire net7016;
 wire net7017;
 wire net7018;
 wire net7019;
 wire net7020;
 wire net7021;
 wire net7022;
 wire net7023;
 wire net7024;
 wire net7025;
 wire net7026;
 wire net7027;
 wire net7028;
 wire net7029;
 wire net7030;
 wire net7031;
 wire net7032;
 wire net7033;
 wire net7034;
 wire net7035;
 wire net7036;
 wire net7037;
 wire net7038;
 wire net7039;
 wire net7040;
 wire net7041;
 wire net7042;
 wire net7043;
 wire net7044;
 wire net7045;
 wire net7046;
 wire net7047;
 wire net7048;
 wire net7049;
 wire net7050;
 wire net7051;
 wire net7052;
 wire net7053;
 wire net7054;
 wire net7055;
 wire net7056;
 wire net7057;
 wire net7058;
 wire net7059;
 wire net7060;
 wire net7061;
 wire net7062;
 wire net7063;
 wire net7064;
 wire net7065;
 wire net7066;
 wire net7067;
 wire net7068;
 wire net7069;
 wire net7070;
 wire net7071;
 wire net7072;
 wire net7073;
 wire net7074;
 wire net7075;
 wire net7076;
 wire net7077;
 wire net7078;
 wire net7079;
 wire net7080;
 wire net7081;
 wire net7082;
 wire net7083;
 wire net7084;
 wire net7085;
 wire net7086;
 wire net7087;
 wire net7088;
 wire net7089;
 wire net7090;
 wire net7091;
 wire net7092;
 wire net7093;
 wire net7094;
 wire net7095;
 wire net7096;
 wire net7097;
 wire net7098;
 wire net7099;
 wire net7100;
 wire net7101;
 wire net7102;
 wire net7103;
 wire net7104;
 wire net7105;
 wire net7106;
 wire net7107;
 wire net7108;
 wire net7109;
 wire net7110;
 wire net7111;
 wire net7112;
 wire net7113;
 wire net7114;
 wire net7115;
 wire net7116;
 wire net7117;
 wire net7118;
 wire net7119;
 wire net7120;
 wire net7121;
 wire net7122;
 wire net7123;
 wire net7124;
 wire net7125;
 wire net7126;
 wire net7127;
 wire net7128;
 wire net7129;
 wire net7130;
 wire net7131;
 wire net7132;
 wire net7133;
 wire net7134;
 wire net7135;
 wire net7136;
 wire net7137;
 wire net7138;
 wire net7139;
 wire net7140;
 wire net7141;
 wire net7142;
 wire net7143;
 wire net7144;
 wire net7145;
 wire net7146;
 wire net7147;
 wire net7148;
 wire net7149;
 wire net7150;
 wire net7151;
 wire net7152;
 wire net7153;
 wire net7154;
 wire net7155;
 wire net7156;
 wire net7157;
 wire net7158;
 wire net7159;
 wire net7160;
 wire net7161;
 wire net7162;
 wire net7163;
 wire net7164;
 wire net7165;
 wire net7166;
 wire net7167;
 wire net7168;
 wire net7169;
 wire net7170;
 wire net7171;
 wire net7172;
 wire net7173;
 wire net7174;
 wire net7175;
 wire net7176;
 wire net7177;
 wire net7178;
 wire net7179;
 wire net7180;
 wire net7181;
 wire net7182;
 wire net7183;
 wire net7184;
 wire net7185;
 wire net7186;
 wire net7187;
 wire net7188;
 wire net7189;
 wire net7190;
 wire net7191;
 wire net7192;
 wire net7193;
 wire net7194;
 wire net7195;
 wire net7196;
 wire net7197;
 wire net7198;
 wire net7199;
 wire net7200;
 wire net7201;
 wire net7202;
 wire net7203;
 wire net7204;
 wire net7205;
 wire net7206;
 wire net7207;
 wire net7208;
 wire net7209;
 wire net7210;
 wire net7211;
 wire net7212;
 wire net7213;
 wire net7214;
 wire net7215;
 wire net7216;
 wire net7217;
 wire net7218;
 wire net7219;
 wire net7220;
 wire net7221;
 wire net7222;
 wire net7223;
 wire net7224;
 wire net7225;
 wire net7226;
 wire net7227;
 wire net7228;
 wire net7229;
 wire net7230;
 wire net7231;
 wire net7232;
 wire net7233;
 wire net7234;
 wire net7235;
 wire net7236;
 wire net7237;
 wire net7238;
 wire net7239;
 wire net7240;
 wire net7241;
 wire net7242;
 wire net7243;
 wire net7244;
 wire net7245;
 wire net7246;
 wire net7247;
 wire net7248;
 wire net7249;
 wire net7250;
 wire net7251;
 wire net7252;
 wire net7253;
 wire net7254;
 wire net7255;
 wire net7256;
 wire net7257;
 wire net7258;
 wire net7259;
 wire net7260;
 wire net7261;
 wire net7262;
 wire net7263;
 wire net7264;
 wire net7265;
 wire net7266;
 wire net7267;
 wire net7268;
 wire net7269;
 wire net7270;
 wire net7271;
 wire net7272;
 wire net7273;
 wire net7274;
 wire net7275;
 wire net7276;
 wire net7277;
 wire net7278;
 wire net7279;
 wire net7280;
 wire net7281;
 wire net7282;
 wire net7283;
 wire net7284;
 wire net7285;
 wire net7286;
 wire net7287;
 wire net7288;
 wire net7289;
 wire net7290;
 wire net7291;
 wire net7292;
 wire net7293;
 wire net7294;
 wire net7295;
 wire net7296;
 wire net7297;
 wire net7298;
 wire net7299;
 wire net7300;
 wire net7301;
 wire net7302;
 wire net7303;
 wire net7304;
 wire net7305;
 wire net7306;
 wire net7307;
 wire net7308;
 wire net7309;
 wire net7310;
 wire net7311;
 wire net7312;
 wire net7313;
 wire net7314;
 wire net7315;
 wire net7316;
 wire net7317;
 wire net7318;
 wire net7319;
 wire net7320;
 wire net7321;
 wire net7322;
 wire net7323;
 wire net7324;
 wire net7325;
 wire net7326;
 wire net7327;
 wire net7328;
 wire net7329;
 wire net7330;
 wire net7331;
 wire net7332;
 wire net7333;
 wire net7334;
 wire net7335;
 wire net7336;
 wire net7337;
 wire net7338;
 wire net7339;
 wire net7340;
 wire net7341;
 wire net7342;
 wire net7343;
 wire net7344;
 wire net7345;
 wire net7346;
 wire net7347;
 wire net7348;
 wire net7349;
 wire net7350;
 wire net7351;
 wire net7352;
 wire net7353;
 wire net7354;
 wire net7355;
 wire net7356;
 wire net7357;
 wire net7358;
 wire net7359;
 wire net7360;
 wire net7361;
 wire net7362;
 wire net7363;
 wire net7364;
 wire net7365;
 wire net7366;
 wire net7367;
 wire net7368;
 wire net7369;
 wire net7370;
 wire net7371;
 wire net7372;
 wire net7373;
 wire net7374;
 wire net7375;
 wire net7376;
 wire net7377;
 wire net7378;
 wire net7379;
 wire net7380;
 wire net7381;
 wire net7382;
 wire net7383;
 wire net7384;
 wire net7385;
 wire net7386;
 wire net7387;
 wire net7388;
 wire net7389;
 wire net7390;
 wire net7391;
 wire net7392;
 wire net7393;
 wire net7394;
 wire net7395;
 wire net7396;
 wire net7397;
 wire net7398;
 wire net7399;
 wire net7400;
 wire net7401;
 wire net7402;
 wire net7403;
 wire net7404;
 wire net7405;
 wire net7406;
 wire net7407;
 wire net7408;
 wire net7409;
 wire net7410;
 wire net7411;
 wire net7412;
 wire net7413;
 wire net7414;
 wire net7415;
 wire net7416;
 wire net7417;
 wire net7418;
 wire net7419;
 wire net7420;
 wire net7421;
 wire net7422;
 wire net7423;
 wire net7424;
 wire net7425;
 wire net7426;
 wire net7427;
 wire net7428;
 wire net7429;
 wire net7430;
 wire net7431;
 wire net7432;
 wire net7433;
 wire net7434;
 wire net7435;
 wire net7436;
 wire net7437;
 wire net7438;
 wire net7439;
 wire net7440;
 wire net7441;
 wire net7442;
 wire net7443;
 wire net7444;
 wire net7445;
 wire net7446;
 wire net7447;
 wire net7448;
 wire net7449;
 wire net7450;
 wire net7451;
 wire net7452;
 wire net7453;
 wire net7454;
 wire net7455;
 wire net7456;
 wire net7457;
 wire net7458;
 wire net7459;
 wire net7460;
 wire net7461;
 wire net7462;
 wire net7463;
 wire net7464;
 wire net7465;
 wire net7466;
 wire net7467;
 wire net7468;
 wire net7469;
 wire net7470;
 wire net7471;
 wire net7472;
 wire net7473;
 wire net7474;
 wire net7475;
 wire net7476;
 wire net7477;
 wire net7478;
 wire net7479;
 wire net7480;
 wire net7481;
 wire net7482;
 wire net7483;
 wire net7484;
 wire net7485;
 wire net7486;
 wire net7487;
 wire net7488;
 wire net7489;
 wire net7490;
 wire net7491;
 wire net7492;
 wire net7493;
 wire net7494;
 wire net7495;
 wire net7496;
 wire net7497;
 wire net7498;
 wire net7499;
 wire net7500;
 wire net7501;
 wire net7502;
 wire net7503;
 wire net7504;
 wire net7505;
 wire net7506;
 wire net7507;
 wire net7508;
 wire net7509;
 wire net7510;
 wire net7511;
 wire net7512;
 wire net7513;
 wire net7514;
 wire net7515;
 wire net7516;
 wire net7517;
 wire net7518;
 wire net7519;
 wire net7520;
 wire net7521;
 wire net7522;
 wire net7523;
 wire net7524;
 wire net7525;
 wire net7526;
 wire net7527;
 wire net7528;
 wire net7529;
 wire net7530;
 wire net7531;
 wire net7532;
 wire net7533;
 wire net7534;
 wire net7535;
 wire net7536;
 wire net7537;
 wire net7538;
 wire net7539;
 wire net7540;
 wire net7541;
 wire net7542;
 wire net7543;
 wire net7544;
 wire net7545;
 wire net7546;
 wire net7547;
 wire net7548;
 wire net7549;
 wire net7550;
 wire net7551;
 wire net7552;
 wire net7553;
 wire net7554;
 wire net7555;
 wire net7556;
 wire net7557;
 wire net7558;
 wire net7559;
 wire net7560;
 wire net7561;
 wire net7562;
 wire net7563;
 wire net7564;
 wire net7565;
 wire net7566;
 wire net7567;
 wire net7568;
 wire net7569;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_5_0_0_clk;
 wire clknet_5_1_0_clk;
 wire clknet_5_2_0_clk;
 wire clknet_5_3_0_clk;
 wire clknet_5_4_0_clk;
 wire clknet_5_5_0_clk;
 wire clknet_5_6_0_clk;
 wire clknet_5_7_0_clk;
 wire clknet_5_8_0_clk;
 wire clknet_5_9_0_clk;
 wire clknet_5_10_0_clk;
 wire clknet_5_11_0_clk;
 wire clknet_5_12_0_clk;
 wire clknet_5_13_0_clk;
 wire clknet_5_14_0_clk;
 wire clknet_5_15_0_clk;
 wire clknet_5_16_0_clk;
 wire clknet_5_17_0_clk;
 wire clknet_5_18_0_clk;
 wire clknet_5_19_0_clk;
 wire clknet_5_20_0_clk;
 wire clknet_5_21_0_clk;
 wire clknet_5_22_0_clk;
 wire clknet_5_23_0_clk;
 wire clknet_5_24_0_clk;
 wire clknet_5_25_0_clk;
 wire clknet_5_26_0_clk;
 wire clknet_5_27_0_clk;
 wire clknet_5_28_0_clk;
 wire clknet_5_29_0_clk;
 wire clknet_5_30_0_clk;
 wire clknet_5_31_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire [0:0] _24689_;
 wire [0:0] _24690_;

 sg13g2_nand3_1 _24691_ (.B(net7135),
    .C(net6162),
    .A(net3252),
    .Y(_17140_));
 sg13g2_o21ai_1 _24692_ (.B1(_17140_),
    .Y(_01364_),
    .A1(_18500_),
    .A2(net6163));
 sg13g2_nand3_1 _24693_ (.B(net7135),
    .C(net6161),
    .A(net2328),
    .Y(_17141_));
 sg13g2_o21ai_1 _24694_ (.B1(_17141_),
    .Y(_01365_),
    .A1(_18499_),
    .A2(net6161));
 sg13g2_nand3_1 _24695_ (.B(net7135),
    .C(net6160),
    .A(net2980),
    .Y(_17142_));
 sg13g2_o21ai_1 _24696_ (.B1(_17142_),
    .Y(_01366_),
    .A1(_18498_),
    .A2(net6160));
 sg13g2_nand3_1 _24697_ (.B(net7135),
    .C(net6161),
    .A(net2877),
    .Y(_17143_));
 sg13g2_o21ai_1 _24698_ (.B1(_17143_),
    .Y(_01367_),
    .A1(_18497_),
    .A2(net6161));
 sg13g2_nand3_1 _24699_ (.B(net7135),
    .C(net6162),
    .A(net2361),
    .Y(_17144_));
 sg13g2_o21ai_1 _24700_ (.B1(_17144_),
    .Y(_01368_),
    .A1(_18496_),
    .A2(net6162));
 sg13g2_nand3_1 _24701_ (.B(net7136),
    .C(net6162),
    .A(net2890),
    .Y(_17145_));
 sg13g2_o21ai_1 _24702_ (.B1(_17145_),
    .Y(_01369_),
    .A1(_18495_),
    .A2(net6162));
 sg13g2_nand3_1 _24703_ (.B(net7137),
    .C(net6156),
    .A(net2225),
    .Y(_17146_));
 sg13g2_o21ai_1 _24704_ (.B1(_17146_),
    .Y(_01370_),
    .A1(_18494_),
    .A2(net6156));
 sg13g2_nand3_1 _24705_ (.B(net7137),
    .C(net6156),
    .A(net3128),
    .Y(_17147_));
 sg13g2_o21ai_1 _24706_ (.B1(_17147_),
    .Y(_01371_),
    .A1(_18493_),
    .A2(net6164));
 sg13g2_nand3_1 _24707_ (.B(net7126),
    .C(net6139),
    .A(net3157),
    .Y(_17148_));
 sg13g2_o21ai_1 _24708_ (.B1(_17148_),
    .Y(_01372_),
    .A1(_18492_),
    .A2(net6139));
 sg13g2_nand3_1 _24709_ (.B(net7137),
    .C(net6156),
    .A(net2397),
    .Y(_17149_));
 sg13g2_o21ai_1 _24710_ (.B1(_17149_),
    .Y(_01373_),
    .A1(_18491_),
    .A2(net6156));
 sg13g2_nand3_1 _24711_ (.B(net7126),
    .C(net6139),
    .A(net2437),
    .Y(_17150_));
 sg13g2_o21ai_1 _24712_ (.B1(_17150_),
    .Y(_01374_),
    .A1(_18490_),
    .A2(net6139));
 sg13g2_nand3_1 _24713_ (.B(net7126),
    .C(net6139),
    .A(net3360),
    .Y(_17151_));
 sg13g2_o21ai_1 _24714_ (.B1(_17151_),
    .Y(_01375_),
    .A1(_18489_),
    .A2(net6139));
 sg13g2_nand3_1 _24715_ (.B(net7126),
    .C(net6156),
    .A(net2401),
    .Y(_17152_));
 sg13g2_o21ai_1 _24716_ (.B1(_17152_),
    .Y(_01376_),
    .A1(_18488_),
    .A2(net6141));
 sg13g2_nand3_1 _24717_ (.B(net7127),
    .C(net6139),
    .A(net3585),
    .Y(_17153_));
 sg13g2_o21ai_1 _24718_ (.B1(_17153_),
    .Y(_01377_),
    .A1(_18487_),
    .A2(net6139));
 sg13g2_nand3_1 _24719_ (.B(net7126),
    .C(net6140),
    .A(net2587),
    .Y(_17154_));
 sg13g2_o21ai_1 _24720_ (.B1(_17154_),
    .Y(_01378_),
    .A1(_18486_),
    .A2(net6140));
 sg13g2_nand3_1 _24721_ (.B(net7126),
    .C(net6140),
    .A(net3299),
    .Y(_17155_));
 sg13g2_o21ai_1 _24722_ (.B1(_17155_),
    .Y(_01379_),
    .A1(_18485_),
    .A2(net6140));
 sg13g2_nand3_1 _24723_ (.B(net7126),
    .C(net6140),
    .A(\u_inv.d_next[130] ),
    .Y(_17156_));
 sg13g2_o21ai_1 _24724_ (.B1(net1242),
    .Y(_01380_),
    .A1(_18484_),
    .A2(net6140));
 sg13g2_nand3_1 _24725_ (.B(net7128),
    .C(net6140),
    .A(net3363),
    .Y(_17157_));
 sg13g2_o21ai_1 _24726_ (.B1(_17157_),
    .Y(_01381_),
    .A1(_18483_),
    .A2(net6140));
 sg13g2_nand3_1 _24727_ (.B(net7128),
    .C(net6134),
    .A(net3413),
    .Y(_17158_));
 sg13g2_o21ai_1 _24728_ (.B1(_17158_),
    .Y(_01382_),
    .A1(_18482_),
    .A2(net6135));
 sg13g2_nand3_1 _24729_ (.B(net7128),
    .C(net6134),
    .A(net3296),
    .Y(_17159_));
 sg13g2_o21ai_1 _24730_ (.B1(_17159_),
    .Y(_01383_),
    .A1(net3556),
    .A2(net6135));
 sg13g2_nand3_1 _24731_ (.B(net7128),
    .C(net6134),
    .A(net3225),
    .Y(_17160_));
 sg13g2_o21ai_1 _24732_ (.B1(_17160_),
    .Y(_01384_),
    .A1(_18480_),
    .A2(net6134));
 sg13g2_nand3_1 _24733_ (.B(net7128),
    .C(net6135),
    .A(net3475),
    .Y(_17161_));
 sg13g2_o21ai_1 _24734_ (.B1(_17161_),
    .Y(_01385_),
    .A1(_18479_),
    .A2(net6135));
 sg13g2_nand3_1 _24735_ (.B(net7119),
    .C(net6116),
    .A(net2826),
    .Y(_17162_));
 sg13g2_o21ai_1 _24736_ (.B1(_17162_),
    .Y(_01386_),
    .A1(_18478_),
    .A2(net6116));
 sg13g2_nand3_1 _24737_ (.B(net7119),
    .C(net6116),
    .A(net3307),
    .Y(_17163_));
 sg13g2_o21ai_1 _24738_ (.B1(_17163_),
    .Y(_01387_),
    .A1(_18477_),
    .A2(net6116));
 sg13g2_nand3_1 _24739_ (.B(net7119),
    .C(net6115),
    .A(net2082),
    .Y(_17164_));
 sg13g2_o21ai_1 _24740_ (.B1(_17164_),
    .Y(_01388_),
    .A1(net2675),
    .A2(net6115));
 sg13g2_nand3_1 _24741_ (.B(net7119),
    .C(net6116),
    .A(net3568),
    .Y(_17165_));
 sg13g2_o21ai_1 _24742_ (.B1(_17165_),
    .Y(_01389_),
    .A1(_18475_),
    .A2(net6116));
 sg13g2_nand3_1 _24743_ (.B(net7119),
    .C(net6115),
    .A(net2606),
    .Y(_17166_));
 sg13g2_o21ai_1 _24744_ (.B1(_17166_),
    .Y(_01390_),
    .A1(_18474_),
    .A2(net6115));
 sg13g2_nand3_1 _24745_ (.B(net7119),
    .C(net6115),
    .A(net3253),
    .Y(_17167_));
 sg13g2_o21ai_1 _24746_ (.B1(_17167_),
    .Y(_01391_),
    .A1(_18473_),
    .A2(net6117));
 sg13g2_nand3_1 _24747_ (.B(net7119),
    .C(net6117),
    .A(net2744),
    .Y(_17168_));
 sg13g2_o21ai_1 _24748_ (.B1(_17168_),
    .Y(_01392_),
    .A1(_18472_),
    .A2(net6117));
 sg13g2_nand3_1 _24749_ (.B(net7119),
    .C(net6116),
    .A(net3396),
    .Y(_17169_));
 sg13g2_o21ai_1 _24750_ (.B1(_17169_),
    .Y(_01393_),
    .A1(_18471_),
    .A2(net6116));
 sg13g2_nand3_1 _24751_ (.B(net7118),
    .C(net6115),
    .A(net2726),
    .Y(_17170_));
 sg13g2_o21ai_1 _24752_ (.B1(_17170_),
    .Y(_01394_),
    .A1(_18470_),
    .A2(net6115));
 sg13g2_nand3_1 _24753_ (.B(net7118),
    .C(net6114),
    .A(net2835),
    .Y(_17171_));
 sg13g2_o21ai_1 _24754_ (.B1(_17171_),
    .Y(_01395_),
    .A1(_18469_),
    .A2(net6114));
 sg13g2_nand3_1 _24755_ (.B(net7118),
    .C(net6114),
    .A(net2694),
    .Y(_17172_));
 sg13g2_o21ai_1 _24756_ (.B1(_17172_),
    .Y(_01396_),
    .A1(_18468_),
    .A2(net6115));
 sg13g2_nand3_1 _24757_ (.B(net7118),
    .C(net6114),
    .A(net3625),
    .Y(_17173_));
 sg13g2_o21ai_1 _24758_ (.B1(_17173_),
    .Y(_01397_),
    .A1(_18467_),
    .A2(net6114));
 sg13g2_nand3_1 _24759_ (.B(net7118),
    .C(net6113),
    .A(net3366),
    .Y(_17174_));
 sg13g2_o21ai_1 _24760_ (.B1(_17174_),
    .Y(_01398_),
    .A1(_18466_),
    .A2(net6112));
 sg13g2_nand3_1 _24761_ (.B(net7118),
    .C(net6113),
    .A(net1902),
    .Y(_17175_));
 sg13g2_o21ai_1 _24762_ (.B1(_17175_),
    .Y(_01399_),
    .A1(_18465_),
    .A2(net6113));
 sg13g2_nand3_1 _24763_ (.B(net7118),
    .C(net6113),
    .A(net2581),
    .Y(_17176_));
 sg13g2_o21ai_1 _24764_ (.B1(_17176_),
    .Y(_01400_),
    .A1(_18464_),
    .A2(net6112));
 sg13g2_nand3_1 _24765_ (.B(net7118),
    .C(net6114),
    .A(net3285),
    .Y(_17177_));
 sg13g2_o21ai_1 _24766_ (.B1(_17177_),
    .Y(_01401_),
    .A1(_18463_),
    .A2(net6113));
 sg13g2_nand3_1 _24767_ (.B(net7111),
    .C(net6113),
    .A(net2589),
    .Y(_17178_));
 sg13g2_o21ai_1 _24768_ (.B1(_17178_),
    .Y(_01402_),
    .A1(_18462_),
    .A2(net6111));
 sg13g2_nand3_1 _24769_ (.B(net7111),
    .C(net6113),
    .A(net2490),
    .Y(_17179_));
 sg13g2_o21ai_1 _24770_ (.B1(_17179_),
    .Y(_01403_),
    .A1(_18461_),
    .A2(net6111));
 sg13g2_nand3_1 _24771_ (.B(net7110),
    .C(net6111),
    .A(net2886),
    .Y(_17180_));
 sg13g2_o21ai_1 _24772_ (.B1(_17180_),
    .Y(_01404_),
    .A1(_18460_),
    .A2(net6111));
 sg13g2_nand3_1 _24773_ (.B(net7110),
    .C(net6112),
    .A(net2950),
    .Y(_17181_));
 sg13g2_o21ai_1 _24774_ (.B1(_17181_),
    .Y(_01405_),
    .A1(_18459_),
    .A2(net6111));
 sg13g2_nand3_1 _24775_ (.B(net7111),
    .C(net6113),
    .A(net2669),
    .Y(_17182_));
 sg13g2_o21ai_1 _24776_ (.B1(_17182_),
    .Y(_01406_),
    .A1(_18458_),
    .A2(net6111));
 sg13g2_nand3_1 _24777_ (.B(net7110),
    .C(net6111),
    .A(net3220),
    .Y(_17183_));
 sg13g2_o21ai_1 _24778_ (.B1(_17183_),
    .Y(_01407_),
    .A1(_18457_),
    .A2(net6111));
 sg13g2_nand3_1 _24779_ (.B(net7111),
    .C(net6095),
    .A(net2471),
    .Y(_17184_));
 sg13g2_o21ai_1 _24780_ (.B1(_17184_),
    .Y(_01408_),
    .A1(_18456_),
    .A2(net6094));
 sg13g2_nand3_1 _24781_ (.B(net7111),
    .C(net6095),
    .A(net3314),
    .Y(_17185_));
 sg13g2_o21ai_1 _24782_ (.B1(_17185_),
    .Y(_01409_),
    .A1(_18455_),
    .A2(net6094));
 sg13g2_nand3_1 _24783_ (.B(net7111),
    .C(net6095),
    .A(net3105),
    .Y(_17186_));
 sg13g2_o21ai_1 _24784_ (.B1(_17186_),
    .Y(_01410_),
    .A1(_18454_),
    .A2(net6095));
 sg13g2_nand3_1 _24785_ (.B(net7110),
    .C(net6093),
    .A(net2266),
    .Y(_17187_));
 sg13g2_o21ai_1 _24786_ (.B1(_17187_),
    .Y(_01411_),
    .A1(_18453_),
    .A2(net6093));
 sg13g2_nand3_1 _24787_ (.B(net7110),
    .C(net6093),
    .A(net2006),
    .Y(_17188_));
 sg13g2_o21ai_1 _24788_ (.B1(_17188_),
    .Y(_01412_),
    .A1(_18452_),
    .A2(net6093));
 sg13g2_nand3_1 _24789_ (.B(net7110),
    .C(net6093),
    .A(net1496),
    .Y(_17189_));
 sg13g2_o21ai_1 _24790_ (.B1(_17189_),
    .Y(_01413_),
    .A1(_18451_),
    .A2(net6093));
 sg13g2_nand3_1 _24791_ (.B(net7110),
    .C(net6093),
    .A(net2712),
    .Y(_17190_));
 sg13g2_o21ai_1 _24792_ (.B1(_17190_),
    .Y(_01414_),
    .A1(_18450_),
    .A2(net6093));
 sg13g2_nand3_1 _24793_ (.B(net7108),
    .C(net6091),
    .A(net1539),
    .Y(_17191_));
 sg13g2_o21ai_1 _24794_ (.B1(_17191_),
    .Y(_01415_),
    .A1(_18449_),
    .A2(net6091));
 sg13g2_nand3_1 _24795_ (.B(net7109),
    .C(net6092),
    .A(net2991),
    .Y(_17192_));
 sg13g2_o21ai_1 _24796_ (.B1(_17192_),
    .Y(_01416_),
    .A1(_18448_),
    .A2(net6092));
 sg13g2_nand3_1 _24797_ (.B(net7109),
    .C(net6091),
    .A(net3181),
    .Y(_17193_));
 sg13g2_o21ai_1 _24798_ (.B1(_17193_),
    .Y(_01417_),
    .A1(_18447_),
    .A2(net6091));
 sg13g2_nand3_1 _24799_ (.B(net7108),
    .C(net6091),
    .A(net3058),
    .Y(_17194_));
 sg13g2_o21ai_1 _24800_ (.B1(_17194_),
    .Y(_01418_),
    .A1(_18446_),
    .A2(net6091));
 sg13g2_nand3_1 _24801_ (.B(net7109),
    .C(net6091),
    .A(net3561),
    .Y(_17195_));
 sg13g2_o21ai_1 _24802_ (.B1(_17195_),
    .Y(_01419_),
    .A1(_18445_),
    .A2(net6091));
 sg13g2_nand3_1 _24803_ (.B(net7109),
    .C(net6089),
    .A(net2427),
    .Y(_17196_));
 sg13g2_o21ai_1 _24804_ (.B1(_17196_),
    .Y(_01420_),
    .A1(_18444_),
    .A2(net6090));
 sg13g2_nand3_1 _24805_ (.B(net7108),
    .C(net6089),
    .A(net2196),
    .Y(_17197_));
 sg13g2_o21ai_1 _24806_ (.B1(_17197_),
    .Y(_01421_),
    .A1(_18443_),
    .A2(net6090));
 sg13g2_nand3_1 _24807_ (.B(net7108),
    .C(net6089),
    .A(net3065),
    .Y(_17198_));
 sg13g2_o21ai_1 _24808_ (.B1(_17198_),
    .Y(_01422_),
    .A1(_18442_),
    .A2(net6089));
 sg13g2_nand3_1 _24809_ (.B(net7109),
    .C(net6092),
    .A(net2191),
    .Y(_17199_));
 sg13g2_o21ai_1 _24810_ (.B1(_17199_),
    .Y(_01423_),
    .A1(_18441_),
    .A2(net6092));
 sg13g2_nand3_1 _24811_ (.B(net7108),
    .C(net6089),
    .A(net1782),
    .Y(_17200_));
 sg13g2_o21ai_1 _24812_ (.B1(_17200_),
    .Y(_01424_),
    .A1(_18440_),
    .A2(net6089));
 sg13g2_nand3_1 _24813_ (.B(net7108),
    .C(net6089),
    .A(net2578),
    .Y(_17201_));
 sg13g2_o21ai_1 _24814_ (.B1(_17201_),
    .Y(_01425_),
    .A1(_18439_),
    .A2(net6089));
 sg13g2_nand3_1 _24815_ (.B(net7108),
    .C(net6088),
    .A(net3111),
    .Y(_17202_));
 sg13g2_o21ai_1 _24816_ (.B1(_17202_),
    .Y(_01426_),
    .A1(_18438_),
    .A2(net6088));
 sg13g2_nand3_1 _24817_ (.B(net7108),
    .C(net6087),
    .A(net2707),
    .Y(_17203_));
 sg13g2_o21ai_1 _24818_ (.B1(_17203_),
    .Y(_01427_),
    .A1(_18437_),
    .A2(net6088));
 sg13g2_nand3_1 _24819_ (.B(net7102),
    .C(net6088),
    .A(net2074),
    .Y(_17204_));
 sg13g2_o21ai_1 _24820_ (.B1(_17204_),
    .Y(_01428_),
    .A1(_18436_),
    .A2(net6088));
 sg13g2_nand3_1 _24821_ (.B(net7102),
    .C(net6088),
    .A(net2240),
    .Y(_17205_));
 sg13g2_o21ai_1 _24822_ (.B1(_17205_),
    .Y(_01429_),
    .A1(_18435_),
    .A2(net6088));
 sg13g2_nand3_1 _24823_ (.B(net7102),
    .C(net6087),
    .A(net2031),
    .Y(_17206_));
 sg13g2_o21ai_1 _24824_ (.B1(_17206_),
    .Y(_01430_),
    .A1(_18434_),
    .A2(net6087));
 sg13g2_nand3_1 _24825_ (.B(net7102),
    .C(net6087),
    .A(net1982),
    .Y(_17207_));
 sg13g2_o21ai_1 _24826_ (.B1(_17207_),
    .Y(_01431_),
    .A1(_18433_),
    .A2(net6087));
 sg13g2_nand3_1 _24827_ (.B(net7102),
    .C(net6087),
    .A(net2095),
    .Y(_17208_));
 sg13g2_o21ai_1 _24828_ (.B1(_17208_),
    .Y(_01432_),
    .A1(_18432_),
    .A2(net6087));
 sg13g2_nand3_1 _24829_ (.B(net7102),
    .C(net6090),
    .A(net2654),
    .Y(_17209_));
 sg13g2_o21ai_1 _24830_ (.B1(_17209_),
    .Y(_01433_),
    .A1(_18431_),
    .A2(net6087));
 sg13g2_nand3_1 _24831_ (.B(net7101),
    .C(net6073),
    .A(net2314),
    .Y(_17210_));
 sg13g2_o21ai_1 _24832_ (.B1(_17210_),
    .Y(_01434_),
    .A1(_18430_),
    .A2(net6073));
 sg13g2_nand3_1 _24833_ (.B(net7101),
    .C(net6073),
    .A(net3374),
    .Y(_17211_));
 sg13g2_o21ai_1 _24834_ (.B1(_17211_),
    .Y(_01435_),
    .A1(_18429_),
    .A2(net6073));
 sg13g2_nand3_1 _24835_ (.B(net7101),
    .C(net6073),
    .A(net2440),
    .Y(_17212_));
 sg13g2_o21ai_1 _24836_ (.B1(_17212_),
    .Y(_01436_),
    .A1(_18428_),
    .A2(net6073));
 sg13g2_nand3_1 _24837_ (.B(net7101),
    .C(net6074),
    .A(net1483),
    .Y(_17213_));
 sg13g2_o21ai_1 _24838_ (.B1(_17213_),
    .Y(_01437_),
    .A1(_18427_),
    .A2(net6073));
 sg13g2_nand3_1 _24839_ (.B(net7101),
    .C(net6074),
    .A(net2687),
    .Y(_17214_));
 sg13g2_o21ai_1 _24840_ (.B1(_17214_),
    .Y(_01438_),
    .A1(_18426_),
    .A2(net6074));
 sg13g2_nand3_1 _24841_ (.B(net7101),
    .C(net6074),
    .A(\u_inv.d_next[189] ),
    .Y(_17215_));
 sg13g2_o21ai_1 _24842_ (.B1(_17215_),
    .Y(_01439_),
    .A1(_18425_),
    .A2(net6074));
 sg13g2_nand3_1 _24843_ (.B(net7101),
    .C(net6074),
    .A(net2548),
    .Y(_17216_));
 sg13g2_o21ai_1 _24844_ (.B1(_17216_),
    .Y(_01440_),
    .A1(_18424_),
    .A2(net6075));
 sg13g2_nand3_1 _24845_ (.B(net7101),
    .C(net6074),
    .A(net3539),
    .Y(_17217_));
 sg13g2_o21ai_1 _24846_ (.B1(_17217_),
    .Y(_01441_),
    .A1(_18423_),
    .A2(net6073));
 sg13g2_nand3_1 _24847_ (.B(net7100),
    .C(net6072),
    .A(net2925),
    .Y(_17218_));
 sg13g2_o21ai_1 _24848_ (.B1(_17218_),
    .Y(_01442_),
    .A1(_18422_),
    .A2(net6072));
 sg13g2_nand3_1 _24849_ (.B(net7100),
    .C(net6071),
    .A(net3547),
    .Y(_17219_));
 sg13g2_o21ai_1 _24850_ (.B1(_17219_),
    .Y(_01443_),
    .A1(_18421_),
    .A2(net6072));
 sg13g2_nand3_1 _24851_ (.B(net7100),
    .C(net6072),
    .A(net2447),
    .Y(_17220_));
 sg13g2_o21ai_1 _24852_ (.B1(_17220_),
    .Y(_01444_),
    .A1(_18420_),
    .A2(net6072));
 sg13g2_nand3_1 _24853_ (.B(net7100),
    .C(net6071),
    .A(net3389),
    .Y(_17221_));
 sg13g2_o21ai_1 _24854_ (.B1(_17221_),
    .Y(_01445_),
    .A1(_18419_),
    .A2(net6072));
 sg13g2_nand3_1 _24855_ (.B(net7100),
    .C(net6071),
    .A(net3549),
    .Y(_17222_));
 sg13g2_o21ai_1 _24856_ (.B1(_17222_),
    .Y(_01446_),
    .A1(_18418_),
    .A2(net6071));
 sg13g2_nand3_1 _24857_ (.B(net7100),
    .C(net6071),
    .A(net3438),
    .Y(_17223_));
 sg13g2_o21ai_1 _24858_ (.B1(_17223_),
    .Y(_01447_),
    .A1(_18417_),
    .A2(net6071));
 sg13g2_nand3_1 _24859_ (.B(net7100),
    .C(net6069),
    .A(net2561),
    .Y(_17224_));
 sg13g2_o21ai_1 _24860_ (.B1(_17224_),
    .Y(_01448_),
    .A1(_18416_),
    .A2(net6069));
 sg13g2_nand3_1 _24861_ (.B(net7100),
    .C(net6071),
    .A(net3027),
    .Y(_17225_));
 sg13g2_o21ai_1 _24862_ (.B1(_17225_),
    .Y(_01449_),
    .A1(_18415_),
    .A2(net6071));
 sg13g2_nand3_1 _24863_ (.B(net7099),
    .C(net6069),
    .A(net2691),
    .Y(_17226_));
 sg13g2_o21ai_1 _24864_ (.B1(_17226_),
    .Y(_01450_),
    .A1(_18414_),
    .A2(net6069));
 sg13g2_nand3_1 _24865_ (.B(net7099),
    .C(net6068),
    .A(net2772),
    .Y(_17227_));
 sg13g2_o21ai_1 _24866_ (.B1(_17227_),
    .Y(_01451_),
    .A1(_18413_),
    .A2(net6068));
 sg13g2_nand3_1 _24867_ (.B(net7099),
    .C(net6068),
    .A(net2693),
    .Y(_17228_));
 sg13g2_o21ai_1 _24868_ (.B1(_17228_),
    .Y(_01452_),
    .A1(_18412_),
    .A2(net6068));
 sg13g2_nand3_1 _24869_ (.B(net7099),
    .C(net6068),
    .A(net3455),
    .Y(_17229_));
 sg13g2_o21ai_1 _24870_ (.B1(_17229_),
    .Y(_01453_),
    .A1(_18411_),
    .A2(net6068));
 sg13g2_nand3_1 _24871_ (.B(net7099),
    .C(net6069),
    .A(net2456),
    .Y(_17230_));
 sg13g2_o21ai_1 _24872_ (.B1(_17230_),
    .Y(_01454_),
    .A1(_18410_),
    .A2(net6068));
 sg13g2_nand3_1 _24873_ (.B(net7099),
    .C(net6070),
    .A(net2824),
    .Y(_17231_));
 sg13g2_o21ai_1 _24874_ (.B1(_17231_),
    .Y(_01455_),
    .A1(_18409_),
    .A2(net6070));
 sg13g2_nand3_1 _24875_ (.B(net7099),
    .C(net6068),
    .A(net2922),
    .Y(_17232_));
 sg13g2_o21ai_1 _24876_ (.B1(_17232_),
    .Y(_01456_),
    .A1(_18408_),
    .A2(net6066));
 sg13g2_nand3_1 _24877_ (.B(net7099),
    .C(net6069),
    .A(net2721),
    .Y(_17233_));
 sg13g2_o21ai_1 _24878_ (.B1(_17233_),
    .Y(_01457_),
    .A1(_18407_),
    .A2(net6069));
 sg13g2_nand3_1 _24879_ (.B(net7092),
    .C(net6066),
    .A(net3425),
    .Y(_17234_));
 sg13g2_o21ai_1 _24880_ (.B1(_17234_),
    .Y(_01458_),
    .A1(_18406_),
    .A2(net6065));
 sg13g2_nand3_1 _24881_ (.B(net7092),
    .C(net6066),
    .A(net3271),
    .Y(_17235_));
 sg13g2_o21ai_1 _24882_ (.B1(_17235_),
    .Y(_01459_),
    .A1(_18405_),
    .A2(net6066));
 sg13g2_nand3_1 _24883_ (.B(net7092),
    .C(net6065),
    .A(net2871),
    .Y(_17236_));
 sg13g2_o21ai_1 _24884_ (.B1(_17236_),
    .Y(_01460_),
    .A1(_18404_),
    .A2(net6065));
 sg13g2_nand3_1 _24885_ (.B(net7092),
    .C(net6065),
    .A(net2787),
    .Y(_17237_));
 sg13g2_o21ai_1 _24886_ (.B1(_17237_),
    .Y(_01461_),
    .A1(_18403_),
    .A2(net6066));
 sg13g2_nand3_1 _24887_ (.B(net7092),
    .C(net6065),
    .A(net2283),
    .Y(_17238_));
 sg13g2_o21ai_1 _24888_ (.B1(_17238_),
    .Y(_01462_),
    .A1(_18402_),
    .A2(net6065));
 sg13g2_nand3_1 _24889_ (.B(net7092),
    .C(net6067),
    .A(net3620),
    .Y(_17239_));
 sg13g2_o21ai_1 _24890_ (.B1(_17239_),
    .Y(_01463_),
    .A1(_18401_),
    .A2(net6067));
 sg13g2_nand3_1 _24891_ (.B(net7091),
    .C(net6067),
    .A(net2920),
    .Y(_17240_));
 sg13g2_o21ai_1 _24892_ (.B1(_17240_),
    .Y(_01464_),
    .A1(_18400_),
    .A2(net6067));
 sg13g2_nand3_1 _24893_ (.B(net7092),
    .C(net6065),
    .A(net3581),
    .Y(_17241_));
 sg13g2_o21ai_1 _24894_ (.B1(_17241_),
    .Y(_01465_),
    .A1(_18399_),
    .A2(net6065));
 sg13g2_nand3_1 _24895_ (.B(net7091),
    .C(net6052),
    .A(net2298),
    .Y(_17242_));
 sg13g2_o21ai_1 _24896_ (.B1(_17242_),
    .Y(_01466_),
    .A1(_18398_),
    .A2(net6053));
 sg13g2_nand3_1 _24897_ (.B(net7091),
    .C(net6052),
    .A(net3506),
    .Y(_17243_));
 sg13g2_o21ai_1 _24898_ (.B1(_17243_),
    .Y(_01467_),
    .A1(_18397_),
    .A2(net6052));
 sg13g2_nand3_1 _24899_ (.B(net7091),
    .C(net6051),
    .A(net2368),
    .Y(_17244_));
 sg13g2_o21ai_1 _24900_ (.B1(_17244_),
    .Y(_01468_),
    .A1(_18396_),
    .A2(net6051));
 sg13g2_nand3_1 _24901_ (.B(net7091),
    .C(net6051),
    .A(net2122),
    .Y(_17245_));
 sg13g2_o21ai_1 _24902_ (.B1(_17245_),
    .Y(_01469_),
    .A1(_18395_),
    .A2(net6051));
 sg13g2_nand3_1 _24903_ (.B(net7091),
    .C(net6051),
    .A(net1987),
    .Y(_17246_));
 sg13g2_o21ai_1 _24904_ (.B1(_17246_),
    .Y(_01470_),
    .A1(_18394_),
    .A2(net6053));
 sg13g2_nand3_1 _24905_ (.B(net7093),
    .C(net6053),
    .A(net2417),
    .Y(_17247_));
 sg13g2_o21ai_1 _24906_ (.B1(_17247_),
    .Y(_01471_),
    .A1(_18393_),
    .A2(net6053));
 sg13g2_nand3_1 _24907_ (.B(net7091),
    .C(net6051),
    .A(net2033),
    .Y(_17248_));
 sg13g2_o21ai_1 _24908_ (.B1(_17248_),
    .Y(_01472_),
    .A1(_18392_),
    .A2(net6051));
 sg13g2_nand3_1 _24909_ (.B(net7091),
    .C(net6051),
    .A(net3070),
    .Y(_17249_));
 sg13g2_o21ai_1 _24910_ (.B1(_17249_),
    .Y(_01473_),
    .A1(_18391_),
    .A2(net6052));
 sg13g2_nand3_1 _24911_ (.B(net7086),
    .C(net6030),
    .A(net2989),
    .Y(_17250_));
 sg13g2_o21ai_1 _24912_ (.B1(_17250_),
    .Y(_01474_),
    .A1(_18390_),
    .A2(net6030));
 sg13g2_nand3_1 _24913_ (.B(net7086),
    .C(net6030),
    .A(net2533),
    .Y(_17251_));
 sg13g2_o21ai_1 _24914_ (.B1(_17251_),
    .Y(_01475_),
    .A1(_18389_),
    .A2(net6030));
 sg13g2_nand3_1 _24915_ (.B(net7086),
    .C(net6049),
    .A(net2591),
    .Y(_17252_));
 sg13g2_o21ai_1 _24916_ (.B1(_17252_),
    .Y(_01476_),
    .A1(_18388_),
    .A2(net6031));
 sg13g2_nand3_1 _24917_ (.B(net7086),
    .C(net6049),
    .A(net3376),
    .Y(_17253_));
 sg13g2_o21ai_1 _24918_ (.B1(_17253_),
    .Y(_01477_),
    .A1(_18387_),
    .A2(net6030));
 sg13g2_nand3_1 _24919_ (.B(net7085),
    .C(net6049),
    .A(net3231),
    .Y(_17254_));
 sg13g2_o21ai_1 _24920_ (.B1(_17254_),
    .Y(_01478_),
    .A1(_18386_),
    .A2(net6049));
 sg13g2_nand3_1 _24921_ (.B(net7085),
    .C(net6050),
    .A(net3445),
    .Y(_17255_));
 sg13g2_o21ai_1 _24922_ (.B1(_17255_),
    .Y(_01479_),
    .A1(_18385_),
    .A2(net6049));
 sg13g2_nand3_1 _24923_ (.B(net7085),
    .C(net6049),
    .A(net2786),
    .Y(_17256_));
 sg13g2_o21ai_1 _24924_ (.B1(_17256_),
    .Y(_01480_),
    .A1(_18384_),
    .A2(net6050));
 sg13g2_nand3_1 _24925_ (.B(net7086),
    .C(net6049),
    .A(net3149),
    .Y(_17257_));
 sg13g2_o21ai_1 _24926_ (.B1(_17257_),
    .Y(_01481_),
    .A1(_18383_),
    .A2(net6049));
 sg13g2_nand3_1 _24927_ (.B(net7085),
    .C(net6048),
    .A(net3273),
    .Y(_17258_));
 sg13g2_o21ai_1 _24928_ (.B1(_17258_),
    .Y(_01482_),
    .A1(_18382_),
    .A2(net6048));
 sg13g2_nand3_1 _24929_ (.B(net7085),
    .C(net6048),
    .A(net3161),
    .Y(_17259_));
 sg13g2_o21ai_1 _24930_ (.B1(_17259_),
    .Y(_01483_),
    .A1(_18381_),
    .A2(net6050));
 sg13g2_nand3_1 _24931_ (.B(net7085),
    .C(net6048),
    .A(net2620),
    .Y(_17260_));
 sg13g2_o21ai_1 _24932_ (.B1(_17260_),
    .Y(_01484_),
    .A1(_18380_),
    .A2(net6048));
 sg13g2_nand3_1 _24933_ (.B(net7085),
    .C(net6048),
    .A(net3593),
    .Y(_17261_));
 sg13g2_o21ai_1 _24934_ (.B1(_17261_),
    .Y(_01485_),
    .A1(_18379_),
    .A2(net6048));
 sg13g2_nand3_1 _24935_ (.B(net7087),
    .C(net6044),
    .A(net2376),
    .Y(_17262_));
 sg13g2_o21ai_1 _24936_ (.B1(_17262_),
    .Y(_01486_),
    .A1(_18378_),
    .A2(net6044));
 sg13g2_nand3_1 _24937_ (.B(net7085),
    .C(net6050),
    .A(net2126),
    .Y(_17263_));
 sg13g2_o21ai_1 _24938_ (.B1(_17263_),
    .Y(_01487_),
    .A1(_18377_),
    .A2(net6048));
 sg13g2_nand3_1 _24939_ (.B(net7087),
    .C(net6045),
    .A(net2671),
    .Y(_17264_));
 sg13g2_o21ai_1 _24940_ (.B1(_17264_),
    .Y(_01488_),
    .A1(_18376_),
    .A2(net6045));
 sg13g2_nand3_1 _24941_ (.B(net7087),
    .C(net6044),
    .A(net2235),
    .Y(_17265_));
 sg13g2_o21ai_1 _24942_ (.B1(_17265_),
    .Y(_01489_),
    .A1(_18375_),
    .A2(net6044));
 sg13g2_nand3_1 _24943_ (.B(net7093),
    .C(net6045),
    .A(net3606),
    .Y(_17266_));
 sg13g2_o21ai_1 _24944_ (.B1(_17266_),
    .Y(_01490_),
    .A1(_18374_),
    .A2(net6043));
 sg13g2_nand3_1 _24945_ (.B(net7093),
    .C(net6046),
    .A(net3575),
    .Y(_17267_));
 sg13g2_o21ai_1 _24946_ (.B1(_17267_),
    .Y(_01491_),
    .A1(_18373_),
    .A2(net6045));
 sg13g2_nand3_1 _24947_ (.B(net7093),
    .C(net6045),
    .A(net3601),
    .Y(_17268_));
 sg13g2_o21ai_1 _24948_ (.B1(_17268_),
    .Y(_01492_),
    .A1(_18372_),
    .A2(net6045));
 sg13g2_nand3_1 _24949_ (.B(net7093),
    .C(net6045),
    .A(net2310),
    .Y(_17269_));
 sg13g2_o21ai_1 _24950_ (.B1(_17269_),
    .Y(_01493_),
    .A1(_18371_),
    .A2(net6045));
 sg13g2_nand3_1 _24951_ (.B(net7087),
    .C(net6043),
    .A(net2633),
    .Y(_17270_));
 sg13g2_o21ai_1 _24952_ (.B1(_17270_),
    .Y(_01494_),
    .A1(_18370_),
    .A2(net6043));
 sg13g2_nand3_1 _24953_ (.B(net7087),
    .C(net6043),
    .A(net7295),
    .Y(_17271_));
 sg13g2_o21ai_1 _24954_ (.B1(_17271_),
    .Y(_01495_),
    .A1(_18369_),
    .A2(net6043));
 sg13g2_nand3_1 _24955_ (.B(net7087),
    .C(net6043),
    .A(net2450),
    .Y(_17272_));
 sg13g2_o21ai_1 _24956_ (.B1(_17272_),
    .Y(_01496_),
    .A1(_18368_),
    .A2(net6043));
 sg13g2_nand3_1 _24957_ (.B(net7087),
    .C(net6046),
    .A(net3017),
    .Y(_17273_));
 sg13g2_o21ai_1 _24958_ (.B1(_17273_),
    .Y(_01497_),
    .A1(_18367_),
    .A2(net6043));
 sg13g2_nand3_1 _24959_ (.B(net7093),
    .C(net6046),
    .A(net3543),
    .Y(_17274_));
 sg13g2_o21ai_1 _24960_ (.B1(_17274_),
    .Y(_01498_),
    .A1(_18366_),
    .A2(net6046));
 sg13g2_nand3_1 _24961_ (.B(net7081),
    .C(net6037),
    .A(net3504),
    .Y(_17275_));
 sg13g2_o21ai_1 _24962_ (.B1(_17275_),
    .Y(_01499_),
    .A1(_18365_),
    .A2(net6036));
 sg13g2_nand3_1 _24963_ (.B(net7081),
    .C(net6036),
    .A(net2880),
    .Y(_17276_));
 sg13g2_o21ai_1 _24964_ (.B1(_17276_),
    .Y(_01500_),
    .A1(_18364_),
    .A2(net6036));
 sg13g2_nand3_1 _24965_ (.B(net7090),
    .C(net6036),
    .A(net2809),
    .Y(_17277_));
 sg13g2_o21ai_1 _24966_ (.B1(_17277_),
    .Y(_01501_),
    .A1(_18363_),
    .A2(net6037));
 sg13g2_nand3_1 _24967_ (.B(net7088),
    .C(net6036),
    .A(net3347),
    .Y(_17278_));
 sg13g2_o21ai_1 _24968_ (.B1(_17278_),
    .Y(_01502_),
    .A1(_18362_),
    .A2(net6036));
 sg13g2_nand3_1 _24969_ (.B(net7088),
    .C(net6036),
    .A(net3493),
    .Y(_17279_));
 sg13g2_o21ai_1 _24970_ (.B1(_17279_),
    .Y(_01503_),
    .A1(_18361_),
    .A2(net6036));
 sg13g2_nand3_1 _24971_ (.B(net7088),
    .C(net6046),
    .A(net2888),
    .Y(_17280_));
 sg13g2_o21ai_1 _24972_ (.B1(_17280_),
    .Y(_01504_),
    .A1(_18360_),
    .A2(net6046));
 sg13g2_nand3_1 _24973_ (.B(net7093),
    .C(net6046),
    .A(net3405),
    .Y(_17281_));
 sg13g2_o21ai_1 _24974_ (.B1(_17281_),
    .Y(_01505_),
    .A1(_18359_),
    .A2(net6046));
 sg13g2_nand3_1 _24975_ (.B(net7090),
    .C(net6059),
    .A(net2988),
    .Y(_17282_));
 sg13g2_o21ai_1 _24976_ (.B1(_17282_),
    .Y(_01506_),
    .A1(_18358_),
    .A2(net6059));
 sg13g2_or2_1 _24977_ (.X(_01507_),
    .B(net6035),
    .A(net2497));
 sg13g2_nor2_1 _24978_ (.A(\u_inv.f_next[1] ),
    .B(net7017),
    .Y(_17283_));
 sg13g2_nor2_1 _24979_ (.A(net2181),
    .B(net6033),
    .Y(_17284_));
 sg13g2_a21oi_1 _24980_ (.A1(net6033),
    .A2(_17283_),
    .Y(_01508_),
    .B1(_17284_));
 sg13g2_nor2_1 _24981_ (.A(\u_inv.f_next[2] ),
    .B(net7017),
    .Y(_17285_));
 sg13g2_nor2_1 _24982_ (.A(net1347),
    .B(net6033),
    .Y(_17286_));
 sg13g2_a21oi_1 _24983_ (.A1(net6033),
    .A2(_17285_),
    .Y(_01509_),
    .B1(_17286_));
 sg13g2_nor2_1 _24984_ (.A(\u_inv.f_next[3] ),
    .B(net7017),
    .Y(_17287_));
 sg13g2_nor2_1 _24985_ (.A(net1722),
    .B(net6033),
    .Y(_17288_));
 sg13g2_a21oi_1 _24986_ (.A1(net6034),
    .A2(_17287_),
    .Y(_01510_),
    .B1(_17288_));
 sg13g2_nand3_1 _24987_ (.B(net7088),
    .C(net6038),
    .A(net1753),
    .Y(_17289_));
 sg13g2_o21ai_1 _24988_ (.B1(_17289_),
    .Y(_01511_),
    .A1(_18191_),
    .A2(net6038));
 sg13g2_nor2_1 _24989_ (.A(\u_inv.f_next[5] ),
    .B(net7021),
    .Y(_17290_));
 sg13g2_nor2_1 _24990_ (.A(net1442),
    .B(net6038),
    .Y(_17291_));
 sg13g2_a21oi_1 _24991_ (.A1(net6038),
    .A2(_17290_),
    .Y(_01512_),
    .B1(_17291_));
 sg13g2_nand3_1 _24992_ (.B(net7088),
    .C(net6039),
    .A(\u_inv.f_next[6] ),
    .Y(_17292_));
 sg13g2_o21ai_1 _24993_ (.B1(_17292_),
    .Y(_01513_),
    .A1(_18192_),
    .A2(net6039));
 sg13g2_nand3_1 _24994_ (.B(net7089),
    .C(net6040),
    .A(net2132),
    .Y(_17293_));
 sg13g2_o21ai_1 _24995_ (.B1(_17293_),
    .Y(_01514_),
    .A1(_18193_),
    .A2(net6040));
 sg13g2_nand3_1 _24996_ (.B(net7089),
    .C(net6040),
    .A(\u_inv.f_next[8] ),
    .Y(_17294_));
 sg13g2_o21ai_1 _24997_ (.B1(_17294_),
    .Y(_01515_),
    .A1(_18194_),
    .A2(net6040));
 sg13g2_nand3_1 _24998_ (.B(net7089),
    .C(net6055),
    .A(\u_inv.f_next[9] ),
    .Y(_17295_));
 sg13g2_o21ai_1 _24999_ (.B1(_17295_),
    .Y(_01516_),
    .A1(_18195_),
    .A2(net6055));
 sg13g2_nor2_1 _25000_ (.A(\u_inv.f_next[10] ),
    .B(net7024),
    .Y(_17296_));
 sg13g2_nor2_1 _25001_ (.A(net2025),
    .B(net6055),
    .Y(_17297_));
 sg13g2_a21oi_1 _25002_ (.A1(net6056),
    .A2(_17296_),
    .Y(_01517_),
    .B1(_17297_));
 sg13g2_nor2_1 _25003_ (.A(net1684),
    .B(net7024),
    .Y(_17298_));
 sg13g2_nor2_1 _25004_ (.A(net2224),
    .B(net6058),
    .Y(_17299_));
 sg13g2_a21oi_1 _25005_ (.A1(net6055),
    .A2(_17298_),
    .Y(_01518_),
    .B1(_17299_));
 sg13g2_nor2_1 _25006_ (.A(\u_inv.f_next[12] ),
    .B(net7025),
    .Y(_17300_));
 sg13g2_nor2_1 _25007_ (.A(net1696),
    .B(net6058),
    .Y(_17301_));
 sg13g2_a21oi_1 _25008_ (.A1(net6058),
    .A2(_17300_),
    .Y(_01519_),
    .B1(_17301_));
 sg13g2_nor2_1 _25009_ (.A(\u_inv.f_next[13] ),
    .B(net7025),
    .Y(_17302_));
 sg13g2_nor2_1 _25010_ (.A(net2839),
    .B(net6058),
    .Y(_17303_));
 sg13g2_a21oi_1 _25011_ (.A1(net6058),
    .A2(_17302_),
    .Y(_01520_),
    .B1(_17303_));
 sg13g2_nor2_1 _25012_ (.A(\u_inv.f_next[14] ),
    .B(net7029),
    .Y(_17304_));
 sg13g2_nor2_1 _25013_ (.A(net1831),
    .B(net6061),
    .Y(_17305_));
 sg13g2_a21oi_1 _25014_ (.A1(net6061),
    .A2(_17304_),
    .Y(_01521_),
    .B1(_17305_));
 sg13g2_nor2_1 _25015_ (.A(net2124),
    .B(net7030),
    .Y(_17306_));
 sg13g2_nor2_1 _25016_ (.A(net2243),
    .B(net6064),
    .Y(_17307_));
 sg13g2_a21oi_1 _25017_ (.A1(net6061),
    .A2(_17306_),
    .Y(_01522_),
    .B1(_17307_));
 sg13g2_nor2_1 _25018_ (.A(\u_inv.f_next[16] ),
    .B(net7031),
    .Y(_17308_));
 sg13g2_nor2_1 _25019_ (.A(net1646),
    .B(net6077),
    .Y(_17309_));
 sg13g2_a21oi_1 _25020_ (.A1(net6077),
    .A2(_17308_),
    .Y(_01523_),
    .B1(_17309_));
 sg13g2_nor2_1 _25021_ (.A(\u_inv.f_next[17] ),
    .B(net7031),
    .Y(_17310_));
 sg13g2_nor2_1 _25022_ (.A(net1717),
    .B(net6077),
    .Y(_17311_));
 sg13g2_a21oi_1 _25023_ (.A1(net6077),
    .A2(_17310_),
    .Y(_01524_),
    .B1(_17311_));
 sg13g2_nor2_1 _25024_ (.A(\u_inv.f_next[18] ),
    .B(net7033),
    .Y(_17312_));
 sg13g2_nor2_1 _25025_ (.A(net2656),
    .B(net6083),
    .Y(_17313_));
 sg13g2_a21oi_1 _25026_ (.A1(net6078),
    .A2(_17312_),
    .Y(_01525_),
    .B1(_17313_));
 sg13g2_nor2_1 _25027_ (.A(net7300),
    .B(net7033),
    .Y(_17314_));
 sg13g2_nor2_1 _25028_ (.A(net3197),
    .B(net6083),
    .Y(_17315_));
 sg13g2_a21oi_1 _25029_ (.A1(net6083),
    .A2(_17314_),
    .Y(_01526_),
    .B1(_17315_));
 sg13g2_nor2_1 _25030_ (.A(\u_inv.f_next[20] ),
    .B(net7033),
    .Y(_17316_));
 sg13g2_nor2_1 _25031_ (.A(net1750),
    .B(net6082),
    .Y(_17317_));
 sg13g2_a21oi_1 _25032_ (.A1(net6082),
    .A2(_17316_),
    .Y(_01527_),
    .B1(_17317_));
 sg13g2_nor2_1 _25033_ (.A(\u_inv.f_next[21] ),
    .B(net7034),
    .Y(_17318_));
 sg13g2_nor2_1 _25034_ (.A(net2169),
    .B(net6082),
    .Y(_17319_));
 sg13g2_a21oi_1 _25035_ (.A1(net6082),
    .A2(_17318_),
    .Y(_01528_),
    .B1(_17319_));
 sg13g2_nor2_1 _25036_ (.A(\u_inv.f_next[22] ),
    .B(net7034),
    .Y(_17320_));
 sg13g2_nor2_1 _25037_ (.A(net2007),
    .B(net6082),
    .Y(_17321_));
 sg13g2_a21oi_1 _25038_ (.A1(net6082),
    .A2(_17320_),
    .Y(_01529_),
    .B1(_17321_));
 sg13g2_nor2_1 _25039_ (.A(\u_inv.f_next[23] ),
    .B(net7036),
    .Y(_17322_));
 sg13g2_nor2_1 _25040_ (.A(net2896),
    .B(net6097),
    .Y(_17323_));
 sg13g2_a21oi_1 _25041_ (.A1(net6097),
    .A2(_17322_),
    .Y(_01530_),
    .B1(_17323_));
 sg13g2_nor2_1 _25042_ (.A(\u_inv.f_next[24] ),
    .B(net7036),
    .Y(_17324_));
 sg13g2_nor2_1 _25043_ (.A(net2076),
    .B(net6097),
    .Y(_17325_));
 sg13g2_a21oi_1 _25044_ (.A1(net6097),
    .A2(_17324_),
    .Y(_01531_),
    .B1(_17325_));
 sg13g2_nor2_1 _25045_ (.A(\u_inv.f_next[25] ),
    .B(net7039),
    .Y(_17326_));
 sg13g2_nor2_1 _25046_ (.A(net3289),
    .B(net6103),
    .Y(_17327_));
 sg13g2_a21oi_1 _25047_ (.A1(net6103),
    .A2(_17326_),
    .Y(_01532_),
    .B1(_17327_));
 sg13g2_nor2_1 _25048_ (.A(\u_inv.f_next[26] ),
    .B(net7041),
    .Y(_17328_));
 sg13g2_nor2_1 _25049_ (.A(net1588),
    .B(net6104),
    .Y(_17329_));
 sg13g2_a21oi_1 _25050_ (.A1(net6104),
    .A2(_17328_),
    .Y(_01533_),
    .B1(_17329_));
 sg13g2_nor2_1 _25051_ (.A(\u_inv.f_next[27] ),
    .B(net7045),
    .Y(_17330_));
 sg13g2_nor2_1 _25052_ (.A(net1920),
    .B(net6104),
    .Y(_17331_));
 sg13g2_a21oi_1 _25053_ (.A1(net6104),
    .A2(_17330_),
    .Y(_01534_),
    .B1(_17331_));
 sg13g2_nor2_1 _25054_ (.A(\u_inv.f_next[28] ),
    .B(net7045),
    .Y(_17332_));
 sg13g2_nor2_1 _25055_ (.A(net2244),
    .B(net6119),
    .Y(_17333_));
 sg13g2_a21oi_1 _25056_ (.A1(net6119),
    .A2(_17332_),
    .Y(_01535_),
    .B1(_17333_));
 sg13g2_nor2_1 _25057_ (.A(\u_inv.f_next[29] ),
    .B(net7047),
    .Y(_17334_));
 sg13g2_nor2_1 _25058_ (.A(net3042),
    .B(net6119),
    .Y(_17335_));
 sg13g2_a21oi_1 _25059_ (.A1(net6119),
    .A2(_17334_),
    .Y(_01536_),
    .B1(_17335_));
 sg13g2_nor2_1 _25060_ (.A(\u_inv.f_next[30] ),
    .B(net7045),
    .Y(_17336_));
 sg13g2_nor2_1 _25061_ (.A(net1708),
    .B(net6125),
    .Y(_17337_));
 sg13g2_a21oi_1 _25062_ (.A1(net6120),
    .A2(_17336_),
    .Y(_01537_),
    .B1(_17337_));
 sg13g2_nor2_1 _25063_ (.A(\u_inv.f_next[31] ),
    .B(net7045),
    .Y(_17338_));
 sg13g2_nor2_1 _25064_ (.A(net2393),
    .B(net6120),
    .Y(_17339_));
 sg13g2_a21oi_1 _25065_ (.A1(net6120),
    .A2(_17338_),
    .Y(_01538_),
    .B1(_17339_));
 sg13g2_nand3_1 _25066_ (.B(net7123),
    .C(net6126),
    .A(net2760),
    .Y(_17340_));
 sg13g2_o21ai_1 _25067_ (.B1(_17340_),
    .Y(_01539_),
    .A1(_18200_),
    .A2(net6126));
 sg13g2_nor2_1 _25068_ (.A(\u_inv.f_next[33] ),
    .B(net7048),
    .Y(_17341_));
 sg13g2_nor2_1 _25069_ (.A(net2055),
    .B(net6126),
    .Y(_17342_));
 sg13g2_a21oi_1 _25070_ (.A1(net6126),
    .A2(_17341_),
    .Y(_01540_),
    .B1(_17342_));
 sg13g2_nor2_1 _25071_ (.A(\u_inv.f_next[34] ),
    .B(net7048),
    .Y(_17343_));
 sg13g2_nor2_1 _25072_ (.A(net1486),
    .B(net6126),
    .Y(_17344_));
 sg13g2_a21oi_1 _25073_ (.A1(net6126),
    .A2(_17343_),
    .Y(_01541_),
    .B1(_17344_));
 sg13g2_nor2_1 _25074_ (.A(\u_inv.f_next[35] ),
    .B(net7049),
    .Y(_17345_));
 sg13g2_nor2_1 _25075_ (.A(net2070),
    .B(net6127),
    .Y(_17346_));
 sg13g2_a21oi_1 _25076_ (.A1(net6127),
    .A2(_17345_),
    .Y(_01542_),
    .B1(_17346_));
 sg13g2_nor2_1 _25077_ (.A(\u_inv.f_next[36] ),
    .B(net7049),
    .Y(_17347_));
 sg13g2_nor2_1 _25078_ (.A(net1579),
    .B(net6127),
    .Y(_17348_));
 sg13g2_a21oi_1 _25079_ (.A1(net6128),
    .A2(_17347_),
    .Y(_01543_),
    .B1(_17348_));
 sg13g2_nor2_1 _25080_ (.A(\u_inv.f_next[37] ),
    .B(net7049),
    .Y(_17349_));
 sg13g2_nor2_1 _25081_ (.A(net1353),
    .B(net6127),
    .Y(_17350_));
 sg13g2_a21oi_1 _25082_ (.A1(net6128),
    .A2(_17349_),
    .Y(_01544_),
    .B1(_17350_));
 sg13g2_nor2_1 _25083_ (.A(\u_inv.f_next[38] ),
    .B(net7048),
    .Y(_17351_));
 sg13g2_nor2_1 _25084_ (.A(net1654),
    .B(net6127),
    .Y(_17352_));
 sg13g2_a21oi_1 _25085_ (.A1(net6127),
    .A2(_17351_),
    .Y(_01545_),
    .B1(_17352_));
 sg13g2_nor2_1 _25086_ (.A(\u_inv.f_next[39] ),
    .B(net7049),
    .Y(_17353_));
 sg13g2_nor2_1 _25087_ (.A(net2035),
    .B(net6127),
    .Y(_17354_));
 sg13g2_a21oi_1 _25088_ (.A1(net6127),
    .A2(_17353_),
    .Y(_01546_),
    .B1(_17354_));
 sg13g2_nor2_1 _25089_ (.A(\u_inv.f_next[40] ),
    .B(net7053),
    .Y(_17355_));
 sg13g2_nor2_1 _25090_ (.A(net2117),
    .B(net6145),
    .Y(_17356_));
 sg13g2_a21oi_1 _25091_ (.A1(net6145),
    .A2(_17355_),
    .Y(_01547_),
    .B1(_17356_));
 sg13g2_nor2_1 _25092_ (.A(net2439),
    .B(net7053),
    .Y(_17357_));
 sg13g2_nor2_1 _25093_ (.A(net2659),
    .B(net6145),
    .Y(_17358_));
 sg13g2_a21oi_1 _25094_ (.A1(net6145),
    .A2(_17357_),
    .Y(_01548_),
    .B1(_17358_));
 sg13g2_nor2_1 _25095_ (.A(\u_inv.f_next[42] ),
    .B(net7054),
    .Y(_17359_));
 sg13g2_nor2_1 _25096_ (.A(net2685),
    .B(net6144),
    .Y(_17360_));
 sg13g2_a21oi_1 _25097_ (.A1(net6144),
    .A2(_17359_),
    .Y(_01549_),
    .B1(_17360_));
 sg13g2_nor2_1 _25098_ (.A(\u_inv.f_next[43] ),
    .B(net7053),
    .Y(_17361_));
 sg13g2_nor2_1 _25099_ (.A(net2941),
    .B(net6145),
    .Y(_17362_));
 sg13g2_a21oi_1 _25100_ (.A1(net6145),
    .A2(_17361_),
    .Y(_01550_),
    .B1(_17362_));
 sg13g2_nor2_1 _25101_ (.A(\u_inv.f_next[44] ),
    .B(net7054),
    .Y(_17363_));
 sg13g2_nor2_1 _25102_ (.A(net1444),
    .B(net6144),
    .Y(_17364_));
 sg13g2_a21oi_1 _25103_ (.A1(net6144),
    .A2(_17363_),
    .Y(_01551_),
    .B1(_17364_));
 sg13g2_nor2_1 _25104_ (.A(net1284),
    .B(net7054),
    .Y(_17365_));
 sg13g2_nor2_1 _25105_ (.A(net2137),
    .B(net6143),
    .Y(_17366_));
 sg13g2_a21oi_1 _25106_ (.A1(net6143),
    .A2(_17365_),
    .Y(_01552_),
    .B1(_17366_));
 sg13g2_nor2_1 _25107_ (.A(\u_inv.f_next[46] ),
    .B(net7058),
    .Y(_17367_));
 sg13g2_nor2_1 _25108_ (.A(net2079),
    .B(net6150),
    .Y(_17368_));
 sg13g2_a21oi_1 _25109_ (.A1(net6150),
    .A2(_17367_),
    .Y(_01553_),
    .B1(_17368_));
 sg13g2_nor2_1 _25110_ (.A(\u_inv.f_next[47] ),
    .B(net7058),
    .Y(_17369_));
 sg13g2_nor2_1 _25111_ (.A(net2598),
    .B(net6150),
    .Y(_17370_));
 sg13g2_a21oi_1 _25112_ (.A1(net6150),
    .A2(_17369_),
    .Y(_01554_),
    .B1(_17370_));
 sg13g2_nor2_1 _25113_ (.A(\u_inv.f_next[48] ),
    .B(net7053),
    .Y(_17371_));
 sg13g2_nor2_1 _25114_ (.A(net1506),
    .B(net6143),
    .Y(_17372_));
 sg13g2_a21oi_1 _25115_ (.A1(net6143),
    .A2(_17371_),
    .Y(_01555_),
    .B1(_17372_));
 sg13g2_nor2_1 _25116_ (.A(net1669),
    .B(net7054),
    .Y(_17373_));
 sg13g2_nor2_1 _25117_ (.A(net2030),
    .B(net6143),
    .Y(_17374_));
 sg13g2_a21oi_1 _25118_ (.A1(net6143),
    .A2(_17373_),
    .Y(_01556_),
    .B1(_17374_));
 sg13g2_nor2_1 _25119_ (.A(\u_inv.f_next[50] ),
    .B(net7053),
    .Y(_17375_));
 sg13g2_nor2_1 _25120_ (.A(net1894),
    .B(net6143),
    .Y(_17376_));
 sg13g2_a21oi_1 _25121_ (.A1(net6143),
    .A2(_17375_),
    .Y(_01557_),
    .B1(_17376_));
 sg13g2_nor2_1 _25122_ (.A(\u_inv.f_next[51] ),
    .B(net7058),
    .Y(_17377_));
 sg13g2_nor2_1 _25123_ (.A(net2344),
    .B(net6152),
    .Y(_17378_));
 sg13g2_a21oi_1 _25124_ (.A1(net6150),
    .A2(_17377_),
    .Y(_01558_),
    .B1(_17378_));
 sg13g2_nor2_1 _25125_ (.A(\u_inv.f_next[52] ),
    .B(net7058),
    .Y(_17379_));
 sg13g2_nor2_1 _25126_ (.A(net2453),
    .B(net6150),
    .Y(_17380_));
 sg13g2_a21oi_1 _25127_ (.A1(net6150),
    .A2(_17379_),
    .Y(_01559_),
    .B1(_17380_));
 sg13g2_nor2_1 _25128_ (.A(\u_inv.f_next[53] ),
    .B(net7059),
    .Y(_17381_));
 sg13g2_nor2_1 _25129_ (.A(net2841),
    .B(net6151),
    .Y(_17382_));
 sg13g2_a21oi_1 _25130_ (.A1(net6151),
    .A2(_17381_),
    .Y(_01560_),
    .B1(_17382_));
 sg13g2_nor2_1 _25131_ (.A(\u_inv.f_next[54] ),
    .B(net7065),
    .Y(_17383_));
 sg13g2_nor2_1 _25132_ (.A(net2875),
    .B(net6166),
    .Y(_17384_));
 sg13g2_a21oi_1 _25133_ (.A1(net6166),
    .A2(_17383_),
    .Y(_01561_),
    .B1(_17384_));
 sg13g2_nor2_1 _25134_ (.A(\u_inv.f_next[55] ),
    .B(net7059),
    .Y(_17385_));
 sg13g2_nor2_1 _25135_ (.A(net1785),
    .B(net6151),
    .Y(_17386_));
 sg13g2_a21oi_1 _25136_ (.A1(net6151),
    .A2(_17385_),
    .Y(_01562_),
    .B1(_17386_));
 sg13g2_nor2_1 _25137_ (.A(\u_inv.f_next[56] ),
    .B(net7065),
    .Y(_17387_));
 sg13g2_nor2_1 _25138_ (.A(net2425),
    .B(net6165),
    .Y(_17388_));
 sg13g2_a21oi_1 _25139_ (.A1(net6166),
    .A2(_17387_),
    .Y(_01563_),
    .B1(_17388_));
 sg13g2_nor2_1 _25140_ (.A(\u_inv.f_next[57] ),
    .B(net7066),
    .Y(_17389_));
 sg13g2_nor2_1 _25141_ (.A(net3109),
    .B(net6152),
    .Y(_17390_));
 sg13g2_a21oi_1 _25142_ (.A1(net6152),
    .A2(_17389_),
    .Y(_01564_),
    .B1(_17390_));
 sg13g2_nor2_1 _25143_ (.A(\u_inv.f_next[58] ),
    .B(net7058),
    .Y(_17391_));
 sg13g2_nor2_1 _25144_ (.A(net2388),
    .B(net6151),
    .Y(_17392_));
 sg13g2_a21oi_1 _25145_ (.A1(net6151),
    .A2(_17391_),
    .Y(_01565_),
    .B1(_17392_));
 sg13g2_nor2_1 _25146_ (.A(\u_inv.f_next[59] ),
    .B(net7065),
    .Y(_17393_));
 sg13g2_nor2_1 _25147_ (.A(net1865),
    .B(net6165),
    .Y(_17394_));
 sg13g2_a21oi_1 _25148_ (.A1(net6165),
    .A2(_17393_),
    .Y(_01566_),
    .B1(_17394_));
 sg13g2_nor2_1 _25149_ (.A(\u_inv.f_next[60] ),
    .B(net7065),
    .Y(_17395_));
 sg13g2_nor2_1 _25150_ (.A(net1687),
    .B(net6165),
    .Y(_17396_));
 sg13g2_a21oi_1 _25151_ (.A1(net6165),
    .A2(_17395_),
    .Y(_01567_),
    .B1(_17396_));
 sg13g2_nor2_1 _25152_ (.A(\u_inv.f_next[61] ),
    .B(net7065),
    .Y(_17397_));
 sg13g2_nor2_1 _25153_ (.A(net2198),
    .B(net6165),
    .Y(_17398_));
 sg13g2_a21oi_1 _25154_ (.A1(net6165),
    .A2(_17397_),
    .Y(_01568_),
    .B1(_17398_));
 sg13g2_nor2_1 _25155_ (.A(\u_inv.f_next[62] ),
    .B(net7065),
    .Y(_17399_));
 sg13g2_nor2_1 _25156_ (.A(net1949),
    .B(net6167),
    .Y(_17400_));
 sg13g2_a21oi_1 _25157_ (.A1(net6167),
    .A2(_17399_),
    .Y(_01569_),
    .B1(_17400_));
 sg13g2_nor2_1 _25158_ (.A(\u_inv.f_next[63] ),
    .B(net7065),
    .Y(_17401_));
 sg13g2_nor2_1 _25159_ (.A(net2810),
    .B(net6165),
    .Y(_17402_));
 sg13g2_a21oi_1 _25160_ (.A1(net6151),
    .A2(_17401_),
    .Y(_01570_),
    .B1(_17402_));
 sg13g2_nor2_1 _25161_ (.A(\u_inv.f_next[64] ),
    .B(net7067),
    .Y(_17403_));
 sg13g2_nor2_1 _25162_ (.A(net1857),
    .B(net6167),
    .Y(_17404_));
 sg13g2_a21oi_1 _25163_ (.A1(net6167),
    .A2(_17403_),
    .Y(_01571_),
    .B1(_17404_));
 sg13g2_nor2_1 _25164_ (.A(\u_inv.f_next[65] ),
    .B(net7067),
    .Y(_17405_));
 sg13g2_nor2_1 _25165_ (.A(net2295),
    .B(net6166),
    .Y(_17406_));
 sg13g2_a21oi_1 _25166_ (.A1(net6166),
    .A2(_17405_),
    .Y(_01572_),
    .B1(_17406_));
 sg13g2_nor2_1 _25167_ (.A(\u_inv.f_next[66] ),
    .B(net7067),
    .Y(_17407_));
 sg13g2_nor2_1 _25168_ (.A(net2341),
    .B(net6167),
    .Y(_17408_));
 sg13g2_a21oi_1 _25169_ (.A1(net6167),
    .A2(_17407_),
    .Y(_01573_),
    .B1(_17408_));
 sg13g2_nor2_1 _25170_ (.A(\u_inv.f_next[67] ),
    .B(net7068),
    .Y(_17409_));
 sg13g2_nor2_1 _25171_ (.A(net2113),
    .B(net6170),
    .Y(_17410_));
 sg13g2_a21oi_1 _25172_ (.A1(net6170),
    .A2(_17409_),
    .Y(_01574_),
    .B1(_17410_));
 sg13g2_nor2_1 _25173_ (.A(\u_inv.f_next[68] ),
    .B(net7070),
    .Y(_17411_));
 sg13g2_nor2_1 _25174_ (.A(net2501),
    .B(net6172),
    .Y(_17412_));
 sg13g2_a21oi_1 _25175_ (.A1(net6170),
    .A2(_17411_),
    .Y(_01575_),
    .B1(_17412_));
 sg13g2_nor2_1 _25176_ (.A(\u_inv.f_next[69] ),
    .B(net7070),
    .Y(_17413_));
 sg13g2_nor2_1 _25177_ (.A(net3344),
    .B(net6171),
    .Y(_17414_));
 sg13g2_a21oi_1 _25178_ (.A1(net6171),
    .A2(_17413_),
    .Y(_01576_),
    .B1(_17414_));
 sg13g2_nor2_1 _25179_ (.A(\u_inv.f_next[70] ),
    .B(net7068),
    .Y(_17415_));
 sg13g2_nor2_1 _25180_ (.A(net1900),
    .B(net6170),
    .Y(_17416_));
 sg13g2_a21oi_1 _25181_ (.A1(net6170),
    .A2(_17415_),
    .Y(_01577_),
    .B1(_17416_));
 sg13g2_nor2_1 _25182_ (.A(\u_inv.f_next[71] ),
    .B(net7068),
    .Y(_17417_));
 sg13g2_nor2_1 _25183_ (.A(net2776),
    .B(net6170),
    .Y(_17418_));
 sg13g2_a21oi_1 _25184_ (.A1(net6170),
    .A2(_17417_),
    .Y(_01578_),
    .B1(_17418_));
 sg13g2_nor2_1 _25185_ (.A(\u_inv.f_next[72] ),
    .B(net7070),
    .Y(_17419_));
 sg13g2_nor2_1 _25186_ (.A(net1586),
    .B(net6172),
    .Y(_17420_));
 sg13g2_a21oi_1 _25187_ (.A1(net6172),
    .A2(_17419_),
    .Y(_01579_),
    .B1(_17420_));
 sg13g2_nor2_1 _25188_ (.A(\u_inv.f_next[73] ),
    .B(net7070),
    .Y(_17421_));
 sg13g2_nor2_1 _25189_ (.A(net1947),
    .B(net6171),
    .Y(_17422_));
 sg13g2_a21oi_1 _25190_ (.A1(net6171),
    .A2(_17421_),
    .Y(_01580_),
    .B1(_17422_));
 sg13g2_nor2_1 _25191_ (.A(\u_inv.f_next[74] ),
    .B(net7070),
    .Y(_17423_));
 sg13g2_nor2_1 _25192_ (.A(net2738),
    .B(net6172),
    .Y(_17424_));
 sg13g2_a21oi_1 _25193_ (.A1(net6172),
    .A2(_17423_),
    .Y(_01581_),
    .B1(_17424_));
 sg13g2_nor2_1 _25194_ (.A(\u_inv.f_next[75] ),
    .B(net7070),
    .Y(_17425_));
 sg13g2_nor2_1 _25195_ (.A(net3004),
    .B(net6171),
    .Y(_17426_));
 sg13g2_a21oi_1 _25196_ (.A1(net6171),
    .A2(_17425_),
    .Y(_01582_),
    .B1(_17426_));
 sg13g2_nor2_1 _25197_ (.A(\u_inv.f_next[76] ),
    .B(net7070),
    .Y(_17427_));
 sg13g2_nor2_1 _25198_ (.A(net2415),
    .B(net6171),
    .Y(_17428_));
 sg13g2_a21oi_1 _25199_ (.A1(net6171),
    .A2(_17427_),
    .Y(_01583_),
    .B1(_17428_));
 sg13g2_nor2_1 _25200_ (.A(\u_inv.f_next[77] ),
    .B(net7071),
    .Y(_17429_));
 sg13g2_nor2_1 _25201_ (.A(net1665),
    .B(net6173),
    .Y(_17430_));
 sg13g2_a21oi_1 _25202_ (.A1(net6173),
    .A2(_17429_),
    .Y(_01584_),
    .B1(_17430_));
 sg13g2_nor2_1 _25203_ (.A(\u_inv.f_next[78] ),
    .B(net7071),
    .Y(_17431_));
 sg13g2_nor2_1 _25204_ (.A(net2194),
    .B(net6173),
    .Y(_17432_));
 sg13g2_a21oi_1 _25205_ (.A1(net6173),
    .A2(_17431_),
    .Y(_01585_),
    .B1(_17432_));
 sg13g2_nor2_1 _25206_ (.A(\u_inv.f_next[79] ),
    .B(net7070),
    .Y(_17433_));
 sg13g2_nor2_1 _25207_ (.A(net2364),
    .B(net6174),
    .Y(_17434_));
 sg13g2_a21oi_1 _25208_ (.A1(net6174),
    .A2(_17433_),
    .Y(_01586_),
    .B1(_17434_));
 sg13g2_nor2_1 _25209_ (.A(\u_inv.f_next[80] ),
    .B(net7069),
    .Y(_17435_));
 sg13g2_nor2_1 _25210_ (.A(net2129),
    .B(net6170),
    .Y(_17436_));
 sg13g2_a21oi_1 _25211_ (.A1(net6175),
    .A2(_17435_),
    .Y(_01587_),
    .B1(_17436_));
 sg13g2_nor2_1 _25212_ (.A(\u_inv.f_next[81] ),
    .B(net7071),
    .Y(_17437_));
 sg13g2_nor2_1 _25213_ (.A(net2460),
    .B(net6173),
    .Y(_17438_));
 sg13g2_a21oi_1 _25214_ (.A1(net6173),
    .A2(_17437_),
    .Y(_01588_),
    .B1(_17438_));
 sg13g2_nor2_1 _25215_ (.A(\u_inv.f_next[82] ),
    .B(net7073),
    .Y(_17439_));
 sg13g2_nor2_1 _25216_ (.A(net2107),
    .B(net6173),
    .Y(_17440_));
 sg13g2_a21oi_1 _25217_ (.A1(net6173),
    .A2(_17439_),
    .Y(_01589_),
    .B1(_17440_));
 sg13g2_nor2_1 _25218_ (.A(\u_inv.f_next[83] ),
    .B(net7073),
    .Y(_17441_));
 sg13g2_nor2_1 _25219_ (.A(net1711),
    .B(net6176),
    .Y(_17442_));
 sg13g2_a21oi_1 _25220_ (.A1(net6176),
    .A2(_17441_),
    .Y(_01590_),
    .B1(_17442_));
 sg13g2_nor2_1 _25221_ (.A(\u_inv.f_next[84] ),
    .B(net7073),
    .Y(_17443_));
 sg13g2_nor2_1 _25222_ (.A(net3093),
    .B(net6174),
    .Y(_17444_));
 sg13g2_a21oi_1 _25223_ (.A1(net6174),
    .A2(_17443_),
    .Y(_01591_),
    .B1(_17444_));
 sg13g2_nor2_1 _25224_ (.A(\u_inv.f_next[85] ),
    .B(net7073),
    .Y(_17445_));
 sg13g2_nor2_1 _25225_ (.A(net2395),
    .B(net6178),
    .Y(_17446_));
 sg13g2_a21oi_1 _25226_ (.A1(net6178),
    .A2(_17445_),
    .Y(_01592_),
    .B1(_17446_));
 sg13g2_nor2_1 _25227_ (.A(\u_inv.f_next[86] ),
    .B(net7073),
    .Y(_17447_));
 sg13g2_nor2_1 _25228_ (.A(net2740),
    .B(net6176),
    .Y(_17448_));
 sg13g2_a21oi_1 _25229_ (.A1(net6176),
    .A2(_17447_),
    .Y(_01593_),
    .B1(_17448_));
 sg13g2_nor2_1 _25230_ (.A(net1576),
    .B(net7072),
    .Y(_17449_));
 sg13g2_nor2_1 _25231_ (.A(net2050),
    .B(net6181),
    .Y(_17450_));
 sg13g2_a21oi_1 _25232_ (.A1(net6181),
    .A2(_17449_),
    .Y(_01594_),
    .B1(_17450_));
 sg13g2_nor2_1 _25233_ (.A(\u_inv.f_next[88] ),
    .B(net7074),
    .Y(_17451_));
 sg13g2_nor2_1 _25234_ (.A(net2091),
    .B(net6176),
    .Y(_17452_));
 sg13g2_a21oi_1 _25235_ (.A1(net6176),
    .A2(_17451_),
    .Y(_01595_),
    .B1(_17452_));
 sg13g2_nor2_1 _25236_ (.A(\u_inv.f_next[89] ),
    .B(net7074),
    .Y(_17453_));
 sg13g2_nor2_1 _25237_ (.A(net3068),
    .B(net6180),
    .Y(_17454_));
 sg13g2_a21oi_1 _25238_ (.A1(net6180),
    .A2(_17453_),
    .Y(_01596_),
    .B1(_17454_));
 sg13g2_nor2_1 _25239_ (.A(\u_inv.f_next[90] ),
    .B(net7074),
    .Y(_17455_));
 sg13g2_nor2_1 _25240_ (.A(net2023),
    .B(net6179),
    .Y(_17456_));
 sg13g2_a21oi_1 _25241_ (.A1(net6179),
    .A2(_17455_),
    .Y(_01597_),
    .B1(_17456_));
 sg13g2_nor2_1 _25242_ (.A(\u_inv.f_next[91] ),
    .B(net7074),
    .Y(_17457_));
 sg13g2_nor2_1 _25243_ (.A(net2359),
    .B(net6179),
    .Y(_17458_));
 sg13g2_a21oi_1 _25244_ (.A1(net6179),
    .A2(_17457_),
    .Y(_01598_),
    .B1(_17458_));
 sg13g2_nor2_1 _25245_ (.A(\u_inv.f_next[92] ),
    .B(net7073),
    .Y(_17459_));
 sg13g2_nor2_1 _25246_ (.A(net1632),
    .B(net6176),
    .Y(_17460_));
 sg13g2_a21oi_1 _25247_ (.A1(net6176),
    .A2(_17459_),
    .Y(_01599_),
    .B1(_17460_));
 sg13g2_nor2_1 _25248_ (.A(\u_inv.f_next[93] ),
    .B(net7073),
    .Y(_17461_));
 sg13g2_nor2_1 _25249_ (.A(net2027),
    .B(net6177),
    .Y(_17462_));
 sg13g2_a21oi_1 _25250_ (.A1(net6177),
    .A2(_17461_),
    .Y(_01600_),
    .B1(_17462_));
 sg13g2_nor2_1 _25251_ (.A(\u_inv.f_next[94] ),
    .B(net7073),
    .Y(_17463_));
 sg13g2_nor2_1 _25252_ (.A(net2220),
    .B(net6177),
    .Y(_17464_));
 sg13g2_a21oi_1 _25253_ (.A1(net6177),
    .A2(_17463_),
    .Y(_01601_),
    .B1(_17464_));
 sg13g2_nor2_1 _25254_ (.A(\u_inv.f_next[95] ),
    .B(net7074),
    .Y(_17465_));
 sg13g2_nor2_1 _25255_ (.A(net2214),
    .B(net6177),
    .Y(_17466_));
 sg13g2_a21oi_1 _25256_ (.A1(net6177),
    .A2(_17465_),
    .Y(_01602_),
    .B1(_17466_));
 sg13g2_nor2_1 _25257_ (.A(\u_inv.f_next[96] ),
    .B(net7076),
    .Y(_17467_));
 sg13g2_nor2_1 _25258_ (.A(net2491),
    .B(net6168),
    .Y(_17468_));
 sg13g2_a21oi_1 _25259_ (.A1(net6168),
    .A2(_17467_),
    .Y(_01603_),
    .B1(_17468_));
 sg13g2_nor2_1 _25260_ (.A(\u_inv.f_next[97] ),
    .B(net7067),
    .Y(_17469_));
 sg13g2_nor2_1 _25261_ (.A(net2072),
    .B(net6168),
    .Y(_17470_));
 sg13g2_a21oi_1 _25262_ (.A1(net6168),
    .A2(_17469_),
    .Y(_01604_),
    .B1(_17470_));
 sg13g2_nor2_1 _25263_ (.A(\u_inv.f_next[98] ),
    .B(net7061),
    .Y(_17471_));
 sg13g2_nor2_1 _25264_ (.A(net2683),
    .B(net6153),
    .Y(_17472_));
 sg13g2_a21oi_1 _25265_ (.A1(net6154),
    .A2(_17471_),
    .Y(_01605_),
    .B1(_17472_));
 sg13g2_nor2_1 _25266_ (.A(\u_inv.f_next[99] ),
    .B(net7061),
    .Y(_17473_));
 sg13g2_nor2_1 _25267_ (.A(net2222),
    .B(net6154),
    .Y(_17474_));
 sg13g2_a21oi_1 _25268_ (.A1(net6154),
    .A2(_17473_),
    .Y(_01606_),
    .B1(_17474_));
 sg13g2_nor2_1 _25269_ (.A(\u_inv.f_next[100] ),
    .B(net7060),
    .Y(_17475_));
 sg13g2_nor2_1 _25270_ (.A(net2200),
    .B(net6151),
    .Y(_17476_));
 sg13g2_a21oi_1 _25271_ (.A1(net6150),
    .A2(_17475_),
    .Y(_01607_),
    .B1(_17476_));
 sg13g2_nor2_1 _25272_ (.A(\u_inv.f_next[101] ),
    .B(net7060),
    .Y(_17477_));
 sg13g2_nor2_1 _25273_ (.A(net2241),
    .B(net6153),
    .Y(_17478_));
 sg13g2_a21oi_1 _25274_ (.A1(net6153),
    .A2(_17477_),
    .Y(_01608_),
    .B1(_17478_));
 sg13g2_nor2_1 _25275_ (.A(\u_inv.f_next[102] ),
    .B(net7061),
    .Y(_17479_));
 sg13g2_nor2_1 _25276_ (.A(net2405),
    .B(net6154),
    .Y(_17480_));
 sg13g2_a21oi_1 _25277_ (.A1(net6154),
    .A2(_17479_),
    .Y(_01609_),
    .B1(_17480_));
 sg13g2_nor2_1 _25278_ (.A(\u_inv.f_next[103] ),
    .B(net7060),
    .Y(_17481_));
 sg13g2_nor2_1 _25279_ (.A(net2812),
    .B(net6153),
    .Y(_17482_));
 sg13g2_a21oi_1 _25280_ (.A1(net6153),
    .A2(_17481_),
    .Y(_01610_),
    .B1(_17482_));
 sg13g2_nor2_1 _25281_ (.A(\u_inv.f_next[104] ),
    .B(net7056),
    .Y(_17483_));
 sg13g2_nor2_1 _25282_ (.A(net1642),
    .B(net6148),
    .Y(_17484_));
 sg13g2_a21oi_1 _25283_ (.A1(net6148),
    .A2(_17483_),
    .Y(_01611_),
    .B1(_17484_));
 sg13g2_nor2_1 _25284_ (.A(net1419),
    .B(net7060),
    .Y(_17485_));
 sg13g2_nor2_1 _25285_ (.A(net2573),
    .B(net6153),
    .Y(_17486_));
 sg13g2_a21oi_1 _25286_ (.A1(net6153),
    .A2(_17485_),
    .Y(_01612_),
    .B1(_17486_));
 sg13g2_nor2_1 _25287_ (.A(\u_inv.f_next[106] ),
    .B(net7056),
    .Y(_17487_));
 sg13g2_nor2_1 _25288_ (.A(net2917),
    .B(net6148),
    .Y(_17488_));
 sg13g2_a21oi_1 _25289_ (.A1(net6148),
    .A2(_17487_),
    .Y(_01613_),
    .B1(_17488_));
 sg13g2_nor2_1 _25290_ (.A(\u_inv.f_next[107] ),
    .B(net7056),
    .Y(_17489_));
 sg13g2_nor2_1 _25291_ (.A(net1854),
    .B(net6146),
    .Y(_17490_));
 sg13g2_a21oi_1 _25292_ (.A1(net6146),
    .A2(_17489_),
    .Y(_01614_),
    .B1(_17490_));
 sg13g2_nor2_1 _25293_ (.A(\u_inv.f_next[108] ),
    .B(net7056),
    .Y(_17491_));
 sg13g2_nor2_1 _25294_ (.A(net2709),
    .B(net6147),
    .Y(_17492_));
 sg13g2_a21oi_1 _25295_ (.A1(net6147),
    .A2(_17491_),
    .Y(_01615_),
    .B1(_17492_));
 sg13g2_nor2_1 _25296_ (.A(\u_inv.f_next[109] ),
    .B(net7057),
    .Y(_17493_));
 sg13g2_nor2_1 _25297_ (.A(net1431),
    .B(net6148),
    .Y(_17494_));
 sg13g2_a21oi_1 _25298_ (.A1(net6148),
    .A2(_17493_),
    .Y(_01616_),
    .B1(_17494_));
 sg13g2_nor2_1 _25299_ (.A(\u_inv.f_next[110] ),
    .B(net7057),
    .Y(_17495_));
 sg13g2_nor2_1 _25300_ (.A(net1874),
    .B(net6148),
    .Y(_17496_));
 sg13g2_a21oi_1 _25301_ (.A1(net6149),
    .A2(_17495_),
    .Y(_01617_),
    .B1(_17496_));
 sg13g2_nor2_1 _25302_ (.A(\u_inv.f_next[111] ),
    .B(net7056),
    .Y(_17497_));
 sg13g2_nor2_1 _25303_ (.A(net3208),
    .B(net6149),
    .Y(_17498_));
 sg13g2_a21oi_1 _25304_ (.A1(net6148),
    .A2(_17497_),
    .Y(_01618_),
    .B1(_17498_));
 sg13g2_nor2_1 _25305_ (.A(\u_inv.f_next[112] ),
    .B(net7055),
    .Y(_17499_));
 sg13g2_nor2_1 _25306_ (.A(net2339),
    .B(net6146),
    .Y(_17500_));
 sg13g2_a21oi_1 _25307_ (.A1(net6132),
    .A2(_17499_),
    .Y(_01619_),
    .B1(_17500_));
 sg13g2_nor2_1 _25308_ (.A(\u_inv.f_next[113] ),
    .B(net7055),
    .Y(_17501_));
 sg13g2_nor2_1 _25309_ (.A(net2009),
    .B(net6146),
    .Y(_17502_));
 sg13g2_a21oi_1 _25310_ (.A1(net6132),
    .A2(_17501_),
    .Y(_01620_),
    .B1(_17502_));
 sg13g2_nor2_1 _25311_ (.A(\u_inv.f_next[114] ),
    .B(net7057),
    .Y(_17503_));
 sg13g2_nor2_1 _25312_ (.A(net2413),
    .B(net6146),
    .Y(_17504_));
 sg13g2_a21oi_1 _25313_ (.A1(net6146),
    .A2(_17503_),
    .Y(_01621_),
    .B1(_17504_));
 sg13g2_nor2_1 _25314_ (.A(\u_inv.f_next[115] ),
    .B(net7057),
    .Y(_17505_));
 sg13g2_nor2_1 _25315_ (.A(net3050),
    .B(net6147),
    .Y(_17506_));
 sg13g2_a21oi_1 _25316_ (.A1(net6147),
    .A2(_17505_),
    .Y(_01622_),
    .B1(_17506_));
 sg13g2_nor2_1 _25317_ (.A(net2143),
    .B(net7050),
    .Y(_17507_));
 sg13g2_nor2_1 _25318_ (.A(net2173),
    .B(net6132),
    .Y(_17508_));
 sg13g2_a21oi_1 _25319_ (.A1(net6132),
    .A2(_17507_),
    .Y(_01623_),
    .B1(_17508_));
 sg13g2_nor2_1 _25320_ (.A(\u_inv.f_next[117] ),
    .B(net7055),
    .Y(_17509_));
 sg13g2_nor2_1 _25321_ (.A(net2306),
    .B(net6146),
    .Y(_17510_));
 sg13g2_a21oi_1 _25322_ (.A1(net6146),
    .A2(_17509_),
    .Y(_01624_),
    .B1(_17510_));
 sg13g2_nor2_1 _25323_ (.A(\u_inv.f_next[118] ),
    .B(net7050),
    .Y(_17511_));
 sg13g2_nor2_1 _25324_ (.A(net1433),
    .B(net6132),
    .Y(_17512_));
 sg13g2_a21oi_1 _25325_ (.A1(net6132),
    .A2(_17511_),
    .Y(_01625_),
    .B1(_17512_));
 sg13g2_nor2_1 _25326_ (.A(\u_inv.f_next[119] ),
    .B(net7050),
    .Y(_17513_));
 sg13g2_nor2_1 _25327_ (.A(net1908),
    .B(net6128),
    .Y(_17514_));
 sg13g2_a21oi_1 _25328_ (.A1(net6128),
    .A2(_17513_),
    .Y(_01626_),
    .B1(_17514_));
 sg13g2_nor2_1 _25329_ (.A(\u_inv.f_next[120] ),
    .B(net7051),
    .Y(_17515_));
 sg13g2_nor2_1 _25330_ (.A(net1992),
    .B(net6130),
    .Y(_17516_));
 sg13g2_a21oi_1 _25331_ (.A1(net6130),
    .A2(_17515_),
    .Y(_01627_),
    .B1(_17516_));
 sg13g2_nor2_1 _25332_ (.A(\u_inv.f_next[121] ),
    .B(net7051),
    .Y(_17517_));
 sg13g2_nor2_1 _25333_ (.A(net1739),
    .B(net6130),
    .Y(_17518_));
 sg13g2_a21oi_1 _25334_ (.A1(net6130),
    .A2(_17517_),
    .Y(_01628_),
    .B1(_17518_));
 sg13g2_nor2_1 _25335_ (.A(\u_inv.f_next[122] ),
    .B(net7052),
    .Y(_17519_));
 sg13g2_nor2_1 _25336_ (.A(net2955),
    .B(net6133),
    .Y(_17520_));
 sg13g2_a21oi_1 _25337_ (.A1(net6133),
    .A2(_17519_),
    .Y(_01629_),
    .B1(_17520_));
 sg13g2_nor2_1 _25338_ (.A(\u_inv.f_next[123] ),
    .B(net7051),
    .Y(_17521_));
 sg13g2_nor2_1 _25339_ (.A(net1897),
    .B(net6131),
    .Y(_17522_));
 sg13g2_a21oi_1 _25340_ (.A1(net6131),
    .A2(_17521_),
    .Y(_01630_),
    .B1(_17522_));
 sg13g2_nor2_1 _25341_ (.A(\u_inv.f_next[124] ),
    .B(net7050),
    .Y(_17523_));
 sg13g2_nor2_1 _25342_ (.A(net3153),
    .B(net6128),
    .Y(_17524_));
 sg13g2_a21oi_1 _25343_ (.A1(net6128),
    .A2(_17523_),
    .Y(_01631_),
    .B1(_17524_));
 sg13g2_nor2_1 _25344_ (.A(\u_inv.f_next[125] ),
    .B(net7051),
    .Y(_17525_));
 sg13g2_nor2_1 _25345_ (.A(net2227),
    .B(net6128),
    .Y(_17526_));
 sg13g2_a21oi_1 _25346_ (.A1(net6129),
    .A2(_17525_),
    .Y(_01632_),
    .B1(_17526_));
 sg13g2_nor2_1 _25347_ (.A(\u_inv.f_next[126] ),
    .B(net7048),
    .Y(_17527_));
 sg13g2_nor2_1 _25348_ (.A(net3232),
    .B(net6129),
    .Y(_17528_));
 sg13g2_a21oi_1 _25349_ (.A1(net6126),
    .A2(_17527_),
    .Y(_01633_),
    .B1(_17528_));
 sg13g2_nor2_1 _25350_ (.A(\u_inv.f_next[127] ),
    .B(net7048),
    .Y(_17529_));
 sg13g2_nor2_1 _25351_ (.A(net2667),
    .B(net6129),
    .Y(_17530_));
 sg13g2_a21oi_1 _25352_ (.A1(net6126),
    .A2(_17529_),
    .Y(_01634_),
    .B1(_17530_));
 sg13g2_nor2_1 _25353_ (.A(\u_inv.f_next[128] ),
    .B(net7046),
    .Y(_17531_));
 sg13g2_nor2_1 _25354_ (.A(net2766),
    .B(net6124),
    .Y(_17532_));
 sg13g2_a21oi_1 _25355_ (.A1(net6125),
    .A2(_17531_),
    .Y(_01635_),
    .B1(_17532_));
 sg13g2_nor2_1 _25356_ (.A(\u_inv.f_next[129] ),
    .B(net7046),
    .Y(_17533_));
 sg13g2_nor2_1 _25357_ (.A(net2503),
    .B(net6123),
    .Y(_17534_));
 sg13g2_a21oi_1 _25358_ (.A1(net6123),
    .A2(_17533_),
    .Y(_01636_),
    .B1(_17534_));
 sg13g2_nor2_1 _25359_ (.A(\u_inv.f_next[130] ),
    .B(net7046),
    .Y(_17535_));
 sg13g2_nor2_1 _25360_ (.A(net1623),
    .B(net6120),
    .Y(_17536_));
 sg13g2_a21oi_1 _25361_ (.A1(net6119),
    .A2(_17535_),
    .Y(_01637_),
    .B1(_17536_));
 sg13g2_nor2_1 _25362_ (.A(\u_inv.f_next[131] ),
    .B(net7047),
    .Y(_17537_));
 sg13g2_nor2_1 _25363_ (.A(net2149),
    .B(net6120),
    .Y(_17538_));
 sg13g2_a21oi_1 _25364_ (.A1(net6120),
    .A2(_17537_),
    .Y(_01638_),
    .B1(_17538_));
 sg13g2_nor2_1 _25365_ (.A(\u_inv.f_next[132] ),
    .B(net7045),
    .Y(_17539_));
 sg13g2_nor2_1 _25366_ (.A(net2043),
    .B(net6119),
    .Y(_17540_));
 sg13g2_a21oi_1 _25367_ (.A1(net6119),
    .A2(_17539_),
    .Y(_01639_),
    .B1(_17540_));
 sg13g2_nor2_1 _25368_ (.A(\u_inv.f_next[133] ),
    .B(net7045),
    .Y(_17541_));
 sg13g2_nor2_1 _25369_ (.A(net3084),
    .B(net6119),
    .Y(_17542_));
 sg13g2_a21oi_1 _25370_ (.A1(net6120),
    .A2(_17541_),
    .Y(_01640_),
    .B1(_17542_));
 sg13g2_nor2_1 _25371_ (.A(\u_inv.f_next[134] ),
    .B(net7040),
    .Y(_17543_));
 sg13g2_nor2_1 _25372_ (.A(net2714),
    .B(net6105),
    .Y(_17544_));
 sg13g2_a21oi_1 _25373_ (.A1(net6105),
    .A2(_17543_),
    .Y(_01641_),
    .B1(_17544_));
 sg13g2_nor2_1 _25374_ (.A(\u_inv.f_next[135] ),
    .B(net7043),
    .Y(_17545_));
 sg13g2_nor2_1 _25375_ (.A(net3103),
    .B(net6105),
    .Y(_17546_));
 sg13g2_a21oi_1 _25376_ (.A1(net6105),
    .A2(_17545_),
    .Y(_01642_),
    .B1(_17546_));
 sg13g2_nor2_1 _25377_ (.A(\u_inv.f_next[136] ),
    .B(net7042),
    .Y(_17547_));
 sg13g2_nor2_1 _25378_ (.A(net2102),
    .B(net6107),
    .Y(_17548_));
 sg13g2_a21oi_1 _25379_ (.A1(net6107),
    .A2(_17547_),
    .Y(_01643_),
    .B1(_17548_));
 sg13g2_nor2_1 _25380_ (.A(\u_inv.f_next[137] ),
    .B(net7042),
    .Y(_17549_));
 sg13g2_nor2_1 _25381_ (.A(net1972),
    .B(net6107),
    .Y(_17550_));
 sg13g2_a21oi_1 _25382_ (.A1(net6107),
    .A2(_17549_),
    .Y(_01644_),
    .B1(_17550_));
 sg13g2_nor2_1 _25383_ (.A(\u_inv.f_next[138] ),
    .B(net7042),
    .Y(_17551_));
 sg13g2_nor2_1 _25384_ (.A(net1621),
    .B(net6107),
    .Y(_17552_));
 sg13g2_a21oi_1 _25385_ (.A1(net6110),
    .A2(_17551_),
    .Y(_01645_),
    .B1(_17552_));
 sg13g2_nor2_1 _25386_ (.A(\u_inv.f_next[139] ),
    .B(net7043),
    .Y(_17553_));
 sg13g2_nor2_1 _25387_ (.A(net3159),
    .B(net6110),
    .Y(_17554_));
 sg13g2_a21oi_1 _25388_ (.A1(net6110),
    .A2(_17553_),
    .Y(_01646_),
    .B1(_17554_));
 sg13g2_nor2_1 _25389_ (.A(\u_inv.f_next[140] ),
    .B(net7038),
    .Y(_17555_));
 sg13g2_nor2_1 _25390_ (.A(net2374),
    .B(net6101),
    .Y(_17556_));
 sg13g2_a21oi_1 _25391_ (.A1(net6101),
    .A2(_17555_),
    .Y(_01647_),
    .B1(_17556_));
 sg13g2_nor2_1 _25392_ (.A(\u_inv.f_next[141] ),
    .B(net7038),
    .Y(_17557_));
 sg13g2_nor2_1 _25393_ (.A(net2488),
    .B(net6101),
    .Y(_17558_));
 sg13g2_a21oi_1 _25394_ (.A1(net6101),
    .A2(_17557_),
    .Y(_01648_),
    .B1(_17558_));
 sg13g2_nor2_1 _25395_ (.A(\u_inv.f_next[142] ),
    .B(net7038),
    .Y(_17559_));
 sg13g2_nor2_1 _25396_ (.A(net2274),
    .B(net6101),
    .Y(_17560_));
 sg13g2_a21oi_1 _25397_ (.A1(net6101),
    .A2(_17559_),
    .Y(_01649_),
    .B1(_17560_));
 sg13g2_nor2_1 _25398_ (.A(\u_inv.f_next[143] ),
    .B(net7042),
    .Y(_17561_));
 sg13g2_nor2_1 _25399_ (.A(net3013),
    .B(net6107),
    .Y(_17562_));
 sg13g2_a21oi_1 _25400_ (.A1(net6103),
    .A2(_17561_),
    .Y(_01650_),
    .B1(_17562_));
 sg13g2_nor2_1 _25401_ (.A(\u_inv.f_next[144] ),
    .B(net7040),
    .Y(_17563_));
 sg13g2_nor2_1 _25402_ (.A(net1860),
    .B(net6105),
    .Y(_17564_));
 sg13g2_a21oi_1 _25403_ (.A1(net6105),
    .A2(_17563_),
    .Y(_01651_),
    .B1(_17564_));
 sg13g2_nor2_1 _25404_ (.A(net1473),
    .B(net7041),
    .Y(_17565_));
 sg13g2_nor2_1 _25405_ (.A(net1504),
    .B(net6105),
    .Y(_17566_));
 sg13g2_a21oi_1 _25406_ (.A1(net6105),
    .A2(_17565_),
    .Y(_01652_),
    .B1(_17566_));
 sg13g2_nor2_1 _25407_ (.A(\u_inv.f_next[146] ),
    .B(net7041),
    .Y(_17567_));
 sg13g2_nor2_1 _25408_ (.A(net1667),
    .B(net6104),
    .Y(_17568_));
 sg13g2_a21oi_1 _25409_ (.A1(net6104),
    .A2(_17567_),
    .Y(_01653_),
    .B1(_17568_));
 sg13g2_nor2_1 _25410_ (.A(\u_inv.f_next[147] ),
    .B(net7041),
    .Y(_17569_));
 sg13g2_nor2_1 _25411_ (.A(net3113),
    .B(net6104),
    .Y(_17570_));
 sg13g2_a21oi_1 _25412_ (.A1(net6104),
    .A2(_17569_),
    .Y(_01654_),
    .B1(_17570_));
 sg13g2_nor2_1 _25413_ (.A(\u_inv.f_next[148] ),
    .B(net7039),
    .Y(_17571_));
 sg13g2_nor2_1 _25414_ (.A(net2768),
    .B(net6103),
    .Y(_17572_));
 sg13g2_a21oi_1 _25415_ (.A1(net6103),
    .A2(_17571_),
    .Y(_01655_),
    .B1(_17572_));
 sg13g2_nor2_1 _25416_ (.A(\u_inv.f_next[149] ),
    .B(net7039),
    .Y(_17573_));
 sg13g2_nor2_1 _25417_ (.A(net2904),
    .B(net6103),
    .Y(_17574_));
 sg13g2_a21oi_1 _25418_ (.A1(net6103),
    .A2(_17573_),
    .Y(_01656_),
    .B1(_17574_));
 sg13g2_nor2_1 _25419_ (.A(\u_inv.f_next[150] ),
    .B(net7040),
    .Y(_17575_));
 sg13g2_nor2_1 _25420_ (.A(net1820),
    .B(net6103),
    .Y(_17576_));
 sg13g2_a21oi_1 _25421_ (.A1(net6106),
    .A2(_17575_),
    .Y(_01657_),
    .B1(_17576_));
 sg13g2_nor2_1 _25422_ (.A(net3230),
    .B(net7040),
    .Y(_17577_));
 sg13g2_nor2_1 _25423_ (.A(net3270),
    .B(net6106),
    .Y(_17578_));
 sg13g2_a21oi_1 _25424_ (.A1(net6106),
    .A2(_17577_),
    .Y(_01658_),
    .B1(_17578_));
 sg13g2_nor2_1 _25425_ (.A(\u_inv.f_next[152] ),
    .B(net7037),
    .Y(_17579_));
 sg13g2_nor2_1 _25426_ (.A(net2748),
    .B(net6099),
    .Y(_17580_));
 sg13g2_a21oi_1 _25427_ (.A1(net6099),
    .A2(_17579_),
    .Y(_01659_),
    .B1(_17580_));
 sg13g2_nor2_1 _25428_ (.A(\u_inv.f_next[153] ),
    .B(net7037),
    .Y(_17581_));
 sg13g2_nor2_1 _25429_ (.A(net2881),
    .B(net6099),
    .Y(_17582_));
 sg13g2_a21oi_1 _25430_ (.A1(net6099),
    .A2(_17581_),
    .Y(_01660_),
    .B1(_17582_));
 sg13g2_nor2_1 _25431_ (.A(\u_inv.f_next[154] ),
    .B(net7038),
    .Y(_17583_));
 sg13g2_nor2_1 _25432_ (.A(net1787),
    .B(net6099),
    .Y(_17584_));
 sg13g2_a21oi_1 _25433_ (.A1(net6099),
    .A2(_17583_),
    .Y(_01661_),
    .B1(_17584_));
 sg13g2_nor2_1 _25434_ (.A(\u_inv.f_next[155] ),
    .B(net7038),
    .Y(_17585_));
 sg13g2_nor2_1 _25435_ (.A(net2177),
    .B(net6102),
    .Y(_17586_));
 sg13g2_a21oi_1 _25436_ (.A1(net6102),
    .A2(_17585_),
    .Y(_01662_),
    .B1(_17586_));
 sg13g2_nor2_1 _25437_ (.A(\u_inv.f_next[156] ),
    .B(net7036),
    .Y(_17587_));
 sg13g2_nor2_1 _25438_ (.A(net1634),
    .B(net6097),
    .Y(_17588_));
 sg13g2_a21oi_1 _25439_ (.A1(net6097),
    .A2(_17587_),
    .Y(_01663_),
    .B1(_17588_));
 sg13g2_nor2_1 _25440_ (.A(\u_inv.f_next[157] ),
    .B(net7036),
    .Y(_17589_));
 sg13g2_nor2_1 _25441_ (.A(net2996),
    .B(net6097),
    .Y(_17590_));
 sg13g2_a21oi_1 _25442_ (.A1(net6097),
    .A2(_17589_),
    .Y(_01664_),
    .B1(_17590_));
 sg13g2_nor2_1 _25443_ (.A(\u_inv.f_next[158] ),
    .B(net7037),
    .Y(_17591_));
 sg13g2_nor2_1 _25444_ (.A(net2540),
    .B(net6098),
    .Y(_17592_));
 sg13g2_a21oi_1 _25445_ (.A1(net6098),
    .A2(_17591_),
    .Y(_01665_),
    .B1(_17592_));
 sg13g2_nor2_1 _25446_ (.A(\u_inv.f_next[159] ),
    .B(net7037),
    .Y(_17593_));
 sg13g2_nor2_1 _25447_ (.A(net2355),
    .B(net6098),
    .Y(_17594_));
 sg13g2_a21oi_1 _25448_ (.A1(net6098),
    .A2(_17593_),
    .Y(_01666_),
    .B1(_17594_));
 sg13g2_nor2_1 _25449_ (.A(\u_inv.f_next[160] ),
    .B(net7031),
    .Y(_17595_));
 sg13g2_nor2_1 _25450_ (.A(net2640),
    .B(net6078),
    .Y(_17596_));
 sg13g2_a21oi_1 _25451_ (.A1(net6078),
    .A2(_17595_),
    .Y(_01667_),
    .B1(_17596_));
 sg13g2_nor2_1 _25452_ (.A(\u_inv.f_next[161] ),
    .B(net7032),
    .Y(_17597_));
 sg13g2_nor2_1 _25453_ (.A(net2906),
    .B(net6078),
    .Y(_17598_));
 sg13g2_a21oi_1 _25454_ (.A1(net6078),
    .A2(_17597_),
    .Y(_01668_),
    .B1(_17598_));
 sg13g2_nor2_1 _25455_ (.A(\u_inv.f_next[162] ),
    .B(net7032),
    .Y(_17599_));
 sg13g2_nor2_1 _25456_ (.A(net1844),
    .B(net6078),
    .Y(_17600_));
 sg13g2_a21oi_1 _25457_ (.A1(net6078),
    .A2(_17599_),
    .Y(_01669_),
    .B1(_17600_));
 sg13g2_nor2_1 _25458_ (.A(\u_inv.f_next[163] ),
    .B(net7031),
    .Y(_17601_));
 sg13g2_nor2_1 _25459_ (.A(net1252),
    .B(net6077),
    .Y(_17602_));
 sg13g2_a21oi_1 _25460_ (.A1(net6077),
    .A2(_17601_),
    .Y(_01670_),
    .B1(_17602_));
 sg13g2_nor2_1 _25461_ (.A(\u_inv.f_next[164] ),
    .B(net7030),
    .Y(_17603_));
 sg13g2_nor2_1 _25462_ (.A(net2602),
    .B(net6061),
    .Y(_17604_));
 sg13g2_a21oi_1 _25463_ (.A1(net6061),
    .A2(_17603_),
    .Y(_01671_),
    .B1(_17604_));
 sg13g2_nor2_1 _25464_ (.A(net1511),
    .B(net7030),
    .Y(_17605_));
 sg13g2_nor2_1 _25465_ (.A(net2045),
    .B(net6061),
    .Y(_17606_));
 sg13g2_a21oi_1 _25466_ (.A1(net6061),
    .A2(_17605_),
    .Y(_01672_),
    .B1(_17606_));
 sg13g2_nor2_1 _25467_ (.A(\u_inv.f_next[166] ),
    .B(net7029),
    .Y(_17607_));
 sg13g2_nor2_1 _25468_ (.A(net2377),
    .B(net6060),
    .Y(_17608_));
 sg13g2_a21oi_1 _25469_ (.A1(net6060),
    .A2(_17607_),
    .Y(_01673_),
    .B1(_17608_));
 sg13g2_nor2_1 _25470_ (.A(\u_inv.f_next[167] ),
    .B(net7029),
    .Y(_17609_));
 sg13g2_nor2_1 _25471_ (.A(net2185),
    .B(net6060),
    .Y(_17610_));
 sg13g2_a21oi_1 _25472_ (.A1(net6060),
    .A2(_17609_),
    .Y(_01674_),
    .B1(_17610_));
 sg13g2_nor2_1 _25473_ (.A(\u_inv.f_next[168] ),
    .B(net7029),
    .Y(_17611_));
 sg13g2_nor2_1 _25474_ (.A(net2864),
    .B(net6060),
    .Y(_17612_));
 sg13g2_a21oi_1 _25475_ (.A1(net6060),
    .A2(_17611_),
    .Y(_01675_),
    .B1(_17612_));
 sg13g2_nor2_1 _25476_ (.A(\u_inv.f_next[169] ),
    .B(net7029),
    .Y(_17613_));
 sg13g2_nor2_1 _25477_ (.A(net2432),
    .B(net6060),
    .Y(_17614_));
 sg13g2_a21oi_1 _25478_ (.A1(net6060),
    .A2(_17613_),
    .Y(_01676_),
    .B1(_17614_));
 sg13g2_nor2_1 _25479_ (.A(\u_inv.f_next[170] ),
    .B(net7026),
    .Y(_17615_));
 sg13g2_nor2_1 _25480_ (.A(net2017),
    .B(net6058),
    .Y(_17616_));
 sg13g2_a21oi_1 _25481_ (.A1(net6057),
    .A2(_17615_),
    .Y(_01677_),
    .B1(_17616_));
 sg13g2_nor2_1 _25482_ (.A(net2927),
    .B(net7026),
    .Y(_17617_));
 sg13g2_nor2_1 _25483_ (.A(net3241),
    .B(net6059),
    .Y(_17618_));
 sg13g2_a21oi_1 _25484_ (.A1(net6058),
    .A2(_17617_),
    .Y(_01678_),
    .B1(_17618_));
 sg13g2_nor2_1 _25485_ (.A(\u_inv.f_next[172] ),
    .B(net7026),
    .Y(_17619_));
 sg13g2_nor2_1 _25486_ (.A(net2616),
    .B(net6057),
    .Y(_17620_));
 sg13g2_a21oi_1 _25487_ (.A1(net6057),
    .A2(_17619_),
    .Y(_01679_),
    .B1(_17620_));
 sg13g2_nor2_1 _25488_ (.A(\u_inv.f_next[173] ),
    .B(net7028),
    .Y(_17621_));
 sg13g2_nor2_1 _25489_ (.A(net1789),
    .B(net6057),
    .Y(_17622_));
 sg13g2_a21oi_1 _25490_ (.A1(net6057),
    .A2(_17621_),
    .Y(_01680_),
    .B1(_17622_));
 sg13g2_nor2_1 _25491_ (.A(\u_inv.f_next[174] ),
    .B(net7026),
    .Y(_17623_));
 sg13g2_nor2_1 _25492_ (.A(net1777),
    .B(net6057),
    .Y(_17624_));
 sg13g2_a21oi_1 _25493_ (.A1(net6056),
    .A2(_17623_),
    .Y(_01681_),
    .B1(_17624_));
 sg13g2_nor2_1 _25494_ (.A(net2493),
    .B(net7026),
    .Y(_17625_));
 sg13g2_nor2_1 _25495_ (.A(net2952),
    .B(net6057),
    .Y(_17626_));
 sg13g2_a21oi_1 _25496_ (.A1(net6057),
    .A2(_17625_),
    .Y(_01682_),
    .B1(_17626_));
 sg13g2_nor2_1 _25497_ (.A(\u_inv.f_next[176] ),
    .B(net7024),
    .Y(_17627_));
 sg13g2_nor2_1 _25498_ (.A(net3032),
    .B(net6055),
    .Y(_17628_));
 sg13g2_a21oi_1 _25499_ (.A1(net6055),
    .A2(_17627_),
    .Y(_01683_),
    .B1(_17628_));
 sg13g2_nor2_1 _25500_ (.A(net2064),
    .B(net7024),
    .Y(_17629_));
 sg13g2_nor2_1 _25501_ (.A(net2468),
    .B(net6055),
    .Y(_17630_));
 sg13g2_a21oi_1 _25502_ (.A1(net6055),
    .A2(_17629_),
    .Y(_01684_),
    .B1(_17630_));
 sg13g2_nor2_1 _25503_ (.A(\u_inv.f_next[178] ),
    .B(net7027),
    .Y(_17631_));
 sg13g2_nor2_1 _25504_ (.A(net2789),
    .B(net6056),
    .Y(_17632_));
 sg13g2_a21oi_1 _25505_ (.A1(net6056),
    .A2(_17631_),
    .Y(_01685_),
    .B1(_17632_));
 sg13g2_nor2_1 _25506_ (.A(net2830),
    .B(net7027),
    .Y(_17633_));
 sg13g2_nor2_1 _25507_ (.A(net3190),
    .B(net6056),
    .Y(_17634_));
 sg13g2_a21oi_1 _25508_ (.A1(net6056),
    .A2(_17633_),
    .Y(_01686_),
    .B1(_17634_));
 sg13g2_nor2_1 _25509_ (.A(net2716),
    .B(net7020),
    .Y(_17635_));
 sg13g2_nor2_1 _25510_ (.A(net2831),
    .B(net6041),
    .Y(_17636_));
 sg13g2_a21oi_1 _25511_ (.A1(net6040),
    .A2(_17635_),
    .Y(_01687_),
    .B1(_17636_));
 sg13g2_nor2_1 _25512_ (.A(\u_inv.f_next[181] ),
    .B(net7020),
    .Y(_17637_));
 sg13g2_nor2_1 _25513_ (.A(net2104),
    .B(net6041),
    .Y(_17638_));
 sg13g2_a21oi_1 _25514_ (.A1(net6040),
    .A2(_17637_),
    .Y(_01688_),
    .B1(_17638_));
 sg13g2_nor2_1 _25515_ (.A(\u_inv.f_next[182] ),
    .B(net7022),
    .Y(_17639_));
 sg13g2_nor2_1 _25516_ (.A(net2795),
    .B(net6040),
    .Y(_17640_));
 sg13g2_a21oi_1 _25517_ (.A1(net6041),
    .A2(_17639_),
    .Y(_01689_),
    .B1(_17640_));
 sg13g2_nor2_1 _25518_ (.A(\u_inv.f_next[183] ),
    .B(net7020),
    .Y(_17641_));
 sg13g2_nor2_1 _25519_ (.A(net1185),
    .B(net6041),
    .Y(_17642_));
 sg13g2_a21oi_1 _25520_ (.A1(net6040),
    .A2(_17641_),
    .Y(_01690_),
    .B1(_17642_));
 sg13g2_nor2_1 _25521_ (.A(\u_inv.f_next[184] ),
    .B(net7021),
    .Y(_17643_));
 sg13g2_nor2_1 _25522_ (.A(net1650),
    .B(net6042),
    .Y(_17644_));
 sg13g2_a21oi_1 _25523_ (.A1(net6039),
    .A2(_17643_),
    .Y(_01691_),
    .B1(_17644_));
 sg13g2_nor2_1 _25524_ (.A(\u_inv.f_next[185] ),
    .B(net7021),
    .Y(_17645_));
 sg13g2_nor2_1 _25525_ (.A(net3136),
    .B(net6039),
    .Y(_17646_));
 sg13g2_a21oi_1 _25526_ (.A1(net6038),
    .A2(_17645_),
    .Y(_01692_),
    .B1(_17646_));
 sg13g2_nor2_1 _25527_ (.A(\u_inv.f_next[186] ),
    .B(net7021),
    .Y(_17647_));
 sg13g2_nor2_1 _25528_ (.A(net2559),
    .B(net6038),
    .Y(_17648_));
 sg13g2_a21oi_1 _25529_ (.A1(net6038),
    .A2(_17647_),
    .Y(_01693_),
    .B1(_17648_));
 sg13g2_nor2_1 _25530_ (.A(\u_inv.f_next[187] ),
    .B(net7018),
    .Y(_17649_));
 sg13g2_nor2_1 _25531_ (.A(net2593),
    .B(net6038),
    .Y(_17650_));
 sg13g2_a21oi_1 _25532_ (.A1(net6033),
    .A2(_17649_),
    .Y(_01694_),
    .B1(_17650_));
 sg13g2_nor2_1 _25533_ (.A(\u_inv.f_next[188] ),
    .B(net7018),
    .Y(_17651_));
 sg13g2_nor2_1 _25534_ (.A(net1957),
    .B(net6034),
    .Y(_17652_));
 sg13g2_a21oi_1 _25535_ (.A1(net6034),
    .A2(_17651_),
    .Y(_01695_),
    .B1(_17652_));
 sg13g2_nor2_1 _25536_ (.A(\u_inv.f_next[189] ),
    .B(net7018),
    .Y(_17653_));
 sg13g2_nor2_1 _25537_ (.A(net1996),
    .B(net6034),
    .Y(_17654_));
 sg13g2_a21oi_1 _25538_ (.A1(net6034),
    .A2(_17653_),
    .Y(_01696_),
    .B1(_17654_));
 sg13g2_nor2_1 _25539_ (.A(\u_inv.f_next[190] ),
    .B(net7018),
    .Y(_17655_));
 sg13g2_nor2_1 _25540_ (.A(net2204),
    .B(net6034),
    .Y(_17656_));
 sg13g2_a21oi_1 _25541_ (.A1(net6034),
    .A2(_17655_),
    .Y(_01697_),
    .B1(_17656_));
 sg13g2_nor2_1 _25542_ (.A(\u_inv.f_next[191] ),
    .B(net7017),
    .Y(_17657_));
 sg13g2_nor2_1 _25543_ (.A(net2676),
    .B(net6033),
    .Y(_17658_));
 sg13g2_a21oi_1 _25544_ (.A1(net6033),
    .A2(_17657_),
    .Y(_01698_),
    .B1(_17658_));
 sg13g2_nor2_1 _25545_ (.A(\u_inv.f_next[192] ),
    .B(net7019),
    .Y(_17659_));
 sg13g2_nor2_1 _25546_ (.A(net3090),
    .B(net6035),
    .Y(_17660_));
 sg13g2_a21oi_1 _25547_ (.A1(net6035),
    .A2(_17659_),
    .Y(_01699_),
    .B1(_17660_));
 sg13g2_nor2_1 _25548_ (.A(\u_inv.f_next[193] ),
    .B(net7019),
    .Y(_17661_));
 sg13g2_nor2_1 _25549_ (.A(net2419),
    .B(net6035),
    .Y(_17662_));
 sg13g2_a21oi_1 _25550_ (.A1(net6035),
    .A2(_17661_),
    .Y(_01700_),
    .B1(_17662_));
 sg13g2_nor2_1 _25551_ (.A(\u_inv.f_next[194] ),
    .B(net7019),
    .Y(_17663_));
 sg13g2_nor2_1 _25552_ (.A(net2385),
    .B(net6035),
    .Y(_17664_));
 sg13g2_a21oi_1 _25553_ (.A1(net6035),
    .A2(_17663_),
    .Y(_01701_),
    .B1(_17664_));
 sg13g2_nor2_1 _25554_ (.A(\u_inv.f_next[195] ),
    .B(net7004),
    .Y(_17665_));
 sg13g2_nor2_1 _25555_ (.A(net2567),
    .B(net6021),
    .Y(_17666_));
 sg13g2_a21oi_1 _25556_ (.A1(net6021),
    .A2(_17665_),
    .Y(_01702_),
    .B1(_17666_));
 sg13g2_nor2_1 _25557_ (.A(\u_inv.f_next[196] ),
    .B(net7004),
    .Y(_17667_));
 sg13g2_nor2_1 _25558_ (.A(net3155),
    .B(net6022),
    .Y(_17668_));
 sg13g2_a21oi_1 _25559_ (.A1(net6022),
    .A2(_17667_),
    .Y(_01703_),
    .B1(_17668_));
 sg13g2_nor2_1 _25560_ (.A(\u_inv.f_next[197] ),
    .B(net7004),
    .Y(_17669_));
 sg13g2_nor2_1 _25561_ (.A(net2866),
    .B(net6021),
    .Y(_17670_));
 sg13g2_a21oi_1 _25562_ (.A1(net6021),
    .A2(_17669_),
    .Y(_01704_),
    .B1(_17670_));
 sg13g2_nor2_1 _25563_ (.A(\u_inv.f_next[198] ),
    .B(net7004),
    .Y(_17671_));
 sg13g2_nor2_1 _25564_ (.A(net1953),
    .B(net6021),
    .Y(_17672_));
 sg13g2_a21oi_1 _25565_ (.A1(net6021),
    .A2(_17671_),
    .Y(_01705_),
    .B1(_17672_));
 sg13g2_nor2_1 _25566_ (.A(net2380),
    .B(net7004),
    .Y(_17673_));
 sg13g2_nor2_1 _25567_ (.A(net2384),
    .B(net6021),
    .Y(_17674_));
 sg13g2_a21oi_1 _25568_ (.A1(net6021),
    .A2(_17673_),
    .Y(_01706_),
    .B1(_17674_));
 sg13g2_nor2_1 _25569_ (.A(\u_inv.f_next[200] ),
    .B(net7005),
    .Y(_17675_));
 sg13g2_nor2_1 _25570_ (.A(net2958),
    .B(net6022),
    .Y(_17676_));
 sg13g2_a21oi_1 _25571_ (.A1(net6022),
    .A2(_17675_),
    .Y(_01707_),
    .B1(_17676_));
 sg13g2_nor2_1 _25572_ (.A(\u_inv.f_next[201] ),
    .B(net7003),
    .Y(_17677_));
 sg13g2_nor2_1 _25573_ (.A(net2408),
    .B(net6020),
    .Y(_17678_));
 sg13g2_a21oi_1 _25574_ (.A1(net6020),
    .A2(_17677_),
    .Y(_01708_),
    .B1(_17678_));
 sg13g2_nor2_1 _25575_ (.A(\u_inv.f_next[202] ),
    .B(net7003),
    .Y(_17679_));
 sg13g2_nor2_1 _25576_ (.A(net1810),
    .B(net6020),
    .Y(_17680_));
 sg13g2_a21oi_1 _25577_ (.A1(net6020),
    .A2(_17679_),
    .Y(_01709_),
    .B1(_17680_));
 sg13g2_nor2_1 _25578_ (.A(\u_inv.f_next[203] ),
    .B(net7003),
    .Y(_17681_));
 sg13g2_nor2_1 _25579_ (.A(net2984),
    .B(net6020),
    .Y(_17682_));
 sg13g2_a21oi_1 _25580_ (.A1(net6020),
    .A2(_17681_),
    .Y(_01710_),
    .B1(_17682_));
 sg13g2_nor2_1 _25581_ (.A(\u_inv.f_next[204] ),
    .B(net6996),
    .Y(_17683_));
 sg13g2_nor2_1 _25582_ (.A(net2349),
    .B(net6020),
    .Y(_17684_));
 sg13g2_a21oi_1 _25583_ (.A1(net6020),
    .A2(_17683_),
    .Y(_01711_),
    .B1(_17684_));
 sg13g2_nor2_1 _25584_ (.A(\u_inv.f_next[205] ),
    .B(net6996),
    .Y(_17685_));
 sg13g2_nor2_1 _25585_ (.A(net1773),
    .B(net6011),
    .Y(_17686_));
 sg13g2_a21oi_1 _25586_ (.A1(net6011),
    .A2(_17685_),
    .Y(_01712_),
    .B1(_17686_));
 sg13g2_nor2_1 _25587_ (.A(\u_inv.f_next[206] ),
    .B(net6996),
    .Y(_17687_));
 sg13g2_nor2_1 _25588_ (.A(net2531),
    .B(net6011),
    .Y(_17688_));
 sg13g2_a21oi_1 _25589_ (.A1(net6011),
    .A2(_17687_),
    .Y(_01713_),
    .B1(_17688_));
 sg13g2_nor2_1 _25590_ (.A(\u_inv.f_next[207] ),
    .B(net6996),
    .Y(_17689_));
 sg13g2_nor2_1 _25591_ (.A(net2163),
    .B(net6011),
    .Y(_17690_));
 sg13g2_a21oi_1 _25592_ (.A1(net6011),
    .A2(_17689_),
    .Y(_01714_),
    .B1(_17690_));
 sg13g2_nor2_1 _25593_ (.A(\u_inv.f_next[208] ),
    .B(net6997),
    .Y(_17691_));
 sg13g2_nor2_1 _25594_ (.A(net3244),
    .B(net6011),
    .Y(_17692_));
 sg13g2_a21oi_1 _25595_ (.A1(net6011),
    .A2(_17691_),
    .Y(_01715_),
    .B1(_17692_));
 sg13g2_nor2_1 _25596_ (.A(\u_inv.f_next[209] ),
    .B(net6997),
    .Y(_17693_));
 sg13g2_nor2_1 _25597_ (.A(net2308),
    .B(net6009),
    .Y(_17694_));
 sg13g2_a21oi_1 _25598_ (.A1(net6009),
    .A2(_17693_),
    .Y(_01716_),
    .B1(_17694_));
 sg13g2_nor2_1 _25599_ (.A(\u_inv.f_next[210] ),
    .B(net6997),
    .Y(_17695_));
 sg13g2_nor2_1 _25600_ (.A(net3131),
    .B(net6009),
    .Y(_17696_));
 sg13g2_a21oi_1 _25601_ (.A1(net6009),
    .A2(_17695_),
    .Y(_01717_),
    .B1(_17696_));
 sg13g2_nor2_1 _25602_ (.A(\u_inv.f_next[211] ),
    .B(net6997),
    .Y(_17697_));
 sg13g2_nor2_1 _25603_ (.A(net2462),
    .B(net6009),
    .Y(_17698_));
 sg13g2_a21oi_1 _25604_ (.A1(net6009),
    .A2(_17697_),
    .Y(_01718_),
    .B1(_17698_));
 sg13g2_nor2_1 _25605_ (.A(\u_inv.f_next[212] ),
    .B(net6997),
    .Y(_17699_));
 sg13g2_nor2_1 _25606_ (.A(net2943),
    .B(net6009),
    .Y(_17700_));
 sg13g2_a21oi_1 _25607_ (.A1(net6009),
    .A2(_17699_),
    .Y(_01719_),
    .B1(_17700_));
 sg13g2_nor2_1 _25608_ (.A(\u_inv.f_next[213] ),
    .B(net6997),
    .Y(_17701_));
 sg13g2_nor2_1 _25609_ (.A(net2753),
    .B(net6010),
    .Y(_17702_));
 sg13g2_a21oi_1 _25610_ (.A1(net6010),
    .A2(_17701_),
    .Y(_01720_),
    .B1(_17702_));
 sg13g2_nor2_1 _25611_ (.A(\u_inv.f_next[214] ),
    .B(net6997),
    .Y(_17703_));
 sg13g2_nor2_1 _25612_ (.A(net2516),
    .B(net6010),
    .Y(_17704_));
 sg13g2_a21oi_1 _25613_ (.A1(net6010),
    .A2(_17703_),
    .Y(_01721_),
    .B1(_17704_));
 sg13g2_nor2_1 _25614_ (.A(\u_inv.f_next[215] ),
    .B(net6998),
    .Y(_17705_));
 sg13g2_nor2_1 _25615_ (.A(net2445),
    .B(net6010),
    .Y(_17706_));
 sg13g2_a21oi_1 _25616_ (.A1(net6010),
    .A2(_17705_),
    .Y(_01722_),
    .B1(_17706_));
 sg13g2_nor2_1 _25617_ (.A(net2052),
    .B(net7000),
    .Y(_17707_));
 sg13g2_nor2_1 _25618_ (.A(net2387),
    .B(net6012),
    .Y(_17708_));
 sg13g2_a21oi_1 _25619_ (.A1(net6012),
    .A2(_17707_),
    .Y(_01723_),
    .B1(_17708_));
 sg13g2_nor2_1 _25620_ (.A(net2634),
    .B(net7007),
    .Y(_17709_));
 sg13g2_nor2_1 _25621_ (.A(net2960),
    .B(net6012),
    .Y(_17710_));
 sg13g2_a21oi_1 _25622_ (.A1(net6012),
    .A2(_17709_),
    .Y(_01724_),
    .B1(_17710_));
 sg13g2_nor2_1 _25623_ (.A(\u_inv.f_next[218] ),
    .B(net7000),
    .Y(_17711_));
 sg13g2_nor2_1 _25624_ (.A(net2699),
    .B(net6019),
    .Y(_17712_));
 sg13g2_a21oi_1 _25625_ (.A1(net6019),
    .A2(_17711_),
    .Y(_01725_),
    .B1(_17712_));
 sg13g2_nor2_1 _25626_ (.A(net1726),
    .B(net7000),
    .Y(_17713_));
 sg13g2_nor2_1 _25627_ (.A(net2160),
    .B(net6019),
    .Y(_17714_));
 sg13g2_a21oi_1 _25628_ (.A1(net6019),
    .A2(_17713_),
    .Y(_01726_),
    .B1(_17714_));
 sg13g2_nor2_1 _25629_ (.A(\u_inv.f_next[220] ),
    .B(net6998),
    .Y(_17715_));
 sg13g2_nor2_1 _25630_ (.A(net2966),
    .B(net6015),
    .Y(_17716_));
 sg13g2_a21oi_1 _25631_ (.A1(net6015),
    .A2(_17715_),
    .Y(_01727_),
    .B1(_17716_));
 sg13g2_nor2_1 _25632_ (.A(\u_inv.f_next[221] ),
    .B(net6998),
    .Y(_17717_));
 sg13g2_nor2_1 _25633_ (.A(net3034),
    .B(net6015),
    .Y(_17718_));
 sg13g2_a21oi_1 _25634_ (.A1(net6015),
    .A2(_17717_),
    .Y(_01728_),
    .B1(_17718_));
 sg13g2_nor2_1 _25635_ (.A(\u_inv.f_next[222] ),
    .B(net6998),
    .Y(_17719_));
 sg13g2_nor2_1 _25636_ (.A(net2695),
    .B(net6014),
    .Y(_17720_));
 sg13g2_a21oi_1 _25637_ (.A1(net6014),
    .A2(_17719_),
    .Y(_01729_),
    .B1(_17720_));
 sg13g2_nor2_1 _25638_ (.A(\u_inv.f_next[223] ),
    .B(net6998),
    .Y(_17721_));
 sg13g2_nor2_1 _25639_ (.A(net2206),
    .B(net6014),
    .Y(_17722_));
 sg13g2_a21oi_1 _25640_ (.A1(net6014),
    .A2(_17721_),
    .Y(_01730_),
    .B1(_17722_));
 sg13g2_nor2_1 _25641_ (.A(\u_inv.f_next[224] ),
    .B(net6998),
    .Y(_17723_));
 sg13g2_nor2_1 _25642_ (.A(net1577),
    .B(net6014),
    .Y(_17724_));
 sg13g2_a21oi_1 _25643_ (.A1(net6014),
    .A2(_17723_),
    .Y(_01731_),
    .B1(_17724_));
 sg13g2_nor2_1 _25644_ (.A(\u_inv.f_next[225] ),
    .B(net6998),
    .Y(_17725_));
 sg13g2_nor2_1 _25645_ (.A(net3203),
    .B(net6014),
    .Y(_17726_));
 sg13g2_a21oi_1 _25646_ (.A1(net6014),
    .A2(_17725_),
    .Y(_01732_),
    .B1(_17726_));
 sg13g2_nor2_1 _25647_ (.A(\u_inv.f_next[226] ),
    .B(net6999),
    .Y(_17727_));
 sg13g2_nor2_1 _25648_ (.A(net1746),
    .B(net6016),
    .Y(_17728_));
 sg13g2_a21oi_1 _25649_ (.A1(net6016),
    .A2(_17727_),
    .Y(_01733_),
    .B1(_17728_));
 sg13g2_nor2_1 _25650_ (.A(\u_inv.f_next[227] ),
    .B(net6999),
    .Y(_17729_));
 sg13g2_nor2_1 _25651_ (.A(net2167),
    .B(net6016),
    .Y(_17730_));
 sg13g2_a21oi_1 _25652_ (.A1(net6016),
    .A2(_17729_),
    .Y(_01734_),
    .B1(_17730_));
 sg13g2_nor2_1 _25653_ (.A(\u_inv.f_next[228] ),
    .B(net6999),
    .Y(_17731_));
 sg13g2_nor2_1 _25654_ (.A(net2902),
    .B(net6018),
    .Y(_17732_));
 sg13g2_a21oi_1 _25655_ (.A1(net6018),
    .A2(_17731_),
    .Y(_01735_),
    .B1(_17732_));
 sg13g2_nor2_1 _25656_ (.A(\u_inv.f_next[229] ),
    .B(net6999),
    .Y(_17733_));
 sg13g2_nor2_1 _25657_ (.A(net1842),
    .B(net6018),
    .Y(_17734_));
 sg13g2_a21oi_1 _25658_ (.A1(net6015),
    .A2(_17733_),
    .Y(_01736_),
    .B1(_17734_));
 sg13g2_nor2_1 _25659_ (.A(\u_inv.f_next[230] ),
    .B(net6999),
    .Y(_17735_));
 sg13g2_nor2_1 _25660_ (.A(net2855),
    .B(net6016),
    .Y(_17736_));
 sg13g2_a21oi_1 _25661_ (.A1(net6016),
    .A2(_17735_),
    .Y(_01737_),
    .B1(_17736_));
 sg13g2_nor2_1 _25662_ (.A(net3130),
    .B(net6998),
    .Y(_17737_));
 sg13g2_nor2_1 _25663_ (.A(net3196),
    .B(net6016),
    .Y(_17738_));
 sg13g2_a21oi_1 _25664_ (.A1(net6017),
    .A2(_17737_),
    .Y(_01738_),
    .B1(_17738_));
 sg13g2_nor2_1 _25665_ (.A(\u_inv.f_next[232] ),
    .B(net7008),
    .Y(_17739_));
 sg13g2_nor2_1 _25666_ (.A(net2884),
    .B(net6017),
    .Y(_17740_));
 sg13g2_a21oi_1 _25667_ (.A1(net6017),
    .A2(_17739_),
    .Y(_01739_),
    .B1(_17740_));
 sg13g2_nor2_1 _25668_ (.A(net2818),
    .B(net7008),
    .Y(_17741_));
 sg13g2_nor2_1 _25669_ (.A(net2919),
    .B(net6016),
    .Y(_17742_));
 sg13g2_a21oi_1 _25670_ (.A1(net6017),
    .A2(_17741_),
    .Y(_01740_),
    .B1(_17742_));
 sg13g2_nor2_1 _25671_ (.A(\u_inv.f_next[234] ),
    .B(net7008),
    .Y(_17743_));
 sg13g2_nor2_1 _25672_ (.A(net3276),
    .B(net6023),
    .Y(_17744_));
 sg13g2_a21oi_1 _25673_ (.A1(net6023),
    .A2(_17743_),
    .Y(_01741_),
    .B1(_17744_));
 sg13g2_nor2_1 _25674_ (.A(\u_inv.f_next[235] ),
    .B(net7008),
    .Y(_17745_));
 sg13g2_nor2_1 _25675_ (.A(net2146),
    .B(net6023),
    .Y(_17746_));
 sg13g2_a21oi_1 _25676_ (.A1(net6023),
    .A2(_17745_),
    .Y(_01742_),
    .B1(_17746_));
 sg13g2_nor2_1 _25677_ (.A(\u_inv.f_next[236] ),
    .B(net7008),
    .Y(_17747_));
 sg13g2_nor2_1 _25678_ (.A(net3029),
    .B(net6023),
    .Y(_17748_));
 sg13g2_a21oi_1 _25679_ (.A1(net6024),
    .A2(_17747_),
    .Y(_01743_),
    .B1(_17748_));
 sg13g2_nor2_1 _25680_ (.A(\u_inv.f_next[237] ),
    .B(net7008),
    .Y(_17749_));
 sg13g2_nor2_1 _25681_ (.A(net2140),
    .B(net6023),
    .Y(_17750_));
 sg13g2_a21oi_1 _25682_ (.A1(net6024),
    .A2(_17749_),
    .Y(_01744_),
    .B1(_17750_));
 sg13g2_nor2_1 _25683_ (.A(\u_inv.f_next[238] ),
    .B(net7010),
    .Y(_17751_));
 sg13g2_nor2_1 _25684_ (.A(net1940),
    .B(net6024),
    .Y(_17752_));
 sg13g2_a21oi_1 _25685_ (.A1(net6023),
    .A2(_17751_),
    .Y(_01745_),
    .B1(_17752_));
 sg13g2_nor2_1 _25686_ (.A(\u_inv.f_next[239] ),
    .B(net7008),
    .Y(_17753_));
 sg13g2_nor2_1 _25687_ (.A(net2908),
    .B(net6023),
    .Y(_17754_));
 sg13g2_a21oi_1 _25688_ (.A1(net6024),
    .A2(_17753_),
    .Y(_01746_),
    .B1(_17754_));
 sg13g2_nor2_1 _25689_ (.A(\u_inv.f_next[240] ),
    .B(net7010),
    .Y(_17755_));
 sg13g2_nor2_1 _25690_ (.A(net2642),
    .B(net6025),
    .Y(_17756_));
 sg13g2_a21oi_1 _25691_ (.A1(net6025),
    .A2(_17755_),
    .Y(_01747_),
    .B1(_17756_));
 sg13g2_nor2_1 _25692_ (.A(\u_inv.f_next[241] ),
    .B(net7008),
    .Y(_17757_));
 sg13g2_nor2_1 _25693_ (.A(net2332),
    .B(net6025),
    .Y(_17758_));
 sg13g2_a21oi_1 _25694_ (.A1(net6025),
    .A2(_17757_),
    .Y(_01748_),
    .B1(_17758_));
 sg13g2_nor2_1 _25695_ (.A(\u_inv.f_next[242] ),
    .B(net7011),
    .Y(_17759_));
 sg13g2_nor2_1 _25696_ (.A(net2724),
    .B(net6025),
    .Y(_17760_));
 sg13g2_a21oi_1 _25697_ (.A1(net6025),
    .A2(_17759_),
    .Y(_01749_),
    .B1(_17760_));
 sg13g2_nor2_1 _25698_ (.A(net1691),
    .B(net7011),
    .Y(_17761_));
 sg13g2_nor2_1 _25699_ (.A(net2697),
    .B(net6026),
    .Y(_17762_));
 sg13g2_a21oi_1 _25700_ (.A1(net6026),
    .A2(_17761_),
    .Y(_01750_),
    .B1(_17762_));
 sg13g2_nor2_1 _25701_ (.A(\u_inv.f_next[244] ),
    .B(net7011),
    .Y(_17763_));
 sg13g2_nor2_1 _25702_ (.A(net2680),
    .B(net6025),
    .Y(_17764_));
 sg13g2_a21oi_1 _25703_ (.A1(net6025),
    .A2(_17763_),
    .Y(_01751_),
    .B1(_17764_));
 sg13g2_nor2_1 _25704_ (.A(\u_inv.f_next[245] ),
    .B(net7011),
    .Y(_17765_));
 sg13g2_nor2_1 _25705_ (.A(net2231),
    .B(net6027),
    .Y(_17766_));
 sg13g2_a21oi_1 _25706_ (.A1(net6027),
    .A2(_17765_),
    .Y(_01752_),
    .B1(_17766_));
 sg13g2_nor2_1 _25707_ (.A(\u_inv.f_next[246] ),
    .B(net7012),
    .Y(_17767_));
 sg13g2_nor2_1 _25708_ (.A(net1913),
    .B(net6027),
    .Y(_17768_));
 sg13g2_a21oi_1 _25709_ (.A1(net6027),
    .A2(_17767_),
    .Y(_01753_),
    .B1(_17768_));
 sg13g2_nor2_1 _25710_ (.A(\u_inv.f_next[247] ),
    .B(net7011),
    .Y(_17769_));
 sg13g2_nor2_1 _25711_ (.A(net3055),
    .B(net6027),
    .Y(_17770_));
 sg13g2_a21oi_1 _25712_ (.A1(net6027),
    .A2(_17769_),
    .Y(_01754_),
    .B1(_17770_));
 sg13g2_nor2_1 _25713_ (.A(\u_inv.f_next[248] ),
    .B(net7011),
    .Y(_17771_));
 sg13g2_nor2_1 _25714_ (.A(net2688),
    .B(net6028),
    .Y(_17772_));
 sg13g2_a21oi_1 _25715_ (.A1(net6028),
    .A2(_17771_),
    .Y(_01755_),
    .B1(_17772_));
 sg13g2_nor2_1 _25716_ (.A(\u_inv.f_next[249] ),
    .B(net7012),
    .Y(_17773_));
 sg13g2_nor2_1 _25717_ (.A(net2857),
    .B(net6028),
    .Y(_17774_));
 sg13g2_a21oi_1 _25718_ (.A1(net6029),
    .A2(_17773_),
    .Y(_01756_),
    .B1(_17774_));
 sg13g2_nor2_1 _25719_ (.A(\u_inv.f_next[250] ),
    .B(net7012),
    .Y(_17775_));
 sg13g2_nor2_1 _25720_ (.A(net2165),
    .B(net6028),
    .Y(_17776_));
 sg13g2_a21oi_1 _25721_ (.A1(net6028),
    .A2(_17775_),
    .Y(_01757_),
    .B1(_17776_));
 sg13g2_nor2_1 _25722_ (.A(\u_inv.f_next[251] ),
    .B(net7012),
    .Y(_17777_));
 sg13g2_nor2_1 _25723_ (.A(net2623),
    .B(net6029),
    .Y(_17778_));
 sg13g2_a21oi_1 _25724_ (.A1(net6028),
    .A2(_17777_),
    .Y(_01758_),
    .B1(_17778_));
 sg13g2_nor2_1 _25725_ (.A(\u_inv.f_next[252] ),
    .B(net7013),
    .Y(_17779_));
 sg13g2_nor2_1 _25726_ (.A(net2526),
    .B(net6029),
    .Y(_17780_));
 sg13g2_a21oi_1 _25727_ (.A1(net6029),
    .A2(_17779_),
    .Y(_01759_),
    .B1(_17780_));
 sg13g2_nor2_1 _25728_ (.A(\u_inv.f_next[253] ),
    .B(net7016),
    .Y(_17781_));
 sg13g2_nor2_1 _25729_ (.A(net3072),
    .B(net6030),
    .Y(_17782_));
 sg13g2_a21oi_1 _25730_ (.A1(net6030),
    .A2(_17781_),
    .Y(_01760_),
    .B1(_17782_));
 sg13g2_nor2_1 _25731_ (.A(\u_inv.f_next[254] ),
    .B(net7011),
    .Y(_17783_));
 sg13g2_nor2_1 _25732_ (.A(net2660),
    .B(net6027),
    .Y(_17784_));
 sg13g2_a21oi_1 _25733_ (.A1(net6027),
    .A2(_17783_),
    .Y(_01761_),
    .B1(_17784_));
 sg13g2_nor2_1 _25734_ (.A(\u_inv.f_next[255] ),
    .B(net7011),
    .Y(_17785_));
 sg13g2_nor2_1 _25735_ (.A(net3214),
    .B(net6029),
    .Y(_17786_));
 sg13g2_a21oi_1 _25736_ (.A1(net6028),
    .A2(_17785_),
    .Y(_01762_),
    .B1(_17786_));
 sg13g2_nand3_1 _25737_ (.B(net7084),
    .C(net6030),
    .A(net2730),
    .Y(_17787_));
 sg13g2_o21ai_1 _25738_ (.B1(_17787_),
    .Y(_01763_),
    .A1(net7163),
    .A2(net6031));
 sg13g2_nor3_1 _25739_ (.A(net7246),
    .B(\u_inv.counter[4] ),
    .C(_02337_),
    .Y(_17788_));
 sg13g2_nor3_1 _25740_ (.A(\u_inv.counter[3] ),
    .B(\u_inv.counter[2] ),
    .C(_18255_),
    .Y(_17789_));
 sg13g2_nand4_1 _25741_ (.B(_19841_),
    .C(_17788_),
    .A(\u_inv.counter[1] ),
    .Y(_17790_),
    .D(_17789_));
 sg13g2_nor2_1 _25742_ (.A(\u_inv.counter[1] ),
    .B(_18255_),
    .Y(_17791_));
 sg13g2_nand4_1 _25743_ (.B(\u_inv.counter[2] ),
    .C(_17788_),
    .A(_18190_),
    .Y(_17792_),
    .D(_17791_));
 sg13g2_a22oi_1 _25744_ (.Y(_17793_),
    .B1(_17792_),
    .B2(net5976),
    .A2(_17790_),
    .A1(_02353_));
 sg13g2_nand2b_1 _25745_ (.Y(_17794_),
    .B(net5235),
    .A_N(_17793_));
 sg13g2_inv_1 _25746_ (.Y(_17795_),
    .A(_17794_));
 sg13g2_nand2_1 _25747_ (.Y(_01764_),
    .A(net6606),
    .B(_17794_));
 sg13g2_a21oi_1 _25748_ (.A1(net3669),
    .A2(net7016),
    .Y(_01765_),
    .B1(_17795_));
 sg13g2_nor2_2 _25749_ (.A(_24689_[0]),
    .B(net5132),
    .Y(_17796_));
 sg13g2_o21ai_1 _25750_ (.B1(net3412),
    .Y(_17797_),
    .A1(_24689_[0]),
    .A2(net5133));
 sg13g2_mux2_1 _25751_ (.A0(net5133),
    .A1(_17796_),
    .S(net3412),
    .X(_01766_));
 sg13g2_and2_1 _25752_ (.A(net3412),
    .B(net1221),
    .X(_17798_));
 sg13g2_nor2_1 _25753_ (.A(net7016),
    .B(_17798_),
    .Y(_17799_));
 sg13g2_nor2_1 _25754_ (.A(_17796_),
    .B(_17799_),
    .Y(_17800_));
 sg13g2_a21oi_1 _25755_ (.A1(_18340_),
    .A2(_17797_),
    .Y(_01767_),
    .B1(_17800_));
 sg13g2_a21oi_1 _25756_ (.A1(net5133),
    .A2(_17798_),
    .Y(_17801_),
    .B1(net1163));
 sg13g2_a21oi_1 _25757_ (.A1(net1163),
    .A2(_17800_),
    .Y(_01768_),
    .B1(_17801_));
 sg13g2_a21oi_1 _25758_ (.A1(net1163),
    .A2(_17798_),
    .Y(_17802_),
    .B1(net3121));
 sg13g2_nand3_1 _25759_ (.B(net3121),
    .C(_17798_),
    .A(net1163),
    .Y(_17803_));
 sg13g2_nor2b_1 _25760_ (.A(_17802_),
    .B_N(_17803_),
    .Y(_17804_));
 sg13g2_a22oi_1 _25761_ (.Y(_17805_),
    .B1(_17804_),
    .B2(net5133),
    .A2(_17796_),
    .A1(net3121));
 sg13g2_inv_1 _25762_ (.Y(_01769_),
    .A(_17805_));
 sg13g2_nor2_1 _25763_ (.A(_18342_),
    .B(_17803_),
    .Y(_17806_));
 sg13g2_xnor2_1 _25764_ (.Y(_17807_),
    .A(net2672),
    .B(_17803_));
 sg13g2_a22oi_1 _25765_ (.Y(_17808_),
    .B1(_17807_),
    .B2(net5131),
    .A2(_17796_),
    .A1(net2672));
 sg13g2_inv_1 _25766_ (.Y(_01770_),
    .A(_17808_));
 sg13g2_xnor2_1 _25767_ (.Y(_17809_),
    .A(_18343_),
    .B(_17806_));
 sg13g2_a22oi_1 _25768_ (.Y(_17810_),
    .B1(_17809_),
    .B2(net5131),
    .A2(_17796_),
    .A1(net3284));
 sg13g2_inv_1 _25769_ (.Y(_01771_),
    .A(_17810_));
 sg13g2_a21oi_1 _25770_ (.A1(net3284),
    .A2(_17806_),
    .Y(_17811_),
    .B1(net2421));
 sg13g2_and3_2 _25771_ (.X(_17812_),
    .A(net3284),
    .B(net2421),
    .C(_17806_));
 sg13g2_nor2_1 _25772_ (.A(_17811_),
    .B(_17812_),
    .Y(_17813_));
 sg13g2_a22oi_1 _25773_ (.Y(_17814_),
    .B1(_17813_),
    .B2(net5131),
    .A2(_17796_),
    .A1(net2421));
 sg13g2_inv_1 _25774_ (.Y(_01772_),
    .A(_17814_));
 sg13g2_nand2_1 _25775_ (.Y(_17815_),
    .A(net2592),
    .B(_17812_));
 sg13g2_xnor2_1 _25776_ (.Y(_17816_),
    .A(_18344_),
    .B(_17812_));
 sg13g2_a22oi_1 _25777_ (.Y(_17817_),
    .B1(_17816_),
    .B2(net5131),
    .A2(_17796_),
    .A1(net2592));
 sg13g2_inv_1 _25778_ (.Y(_01773_),
    .A(_17817_));
 sg13g2_xnor2_1 _25779_ (.Y(_17818_),
    .A(net3356),
    .B(_17815_));
 sg13g2_a22oi_1 _25780_ (.Y(_17819_),
    .B1(_17818_),
    .B2(net5131),
    .A2(_17796_),
    .A1(net3356));
 sg13g2_inv_1 _25781_ (.Y(_01774_),
    .A(_17819_));
 sg13g2_nand4_1 _25782_ (.B(net3356),
    .C(net5131),
    .A(net2592),
    .Y(_17820_),
    .D(_17812_));
 sg13g2_o21ai_1 _25783_ (.B1(net6606),
    .Y(_17821_),
    .A1(_18345_),
    .A2(_17820_));
 sg13g2_a21oi_1 _25784_ (.A1(_18345_),
    .A2(_17820_),
    .Y(_01775_),
    .B1(_17821_));
 sg13g2_xnor2_1 _25785_ (.Y(_17822_),
    .A(_18184_),
    .B(net5212));
 sg13g2_a22oi_1 _25786_ (.Y(_01776_),
    .B1(net6882),
    .B2(_17822_),
    .A2(net6442),
    .A1(_18184_));
 sg13g2_o21ai_1 _25787_ (.B1(net5242),
    .Y(_17823_),
    .A1(_18184_),
    .A2(net5956));
 sg13g2_nand2_1 _25788_ (.Y(_17824_),
    .A(\u_inv.delta_double[0] ),
    .B(_19813_));
 sg13g2_xor2_1 _25789_ (.B(_17824_),
    .A(net3420),
    .X(_17825_));
 sg13g2_or2_1 _25790_ (.X(_17826_),
    .B(_17825_),
    .A(_17823_));
 sg13g2_a21oi_1 _25791_ (.A1(_17823_),
    .A2(_17825_),
    .Y(_17827_),
    .B1(net6855));
 sg13g2_a22oi_1 _25792_ (.Y(_17828_),
    .B1(_17826_),
    .B2(_17827_),
    .A2(net6442),
    .A1(net3420));
 sg13g2_inv_1 _25793_ (.Y(_01777_),
    .A(_17828_));
 sg13g2_nand2_1 _25794_ (.Y(_17829_),
    .A(net1211),
    .B(net6443));
 sg13g2_o21ai_1 _25795_ (.B1(\u_inv.delta_reg[1] ),
    .Y(_17830_),
    .A1(\u_inv.delta_double[0] ),
    .A2(_19819_));
 sg13g2_xor2_1 _25796_ (.B(_17830_),
    .A(net1211),
    .X(_17831_));
 sg13g2_nor2_1 _25797_ (.A(_17826_),
    .B(_17831_),
    .Y(_17832_));
 sg13g2_a21o_1 _25798_ (.A2(_17831_),
    .A1(_17826_),
    .B1(net6855),
    .X(_17833_));
 sg13g2_o21ai_1 _25799_ (.B1(_17829_),
    .Y(_01778_),
    .A1(_17832_),
    .A2(_17833_));
 sg13g2_nand2_1 _25800_ (.Y(_17834_),
    .A(net1215),
    .B(net6443));
 sg13g2_nand3_1 _25801_ (.B(\u_inv.delta_reg[1] ),
    .C(\u_inv.delta_reg[2] ),
    .A(\u_inv.delta_double[0] ),
    .Y(_17835_));
 sg13g2_o21ai_1 _25802_ (.B1(_17835_),
    .Y(_17836_),
    .A1(_19814_),
    .A2(net6248));
 sg13g2_xnor2_1 _25803_ (.Y(_17837_),
    .A(net1215),
    .B(_17836_));
 sg13g2_nor2_1 _25804_ (.A(_17831_),
    .B(_17837_),
    .Y(_17838_));
 sg13g2_nor2b_1 _25805_ (.A(_17826_),
    .B_N(_17838_),
    .Y(_17839_));
 sg13g2_xor2_1 _25806_ (.B(_17837_),
    .A(_17832_),
    .X(_17840_));
 sg13g2_o21ai_1 _25807_ (.B1(_17834_),
    .Y(_01779_),
    .A1(net6856),
    .A2(_17840_));
 sg13g2_nand2_1 _25808_ (.Y(_17841_),
    .A(net1672),
    .B(net6442));
 sg13g2_nor2_1 _25809_ (.A(_18185_),
    .B(_17835_),
    .Y(_17842_));
 sg13g2_o21ai_1 _25810_ (.B1(_19815_),
    .Y(_17843_),
    .A1(net6341),
    .A2(_17842_));
 sg13g2_xnor2_1 _25811_ (.Y(_17844_),
    .A(net1672),
    .B(_17843_));
 sg13g2_nand2_1 _25812_ (.Y(_17845_),
    .A(_17838_),
    .B(_17844_));
 sg13g2_nor2_1 _25813_ (.A(_17826_),
    .B(_17845_),
    .Y(_17846_));
 sg13g2_o21ai_1 _25814_ (.B1(net6882),
    .Y(_17847_),
    .A1(_17839_),
    .A2(_17844_));
 sg13g2_o21ai_1 _25815_ (.B1(_17841_),
    .Y(_01780_),
    .A1(_17846_),
    .A2(_17847_));
 sg13g2_nand2_1 _25816_ (.Y(_17848_),
    .A(net1225),
    .B(net6442));
 sg13g2_a21oi_1 _25817_ (.A1(\u_inv.delta_reg[4] ),
    .A2(_17842_),
    .Y(_17849_),
    .B1(\u_inv.delta_reg[5] ));
 sg13g2_nand3_1 _25818_ (.B(\u_inv.delta_reg[4] ),
    .C(_17842_),
    .A(\u_inv.delta_reg[5] ),
    .Y(_17850_));
 sg13g2_nor2b_1 _25819_ (.A(_17849_),
    .B_N(_17850_),
    .Y(_17851_));
 sg13g2_o21ai_1 _25820_ (.B1(net1225),
    .Y(_17852_),
    .A1(\u_inv.delta_reg[4] ),
    .A2(_19815_));
 sg13g2_nor2_1 _25821_ (.A(_19813_),
    .B(_19816_),
    .Y(_17853_));
 sg13g2_a22oi_1 _25822_ (.Y(_17854_),
    .B1(_17852_),
    .B2(_17853_),
    .A2(_17851_),
    .A1(net6248));
 sg13g2_or3_1 _25823_ (.A(_17825_),
    .B(_17845_),
    .C(_17854_),
    .X(_17855_));
 sg13g2_xor2_1 _25824_ (.B(_17854_),
    .A(_17846_),
    .X(_17856_));
 sg13g2_o21ai_1 _25825_ (.B1(_17848_),
    .Y(_01781_),
    .A1(net6855),
    .A2(_17856_));
 sg13g2_nand2_1 _25826_ (.Y(_17857_),
    .A(net1171),
    .B(net6442));
 sg13g2_o21ai_1 _25827_ (.B1(_17850_),
    .Y(_17858_),
    .A1(_19813_),
    .A2(_19816_));
 sg13g2_xnor2_1 _25828_ (.Y(_17859_),
    .A(_18186_),
    .B(_17858_));
 sg13g2_nand2_1 _25829_ (.Y(_17860_),
    .A(_18184_),
    .B(\u_inv.delta_reg[1] ));
 sg13g2_nor4_1 _25830_ (.A(net5991),
    .B(_17845_),
    .C(_17854_),
    .D(_17860_),
    .Y(_17861_));
 sg13g2_a21oi_1 _25831_ (.A1(_17859_),
    .A2(_17861_),
    .Y(_17862_),
    .B1(net5956));
 sg13g2_nand2b_1 _25832_ (.Y(_17863_),
    .B(_17859_),
    .A_N(_17855_));
 sg13g2_a21oi_1 _25833_ (.A1(net5957),
    .A2(_17863_),
    .Y(_17864_),
    .B1(_17862_));
 sg13g2_inv_1 _25834_ (.Y(_17865_),
    .A(_17864_));
 sg13g2_nor3_1 _25835_ (.A(net5928),
    .B(_17855_),
    .C(_17859_),
    .Y(_17866_));
 sg13g2_a21oi_1 _25836_ (.A1(_17859_),
    .A2(_17865_),
    .Y(_17867_),
    .B1(_17866_));
 sg13g2_nand2_1 _25837_ (.Y(_17868_),
    .A(net5285),
    .B(_17867_));
 sg13g2_a21oi_1 _25838_ (.A1(_17861_),
    .A2(_17862_),
    .Y(_17869_),
    .B1(_17868_));
 sg13g2_o21ai_1 _25839_ (.B1(net6882),
    .Y(_17870_),
    .A1(net5285),
    .A2(_17859_));
 sg13g2_o21ai_1 _25840_ (.B1(_17857_),
    .Y(_01782_),
    .A1(_17869_),
    .A2(_17870_));
 sg13g2_a21oi_1 _25841_ (.A1(net5321),
    .A2(net5317),
    .Y(_17871_),
    .B1(_17865_));
 sg13g2_nor2_1 _25842_ (.A(_18186_),
    .B(_17850_),
    .Y(_17872_));
 sg13g2_a21oi_1 _25843_ (.A1(_19812_),
    .A2(_19817_),
    .Y(_17873_),
    .B1(_17872_));
 sg13g2_xnor2_1 _25844_ (.Y(_17874_),
    .A(net3095),
    .B(_17873_));
 sg13g2_nor2_1 _25845_ (.A(_17871_),
    .B(_17874_),
    .Y(_17875_));
 sg13g2_nand2_1 _25846_ (.Y(_17876_),
    .A(_17871_),
    .B(_17874_));
 sg13g2_nor2_1 _25847_ (.A(net6855),
    .B(_17875_),
    .Y(_17877_));
 sg13g2_a22oi_1 _25848_ (.Y(_17878_),
    .B1(_17876_),
    .B2(_17877_),
    .A2(net6442),
    .A1(net3095));
 sg13g2_inv_1 _25849_ (.Y(_01783_),
    .A(_17878_));
 sg13g2_nand2_1 _25850_ (.Y(_17879_),
    .A(net1342),
    .B(net6443));
 sg13g2_and2_1 _25851_ (.A(\u_inv.delta_reg[7] ),
    .B(_17872_),
    .X(_17880_));
 sg13g2_nor2_1 _25852_ (.A(_19813_),
    .B(_19818_),
    .Y(_17881_));
 sg13g2_nor2_1 _25853_ (.A(_17880_),
    .B(_17881_),
    .Y(_17882_));
 sg13g2_xnor2_1 _25854_ (.Y(_17883_),
    .A(net1342),
    .B(_17882_));
 sg13g2_nand3_1 _25855_ (.B(_17874_),
    .C(_17883_),
    .A(_17871_),
    .Y(_17884_));
 sg13g2_xor2_1 _25856_ (.B(_17883_),
    .A(_17876_),
    .X(_17885_));
 sg13g2_o21ai_1 _25857_ (.B1(_17879_),
    .Y(_01784_),
    .A1(net6855),
    .A2(_17885_));
 sg13g2_nand2_1 _25858_ (.Y(_17886_),
    .A(net1249),
    .B(net6443));
 sg13g2_a21oi_1 _25859_ (.A1(\u_inv.delta_reg[8] ),
    .A2(_17880_),
    .Y(_17887_),
    .B1(net1249));
 sg13g2_nand3_1 _25860_ (.B(net1249),
    .C(_17880_),
    .A(\u_inv.delta_reg[8] ),
    .Y(_17888_));
 sg13g2_nor2_1 _25861_ (.A(net6341),
    .B(_17887_),
    .Y(_17889_));
 sg13g2_a21oi_1 _25862_ (.A1(_17888_),
    .A2(_17889_),
    .Y(_17890_),
    .B1(_19819_));
 sg13g2_xnor2_1 _25863_ (.Y(_17891_),
    .A(_17884_),
    .B(_17890_));
 sg13g2_o21ai_1 _25864_ (.B1(_17886_),
    .Y(_01785_),
    .A1(net6855),
    .A2(_17891_));
 sg13g2_nor2_1 _25865_ (.A(_19808_),
    .B(net5197),
    .Y(_17892_));
 sg13g2_o21ai_1 _25866_ (.B1(net6608),
    .Y(_17893_),
    .A1(net7251),
    .A2(_17892_));
 sg13g2_a21oi_1 _25867_ (.A1(net7251),
    .A2(_17892_),
    .Y(_01786_),
    .B1(_17893_));
 sg13g2_nor2_1 _25868_ (.A(net1233),
    .B(net6679),
    .Y(_17894_));
 sg13g2_a21oi_1 _25869_ (.A1(_18255_),
    .A2(net6679),
    .Y(_01787_),
    .B1(_17894_));
 sg13g2_mux2_1 _25870_ (.A0(net2202),
    .A1(\u_inv.counter[1] ),
    .S(net6681),
    .X(_01788_));
 sg13g2_mux2_1 _25871_ (.A0(net2304),
    .A1(\u_inv.counter[2] ),
    .S(net6679),
    .X(_01789_));
 sg13g2_nor2_1 _25872_ (.A(net1212),
    .B(net6679),
    .Y(_17895_));
 sg13g2_a21oi_1 _25873_ (.A1(_18190_),
    .A2(net6679),
    .Y(_01790_),
    .B1(_17895_));
 sg13g2_nor2_1 _25874_ (.A(net1203),
    .B(net6678),
    .Y(_17896_));
 sg13g2_a21oi_1 _25875_ (.A1(_18189_),
    .A2(net6678),
    .Y(_01791_),
    .B1(_17896_));
 sg13g2_nor2_1 _25876_ (.A(net1188),
    .B(net6678),
    .Y(_17897_));
 sg13g2_a21oi_1 _25877_ (.A1(_18188_),
    .A2(net6678),
    .Y(_01792_),
    .B1(_17897_));
 sg13g2_mux2_1 _25878_ (.A0(net1878),
    .A1(net7249),
    .S(net6678),
    .X(_01793_));
 sg13g2_mux2_1 _25879_ (.A0(net1766),
    .A1(net7247),
    .S(net6678),
    .X(_01794_));
 sg13g2_mux2_1 _25880_ (.A0(net1735),
    .A1(net7246),
    .S(net6678),
    .X(_01795_));
 sg13g2_mux2_1 _25881_ (.A0(net1415),
    .A1(\u_inv.counter[9] ),
    .S(net6680),
    .X(_01796_));
 sg13g2_nand2_1 _25882_ (.Y(_17898_),
    .A(net7251),
    .B(net5223));
 sg13g2_a21oi_1 _25883_ (.A1(_18255_),
    .A2(net5155),
    .Y(_17899_),
    .B1(net7006));
 sg13g2_nand2_1 _25884_ (.Y(_17900_),
    .A(_17898_),
    .B(_17899_));
 sg13g2_nand2_1 _25885_ (.Y(_17901_),
    .A(net3692),
    .B(net6608));
 sg13g2_mux2_1 _25886_ (.A0(net3692),
    .A1(_17901_),
    .S(_17900_),
    .X(_17902_));
 sg13g2_inv_1 _25887_ (.Y(_01797_),
    .A(_17902_));
 sg13g2_o21ai_1 _25888_ (.B1(net3692),
    .Y(_17903_),
    .A1(net7251),
    .A2(net5239));
 sg13g2_a21oi_1 _25889_ (.A1(_17898_),
    .A2(_17903_),
    .Y(_17904_),
    .B1(net7006));
 sg13g2_nand2_1 _25890_ (.Y(_17905_),
    .A(net3756),
    .B(_17904_));
 sg13g2_and2_1 _25891_ (.A(net3756),
    .B(net6608),
    .X(_17906_));
 sg13g2_o21ai_1 _25892_ (.B1(_17905_),
    .Y(_17907_),
    .A1(_17904_),
    .A2(_17906_));
 sg13g2_inv_1 _25893_ (.Y(_01798_),
    .A(_17907_));
 sg13g2_nand3_1 _25894_ (.B(net6608),
    .C(_17905_),
    .A(net1618),
    .Y(_17908_));
 sg13g2_o21ai_1 _25895_ (.B1(_17908_),
    .Y(_01799_),
    .A1(net1618),
    .A2(_17905_));
 sg13g2_nand3_1 _25896_ (.B(\u_inv.counter[2] ),
    .C(\u_inv.counter[1] ),
    .A(\u_inv.counter[3] ),
    .Y(_17909_));
 sg13g2_nor2_1 _25897_ (.A(_18189_),
    .B(_17909_),
    .Y(_17910_));
 sg13g2_and2_1 _25898_ (.A(_18189_),
    .B(_17909_),
    .X(_17911_));
 sg13g2_nor3_1 _25899_ (.A(net5880),
    .B(_17910_),
    .C(_17911_),
    .Y(_17912_));
 sg13g2_or2_1 _25900_ (.X(_17913_),
    .B(_17909_),
    .A(_18255_));
 sg13g2_xnor2_1 _25901_ (.Y(_17914_),
    .A(net3636),
    .B(_17913_));
 sg13g2_nor2_1 _25902_ (.A(_18190_),
    .B(_02338_),
    .Y(_17915_));
 sg13g2_nor3_1 _25903_ (.A(_18189_),
    .B(_18190_),
    .C(_02338_),
    .Y(_17916_));
 sg13g2_xnor2_1 _25904_ (.Y(_17917_),
    .A(_18189_),
    .B(_17915_));
 sg13g2_a221oi_1 _25905_ (.B2(net5937),
    .C1(_17912_),
    .B1(_17917_),
    .A1(net5976),
    .Y(_17918_),
    .A2(_17914_));
 sg13g2_a21oi_1 _25906_ (.A1(net5245),
    .A2(_17918_),
    .Y(_17919_),
    .B1(net7006));
 sg13g2_o21ai_1 _25907_ (.B1(_17919_),
    .Y(_17920_),
    .A1(net5245),
    .A2(_17914_));
 sg13g2_o21ai_1 _25908_ (.B1(_17920_),
    .Y(_01800_),
    .A1(_18189_),
    .A2(_19809_));
 sg13g2_nor3_2 _25909_ (.A(_18188_),
    .B(_18189_),
    .C(_17909_),
    .Y(_17921_));
 sg13g2_o21ai_1 _25910_ (.B1(_17921_),
    .Y(_17922_),
    .A1(net7250),
    .A2(net6003));
 sg13g2_nand2_1 _25911_ (.Y(_17923_),
    .A(net5918),
    .B(_17922_));
 sg13g2_o21ai_1 _25912_ (.B1(_17910_),
    .Y(_17924_),
    .A1(net7250),
    .A2(net6003));
 sg13g2_nor3_1 _25913_ (.A(_18188_),
    .B(_18189_),
    .C(_17913_),
    .Y(_17925_));
 sg13g2_a21oi_1 _25914_ (.A1(net7250),
    .A2(_17910_),
    .Y(_17926_),
    .B1(net3639));
 sg13g2_nor2_1 _25915_ (.A(_17925_),
    .B(_17926_),
    .Y(_17927_));
 sg13g2_a21oi_1 _25916_ (.A1(_18188_),
    .A2(_17924_),
    .Y(_17928_),
    .B1(_17923_));
 sg13g2_nor2_1 _25917_ (.A(\u_inv.counter[5] ),
    .B(_17916_),
    .Y(_17929_));
 sg13g2_and2_1 _25918_ (.A(net3639),
    .B(_17916_),
    .X(_17930_));
 sg13g2_nor3_1 _25919_ (.A(net5919),
    .B(_17929_),
    .C(_17930_),
    .Y(_17931_));
 sg13g2_nor2_1 _25920_ (.A(_17928_),
    .B(_17931_),
    .Y(_17932_));
 sg13g2_a21oi_1 _25921_ (.A1(net5245),
    .A2(_17932_),
    .Y(_17933_),
    .B1(net7006));
 sg13g2_o21ai_1 _25922_ (.B1(_17933_),
    .Y(_17934_),
    .A1(net5245),
    .A2(_17927_));
 sg13g2_o21ai_1 _25923_ (.B1(_17934_),
    .Y(_01801_),
    .A1(_18188_),
    .A2(_19809_));
 sg13g2_nand2_1 _25924_ (.Y(_17935_),
    .A(net7248),
    .B(_19808_));
 sg13g2_nand3_1 _25925_ (.B(net7250),
    .C(_17921_),
    .A(net7248),
    .Y(_17936_));
 sg13g2_o21ai_1 _25926_ (.B1(_17936_),
    .Y(_17937_),
    .A1(net7248),
    .A2(_17925_));
 sg13g2_o21ai_1 _25927_ (.B1(_17923_),
    .Y(_17938_),
    .A1(net5919),
    .A2(_17930_));
 sg13g2_xor2_1 _25928_ (.B(_17938_),
    .A(net7248),
    .X(_17939_));
 sg13g2_mux2_1 _25929_ (.A0(_17937_),
    .A1(_17939_),
    .S(net5245),
    .X(_17940_));
 sg13g2_o21ai_1 _25930_ (.B1(_17935_),
    .Y(_01802_),
    .A1(net7007),
    .A2(_17940_));
 sg13g2_nand3_1 _25931_ (.B(net7249),
    .C(_17930_),
    .A(net7247),
    .Y(_17941_));
 sg13g2_a21o_1 _25932_ (.A2(_17930_),
    .A1(net7248),
    .B1(net7247),
    .X(_17942_));
 sg13g2_nand2_1 _25933_ (.Y(_17943_),
    .A(_17941_),
    .B(_17942_));
 sg13g2_and3_2 _25934_ (.X(_17944_),
    .A(net7247),
    .B(net7248),
    .C(_17921_));
 sg13g2_xor2_1 _25935_ (.B(_17936_),
    .A(net7247),
    .X(_17945_));
 sg13g2_a21oi_1 _25936_ (.A1(net7248),
    .A2(_17921_),
    .Y(_17946_),
    .B1(net7247));
 sg13g2_o21ai_1 _25937_ (.B1(net5884),
    .Y(_17947_),
    .A1(_17944_),
    .A2(_17946_));
 sg13g2_nand2_1 _25938_ (.Y(_17948_),
    .A(net7081),
    .B(_17947_));
 sg13g2_a221oi_1 _25939_ (.B2(net5155),
    .C1(_17948_),
    .B1(_17945_),
    .A1(net5223),
    .Y(_17949_),
    .A2(_17943_));
 sg13g2_a21o_1 _25940_ (.A2(_19808_),
    .A1(net7247),
    .B1(_17949_),
    .X(_01803_));
 sg13g2_nand4_1 _25941_ (.B(net7247),
    .C(net7249),
    .A(net7246),
    .Y(_17950_),
    .D(_17930_));
 sg13g2_xor2_1 _25942_ (.B(_17941_),
    .A(net7246),
    .X(_17951_));
 sg13g2_a21oi_1 _25943_ (.A1(net7250),
    .A2(_17944_),
    .Y(_17952_),
    .B1(net7246));
 sg13g2_nand3_1 _25944_ (.B(net7250),
    .C(_17944_),
    .A(\u_inv.counter[8] ),
    .Y(_17953_));
 sg13g2_nor2b_1 _25945_ (.A(_17952_),
    .B_N(_17953_),
    .Y(_17954_));
 sg13g2_xor2_1 _25946_ (.B(_17944_),
    .A(net7246),
    .X(_17955_));
 sg13g2_and3_1 _25947_ (.X(_17956_),
    .A(net5235),
    .B(net5884),
    .C(_17955_));
 sg13g2_a221oi_1 _25948_ (.B2(_17954_),
    .C1(_17956_),
    .B1(net5110),
    .A1(net7246),
    .Y(_17957_),
    .A2(_19808_));
 sg13g2_o21ai_1 _25949_ (.B1(_17957_),
    .Y(_01804_),
    .A1(net5124),
    .A2(net3758));
 sg13g2_xnor2_1 _25950_ (.Y(_17958_),
    .A(net3741),
    .B(_17953_));
 sg13g2_and3_1 _25951_ (.X(_17959_),
    .A(net7246),
    .B(_02346_),
    .C(_17944_));
 sg13g2_a221oi_1 _25952_ (.B2(net7081),
    .C1(_17959_),
    .B1(_17958_),
    .A1(net3741),
    .Y(_17960_),
    .A2(_19808_));
 sg13g2_o21ai_1 _25953_ (.B1(net3742),
    .Y(_01805_),
    .A1(net5124),
    .A2(_17950_));
 sg13g2_mux2_1 _25954_ (.A0(net1306),
    .A1(\shift_reg[16] ),
    .S(net6952),
    .X(_01806_));
 sg13g2_mux2_1 _25955_ (.A0(net1924),
    .A1(\shift_reg[17] ),
    .S(net6958),
    .X(_01807_));
 sg13g2_mux2_1 _25956_ (.A0(net1537),
    .A1(\shift_reg[18] ),
    .S(net6958),
    .X(_01808_));
 sg13g2_mux2_1 _25957_ (.A0(net1648),
    .A1(\shift_reg[19] ),
    .S(net6959),
    .X(_01809_));
 sg13g2_mux2_1 _25958_ (.A0(net1295),
    .A1(\shift_reg[20] ),
    .S(net6959),
    .X(_01810_));
 sg13g2_mux2_1 _25959_ (.A0(net1888),
    .A1(\shift_reg[21] ),
    .S(net6959),
    .X(_01811_));
 sg13g2_mux2_1 _25960_ (.A0(net1567),
    .A1(\shift_reg[22] ),
    .S(net6959),
    .X(_01812_));
 sg13g2_mux2_1 _25961_ (.A0(net1760),
    .A1(\shift_reg[23] ),
    .S(net6962),
    .X(_01813_));
 sg13g2_mux2_1 _25962_ (.A0(net1293),
    .A1(\shift_reg[24] ),
    .S(net6962),
    .X(_01814_));
 sg13g2_mux2_1 _25963_ (.A0(net1391),
    .A1(\shift_reg[25] ),
    .S(net6962),
    .X(_01815_));
 sg13g2_mux2_1 _25964_ (.A0(net1331),
    .A1(\shift_reg[26] ),
    .S(net6962),
    .X(_01816_));
 sg13g2_mux2_1 _25965_ (.A0(net1448),
    .A1(\shift_reg[27] ),
    .S(net6962),
    .X(_01817_));
 sg13g2_mux2_1 _25966_ (.A0(net1274),
    .A1(\shift_reg[28] ),
    .S(net6962),
    .X(_01818_));
 sg13g2_mux2_1 _25967_ (.A0(net1694),
    .A1(\shift_reg[29] ),
    .S(net6964),
    .X(_01819_));
 sg13g2_mux2_1 _25968_ (.A0(net1302),
    .A1(\shift_reg[30] ),
    .S(net6964),
    .X(_01820_));
 sg13g2_mux2_1 _25969_ (.A0(net1612),
    .A1(\shift_reg[31] ),
    .S(net6965),
    .X(_01821_));
 sg13g2_mux2_1 _25970_ (.A0(net1870),
    .A1(\shift_reg[32] ),
    .S(net6965),
    .X(_01822_));
 sg13g2_mux2_1 _25971_ (.A0(net1452),
    .A1(\shift_reg[33] ),
    .S(net6965),
    .X(_01823_));
 sg13g2_mux2_1 _25972_ (.A0(net1369),
    .A1(\shift_reg[34] ),
    .S(net6965),
    .X(_01824_));
 sg13g2_mux2_1 _25973_ (.A0(net2053),
    .A1(\shift_reg[35] ),
    .S(net6966),
    .X(_01825_));
 sg13g2_mux2_1 _25974_ (.A0(net1375),
    .A1(\shift_reg[36] ),
    .S(net6966),
    .X(_01826_));
 sg13g2_mux2_1 _25975_ (.A0(net1692),
    .A1(\shift_reg[37] ),
    .S(net6966),
    .X(_01827_));
 sg13g2_mux2_1 _25976_ (.A0(net1509),
    .A1(\shift_reg[38] ),
    .S(net6967),
    .X(_01828_));
 sg13g2_mux2_1 _25977_ (.A0(net1335),
    .A1(\shift_reg[39] ),
    .S(net6968),
    .X(_01829_));
 sg13g2_mux2_1 _25978_ (.A0(net1450),
    .A1(\shift_reg[40] ),
    .S(net6966),
    .X(_01830_));
 sg13g2_mux2_1 _25979_ (.A0(net1557),
    .A1(\shift_reg[41] ),
    .S(net6969),
    .X(_01831_));
 sg13g2_mux2_1 _25980_ (.A0(net1343),
    .A1(\shift_reg[42] ),
    .S(net6970),
    .X(_01832_));
 sg13g2_mux2_1 _25981_ (.A0(net1318),
    .A1(\shift_reg[43] ),
    .S(net6975),
    .X(_01833_));
 sg13g2_mux2_1 _25982_ (.A0(net1379),
    .A1(\shift_reg[44] ),
    .S(net6975),
    .X(_01834_));
 sg13g2_mux2_1 _25983_ (.A0(net1299),
    .A1(\shift_reg[45] ),
    .S(net6975),
    .X(_01835_));
 sg13g2_mux2_1 _25984_ (.A0(net1744),
    .A1(\shift_reg[46] ),
    .S(net6973),
    .X(_01836_));
 sg13g2_mux2_1 _25985_ (.A0(net1500),
    .A1(\shift_reg[47] ),
    .S(net6973),
    .X(_01837_));
 sg13g2_mux2_1 _25986_ (.A0(net1268),
    .A1(\shift_reg[48] ),
    .S(net6973),
    .X(_01838_));
 sg13g2_mux2_1 _25987_ (.A0(net1420),
    .A1(\shift_reg[49] ),
    .S(net6973),
    .X(_01839_));
 sg13g2_mux2_1 _25988_ (.A0(net1345),
    .A1(\shift_reg[50] ),
    .S(net6973),
    .X(_01840_));
 sg13g2_mux2_1 _25989_ (.A0(net1256),
    .A1(\shift_reg[51] ),
    .S(net6973),
    .X(_01841_));
 sg13g2_mux2_1 _25990_ (.A0(net1264),
    .A1(\shift_reg[52] ),
    .S(net6973),
    .X(_01842_));
 sg13g2_mux2_1 _25991_ (.A0(net1808),
    .A1(\shift_reg[53] ),
    .S(net6974),
    .X(_01843_));
 sg13g2_mux2_1 _25992_ (.A0(net1351),
    .A1(\shift_reg[54] ),
    .S(net6977),
    .X(_01844_));
 sg13g2_mux2_1 _25993_ (.A0(net1304),
    .A1(\shift_reg[55] ),
    .S(net6977),
    .X(_01845_));
 sg13g2_mux2_1 _25994_ (.A0(net1590),
    .A1(\shift_reg[56] ),
    .S(net6977),
    .X(_01846_));
 sg13g2_mux2_1 _25995_ (.A0(net2151),
    .A1(\shift_reg[57] ),
    .S(net6973),
    .X(_01847_));
 sg13g2_mux2_1 _25996_ (.A0(net1755),
    .A1(\shift_reg[58] ),
    .S(net6977),
    .X(_01848_));
 sg13g2_mux2_1 _25997_ (.A0(net1599),
    .A1(\shift_reg[59] ),
    .S(net6977),
    .X(_01849_));
 sg13g2_mux2_1 _25998_ (.A0(net1411),
    .A1(\shift_reg[60] ),
    .S(net6977),
    .X(_01850_));
 sg13g2_mux2_1 _25999_ (.A0(net1876),
    .A1(\shift_reg[61] ),
    .S(net6977),
    .X(_01851_));
 sg13g2_mux2_1 _26000_ (.A0(net1349),
    .A1(\shift_reg[62] ),
    .S(net6978),
    .X(_01852_));
 sg13g2_mux2_1 _26001_ (.A0(net1523),
    .A1(\shift_reg[63] ),
    .S(net6978),
    .X(_01853_));
 sg13g2_mux2_1 _26002_ (.A0(net1262),
    .A1(\shift_reg[64] ),
    .S(net6978),
    .X(_01854_));
 sg13g2_mux2_1 _26003_ (.A0(net1477),
    .A1(\shift_reg[65] ),
    .S(net6978),
    .X(_01855_));
 sg13g2_mux2_1 _26004_ (.A0(net1492),
    .A1(\shift_reg[66] ),
    .S(net6978),
    .X(_01856_));
 sg13g2_mux2_1 _26005_ (.A0(net1490),
    .A1(\shift_reg[67] ),
    .S(net6979),
    .X(_01857_));
 sg13g2_mux2_1 _26006_ (.A0(net1541),
    .A1(\shift_reg[68] ),
    .S(net6979),
    .X(_01858_));
 sg13g2_mux2_1 _26007_ (.A0(net1890),
    .A1(\shift_reg[69] ),
    .S(net6978),
    .X(_01859_));
 sg13g2_mux2_1 _26008_ (.A0(net1467),
    .A1(\shift_reg[70] ),
    .S(net6979),
    .X(_01860_));
 sg13g2_mux2_1 _26009_ (.A0(net1966),
    .A1(\shift_reg[71] ),
    .S(net6990),
    .X(_01861_));
 sg13g2_mux2_1 _26010_ (.A0(net1373),
    .A1(\shift_reg[72] ),
    .S(net6990),
    .X(_01862_));
 sg13g2_mux2_1 _26011_ (.A0(net1597),
    .A1(\shift_reg[73] ),
    .S(net6990),
    .X(_01863_));
 sg13g2_mux2_1 _26012_ (.A0(net1572),
    .A1(\shift_reg[74] ),
    .S(net6979),
    .X(_01864_));
 sg13g2_mux2_1 _26013_ (.A0(net1465),
    .A1(\shift_reg[75] ),
    .S(net6990),
    .X(_01865_));
 sg13g2_mux2_1 _26014_ (.A0(net1670),
    .A1(\shift_reg[76] ),
    .S(net6978),
    .X(_01866_));
 sg13g2_mux2_1 _26015_ (.A0(net1594),
    .A1(\shift_reg[77] ),
    .S(net6990),
    .X(_01867_));
 sg13g2_mux2_1 _26016_ (.A0(net1825),
    .A1(\shift_reg[78] ),
    .S(net6990),
    .X(_01868_));
 sg13g2_mux2_1 _26017_ (.A0(net1417),
    .A1(\shift_reg[79] ),
    .S(net6990),
    .X(_01869_));
 sg13g2_mux2_1 _26018_ (.A0(net1616),
    .A1(\shift_reg[80] ),
    .S(net6985),
    .X(_01870_));
 sg13g2_mux2_1 _26019_ (.A0(net1737),
    .A1(\shift_reg[81] ),
    .S(net6987),
    .X(_01871_));
 sg13g2_mux2_1 _26020_ (.A0(net1601),
    .A1(\shift_reg[82] ),
    .S(net6985),
    .X(_01872_));
 sg13g2_mux2_1 _26021_ (.A0(net1757),
    .A1(\shift_reg[83] ),
    .S(net6985),
    .X(_01873_));
 sg13g2_mux2_1 _26022_ (.A0(net1951),
    .A1(\shift_reg[84] ),
    .S(net6985),
    .X(_01874_));
 sg13g2_mux2_1 _26023_ (.A0(net1780),
    .A1(\shift_reg[85] ),
    .S(net6987),
    .X(_01875_));
 sg13g2_mux2_1 _26024_ (.A0(net1829),
    .A1(\shift_reg[86] ),
    .S(net6985),
    .X(_01876_));
 sg13g2_mux2_1 _26025_ (.A0(net1584),
    .A1(\shift_reg[87] ),
    .S(net6985),
    .X(_01877_));
 sg13g2_mux2_1 _26026_ (.A0(net2085),
    .A1(\shift_reg[88] ),
    .S(net6986),
    .X(_01878_));
 sg13g2_mux2_1 _26027_ (.A0(net1471),
    .A1(\shift_reg[89] ),
    .S(net6986),
    .X(_01879_));
 sg13g2_mux2_1 _26028_ (.A0(net2153),
    .A1(\shift_reg[90] ),
    .S(net6986),
    .X(_01880_));
 sg13g2_mux2_1 _26029_ (.A0(net1675),
    .A1(\shift_reg[91] ),
    .S(net6986),
    .X(_01881_));
 sg13g2_mux2_1 _26030_ (.A0(net2188),
    .A1(\shift_reg[92] ),
    .S(net6985),
    .X(_01882_));
 sg13g2_mux2_1 _26031_ (.A0(net1827),
    .A1(\shift_reg[93] ),
    .S(net6986),
    .X(_01883_));
 sg13g2_mux2_1 _26032_ (.A0(net2003),
    .A1(\shift_reg[94] ),
    .S(net6987),
    .X(_01884_));
 sg13g2_mux2_1 _26033_ (.A0(net1553),
    .A1(\shift_reg[95] ),
    .S(net6985),
    .X(_01885_));
 sg13g2_mux2_1 _26034_ (.A0(net1791),
    .A1(\shift_reg[96] ),
    .S(net6986),
    .X(_01886_));
 sg13g2_mux2_1 _26035_ (.A0(net1815),
    .A1(\shift_reg[97] ),
    .S(net6986),
    .X(_01887_));
 sg13g2_mux2_1 _26036_ (.A0(net1771),
    .A1(\shift_reg[98] ),
    .S(net6986),
    .X(_01888_));
 sg13g2_mux2_1 _26037_ (.A0(net1423),
    .A1(\shift_reg[99] ),
    .S(net6988),
    .X(_01889_));
 sg13g2_mux2_1 _26038_ (.A0(net1358),
    .A1(\shift_reg[100] ),
    .S(net6988),
    .X(_01890_));
 sg13g2_mux2_1 _26039_ (.A0(net1934),
    .A1(\shift_reg[101] ),
    .S(net6989),
    .X(_01891_));
 sg13g2_mux2_1 _26040_ (.A0(net1614),
    .A1(\shift_reg[102] ),
    .S(net6989),
    .X(_01892_));
 sg13g2_mux2_1 _26041_ (.A0(net1371),
    .A1(\shift_reg[103] ),
    .S(net6989),
    .X(_01893_));
 sg13g2_mux2_1 _26042_ (.A0(net1460),
    .A1(\shift_reg[104] ),
    .S(net6989),
    .X(_01894_));
 sg13g2_mux2_1 _26043_ (.A0(net1435),
    .A1(\shift_reg[105] ),
    .S(net6988),
    .X(_01895_));
 sg13g2_mux2_1 _26044_ (.A0(net1719),
    .A1(\shift_reg[106] ),
    .S(net6989),
    .X(_01896_));
 sg13g2_mux2_1 _26045_ (.A0(net1526),
    .A1(\shift_reg[107] ),
    .S(net6988),
    .X(_01897_));
 sg13g2_mux2_1 _26046_ (.A0(net1533),
    .A1(\shift_reg[108] ),
    .S(net6988),
    .X(_01898_));
 sg13g2_mux2_1 _26047_ (.A0(net2087),
    .A1(\shift_reg[109] ),
    .S(net6988),
    .X(_01899_));
 sg13g2_mux2_1 _26048_ (.A0(net1608),
    .A1(\shift_reg[110] ),
    .S(net6988),
    .X(_01900_));
 sg13g2_inv_1 _26049_ (.Y(_17961_),
    .A(net3677));
 sg13g2_inv_1 _26050_ (.Y(_17962_),
    .A(net3633));
 sg13g2_inv_2 _26051_ (.Y(_17963_),
    .A(net3368));
 sg13g2_inv_1 _26052_ (.Y(_17964_),
    .A(net3409));
 sg13g2_inv_1 _26053_ (.Y(_17965_),
    .A(net3691));
 sg13g2_inv_1 _26054_ (.Y(_17966_),
    .A(net3683));
 sg13g2_inv_1 _26055_ (.Y(_17967_),
    .A(net3674));
 sg13g2_inv_1 _26056_ (.Y(_17968_),
    .A(\u_inv.f_next[243] ));
 sg13g2_inv_1 _26057_ (.Y(_17969_),
    .A(net3722));
 sg13g2_inv_1 _26058_ (.Y(_17970_),
    .A(\u_inv.f_next[241] ));
 sg13g2_inv_1 _26059_ (.Y(_17971_),
    .A(\u_inv.f_next[238] ));
 sg13g2_inv_1 _26060_ (.Y(_17972_),
    .A(net3535));
 sg13g2_inv_1 _26061_ (.Y(_17973_),
    .A(\u_inv.f_next[235] ));
 sg13g2_inv_1 _26062_ (.Y(_17974_),
    .A(net3491));
 sg13g2_inv_1 _26063_ (.Y(_17975_),
    .A(\u_inv.f_next[228] ));
 sg13g2_inv_1 _26064_ (.Y(_17976_),
    .A(\u_inv.f_next[225] ));
 sg13g2_inv_1 _26065_ (.Y(_17977_),
    .A(net3613));
 sg13g2_inv_1 _26066_ (.Y(_17978_),
    .A(net3676));
 sg13g2_inv_1 _26067_ (.Y(_17979_),
    .A(\u_inv.f_next[219] ));
 sg13g2_inv_2 _26068_ (.Y(_17980_),
    .A(net2634));
 sg13g2_inv_1 _26069_ (.Y(_17981_),
    .A(\u_inv.f_next[216] ));
 sg13g2_inv_1 _26070_ (.Y(_17982_),
    .A(net3634));
 sg13g2_inv_1 _26071_ (.Y(_17983_),
    .A(\u_inv.f_next[213] ));
 sg13g2_inv_1 _26072_ (.Y(_17984_),
    .A(net3586));
 sg13g2_inv_1 _26073_ (.Y(_17985_),
    .A(net3655));
 sg13g2_inv_1 _26074_ (.Y(_17986_),
    .A(net3703));
 sg13g2_inv_1 _26075_ (.Y(_17987_),
    .A(\u_inv.f_next[207] ));
 sg13g2_inv_1 _26076_ (.Y(_17988_),
    .A(\u_inv.f_next[205] ));
 sg13g2_inv_1 _26077_ (.Y(_17989_),
    .A(\u_inv.f_next[203] ));
 sg13g2_inv_1 _26078_ (.Y(_17990_),
    .A(net3313));
 sg13g2_inv_1 _26079_ (.Y(_17991_),
    .A(net3596));
 sg13g2_inv_1 _26080_ (.Y(_17992_),
    .A(\u_inv.f_next[198] ));
 sg13g2_inv_1 _26081_ (.Y(_17993_),
    .A(net3662));
 sg13g2_inv_1 _26082_ (.Y(_17994_),
    .A(net3670));
 sg13g2_inv_2 _26083_ (.Y(_17995_),
    .A(net3612));
 sg13g2_inv_1 _26084_ (.Y(_17996_),
    .A(net3546));
 sg13g2_inv_1 _26085_ (.Y(_17997_),
    .A(net3682));
 sg13g2_inv_1 _26086_ (.Y(_17998_),
    .A(\u_inv.f_next[191] ));
 sg13g2_inv_1 _26087_ (.Y(_17999_),
    .A(\u_inv.f_next[190] ));
 sg13g2_inv_1 _26088_ (.Y(_18000_),
    .A(net3350));
 sg13g2_inv_1 _26089_ (.Y(_18001_),
    .A(net3502));
 sg13g2_inv_1 _26090_ (.Y(_18002_),
    .A(net3513));
 sg13g2_inv_1 _26091_ (.Y(_18003_),
    .A(net3698));
 sg13g2_inv_1 _26092_ (.Y(_18004_),
    .A(net2883));
 sg13g2_inv_2 _26093_ (.Y(_18005_),
    .A(net2850));
 sg13g2_inv_1 _26094_ (.Y(_18006_),
    .A(net2716));
 sg13g2_inv_1 _26095_ (.Y(_18007_),
    .A(\u_inv.f_next[179] ));
 sg13g2_inv_1 _26096_ (.Y(_18008_),
    .A(net2064));
 sg13g2_inv_1 _26097_ (.Y(_18009_),
    .A(net3729));
 sg13g2_inv_1 _26098_ (.Y(_18010_),
    .A(net2493));
 sg13g2_inv_1 _26099_ (.Y(_18011_),
    .A(net3348));
 sg13g2_inv_1 _26100_ (.Y(_18012_),
    .A(net3217));
 sg13g2_inv_1 _26101_ (.Y(_18013_),
    .A(\u_inv.f_next[171] ));
 sg13g2_inv_1 _26102_ (.Y(_18014_),
    .A(net2848));
 sg13g2_inv_1 _26103_ (.Y(_18015_),
    .A(net3460));
 sg13g2_inv_1 _26104_ (.Y(_18016_),
    .A(\u_inv.f_next[165] ));
 sg13g2_inv_1 _26105_ (.Y(_18017_),
    .A(net3006));
 sg13g2_inv_1 _26106_ (.Y(_18018_),
    .A(net3619));
 sg13g2_inv_1 _26107_ (.Y(_18019_),
    .A(net3694));
 sg13g2_inv_1 _26108_ (.Y(_18020_),
    .A(net3000));
 sg13g2_inv_1 _26109_ (.Y(_18021_),
    .A(net3624));
 sg13g2_inv_1 _26110_ (.Y(_18022_),
    .A(\u_inv.f_next[153] ));
 sg13g2_inv_1 _26111_ (.Y(_18023_),
    .A(net3554));
 sg13g2_inv_1 _26112_ (.Y(_18024_),
    .A(\u_inv.f_next[150] ));
 sg13g2_inv_2 _26113_ (.Y(_18025_),
    .A(net3689));
 sg13g2_inv_1 _26114_ (.Y(_18026_),
    .A(net3706));
 sg13g2_inv_1 _26115_ (.Y(_18027_),
    .A(net3386));
 sg13g2_inv_1 _26116_ (.Y(_18028_),
    .A(net3435));
 sg13g2_inv_1 _26117_ (.Y(_18029_),
    .A(net3645));
 sg13g2_inv_1 _26118_ (.Y(_18030_),
    .A(\u_inv.f_next[139] ));
 sg13g2_inv_1 _26119_ (.Y(_18031_),
    .A(net3617));
 sg13g2_inv_1 _26120_ (.Y(_18032_),
    .A(net3349));
 sg13g2_inv_1 _26121_ (.Y(_18033_),
    .A(net3187));
 sg13g2_inv_1 _26122_ (.Y(_18034_),
    .A(net3679));
 sg13g2_inv_1 _26123_ (.Y(_18035_),
    .A(net3646));
 sg13g2_inv_1 _26124_ (.Y(_18036_),
    .A(net3686));
 sg13g2_inv_1 _26125_ (.Y(_18037_),
    .A(net3599));
 sg13g2_inv_1 _26126_ (.Y(_18038_),
    .A(net3603));
 sg13g2_inv_1 _26127_ (.Y(_18039_),
    .A(\u_inv.f_next[121] ));
 sg13g2_inv_1 _26128_ (.Y(_18040_),
    .A(net3037));
 sg13g2_inv_2 _26129_ (.Y(_18041_),
    .A(net3473));
 sg13g2_inv_1 _26130_ (.Y(_18042_),
    .A(net3509));
 sg13g2_inv_1 _26131_ (.Y(_18043_),
    .A(net3266));
 sg13g2_inv_1 _26132_ (.Y(_18044_),
    .A(net3656));
 sg13g2_inv_1 _26133_ (.Y(_18045_),
    .A(net3298));
 sg13g2_inv_1 _26134_ (.Y(_18046_),
    .A(net3054));
 sg13g2_inv_1 _26135_ (.Y(_18047_),
    .A(net3553));
 sg13g2_inv_1 _26136_ (.Y(_18048_),
    .A(net3684));
 sg13g2_inv_1 _26137_ (.Y(_18049_),
    .A(\u_inv.f_next[105] ));
 sg13g2_inv_1 _26138_ (.Y(_18050_),
    .A(net2580));
 sg13g2_inv_1 _26139_ (.Y(_18051_),
    .A(net3292));
 sg13g2_inv_1 _26140_ (.Y(_18052_),
    .A(net2846));
 sg13g2_inv_1 _26141_ (.Y(_18053_),
    .A(\u_inv.f_next[91] ));
 sg13g2_inv_1 _26142_ (.Y(_18054_),
    .A(net2939));
 sg13g2_inv_1 _26143_ (.Y(_18055_),
    .A(net3701));
 sg13g2_inv_1 _26144_ (.Y(_18056_),
    .A(\u_inv.f_next[87] ));
 sg13g2_inv_1 _26145_ (.Y(_18057_),
    .A(net3481));
 sg13g2_inv_1 _26146_ (.Y(_18058_),
    .A(net3726));
 sg13g2_inv_1 _26147_ (.Y(_18059_),
    .A(net3392));
 sg13g2_inv_1 _26148_ (.Y(_18060_),
    .A(\u_inv.f_next[81] ));
 sg13g2_inv_1 _26149_ (.Y(_18061_),
    .A(\u_inv.f_next[80] ));
 sg13g2_inv_1 _26150_ (.Y(_18062_),
    .A(net3650));
 sg13g2_inv_1 _26151_ (.Y(_18063_),
    .A(net3434));
 sg13g2_inv_1 _26152_ (.Y(_18064_),
    .A(net3718));
 sg13g2_inv_1 _26153_ (.Y(_18065_),
    .A(net3614));
 sg13g2_inv_1 _26154_ (.Y(_18066_),
    .A(net3651));
 sg13g2_inv_1 _26155_ (.Y(_18067_),
    .A(net3658));
 sg13g2_inv_1 _26156_ (.Y(_18068_),
    .A(net3372));
 sg13g2_inv_1 _26157_ (.Y(_18069_),
    .A(net3560));
 sg13g2_inv_1 _26158_ (.Y(_18070_),
    .A(net3488));
 sg13g2_inv_1 _26159_ (.Y(_18071_),
    .A(net3649));
 sg13g2_inv_1 _26160_ (.Y(_18072_),
    .A(net3715));
 sg13g2_inv_1 _26161_ (.Y(_18073_),
    .A(net3589));
 sg13g2_inv_1 _26162_ (.Y(_18074_),
    .A(\u_inv.f_next[55] ));
 sg13g2_inv_1 _26163_ (.Y(_18075_),
    .A(net3667));
 sg13g2_inv_1 _26164_ (.Y(_18076_),
    .A(net3485));
 sg13g2_inv_1 _26165_ (.Y(_18077_),
    .A(net3135));
 sg13g2_inv_2 _26166_ (.Y(_18078_),
    .A(net3588));
 sg13g2_inv_1 _26167_ (.Y(_18079_),
    .A(\u_inv.f_next[45] ));
 sg13g2_inv_1 _26168_ (.Y(_18080_),
    .A(net2783));
 sg13g2_inv_1 _26169_ (.Y(_18081_),
    .A(net2216));
 sg13g2_inv_1 _26170_ (.Y(_18082_),
    .A(net3436));
 sg13g2_inv_1 _26171_ (.Y(_18083_),
    .A(net3083));
 sg13g2_inv_1 _26172_ (.Y(_18084_),
    .A(net3312));
 sg13g2_inv_1 _26173_ (.Y(_18085_),
    .A(net2760));
 sg13g2_inv_1 _26174_ (.Y(_18086_),
    .A(net3411));
 sg13g2_inv_1 _26175_ (.Y(_18087_),
    .A(net3719));
 sg13g2_inv_1 _26176_ (.Y(_18088_),
    .A(net3642));
 sg13g2_inv_1 _26177_ (.Y(_18089_),
    .A(net3595));
 sg13g2_inv_1 _26178_ (.Y(_18090_),
    .A(net3628));
 sg13g2_inv_1 _26179_ (.Y(_18091_),
    .A(\u_inv.f_next[15] ));
 sg13g2_inv_1 _26180_ (.Y(_18092_),
    .A(net3047));
 sg13g2_inv_1 _26181_ (.Y(_18093_),
    .A(net3709));
 sg13g2_inv_1 _26182_ (.Y(_18094_),
    .A(net3022));
 sg13g2_inv_1 _26183_ (.Y(_18095_),
    .A(\u_inv.f_next[9] ));
 sg13g2_inv_2 _26184_ (.Y(_18096_),
    .A(net1753));
 sg13g2_inv_1 _26185_ (.Y(_18097_),
    .A(net3331));
 sg13g2_inv_1 _26186_ (.Y(_18098_),
    .A(net3564));
 sg13g2_inv_8 _26187_ (.Y(_18099_),
    .A(net7308));
 sg13g2_inv_1 _26188_ (.Y(_18100_),
    .A(\u_inv.d_next[256] ));
 sg13g2_inv_1 _26189_ (.Y(_18101_),
    .A(\u_inv.d_next[255] ));
 sg13g2_inv_1 _26190_ (.Y(_18102_),
    .A(\u_inv.d_next[251] ));
 sg13g2_inv_1 _26191_ (.Y(_18103_),
    .A(\u_inv.d_next[247] ));
 sg13g2_inv_1 _26192_ (.Y(_18104_),
    .A(net7295));
 sg13g2_inv_1 _26193_ (.Y(_18105_),
    .A(\u_inv.d_next[242] ));
 sg13g2_inv_1 _26194_ (.Y(_18106_),
    .A(net2126));
 sg13g2_inv_1 _26195_ (.Y(_18107_),
    .A(\u_inv.d_next[227] ));
 sg13g2_inv_2 _26196_ (.Y(_18108_),
    .A(net3070));
 sg13g2_inv_1 _26197_ (.Y(_18109_),
    .A(\u_inv.d_next[221] ));
 sg13g2_inv_1 _26198_ (.Y(_18110_),
    .A(\u_inv.d_next[217] ));
 sg13g2_inv_1 _26199_ (.Y(_18111_),
    .A(\u_inv.d_next[215] ));
 sg13g2_inv_1 _26200_ (.Y(_18112_),
    .A(\u_inv.d_next[213] ));
 sg13g2_inv_1 _26201_ (.Y(_18113_),
    .A(\u_inv.d_next[210] ));
 sg13g2_inv_2 _26202_ (.Y(_18114_),
    .A(\u_inv.d_next[209] ));
 sg13g2_inv_1 _26203_ (.Y(_18115_),
    .A(\u_inv.d_next[207] ));
 sg13g2_inv_1 _26204_ (.Y(_18116_),
    .A(\u_inv.d_next[203] ));
 sg13g2_inv_1 _26205_ (.Y(_18117_),
    .A(net3374));
 sg13g2_inv_1 _26206_ (.Y(_18118_),
    .A(\u_inv.d_next[183] ));
 sg13g2_inv_1 _26207_ (.Y(_18119_),
    .A(net1982));
 sg13g2_inv_1 _26208_ (.Y(_18120_),
    .A(net2240));
 sg13g2_inv_1 _26209_ (.Y(_18121_),
    .A(\u_inv.d_next[177] ));
 sg13g2_inv_1 _26210_ (.Y(_18122_),
    .A(net2578));
 sg13g2_inv_1 _26211_ (.Y(_18123_),
    .A(\u_inv.d_next[168] ));
 sg13g2_inv_2 _26212_ (.Y(_18124_),
    .A(net1539));
 sg13g2_inv_1 _26213_ (.Y(_18125_),
    .A(net1496));
 sg13g2_inv_1 _26214_ (.Y(_18126_),
    .A(\u_inv.d_next[159] ));
 sg13g2_inv_1 _26215_ (.Y(_18127_),
    .A(\u_inv.d_next[151] ));
 sg13g2_inv_1 _26216_ (.Y(_18128_),
    .A(\u_inv.d_next[150] ));
 sg13g2_inv_1 _26217_ (.Y(_18129_),
    .A(net1902));
 sg13g2_inv_1 _26218_ (.Y(_18130_),
    .A(\u_inv.d_next[143] ));
 sg13g2_inv_1 _26219_ (.Y(_18131_),
    .A(\u_inv.d_next[141] ));
 sg13g2_inv_1 _26220_ (.Y(_18132_),
    .A(\u_inv.d_next[137] ));
 sg13g2_inv_1 _26221_ (.Y(_18133_),
    .A(net3475));
 sg13g2_inv_1 _26222_ (.Y(_18134_),
    .A(\u_inv.d_next[133] ));
 sg13g2_inv_1 _26223_ (.Y(_18135_),
    .A(\u_inv.d_next[131] ));
 sg13g2_inv_1 _26224_ (.Y(_18136_),
    .A(net2587));
 sg13g2_inv_1 _26225_ (.Y(_18137_),
    .A(\u_inv.d_next[125] ));
 sg13g2_inv_1 _26226_ (.Y(_18138_),
    .A(net2397));
 sg13g2_inv_1 _26227_ (.Y(_18139_),
    .A(\u_inv.d_next[119] ));
 sg13g2_inv_1 _26228_ (.Y(_18140_),
    .A(net2328));
 sg13g2_inv_1 _26229_ (.Y(_18141_),
    .A(\u_inv.d_next[111] ));
 sg13g2_inv_1 _26230_ (.Y(_18142_),
    .A(net2665));
 sg13g2_inv_1 _26231_ (.Y(_18143_),
    .A(net2869));
 sg13g2_inv_1 _26232_ (.Y(_18144_),
    .A(net2663));
 sg13g2_inv_1 _26233_ (.Y(_18145_),
    .A(\u_inv.d_next[105] ));
 sg13g2_inv_1 _26234_ (.Y(_18146_),
    .A(net2862));
 sg13g2_inv_1 _26235_ (.Y(_18147_),
    .A(\u_inv.d_next[95] ));
 sg13g2_inv_1 _26236_ (.Y(_18148_),
    .A(\u_inv.d_next[93] ));
 sg13g2_inv_1 _26237_ (.Y(_18149_),
    .A(\u_inv.d_next[89] ));
 sg13g2_inv_1 _26238_ (.Y(_18150_),
    .A(\u_inv.d_next[85] ));
 sg13g2_inv_1 _26239_ (.Y(_18151_),
    .A(\u_inv.d_next[83] ));
 sg13g2_inv_1 _26240_ (.Y(_18152_),
    .A(net3659));
 sg13g2_inv_1 _26241_ (.Y(_18153_),
    .A(net2366));
 sg13g2_inv_1 _26242_ (.Y(_18154_),
    .A(net1849));
 sg13g2_inv_1 _26243_ (.Y(_18155_),
    .A(net2585));
 sg13g2_inv_1 _26244_ (.Y(_18156_),
    .A(\u_inv.d_next[75] ));
 sg13g2_inv_1 _26245_ (.Y(_18157_),
    .A(net3523));
 sg13g2_inv_1 _26246_ (.Y(_18158_),
    .A(\u_inv.d_next[67] ));
 sg13g2_inv_1 _26247_ (.Y(_18159_),
    .A(net2521));
 sg13g2_inv_1 _26248_ (.Y(_18160_),
    .A(net3009));
 sg13g2_inv_1 _26249_ (.Y(_18161_),
    .A(\u_inv.d_next[61] ));
 sg13g2_inv_1 _26250_ (.Y(_18162_),
    .A(\u_inv.d_next[55] ));
 sg13g2_inv_1 _26251_ (.Y(_18163_),
    .A(net2910));
 sg13g2_inv_1 _26252_ (.Y(_18164_),
    .A(\u_inv.d_next[49] ));
 sg13g2_inv_1 _26253_ (.Y(_18165_),
    .A(\u_inv.d_next[47] ));
 sg13g2_inv_1 _26254_ (.Y(_18166_),
    .A(net3353));
 sg13g2_inv_1 _26255_ (.Y(_18167_),
    .A(net3124));
 sg13g2_inv_1 _26256_ (.Y(_18168_),
    .A(\u_inv.d_next[43] ));
 sg13g2_inv_1 _26257_ (.Y(_18169_),
    .A(net1724));
 sg13g2_inv_1 _26258_ (.Y(_18170_),
    .A(net2762));
 sg13g2_inv_1 _26259_ (.Y(_18171_),
    .A(net2705));
 sg13g2_inv_1 _26260_ (.Y(_18172_),
    .A(net1955));
 sg13g2_inv_1 _26261_ (.Y(_18173_),
    .A(\u_inv.d_next[33] ));
 sg13g2_inv_1 _26262_ (.Y(_18174_),
    .A(net1742));
 sg13g2_inv_1 _26263_ (.Y(_18175_),
    .A(\u_inv.d_next[29] ));
 sg13g2_inv_1 _26264_ (.Y(_18176_),
    .A(net2268));
 sg13g2_inv_1 _26265_ (.Y(_18177_),
    .A(net2038));
 sg13g2_inv_1 _26266_ (.Y(_18178_),
    .A(\u_inv.d_next[19] ));
 sg13g2_inv_1 _26267_ (.Y(_18179_),
    .A(net2945));
 sg13g2_inv_1 _26268_ (.Y(_18180_),
    .A(\u_inv.d_next[9] ));
 sg13g2_inv_1 _26269_ (.Y(_18181_),
    .A(inv_go));
 sg13g2_inv_1 _26270_ (.Y(_18182_),
    .A(\u_inv.input_valid ));
 sg13g2_inv_1 _26271_ (.Y(_18183_),
    .A(\u_inv.f_reg[0] ));
 sg13g2_inv_2 _26272_ (.Y(_18184_),
    .A(net3602));
 sg13g2_inv_1 _26273_ (.Y(_18185_),
    .A(\u_inv.delta_reg[3] ));
 sg13g2_inv_1 _26274_ (.Y(_18186_),
    .A(\u_inv.delta_reg[6] ));
 sg13g2_inv_1 _26275_ (.Y(_18187_),
    .A(\u_inv.delta_reg[8] ));
 sg13g2_inv_2 _26276_ (.Y(_18188_),
    .A(net3639));
 sg13g2_inv_4 _26277_ (.A(net3636),
    .Y(_18189_));
 sg13g2_inv_2 _26278_ (.Y(_18190_),
    .A(\u_inv.counter[3] ));
 sg13g2_inv_1 _26279_ (.Y(_18191_),
    .A(\u_inv.f_reg[4] ));
 sg13g2_inv_1 _26280_ (.Y(_18192_),
    .A(net1636));
 sg13g2_inv_1 _26281_ (.Y(_18193_),
    .A(\u_inv.f_reg[7] ));
 sg13g2_inv_1 _26282_ (.Y(_18194_),
    .A(net1549));
 sg13g2_inv_2 _26283_ (.Y(_18195_),
    .A(net2628));
 sg13g2_inv_1 _26284_ (.Y(_18196_),
    .A(\u_inv.f_reg[20] ));
 sg13g2_inv_1 _26285_ (.Y(_18197_),
    .A(\u_inv.f_reg[21] ));
 sg13g2_inv_1 _26286_ (.Y(_18198_),
    .A(\u_inv.f_reg[22] ));
 sg13g2_inv_1 _26287_ (.Y(_18199_),
    .A(\u_inv.f_reg[30] ));
 sg13g2_inv_1 _26288_ (.Y(_18200_),
    .A(\u_inv.f_reg[32] ));
 sg13g2_inv_1 _26289_ (.Y(_18201_),
    .A(\u_inv.f_reg[33] ));
 sg13g2_inv_1 _26290_ (.Y(_18202_),
    .A(\u_inv.f_reg[39] ));
 sg13g2_inv_1 _26291_ (.Y(_18203_),
    .A(\u_inv.f_reg[47] ));
 sg13g2_inv_1 _26292_ (.Y(_18204_),
    .A(\u_inv.f_reg[54] ));
 sg13g2_inv_1 _26293_ (.Y(_18205_),
    .A(\u_inv.f_reg[55] ));
 sg13g2_inv_1 _26294_ (.Y(_18206_),
    .A(\u_inv.f_reg[59] ));
 sg13g2_inv_1 _26295_ (.Y(_18207_),
    .A(\u_inv.f_reg[63] ));
 sg13g2_inv_1 _26296_ (.Y(_18208_),
    .A(\u_inv.f_reg[69] ));
 sg13g2_inv_1 _26297_ (.Y(_18209_),
    .A(\u_inv.f_reg[73] ));
 sg13g2_inv_1 _26298_ (.Y(_18210_),
    .A(\u_inv.f_reg[77] ));
 sg13g2_inv_1 _26299_ (.Y(_18211_),
    .A(\u_inv.f_reg[81] ));
 sg13g2_inv_1 _26300_ (.Y(_18212_),
    .A(\u_inv.f_reg[88] ));
 sg13g2_inv_1 _26301_ (.Y(_18213_),
    .A(\u_inv.f_reg[91] ));
 sg13g2_inv_1 _26302_ (.Y(_18214_),
    .A(\u_inv.f_reg[93] ));
 sg13g2_inv_1 _26303_ (.Y(_18215_),
    .A(\u_inv.f_reg[97] ));
 sg13g2_inv_1 _26304_ (.Y(_18216_),
    .A(\u_inv.f_reg[105] ));
 sg13g2_inv_1 _26305_ (.Y(_18217_),
    .A(\u_inv.f_reg[107] ));
 sg13g2_inv_1 _26306_ (.Y(_18218_),
    .A(\u_inv.f_reg[111] ));
 sg13g2_inv_1 _26307_ (.Y(_18219_),
    .A(\u_inv.f_reg[117] ));
 sg13g2_inv_1 _26308_ (.Y(_18220_),
    .A(\u_inv.f_reg[119] ));
 sg13g2_inv_1 _26309_ (.Y(_18221_),
    .A(\u_inv.f_reg[121] ));
 sg13g2_inv_1 _26310_ (.Y(_18222_),
    .A(\u_inv.f_reg[123] ));
 sg13g2_inv_1 _26311_ (.Y(_18223_),
    .A(\u_inv.f_reg[125] ));
 sg13g2_inv_1 _26312_ (.Y(_18224_),
    .A(\u_inv.f_reg[139] ));
 sg13g2_inv_1 _26313_ (.Y(_18225_),
    .A(\u_inv.f_reg[141] ));
 sg13g2_inv_1 _26314_ (.Y(_18226_),
    .A(\u_inv.f_reg[142] ));
 sg13g2_inv_1 _26315_ (.Y(_18227_),
    .A(\u_inv.f_reg[147] ));
 sg13g2_inv_1 _26316_ (.Y(_18228_),
    .A(\u_inv.f_reg[149] ));
 sg13g2_inv_1 _26317_ (.Y(_18229_),
    .A(\u_inv.f_reg[155] ));
 sg13g2_inv_1 _26318_ (.Y(_18230_),
    .A(\u_inv.f_reg[161] ));
 sg13g2_inv_1 _26319_ (.Y(_18231_),
    .A(\u_inv.f_reg[163] ));
 sg13g2_inv_1 _26320_ (.Y(_18232_),
    .A(\u_inv.f_reg[167] ));
 sg13g2_inv_1 _26321_ (.Y(_18233_),
    .A(\u_inv.f_reg[171] ));
 sg13g2_inv_1 _26322_ (.Y(_18234_),
    .A(\u_inv.f_reg[173] ));
 sg13g2_inv_1 _26323_ (.Y(_18235_),
    .A(\u_inv.f_reg[175] ));
 sg13g2_inv_1 _26324_ (.Y(_18236_),
    .A(\u_inv.f_reg[177] ));
 sg13g2_inv_1 _26325_ (.Y(_18237_),
    .A(\u_inv.f_reg[179] ));
 sg13g2_inv_1 _26326_ (.Y(_18238_),
    .A(\u_inv.f_reg[183] ));
 sg13g2_inv_1 _26327_ (.Y(_18239_),
    .A(\u_inv.f_reg[185] ));
 sg13g2_inv_1 _26328_ (.Y(_18240_),
    .A(\u_inv.f_reg[187] ));
 sg13g2_inv_1 _26329_ (.Y(_18241_),
    .A(\u_inv.f_reg[191] ));
 sg13g2_inv_1 _26330_ (.Y(_18242_),
    .A(\u_inv.f_reg[192] ));
 sg13g2_inv_1 _26331_ (.Y(_18243_),
    .A(\u_inv.f_reg[195] ));
 sg13g2_inv_1 _26332_ (.Y(_18244_),
    .A(\u_inv.f_reg[196] ));
 sg13g2_inv_1 _26333_ (.Y(_18245_),
    .A(\u_inv.f_reg[201] ));
 sg13g2_inv_1 _26334_ (.Y(_18246_),
    .A(\u_inv.f_reg[205] ));
 sg13g2_inv_1 _26335_ (.Y(_18247_),
    .A(\u_inv.f_reg[207] ));
 sg13g2_inv_1 _26336_ (.Y(_18248_),
    .A(\u_inv.f_reg[213] ));
 sg13g2_inv_1 _26337_ (.Y(_18249_),
    .A(\u_inv.f_reg[219] ));
 sg13g2_inv_1 _26338_ (.Y(_18250_),
    .A(\u_inv.f_reg[225] ));
 sg13g2_inv_1 _26339_ (.Y(_18251_),
    .A(\u_inv.f_reg[229] ));
 sg13g2_inv_1 _26340_ (.Y(_18252_),
    .A(\u_inv.f_reg[235] ));
 sg13g2_inv_1 _26341_ (.Y(_18253_),
    .A(\u_inv.f_reg[251] ));
 sg13g2_inv_1 _26342_ (.Y(_18254_),
    .A(net7269));
 sg13g2_inv_2 _26343_ (.Y(_18255_),
    .A(net7250));
 sg13g2_inv_1 _26344_ (.Y(_18256_),
    .A(net1166));
 sg13g2_inv_1 _26345_ (.Y(_18257_),
    .A(net13));
 sg13g2_inv_1 _26346_ (.Y(_18258_),
    .A(net1730));
 sg13g2_inv_1 _26347_ (.Y(_18259_),
    .A(net1969));
 sg13g2_inv_1 _26348_ (.Y(_18260_),
    .A(net1521));
 sg13g2_inv_1 _26349_ (.Y(_18261_),
    .A(net1574));
 sg13g2_inv_1 _26350_ (.Y(_18262_),
    .A(net3402));
 sg13g2_inv_1 _26351_ (.Y(_18263_),
    .A(net3671));
 sg13g2_inv_1 _26352_ (.Y(_18264_),
    .A(net3450));
 sg13g2_inv_1 _26353_ (.Y(_18265_),
    .A(parity_error));
 sg13g2_inv_1 _26354_ (.Y(_18266_),
    .A(net1192));
 sg13g2_inv_1 _26355_ (.Y(_18267_),
    .A(net2179));
 sg13g2_inv_1 _26356_ (.Y(_18268_),
    .A(net2336));
 sg13g2_inv_1 _26357_ (.Y(_18269_),
    .A(net1488));
 sg13g2_inv_1 _26358_ (.Y(_18270_),
    .A(net2469));
 sg13g2_inv_1 _26359_ (.Y(_18271_),
    .A(net1548));
 sg13g2_inv_1 _26360_ (.Y(_18272_),
    .A(net1298));
 sg13g2_inv_1 _26361_ (.Y(_18273_),
    .A(net1220));
 sg13g2_inv_1 _26362_ (.Y(_18274_),
    .A(net1326));
 sg13g2_inv_1 _26363_ (.Y(_18275_),
    .A(net1245));
 sg13g2_inv_1 _26364_ (.Y(_18276_),
    .A(net1254));
 sg13g2_inv_1 _26365_ (.Y(_18277_),
    .A(net1403));
 sg13g2_inv_1 _26366_ (.Y(_18278_),
    .A(net1270));
 sg13g2_inv_1 _26367_ (.Y(_18279_),
    .A(net1273));
 sg13g2_inv_1 _26368_ (.Y(_18280_),
    .A(net1232));
 sg13g2_inv_1 _26369_ (.Y(_18281_),
    .A(net1230));
 sg13g2_inv_1 _26370_ (.Y(_18282_),
    .A(net1458));
 sg13g2_inv_1 _26371_ (.Y(_18283_),
    .A(net1297));
 sg13g2_inv_1 _26372_ (.Y(_18284_),
    .A(net1260));
 sg13g2_inv_1 _26373_ (.Y(_18285_),
    .A(net1227));
 sg13g2_inv_1 _26374_ (.Y(_18286_),
    .A(net1479));
 sg13g2_inv_1 _26375_ (.Y(_18287_),
    .A(net1261));
 sg13g2_inv_1 _26376_ (.Y(_18288_),
    .A(net1219));
 sg13g2_inv_1 _26377_ (.Y(_18289_),
    .A(net1292));
 sg13g2_inv_1 _26378_ (.Y(_18290_),
    .A(net2012));
 sg13g2_inv_1 _26379_ (.Y(_18291_),
    .A(net1710));
 sg13g2_inv_1 _26380_ (.Y(_18292_),
    .A(net1355));
 sg13g2_inv_1 _26381_ (.Y(_18293_),
    .A(net1228));
 sg13g2_inv_1 _26382_ (.Y(_18294_),
    .A(net1464));
 sg13g2_inv_1 _26383_ (.Y(_18295_),
    .A(net2343));
 sg13g2_inv_1 _26384_ (.Y(_18296_),
    .A(net1237));
 sg13g2_inv_1 _26385_ (.Y(_18297_),
    .A(net1919));
 sg13g2_inv_1 _26386_ (.Y(_18298_),
    .A(net1248));
 sg13g2_inv_1 _26387_ (.Y(_18299_),
    .A(\inv_result[214] ));
 sg13g2_inv_1 _26388_ (.Y(_18300_),
    .A(net1543));
 sg13g2_inv_1 _26389_ (.Y(_18301_),
    .A(net1246));
 sg13g2_inv_1 _26390_ (.Y(_18302_),
    .A(net1899));
 sg13g2_inv_1 _26391_ (.Y(_18303_),
    .A(\inv_result[221] ));
 sg13g2_inv_1 _26392_ (.Y(_18304_),
    .A(net2029));
 sg13g2_inv_1 _26393_ (.Y(_18305_),
    .A(net1663));
 sg13g2_inv_1 _26394_ (.Y(_18306_),
    .A(net1606));
 sg13g2_inv_1 _26395_ (.Y(_18307_),
    .A(\inv_result[225] ));
 sg13g2_inv_1 _26396_ (.Y(_18308_),
    .A(net1231));
 sg13g2_inv_1 _26397_ (.Y(_18309_),
    .A(net1664));
 sg13g2_inv_1 _26398_ (.Y(_18310_),
    .A(net1226));
 sg13g2_inv_1 _26399_ (.Y(_18311_),
    .A(net1182));
 sg13g2_inv_1 _26400_ (.Y(_18312_),
    .A(net1518));
 sg13g2_inv_1 _26401_ (.Y(_18313_),
    .A(net1301));
 sg13g2_inv_1 _26402_ (.Y(_18314_),
    .A(net1384));
 sg13g2_inv_1 _26403_ (.Y(_18315_),
    .A(net2530));
 sg13g2_inv_1 _26404_ (.Y(_18316_),
    .A(net2148));
 sg13g2_inv_1 _26405_ (.Y(_18317_),
    .A(net2276));
 sg13g2_inv_1 _26406_ (.Y(_18318_),
    .A(net1933));
 sg13g2_inv_1 _26407_ (.Y(_18319_),
    .A(net1278));
 sg13g2_inv_1 _26408_ (.Y(_18320_),
    .A(net1880));
 sg13g2_inv_1 _26409_ (.Y(_18321_),
    .A(net3186));
 sg13g2_inv_1 _26410_ (.Y(_18322_),
    .A(net2259));
 sg13g2_inv_1 _26411_ (.Y(_18323_),
    .A(\inv_result[247] ));
 sg13g2_inv_1 _26412_ (.Y(_18324_),
    .A(net2098));
 sg13g2_inv_1 _26413_ (.Y(_18325_),
    .A(net2002));
 sg13g2_inv_1 _26414_ (.Y(_18326_),
    .A(net2723));
 sg13g2_inv_1 _26415_ (.Y(_18327_),
    .A(net3371));
 sg13g2_inv_1 _26416_ (.Y(_18328_),
    .A(net1644));
 sg13g2_inv_2 _26417_ (.Y(_18329_),
    .A(net3304));
 sg13g2_inv_1 _26418_ (.Y(_18330_),
    .A(net1965));
 sg13g2_inv_1 _26419_ (.Y(_18331_),
    .A(net1508));
 sg13g2_inv_1 _26420_ (.Y(_18332_),
    .A(net2193));
 sg13g2_inv_1 _26421_ (.Y(_18333_),
    .A(net1494));
 sg13g2_inv_1 _26422_ (.Y(_18334_),
    .A(net1324));
 sg13g2_inv_1 _26423_ (.Y(_18335_),
    .A(net2658));
 sg13g2_inv_1 _26424_ (.Y(_18336_),
    .A(net1814));
 sg13g2_inv_1 _26425_ (.Y(_18337_),
    .A(net2466));
 sg13g2_inv_1 _26426_ (.Y(_18338_),
    .A(net1199));
 sg13g2_inv_1 _26427_ (.Y(_18339_),
    .A(net1212));
 sg13g2_inv_1 _26428_ (.Y(_18340_),
    .A(net1221));
 sg13g2_inv_1 _26429_ (.Y(_18341_),
    .A(\perf_triple[3] ));
 sg13g2_inv_1 _26430_ (.Y(_18342_),
    .A(net2672));
 sg13g2_inv_1 _26431_ (.Y(_18343_),
    .A(net3284));
 sg13g2_inv_1 _26432_ (.Y(_18344_),
    .A(net2592));
 sg13g2_inv_1 _26433_ (.Y(_18345_),
    .A(net1216));
 sg13g2_inv_1 _26434_ (.Y(_18346_),
    .A(net1387));
 sg13g2_inv_2 _26435_ (.Y(_18347_),
    .A(net1164));
 sg13g2_inv_1 _26436_ (.Y(_18348_),
    .A(net1251));
 sg13g2_inv_2 _26437_ (.Y(_18349_),
    .A(net1169));
 sg13g2_inv_1 _26438_ (.Y(_18350_),
    .A(net1149));
 sg13g2_inv_1 _26439_ (.Y(_18351_),
    .A(net1266));
 sg13g2_inv_1 _26440_ (.Y(_18352_),
    .A(net1155));
 sg13g2_inv_1 _26441_ (.Y(_18353_),
    .A(net1279));
 sg13g2_inv_1 _26442_ (.Y(_18354_),
    .A(net2069));
 sg13g2_inv_1 _26443_ (.Y(_18355_),
    .A(\perf_total[9] ));
 sg13g2_inv_1 _26444_ (.Y(_18356_),
    .A(net1151));
 sg13g2_inv_2 _26445_ (.Y(_18357_),
    .A(net7294));
 sg13g2_inv_2 _26446_ (.Y(_18358_),
    .A(net3388));
 sg13g2_inv_1 _26447_ (.Y(_18359_),
    .A(\u_inv.d_reg[255] ));
 sg13g2_inv_2 _26448_ (.Y(_18360_),
    .A(\u_inv.d_reg[254] ));
 sg13g2_inv_2 _26449_ (.Y(_18361_),
    .A(net3525));
 sg13g2_inv_2 _26450_ (.Y(_18362_),
    .A(net3574));
 sg13g2_inv_2 _26451_ (.Y(_18363_),
    .A(net3064));
 sg13g2_inv_1 _26452_ (.Y(_18364_),
    .A(net2894));
 sg13g2_inv_2 _26453_ (.Y(_18365_),
    .A(\u_inv.d_reg[249] ));
 sg13g2_inv_2 _26454_ (.Y(_18366_),
    .A(\u_inv.d_reg[248] ));
 sg13g2_inv_2 _26455_ (.Y(_18367_),
    .A(\u_inv.d_reg[247] ));
 sg13g2_inv_2 _26456_ (.Y(_18368_),
    .A(net3044));
 sg13g2_inv_2 _26457_ (.Y(_18369_),
    .A(net3675));
 sg13g2_inv_2 _26458_ (.Y(_18370_),
    .A(net3138));
 sg13g2_inv_1 _26459_ (.Y(_18371_),
    .A(\u_inv.d_reg[243] ));
 sg13g2_inv_1 _26460_ (.Y(_18372_),
    .A(net3611));
 sg13g2_inv_1 _26461_ (.Y(_18373_),
    .A(net7287));
 sg13g2_inv_1 _26462_ (.Y(_18374_),
    .A(net7288));
 sg13g2_inv_1 _26463_ (.Y(_18375_),
    .A(net3025));
 sg13g2_inv_1 _26464_ (.Y(_18376_),
    .A(net3201));
 sg13g2_inv_1 _26465_ (.Y(_18377_),
    .A(\u_inv.d_reg[237] ));
 sg13g2_inv_1 _26466_ (.Y(_18378_),
    .A(net3404));
 sg13g2_inv_1 _26467_ (.Y(_18379_),
    .A(\u_inv.d_reg[235] ));
 sg13g2_inv_1 _26468_ (.Y(_18380_),
    .A(net2963));
 sg13g2_inv_2 _26469_ (.Y(_18381_),
    .A(\u_inv.d_reg[233] ));
 sg13g2_inv_2 _26470_ (.Y(_18382_),
    .A(net3309));
 sg13g2_inv_1 _26471_ (.Y(_18383_),
    .A(\u_inv.d_reg[231] ));
 sg13g2_inv_1 _26472_ (.Y(_18384_),
    .A(net3483));
 sg13g2_inv_1 _26473_ (.Y(_18385_),
    .A(\u_inv.d_reg[229] ));
 sg13g2_inv_2 _26474_ (.Y(_18386_),
    .A(net3542));
 sg13g2_inv_4 _26475_ (.A(\u_inv.d_reg[227] ),
    .Y(_18387_));
 sg13g2_inv_2 _26476_ (.Y(_18388_),
    .A(net3291));
 sg13g2_inv_2 _26477_ (.Y(_18389_),
    .A(net2745));
 sg13g2_inv_1 _26478_ (.Y(_18390_),
    .A(\u_inv.d_reg[224] ));
 sg13g2_inv_2 _26479_ (.Y(_18391_),
    .A(\u_inv.d_reg[223] ));
 sg13g2_inv_2 _26480_ (.Y(_18392_),
    .A(\u_inv.d_reg[222] ));
 sg13g2_inv_1 _26481_ (.Y(_18393_),
    .A(\u_inv.d_reg[221] ));
 sg13g2_inv_1 _26482_ (.Y(_18394_),
    .A(\u_inv.d_reg[220] ));
 sg13g2_inv_2 _26483_ (.Y(_18395_),
    .A(\u_inv.d_reg[219] ));
 sg13g2_inv_1 _26484_ (.Y(_18396_),
    .A(\u_inv.d_reg[218] ));
 sg13g2_inv_1 _26485_ (.Y(_18397_),
    .A(\u_inv.d_reg[217] ));
 sg13g2_inv_2 _26486_ (.Y(_18398_),
    .A(\u_inv.d_reg[216] ));
 sg13g2_inv_2 _26487_ (.Y(_18399_),
    .A(\u_inv.d_reg[215] ));
 sg13g2_inv_1 _26488_ (.Y(_18400_),
    .A(\u_inv.d_reg[214] ));
 sg13g2_inv_2 _26489_ (.Y(_18401_),
    .A(\u_inv.d_reg[213] ));
 sg13g2_inv_2 _26490_ (.Y(_18402_),
    .A(\u_inv.d_reg[212] ));
 sg13g2_inv_2 _26491_ (.Y(_18403_),
    .A(\u_inv.d_reg[211] ));
 sg13g2_inv_2 _26492_ (.Y(_18404_),
    .A(\u_inv.d_reg[210] ));
 sg13g2_inv_2 _26493_ (.Y(_18405_),
    .A(\u_inv.d_reg[209] ));
 sg13g2_inv_2 _26494_ (.Y(_18406_),
    .A(\u_inv.d_reg[208] ));
 sg13g2_inv_1 _26495_ (.Y(_18407_),
    .A(\u_inv.d_reg[207] ));
 sg13g2_inv_2 _26496_ (.Y(_18408_),
    .A(net3038));
 sg13g2_inv_2 _26497_ (.Y(_18409_),
    .A(\u_inv.d_reg[205] ));
 sg13g2_inv_2 _26498_ (.Y(_18410_),
    .A(net2833));
 sg13g2_inv_1 _26499_ (.Y(_18411_),
    .A(\u_inv.d_reg[203] ));
 sg13g2_inv_1 _26500_ (.Y(_18412_),
    .A(net3144));
 sg13g2_inv_2 _26501_ (.Y(_18413_),
    .A(\u_inv.d_reg[201] ));
 sg13g2_inv_2 _26502_ (.Y(_18414_),
    .A(\u_inv.d_reg[200] ));
 sg13g2_inv_2 _26503_ (.Y(_18415_),
    .A(\u_inv.d_reg[199] ));
 sg13g2_inv_2 _26504_ (.Y(_18416_),
    .A(net3213));
 sg13g2_inv_1 _26505_ (.Y(_18417_),
    .A(net3590));
 sg13g2_inv_2 _26506_ (.Y(_18418_),
    .A(\u_inv.d_reg[196] ));
 sg13g2_inv_1 _26507_ (.Y(_18419_),
    .A(\u_inv.d_reg[195] ));
 sg13g2_inv_1 _26508_ (.Y(_18420_),
    .A(\u_inv.d_reg[194] ));
 sg13g2_inv_1 _26509_ (.Y(_18421_),
    .A(net3610));
 sg13g2_inv_2 _26510_ (.Y(_18422_),
    .A(\u_inv.d_reg[192] ));
 sg13g2_inv_2 _26511_ (.Y(_18423_),
    .A(\u_inv.d_reg[191] ));
 sg13g2_inv_1 _26512_ (.Y(_18424_),
    .A(net2834));
 sg13g2_inv_2 _26513_ (.Y(_18425_),
    .A(net3465));
 sg13g2_inv_1 _26514_ (.Y(_18426_),
    .A(net2932));
 sg13g2_inv_1 _26515_ (.Y(_18427_),
    .A(\u_inv.d_reg[187] ));
 sg13g2_inv_1 _26516_ (.Y(_18428_),
    .A(\u_inv.d_reg[186] ));
 sg13g2_inv_2 _26517_ (.Y(_18429_),
    .A(\u_inv.d_reg[185] ));
 sg13g2_inv_1 _26518_ (.Y(_18430_),
    .A(net2940));
 sg13g2_inv_1 _26519_ (.Y(_18431_),
    .A(\u_inv.d_reg[183] ));
 sg13g2_inv_1 _26520_ (.Y(_18432_),
    .A(net2142));
 sg13g2_inv_2 _26521_ (.Y(_18433_),
    .A(\u_inv.d_reg[181] ));
 sg13g2_inv_1 _26522_ (.Y(_18434_),
    .A(\u_inv.d_reg[180] ));
 sg13g2_inv_1 _26523_ (.Y(_18435_),
    .A(net2455));
 sg13g2_inv_1 _26524_ (.Y(_18436_),
    .A(\u_inv.d_reg[178] ));
 sg13g2_inv_2 _26525_ (.Y(_18437_),
    .A(\u_inv.d_reg[177] ));
 sg13g2_inv_2 _26526_ (.Y(_18438_),
    .A(\u_inv.d_reg[176] ));
 sg13g2_inv_2 _26527_ (.Y(_18439_),
    .A(\u_inv.d_reg[175] ));
 sg13g2_inv_1 _26528_ (.Y(_18440_),
    .A(net2837));
 sg13g2_inv_1 _26529_ (.Y(_18441_),
    .A(\u_inv.d_reg[173] ));
 sg13g2_inv_1 _26530_ (.Y(_18442_),
    .A(\u_inv.d_reg[172] ));
 sg13g2_inv_1 _26531_ (.Y(_18443_),
    .A(\u_inv.d_reg[171] ));
 sg13g2_inv_1 _26532_ (.Y(_18444_),
    .A(net2720));
 sg13g2_inv_1 _26533_ (.Y(_18445_),
    .A(\u_inv.d_reg[169] ));
 sg13g2_inv_2 _26534_ (.Y(_18446_),
    .A(\u_inv.d_reg[168] ));
 sg13g2_inv_2 _26535_ (.Y(_18447_),
    .A(\u_inv.d_reg[167] ));
 sg13g2_inv_1 _26536_ (.Y(_18448_),
    .A(net3533));
 sg13g2_inv_1 _26537_ (.Y(_18449_),
    .A(\u_inv.d_reg[165] ));
 sg13g2_inv_1 _26538_ (.Y(_18450_),
    .A(\u_inv.d_reg[164] ));
 sg13g2_inv_1 _26539_ (.Y(_18451_),
    .A(\u_inv.d_reg[163] ));
 sg13g2_inv_1 _26540_ (.Y(_18452_),
    .A(net3008));
 sg13g2_inv_2 _26541_ (.Y(_18453_),
    .A(\u_inv.d_reg[161] ));
 sg13g2_inv_1 _26542_ (.Y(_18454_),
    .A(\u_inv.d_reg[160] ));
 sg13g2_inv_2 _26543_ (.Y(_18455_),
    .A(\u_inv.d_reg[159] ));
 sg13g2_inv_2 _26544_ (.Y(_18456_),
    .A(\u_inv.d_reg[158] ));
 sg13g2_inv_1 _26545_ (.Y(_18457_),
    .A(\u_inv.d_reg[157] ));
 sg13g2_inv_1 _26546_ (.Y(_18458_),
    .A(\u_inv.d_reg[156] ));
 sg13g2_inv_2 _26547_ (.Y(_18459_),
    .A(\u_inv.d_reg[155] ));
 sg13g2_inv_2 _26548_ (.Y(_18460_),
    .A(\u_inv.d_reg[154] ));
 sg13g2_inv_1 _26549_ (.Y(_18461_),
    .A(net2613));
 sg13g2_inv_2 _26550_ (.Y(_18462_),
    .A(\u_inv.d_reg[152] ));
 sg13g2_inv_2 _26551_ (.Y(_18463_),
    .A(net3608));
 sg13g2_inv_1 _26552_ (.Y(_18464_),
    .A(net3422));
 sg13g2_inv_1 _26553_ (.Y(_18465_),
    .A(\u_inv.d_reg[149] ));
 sg13g2_inv_1 _26554_ (.Y(_18466_),
    .A(\u_inv.d_reg[148] ));
 sg13g2_inv_1 _26555_ (.Y(_18467_),
    .A(\u_inv.d_reg[147] ));
 sg13g2_inv_1 _26556_ (.Y(_18468_),
    .A(net3338));
 sg13g2_inv_2 _26557_ (.Y(_18469_),
    .A(\u_inv.d_reg[145] ));
 sg13g2_inv_2 _26558_ (.Y(_18470_),
    .A(\u_inv.d_reg[144] ));
 sg13g2_inv_1 _26559_ (.Y(_18471_),
    .A(\u_inv.d_reg[143] ));
 sg13g2_inv_2 _26560_ (.Y(_18472_),
    .A(net3618));
 sg13g2_inv_1 _26561_ (.Y(_18473_),
    .A(\u_inv.d_reg[141] ));
 sg13g2_inv_1 _26562_ (.Y(_18474_),
    .A(\u_inv.d_reg[140] ));
 sg13g2_inv_1 _26563_ (.Y(_18475_),
    .A(\u_inv.d_reg[139] ));
 sg13g2_inv_1 _26564_ (.Y(_18476_),
    .A(\u_inv.d_reg[138] ));
 sg13g2_inv_2 _26565_ (.Y(_18477_),
    .A(\u_inv.d_reg[137] ));
 sg13g2_inv_2 _26566_ (.Y(_18478_),
    .A(\u_inv.d_reg[136] ));
 sg13g2_inv_1 _26567_ (.Y(_18479_),
    .A(\u_inv.d_reg[135] ));
 sg13g2_inv_1 _26568_ (.Y(_18480_),
    .A(net3571));
 sg13g2_inv_2 _26569_ (.Y(_18481_),
    .A(\u_inv.d_reg[133] ));
 sg13g2_inv_1 _26570_ (.Y(_18482_),
    .A(\u_inv.d_reg[132] ));
 sg13g2_inv_2 _26571_ (.Y(_18483_),
    .A(\u_inv.d_reg[131] ));
 sg13g2_inv_1 _26572_ (.Y(_18484_),
    .A(\u_inv.d_reg[130] ));
 sg13g2_inv_2 _26573_ (.Y(_18485_),
    .A(\u_inv.d_reg[129] ));
 sg13g2_inv_1 _26574_ (.Y(_18486_),
    .A(\u_inv.d_reg[128] ));
 sg13g2_inv_1 _26575_ (.Y(_18487_),
    .A(net3616));
 sg13g2_inv_1 _26576_ (.Y(_18488_),
    .A(\u_inv.d_reg[126] ));
 sg13g2_inv_2 _26577_ (.Y(_18489_),
    .A(\u_inv.d_reg[125] ));
 sg13g2_inv_1 _26578_ (.Y(_18490_),
    .A(\u_inv.d_reg[124] ));
 sg13g2_inv_2 _26579_ (.Y(_18491_),
    .A(\u_inv.d_reg[123] ));
 sg13g2_inv_2 _26580_ (.Y(_18492_),
    .A(\u_inv.d_reg[122] ));
 sg13g2_inv_1 _26581_ (.Y(_18493_),
    .A(\u_inv.d_reg[121] ));
 sg13g2_inv_1 _26582_ (.Y(_18494_),
    .A(\u_inv.d_reg[120] ));
 sg13g2_inv_2 _26583_ (.Y(_18495_),
    .A(\u_inv.d_reg[119] ));
 sg13g2_inv_2 _26584_ (.Y(_18496_),
    .A(net2637));
 sg13g2_inv_2 _26585_ (.Y(_18497_),
    .A(\u_inv.d_reg[117] ));
 sg13g2_inv_2 _26586_ (.Y(_18498_),
    .A(\u_inv.d_reg[116] ));
 sg13g2_inv_1 _26587_ (.Y(_18499_),
    .A(\u_inv.d_reg[115] ));
 sg13g2_inv_1 _26588_ (.Y(_18500_),
    .A(net3264));
 sg13g2_inv_2 _26589_ (.Y(_18501_),
    .A(\u_inv.d_reg[113] ));
 sg13g2_inv_1 _26590_ (.Y(_18502_),
    .A(net3680));
 sg13g2_inv_2 _26591_ (.Y(_18503_),
    .A(net3604));
 sg13g2_inv_1 _26592_ (.Y(_18504_),
    .A(net2383));
 sg13g2_inv_2 _26593_ (.Y(_18505_),
    .A(\u_inv.d_reg[109] ));
 sg13g2_inv_2 _26594_ (.Y(_18506_),
    .A(\u_inv.d_reg[108] ));
 sg13g2_inv_8 _26595_ (.Y(_18507_),
    .A(\u_inv.d_reg[107] ));
 sg13g2_inv_4 _26596_ (.A(\u_inv.d_reg[106] ),
    .Y(_18508_));
 sg13g2_inv_2 _26597_ (.Y(_18509_),
    .A(\u_inv.d_reg[105] ));
 sg13g2_inv_2 _26598_ (.Y(_18510_),
    .A(\u_inv.d_reg[104] ));
 sg13g2_inv_1 _26599_ (.Y(_18511_),
    .A(\u_inv.d_reg[103] ));
 sg13g2_inv_2 _26600_ (.Y(_18512_),
    .A(net3255));
 sg13g2_inv_1 _26601_ (.Y(_18513_),
    .A(\u_inv.d_reg[101] ));
 sg13g2_inv_1 _26602_ (.Y(_18514_),
    .A(\u_inv.d_reg[100] ));
 sg13g2_inv_1 _26603_ (.Y(_18515_),
    .A(\u_inv.d_reg[99] ));
 sg13g2_inv_1 _26604_ (.Y(_18516_),
    .A(\u_inv.d_reg[98] ));
 sg13g2_inv_2 _26605_ (.Y(_18517_),
    .A(\u_inv.d_reg[97] ));
 sg13g2_inv_1 _26606_ (.Y(_18518_),
    .A(\u_inv.d_reg[96] ));
 sg13g2_inv_2 _26607_ (.Y(_18519_),
    .A(net3640));
 sg13g2_inv_2 _26608_ (.Y(_18520_),
    .A(\u_inv.d_reg[94] ));
 sg13g2_inv_1 _26609_ (.Y(_18521_),
    .A(\u_inv.d_reg[93] ));
 sg13g2_inv_1 _26610_ (.Y(_18522_),
    .A(\u_inv.d_reg[92] ));
 sg13g2_inv_1 _26611_ (.Y(_18523_),
    .A(\u_inv.d_reg[91] ));
 sg13g2_inv_1 _26612_ (.Y(_18524_),
    .A(net3280));
 sg13g2_inv_2 _26613_ (.Y(_18525_),
    .A(\u_inv.d_reg[89] ));
 sg13g2_inv_1 _26614_ (.Y(_18526_),
    .A(\u_inv.d_reg[88] ));
 sg13g2_inv_1 _26615_ (.Y(_18527_),
    .A(\u_inv.d_reg[87] ));
 sg13g2_inv_1 _26616_ (.Y(_18528_),
    .A(\u_inv.d_reg[86] ));
 sg13g2_inv_2 _26617_ (.Y(_18529_),
    .A(net2895));
 sg13g2_inv_2 _26618_ (.Y(_18530_),
    .A(\u_inv.d_reg[84] ));
 sg13g2_inv_1 _26619_ (.Y(_18531_),
    .A(\u_inv.d_reg[83] ));
 sg13g2_inv_1 _26620_ (.Y(_18532_),
    .A(\u_inv.d_reg[82] ));
 sg13g2_inv_2 _26621_ (.Y(_18533_),
    .A(net2731));
 sg13g2_inv_2 _26622_ (.Y(_18534_),
    .A(\u_inv.d_reg[80] ));
 sg13g2_inv_1 _26623_ (.Y(_18535_),
    .A(\u_inv.d_reg[79] ));
 sg13g2_inv_1 _26624_ (.Y(_18536_),
    .A(\u_inv.d_reg[78] ));
 sg13g2_inv_2 _26625_ (.Y(_18537_),
    .A(\u_inv.d_reg[77] ));
 sg13g2_inv_2 _26626_ (.Y(_18538_),
    .A(\u_inv.d_reg[76] ));
 sg13g2_inv_2 _26627_ (.Y(_18539_),
    .A(\u_inv.d_reg[75] ));
 sg13g2_inv_2 _26628_ (.Y(_18540_),
    .A(\u_inv.d_reg[74] ));
 sg13g2_inv_2 _26629_ (.Y(_18541_),
    .A(net3515));
 sg13g2_inv_2 _26630_ (.Y(_18542_),
    .A(\u_inv.d_reg[72] ));
 sg13g2_inv_1 _26631_ (.Y(_18543_),
    .A(net3480));
 sg13g2_inv_2 _26632_ (.Y(_18544_),
    .A(net3673));
 sg13g2_inv_1 _26633_ (.Y(_18545_),
    .A(\u_inv.d_reg[69] ));
 sg13g2_inv_2 _26634_ (.Y(_18546_),
    .A(\u_inv.d_reg[68] ));
 sg13g2_inv_1 _26635_ (.Y(_18547_),
    .A(\u_inv.d_reg[67] ));
 sg13g2_inv_1 _26636_ (.Y(_18548_),
    .A(\u_inv.d_reg[66] ));
 sg13g2_inv_1 _26637_ (.Y(_18549_),
    .A(\u_inv.d_reg[65] ));
 sg13g2_inv_1 _26638_ (.Y(_18550_),
    .A(\u_inv.d_reg[64] ));
 sg13g2_inv_1 _26639_ (.Y(_18551_),
    .A(\u_inv.d_reg[63] ));
 sg13g2_inv_1 _26640_ (.Y(_18552_),
    .A(net3287));
 sg13g2_inv_1 _26641_ (.Y(_18553_),
    .A(\u_inv.d_reg[61] ));
 sg13g2_inv_2 _26642_ (.Y(_18554_),
    .A(\u_inv.d_reg[60] ));
 sg13g2_inv_2 _26643_ (.Y(_18555_),
    .A(net3258));
 sg13g2_inv_2 _26644_ (.Y(_18556_),
    .A(\u_inv.d_reg[58] ));
 sg13g2_inv_1 _26645_ (.Y(_18557_),
    .A(net2443));
 sg13g2_inv_2 _26646_ (.Y(_18558_),
    .A(\u_inv.d_reg[56] ));
 sg13g2_inv_1 _26647_ (.Y(_18559_),
    .A(net2775));
 sg13g2_inv_2 _26648_ (.Y(_18560_),
    .A(\u_inv.d_reg[54] ));
 sg13g2_inv_1 _26649_ (.Y(_18561_),
    .A(\u_inv.d_reg[53] ));
 sg13g2_inv_2 _26650_ (.Y(_18562_),
    .A(net3536));
 sg13g2_inv_2 _26651_ (.Y(_18563_),
    .A(\u_inv.d_reg[51] ));
 sg13g2_inv_2 _26652_ (.Y(_18564_),
    .A(\u_inv.d_reg[50] ));
 sg13g2_inv_2 _26653_ (.Y(_18565_),
    .A(net3179));
 sg13g2_inv_2 _26654_ (.Y(_18566_),
    .A(\u_inv.d_reg[48] ));
 sg13g2_inv_1 _26655_ (.Y(_18567_),
    .A(\u_inv.d_reg[47] ));
 sg13g2_inv_1 _26656_ (.Y(_18568_),
    .A(net2971));
 sg13g2_inv_2 _26657_ (.Y(_18569_),
    .A(\u_inv.d_reg[45] ));
 sg13g2_inv_1 _26658_ (.Y(_18570_),
    .A(\u_inv.d_reg[44] ));
 sg13g2_inv_2 _26659_ (.Y(_18571_),
    .A(\u_inv.d_reg[43] ));
 sg13g2_inv_2 _26660_ (.Y(_18572_),
    .A(\u_inv.d_reg[42] ));
 sg13g2_inv_1 _26661_ (.Y(_18573_),
    .A(\u_inv.d_reg[41] ));
 sg13g2_inv_1 _26662_ (.Y(_18574_),
    .A(\u_inv.d_reg[40] ));
 sg13g2_inv_1 _26663_ (.Y(_18575_),
    .A(\u_inv.d_reg[39] ));
 sg13g2_inv_2 _26664_ (.Y(_18576_),
    .A(\u_inv.d_reg[38] ));
 sg13g2_inv_2 _26665_ (.Y(_18577_),
    .A(\u_inv.d_reg[37] ));
 sg13g2_inv_2 _26666_ (.Y(_18578_),
    .A(\u_inv.d_reg[36] ));
 sg13g2_inv_2 _26667_ (.Y(_18579_),
    .A(\u_inv.d_reg[35] ));
 sg13g2_inv_2 _26668_ (.Y(_18580_),
    .A(\u_inv.d_reg[34] ));
 sg13g2_inv_2 _26669_ (.Y(_18581_),
    .A(\u_inv.d_reg[33] ));
 sg13g2_inv_1 _26670_ (.Y(_18582_),
    .A(\u_inv.d_reg[32] ));
 sg13g2_inv_2 _26671_ (.Y(_18583_),
    .A(\u_inv.d_reg[31] ));
 sg13g2_inv_1 _26672_ (.Y(_18584_),
    .A(\u_inv.d_reg[30] ));
 sg13g2_inv_1 _26673_ (.Y(_18585_),
    .A(\u_inv.d_reg[29] ));
 sg13g2_inv_2 _26674_ (.Y(_18586_),
    .A(\u_inv.d_reg[28] ));
 sg13g2_inv_1 _26675_ (.Y(_18587_),
    .A(\u_inv.d_reg[27] ));
 sg13g2_inv_2 _26676_ (.Y(_18588_),
    .A(\u_inv.d_reg[26] ));
 sg13g2_inv_1 _26677_ (.Y(_18589_),
    .A(\u_inv.d_reg[25] ));
 sg13g2_inv_1 _26678_ (.Y(_18590_),
    .A(net3039));
 sg13g2_inv_1 _26679_ (.Y(_18591_),
    .A(\u_inv.d_reg[23] ));
 sg13g2_inv_2 _26680_ (.Y(_18592_),
    .A(net7291));
 sg13g2_inv_1 _26681_ (.Y(_18593_),
    .A(\u_inv.d_reg[21] ));
 sg13g2_inv_2 _26682_ (.Y(_18594_),
    .A(\u_inv.d_reg[20] ));
 sg13g2_inv_2 _26683_ (.Y(_18595_),
    .A(\u_inv.d_reg[19] ));
 sg13g2_inv_2 _26684_ (.Y(_18596_),
    .A(net3598));
 sg13g2_inv_1 _26685_ (.Y(_18597_),
    .A(net3551));
 sg13g2_inv_2 _26686_ (.Y(_18598_),
    .A(\u_inv.d_reg[16] ));
 sg13g2_inv_1 _26687_ (.Y(_18599_),
    .A(\u_inv.d_reg[15] ));
 sg13g2_inv_2 _26688_ (.Y(_18600_),
    .A(\u_inv.d_reg[14] ));
 sg13g2_inv_2 _26689_ (.Y(_18601_),
    .A(net2583));
 sg13g2_inv_1 _26690_ (.Y(_18602_),
    .A(\u_inv.d_reg[12] ));
 sg13g2_inv_1 _26691_ (.Y(_18603_),
    .A(\u_inv.d_reg[11] ));
 sg13g2_inv_1 _26692_ (.Y(_18604_),
    .A(net7292));
 sg13g2_inv_2 _26693_ (.Y(_18605_),
    .A(\u_inv.d_reg[9] ));
 sg13g2_inv_1 _26694_ (.Y(_18606_),
    .A(\u_inv.d_reg[8] ));
 sg13g2_inv_2 _26695_ (.Y(_18607_),
    .A(\u_inv.d_reg[7] ));
 sg13g2_inv_1 _26696_ (.Y(_18608_),
    .A(\u_inv.d_reg[6] ));
 sg13g2_inv_1 _26697_ (.Y(_18609_),
    .A(\u_inv.d_reg[5] ));
 sg13g2_inv_2 _26698_ (.Y(_18610_),
    .A(\u_inv.d_reg[4] ));
 sg13g2_inv_1 _26699_ (.Y(_18611_),
    .A(\u_inv.d_reg[3] ));
 sg13g2_inv_1 _26700_ (.Y(_18612_),
    .A(\u_inv.d_reg[2] ));
 sg13g2_inv_1 _26701_ (.Y(_18613_),
    .A(net2562));
 sg13g2_inv_1 _26702_ (.Y(_18614_),
    .A(net1217));
 sg13g2_nor2b_2 _26703_ (.A(net7413),
    .B_N(net7412),
    .Y(uio_out[1]));
 sg13g2_nor2_1 _26704_ (.A(net7412),
    .B(net7413),
    .Y(_18615_));
 sg13g2_a21oi_1 _26705_ (.A1(net7413),
    .A2(net1179),
    .Y(accepting),
    .B1(net7412));
 sg13g2_nor3_1 _26706_ (.A(net1153),
    .B(net1840),
    .C(net1174),
    .Y(_18616_));
 sg13g2_nand4_1 _26707_ (.B(_18256_),
    .C(net2486),
    .A(net2976),
    .Y(_18617_),
    .D(_18616_));
 sg13g2_nor2b_2 _26708_ (.A(net2610),
    .B_N(net10),
    .Y(_18618_));
 sg13g2_nand2_1 _26709_ (.Y(_18619_),
    .A(inv_done),
    .B(net7413));
 sg13g2_nand3_1 _26710_ (.B(_18618_),
    .C(_18619_),
    .A(accepting),
    .Y(_18620_));
 sg13g2_nor2_1 _26711_ (.A(_18617_),
    .B(net2611),
    .Y(_24690_[0]));
 sg13g2_nand3b_1 _26712_ (.B(uio_out[1]),
    .C(net13),
    .Y(_18621_),
    .A_N(net12));
 sg13g2_mux2_1 _26713_ (.A0(\trng_data[0] ),
    .A1(\shift_reg[264] ),
    .S(net6993),
    .X(uo_out[0]));
 sg13g2_mux2_1 _26714_ (.A0(\trng_data[1] ),
    .A1(\shift_reg[265] ),
    .S(net6993),
    .X(uo_out[1]));
 sg13g2_mux2_1 _26715_ (.A0(\trng_data[2] ),
    .A1(\shift_reg[266] ),
    .S(net6993),
    .X(uo_out[2]));
 sg13g2_mux2_1 _26716_ (.A0(\trng_data[3] ),
    .A1(\shift_reg[267] ),
    .S(net6993),
    .X(uo_out[3]));
 sg13g2_mux2_1 _26717_ (.A0(\trng_data[4] ),
    .A1(\shift_reg[268] ),
    .S(net6993),
    .X(uo_out[4]));
 sg13g2_mux2_1 _26718_ (.A0(\trng_data[5] ),
    .A1(\shift_reg[269] ),
    .S(net6993),
    .X(uo_out[5]));
 sg13g2_mux2_1 _26719_ (.A0(\trng_data[6] ),
    .A1(\shift_reg[270] ),
    .S(net6993),
    .X(uo_out[6]));
 sg13g2_mux2_1 _26720_ (.A0(\trng_data[7] ),
    .A1(\shift_reg[271] ),
    .S(_18621_),
    .X(uo_out[7]));
 sg13g2_nor2b_1 _26721_ (.A(\u_inv.state[0] ),
    .B_N(net1768),
    .Y(_18622_));
 sg13g2_nand2b_1 _26722_ (.Y(_18623_),
    .B(net1768),
    .A_N(\u_inv.state[0] ));
 sg13g2_nor2b_1 _26723_ (.A(net7412),
    .B_N(net7413),
    .Y(_18624_));
 sg13g2_nand2b_2 _26724_ (.Y(_18625_),
    .B(net3747),
    .A_N(net7412));
 sg13g2_nand2_1 _26725_ (.Y(_18626_),
    .A(inv_done),
    .B(_18625_));
 sg13g2_nand3_1 _26726_ (.B(_18622_),
    .C(_18625_),
    .A(net3668),
    .Y(_18627_));
 sg13g2_nand2_1 _26727_ (.Y(_18628_),
    .A(\u_inv.input_valid ),
    .B(_18627_));
 sg13g2_or2_1 _26728_ (.X(_18629_),
    .B(_18628_),
    .A(\u_inv.state[0] ));
 sg13g2_inv_8 _26729_ (.Y(_24689_[0]),
    .A(net6607));
 sg13g2_nand2b_1 _26730_ (.Y(_18630_),
    .B(net2256),
    .A_N(trng_ready));
 sg13g2_a21oi_1 _26731_ (.A1(\u_trng.entropy_bit ),
    .A2(\u_trng.prev_sample ),
    .Y(_18631_),
    .B1(_18630_));
 sg13g2_o21ai_1 _26732_ (.B1(_18631_),
    .Y(_18632_),
    .A1(\u_trng.entropy_bit ),
    .A2(net3514));
 sg13g2_inv_1 _26733_ (.Y(_18633_),
    .A(net6677));
 sg13g2_nand3_1 _26734_ (.B(net1173),
    .C(_18633_),
    .A(net1222),
    .Y(_18634_));
 sg13g2_nand2b_2 _26735_ (.Y(_18635_),
    .B(net11),
    .A_N(rd_prev));
 sg13g2_o21ai_1 _26736_ (.B1(trng_ready),
    .Y(_18636_),
    .A1(net6993),
    .A2(_18635_));
 sg13g2_o21ai_1 _26737_ (.B1(_18636_),
    .Y(_00001_),
    .A1(_18356_),
    .A2(_18634_));
 sg13g2_nand2_1 _26738_ (.Y(_00000_),
    .A(net1769),
    .B(_18626_));
 sg13g2_xnor2_1 _26739_ (.Y(_18637_),
    .A(\u_trng.u_ro5.c[4] ),
    .B(\u_trng.u_ro9.c[8] ));
 sg13g2_xnor2_1 _26740_ (.Y(\u_trng.entropy_raw ),
    .A(\u_trng.u_ro7.c[6] ),
    .B(_18637_));
 sg13g2_nor3_1 _26741_ (.A(\u_inv.load_input ),
    .B(_18181_),
    .C(\u_inv.input_valid ),
    .Y(_18638_));
 sg13g2_mux2_1 _26742_ (.A0(net1797),
    .A1(\shift_reg[111] ),
    .S(net6988),
    .X(_00002_));
 sg13g2_mux2_1 _26743_ (.A0(net1546),
    .A1(\shift_reg[112] ),
    .S(net6980),
    .X(_00003_));
 sg13g2_mux2_1 _26744_ (.A0(net1365),
    .A1(\shift_reg[113] ),
    .S(net6980),
    .X(_00004_));
 sg13g2_mux2_1 _26745_ (.A0(net1658),
    .A1(\shift_reg[114] ),
    .S(net6980),
    .X(_00005_));
 sg13g2_mux2_1 _26746_ (.A0(net1322),
    .A1(\shift_reg[115] ),
    .S(net6980),
    .X(_00006_));
 sg13g2_mux2_1 _26747_ (.A0(net1945),
    .A1(\shift_reg[116] ),
    .S(net6981),
    .X(_00007_));
 sg13g2_mux2_1 _26748_ (.A0(net1800),
    .A1(\shift_reg[117] ),
    .S(net6984),
    .X(_00008_));
 sg13g2_mux2_1 _26749_ (.A0(net1863),
    .A1(\shift_reg[118] ),
    .S(net6981),
    .X(_00009_));
 sg13g2_mux2_1 _26750_ (.A0(net1409),
    .A1(\shift_reg[119] ),
    .S(net6978),
    .X(_00010_));
 sg13g2_mux2_1 _26751_ (.A0(net1682),
    .A1(\shift_reg[120] ),
    .S(net6984),
    .X(_00011_));
 sg13g2_mux2_1 _26752_ (.A0(net1363),
    .A1(\shift_reg[121] ),
    .S(net6980),
    .X(_00012_));
 sg13g2_mux2_1 _26753_ (.A0(net2370),
    .A1(\shift_reg[122] ),
    .S(net6980),
    .X(_00013_));
 sg13g2_mux2_1 _26754_ (.A0(net1276),
    .A1(\shift_reg[123] ),
    .S(net6984),
    .X(_00014_));
 sg13g2_mux2_1 _26755_ (.A0(net1689),
    .A1(\shift_reg[124] ),
    .S(net6982),
    .X(_00015_));
 sg13g2_mux2_1 _26756_ (.A0(net1762),
    .A1(\shift_reg[125] ),
    .S(net6982),
    .X(_00016_));
 sg13g2_mux2_1 _26757_ (.A0(net1592),
    .A1(\shift_reg[126] ),
    .S(net6982),
    .X(_00017_));
 sg13g2_mux2_1 _26758_ (.A0(net1733),
    .A1(\shift_reg[127] ),
    .S(net6982),
    .X(_00018_));
 sg13g2_mux2_1 _26759_ (.A0(net1397),
    .A1(\shift_reg[128] ),
    .S(net6983),
    .X(_00019_));
 sg13g2_mux2_1 _26760_ (.A0(net1535),
    .A1(\shift_reg[129] ),
    .S(net6982),
    .X(_00020_));
 sg13g2_mux2_1 _26761_ (.A0(net1748),
    .A1(\shift_reg[130] ),
    .S(net6981),
    .X(_00021_));
 sg13g2_mux2_1 _26762_ (.A0(net2015),
    .A1(\shift_reg[131] ),
    .S(net6982),
    .X(_00022_));
 sg13g2_mux2_1 _26763_ (.A0(net2512),
    .A1(\shift_reg[132] ),
    .S(net6983),
    .X(_00023_));
 sg13g2_mux2_1 _26764_ (.A0(net1429),
    .A1(\shift_reg[133] ),
    .S(net6976),
    .X(_00024_));
 sg13g2_mux2_1 _26765_ (.A0(net1728),
    .A1(\shift_reg[134] ),
    .S(net6982),
    .X(_00025_));
 sg13g2_mux2_1 _26766_ (.A0(net2569),
    .A1(net2303),
    .S(net6982),
    .X(_00026_));
 sg13g2_mux2_1 _26767_ (.A0(net1316),
    .A1(\shift_reg[136] ),
    .S(net6983),
    .X(_00027_));
 sg13g2_mux2_1 _26768_ (.A0(net2346),
    .A1(net2291),
    .S(net6983),
    .X(_00028_));
 sg13g2_mux2_1 _26769_ (.A0(net1656),
    .A1(\shift_reg[138] ),
    .S(net6977),
    .X(_00029_));
 sg13g2_mux2_1 _26770_ (.A0(net1258),
    .A1(\shift_reg[139] ),
    .S(net6976),
    .X(_00030_));
 sg13g2_mux2_1 _26771_ (.A0(net3170),
    .A1(\shift_reg[140] ),
    .S(net6976),
    .X(_00031_));
 sg13g2_mux2_1 _26772_ (.A0(net3165),
    .A1(\shift_reg[141] ),
    .S(net6976),
    .X(_00032_));
 sg13g2_mux2_1 _26773_ (.A0(net2998),
    .A1(\shift_reg[142] ),
    .S(net6981),
    .X(_00033_));
 sg13g2_mux2_1 _26774_ (.A0(net1906),
    .A1(\shift_reg[143] ),
    .S(net6974),
    .X(_00034_));
 sg13g2_mux2_1 _26775_ (.A0(net2317),
    .A1(\shift_reg[144] ),
    .S(net6974),
    .X(_00035_));
 sg13g2_mux2_1 _26776_ (.A0(net1640),
    .A1(\shift_reg[145] ),
    .S(net6974),
    .X(_00036_));
 sg13g2_mux2_1 _26777_ (.A0(net2399),
    .A1(\shift_reg[146] ),
    .S(net6974),
    .X(_00037_));
 sg13g2_mux2_1 _26778_ (.A0(net1381),
    .A1(\shift_reg[147] ),
    .S(net6974),
    .X(_00038_));
 sg13g2_mux2_1 _26779_ (.A0(net1271),
    .A1(\shift_reg[148] ),
    .S(net6975),
    .X(_00039_));
 sg13g2_mux2_1 _26780_ (.A0(net1531),
    .A1(\shift_reg[149] ),
    .S(net6970),
    .X(_00040_));
 sg13g2_mux2_1 _26781_ (.A0(net1685),
    .A1(\shift_reg[150] ),
    .S(net6970),
    .X(_00041_));
 sg13g2_mux2_1 _26782_ (.A0(net2552),
    .A1(\shift_reg[151] ),
    .S(net6971),
    .X(_00042_));
 sg13g2_mux2_1 _26783_ (.A0(net2600),
    .A1(\shift_reg[152] ),
    .S(net6972),
    .X(_00043_));
 sg13g2_mux2_1 _26784_ (.A0(net2969),
    .A1(\shift_reg[153] ),
    .S(net6972),
    .X(_00044_));
 sg13g2_mux2_1 _26785_ (.A0(net2229),
    .A1(\shift_reg[154] ),
    .S(net6971),
    .X(_00045_));
 sg13g2_mux2_1 _26786_ (.A0(net2473),
    .A1(\shift_reg[155] ),
    .S(net6972),
    .X(_00046_));
 sg13g2_mux2_1 _26787_ (.A0(net1911),
    .A1(\shift_reg[156] ),
    .S(net6972),
    .X(_00047_));
 sg13g2_mux2_1 _26788_ (.A0(net2262),
    .A1(\shift_reg[157] ),
    .S(net6972),
    .X(_00048_));
 sg13g2_mux2_1 _26789_ (.A0(net1960),
    .A1(\shift_reg[158] ),
    .S(net6969),
    .X(_00049_));
 sg13g2_mux2_1 _26790_ (.A0(net1337),
    .A1(\shift_reg[159] ),
    .S(net6969),
    .X(_00050_));
 sg13g2_mux2_1 _26791_ (.A0(net2362),
    .A1(\shift_reg[160] ),
    .S(net6968),
    .X(_00051_));
 sg13g2_mux2_1 _26792_ (.A0(net2357),
    .A1(\shift_reg[161] ),
    .S(net6970),
    .X(_00052_));
 sg13g2_mux2_1 _26793_ (.A0(net2791),
    .A1(\shift_reg[162] ),
    .S(net6970),
    .X(_00053_));
 sg13g2_mux2_1 _26794_ (.A0(net2495),
    .A1(\shift_reg[163] ),
    .S(net6970),
    .X(_00054_));
 sg13g2_mux2_1 _26795_ (.A0(net1885),
    .A1(\shift_reg[164] ),
    .S(net6970),
    .X(_00055_));
 sg13g2_mux2_1 _26796_ (.A0(net2892),
    .A1(\shift_reg[165] ),
    .S(net6968),
    .X(_00056_));
 sg13g2_mux2_1 _26797_ (.A0(net1804),
    .A1(\shift_reg[166] ),
    .S(net6969),
    .X(_00057_));
 sg13g2_mux2_1 _26798_ (.A0(net2238),
    .A1(\shift_reg[167] ),
    .S(net6969),
    .X(_00058_));
 sg13g2_mux2_1 _26799_ (.A0(net1498),
    .A1(\shift_reg[168] ),
    .S(net6970),
    .X(_00059_));
 sg13g2_mux2_1 _26800_ (.A0(net1555),
    .A1(\shift_reg[169] ),
    .S(net6969),
    .X(_00060_));
 sg13g2_mux2_1 _26801_ (.A0(net2041),
    .A1(\shift_reg[170] ),
    .S(net6968),
    .X(_00061_));
 sg13g2_mux2_1 _26802_ (.A0(net2089),
    .A1(\shift_reg[171] ),
    .S(net6966),
    .X(_00062_));
 sg13g2_mux2_1 _26803_ (.A0(net1413),
    .A1(\shift_reg[172] ),
    .S(net6968),
    .X(_00063_));
 sg13g2_mux2_1 _26804_ (.A0(net2021),
    .A1(\shift_reg[173] ),
    .S(net6968),
    .X(_00064_));
 sg13g2_mux2_1 _26805_ (.A0(net1502),
    .A1(\shift_reg[174] ),
    .S(net6968),
    .X(_00065_));
 sg13g2_mux2_1 _26806_ (.A0(net2048),
    .A1(\shift_reg[175] ),
    .S(net6968),
    .X(_00066_));
 sg13g2_mux2_1 _26807_ (.A0(net2477),
    .A1(\shift_reg[176] ),
    .S(net6966),
    .X(_00067_));
 sg13g2_mux2_1 _26808_ (.A0(net1561),
    .A1(\shift_reg[177] ),
    .S(net6965),
    .X(_00068_));
 sg13g2_mux2_1 _26809_ (.A0(net1454),
    .A1(\shift_reg[178] ),
    .S(net6965),
    .X(_00069_));
 sg13g2_mux2_1 _26810_ (.A0(net3019),
    .A1(net2793),
    .S(net6966),
    .X(_00070_));
 sg13g2_mux2_1 _26811_ (.A0(net1980),
    .A1(\shift_reg[180] ),
    .S(net6965),
    .X(_00071_));
 sg13g2_mux2_1 _26812_ (.A0(net1883),
    .A1(\shift_reg[181] ),
    .S(net6965),
    .X(_00072_));
 sg13g2_mux2_1 _26813_ (.A0(net1356),
    .A1(\shift_reg[182] ),
    .S(net6964),
    .X(_00073_));
 sg13g2_mux2_1 _26814_ (.A0(net1516),
    .A1(\shift_reg[183] ),
    .S(net6964),
    .X(_00074_));
 sg13g2_mux2_1 _26815_ (.A0(net2353),
    .A1(\shift_reg[184] ),
    .S(net6962),
    .X(_00075_));
 sg13g2_mux2_1 _26816_ (.A0(net2639),
    .A1(net2282),
    .S(net6963),
    .X(_00076_));
 sg13g2_mux2_1 _26817_ (.A0(net1930),
    .A1(\shift_reg[186] ),
    .S(net6963),
    .X(_00077_));
 sg13g2_mux2_1 _26818_ (.A0(net1519),
    .A1(\shift_reg[187] ),
    .S(net6963),
    .X(_00078_));
 sg13g2_mux2_1 _26819_ (.A0(net1329),
    .A1(\shift_reg[188] ),
    .S(net6962),
    .X(_00079_));
 sg13g2_mux2_1 _26820_ (.A0(net1287),
    .A1(\shift_reg[189] ),
    .S(net6963),
    .X(_00080_));
 sg13g2_mux2_1 _26821_ (.A0(net1630),
    .A1(\shift_reg[190] ),
    .S(net6963),
    .X(_00081_));
 sg13g2_mux2_1 _26822_ (.A0(net1978),
    .A1(\shift_reg[191] ),
    .S(net6963),
    .X(_00082_));
 sg13g2_mux2_1 _26823_ (.A0(net1551),
    .A1(\shift_reg[192] ),
    .S(net6959),
    .X(_00083_));
 sg13g2_mux2_1 _26824_ (.A0(net1570),
    .A1(\shift_reg[193] ),
    .S(net6959),
    .X(_00084_));
 sg13g2_mux2_1 _26825_ (.A0(net1404),
    .A1(\shift_reg[194] ),
    .S(net6959),
    .X(_00085_));
 sg13g2_mux2_1 _26826_ (.A0(net1581),
    .A1(\shift_reg[195] ),
    .S(net6960),
    .X(_00086_));
 sg13g2_mux2_1 _26827_ (.A0(net1544),
    .A1(\shift_reg[196] ),
    .S(net6960),
    .X(_00087_));
 sg13g2_mux2_1 _26828_ (.A0(net1393),
    .A1(\shift_reg[197] ),
    .S(net6960),
    .X(_00088_));
 sg13g2_mux2_1 _26829_ (.A0(net1835),
    .A1(\shift_reg[198] ),
    .S(net6960),
    .X(_00089_));
 sg13g2_mux2_1 _26830_ (.A0(net2289),
    .A1(\shift_reg[199] ),
    .S(net6960),
    .X(_00090_));
 sg13g2_mux2_1 _26831_ (.A0(net1812),
    .A1(\shift_reg[200] ),
    .S(net6958),
    .X(_00091_));
 sg13g2_mux2_1 _26832_ (.A0(net1817),
    .A1(\shift_reg[201] ),
    .S(net6958),
    .X(_00092_));
 sg13g2_mux2_1 _26833_ (.A0(net2059),
    .A1(\shift_reg[202] ),
    .S(net6958),
    .X(_00093_));
 sg13g2_mux2_1 _26834_ (.A0(net2312),
    .A1(net2277),
    .S(net6959),
    .X(_00094_));
 sg13g2_mux2_1 _26835_ (.A0(net1872),
    .A1(\shift_reg[204] ),
    .S(net6961),
    .X(_00095_));
 sg13g2_mux2_1 _26836_ (.A0(net2382),
    .A1(net2248),
    .S(net6958),
    .X(_00096_));
 sg13g2_mux2_1 _26837_ (.A0(net1999),
    .A1(\shift_reg[206] ),
    .S(net6958),
    .X(_00097_));
 sg13g2_mux2_1 _26838_ (.A0(net1462),
    .A1(\shift_reg[207] ),
    .S(net6958),
    .X(_00098_));
 sg13g2_mux2_1 _26839_ (.A0(net1282),
    .A1(\shift_reg[208] ),
    .S(net6951),
    .X(_00099_));
 sg13g2_mux2_1 _26840_ (.A0(net1806),
    .A1(\shift_reg[209] ),
    .S(net6952),
    .X(_00100_));
 sg13g2_mux2_1 _26841_ (.A0(net1713),
    .A1(\shift_reg[210] ),
    .S(net6951),
    .X(_00101_));
 sg13g2_mux2_1 _26842_ (.A0(net1783),
    .A1(\shift_reg[211] ),
    .S(net6951),
    .X(_00102_));
 sg13g2_mux2_1 _26843_ (.A0(net1704),
    .A1(\shift_reg[212] ),
    .S(net6951),
    .X(_00103_));
 sg13g2_mux2_1 _26844_ (.A0(net1833),
    .A1(\shift_reg[213] ),
    .S(net6951),
    .X(_00104_));
 sg13g2_mux2_1 _26845_ (.A0(net1456),
    .A1(\shift_reg[214] ),
    .S(net6951),
    .X(_00105_));
 sg13g2_mux2_1 _26846_ (.A0(net1425),
    .A1(\shift_reg[215] ),
    .S(net6951),
    .X(_00106_));
 sg13g2_mux2_1 _26847_ (.A0(net1340),
    .A1(\shift_reg[216] ),
    .S(net6946),
    .X(_00107_));
 sg13g2_mux2_1 _26848_ (.A0(net2759),
    .A1(net2171),
    .S(net6952),
    .X(_00108_));
 sg13g2_mux2_1 _26849_ (.A0(net1660),
    .A1(\shift_reg[218] ),
    .S(net6946),
    .X(_00109_));
 sg13g2_mux2_1 _26850_ (.A0(net2785),
    .A1(net2728),
    .S(net6952),
    .X(_00110_));
 sg13g2_mux2_1 _26851_ (.A0(net2484),
    .A1(\shift_reg[220] ),
    .S(net6947),
    .X(_00111_));
 sg13g2_mux2_1 _26852_ (.A0(net2260),
    .A1(\shift_reg[221] ),
    .S(net6946),
    .X(_00112_));
 sg13g2_mux2_1 _26853_ (.A0(net1928),
    .A1(\shift_reg[222] ),
    .S(net6947),
    .X(_00113_));
 sg13g2_mux2_1 _26854_ (.A0(net2718),
    .A1(\shift_reg[223] ),
    .S(net6951),
    .X(_00114_));
 sg13g2_mux2_1 _26855_ (.A0(net1481),
    .A1(\shift_reg[224] ),
    .S(net6946),
    .X(_00115_));
 sg13g2_mux2_1 _26856_ (.A0(net2301),
    .A1(\shift_reg[225] ),
    .S(net6946),
    .X(_00116_));
 sg13g2_mux2_1 _26857_ (.A0(net1528),
    .A1(\shift_reg[226] ),
    .S(net6946),
    .X(_00117_));
 sg13g2_nand2_1 _26858_ (.Y(_18639_),
    .A(\shift_reg[227] ),
    .B(net6948));
 sg13g2_o21ai_1 _26859_ (.B1(_18639_),
    .Y(_00118_),
    .A1(_18614_),
    .A2(net6946));
 sg13g2_mux2_1 _26860_ (.A0(net1699),
    .A1(\shift_reg[228] ),
    .S(net6948),
    .X(_00119_));
 sg13g2_mux2_1 _26861_ (.A0(net2457),
    .A1(\shift_reg[229] ),
    .S(net6947),
    .X(_00120_));
 sg13g2_mux2_1 _26862_ (.A0(net2272),
    .A1(\shift_reg[230] ),
    .S(net6946),
    .X(_00121_));
 sg13g2_mux2_1 _26863_ (.A0(net1628),
    .A1(\shift_reg[231] ),
    .S(net6948),
    .X(_00122_));
 sg13g2_mux2_1 _26864_ (.A0(net1625),
    .A1(\shift_reg[232] ),
    .S(net6948),
    .X(_00123_));
 sg13g2_mux2_1 _26865_ (.A0(net1310),
    .A1(\shift_reg[233] ),
    .S(net6948),
    .X(_00124_));
 sg13g2_mux2_1 _26866_ (.A0(net1469),
    .A1(\shift_reg[234] ),
    .S(net6948),
    .X(_00125_));
 sg13g2_mux2_1 _26867_ (.A0(net2523),
    .A1(\shift_reg[235] ),
    .S(net6948),
    .X(_00126_));
 sg13g2_mux2_1 _26868_ (.A0(net1312),
    .A1(\shift_reg[236] ),
    .S(net6948),
    .X(_00127_));
 sg13g2_mux2_1 _26869_ (.A0(net1868),
    .A1(\shift_reg[237] ),
    .S(net6949),
    .X(_00128_));
 sg13g2_mux2_1 _26870_ (.A0(net1795),
    .A1(\shift_reg[238] ),
    .S(net6950),
    .X(_00129_));
 sg13g2_mux2_1 _26871_ (.A0(net2673),
    .A1(net1851),
    .S(net6949),
    .X(_00130_));
 sg13g2_mux2_1 _26872_ (.A0(net1399),
    .A1(\shift_reg[240] ),
    .S(net6949),
    .X(_00131_));
 sg13g2_mux2_1 _26873_ (.A0(net1838),
    .A1(\shift_reg[241] ),
    .S(net6949),
    .X(_00132_));
 sg13g2_mux2_1 _26874_ (.A0(net1395),
    .A1(\shift_reg[242] ),
    .S(net6949),
    .X(_00133_));
 sg13g2_mux2_1 _26875_ (.A0(net1652),
    .A1(\shift_reg[243] ),
    .S(net6949),
    .X(_00134_));
 sg13g2_mux2_1 _26876_ (.A0(net1559),
    .A1(\shift_reg[244] ),
    .S(net6949),
    .X(_00135_));
 sg13g2_mux2_1 _26877_ (.A0(net1610),
    .A1(\shift_reg[245] ),
    .S(net6949),
    .X(_00136_));
 sg13g2_mux2_1 _26878_ (.A0(net1401),
    .A1(\shift_reg[246] ),
    .S(net6953),
    .X(_00137_));
 sg13g2_mux2_1 _26879_ (.A0(net2093),
    .A1(\shift_reg[247] ),
    .S(net6953),
    .X(_00138_));
 sg13g2_mux2_1 _26880_ (.A0(net1385),
    .A1(\shift_reg[248] ),
    .S(net6953),
    .X(_00139_));
 sg13g2_mux2_1 _26881_ (.A0(net1377),
    .A1(\shift_reg[249] ),
    .S(net6953),
    .X(_00140_));
 sg13g2_mux2_1 _26882_ (.A0(net1514),
    .A1(\shift_reg[250] ),
    .S(net6953),
    .X(_00141_));
 sg13g2_mux2_1 _26883_ (.A0(net1942),
    .A1(\shift_reg[251] ),
    .S(net6954),
    .X(_00142_));
 sg13g2_mux2_1 _26884_ (.A0(net1438),
    .A1(\shift_reg[252] ),
    .S(net6953),
    .X(_00143_));
 sg13g2_mux2_1 _26885_ (.A0(net1289),
    .A1(\shift_reg[253] ),
    .S(net6953),
    .X(_00144_));
 sg13g2_mux2_1 _26886_ (.A0(net1604),
    .A1(\shift_reg[254] ),
    .S(net6954),
    .X(_00145_));
 sg13g2_mux2_1 _26887_ (.A0(net1333),
    .A1(\shift_reg[255] ),
    .S(net6954),
    .X(_00146_));
 sg13g2_mux2_1 _26888_ (.A0(net1327),
    .A1(\shift_reg[256] ),
    .S(net6954),
    .X(_00147_));
 sg13g2_mux2_1 _26889_ (.A0(net1320),
    .A1(\shift_reg[257] ),
    .S(net6953),
    .X(_00148_));
 sg13g2_mux2_1 _26890_ (.A0(net1475),
    .A1(\shift_reg[258] ),
    .S(net6954),
    .X(_00149_));
 sg13g2_mux2_1 _26891_ (.A0(net1427),
    .A1(\shift_reg[259] ),
    .S(net6955),
    .X(_00150_));
 sg13g2_mux2_1 _26892_ (.A0(net1706),
    .A1(\shift_reg[260] ),
    .S(net6955),
    .X(_00151_));
 sg13g2_mux2_1 _26893_ (.A0(net1564),
    .A1(\shift_reg[261] ),
    .S(net6956),
    .X(_00152_));
 sg13g2_mux2_1 _26894_ (.A0(net1367),
    .A1(\shift_reg[262] ),
    .S(net6955),
    .X(_00153_));
 sg13g2_mux2_1 _26895_ (.A0(net1308),
    .A1(\shift_reg[263] ),
    .S(net6956),
    .X(_00154_));
 sg13g2_mux2_1 _26896_ (.A0(net1715),
    .A1(\shift_reg[264] ),
    .S(net6955),
    .X(_00155_));
 sg13g2_mux2_1 _26897_ (.A0(net1989),
    .A1(\shift_reg[265] ),
    .S(net6955),
    .X(_00156_));
 sg13g2_mux2_1 _26898_ (.A0(net2323),
    .A1(\shift_reg[266] ),
    .S(net6955),
    .X(_00157_));
 sg13g2_mux2_1 _26899_ (.A0(net1963),
    .A1(\shift_reg[267] ),
    .S(net6955),
    .X(_00158_));
 sg13g2_mux2_1 _26900_ (.A0(net2505),
    .A1(\shift_reg[268] ),
    .S(net6955),
    .X(_00159_));
 sg13g2_mux2_1 _26901_ (.A0(net1314),
    .A1(\shift_reg[269] ),
    .S(net6956),
    .X(_00160_));
 sg13g2_mux2_1 _26902_ (.A0(net1775),
    .A1(\shift_reg[270] ),
    .S(net6956),
    .X(_00161_));
 sg13g2_mux2_1 _26903_ (.A0(net1802),
    .A1(\shift_reg[271] ),
    .S(net6956),
    .X(_00162_));
 sg13g2_nor2_1 _26904_ (.A(net1159),
    .B(parity_error),
    .Y(_18640_));
 sg13g2_xnor2_1 _26905_ (.Y(_18641_),
    .A(\shift_reg[90] ),
    .B(\shift_reg[91] ));
 sg13g2_xor2_1 _26906_ (.B(\shift_reg[89] ),
    .A(\shift_reg[88] ),
    .X(_18642_));
 sg13g2_xnor2_1 _26907_ (.Y(_18643_),
    .A(_18641_),
    .B(_18642_));
 sg13g2_xnor2_1 _26908_ (.Y(_18644_),
    .A(\shift_reg[94] ),
    .B(\shift_reg[95] ));
 sg13g2_xor2_1 _26909_ (.B(\shift_reg[93] ),
    .A(\shift_reg[92] ),
    .X(_18645_));
 sg13g2_xnor2_1 _26910_ (.Y(_18646_),
    .A(_18644_),
    .B(_18645_));
 sg13g2_xnor2_1 _26911_ (.Y(_18647_),
    .A(_18643_),
    .B(_18646_));
 sg13g2_xor2_1 _26912_ (.B(\shift_reg[83] ),
    .A(\shift_reg[82] ),
    .X(_18648_));
 sg13g2_xor2_1 _26913_ (.B(\shift_reg[81] ),
    .A(\shift_reg[80] ),
    .X(_18649_));
 sg13g2_xnor2_1 _26914_ (.Y(_18650_),
    .A(_18648_),
    .B(_18649_));
 sg13g2_xnor2_1 _26915_ (.Y(_18651_),
    .A(\shift_reg[86] ),
    .B(\shift_reg[87] ));
 sg13g2_xor2_1 _26916_ (.B(\shift_reg[85] ),
    .A(\shift_reg[84] ),
    .X(_18652_));
 sg13g2_xnor2_1 _26917_ (.Y(_18653_),
    .A(_18651_),
    .B(_18652_));
 sg13g2_xnor2_1 _26918_ (.Y(_18654_),
    .A(_18650_),
    .B(_18653_));
 sg13g2_xnor2_1 _26919_ (.Y(_18655_),
    .A(_18647_),
    .B(_18654_));
 sg13g2_xnor2_1 _26920_ (.Y(_18656_),
    .A(\shift_reg[26] ),
    .B(\shift_reg[27] ));
 sg13g2_xor2_1 _26921_ (.B(\shift_reg[25] ),
    .A(\shift_reg[24] ),
    .X(_18657_));
 sg13g2_xnor2_1 _26922_ (.Y(_18658_),
    .A(_18656_),
    .B(_18657_));
 sg13g2_xnor2_1 _26923_ (.Y(_18659_),
    .A(\shift_reg[30] ),
    .B(\shift_reg[31] ));
 sg13g2_xor2_1 _26924_ (.B(\shift_reg[29] ),
    .A(\shift_reg[28] ),
    .X(_18660_));
 sg13g2_xnor2_1 _26925_ (.Y(_18661_),
    .A(_18659_),
    .B(_18660_));
 sg13g2_xnor2_1 _26926_ (.Y(_18662_),
    .A(_18658_),
    .B(_18661_));
 sg13g2_xor2_1 _26927_ (.B(\shift_reg[19] ),
    .A(\shift_reg[18] ),
    .X(_18663_));
 sg13g2_xor2_1 _26928_ (.B(\shift_reg[17] ),
    .A(\shift_reg[16] ),
    .X(_18664_));
 sg13g2_xnor2_1 _26929_ (.Y(_18665_),
    .A(_18663_),
    .B(_18664_));
 sg13g2_xnor2_1 _26930_ (.Y(_18666_),
    .A(\shift_reg[22] ),
    .B(\shift_reg[23] ));
 sg13g2_xor2_1 _26931_ (.B(\shift_reg[21] ),
    .A(\shift_reg[20] ),
    .X(_18667_));
 sg13g2_xnor2_1 _26932_ (.Y(_18668_),
    .A(_18666_),
    .B(_18667_));
 sg13g2_xnor2_1 _26933_ (.Y(_18669_),
    .A(_18665_),
    .B(_18668_));
 sg13g2_xnor2_1 _26934_ (.Y(_18670_),
    .A(_18662_),
    .B(_18669_));
 sg13g2_xnor2_1 _26935_ (.Y(_18671_),
    .A(\shift_reg[106] ),
    .B(\shift_reg[107] ));
 sg13g2_xor2_1 _26936_ (.B(\shift_reg[105] ),
    .A(\shift_reg[104] ),
    .X(_18672_));
 sg13g2_xnor2_1 _26937_ (.Y(_18673_),
    .A(_18671_),
    .B(_18672_));
 sg13g2_xnor2_1 _26938_ (.Y(_18674_),
    .A(\shift_reg[110] ),
    .B(\shift_reg[111] ));
 sg13g2_xor2_1 _26939_ (.B(\shift_reg[109] ),
    .A(\shift_reg[108] ),
    .X(_18675_));
 sg13g2_xnor2_1 _26940_ (.Y(_18676_),
    .A(_18674_),
    .B(_18675_));
 sg13g2_xnor2_1 _26941_ (.Y(_18677_),
    .A(_18673_),
    .B(_18676_));
 sg13g2_xor2_1 _26942_ (.B(\shift_reg[99] ),
    .A(\shift_reg[98] ),
    .X(_18678_));
 sg13g2_xor2_1 _26943_ (.B(\shift_reg[97] ),
    .A(\shift_reg[96] ),
    .X(_18679_));
 sg13g2_xnor2_1 _26944_ (.Y(_18680_),
    .A(_18678_),
    .B(_18679_));
 sg13g2_xnor2_1 _26945_ (.Y(_18681_),
    .A(\shift_reg[102] ),
    .B(\shift_reg[103] ));
 sg13g2_xor2_1 _26946_ (.B(\shift_reg[101] ),
    .A(\shift_reg[100] ),
    .X(_18682_));
 sg13g2_xnor2_1 _26947_ (.Y(_18683_),
    .A(_18681_),
    .B(_18682_));
 sg13g2_xnor2_1 _26948_ (.Y(_18684_),
    .A(_18680_),
    .B(_18683_));
 sg13g2_xnor2_1 _26949_ (.Y(_18685_),
    .A(_18677_),
    .B(_18684_));
 sg13g2_xnor2_1 _26950_ (.Y(_18686_),
    .A(\shift_reg[58] ),
    .B(\shift_reg[59] ));
 sg13g2_xor2_1 _26951_ (.B(\shift_reg[57] ),
    .A(\shift_reg[56] ),
    .X(_18687_));
 sg13g2_xnor2_1 _26952_ (.Y(_18688_),
    .A(_18686_),
    .B(_18687_));
 sg13g2_xnor2_1 _26953_ (.Y(_18689_),
    .A(\shift_reg[62] ),
    .B(\shift_reg[63] ));
 sg13g2_xor2_1 _26954_ (.B(\shift_reg[61] ),
    .A(\shift_reg[60] ),
    .X(_18690_));
 sg13g2_xnor2_1 _26955_ (.Y(_18691_),
    .A(_18689_),
    .B(_18690_));
 sg13g2_xnor2_1 _26956_ (.Y(_18692_),
    .A(_18688_),
    .B(_18691_));
 sg13g2_xor2_1 _26957_ (.B(\shift_reg[51] ),
    .A(\shift_reg[50] ),
    .X(_18693_));
 sg13g2_xor2_1 _26958_ (.B(\shift_reg[49] ),
    .A(\shift_reg[48] ),
    .X(_18694_));
 sg13g2_xnor2_1 _26959_ (.Y(_18695_),
    .A(_18693_),
    .B(_18694_));
 sg13g2_xnor2_1 _26960_ (.Y(_18696_),
    .A(\shift_reg[54] ),
    .B(\shift_reg[55] ));
 sg13g2_xor2_1 _26961_ (.B(\shift_reg[53] ),
    .A(\shift_reg[52] ),
    .X(_18697_));
 sg13g2_xnor2_1 _26962_ (.Y(_18698_),
    .A(_18696_),
    .B(_18697_));
 sg13g2_xnor2_1 _26963_ (.Y(_18699_),
    .A(_18695_),
    .B(_18698_));
 sg13g2_xnor2_1 _26964_ (.Y(_18700_),
    .A(_18692_),
    .B(_18699_));
 sg13g2_xnor2_1 _26965_ (.Y(_18701_),
    .A(_18655_),
    .B(_18685_));
 sg13g2_xnor2_1 _26966_ (.Y(_18702_),
    .A(_18670_),
    .B(_18700_));
 sg13g2_xnor2_1 _26967_ (.Y(_18703_),
    .A(_18701_),
    .B(_18702_));
 sg13g2_xor2_1 _26968_ (.B(\shift_reg[43] ),
    .A(\shift_reg[42] ),
    .X(_18704_));
 sg13g2_xor2_1 _26969_ (.B(\shift_reg[41] ),
    .A(\shift_reg[40] ),
    .X(_18705_));
 sg13g2_xnor2_1 _26970_ (.Y(_18706_),
    .A(_18704_),
    .B(_18705_));
 sg13g2_xnor2_1 _26971_ (.Y(_18707_),
    .A(\shift_reg[46] ),
    .B(\shift_reg[47] ));
 sg13g2_xor2_1 _26972_ (.B(\shift_reg[45] ),
    .A(\shift_reg[44] ),
    .X(_18708_));
 sg13g2_xnor2_1 _26973_ (.Y(_18709_),
    .A(_18707_),
    .B(_18708_));
 sg13g2_xnor2_1 _26974_ (.Y(_18710_),
    .A(_18706_),
    .B(_18709_));
 sg13g2_xor2_1 _26975_ (.B(\shift_reg[35] ),
    .A(\shift_reg[34] ),
    .X(_18711_));
 sg13g2_xor2_1 _26976_ (.B(\shift_reg[33] ),
    .A(\shift_reg[32] ),
    .X(_18712_));
 sg13g2_xnor2_1 _26977_ (.Y(_18713_),
    .A(_18711_),
    .B(_18712_));
 sg13g2_xnor2_1 _26978_ (.Y(_18714_),
    .A(\shift_reg[38] ),
    .B(\shift_reg[39] ));
 sg13g2_xor2_1 _26979_ (.B(\shift_reg[37] ),
    .A(\shift_reg[36] ),
    .X(_18715_));
 sg13g2_xnor2_1 _26980_ (.Y(_18716_),
    .A(_18714_),
    .B(_18715_));
 sg13g2_xnor2_1 _26981_ (.Y(_18717_),
    .A(_18713_),
    .B(_18716_));
 sg13g2_xnor2_1 _26982_ (.Y(_18718_),
    .A(_18710_),
    .B(_18717_));
 sg13g2_xnor2_1 _26983_ (.Y(_18719_),
    .A(\shift_reg[66] ),
    .B(\shift_reg[67] ));
 sg13g2_xor2_1 _26984_ (.B(\shift_reg[65] ),
    .A(\shift_reg[64] ),
    .X(_18720_));
 sg13g2_xnor2_1 _26985_ (.Y(_18721_),
    .A(_18719_),
    .B(_18720_));
 sg13g2_xnor2_1 _26986_ (.Y(_18722_),
    .A(\shift_reg[70] ),
    .B(\shift_reg[71] ));
 sg13g2_xor2_1 _26987_ (.B(\shift_reg[69] ),
    .A(\shift_reg[68] ),
    .X(_18723_));
 sg13g2_xnor2_1 _26988_ (.Y(_18724_),
    .A(_18722_),
    .B(_18723_));
 sg13g2_xnor2_1 _26989_ (.Y(_18725_),
    .A(_18721_),
    .B(_18724_));
 sg13g2_xnor2_1 _26990_ (.Y(_18726_),
    .A(\shift_reg[124] ),
    .B(\shift_reg[125] ));
 sg13g2_xor2_1 _26991_ (.B(\shift_reg[123] ),
    .A(\shift_reg[122] ),
    .X(_18727_));
 sg13g2_xor2_1 _26992_ (.B(\shift_reg[121] ),
    .A(\shift_reg[120] ),
    .X(_18728_));
 sg13g2_xnor2_1 _26993_ (.Y(_18729_),
    .A(_18727_),
    .B(_18728_));
 sg13g2_xnor2_1 _26994_ (.Y(_18730_),
    .A(\shift_reg[126] ),
    .B(\shift_reg[127] ));
 sg13g2_xnor2_1 _26995_ (.Y(_18731_),
    .A(_18726_),
    .B(_18730_));
 sg13g2_xnor2_1 _26996_ (.Y(_18732_),
    .A(_18729_),
    .B(_18731_));
 sg13g2_xnor2_1 _26997_ (.Y(_18733_),
    .A(\shift_reg[118] ),
    .B(\shift_reg[119] ));
 sg13g2_xor2_1 _26998_ (.B(\shift_reg[117] ),
    .A(\shift_reg[116] ),
    .X(_18734_));
 sg13g2_xnor2_1 _26999_ (.Y(_18735_),
    .A(_18733_),
    .B(_18734_));
 sg13g2_xor2_1 _27000_ (.B(\shift_reg[115] ),
    .A(\shift_reg[114] ),
    .X(_18736_));
 sg13g2_xor2_1 _27001_ (.B(\shift_reg[113] ),
    .A(\shift_reg[112] ),
    .X(_18737_));
 sg13g2_xnor2_1 _27002_ (.Y(_18738_),
    .A(_18736_),
    .B(_18737_));
 sg13g2_xor2_1 _27003_ (.B(\shift_reg[139] ),
    .A(\shift_reg[138] ),
    .X(_18739_));
 sg13g2_xor2_1 _27004_ (.B(\shift_reg[137] ),
    .A(\shift_reg[136] ),
    .X(_18740_));
 sg13g2_xnor2_1 _27005_ (.Y(_18741_),
    .A(_18739_),
    .B(_18740_));
 sg13g2_xnor2_1 _27006_ (.Y(_18742_),
    .A(_18735_),
    .B(_18738_));
 sg13g2_xnor2_1 _27007_ (.Y(_18743_),
    .A(_18732_),
    .B(_18742_));
 sg13g2_xnor2_1 _27008_ (.Y(_18744_),
    .A(\shift_reg[134] ),
    .B(\shift_reg[135] ));
 sg13g2_xnor2_1 _27009_ (.Y(_18745_),
    .A(\shift_reg[15] ),
    .B(_18744_));
 sg13g2_xnor2_1 _27010_ (.Y(_18746_),
    .A(\shift_reg[128] ),
    .B(\shift_reg[129] ));
 sg13g2_xnor2_1 _27011_ (.Y(_18747_),
    .A(\shift_reg[132] ),
    .B(\shift_reg[133] ));
 sg13g2_xnor2_1 _27012_ (.Y(_18748_),
    .A(_18746_),
    .B(_18747_));
 sg13g2_xor2_1 _27013_ (.B(\shift_reg[131] ),
    .A(\shift_reg[130] ),
    .X(_18749_));
 sg13g2_xor2_1 _27014_ (.B(\shift_reg[143] ),
    .A(\shift_reg[142] ),
    .X(_18750_));
 sg13g2_xor2_1 _27015_ (.B(\shift_reg[141] ),
    .A(\shift_reg[140] ),
    .X(_18751_));
 sg13g2_xnor2_1 _27016_ (.Y(_18752_),
    .A(_18750_),
    .B(_18751_));
 sg13g2_xnor2_1 _27017_ (.Y(_18753_),
    .A(_18748_),
    .B(_18749_));
 sg13g2_xnor2_1 _27018_ (.Y(_18754_),
    .A(_18745_),
    .B(_18753_));
 sg13g2_xnor2_1 _27019_ (.Y(_18755_),
    .A(_18741_),
    .B(_18752_));
 sg13g2_xnor2_1 _27020_ (.Y(_18756_),
    .A(_18743_),
    .B(_18755_));
 sg13g2_xnor2_1 _27021_ (.Y(_18757_),
    .A(_18754_),
    .B(_18756_));
 sg13g2_xor2_1 _27022_ (.B(\shift_reg[251] ),
    .A(\shift_reg[250] ),
    .X(_18758_));
 sg13g2_xor2_1 _27023_ (.B(\shift_reg[249] ),
    .A(\shift_reg[248] ),
    .X(_18759_));
 sg13g2_xnor2_1 _27024_ (.Y(_18760_),
    .A(_18758_),
    .B(_18759_));
 sg13g2_xnor2_1 _27025_ (.Y(_18761_),
    .A(\shift_reg[254] ),
    .B(\shift_reg[255] ));
 sg13g2_xor2_1 _27026_ (.B(\shift_reg[253] ),
    .A(\shift_reg[252] ),
    .X(_18762_));
 sg13g2_xnor2_1 _27027_ (.Y(_18763_),
    .A(_18761_),
    .B(_18762_));
 sg13g2_xnor2_1 _27028_ (.Y(_18764_),
    .A(_18760_),
    .B(_18763_));
 sg13g2_xor2_1 _27029_ (.B(\shift_reg[243] ),
    .A(\shift_reg[242] ),
    .X(_18765_));
 sg13g2_xor2_1 _27030_ (.B(\shift_reg[241] ),
    .A(\shift_reg[240] ),
    .X(_18766_));
 sg13g2_xnor2_1 _27031_ (.Y(_18767_),
    .A(_18765_),
    .B(_18766_));
 sg13g2_xnor2_1 _27032_ (.Y(_18768_),
    .A(\shift_reg[246] ),
    .B(\shift_reg[247] ));
 sg13g2_xor2_1 _27033_ (.B(\shift_reg[245] ),
    .A(\shift_reg[244] ),
    .X(_18769_));
 sg13g2_xnor2_1 _27034_ (.Y(_18770_),
    .A(_18768_),
    .B(_18769_));
 sg13g2_xnor2_1 _27035_ (.Y(_18771_),
    .A(_18767_),
    .B(_18770_));
 sg13g2_xnor2_1 _27036_ (.Y(_18772_),
    .A(_18764_),
    .B(_18771_));
 sg13g2_xor2_1 _27037_ (.B(\shift_reg[267] ),
    .A(\shift_reg[266] ),
    .X(_18773_));
 sg13g2_xor2_1 _27038_ (.B(\shift_reg[265] ),
    .A(\shift_reg[264] ),
    .X(_18774_));
 sg13g2_xnor2_1 _27039_ (.Y(_18775_),
    .A(_18773_),
    .B(_18774_));
 sg13g2_xnor2_1 _27040_ (.Y(_18776_),
    .A(\shift_reg[270] ),
    .B(\shift_reg[271] ));
 sg13g2_xor2_1 _27041_ (.B(\shift_reg[269] ),
    .A(\shift_reg[268] ),
    .X(_18777_));
 sg13g2_xnor2_1 _27042_ (.Y(_18778_),
    .A(_18776_),
    .B(_18777_));
 sg13g2_xnor2_1 _27043_ (.Y(_18779_),
    .A(_18775_),
    .B(_18778_));
 sg13g2_xor2_1 _27044_ (.B(\shift_reg[259] ),
    .A(\shift_reg[258] ),
    .X(_18780_));
 sg13g2_xor2_1 _27045_ (.B(\shift_reg[257] ),
    .A(\shift_reg[256] ),
    .X(_18781_));
 sg13g2_xnor2_1 _27046_ (.Y(_18782_),
    .A(_18780_),
    .B(_18781_));
 sg13g2_xnor2_1 _27047_ (.Y(_18783_),
    .A(\shift_reg[262] ),
    .B(\shift_reg[263] ));
 sg13g2_xor2_1 _27048_ (.B(\shift_reg[261] ),
    .A(\shift_reg[260] ),
    .X(_18784_));
 sg13g2_xnor2_1 _27049_ (.Y(_18785_),
    .A(_18783_),
    .B(_18784_));
 sg13g2_xnor2_1 _27050_ (.Y(_18786_),
    .A(_18782_),
    .B(_18785_));
 sg13g2_xnor2_1 _27051_ (.Y(_18787_),
    .A(_18779_),
    .B(_18786_));
 sg13g2_xnor2_1 _27052_ (.Y(_18788_),
    .A(_18772_),
    .B(_18787_));
 sg13g2_xor2_1 _27053_ (.B(\shift_reg[235] ),
    .A(\shift_reg[234] ),
    .X(_18789_));
 sg13g2_xor2_1 _27054_ (.B(\shift_reg[233] ),
    .A(\shift_reg[232] ),
    .X(_18790_));
 sg13g2_xnor2_1 _27055_ (.Y(_18791_),
    .A(_18789_),
    .B(_18790_));
 sg13g2_xnor2_1 _27056_ (.Y(_18792_),
    .A(\shift_reg[238] ),
    .B(\shift_reg[239] ));
 sg13g2_xor2_1 _27057_ (.B(\shift_reg[237] ),
    .A(\shift_reg[236] ),
    .X(_18793_));
 sg13g2_xnor2_1 _27058_ (.Y(_18794_),
    .A(_18792_),
    .B(_18793_));
 sg13g2_xnor2_1 _27059_ (.Y(_18795_),
    .A(_18791_),
    .B(_18794_));
 sg13g2_xor2_1 _27060_ (.B(\shift_reg[227] ),
    .A(\shift_reg[226] ),
    .X(_18796_));
 sg13g2_xor2_1 _27061_ (.B(\shift_reg[225] ),
    .A(\shift_reg[224] ),
    .X(_18797_));
 sg13g2_xnor2_1 _27062_ (.Y(_18798_),
    .A(_18796_),
    .B(_18797_));
 sg13g2_xnor2_1 _27063_ (.Y(_18799_),
    .A(\shift_reg[230] ),
    .B(\shift_reg[231] ));
 sg13g2_xor2_1 _27064_ (.B(\shift_reg[229] ),
    .A(\shift_reg[228] ),
    .X(_18800_));
 sg13g2_xnor2_1 _27065_ (.Y(_18801_),
    .A(_18799_),
    .B(_18800_));
 sg13g2_xnor2_1 _27066_ (.Y(_18802_),
    .A(_18798_),
    .B(_18801_));
 sg13g2_xnor2_1 _27067_ (.Y(_18803_),
    .A(_18795_),
    .B(_18802_));
 sg13g2_xnor2_1 _27068_ (.Y(_18804_),
    .A(\shift_reg[218] ),
    .B(\shift_reg[219] ));
 sg13g2_xor2_1 _27069_ (.B(\shift_reg[217] ),
    .A(\shift_reg[216] ),
    .X(_18805_));
 sg13g2_xnor2_1 _27070_ (.Y(_18806_),
    .A(_18804_),
    .B(_18805_));
 sg13g2_xnor2_1 _27071_ (.Y(_18807_),
    .A(\shift_reg[222] ),
    .B(\shift_reg[223] ));
 sg13g2_xor2_1 _27072_ (.B(\shift_reg[221] ),
    .A(\shift_reg[220] ),
    .X(_18808_));
 sg13g2_xnor2_1 _27073_ (.Y(_18809_),
    .A(_18807_),
    .B(_18808_));
 sg13g2_xnor2_1 _27074_ (.Y(_18810_),
    .A(_18806_),
    .B(_18809_));
 sg13g2_xor2_1 _27075_ (.B(\shift_reg[211] ),
    .A(\shift_reg[210] ),
    .X(_18811_));
 sg13g2_xor2_1 _27076_ (.B(\shift_reg[209] ),
    .A(\shift_reg[208] ),
    .X(_18812_));
 sg13g2_xnor2_1 _27077_ (.Y(_18813_),
    .A(_18811_),
    .B(_18812_));
 sg13g2_xnor2_1 _27078_ (.Y(_18814_),
    .A(\shift_reg[214] ),
    .B(\shift_reg[215] ));
 sg13g2_xor2_1 _27079_ (.B(\shift_reg[213] ),
    .A(\shift_reg[212] ),
    .X(_18815_));
 sg13g2_xnor2_1 _27080_ (.Y(_18816_),
    .A(_18814_),
    .B(_18815_));
 sg13g2_xnor2_1 _27081_ (.Y(_18817_),
    .A(_18813_),
    .B(_18816_));
 sg13g2_xnor2_1 _27082_ (.Y(_18818_),
    .A(_18810_),
    .B(_18817_));
 sg13g2_xnor2_1 _27083_ (.Y(_18819_),
    .A(_18803_),
    .B(_18818_));
 sg13g2_xnor2_1 _27084_ (.Y(_18820_),
    .A(_18788_),
    .B(_18819_));
 sg13g2_xnor2_1 _27085_ (.Y(_18821_),
    .A(_18757_),
    .B(_18820_));
 sg13g2_xor2_1 _27086_ (.B(\shift_reg[75] ),
    .A(\shift_reg[74] ),
    .X(_18822_));
 sg13g2_xor2_1 _27087_ (.B(\shift_reg[73] ),
    .A(\shift_reg[72] ),
    .X(_18823_));
 sg13g2_xnor2_1 _27088_ (.Y(_18824_),
    .A(_18822_),
    .B(_18823_));
 sg13g2_xnor2_1 _27089_ (.Y(_18825_),
    .A(\shift_reg[78] ),
    .B(\shift_reg[79] ));
 sg13g2_xor2_1 _27090_ (.B(\shift_reg[77] ),
    .A(\shift_reg[76] ),
    .X(_18826_));
 sg13g2_xnor2_1 _27091_ (.Y(_18827_),
    .A(_18825_),
    .B(_18826_));
 sg13g2_xnor2_1 _27092_ (.Y(_18828_),
    .A(_18824_),
    .B(_18827_));
 sg13g2_xor2_1 _27093_ (.B(\shift_reg[187] ),
    .A(\shift_reg[186] ),
    .X(_18829_));
 sg13g2_xor2_1 _27094_ (.B(\shift_reg[185] ),
    .A(\shift_reg[184] ),
    .X(_18830_));
 sg13g2_xnor2_1 _27095_ (.Y(_18831_),
    .A(_18829_),
    .B(_18830_));
 sg13g2_xnor2_1 _27096_ (.Y(_18832_),
    .A(\shift_reg[190] ),
    .B(\shift_reg[191] ));
 sg13g2_xor2_1 _27097_ (.B(\shift_reg[189] ),
    .A(\shift_reg[188] ),
    .X(_18833_));
 sg13g2_xnor2_1 _27098_ (.Y(_18834_),
    .A(_18832_),
    .B(_18833_));
 sg13g2_xnor2_1 _27099_ (.Y(_18835_),
    .A(_18831_),
    .B(_18834_));
 sg13g2_xor2_1 _27100_ (.B(\shift_reg[179] ),
    .A(\shift_reg[178] ),
    .X(_18836_));
 sg13g2_xor2_1 _27101_ (.B(\shift_reg[177] ),
    .A(\shift_reg[176] ),
    .X(_18837_));
 sg13g2_xnor2_1 _27102_ (.Y(_18838_),
    .A(_18836_),
    .B(_18837_));
 sg13g2_xnor2_1 _27103_ (.Y(_18839_),
    .A(\shift_reg[182] ),
    .B(\shift_reg[183] ));
 sg13g2_xor2_1 _27104_ (.B(\shift_reg[181] ),
    .A(\shift_reg[180] ),
    .X(_18840_));
 sg13g2_xnor2_1 _27105_ (.Y(_18841_),
    .A(_18839_),
    .B(_18840_));
 sg13g2_xnor2_1 _27106_ (.Y(_18842_),
    .A(_18838_),
    .B(_18841_));
 sg13g2_xnor2_1 _27107_ (.Y(_18843_),
    .A(_18835_),
    .B(_18842_));
 sg13g2_xor2_1 _27108_ (.B(\shift_reg[203] ),
    .A(\shift_reg[202] ),
    .X(_18844_));
 sg13g2_xor2_1 _27109_ (.B(\shift_reg[201] ),
    .A(\shift_reg[200] ),
    .X(_18845_));
 sg13g2_xnor2_1 _27110_ (.Y(_18846_),
    .A(_18844_),
    .B(_18845_));
 sg13g2_xnor2_1 _27111_ (.Y(_18847_),
    .A(\shift_reg[206] ),
    .B(\shift_reg[207] ));
 sg13g2_xor2_1 _27112_ (.B(\shift_reg[205] ),
    .A(\shift_reg[204] ),
    .X(_18848_));
 sg13g2_xnor2_1 _27113_ (.Y(_18849_),
    .A(_18847_),
    .B(_18848_));
 sg13g2_xnor2_1 _27114_ (.Y(_18850_),
    .A(_18846_),
    .B(_18849_));
 sg13g2_xor2_1 _27115_ (.B(\shift_reg[195] ),
    .A(\shift_reg[194] ),
    .X(_18851_));
 sg13g2_xor2_1 _27116_ (.B(\shift_reg[193] ),
    .A(\shift_reg[192] ),
    .X(_18852_));
 sg13g2_xnor2_1 _27117_ (.Y(_18853_),
    .A(_18851_),
    .B(_18852_));
 sg13g2_xnor2_1 _27118_ (.Y(_18854_),
    .A(\shift_reg[198] ),
    .B(\shift_reg[199] ));
 sg13g2_xor2_1 _27119_ (.B(\shift_reg[197] ),
    .A(\shift_reg[196] ),
    .X(_18855_));
 sg13g2_xnor2_1 _27120_ (.Y(_18856_),
    .A(_18854_),
    .B(_18855_));
 sg13g2_xnor2_1 _27121_ (.Y(_18857_),
    .A(_18853_),
    .B(_18856_));
 sg13g2_xnor2_1 _27122_ (.Y(_18858_),
    .A(_18850_),
    .B(_18857_));
 sg13g2_xnor2_1 _27123_ (.Y(_18859_),
    .A(_18843_),
    .B(_18858_));
 sg13g2_xnor2_1 _27124_ (.Y(_18860_),
    .A(\shift_reg[154] ),
    .B(\shift_reg[155] ));
 sg13g2_xor2_1 _27125_ (.B(\shift_reg[153] ),
    .A(\shift_reg[152] ),
    .X(_18861_));
 sg13g2_xnor2_1 _27126_ (.Y(_18862_),
    .A(_18860_),
    .B(_18861_));
 sg13g2_xnor2_1 _27127_ (.Y(_18863_),
    .A(\shift_reg[158] ),
    .B(\shift_reg[159] ));
 sg13g2_xor2_1 _27128_ (.B(\shift_reg[157] ),
    .A(\shift_reg[156] ),
    .X(_18864_));
 sg13g2_xnor2_1 _27129_ (.Y(_18865_),
    .A(_18863_),
    .B(_18864_));
 sg13g2_xnor2_1 _27130_ (.Y(_18866_),
    .A(_18862_),
    .B(_18865_));
 sg13g2_xor2_1 _27131_ (.B(\shift_reg[147] ),
    .A(\shift_reg[146] ),
    .X(_18867_));
 sg13g2_xor2_1 _27132_ (.B(\shift_reg[145] ),
    .A(\shift_reg[144] ),
    .X(_18868_));
 sg13g2_xnor2_1 _27133_ (.Y(_18869_),
    .A(_18867_),
    .B(_18868_));
 sg13g2_xnor2_1 _27134_ (.Y(_18870_),
    .A(\shift_reg[150] ),
    .B(\shift_reg[151] ));
 sg13g2_xor2_1 _27135_ (.B(\shift_reg[149] ),
    .A(\shift_reg[148] ),
    .X(_18871_));
 sg13g2_xnor2_1 _27136_ (.Y(_18872_),
    .A(_18870_),
    .B(_18871_));
 sg13g2_xnor2_1 _27137_ (.Y(_18873_),
    .A(_18869_),
    .B(_18872_));
 sg13g2_xnor2_1 _27138_ (.Y(_18874_),
    .A(_18866_),
    .B(_18873_));
 sg13g2_xor2_1 _27139_ (.B(\shift_reg[171] ),
    .A(\shift_reg[170] ),
    .X(_18875_));
 sg13g2_xor2_1 _27140_ (.B(\shift_reg[169] ),
    .A(\shift_reg[168] ),
    .X(_18876_));
 sg13g2_xnor2_1 _27141_ (.Y(_18877_),
    .A(_18875_),
    .B(_18876_));
 sg13g2_xnor2_1 _27142_ (.Y(_18878_),
    .A(\shift_reg[174] ),
    .B(\shift_reg[175] ));
 sg13g2_xor2_1 _27143_ (.B(\shift_reg[173] ),
    .A(\shift_reg[172] ),
    .X(_18879_));
 sg13g2_xnor2_1 _27144_ (.Y(_18880_),
    .A(_18878_),
    .B(_18879_));
 sg13g2_xnor2_1 _27145_ (.Y(_18881_),
    .A(_18877_),
    .B(_18880_));
 sg13g2_xor2_1 _27146_ (.B(\shift_reg[163] ),
    .A(\shift_reg[162] ),
    .X(_18882_));
 sg13g2_xor2_1 _27147_ (.B(\shift_reg[161] ),
    .A(\shift_reg[160] ),
    .X(_18883_));
 sg13g2_xnor2_1 _27148_ (.Y(_18884_),
    .A(_18882_),
    .B(_18883_));
 sg13g2_xnor2_1 _27149_ (.Y(_18885_),
    .A(\shift_reg[166] ),
    .B(\shift_reg[167] ));
 sg13g2_xor2_1 _27150_ (.B(\shift_reg[165] ),
    .A(\shift_reg[164] ),
    .X(_18886_));
 sg13g2_xnor2_1 _27151_ (.Y(_18887_),
    .A(_18885_),
    .B(_18886_));
 sg13g2_xnor2_1 _27152_ (.Y(_18888_),
    .A(_18884_),
    .B(_18887_));
 sg13g2_xnor2_1 _27153_ (.Y(_18889_),
    .A(_18881_),
    .B(_18888_));
 sg13g2_xnor2_1 _27154_ (.Y(_18890_),
    .A(_18874_),
    .B(_18889_));
 sg13g2_xnor2_1 _27155_ (.Y(_18891_),
    .A(_18859_),
    .B(_18890_));
 sg13g2_xnor2_1 _27156_ (.Y(_18892_),
    .A(_18725_),
    .B(_18828_));
 sg13g2_xnor2_1 _27157_ (.Y(_18893_),
    .A(_18718_),
    .B(_18892_));
 sg13g2_xnor2_1 _27158_ (.Y(_18894_),
    .A(_18703_),
    .B(_18893_));
 sg13g2_xnor2_1 _27159_ (.Y(_18895_),
    .A(_18891_),
    .B(_18894_));
 sg13g2_xnor2_1 _27160_ (.Y(_18896_),
    .A(_18821_),
    .B(_18895_));
 sg13g2_a21oi_1 _27161_ (.A1(net1159),
    .A2(_18896_),
    .Y(_00163_),
    .B1(_18640_));
 sg13g2_xnor2_1 _27162_ (.Y(_00164_),
    .A(net1173),
    .B(net6677));
 sg13g2_a21o_1 _27163_ (.A2(_18633_),
    .A1(net1173),
    .B1(net1222),
    .X(_18897_));
 sg13g2_and2_1 _27164_ (.A(_18634_),
    .B(_18897_),
    .X(_00165_));
 sg13g2_xnor2_1 _27165_ (.Y(_00166_),
    .A(net1151),
    .B(_18634_));
 sg13g2_nor2_1 _27166_ (.A(net3668),
    .B(_18625_),
    .Y(_18898_));
 sg13g2_inv_1 _27167_ (.Y(_18899_),
    .A(_18898_));
 sg13g2_nand3_1 _27168_ (.B(uio_out[1]),
    .C(_18618_),
    .A(net1678),
    .Y(_18900_));
 sg13g2_nand2b_1 _27169_ (.Y(_18901_),
    .B(net2976),
    .A_N(uio_out[1]));
 sg13g2_nor2_2 _27170_ (.A(net7412),
    .B(_18619_),
    .Y(_18902_));
 sg13g2_nand2_1 _27171_ (.Y(_18903_),
    .A(inv_done),
    .B(_18624_));
 sg13g2_nor2_1 _27172_ (.A(uio_out[1]),
    .B(net6945),
    .Y(_18904_));
 sg13g2_and3_1 _27173_ (.X(_18905_),
    .A(_18900_),
    .B(_18901_),
    .C(net6901));
 sg13g2_or2_1 _27174_ (.X(_18906_),
    .B(_18905_),
    .A(net7413));
 sg13g2_nor2_2 _27175_ (.A(net7413),
    .B(_18618_),
    .Y(_18907_));
 sg13g2_a221oi_1 _27176_ (.B2(_18906_),
    .C1(_18907_),
    .B1(_18899_),
    .A1(_18615_),
    .Y(_00167_),
    .A2(_18617_));
 sg13g2_a21oi_2 _27177_ (.B1(net6945),
    .Y(_18908_),
    .A2(_18907_),
    .A1(net3755));
 sg13g2_inv_1 _27178_ (.Y(_00168_),
    .A(net6676));
 sg13g2_nor2b_1 _27179_ (.A(net1179),
    .B_N(_18618_),
    .Y(_18909_));
 sg13g2_nor2_1 _27180_ (.A(inv_done),
    .B(_18909_),
    .Y(_18910_));
 sg13g2_o21ai_1 _27181_ (.B1(net7413),
    .Y(_18911_),
    .A1(net7412),
    .A2(_18910_));
 sg13g2_nor2b_2 _27182_ (.A(_18907_),
    .B_N(_18911_),
    .Y(_18912_));
 sg13g2_inv_1 _27183_ (.Y(_18913_),
    .A(_18912_));
 sg13g2_mux2_1 _27184_ (.A0(net2976),
    .A1(_18905_),
    .S(_18912_),
    .X(_00169_));
 sg13g2_and3_1 _27185_ (.X(_18914_),
    .A(net3769),
    .B(net1166),
    .C(_18912_));
 sg13g2_nor2_1 _27186_ (.A(_18904_),
    .B(_18913_),
    .Y(_18915_));
 sg13g2_inv_1 _27187_ (.Y(_18916_),
    .A(_18915_));
 sg13g2_a21oi_1 _27188_ (.A1(_18617_),
    .A2(_18904_),
    .Y(_18917_),
    .B1(_18913_));
 sg13g2_a21oi_1 _27189_ (.A1(\byte_cnt[0] ),
    .A2(_18912_),
    .Y(_18918_),
    .B1(net1166));
 sg13g2_nor3_1 _27190_ (.A(_18914_),
    .B(_18917_),
    .C(net1167),
    .Y(_00170_));
 sg13g2_nor2_1 _27191_ (.A(net1840),
    .B(_18914_),
    .Y(_18919_));
 sg13g2_and2_1 _27192_ (.A(net1840),
    .B(_18914_),
    .X(_18920_));
 sg13g2_nor3_1 _27193_ (.A(_18915_),
    .B(net1841),
    .C(_18920_),
    .Y(_00171_));
 sg13g2_a22oi_1 _27194_ (.Y(_18921_),
    .B1(_18920_),
    .B2(_18904_),
    .A2(_18916_),
    .A1(net1153));
 sg13g2_a21oi_1 _27195_ (.A1(net1153),
    .A2(_18920_),
    .Y(_00172_),
    .B1(_18921_));
 sg13g2_a21oi_1 _27196_ (.A1(net1153),
    .A2(_18920_),
    .Y(_18922_),
    .B1(net1174));
 sg13g2_nand3_1 _27197_ (.B(net1174),
    .C(_18920_),
    .A(net1153),
    .Y(_18923_));
 sg13g2_nand2_1 _27198_ (.Y(_18924_),
    .A(_18916_),
    .B(_18923_));
 sg13g2_nor2_1 _27199_ (.A(net1175),
    .B(_18924_),
    .Y(_00173_));
 sg13g2_xor2_1 _27200_ (.B(_18923_),
    .A(net2486),
    .X(_18925_));
 sg13g2_nor2_1 _27201_ (.A(_18917_),
    .B(_18925_),
    .Y(_00174_));
 sg13g2_o21ai_1 _27202_ (.B1(net7412),
    .Y(_18926_),
    .A1(_18257_),
    .A2(net12));
 sg13g2_o21ai_1 _27203_ (.B1(_18907_),
    .Y(_18927_),
    .A1(_18635_),
    .A2(_18926_));
 sg13g2_and3_2 _27204_ (.X(_18928_),
    .A(_18900_),
    .B(_18911_),
    .C(_18927_));
 sg13g2_nand3_1 _27205_ (.B(net6676),
    .C(net6529),
    .A(net2),
    .Y(_18929_));
 sg13g2_o21ai_1 _27206_ (.B1(_18929_),
    .Y(_00175_),
    .A1(_18258_),
    .A2(net6530));
 sg13g2_nand3_1 _27207_ (.B(net6676),
    .C(net6529),
    .A(net3),
    .Y(_18930_));
 sg13g2_o21ai_1 _27208_ (.B1(_18930_),
    .Y(_00176_),
    .A1(_18259_),
    .A2(net6532));
 sg13g2_nand3_1 _27209_ (.B(net6676),
    .C(net6529),
    .A(net4),
    .Y(_18931_));
 sg13g2_o21ai_1 _27210_ (.B1(_18931_),
    .Y(_00177_),
    .A1(_18260_),
    .A2(net6530));
 sg13g2_nand3_1 _27211_ (.B(net6676),
    .C(net6529),
    .A(net5),
    .Y(_18932_));
 sg13g2_o21ai_1 _27212_ (.B1(_18932_),
    .Y(_00178_),
    .A1(_18261_),
    .A2(net6532));
 sg13g2_nand3_1 _27213_ (.B(net6676),
    .C(net6529),
    .A(net6),
    .Y(_18933_));
 sg13g2_o21ai_1 _27214_ (.B1(_18933_),
    .Y(_00179_),
    .A1(_18262_),
    .A2(net6530));
 sg13g2_nand3_1 _27215_ (.B(_18908_),
    .C(net6529),
    .A(net7),
    .Y(_18934_));
 sg13g2_o21ai_1 _27216_ (.B1(_18934_),
    .Y(_00180_),
    .A1(_18263_),
    .A2(net6530));
 sg13g2_nand3_1 _27217_ (.B(net6676),
    .C(net6529),
    .A(net8),
    .Y(_18935_));
 sg13g2_o21ai_1 _27218_ (.B1(_18935_),
    .Y(_00181_),
    .A1(_18264_),
    .A2(net6530));
 sg13g2_nand3_1 _27219_ (.B(net6676),
    .C(net6529),
    .A(net9),
    .Y(_18936_));
 sg13g2_o21ai_1 _27220_ (.B1(_18936_),
    .Y(_00182_),
    .A1(_18266_),
    .A2(net6555));
 sg13g2_nand3_1 _27221_ (.B(net6903),
    .C(net6532),
    .A(\shift_reg[0] ),
    .Y(_18937_));
 sg13g2_o21ai_1 _27222_ (.B1(_18937_),
    .Y(_00183_),
    .A1(_18333_),
    .A2(net6517));
 sg13g2_nand3_1 _27223_ (.B(net6908),
    .C(net6542),
    .A(\shift_reg[1] ),
    .Y(_18938_));
 sg13g2_o21ai_1 _27224_ (.B1(_18938_),
    .Y(_00184_),
    .A1(_18334_),
    .A2(net6535));
 sg13g2_nand3_1 _27225_ (.B(net6903),
    .C(net6532),
    .A(net1521),
    .Y(_18939_));
 sg13g2_o21ai_1 _27226_ (.B1(_18939_),
    .Y(_00185_),
    .A1(_18335_),
    .A2(net6516));
 sg13g2_nand3_1 _27227_ (.B(net6903),
    .C(net6532),
    .A(net1574),
    .Y(_18940_));
 sg13g2_o21ai_1 _27228_ (.B1(_18940_),
    .Y(_00186_),
    .A1(_18336_),
    .A2(net6534));
 sg13g2_nand3_1 _27229_ (.B(net6893),
    .C(net6517),
    .A(\shift_reg[4] ),
    .Y(_18941_));
 sg13g2_o21ai_1 _27230_ (.B1(_18941_),
    .Y(_00187_),
    .A1(_18337_),
    .A2(net6515));
 sg13g2_nand3_1 _27231_ (.B(net6894),
    .C(net6518),
    .A(\shift_reg[5] ),
    .Y(_18942_));
 sg13g2_o21ai_1 _27232_ (.B1(_18942_),
    .Y(_00188_),
    .A1(_18338_),
    .A2(net6537));
 sg13g2_nor2b_2 _27233_ (.A(net13),
    .B_N(net12),
    .Y(_18943_));
 sg13g2_nand2_1 _27234_ (.Y(_18944_),
    .A(_18257_),
    .B(net12));
 sg13g2_nor2_2 _27235_ (.A(net6899),
    .B(_18943_),
    .Y(_18945_));
 sg13g2_a22oi_1 _27236_ (.Y(_18946_),
    .B1(net6637),
    .B2(parity_error),
    .A2(net6893),
    .A1(\shift_reg[6] ));
 sg13g2_nor2_1 _27237_ (.A(net2828),
    .B(net6519),
    .Y(_18947_));
 sg13g2_a21oi_1 _27238_ (.A1(net6519),
    .A2(_18946_),
    .Y(_00189_),
    .B1(_18947_));
 sg13g2_xor2_1 _27239_ (.B(\inv_result[102] ),
    .A(\inv_result[103] ),
    .X(_18948_));
 sg13g2_xor2_1 _27240_ (.B(\inv_result[96] ),
    .A(\inv_result[97] ),
    .X(_18949_));
 sg13g2_xnor2_1 _27241_ (.Y(_18950_),
    .A(_18948_),
    .B(_18949_));
 sg13g2_xnor2_1 _27242_ (.Y(_18951_),
    .A(\inv_result[101] ),
    .B(\inv_result[100] ));
 sg13g2_xor2_1 _27243_ (.B(\inv_result[98] ),
    .A(\inv_result[99] ),
    .X(_18952_));
 sg13g2_xnor2_1 _27244_ (.Y(_18953_),
    .A(_18951_),
    .B(_18952_));
 sg13g2_xnor2_1 _27245_ (.Y(_18954_),
    .A(_18950_),
    .B(_18953_));
 sg13g2_xor2_1 _27246_ (.B(\inv_result[110] ),
    .A(\inv_result[111] ),
    .X(_18955_));
 sg13g2_xor2_1 _27247_ (.B(\inv_result[104] ),
    .A(\inv_result[105] ),
    .X(_18956_));
 sg13g2_xnor2_1 _27248_ (.Y(_18957_),
    .A(_18955_),
    .B(_18956_));
 sg13g2_xnor2_1 _27249_ (.Y(_18958_),
    .A(\inv_result[109] ),
    .B(\inv_result[108] ));
 sg13g2_xor2_1 _27250_ (.B(\inv_result[106] ),
    .A(\inv_result[107] ),
    .X(_18959_));
 sg13g2_xnor2_1 _27251_ (.Y(_18960_),
    .A(_18958_),
    .B(_18959_));
 sg13g2_xnor2_1 _27252_ (.Y(_18961_),
    .A(_18957_),
    .B(_18960_));
 sg13g2_xnor2_1 _27253_ (.Y(_18962_),
    .A(_18954_),
    .B(_18961_));
 sg13g2_xor2_1 _27254_ (.B(\inv_result[66] ),
    .A(\inv_result[67] ),
    .X(_18963_));
 sg13g2_xor2_1 _27255_ (.B(\inv_result[64] ),
    .A(\inv_result[65] ),
    .X(_18964_));
 sg13g2_xnor2_1 _27256_ (.Y(_18965_),
    .A(_18963_),
    .B(_18964_));
 sg13g2_xnor2_1 _27257_ (.Y(_18966_),
    .A(\inv_result[71] ),
    .B(\inv_result[70] ));
 sg13g2_xor2_1 _27258_ (.B(\inv_result[68] ),
    .A(\inv_result[69] ),
    .X(_18967_));
 sg13g2_xnor2_1 _27259_ (.Y(_18968_),
    .A(_18966_),
    .B(_18967_));
 sg13g2_xnor2_1 _27260_ (.Y(_18969_),
    .A(_18965_),
    .B(_18968_));
 sg13g2_xor2_1 _27261_ (.B(\inv_result[78] ),
    .A(\inv_result[79] ),
    .X(_18970_));
 sg13g2_xor2_1 _27262_ (.B(\inv_result[72] ),
    .A(\inv_result[73] ),
    .X(_18971_));
 sg13g2_xnor2_1 _27263_ (.Y(_18972_),
    .A(_18970_),
    .B(_18971_));
 sg13g2_xnor2_1 _27264_ (.Y(_18973_),
    .A(\inv_result[77] ),
    .B(\inv_result[76] ));
 sg13g2_xor2_1 _27265_ (.B(\inv_result[74] ),
    .A(\inv_result[75] ),
    .X(_18974_));
 sg13g2_xnor2_1 _27266_ (.Y(_18975_),
    .A(_18973_),
    .B(_18974_));
 sg13g2_xnor2_1 _27267_ (.Y(_18976_),
    .A(_18972_),
    .B(_18975_));
 sg13g2_xnor2_1 _27268_ (.Y(_18977_),
    .A(_18969_),
    .B(_18976_));
 sg13g2_xnor2_1 _27269_ (.Y(_18978_),
    .A(_18962_),
    .B(_18977_));
 sg13g2_xor2_1 _27270_ (.B(\inv_result[6] ),
    .A(\inv_result[7] ),
    .X(_18979_));
 sg13g2_xor2_1 _27271_ (.B(\inv_result[0] ),
    .A(\inv_result[1] ),
    .X(_18980_));
 sg13g2_xnor2_1 _27272_ (.Y(_18981_),
    .A(_18979_),
    .B(_18980_));
 sg13g2_xnor2_1 _27273_ (.Y(_18982_),
    .A(\inv_result[5] ),
    .B(\inv_result[4] ));
 sg13g2_xor2_1 _27274_ (.B(\inv_result[2] ),
    .A(\inv_result[3] ),
    .X(_18983_));
 sg13g2_xnor2_1 _27275_ (.Y(_18984_),
    .A(_18982_),
    .B(_18983_));
 sg13g2_xnor2_1 _27276_ (.Y(_18985_),
    .A(_18981_),
    .B(_18984_));
 sg13g2_xor2_1 _27277_ (.B(\inv_result[10] ),
    .A(\inv_result[11] ),
    .X(_18986_));
 sg13g2_xor2_1 _27278_ (.B(\inv_result[8] ),
    .A(\inv_result[9] ),
    .X(_18987_));
 sg13g2_xnor2_1 _27279_ (.Y(_18988_),
    .A(_18986_),
    .B(_18987_));
 sg13g2_xnor2_1 _27280_ (.Y(_18989_),
    .A(\inv_result[15] ),
    .B(\inv_result[14] ));
 sg13g2_xor2_1 _27281_ (.B(\inv_result[12] ),
    .A(\inv_result[13] ),
    .X(_18990_));
 sg13g2_xnor2_1 _27282_ (.Y(_18991_),
    .A(_18989_),
    .B(_18990_));
 sg13g2_xnor2_1 _27283_ (.Y(_18992_),
    .A(_18988_),
    .B(_18991_));
 sg13g2_xnor2_1 _27284_ (.Y(_18993_),
    .A(_18985_),
    .B(_18992_));
 sg13g2_xor2_1 _27285_ (.B(\inv_result[42] ),
    .A(\inv_result[43] ),
    .X(_18994_));
 sg13g2_xor2_1 _27286_ (.B(\inv_result[40] ),
    .A(\inv_result[41] ),
    .X(_18995_));
 sg13g2_xnor2_1 _27287_ (.Y(_18996_),
    .A(_18994_),
    .B(_18995_));
 sg13g2_xnor2_1 _27288_ (.Y(_18997_),
    .A(\inv_result[47] ),
    .B(\inv_result[46] ));
 sg13g2_xor2_1 _27289_ (.B(\inv_result[44] ),
    .A(\inv_result[45] ),
    .X(_18998_));
 sg13g2_xnor2_1 _27290_ (.Y(_18999_),
    .A(_18997_),
    .B(_18998_));
 sg13g2_xnor2_1 _27291_ (.Y(_19000_),
    .A(_18996_),
    .B(_18999_));
 sg13g2_xor2_1 _27292_ (.B(\inv_result[34] ),
    .A(\inv_result[35] ),
    .X(_19001_));
 sg13g2_xor2_1 _27293_ (.B(\inv_result[32] ),
    .A(\inv_result[33] ),
    .X(_19002_));
 sg13g2_xnor2_1 _27294_ (.Y(_19003_),
    .A(_19001_),
    .B(_19002_));
 sg13g2_xnor2_1 _27295_ (.Y(_19004_),
    .A(\inv_result[39] ),
    .B(\inv_result[38] ));
 sg13g2_xor2_1 _27296_ (.B(\inv_result[36] ),
    .A(\inv_result[37] ),
    .X(_19005_));
 sg13g2_xnor2_1 _27297_ (.Y(_19006_),
    .A(_19004_),
    .B(_19005_));
 sg13g2_xnor2_1 _27298_ (.Y(_19007_),
    .A(_19003_),
    .B(_19006_));
 sg13g2_xnor2_1 _27299_ (.Y(_19008_),
    .A(_19000_),
    .B(_19007_));
 sg13g2_xnor2_1 _27300_ (.Y(_19009_),
    .A(_18993_),
    .B(_19008_));
 sg13g2_xor2_1 _27301_ (.B(\inv_result[90] ),
    .A(\inv_result[91] ),
    .X(_19010_));
 sg13g2_xor2_1 _27302_ (.B(\inv_result[88] ),
    .A(\inv_result[89] ),
    .X(_19011_));
 sg13g2_xnor2_1 _27303_ (.Y(_19012_),
    .A(_19010_),
    .B(_19011_));
 sg13g2_xnor2_1 _27304_ (.Y(_19013_),
    .A(\inv_result[95] ),
    .B(\inv_result[94] ));
 sg13g2_xor2_1 _27305_ (.B(\inv_result[92] ),
    .A(\inv_result[93] ),
    .X(_19014_));
 sg13g2_xnor2_1 _27306_ (.Y(_19015_),
    .A(_19013_),
    .B(_19014_));
 sg13g2_xnor2_1 _27307_ (.Y(_19016_),
    .A(_19012_),
    .B(_19015_));
 sg13g2_xor2_1 _27308_ (.B(\inv_result[82] ),
    .A(\inv_result[83] ),
    .X(_19017_));
 sg13g2_xor2_1 _27309_ (.B(\inv_result[80] ),
    .A(\inv_result[81] ),
    .X(_19018_));
 sg13g2_xnor2_1 _27310_ (.Y(_19019_),
    .A(_19017_),
    .B(_19018_));
 sg13g2_xnor2_1 _27311_ (.Y(_19020_),
    .A(\inv_result[87] ),
    .B(\inv_result[86] ));
 sg13g2_xor2_1 _27312_ (.B(\inv_result[84] ),
    .A(\inv_result[85] ),
    .X(_19021_));
 sg13g2_xnor2_1 _27313_ (.Y(_19022_),
    .A(_19020_),
    .B(_19021_));
 sg13g2_xnor2_1 _27314_ (.Y(_19023_),
    .A(_19019_),
    .B(_19022_));
 sg13g2_xnor2_1 _27315_ (.Y(_19024_),
    .A(_19016_),
    .B(_19023_));
 sg13g2_xor2_1 _27316_ (.B(\inv_result[122] ),
    .A(\inv_result[123] ),
    .X(_19025_));
 sg13g2_xor2_1 _27317_ (.B(\inv_result[120] ),
    .A(\inv_result[121] ),
    .X(_19026_));
 sg13g2_xnor2_1 _27318_ (.Y(_19027_),
    .A(_19025_),
    .B(_19026_));
 sg13g2_xnor2_1 _27319_ (.Y(_19028_),
    .A(\inv_result[127] ),
    .B(\inv_result[126] ));
 sg13g2_xor2_1 _27320_ (.B(\inv_result[124] ),
    .A(\inv_result[125] ),
    .X(_19029_));
 sg13g2_xnor2_1 _27321_ (.Y(_19030_),
    .A(_19028_),
    .B(_19029_));
 sg13g2_xnor2_1 _27322_ (.Y(_19031_),
    .A(_19027_),
    .B(_19030_));
 sg13g2_xor2_1 _27323_ (.B(\inv_result[114] ),
    .A(\inv_result[115] ),
    .X(_19032_));
 sg13g2_xor2_1 _27324_ (.B(\inv_result[112] ),
    .A(\inv_result[113] ),
    .X(_19033_));
 sg13g2_xnor2_1 _27325_ (.Y(_19034_),
    .A(_19032_),
    .B(_19033_));
 sg13g2_xnor2_1 _27326_ (.Y(_19035_),
    .A(\inv_result[119] ),
    .B(\inv_result[118] ));
 sg13g2_xor2_1 _27327_ (.B(\inv_result[116] ),
    .A(\inv_result[117] ),
    .X(_19036_));
 sg13g2_xnor2_1 _27328_ (.Y(_19037_),
    .A(_19035_),
    .B(_19036_));
 sg13g2_xnor2_1 _27329_ (.Y(_19038_),
    .A(_19034_),
    .B(_19037_));
 sg13g2_xnor2_1 _27330_ (.Y(_19039_),
    .A(_19031_),
    .B(_19038_));
 sg13g2_xnor2_1 _27331_ (.Y(_19040_),
    .A(_19024_),
    .B(_19039_));
 sg13g2_xor2_1 _27332_ (.B(\inv_result[62] ),
    .A(\inv_result[63] ),
    .X(_19041_));
 sg13g2_xor2_1 _27333_ (.B(\inv_result[56] ),
    .A(\inv_result[57] ),
    .X(_19042_));
 sg13g2_xnor2_1 _27334_ (.Y(_19043_),
    .A(_19041_),
    .B(_19042_));
 sg13g2_xnor2_1 _27335_ (.Y(_19044_),
    .A(\inv_result[61] ),
    .B(\inv_result[60] ));
 sg13g2_xor2_1 _27336_ (.B(\inv_result[58] ),
    .A(\inv_result[59] ),
    .X(_19045_));
 sg13g2_xnor2_1 _27337_ (.Y(_19046_),
    .A(_19044_),
    .B(_19045_));
 sg13g2_xnor2_1 _27338_ (.Y(_19047_),
    .A(_19043_),
    .B(_19046_));
 sg13g2_xor2_1 _27339_ (.B(\inv_result[54] ),
    .A(\inv_result[55] ),
    .X(_19048_));
 sg13g2_xor2_1 _27340_ (.B(\inv_result[48] ),
    .A(\inv_result[49] ),
    .X(_19049_));
 sg13g2_xnor2_1 _27341_ (.Y(_19050_),
    .A(_19048_),
    .B(_19049_));
 sg13g2_xnor2_1 _27342_ (.Y(_19051_),
    .A(\inv_result[53] ),
    .B(\inv_result[52] ));
 sg13g2_xor2_1 _27343_ (.B(\inv_result[50] ),
    .A(\inv_result[51] ),
    .X(_19052_));
 sg13g2_xnor2_1 _27344_ (.Y(_19053_),
    .A(_19051_),
    .B(_19052_));
 sg13g2_xnor2_1 _27345_ (.Y(_19054_),
    .A(_19050_),
    .B(_19053_));
 sg13g2_xnor2_1 _27346_ (.Y(_19055_),
    .A(_19047_),
    .B(_19054_));
 sg13g2_xor2_1 _27347_ (.B(\inv_result[26] ),
    .A(\inv_result[27] ),
    .X(_19056_));
 sg13g2_xor2_1 _27348_ (.B(\inv_result[24] ),
    .A(\inv_result[25] ),
    .X(_19057_));
 sg13g2_xnor2_1 _27349_ (.Y(_19058_),
    .A(_19056_),
    .B(_19057_));
 sg13g2_xnor2_1 _27350_ (.Y(_19059_),
    .A(\inv_result[31] ),
    .B(\inv_result[30] ));
 sg13g2_xor2_1 _27351_ (.B(\inv_result[28] ),
    .A(\inv_result[29] ),
    .X(_19060_));
 sg13g2_xnor2_1 _27352_ (.Y(_19061_),
    .A(_19059_),
    .B(_19060_));
 sg13g2_xnor2_1 _27353_ (.Y(_19062_),
    .A(_19058_),
    .B(_19061_));
 sg13g2_xor2_1 _27354_ (.B(\inv_result[18] ),
    .A(\inv_result[19] ),
    .X(_19063_));
 sg13g2_xor2_1 _27355_ (.B(\inv_result[16] ),
    .A(\inv_result[17] ),
    .X(_19064_));
 sg13g2_xnor2_1 _27356_ (.Y(_19065_),
    .A(_19063_),
    .B(_19064_));
 sg13g2_xnor2_1 _27357_ (.Y(_19066_),
    .A(\inv_result[23] ),
    .B(\inv_result[22] ));
 sg13g2_xor2_1 _27358_ (.B(\inv_result[20] ),
    .A(\inv_result[21] ),
    .X(_19067_));
 sg13g2_xnor2_1 _27359_ (.Y(_19068_),
    .A(_19066_),
    .B(_19067_));
 sg13g2_xnor2_1 _27360_ (.Y(_19069_),
    .A(_19065_),
    .B(_19068_));
 sg13g2_xnor2_1 _27361_ (.Y(_19070_),
    .A(_19062_),
    .B(_19069_));
 sg13g2_xnor2_1 _27362_ (.Y(_19071_),
    .A(_19055_),
    .B(_19070_));
 sg13g2_xnor2_1 _27363_ (.Y(_19072_),
    .A(_18978_),
    .B(_19040_));
 sg13g2_xnor2_1 _27364_ (.Y(_19073_),
    .A(_19009_),
    .B(_19071_));
 sg13g2_xnor2_1 _27365_ (.Y(_19074_),
    .A(_19072_),
    .B(_19073_));
 sg13g2_xor2_1 _27366_ (.B(\inv_result[158] ),
    .A(\inv_result[159] ),
    .X(_19075_));
 sg13g2_xor2_1 _27367_ (.B(\inv_result[152] ),
    .A(\inv_result[153] ),
    .X(_19076_));
 sg13g2_xnor2_1 _27368_ (.Y(_19077_),
    .A(_19075_),
    .B(_19076_));
 sg13g2_xnor2_1 _27369_ (.Y(_19078_),
    .A(\inv_result[157] ),
    .B(\inv_result[156] ));
 sg13g2_xor2_1 _27370_ (.B(\inv_result[154] ),
    .A(\inv_result[155] ),
    .X(_19079_));
 sg13g2_xnor2_1 _27371_ (.Y(_19080_),
    .A(_19078_),
    .B(_19079_));
 sg13g2_xnor2_1 _27372_ (.Y(_19081_),
    .A(_19077_),
    .B(_19080_));
 sg13g2_xor2_1 _27373_ (.B(\inv_result[146] ),
    .A(\inv_result[147] ),
    .X(_19082_));
 sg13g2_xor2_1 _27374_ (.B(\inv_result[144] ),
    .A(\inv_result[145] ),
    .X(_19083_));
 sg13g2_xnor2_1 _27375_ (.Y(_19084_),
    .A(_19082_),
    .B(_19083_));
 sg13g2_xnor2_1 _27376_ (.Y(_19085_),
    .A(\inv_result[151] ),
    .B(\inv_result[150] ));
 sg13g2_xor2_1 _27377_ (.B(\inv_result[148] ),
    .A(\inv_result[149] ),
    .X(_19086_));
 sg13g2_xnor2_1 _27378_ (.Y(_19087_),
    .A(_19085_),
    .B(_19086_));
 sg13g2_xnor2_1 _27379_ (.Y(_19088_),
    .A(_19084_),
    .B(_19087_));
 sg13g2_xnor2_1 _27380_ (.Y(_19089_),
    .A(_19081_),
    .B(_19088_));
 sg13g2_xor2_1 _27381_ (.B(\inv_result[250] ),
    .A(\inv_result[251] ),
    .X(_19090_));
 sg13g2_xor2_1 _27382_ (.B(\inv_result[248] ),
    .A(\inv_result[249] ),
    .X(_19091_));
 sg13g2_xnor2_1 _27383_ (.Y(_19092_),
    .A(_19090_),
    .B(_19091_));
 sg13g2_xnor2_1 _27384_ (.Y(_19093_),
    .A(\inv_result[255] ),
    .B(\inv_result[254] ));
 sg13g2_xor2_1 _27385_ (.B(\inv_result[252] ),
    .A(\inv_result[253] ),
    .X(_19094_));
 sg13g2_xnor2_1 _27386_ (.Y(_19095_),
    .A(_19093_),
    .B(_19094_));
 sg13g2_xnor2_1 _27387_ (.Y(_19096_),
    .A(_19092_),
    .B(_19095_));
 sg13g2_xor2_1 _27388_ (.B(\inv_result[242] ),
    .A(\inv_result[243] ),
    .X(_19097_));
 sg13g2_xor2_1 _27389_ (.B(\inv_result[240] ),
    .A(\inv_result[241] ),
    .X(_19098_));
 sg13g2_xnor2_1 _27390_ (.Y(_19099_),
    .A(_19097_),
    .B(_19098_));
 sg13g2_xnor2_1 _27391_ (.Y(_19100_),
    .A(\inv_result[247] ),
    .B(\inv_result[246] ));
 sg13g2_xor2_1 _27392_ (.B(\inv_result[244] ),
    .A(\inv_result[245] ),
    .X(_19101_));
 sg13g2_xnor2_1 _27393_ (.Y(_19102_),
    .A(_19100_),
    .B(_19101_));
 sg13g2_xnor2_1 _27394_ (.Y(_19103_),
    .A(_19099_),
    .B(_19102_));
 sg13g2_xnor2_1 _27395_ (.Y(_19104_),
    .A(_19096_),
    .B(_19103_));
 sg13g2_xnor2_1 _27396_ (.Y(_19105_),
    .A(_19089_),
    .B(_19104_));
 sg13g2_xor2_1 _27397_ (.B(\inv_result[226] ),
    .A(\inv_result[227] ),
    .X(_19106_));
 sg13g2_xor2_1 _27398_ (.B(\inv_result[224] ),
    .A(\inv_result[225] ),
    .X(_19107_));
 sg13g2_xnor2_1 _27399_ (.Y(_19108_),
    .A(_19106_),
    .B(_19107_));
 sg13g2_xnor2_1 _27400_ (.Y(_19109_),
    .A(\inv_result[231] ),
    .B(\inv_result[230] ));
 sg13g2_xor2_1 _27401_ (.B(\inv_result[228] ),
    .A(\inv_result[229] ),
    .X(_19110_));
 sg13g2_xnor2_1 _27402_ (.Y(_19111_),
    .A(_19109_),
    .B(_19110_));
 sg13g2_xnor2_1 _27403_ (.Y(_19112_),
    .A(_19108_),
    .B(_19111_));
 sg13g2_xnor2_1 _27404_ (.Y(_19113_),
    .A(\inv_result[139] ),
    .B(\inv_result[138] ));
 sg13g2_xor2_1 _27405_ (.B(\inv_result[136] ),
    .A(\inv_result[137] ),
    .X(_19114_));
 sg13g2_xnor2_1 _27406_ (.Y(_19115_),
    .A(_19113_),
    .B(_19114_));
 sg13g2_xnor2_1 _27407_ (.Y(_19116_),
    .A(\inv_result[143] ),
    .B(\inv_result[142] ));
 sg13g2_xor2_1 _27408_ (.B(\inv_result[140] ),
    .A(\inv_result[141] ),
    .X(_19117_));
 sg13g2_xnor2_1 _27409_ (.Y(_19118_),
    .A(_19116_),
    .B(_19117_));
 sg13g2_xnor2_1 _27410_ (.Y(_19119_),
    .A(_19115_),
    .B(_19118_));
 sg13g2_xnor2_1 _27411_ (.Y(_19120_),
    .A(\inv_result[239] ),
    .B(\inv_result[238] ));
 sg13g2_xor2_1 _27412_ (.B(\inv_result[232] ),
    .A(\inv_result[233] ),
    .X(_19121_));
 sg13g2_xnor2_1 _27413_ (.Y(_19122_),
    .A(_19120_),
    .B(_19121_));
 sg13g2_xnor2_1 _27414_ (.Y(_19123_),
    .A(\inv_result[237] ),
    .B(\inv_result[236] ));
 sg13g2_xor2_1 _27415_ (.B(\inv_result[234] ),
    .A(\inv_result[235] ),
    .X(_19124_));
 sg13g2_xnor2_1 _27416_ (.Y(_19125_),
    .A(_19123_),
    .B(_19124_));
 sg13g2_xnor2_1 _27417_ (.Y(_19126_),
    .A(_19122_),
    .B(_19125_));
 sg13g2_xnor2_1 _27418_ (.Y(_19127_),
    .A(\inv_result[135] ),
    .B(\inv_result[134] ));
 sg13g2_xor2_1 _27419_ (.B(\inv_result[128] ),
    .A(\inv_result[129] ),
    .X(_19128_));
 sg13g2_xnor2_1 _27420_ (.Y(_19129_),
    .A(_19127_),
    .B(_19128_));
 sg13g2_xnor2_1 _27421_ (.Y(_19130_),
    .A(\inv_result[133] ),
    .B(\inv_result[132] ));
 sg13g2_xor2_1 _27422_ (.B(\inv_result[130] ),
    .A(\inv_result[131] ),
    .X(_19131_));
 sg13g2_xnor2_1 _27423_ (.Y(_19132_),
    .A(_19130_),
    .B(_19131_));
 sg13g2_xnor2_1 _27424_ (.Y(_19133_),
    .A(_19129_),
    .B(_19132_));
 sg13g2_xnor2_1 _27425_ (.Y(_19134_),
    .A(_19112_),
    .B(_19126_));
 sg13g2_xnor2_1 _27426_ (.Y(_19135_),
    .A(_19119_),
    .B(_19133_));
 sg13g2_xnor2_1 _27427_ (.Y(_19136_),
    .A(_19134_),
    .B(_19135_));
 sg13g2_xnor2_1 _27428_ (.Y(_19137_),
    .A(_19105_),
    .B(_19136_));
 sg13g2_xor2_1 _27429_ (.B(\inv_result[170] ),
    .A(\inv_result[171] ),
    .X(_19138_));
 sg13g2_xor2_1 _27430_ (.B(\inv_result[168] ),
    .A(\inv_result[169] ),
    .X(_19139_));
 sg13g2_xnor2_1 _27431_ (.Y(_19140_),
    .A(_19138_),
    .B(_19139_));
 sg13g2_xnor2_1 _27432_ (.Y(_19141_),
    .A(\inv_result[175] ),
    .B(\inv_result[174] ));
 sg13g2_xor2_1 _27433_ (.B(\inv_result[172] ),
    .A(\inv_result[173] ),
    .X(_19142_));
 sg13g2_xnor2_1 _27434_ (.Y(_19143_),
    .A(_19141_),
    .B(_19142_));
 sg13g2_xnor2_1 _27435_ (.Y(_19144_),
    .A(_19140_),
    .B(_19143_));
 sg13g2_xor2_1 _27436_ (.B(\inv_result[162] ),
    .A(\inv_result[163] ),
    .X(_19145_));
 sg13g2_xor2_1 _27437_ (.B(\inv_result[160] ),
    .A(\inv_result[161] ),
    .X(_19146_));
 sg13g2_xnor2_1 _27438_ (.Y(_19147_),
    .A(_19145_),
    .B(_19146_));
 sg13g2_xnor2_1 _27439_ (.Y(_19148_),
    .A(\inv_result[167] ),
    .B(\inv_result[166] ));
 sg13g2_xor2_1 _27440_ (.B(\inv_result[164] ),
    .A(\inv_result[165] ),
    .X(_19149_));
 sg13g2_xnor2_1 _27441_ (.Y(_19150_),
    .A(_19148_),
    .B(_19149_));
 sg13g2_xnor2_1 _27442_ (.Y(_19151_),
    .A(_19147_),
    .B(_19150_));
 sg13g2_xnor2_1 _27443_ (.Y(_19152_),
    .A(_19144_),
    .B(_19151_));
 sg13g2_xor2_1 _27444_ (.B(\inv_result[218] ),
    .A(\inv_result[219] ),
    .X(_19153_));
 sg13g2_xor2_1 _27445_ (.B(\inv_result[216] ),
    .A(\inv_result[217] ),
    .X(_19154_));
 sg13g2_xnor2_1 _27446_ (.Y(_19155_),
    .A(_19153_),
    .B(_19154_));
 sg13g2_xnor2_1 _27447_ (.Y(_19156_),
    .A(\inv_result[223] ),
    .B(\inv_result[222] ));
 sg13g2_xor2_1 _27448_ (.B(\inv_result[220] ),
    .A(\inv_result[221] ),
    .X(_19157_));
 sg13g2_xnor2_1 _27449_ (.Y(_19158_),
    .A(_19156_),
    .B(_19157_));
 sg13g2_xnor2_1 _27450_ (.Y(_19159_),
    .A(_19155_),
    .B(_19158_));
 sg13g2_xor2_1 _27451_ (.B(\inv_result[210] ),
    .A(\inv_result[211] ),
    .X(_19160_));
 sg13g2_xor2_1 _27452_ (.B(\inv_result[208] ),
    .A(\inv_result[209] ),
    .X(_19161_));
 sg13g2_xnor2_1 _27453_ (.Y(_19162_),
    .A(_19160_),
    .B(_19161_));
 sg13g2_xnor2_1 _27454_ (.Y(_19163_),
    .A(\inv_result[215] ),
    .B(\inv_result[214] ));
 sg13g2_xor2_1 _27455_ (.B(\inv_result[212] ),
    .A(\inv_result[213] ),
    .X(_19164_));
 sg13g2_xnor2_1 _27456_ (.Y(_19165_),
    .A(_19163_),
    .B(_19164_));
 sg13g2_xnor2_1 _27457_ (.Y(_19166_),
    .A(_19162_),
    .B(_19165_));
 sg13g2_xnor2_1 _27458_ (.Y(_19167_),
    .A(_19159_),
    .B(_19166_));
 sg13g2_xnor2_1 _27459_ (.Y(_19168_),
    .A(_19152_),
    .B(_19167_));
 sg13g2_xor2_1 _27460_ (.B(\inv_result[198] ),
    .A(\inv_result[199] ),
    .X(_19169_));
 sg13g2_xor2_1 _27461_ (.B(\inv_result[192] ),
    .A(\inv_result[193] ),
    .X(_19170_));
 sg13g2_xnor2_1 _27462_ (.Y(_19171_),
    .A(_19169_),
    .B(_19170_));
 sg13g2_xnor2_1 _27463_ (.Y(_19172_),
    .A(\inv_result[197] ),
    .B(\inv_result[196] ));
 sg13g2_xor2_1 _27464_ (.B(\inv_result[194] ),
    .A(\inv_result[195] ),
    .X(_19173_));
 sg13g2_xnor2_1 _27465_ (.Y(_19174_),
    .A(_19172_),
    .B(_19173_));
 sg13g2_xnor2_1 _27466_ (.Y(_19175_),
    .A(_19171_),
    .B(_19174_));
 sg13g2_xor2_1 _27467_ (.B(\inv_result[202] ),
    .A(\inv_result[203] ),
    .X(_19176_));
 sg13g2_xor2_1 _27468_ (.B(\inv_result[200] ),
    .A(\inv_result[201] ),
    .X(_19177_));
 sg13g2_xnor2_1 _27469_ (.Y(_19178_),
    .A(_19176_),
    .B(_19177_));
 sg13g2_xnor2_1 _27470_ (.Y(_19179_),
    .A(\inv_result[207] ),
    .B(\inv_result[206] ));
 sg13g2_xor2_1 _27471_ (.B(\inv_result[204] ),
    .A(\inv_result[205] ),
    .X(_19180_));
 sg13g2_xnor2_1 _27472_ (.Y(_19181_),
    .A(_19179_),
    .B(_19180_));
 sg13g2_xnor2_1 _27473_ (.Y(_19182_),
    .A(_19178_),
    .B(_19181_));
 sg13g2_xnor2_1 _27474_ (.Y(_19183_),
    .A(_19175_),
    .B(_19182_));
 sg13g2_xnor2_1 _27475_ (.Y(_19184_),
    .A(\inv_result[187] ),
    .B(\inv_result[186] ));
 sg13g2_xor2_1 _27476_ (.B(\inv_result[184] ),
    .A(\inv_result[185] ),
    .X(_19185_));
 sg13g2_xnor2_1 _27477_ (.Y(_19186_),
    .A(_19184_),
    .B(_19185_));
 sg13g2_xnor2_1 _27478_ (.Y(_19187_),
    .A(\inv_result[191] ),
    .B(\inv_result[190] ));
 sg13g2_xor2_1 _27479_ (.B(\inv_result[188] ),
    .A(\inv_result[189] ),
    .X(_19188_));
 sg13g2_xnor2_1 _27480_ (.Y(_19189_),
    .A(_19187_),
    .B(_19188_));
 sg13g2_xnor2_1 _27481_ (.Y(_19190_),
    .A(_19186_),
    .B(_19189_));
 sg13g2_xor2_1 _27482_ (.B(\inv_result[182] ),
    .A(\inv_result[183] ),
    .X(_19191_));
 sg13g2_xor2_1 _27483_ (.B(\inv_result[176] ),
    .A(\inv_result[177] ),
    .X(_19192_));
 sg13g2_xnor2_1 _27484_ (.Y(_19193_),
    .A(_19191_),
    .B(_19192_));
 sg13g2_xnor2_1 _27485_ (.Y(_19194_),
    .A(\inv_result[181] ),
    .B(\inv_result[180] ));
 sg13g2_xor2_1 _27486_ (.B(\inv_result[178] ),
    .A(\inv_result[179] ),
    .X(_19195_));
 sg13g2_xnor2_1 _27487_ (.Y(_19196_),
    .A(_19194_),
    .B(_19195_));
 sg13g2_xnor2_1 _27488_ (.Y(_19197_),
    .A(_19193_),
    .B(_19196_));
 sg13g2_xnor2_1 _27489_ (.Y(_19198_),
    .A(_19190_),
    .B(_19197_));
 sg13g2_xnor2_1 _27490_ (.Y(_19199_),
    .A(_19183_),
    .B(_19198_));
 sg13g2_xnor2_1 _27491_ (.Y(_19200_),
    .A(_19168_),
    .B(_19199_));
 sg13g2_xnor2_1 _27492_ (.Y(_19201_),
    .A(_19137_),
    .B(_19200_));
 sg13g2_o21ai_1 _27493_ (.B1(net6647),
    .Y(_19202_),
    .A1(_19074_),
    .A2(_19201_));
 sg13g2_a21oi_1 _27494_ (.A1(_19074_),
    .A2(_19201_),
    .Y(_19203_),
    .B1(_19202_));
 sg13g2_a21o_1 _27495_ (.A2(net6911),
    .A1(net1192),
    .B1(_19203_),
    .X(_19204_));
 sg13g2_mux2_1 _27496_ (.A0(net3753),
    .A1(_19204_),
    .S(net6548),
    .X(_00190_));
 sg13g2_a22oi_1 _27497_ (.Y(_19205_),
    .B1(net6637),
    .B2(net3591),
    .A2(net6894),
    .A1(net1494));
 sg13g2_nor2_1 _27498_ (.A(net3660),
    .B(net6515),
    .Y(_19206_));
 sg13g2_a21oi_1 _27499_ (.A1(net6515),
    .A2(_19205_),
    .Y(_00191_),
    .B1(_19206_));
 sg13g2_a22oi_1 _27500_ (.Y(_19207_),
    .B1(net6644),
    .B2(net2179),
    .A2(net6906),
    .A1(net1324));
 sg13g2_nor2_1 _27501_ (.A(net3530),
    .B(net6536),
    .Y(_19208_));
 sg13g2_a21oi_1 _27502_ (.A1(net6536),
    .A2(_19207_),
    .Y(_00192_),
    .B1(_19208_));
 sg13g2_a22oi_1 _27503_ (.Y(_19209_),
    .B1(net6644),
    .B2(net1488),
    .A2(net6906),
    .A1(net2658));
 sg13g2_nor2_1 _27504_ (.A(net3629),
    .B(net6541),
    .Y(_19210_));
 sg13g2_a21oi_1 _27505_ (.A1(net6546),
    .A2(_19209_),
    .Y(_00193_),
    .B1(_19210_));
 sg13g2_a22oi_1 _27506_ (.Y(_19211_),
    .B1(net6641),
    .B2(net2336),
    .A2(net6906),
    .A1(net1814));
 sg13g2_nor2_1 _27507_ (.A(net3474),
    .B(net6536),
    .Y(_19212_));
 sg13g2_a21oi_1 _27508_ (.A1(net6536),
    .A2(_19211_),
    .Y(_00194_),
    .B1(_19212_));
 sg13g2_a22oi_1 _27509_ (.Y(_19213_),
    .B1(net6641),
    .B2(net2469),
    .A2(net6906),
    .A1(net2466));
 sg13g2_nor2_1 _27510_ (.A(net3385),
    .B(net6536),
    .Y(_19214_));
 sg13g2_a21oi_1 _27511_ (.A1(net6536),
    .A2(_19213_),
    .Y(_00195_),
    .B1(_19214_));
 sg13g2_a22oi_1 _27512_ (.Y(_19215_),
    .B1(net6641),
    .B2(net2111),
    .A2(net6906),
    .A1(net1199));
 sg13g2_nor2_1 _27513_ (.A(net3265),
    .B(net6537),
    .Y(_19216_));
 sg13g2_a21oi_1 _27514_ (.A1(net6537),
    .A2(_19215_),
    .Y(_00196_),
    .B1(_19216_));
 sg13g2_a22oi_1 _27515_ (.Y(_19217_),
    .B1(net6641),
    .B2(net2551),
    .A2(net6905),
    .A1(net2828));
 sg13g2_nor2_1 _27516_ (.A(net3458),
    .B(net6536),
    .Y(_19218_));
 sg13g2_a21oi_1 _27517_ (.A1(net6536),
    .A2(_19217_),
    .Y(_00197_),
    .B1(_19218_));
 sg13g2_a22oi_1 _27518_ (.Y(_19219_),
    .B1(net6645),
    .B2(net1383),
    .A2(net6911),
    .A1(\shift_reg[15] ));
 sg13g2_nor2_1 _27519_ (.A(net2778),
    .B(net6547),
    .Y(_19220_));
 sg13g2_a21oi_1 _27520_ (.A1(net6547),
    .A2(_19219_),
    .Y(_00198_),
    .B1(_19220_));
 sg13g2_a22oi_1 _27521_ (.Y(_19221_),
    .B1(net6645),
    .B2(net2099),
    .A2(net6915),
    .A1(\shift_reg[16] ));
 sg13g2_nor2_1 _27522_ (.A(net3526),
    .B(net6547),
    .Y(_19222_));
 sg13g2_a21oi_1 _27523_ (.A1(net6547),
    .A2(_19221_),
    .Y(_00199_),
    .B1(_19222_));
 sg13g2_a22oi_1 _27524_ (.Y(_19223_),
    .B1(net6645),
    .B2(net2236),
    .A2(net6910),
    .A1(net3530));
 sg13g2_nor2_1 _27525_ (.A(net3558),
    .B(net6546),
    .Y(_19224_));
 sg13g2_a21oi_1 _27526_ (.A1(net6546),
    .A2(_19223_),
    .Y(_00200_),
    .B1(_19224_));
 sg13g2_a22oi_1 _27527_ (.Y(_19225_),
    .B1(net6646),
    .B2(net3328),
    .A2(net6912),
    .A1(\shift_reg[18] ));
 sg13g2_nor2_1 _27528_ (.A(net3336),
    .B(net6549),
    .Y(_19226_));
 sg13g2_a21oi_1 _27529_ (.A1(net6549),
    .A2(_19225_),
    .Y(_00201_),
    .B1(_19226_));
 sg13g2_a22oi_1 _27530_ (.Y(_19227_),
    .B1(net6646),
    .B2(net1793),
    .A2(net6912),
    .A1(\shift_reg[19] ));
 sg13g2_nor2_1 _27531_ (.A(net3399),
    .B(net6549),
    .Y(_19228_));
 sg13g2_a21oi_1 _27532_ (.A1(net6549),
    .A2(_19227_),
    .Y(_00202_),
    .B1(_19228_));
 sg13g2_a22oi_1 _27533_ (.Y(_19229_),
    .B1(net6645),
    .B2(net1848),
    .A2(net6910),
    .A1(net3385));
 sg13g2_nor2_1 _27534_ (.A(net3538),
    .B(net6546),
    .Y(_19230_));
 sg13g2_a21oi_1 _27535_ (.A1(net6546),
    .A2(_19229_),
    .Y(_00203_),
    .B1(_19230_));
 sg13g2_a22oi_1 _27536_ (.Y(_19231_),
    .B1(net6645),
    .B2(net2136),
    .A2(net6911),
    .A1(\shift_reg[21] ));
 sg13g2_nor2_1 _27537_ (.A(net3246),
    .B(net6547),
    .Y(_19232_));
 sg13g2_a21oi_1 _27538_ (.A1(net6547),
    .A2(_19231_),
    .Y(_00204_),
    .B1(_19232_));
 sg13g2_a22oi_1 _27539_ (.Y(_19233_),
    .B1(net6645),
    .B2(net1910),
    .A2(net6911),
    .A1(\shift_reg[22] ));
 sg13g2_nor2_1 _27540_ (.A(net3206),
    .B(net6547),
    .Y(_19234_));
 sg13g2_a21oi_1 _27541_ (.A1(net6547),
    .A2(_19233_),
    .Y(_00205_),
    .B1(_19234_));
 sg13g2_a22oi_1 _27542_ (.Y(_19235_),
    .B1(net6645),
    .B2(net1485),
    .A2(net6911),
    .A1(net2778));
 sg13g2_nor2_1 _27543_ (.A(net3261),
    .B(net6549),
    .Y(_19236_));
 sg13g2_a21oi_1 _27544_ (.A1(net6548),
    .A2(_19235_),
    .Y(_00206_),
    .B1(_19236_));
 sg13g2_a22oi_1 _27545_ (.Y(_19237_),
    .B1(net6648),
    .B2(net1513),
    .A2(net6914),
    .A1(\shift_reg[24] ));
 sg13g2_nor2_1 _27546_ (.A(net2596),
    .B(net6551),
    .Y(_19238_));
 sg13g2_a21oi_1 _27547_ (.A1(net6551),
    .A2(_19237_),
    .Y(_00207_),
    .B1(_19238_));
 sg13g2_a22oi_1 _27548_ (.Y(_19239_),
    .B1(net6648),
    .B2(net2412),
    .A2(net6914),
    .A1(\shift_reg[25] ));
 sg13g2_nor2_1 _27549_ (.A(net2802),
    .B(net6552),
    .Y(_19240_));
 sg13g2_a21oi_1 _27550_ (.A1(net6552),
    .A2(_19239_),
    .Y(_00208_),
    .B1(_19240_));
 sg13g2_a22oi_1 _27551_ (.Y(_19241_),
    .B1(net6646),
    .B2(net1201),
    .A2(net6912),
    .A1(\shift_reg[26] ));
 sg13g2_nor2_1 _27552_ (.A(net3191),
    .B(net6550),
    .Y(_19242_));
 sg13g2_a21oi_1 _27553_ (.A1(net6549),
    .A2(_19241_),
    .Y(_00209_),
    .B1(_19242_));
 sg13g2_a22oi_1 _27554_ (.Y(_19243_),
    .B1(net6646),
    .B2(net2297),
    .A2(net6912),
    .A1(\shift_reg[27] ));
 sg13g2_nor2_1 _27555_ (.A(net3278),
    .B(net6549),
    .Y(_19244_));
 sg13g2_a21oi_1 _27556_ (.A1(net6549),
    .A2(_19243_),
    .Y(_00210_),
    .B1(_19244_));
 sg13g2_a22oi_1 _27557_ (.Y(_19245_),
    .B1(net6648),
    .B2(net2155),
    .A2(net6913),
    .A1(\shift_reg[28] ));
 sg13g2_nor2_1 _27558_ (.A(net2930),
    .B(net6551),
    .Y(_19246_));
 sg13g2_a21oi_1 _27559_ (.A1(net6551),
    .A2(_19245_),
    .Y(_00211_),
    .B1(_19246_));
 sg13g2_a22oi_1 _27560_ (.Y(_19247_),
    .B1(net6648),
    .B2(net1968),
    .A2(net6913),
    .A1(\shift_reg[29] ));
 sg13g2_nor2_1 _27561_ (.A(net3015),
    .B(net6552),
    .Y(_19248_));
 sg13g2_a21oi_1 _27562_ (.A1(net6552),
    .A2(_19247_),
    .Y(_00212_),
    .B1(_19248_));
 sg13g2_a22oi_1 _27563_ (.Y(_19249_),
    .B1(net6648),
    .B2(net1998),
    .A2(net6912),
    .A1(net3206));
 sg13g2_nor2_1 _27564_ (.A(net3424),
    .B(net6551),
    .Y(_19250_));
 sg13g2_a21oi_1 _27565_ (.A1(net6550),
    .A2(_19249_),
    .Y(_00213_),
    .B1(_19250_));
 sg13g2_a22oi_1 _27566_ (.Y(_19251_),
    .B1(net6648),
    .B2(net2005),
    .A2(net6914),
    .A1(\shift_reg[31] ));
 sg13g2_nor2_1 _27567_ (.A(net2251),
    .B(net6556),
    .Y(_19252_));
 sg13g2_a21oi_1 _27568_ (.A1(net6556),
    .A2(_19251_),
    .Y(_00214_),
    .B1(_19252_));
 sg13g2_a22oi_1 _27569_ (.Y(_19253_),
    .B1(net6648),
    .B2(net1190),
    .A2(net6913),
    .A1(net2596));
 sg13g2_nor2_1 _27570_ (.A(net3286),
    .B(net6551),
    .Y(_19254_));
 sg13g2_a21oi_1 _27571_ (.A1(net6551),
    .A2(_19253_),
    .Y(_00215_),
    .B1(_19254_));
 sg13g2_a22oi_1 _27572_ (.Y(_19255_),
    .B1(net6648),
    .B2(net2128),
    .A2(net6913),
    .A1(net2802));
 sg13g2_nor2_1 _27573_ (.A(net3565),
    .B(net6552),
    .Y(_19256_));
 sg13g2_a21oi_1 _27574_ (.A1(net6551),
    .A2(_19255_),
    .Y(_00216_),
    .B1(_19256_));
 sg13g2_a22oi_1 _27575_ (.Y(_19257_),
    .B1(net6650),
    .B2(net1732),
    .A2(net6920),
    .A1(net3191));
 sg13g2_nor2_1 _27576_ (.A(net3528),
    .B(net6556),
    .Y(_19258_));
 sg13g2_a21oi_1 _27577_ (.A1(net6556),
    .A2(_19257_),
    .Y(_00217_),
    .B1(_19258_));
 sg13g2_a22oi_1 _27578_ (.Y(_19259_),
    .B1(net6650),
    .B2(net3173),
    .A2(net6920),
    .A1(net3278));
 sg13g2_nor2_1 _27579_ (.A(net3492),
    .B(net6556),
    .Y(_19260_));
 sg13g2_a21oi_1 _27580_ (.A1(net6556),
    .A2(_19259_),
    .Y(_00218_),
    .B1(_19260_));
 sg13g2_a22oi_1 _27581_ (.Y(_19261_),
    .B1(net6656),
    .B2(net2058),
    .A2(net6920),
    .A1(\shift_reg[36] ));
 sg13g2_nor2_1 _27582_ (.A(net2781),
    .B(net6567),
    .Y(_19262_));
 sg13g2_a21oi_1 _27583_ (.A1(net6567),
    .A2(_19261_),
    .Y(_00219_),
    .B1(_19262_));
 sg13g2_a22oi_1 _27584_ (.Y(_19263_),
    .B1(net6656),
    .B2(\inv_result[29] ),
    .A2(net6920),
    .A1(\shift_reg[37] ));
 sg13g2_nor2_1 _27585_ (.A(net1764),
    .B(net6568),
    .Y(_19264_));
 sg13g2_a21oi_1 _27586_ (.A1(net6568),
    .A2(_19263_),
    .Y(_00220_),
    .B1(_19264_));
 sg13g2_a22oi_1 _27587_ (.Y(_19265_),
    .B1(net6656),
    .B2(net2037),
    .A2(net6920),
    .A1(net3424));
 sg13g2_nor2_1 _27588_ (.A(net3534),
    .B(net6556),
    .Y(_19266_));
 sg13g2_a21oi_1 _27589_ (.A1(net6575),
    .A2(_19265_),
    .Y(_00221_),
    .B1(_19266_));
 sg13g2_a22oi_1 _27590_ (.Y(_19267_),
    .B1(net6656),
    .B2(net1896),
    .A2(net6920),
    .A1(net2251));
 sg13g2_nor2_1 _27591_ (.A(net3116),
    .B(net6566),
    .Y(_19268_));
 sg13g2_a21oi_1 _27592_ (.A1(net6567),
    .A2(_19267_),
    .Y(_00222_),
    .B1(_19268_));
 sg13g2_a22oi_1 _27593_ (.Y(_19269_),
    .B1(net6656),
    .B2(net2648),
    .A2(net6922),
    .A1(\shift_reg[40] ));
 sg13g2_nor2_1 _27594_ (.A(net2822),
    .B(net6566),
    .Y(_19270_));
 sg13g2_a21oi_1 _27595_ (.A1(net6567),
    .A2(_19269_),
    .Y(_00223_),
    .B1(_19270_));
 sg13g2_a22oi_1 _27596_ (.Y(_19271_),
    .B1(net6656),
    .B2(net1548),
    .A2(net6922),
    .A1(\shift_reg[41] ));
 sg13g2_nor2_1 _27597_ (.A(net3100),
    .B(net6567),
    .Y(_19272_));
 sg13g2_a21oi_1 _27598_ (.A1(net6567),
    .A2(_19271_),
    .Y(_00224_),
    .B1(_19272_));
 sg13g2_a22oi_1 _27599_ (.Y(_19273_),
    .B1(net6658),
    .B2(net1196),
    .A2(net6922),
    .A1(\shift_reg[42] ));
 sg13g2_nor2_1 _27600_ (.A(net2733),
    .B(net6566),
    .Y(_19274_));
 sg13g2_a21oi_1 _27601_ (.A1(net6566),
    .A2(_19273_),
    .Y(_00225_),
    .B1(_19274_));
 sg13g2_a22oi_1 _27602_ (.Y(_19275_),
    .B1(net6658),
    .B2(net1525),
    .A2(net6922),
    .A1(\shift_reg[43] ));
 sg13g2_nor2_1 _27603_ (.A(net2953),
    .B(net6566),
    .Y(_19276_));
 sg13g2_a21oi_1 _27604_ (.A1(net6566),
    .A2(_19275_),
    .Y(_00226_),
    .B1(_19276_));
 sg13g2_a22oi_1 _27605_ (.Y(_19277_),
    .B1(net6658),
    .B2(net1563),
    .A2(net6921),
    .A1(net2781));
 sg13g2_nor2_1 _27606_ (.A(net3295),
    .B(net6568),
    .Y(_19278_));
 sg13g2_a21oi_1 _27607_ (.A1(net6568),
    .A2(_19277_),
    .Y(_00227_),
    .B1(_19278_));
 sg13g2_a22oi_1 _27608_ (.Y(_19279_),
    .B1(net6658),
    .B2(net2313),
    .A2(net6921),
    .A1(net1764));
 sg13g2_nor2_1 _27609_ (.A(net3060),
    .B(net6569),
    .Y(_19280_));
 sg13g2_a21oi_1 _27610_ (.A1(net6569),
    .A2(_19279_),
    .Y(_00228_),
    .B1(_19280_));
 sg13g2_a22oi_1 _27611_ (.Y(_19281_),
    .B1(net6658),
    .B2(net1596),
    .A2(net6922),
    .A1(\shift_reg[46] ));
 sg13g2_nor2_1 _27612_ (.A(net3467),
    .B(net6566),
    .Y(_19282_));
 sg13g2_a21oi_1 _27613_ (.A1(net6566),
    .A2(_19281_),
    .Y(_00229_),
    .B1(_19282_));
 sg13g2_a22oi_1 _27614_ (.Y(_19283_),
    .B1(net6658),
    .B2(net1986),
    .A2(net6922),
    .A1(\shift_reg[47] ));
 sg13g2_nor2_1 _27615_ (.A(net3040),
    .B(net6568),
    .Y(_19284_));
 sg13g2_a21oi_1 _27616_ (.A1(net6568),
    .A2(_19283_),
    .Y(_00230_),
    .B1(_19284_));
 sg13g2_a22oi_1 _27617_ (.Y(_19285_),
    .B1(net6657),
    .B2(net2040),
    .A2(net6922),
    .A1(net2822));
 sg13g2_nor2_1 _27618_ (.A(net3082),
    .B(net6571),
    .Y(_19286_));
 sg13g2_a21oi_1 _27619_ (.A1(net6568),
    .A2(_19285_),
    .Y(_00231_),
    .B1(_19286_));
 sg13g2_a22oi_1 _27620_ (.Y(_19287_),
    .B1(net6657),
    .B2(net2219),
    .A2(net6921),
    .A1(\shift_reg[49] ));
 sg13g2_nor2_1 _27621_ (.A(net2770),
    .B(net6568),
    .Y(_19288_));
 sg13g2_a21oi_1 _27622_ (.A1(net6569),
    .A2(_19287_),
    .Y(_00232_),
    .B1(_19288_));
 sg13g2_a22oi_1 _27623_ (.Y(_19289_),
    .B1(net6657),
    .B2(net1994),
    .A2(net6922),
    .A1(net2733));
 sg13g2_nor2_1 _27624_ (.A(net2933),
    .B(net6571),
    .Y(_19290_));
 sg13g2_a21oi_1 _27625_ (.A1(net6571),
    .A2(_19289_),
    .Y(_00233_),
    .B1(_19290_));
 sg13g2_a22oi_1 _27626_ (.Y(_19291_),
    .B1(net6658),
    .B2(net1407),
    .A2(net6921),
    .A1(net2953));
 sg13g2_nor2_1 _27627_ (.A(net3250),
    .B(net6569),
    .Y(_19292_));
 sg13g2_a21oi_1 _27628_ (.A1(net6569),
    .A2(_19291_),
    .Y(_00234_),
    .B1(_19292_));
 sg13g2_a22oi_1 _27629_ (.Y(_19293_),
    .B1(net6657),
    .B2(net2066),
    .A2(net6921),
    .A1(net3295));
 sg13g2_nor2_1 _27630_ (.A(net3380),
    .B(net6571),
    .Y(_19294_));
 sg13g2_a21oi_1 _27631_ (.A1(net6571),
    .A2(_19293_),
    .Y(_00235_),
    .B1(_19294_));
 sg13g2_a22oi_1 _27632_ (.Y(_19295_),
    .B1(net6657),
    .B2(net2210),
    .A2(net6921),
    .A1(net3060));
 sg13g2_nor2_1 _27633_ (.A(net3387),
    .B(net6571),
    .Y(_19296_));
 sg13g2_a21oi_1 _27634_ (.A1(net6572),
    .A2(_19295_),
    .Y(_00236_),
    .B1(_19296_));
 sg13g2_a22oi_1 _27635_ (.Y(_19297_),
    .B1(net6657),
    .B2(net2217),
    .A2(net6921),
    .A1(\shift_reg[54] ));
 sg13g2_nor2_1 _27636_ (.A(net3452),
    .B(net6570),
    .Y(_19298_));
 sg13g2_a21oi_1 _27637_ (.A1(net6570),
    .A2(_19297_),
    .Y(_00237_),
    .B1(_19298_));
 sg13g2_a22oi_1 _27638_ (.Y(_19299_),
    .B1(net6658),
    .B2(net2379),
    .A2(net6921),
    .A1(net3040));
 sg13g2_nor2_1 _27639_ (.A(net3227),
    .B(net6571),
    .Y(_19300_));
 sg13g2_a21oi_1 _27640_ (.A1(net6571),
    .A2(_19299_),
    .Y(_00238_),
    .B1(_19300_));
 sg13g2_a22oi_1 _27641_ (.Y(_19301_),
    .B1(net6657),
    .B2(net2237),
    .A2(net6926),
    .A1(net3082));
 sg13g2_nor2_1 _27642_ (.A(net3226),
    .B(net6577),
    .Y(_19302_));
 sg13g2_a21oi_1 _27643_ (.A1(net6577),
    .A2(_19301_),
    .Y(_00239_),
    .B1(_19302_));
 sg13g2_a22oi_1 _27644_ (.Y(_19303_),
    .B1(net6657),
    .B2(\inv_result[49] ),
    .A2(net6926),
    .A1(net2770));
 sg13g2_nor2_1 _27645_ (.A(net2900),
    .B(net6577),
    .Y(_19304_));
 sg13g2_a21oi_1 _27646_ (.A1(net6577),
    .A2(_19303_),
    .Y(_00240_),
    .B1(_19304_));
 sg13g2_a22oi_1 _27647_ (.Y(_19305_),
    .B1(net6661),
    .B2(net2218),
    .A2(net6926),
    .A1(net2933));
 sg13g2_nor2_1 _27648_ (.A(net3117),
    .B(net6577),
    .Y(_19306_));
 sg13g2_a21oi_1 _27649_ (.A1(net6577),
    .A2(_19305_),
    .Y(_00241_),
    .B1(_19306_));
 sg13g2_a22oi_1 _27650_ (.Y(_19307_),
    .B1(net6661),
    .B2(net2511),
    .A2(net6926),
    .A1(\shift_reg[59] ));
 sg13g2_nor2_1 _27651_ (.A(net3139),
    .B(net6577),
    .Y(_19308_));
 sg13g2_a21oi_1 _27652_ (.A1(net6577),
    .A2(_19307_),
    .Y(_00242_),
    .B1(_19308_));
 sg13g2_a22oi_1 _27653_ (.Y(_19309_),
    .B1(net6661),
    .B2(net1822),
    .A2(net6926),
    .A1(\shift_reg[60] ));
 sg13g2_nor2_1 _27654_ (.A(net3268),
    .B(net6576),
    .Y(_19310_));
 sg13g2_a21oi_1 _27655_ (.A1(net6576),
    .A2(_19309_),
    .Y(_00243_),
    .B1(_19310_));
 sg13g2_a22oi_1 _27656_ (.Y(_19311_),
    .B1(net6661),
    .B2(\inv_result[53] ),
    .A2(net6926),
    .A1(\shift_reg[61] ));
 sg13g2_nor2_1 _27657_ (.A(net2621),
    .B(net6576),
    .Y(_19312_));
 sg13g2_a21oi_1 _27658_ (.A1(net6576),
    .A2(_19311_),
    .Y(_00244_),
    .B1(_19312_));
 sg13g2_a22oi_1 _27659_ (.Y(_19313_),
    .B1(net6661),
    .B2(net1698),
    .A2(net6925),
    .A1(\shift_reg[62] ));
 sg13g2_nor2_1 _27660_ (.A(net3430),
    .B(net6576),
    .Y(_19314_));
 sg13g2_a21oi_1 _27661_ (.A1(net6576),
    .A2(_19313_),
    .Y(_00245_),
    .B1(_19314_));
 sg13g2_a22oi_1 _27662_ (.Y(_19315_),
    .B1(net6661),
    .B2(net2499),
    .A2(net6926),
    .A1(\shift_reg[63] ));
 sg13g2_nor2_1 _27663_ (.A(net3218),
    .B(net6579),
    .Y(_19316_));
 sg13g2_a21oi_1 _27664_ (.A1(net6582),
    .A2(_19315_),
    .Y(_00246_),
    .B1(_19316_));
 sg13g2_a22oi_1 _27665_ (.Y(_19317_),
    .B1(net6662),
    .B2(net2081),
    .A2(net6925),
    .A1(net3226));
 sg13g2_nor2_1 _27666_ (.A(net3439),
    .B(net6578),
    .Y(_19318_));
 sg13g2_a21oi_1 _27667_ (.A1(net6579),
    .A2(_19317_),
    .Y(_00247_),
    .B1(_19318_));
 sg13g2_a22oi_1 _27668_ (.Y(_19319_),
    .B1(net6662),
    .B2(net2838),
    .A2(net6925),
    .A1(net2900));
 sg13g2_nor2_1 _27669_ (.A(net3031),
    .B(net6578),
    .Y(_19320_));
 sg13g2_a21oi_1 _27670_ (.A1(net6578),
    .A2(_19319_),
    .Y(_00248_),
    .B1(_19320_));
 sg13g2_a22oi_1 _27671_ (.Y(_19321_),
    .B1(net6662),
    .B2(net2873),
    .A2(net6925),
    .A1(net3117));
 sg13g2_nor2_1 _27672_ (.A(net3577),
    .B(net6578),
    .Y(_19322_));
 sg13g2_a21oi_1 _27673_ (.A1(net6579),
    .A2(_19321_),
    .Y(_00249_),
    .B1(_19322_));
 sg13g2_a22oi_1 _27674_ (.Y(_19323_),
    .B1(net6662),
    .B2(net2752),
    .A2(net6925),
    .A1(net3139));
 sg13g2_nor2_1 _27675_ (.A(net3461),
    .B(net6581),
    .Y(_19324_));
 sg13g2_a21oi_1 _27676_ (.A1(net6578),
    .A2(_19323_),
    .Y(_00250_),
    .B1(_19324_));
 sg13g2_a22oi_1 _27677_ (.Y(_19325_),
    .B1(net6661),
    .B2(net2068),
    .A2(net6926),
    .A1(net3268));
 sg13g2_nor2_1 _27678_ (.A(net3442),
    .B(net6576),
    .Y(_19326_));
 sg13g2_a21oi_1 _27679_ (.A1(net6576),
    .A2(_19325_),
    .Y(_00251_),
    .B1(_19326_));
 sg13g2_a22oi_1 _27680_ (.Y(_19327_),
    .B1(net6662),
    .B2(\inv_result[61] ),
    .A2(net6925),
    .A1(net2621));
 sg13g2_nor2_1 _27681_ (.A(net3443),
    .B(net6578),
    .Y(_19328_));
 sg13g2_a21oi_1 _27682_ (.A1(net6579),
    .A2(_19327_),
    .Y(_00252_),
    .B1(_19328_));
 sg13g2_a22oi_1 _27683_ (.Y(_19329_),
    .B1(net6661),
    .B2(net2566),
    .A2(net6925),
    .A1(\shift_reg[70] ));
 sg13g2_nor2_1 _27684_ (.A(net3427),
    .B(net6579),
    .Y(_19330_));
 sg13g2_a21oi_1 _27685_ (.A1(net6579),
    .A2(_19329_),
    .Y(_00253_),
    .B1(_19330_));
 sg13g2_a22oi_1 _27686_ (.Y(_19331_),
    .B1(net6662),
    .B2(net2558),
    .A2(net6925),
    .A1(net3218));
 sg13g2_nor2_1 _27687_ (.A(net3440),
    .B(net6578),
    .Y(_19332_));
 sg13g2_a21oi_1 _27688_ (.A1(net6578),
    .A2(_19331_),
    .Y(_00254_),
    .B1(_19332_));
 sg13g2_a22oi_1 _27689_ (.Y(_19333_),
    .B1(net6672),
    .B2(\inv_result[64] ),
    .A2(net6932),
    .A1(\shift_reg[72] ));
 sg13g2_nor2_1 _27690_ (.A(net2701),
    .B(net6593),
    .Y(_19334_));
 sg13g2_a21oi_1 _27691_ (.A1(net6593),
    .A2(_19333_),
    .Y(_00255_),
    .B1(_19334_));
 sg13g2_a22oi_1 _27692_ (.Y(_19335_),
    .B1(net6672),
    .B2(net2711),
    .A2(net6932),
    .A1(\shift_reg[73] ));
 sg13g2_nor2_1 _27693_ (.A(net2994),
    .B(net6595),
    .Y(_19336_));
 sg13g2_a21oi_1 _27694_ (.A1(net6593),
    .A2(_19335_),
    .Y(_00256_),
    .B1(_19336_));
 sg13g2_a22oi_1 _27695_ (.Y(_19337_),
    .B1(net6672),
    .B2(\inv_result[66] ),
    .A2(net6932),
    .A1(\shift_reg[74] ));
 sg13g2_nor2_1 _27696_ (.A(net2816),
    .B(net6594),
    .Y(_19338_));
 sg13g2_a21oi_1 _27697_ (.A1(net6593),
    .A2(_19337_),
    .Y(_00257_),
    .B1(_19338_));
 sg13g2_a22oi_1 _27698_ (.Y(_19339_),
    .B1(net6668),
    .B2(net2250),
    .A2(net6934),
    .A1(\shift_reg[75] ));
 sg13g2_nor2_1 _27699_ (.A(net2434),
    .B(net6595),
    .Y(_19340_));
 sg13g2_a21oi_1 _27700_ (.A1(net6595),
    .A2(_19339_),
    .Y(_00258_),
    .B1(_19340_));
 sg13g2_a22oi_1 _27701_ (.Y(_19341_),
    .B1(net6672),
    .B2(net1360),
    .A2(net6932),
    .A1(\shift_reg[76] ));
 sg13g2_nor2_1 _27702_ (.A(net2912),
    .B(net6593),
    .Y(_19342_));
 sg13g2_a21oi_1 _27703_ (.A1(net6593),
    .A2(_19341_),
    .Y(_00259_),
    .B1(_19342_));
 sg13g2_a22oi_1 _27704_ (.Y(_19343_),
    .B1(net6672),
    .B2(net3057),
    .A2(net6932),
    .A1(\shift_reg[77] ));
 sg13g2_nor2_1 _27705_ (.A(net3126),
    .B(net6593),
    .Y(_19344_));
 sg13g2_a21oi_1 _27706_ (.A1(net6593),
    .A2(_19343_),
    .Y(_00260_),
    .B1(_19344_));
 sg13g2_a22oi_1 _27707_ (.Y(_19345_),
    .B1(net6668),
    .B2(net1923),
    .A2(net6934),
    .A1(\shift_reg[78] ));
 sg13g2_nor2_1 _27708_ (.A(net3088),
    .B(net6595),
    .Y(_19346_));
 sg13g2_a21oi_1 _27709_ (.A1(net6595),
    .A2(_19345_),
    .Y(_00261_),
    .B1(_19346_));
 sg13g2_a22oi_1 _27710_ (.Y(_19347_),
    .B1(net6668),
    .B2(net2630),
    .A2(net6934),
    .A1(\shift_reg[79] ));
 sg13g2_nor2_1 _27711_ (.A(net3168),
    .B(net6595),
    .Y(_19348_));
 sg13g2_a21oi_1 _27712_ (.A1(net6603),
    .A2(_19347_),
    .Y(_00262_),
    .B1(_19348_));
 sg13g2_a22oi_1 _27713_ (.Y(_19349_),
    .B1(net6671),
    .B2(net1406),
    .A2(net6934),
    .A1(\shift_reg[80] ));
 sg13g2_nor2_1 _27714_ (.A(net2410),
    .B(net6596),
    .Y(_19350_));
 sg13g2_a21oi_1 _27715_ (.A1(net6596),
    .A2(_19349_),
    .Y(_00263_),
    .B1(_19350_));
 sg13g2_a22oi_1 _27716_ (.Y(_19351_),
    .B1(net6671),
    .B2(net3174),
    .A2(net6934),
    .A1(net2994));
 sg13g2_nor2_1 _27717_ (.A(net3297),
    .B(net6596),
    .Y(_19352_));
 sg13g2_a21oi_1 _27718_ (.A1(net6596),
    .A2(_19351_),
    .Y(_00264_),
    .B1(_19352_));
 sg13g2_a22oi_1 _27719_ (.Y(_19353_),
    .B1(net6668),
    .B2(net2373),
    .A2(net6933),
    .A1(net2816));
 sg13g2_nor2_1 _27720_ (.A(net3346),
    .B(net6597),
    .Y(_19354_));
 sg13g2_a21oi_1 _27721_ (.A1(net6597),
    .A2(_19353_),
    .Y(_00265_),
    .B1(_19354_));
 sg13g2_a22oi_1 _27722_ (.Y(_19355_),
    .B1(net6668),
    .B2(net2161),
    .A2(net6933),
    .A1(net2434));
 sg13g2_nor2_1 _27723_ (.A(net2993),
    .B(net6596),
    .Y(_19356_));
 sg13g2_a21oi_1 _27724_ (.A1(net6596),
    .A2(_19355_),
    .Y(_00266_),
    .B1(_19356_));
 sg13g2_a22oi_1 _27725_ (.Y(_19357_),
    .B1(net6668),
    .B2(net1207),
    .A2(net6933),
    .A1(net2912));
 sg13g2_nor2_1 _27726_ (.A(net3118),
    .B(net6597),
    .Y(_19358_));
 sg13g2_a21oi_1 _27727_ (.A1(net6597),
    .A2(_19357_),
    .Y(_00267_),
    .B1(_19358_));
 sg13g2_a22oi_1 _27728_ (.Y(_19359_),
    .B1(net6671),
    .B2(net1298),
    .A2(net6933),
    .A1(\shift_reg[85] ));
 sg13g2_nor2_1 _27729_ (.A(net3086),
    .B(net6595),
    .Y(_19360_));
 sg13g2_a21oi_1 _27730_ (.A1(net6595),
    .A2(_19359_),
    .Y(_00268_),
    .B1(_19360_));
 sg13g2_a22oi_1 _27731_ (.Y(_19361_),
    .B1(net6670),
    .B2(net1627),
    .A2(net6933),
    .A1(net3088));
 sg13g2_nor2_1 _27732_ (.A(net3251),
    .B(net6596),
    .Y(_19362_));
 sg13g2_a21oi_1 _27733_ (.A1(net6596),
    .A2(_19361_),
    .Y(_00269_),
    .B1(_19362_));
 sg13g2_a22oi_1 _27734_ (.Y(_19363_),
    .B1(net6670),
    .B2(net1991),
    .A2(net6933),
    .A1(\shift_reg[87] ));
 sg13g2_nor2_1 _27735_ (.A(net3048),
    .B(net6597),
    .Y(_19364_));
 sg13g2_a21oi_1 _27736_ (.A1(net6597),
    .A2(_19363_),
    .Y(_00270_),
    .B1(_19364_));
 sg13g2_a22oi_1 _27737_ (.Y(_19365_),
    .B1(net6668),
    .B2(net2135),
    .A2(net6933),
    .A1(net2410));
 sg13g2_nor2_1 _27738_ (.A(net3061),
    .B(net6598),
    .Y(_19366_));
 sg13g2_a21oi_1 _27739_ (.A1(net6598),
    .A2(_19365_),
    .Y(_00271_),
    .B1(_19366_));
 sg13g2_a22oi_1 _27740_ (.Y(_19367_),
    .B1(net6668),
    .B2(net2936),
    .A2(net6933),
    .A1(net3297));
 sg13g2_nor2_1 _27741_ (.A(net3423),
    .B(net6598),
    .Y(_19368_));
 sg13g2_a21oi_1 _27742_ (.A1(net6598),
    .A2(_19367_),
    .Y(_00272_),
    .B1(_19368_));
 sg13g2_a22oi_1 _27743_ (.Y(_19369_),
    .B1(net6670),
    .B2(net2046),
    .A2(net6936),
    .A1(\shift_reg[90] ));
 sg13g2_nor2_1 _27744_ (.A(net3122),
    .B(net6599),
    .Y(_19370_));
 sg13g2_a21oi_1 _27745_ (.A1(net6599),
    .A2(_19369_),
    .Y(_00273_),
    .B1(_19370_));
 sg13g2_a22oi_1 _27746_ (.Y(_19371_),
    .B1(net6670),
    .B2(net1220),
    .A2(net6936),
    .A1(\shift_reg[91] ));
 sg13g2_nor2_1 _27747_ (.A(net2571),
    .B(net6602),
    .Y(_19372_));
 sg13g2_a21oi_1 _27748_ (.A1(net6602),
    .A2(_19371_),
    .Y(_00274_),
    .B1(_19372_));
 sg13g2_a22oi_1 _27749_ (.Y(_19373_),
    .B1(net6670),
    .B2(net2131),
    .A2(net6936),
    .A1(\shift_reg[92] ));
 sg13g2_nor2_1 _27750_ (.A(net2853),
    .B(net6601),
    .Y(_19374_));
 sg13g2_a21oi_1 _27751_ (.A1(net6601),
    .A2(_19373_),
    .Y(_00275_),
    .B1(_19374_));
 sg13g2_a22oi_1 _27752_ (.Y(_19375_),
    .B1(net6669),
    .B2(\inv_result[85] ),
    .A2(net6935),
    .A1(\shift_reg[93] ));
 sg13g2_nor2_1 _27753_ (.A(net2934),
    .B(net6599),
    .Y(_19376_));
 sg13g2_a21oi_1 _27754_ (.A1(net6599),
    .A2(_19375_),
    .Y(_00276_),
    .B1(_19376_));
 sg13g2_a22oi_1 _27755_ (.Y(_19377_),
    .B1(net6669),
    .B2(net2449),
    .A2(net6935),
    .A1(\shift_reg[94] ));
 sg13g2_nor2_1 _27756_ (.A(net3193),
    .B(net6599),
    .Y(_19378_));
 sg13g2_a21oi_1 _27757_ (.A1(net6599),
    .A2(_19377_),
    .Y(_00277_),
    .B1(_19378_));
 sg13g2_a22oi_1 _27758_ (.Y(_19379_),
    .B1(net6670),
    .B2(net2315),
    .A2(net6936),
    .A1(net3048));
 sg13g2_nor2_1 _27759_ (.A(net3152),
    .B(net6601),
    .Y(_19380_));
 sg13g2_a21oi_1 _27760_ (.A1(net6601),
    .A2(_19379_),
    .Y(_00278_),
    .B1(_19380_));
 sg13g2_a22oi_1 _27761_ (.Y(_19381_),
    .B1(net6670),
    .B2(net1240),
    .A2(net6936),
    .A1(net3061));
 sg13g2_nor2_1 _27762_ (.A(net3600),
    .B(net6601),
    .Y(_19382_));
 sg13g2_a21oi_1 _27763_ (.A1(net6601),
    .A2(_19381_),
    .Y(_00279_),
    .B1(_19382_));
 sg13g2_a22oi_1 _27764_ (.Y(_19383_),
    .B1(net6670),
    .B2(net2644),
    .A2(net6936),
    .A1(net3423));
 sg13g2_nor2_1 _27765_ (.A(net3441),
    .B(net6601),
    .Y(_19384_));
 sg13g2_a21oi_1 _27766_ (.A1(net6601),
    .A2(_19383_),
    .Y(_00280_),
    .B1(_19384_));
 sg13g2_a22oi_1 _27767_ (.Y(_19385_),
    .B1(net6669),
    .B2(net1566),
    .A2(net6935),
    .A1(net3122));
 sg13g2_nor2_1 _27768_ (.A(net3500),
    .B(net6600),
    .Y(_19386_));
 sg13g2_a21oi_1 _27769_ (.A1(net6600),
    .A2(_19385_),
    .Y(_00281_),
    .B1(_19386_));
 sg13g2_a22oi_1 _27770_ (.Y(_19387_),
    .B1(net6669),
    .B2(net3370),
    .A2(net6935),
    .A1(net2571));
 sg13g2_nor2_1 _27771_ (.A(net3661),
    .B(net6600),
    .Y(_19388_));
 sg13g2_a21oi_1 _27772_ (.A1(net6600),
    .A2(_19387_),
    .Y(_00282_),
    .B1(_19388_));
 sg13g2_a22oi_1 _27773_ (.Y(_19389_),
    .B1(net6669),
    .B2(net1208),
    .A2(net6935),
    .A1(net2853));
 sg13g2_nor2_1 _27774_ (.A(net3373),
    .B(net6600),
    .Y(_19390_));
 sg13g2_a21oi_1 _27775_ (.A1(net6600),
    .A2(_19389_),
    .Y(_00283_),
    .B1(_19390_));
 sg13g2_a22oi_1 _27776_ (.Y(_19391_),
    .B1(net6669),
    .B2(net1326),
    .A2(net6935),
    .A1(net2934));
 sg13g2_nor2_1 _27777_ (.A(net3517),
    .B(net6600),
    .Y(_19392_));
 sg13g2_a21oi_1 _27778_ (.A1(net6599),
    .A2(_19391_),
    .Y(_00284_),
    .B1(_19392_));
 sg13g2_a22oi_1 _27779_ (.Y(_19393_),
    .B1(net6669),
    .B2(net1645),
    .A2(net6935),
    .A1(net3193));
 sg13g2_nor2_1 _27780_ (.A(net3464),
    .B(net6594),
    .Y(_19394_));
 sg13g2_a21oi_1 _27781_ (.A1(net6594),
    .A2(_19393_),
    .Y(_00285_),
    .B1(_19394_));
 sg13g2_a22oi_1 _27782_ (.Y(_19395_),
    .B1(net6669),
    .B2(net2162),
    .A2(net6935),
    .A1(net3152));
 sg13g2_nor2_1 _27783_ (.A(net3216),
    .B(net6600),
    .Y(_19396_));
 sg13g2_a21oi_1 _27784_ (.A1(net6599),
    .A2(_19395_),
    .Y(_00286_),
    .B1(_19396_));
 sg13g2_a22oi_1 _27785_ (.Y(_19397_),
    .B1(net6664),
    .B2(net2061),
    .A2(net6927),
    .A1(\shift_reg[104] ));
 sg13g2_nor2_1 _27786_ (.A(net2554),
    .B(net6580),
    .Y(_19398_));
 sg13g2_a21oi_1 _27787_ (.A1(net6580),
    .A2(_19397_),
    .Y(_00287_),
    .B1(_19398_));
 sg13g2_a22oi_1 _27788_ (.Y(_19399_),
    .B1(net6664),
    .B2(net2258),
    .A2(net6932),
    .A1(\shift_reg[105] ));
 sg13g2_nor2_1 _27789_ (.A(net2651),
    .B(net6580),
    .Y(_19400_));
 sg13g2_a21oi_1 _27790_ (.A1(net6580),
    .A2(_19399_),
    .Y(_00288_),
    .B1(_19400_));
 sg13g2_a22oi_1 _27791_ (.Y(_19401_),
    .B1(net6664),
    .B2(net1202),
    .A2(net6927),
    .A1(\shift_reg[106] ));
 sg13g2_nor2_1 _27792_ (.A(net2914),
    .B(net6580),
    .Y(_19402_));
 sg13g2_a21oi_1 _27793_ (.A1(net6580),
    .A2(_19401_),
    .Y(_00289_),
    .B1(_19402_));
 sg13g2_a22oi_1 _27794_ (.Y(_19403_),
    .B1(net6664),
    .B2(net1721),
    .A2(net6932),
    .A1(\shift_reg[107] ));
 sg13g2_nor2_1 _27795_ (.A(net3147),
    .B(net6580),
    .Y(_19404_));
 sg13g2_a21oi_1 _27796_ (.A1(net6580),
    .A2(_19403_),
    .Y(_00290_),
    .B1(_19404_));
 sg13g2_a22oi_1 _27797_ (.Y(_19405_),
    .B1(net6673),
    .B2(net2544),
    .A2(net6932),
    .A1(\shift_reg[108] ));
 sg13g2_nor2_1 _27798_ (.A(net3183),
    .B(net6594),
    .Y(_19406_));
 sg13g2_a21oi_1 _27799_ (.A1(net6594),
    .A2(_19405_),
    .Y(_00291_),
    .B1(_19406_));
 sg13g2_a22oi_1 _27800_ (.Y(_19407_),
    .B1(net6664),
    .B2(net1245),
    .A2(net6927),
    .A1(\shift_reg[109] ));
 sg13g2_nor2_1 _27801_ (.A(net2115),
    .B(net6581),
    .Y(_19408_));
 sg13g2_a21oi_1 _27802_ (.A1(net6581),
    .A2(_19407_),
    .Y(_00292_),
    .B1(_19408_));
 sg13g2_a22oi_1 _27803_ (.Y(_19409_),
    .B1(net6673),
    .B2(net1244),
    .A2(net6937),
    .A1(\shift_reg[110] ));
 sg13g2_nor2_1 _27804_ (.A(net2923),
    .B(net6594),
    .Y(_19410_));
 sg13g2_a21oi_1 _27805_ (.A1(net6604),
    .A2(_19409_),
    .Y(_00293_),
    .B1(_19410_));
 sg13g2_a22oi_1 _27806_ (.Y(_19411_),
    .B1(net6673),
    .B2(net1752),
    .A2(net6937),
    .A1(net3216));
 sg13g2_nor2_1 _27807_ (.A(net3325),
    .B(net6594),
    .Y(_19412_));
 sg13g2_a21oi_1 _27808_ (.A1(net6604),
    .A2(_19411_),
    .Y(_00294_),
    .B1(_19412_));
 sg13g2_a22oi_1 _27809_ (.Y(_19413_),
    .B1(net6664),
    .B2(net1209),
    .A2(net6928),
    .A1(\shift_reg[112] ));
 sg13g2_nor2_1 _27810_ (.A(net2334),
    .B(net6590),
    .Y(_19414_));
 sg13g2_a21oi_1 _27811_ (.A1(net6590),
    .A2(_19413_),
    .Y(_00295_),
    .B1(_19414_));
 sg13g2_a22oi_1 _27812_ (.Y(_19415_),
    .B1(net6664),
    .B2(net2390),
    .A2(net6928),
    .A1(\shift_reg[113] ));
 sg13g2_nor2_1 _27813_ (.A(net2423),
    .B(net6591),
    .Y(_19416_));
 sg13g2_a21oi_1 _27814_ (.A1(net6591),
    .A2(_19415_),
    .Y(_00296_),
    .B1(_19416_));
 sg13g2_a22oi_1 _27815_ (.Y(_19417_),
    .B1(net6664),
    .B2(net1995),
    .A2(net6928),
    .A1(\shift_reg[114] ));
 sg13g2_nor2_1 _27816_ (.A(net2451),
    .B(net6590),
    .Y(_19418_));
 sg13g2_a21oi_1 _27817_ (.A1(net6590),
    .A2(_19417_),
    .Y(_00297_),
    .B1(_19418_));
 sg13g2_a22oi_1 _27818_ (.Y(_19419_),
    .B1(net6665),
    .B2(net1254),
    .A2(net6938),
    .A1(\shift_reg[115] ));
 sg13g2_nor2_1 _27819_ (.A(net1976),
    .B(net6591),
    .Y(_19420_));
 sg13g2_a21oi_1 _27820_ (.A1(net6591),
    .A2(_19419_),
    .Y(_00298_),
    .B1(_19420_));
 sg13g2_a22oi_1 _27821_ (.Y(_19421_),
    .B1(net6665),
    .B2(net1607),
    .A2(net6928),
    .A1(\shift_reg[116] ));
 sg13g2_nor2_1 _27822_ (.A(net2347),
    .B(net6590),
    .Y(_19422_));
 sg13g2_a21oi_1 _27823_ (.A1(net6590),
    .A2(_19421_),
    .Y(_00299_),
    .B1(_19422_));
 sg13g2_a22oi_1 _27824_ (.Y(_19423_),
    .B1(net6665),
    .B2(net1403),
    .A2(net6928),
    .A1(net2115));
 sg13g2_nor2_1 _27825_ (.A(net2459),
    .B(net6589),
    .Y(_19424_));
 sg13g2_a21oi_1 _27826_ (.A1(net6589),
    .A2(_19423_),
    .Y(_00300_),
    .B1(_19424_));
 sg13g2_a22oi_1 _27827_ (.Y(_19425_),
    .B1(net6665),
    .B2(net1837),
    .A2(net6928),
    .A1(net2923));
 sg13g2_nor2_1 _27828_ (.A(net3092),
    .B(net6589),
    .Y(_19426_));
 sg13g2_a21oi_1 _27829_ (.A1(net6590),
    .A2(_19425_),
    .Y(_00301_),
    .B1(_19426_));
 sg13g2_a22oi_1 _27830_ (.Y(_19427_),
    .B1(net6665),
    .B2(\inv_result[111] ),
    .A2(net6928),
    .A1(\shift_reg[119] ));
 sg13g2_nor2_1 _27831_ (.A(net1936),
    .B(net6589),
    .Y(_19428_));
 sg13g2_a21oi_1 _27832_ (.A1(net6589),
    .A2(_19427_),
    .Y(_00302_),
    .B1(_19428_));
 sg13g2_a22oi_1 _27833_ (.Y(_19429_),
    .B1(net6666),
    .B2(\inv_result[112] ),
    .A2(net6928),
    .A1(\shift_reg[120] ));
 sg13g2_nor2_1 _27834_ (.A(net2019),
    .B(net6588),
    .Y(_19430_));
 sg13g2_a21oi_1 _27835_ (.A1(net6588),
    .A2(_19429_),
    .Y(_00303_),
    .B1(_19430_));
 sg13g2_a22oi_1 _27836_ (.Y(_19431_),
    .B1(net6667),
    .B2(net2281),
    .A2(net6930),
    .A1(net2423));
 sg13g2_nor2_1 _27837_ (.A(net2645),
    .B(net6588),
    .Y(_19432_));
 sg13g2_a21oi_1 _27838_ (.A1(net6588),
    .A2(_19431_),
    .Y(_00304_),
    .B1(_19432_));
 sg13g2_a22oi_1 _27839_ (.Y(_19433_),
    .B1(net6666),
    .B2(net1862),
    .A2(net6930),
    .A1(net2451));
 sg13g2_nor2_1 _27840_ (.A(net2965),
    .B(net6591),
    .Y(_19434_));
 sg13g2_a21oi_1 _27841_ (.A1(net6590),
    .A2(_19433_),
    .Y(_00305_),
    .B1(_19434_));
 sg13g2_a22oi_1 _27842_ (.Y(_19435_),
    .B1(net6666),
    .B2(net1603),
    .A2(net6930),
    .A1(net1976));
 sg13g2_nor2_1 _27843_ (.A(net2286),
    .B(net6589),
    .Y(_19436_));
 sg13g2_a21oi_1 _27844_ (.A1(net6588),
    .A2(_19435_),
    .Y(_00306_),
    .B1(_19436_));
 sg13g2_a22oi_1 _27845_ (.Y(_19437_),
    .B1(net6666),
    .B2(net1214),
    .A2(net6929),
    .A1(net2347));
 sg13g2_nor2_1 _27846_ (.A(net3001),
    .B(net6589),
    .Y(_19438_));
 sg13g2_a21oi_1 _27847_ (.A1(net6588),
    .A2(_19437_),
    .Y(_00307_),
    .B1(_19438_));
 sg13g2_a22oi_1 _27848_ (.Y(_19439_),
    .B1(net6666),
    .B2(\inv_result[117] ),
    .A2(net6930),
    .A1(net2459));
 sg13g2_nor2_1 _27849_ (.A(net2576),
    .B(net6586),
    .Y(_19440_));
 sg13g2_a21oi_1 _27850_ (.A1(net6586),
    .A2(_19439_),
    .Y(_00308_),
    .B1(_19440_));
 sg13g2_a22oi_1 _27851_ (.Y(_19441_),
    .B1(net6666),
    .B2(net2190),
    .A2(net6929),
    .A1(\shift_reg[126] ));
 sg13g2_nor2_1 _27852_ (.A(net2428),
    .B(net6588),
    .Y(_19442_));
 sg13g2_a21oi_1 _27853_ (.A1(net6588),
    .A2(_19441_),
    .Y(_00309_),
    .B1(_19442_));
 sg13g2_a22oi_1 _27854_ (.Y(_19443_),
    .B1(net6663),
    .B2(net2047),
    .A2(net6929),
    .A1(net1936));
 sg13g2_nor2_1 _27855_ (.A(net2303),
    .B(net6584),
    .Y(_19444_));
 sg13g2_a21oi_1 _27856_ (.A1(net6584),
    .A2(_19443_),
    .Y(_00310_),
    .B1(_19444_));
 sg13g2_a22oi_1 _27857_ (.Y(_19445_),
    .B1(net6666),
    .B2(\inv_result[120] ),
    .A2(net6930),
    .A1(\shift_reg[128] ));
 sg13g2_nor2_1 _27858_ (.A(net1974),
    .B(net6586),
    .Y(_19446_));
 sg13g2_a21oi_1 _27859_ (.A1(net6586),
    .A2(_19445_),
    .Y(_00311_),
    .B1(_19446_));
 sg13g2_a22oi_1 _27860_ (.Y(_19447_),
    .B1(net6666),
    .B2(\inv_result[121] ),
    .A2(net6930),
    .A1(\shift_reg[129] ));
 sg13g2_nor2_1 _27861_ (.A(net2291),
    .B(net6586),
    .Y(_19448_));
 sg13g2_a21oi_1 _27862_ (.A1(net6583),
    .A2(_19447_),
    .Y(_00312_),
    .B1(_19448_));
 sg13g2_a22oi_1 _27863_ (.Y(_19449_),
    .B1(net6663),
    .B2(net2057),
    .A2(net6929),
    .A1(net2965));
 sg13g2_nor2_1 _27864_ (.A(net3379),
    .B(net6584),
    .Y(_19450_));
 sg13g2_a21oi_1 _27865_ (.A1(net6583),
    .A2(_19449_),
    .Y(_00313_),
    .B1(_19450_));
 sg13g2_a22oi_1 _27866_ (.Y(_19451_),
    .B1(net6667),
    .B2(net2145),
    .A2(net6929),
    .A1(net2286));
 sg13g2_nor2_1 _27867_ (.A(net3487),
    .B(net6583),
    .Y(_19452_));
 sg13g2_a21oi_1 _27868_ (.A1(net6583),
    .A2(_19451_),
    .Y(_00314_),
    .B1(_19452_));
 sg13g2_a22oi_1 _27869_ (.Y(_19453_),
    .B1(net6663),
    .B2(net1893),
    .A2(net6931),
    .A1(net3001));
 sg13g2_nor2_1 _27870_ (.A(net3429),
    .B(net6585),
    .Y(_19454_));
 sg13g2_a21oi_1 _27871_ (.A1(net6585),
    .A2(_19453_),
    .Y(_00315_),
    .B1(_19454_));
 sg13g2_a22oi_1 _27872_ (.Y(_19455_),
    .B1(net6663),
    .B2(net1270),
    .A2(net6931),
    .A1(net2576));
 sg13g2_nor2_1 _27873_ (.A(net3357),
    .B(net6585),
    .Y(_19456_));
 sg13g2_a21oi_1 _27874_ (.A1(net6585),
    .A2(_19455_),
    .Y(_00316_),
    .B1(_19456_));
 sg13g2_a22oi_1 _27875_ (.Y(_19457_),
    .B1(net6663),
    .B2(net1569),
    .A2(net6929),
    .A1(net2428));
 sg13g2_nor2_1 _27876_ (.A(net3449),
    .B(net6583),
    .Y(_19458_));
 sg13g2_a21oi_1 _27877_ (.A1(net6583),
    .A2(_19457_),
    .Y(_00317_),
    .B1(_19458_));
 sg13g2_a22oi_1 _27878_ (.Y(_19459_),
    .B1(net6663),
    .B2(net1905),
    .A2(net6929),
    .A1(net2303));
 sg13g2_nor2_1 _27879_ (.A(net3398),
    .B(net6583),
    .Y(_19460_));
 sg13g2_a21oi_1 _27880_ (.A1(net6583),
    .A2(_19459_),
    .Y(_00318_),
    .B1(_19460_));
 sg13g2_a22oi_1 _27881_ (.Y(_19461_),
    .B1(net6663),
    .B2(net1339),
    .A2(net6931),
    .A1(net1974));
 sg13g2_nor2_1 _27882_ (.A(net3570),
    .B(net6585),
    .Y(_19462_));
 sg13g2_a21oi_1 _27883_ (.A1(net6585),
    .A2(_19461_),
    .Y(_00319_),
    .B1(_19462_));
 sg13g2_a22oi_1 _27884_ (.Y(_19463_),
    .B1(net6663),
    .B2(net3283),
    .A2(net6931),
    .A1(net2291));
 sg13g2_nor2_1 _27885_ (.A(net3508),
    .B(net6585),
    .Y(_19464_));
 sg13g2_a21oi_1 _27886_ (.A1(net6585),
    .A2(_19463_),
    .Y(_00320_),
    .B1(_19464_));
 sg13g2_a22oi_1 _27887_ (.Y(_19465_),
    .B1(net6659),
    .B2(net1673),
    .A2(net6923),
    .A1(net3379));
 sg13g2_nor2_1 _27888_ (.A(net3615),
    .B(net6574),
    .Y(_19466_));
 sg13g2_a21oi_1 _27889_ (.A1(net6574),
    .A2(_19465_),
    .Y(_00321_),
    .B1(_19466_));
 sg13g2_a22oi_1 _27890_ (.Y(_19467_),
    .B1(net6659),
    .B2(net3067),
    .A2(net6931),
    .A1(net3487));
 sg13g2_nor2_1 _27891_ (.A(net3552),
    .B(net6573),
    .Y(_19468_));
 sg13g2_a21oi_1 _27892_ (.A1(net6587),
    .A2(_19467_),
    .Y(_00322_),
    .B1(_19468_));
 sg13g2_a22oi_1 _27893_ (.Y(_19469_),
    .B1(net6659),
    .B2(net1881),
    .A2(net6923),
    .A1(net3429));
 sg13g2_nor2_1 _27894_ (.A(net3479),
    .B(net6574),
    .Y(_19470_));
 sg13g2_a21oi_1 _27895_ (.A1(net6574),
    .A2(_19469_),
    .Y(_00323_),
    .B1(_19470_));
 sg13g2_a22oi_1 _27896_ (.Y(_19471_),
    .B1(net6659),
    .B2(net1273),
    .A2(net6923),
    .A1(net3357));
 sg13g2_nor2_1 _27897_ (.A(net3573),
    .B(net6573),
    .Y(_19472_));
 sg13g2_a21oi_1 _27898_ (.A1(net6573),
    .A2(_19471_),
    .Y(_00324_),
    .B1(_19472_));
 sg13g2_a22oi_1 _27899_ (.Y(_19473_),
    .B1(net6660),
    .B2(net2582),
    .A2(net6923),
    .A1(net3449));
 sg13g2_nor2_1 _27900_ (.A(net3516),
    .B(net6563),
    .Y(_19474_));
 sg13g2_a21oi_1 _27901_ (.A1(net6573),
    .A2(_19473_),
    .Y(_00325_),
    .B1(_19474_));
 sg13g2_a22oi_1 _27902_ (.Y(_19475_),
    .B1(net6660),
    .B2(net1799),
    .A2(net6924),
    .A1(net3398));
 sg13g2_nor2_1 _27903_ (.A(net3572),
    .B(net6573),
    .Y(_19476_));
 sg13g2_a21oi_1 _27904_ (.A1(net6573),
    .A2(_19475_),
    .Y(_00326_),
    .B1(_19476_));
 sg13g2_a22oi_1 _27905_ (.Y(_19477_),
    .B1(net6659),
    .B2(net1847),
    .A2(net6923),
    .A1(\shift_reg[144] ));
 sg13g2_nor2_1 _27906_ (.A(net3256),
    .B(net6573),
    .Y(_19478_));
 sg13g2_a21oi_1 _27907_ (.A1(net6573),
    .A2(_19477_),
    .Y(_00327_),
    .B1(_19478_));
 sg13g2_a22oi_1 _27908_ (.Y(_19479_),
    .B1(net6659),
    .B2(net1232),
    .A2(net6923),
    .A1(\shift_reg[145] ));
 sg13g2_nor2_1 _27909_ (.A(net3098),
    .B(net6563),
    .Y(_19480_));
 sg13g2_a21oi_1 _27910_ (.A1(net6563),
    .A2(_19479_),
    .Y(_00328_),
    .B1(_19480_));
 sg13g2_a22oi_1 _27911_ (.Y(_19481_),
    .B1(net6659),
    .B2(net1741),
    .A2(net6923),
    .A1(\shift_reg[146] ));
 sg13g2_nor2_1 _27912_ (.A(net3332),
    .B(net6564),
    .Y(_19482_));
 sg13g2_a21oi_1 _27913_ (.A1(net6563),
    .A2(_19481_),
    .Y(_00329_),
    .B1(_19482_));
 sg13g2_a22oi_1 _27914_ (.Y(_19483_),
    .B1(net6659),
    .B2(net1230),
    .A2(net6923),
    .A1(\shift_reg[147] ));
 sg13g2_nor2_1 _27915_ (.A(net2750),
    .B(net6562),
    .Y(_19484_));
 sg13g2_a21oi_1 _27916_ (.A1(net6562),
    .A2(_19483_),
    .Y(_00330_),
    .B1(_19484_));
 sg13g2_a22oi_1 _27917_ (.Y(_19485_),
    .B1(net6655),
    .B2(net2717),
    .A2(net6919),
    .A1(\shift_reg[148] ));
 sg13g2_nor2_1 _27918_ (.A(net3381),
    .B(net6564),
    .Y(_19486_));
 sg13g2_a21oi_1 _27919_ (.A1(net6563),
    .A2(_19485_),
    .Y(_00331_),
    .B1(_19486_));
 sg13g2_a22oi_1 _27920_ (.Y(_19487_),
    .B1(net6655),
    .B2(net1458),
    .A2(net6919),
    .A1(\shift_reg[149] ));
 sg13g2_nor2_1 _27921_ (.A(net2898),
    .B(net6563),
    .Y(_19488_));
 sg13g2_a21oi_1 _27922_ (.A1(net6563),
    .A2(_19487_),
    .Y(_00332_),
    .B1(_19488_));
 sg13g2_a22oi_1 _27923_ (.Y(_19489_),
    .B1(net6655),
    .B2(net1620),
    .A2(net6919),
    .A1(\shift_reg[150] ));
 sg13g2_nor2_1 _27924_ (.A(net3301),
    .B(net6560),
    .Y(_19490_));
 sg13g2_a21oi_1 _27925_ (.A1(net6561),
    .A2(_19489_),
    .Y(_00333_),
    .B1(_19490_));
 sg13g2_a22oi_1 _27926_ (.Y(_19491_),
    .B1(net6655),
    .B2(net1441),
    .A2(net6919),
    .A1(\shift_reg[151] ));
 sg13g2_nor2_1 _27927_ (.A(net3329),
    .B(net6564),
    .Y(_19492_));
 sg13g2_a21oi_1 _27928_ (.A1(net6563),
    .A2(_19491_),
    .Y(_00334_),
    .B1(_19492_));
 sg13g2_a22oi_1 _27929_ (.Y(_19493_),
    .B1(net6654),
    .B2(net1178),
    .A2(net6918),
    .A1(net3256));
 sg13g2_nor2_1 _27930_ (.A(net3447),
    .B(net6562),
    .Y(_19494_));
 sg13g2_a21oi_1 _27931_ (.A1(net6562),
    .A2(_19493_),
    .Y(_00335_),
    .B1(_19494_));
 sg13g2_a22oi_1 _27932_ (.Y(_19495_),
    .B1(net6654),
    .B2(net3212),
    .A2(net6918),
    .A1(net3098));
 sg13g2_nor2_1 _27933_ (.A(net3288),
    .B(net6561),
    .Y(_19496_));
 sg13g2_a21oi_1 _27934_ (.A1(net6561),
    .A2(_19495_),
    .Y(_00336_),
    .B1(_19496_));
 sg13g2_a22oi_1 _27935_ (.Y(_19497_),
    .B1(net6654),
    .B2(net1703),
    .A2(net6919),
    .A1(\shift_reg[154] ));
 sg13g2_nor2_1 _27936_ (.A(net3248),
    .B(net6562),
    .Y(_19498_));
 sg13g2_a21oi_1 _27937_ (.A1(net6561),
    .A2(_19497_),
    .Y(_00337_),
    .B1(_19498_));
 sg13g2_a22oi_1 _27938_ (.Y(_19499_),
    .B1(net6654),
    .B2(net1297),
    .A2(net6919),
    .A1(net2750));
 sg13g2_nor2_1 _27939_ (.A(net3437),
    .B(net6562),
    .Y(_19500_));
 sg13g2_a21oi_1 _27940_ (.A1(net6561),
    .A2(_19499_),
    .Y(_00338_),
    .B1(_19500_));
 sg13g2_a22oi_1 _27941_ (.Y(_19501_),
    .B1(net6653),
    .B2(net1437),
    .A2(net6918),
    .A1(\shift_reg[156] ));
 sg13g2_nor2_1 _27942_ (.A(net3107),
    .B(net6562),
    .Y(_19502_));
 sg13g2_a21oi_1 _27943_ (.A1(net6560),
    .A2(_19501_),
    .Y(_00339_),
    .B1(_19502_));
 sg13g2_a22oi_1 _27944_ (.Y(_19503_),
    .B1(net6654),
    .B2(net1260),
    .A2(net6918),
    .A1(net2898));
 sg13g2_nor2_1 _27945_ (.A(net3339),
    .B(net6561),
    .Y(_19504_));
 sg13g2_a21oi_1 _27946_ (.A1(net6561),
    .A2(_19503_),
    .Y(_00340_),
    .B1(_19504_));
 sg13g2_a22oi_1 _27947_ (.Y(_19505_),
    .B1(net6652),
    .B2(net1583),
    .A2(net6918),
    .A1(net3301));
 sg13g2_nor2_1 _27948_ (.A(net3541),
    .B(net6559),
    .Y(_19506_));
 sg13g2_a21oi_1 _27949_ (.A1(net6559),
    .A2(_19505_),
    .Y(_00341_),
    .B1(_19506_));
 sg13g2_a22oi_1 _27950_ (.Y(_19507_),
    .B1(net6653),
    .B2(net2067),
    .A2(net6918),
    .A1(\shift_reg[159] ));
 sg13g2_nor2_1 _27951_ (.A(net3242),
    .B(net6560),
    .Y(_19508_));
 sg13g2_a21oi_1 _27952_ (.A1(net6560),
    .A2(_19507_),
    .Y(_00342_),
    .B1(_19508_));
 sg13g2_a22oi_1 _27953_ (.Y(_19509_),
    .B1(net6653),
    .B2(net2184),
    .A2(net6918),
    .A1(net3447));
 sg13g2_nor2_1 _27954_ (.A(net3559),
    .B(net6560),
    .Y(_19510_));
 sg13g2_a21oi_1 _27955_ (.A1(net6560),
    .A2(_19509_),
    .Y(_00343_),
    .B1(_19510_));
 sg13g2_a22oi_1 _27956_ (.Y(_19511_),
    .B1(net6653),
    .B2(net3486),
    .A2(net6918),
    .A1(net3288));
 sg13g2_nor2_1 _27957_ (.A(net3529),
    .B(net6560),
    .Y(_19512_));
 sg13g2_a21oi_1 _27958_ (.A1(net6560),
    .A2(_19511_),
    .Y(_00344_),
    .B1(_19512_));
 sg13g2_a22oi_1 _27959_ (.Y(_19513_),
    .B1(net6652),
    .B2(net1759),
    .A2(net6916),
    .A1(net3248));
 sg13g2_nor2_1 _27960_ (.A(net3489),
    .B(net6565),
    .Y(_19514_));
 sg13g2_a21oi_1 _27961_ (.A1(net6559),
    .A2(_19513_),
    .Y(_00345_),
    .B1(_19514_));
 sg13g2_a22oi_1 _27962_ (.Y(_19515_),
    .B1(net6652),
    .B2(net1227),
    .A2(net6916),
    .A1(\shift_reg[163] ));
 sg13g2_nor2_1 _27963_ (.A(net3351),
    .B(net6559),
    .Y(_19516_));
 sg13g2_a21oi_1 _27964_ (.A1(net6559),
    .A2(_19515_),
    .Y(_00346_),
    .B1(_19516_));
 sg13g2_a22oi_1 _27965_ (.Y(_19517_),
    .B1(net6652),
    .B2(net1210),
    .A2(net6916),
    .A1(net3107));
 sg13g2_nor2_1 _27966_ (.A(net3415),
    .B(net6556),
    .Y(_19518_));
 sg13g2_a21oi_1 _27967_ (.A1(net6559),
    .A2(_19517_),
    .Y(_00347_),
    .B1(_19518_));
 sg13g2_a22oi_1 _27968_ (.Y(_19519_),
    .B1(net6652),
    .B2(net1479),
    .A2(net6916),
    .A1(net3339));
 sg13g2_nor2_1 _27969_ (.A(net3545),
    .B(net6557),
    .Y(_19520_));
 sg13g2_a21oi_1 _27970_ (.A1(net6558),
    .A2(_19519_),
    .Y(_00348_),
    .B1(_19520_));
 sg13g2_a22oi_1 _27971_ (.Y(_19521_),
    .B1(net6652),
    .B2(net1846),
    .A2(net6917),
    .A1(net3541));
 sg13g2_nor2_1 _27972_ (.A(net3597),
    .B(net6557),
    .Y(_19522_));
 sg13g2_a21oi_1 _27973_ (.A1(net6558),
    .A2(_19521_),
    .Y(_00349_),
    .B1(_19522_));
 sg13g2_a22oi_1 _27974_ (.Y(_19523_),
    .B1(net6652),
    .B2(net1459),
    .A2(net6917),
    .A1(net3242));
 sg13g2_nor2_1 _27975_ (.A(net3623),
    .B(net6557),
    .Y(_19524_));
 sg13g2_a21oi_1 _27976_ (.A1(net6557),
    .A2(_19523_),
    .Y(_00350_),
    .B1(_19524_));
 sg13g2_a22oi_1 _27977_ (.Y(_19525_),
    .B1(net6652),
    .B2(net1856),
    .A2(net6917),
    .A1(\shift_reg[168] ));
 sg13g2_nor2_1 _27978_ (.A(net3521),
    .B(net6558),
    .Y(_19526_));
 sg13g2_a21oi_1 _27979_ (.A1(net6558),
    .A2(_19525_),
    .Y(_00351_),
    .B1(_19526_));
 sg13g2_a22oi_1 _27980_ (.Y(_19527_),
    .B1(net6649),
    .B2(net1959),
    .A2(net6916),
    .A1(\shift_reg[169] ));
 sg13g2_nor2_1 _27981_ (.A(net3281),
    .B(net6557),
    .Y(_19528_));
 sg13g2_a21oi_1 _27982_ (.A1(net6557),
    .A2(_19527_),
    .Y(_00352_),
    .B1(_19528_));
 sg13g2_a22oi_1 _27983_ (.Y(_19529_),
    .B1(net6649),
    .B2(net2176),
    .A2(net6916),
    .A1(net3489));
 sg13g2_nor2_1 _27984_ (.A(net3557),
    .B(net6554),
    .Y(_19530_));
 sg13g2_a21oi_1 _27985_ (.A1(net6554),
    .A2(_19529_),
    .Y(_00353_),
    .B1(_19530_));
 sg13g2_a22oi_1 _27986_ (.Y(_19531_),
    .B1(net6649),
    .B2(net1261),
    .A2(net6916),
    .A1(\shift_reg[171] ));
 sg13g2_nor2_1 _27987_ (.A(net2793),
    .B(net6554),
    .Y(_19532_));
 sg13g2_a21oi_1 _27988_ (.A1(net6554),
    .A2(_19531_),
    .Y(_00354_),
    .B1(_19532_));
 sg13g2_a22oi_1 _27989_ (.Y(_19533_),
    .B1(net6649),
    .B2(net1440),
    .A2(net6914),
    .A1(\shift_reg[172] ));
 sg13g2_nor2_1 _27990_ (.A(net3310),
    .B(net6550),
    .Y(_19534_));
 sg13g2_a21oi_1 _27991_ (.A1(net6554),
    .A2(_19533_),
    .Y(_00355_),
    .B1(_19534_));
 sg13g2_a22oi_1 _27992_ (.Y(_19535_),
    .B1(net6649),
    .B2(net1219),
    .A2(net6916),
    .A1(\shift_reg[173] ));
 sg13g2_nor2_1 _27993_ (.A(net3498),
    .B(net6557),
    .Y(_19536_));
 sg13g2_a21oi_1 _27994_ (.A1(net6557),
    .A2(_19535_),
    .Y(_00356_),
    .B1(_19536_));
 sg13g2_a22oi_1 _27995_ (.Y(_19537_),
    .B1(net6649),
    .B2(net1819),
    .A2(net6914),
    .A1(\shift_reg[174] ));
 sg13g2_nor2_1 _27996_ (.A(net3223),
    .B(net6553),
    .Y(_19538_));
 sg13g2_a21oi_1 _27997_ (.A1(net6554),
    .A2(_19537_),
    .Y(_00357_),
    .B1(_19538_));
 sg13g2_a22oi_1 _27998_ (.Y(_19539_),
    .B1(net6650),
    .B2(net2065),
    .A2(net6914),
    .A1(\shift_reg[175] ));
 sg13g2_nor2_1 _27999_ (.A(net3177),
    .B(net6553),
    .Y(_19540_));
 sg13g2_a21oi_1 _28000_ (.A1(net6553),
    .A2(_19539_),
    .Y(_00358_),
    .B1(_19540_));
 sg13g2_a22oi_1 _28001_ (.Y(_19541_),
    .B1(net6649),
    .B2(net1922),
    .A2(net6913),
    .A1(\shift_reg[176] ));
 sg13g2_nor2_1 _28002_ (.A(net2442),
    .B(net6545),
    .Y(_19542_));
 sg13g2_a21oi_1 _28003_ (.A1(net6545),
    .A2(_19541_),
    .Y(_00359_),
    .B1(_19542_));
 sg13g2_a22oi_1 _28004_ (.Y(_19543_),
    .B1(net6649),
    .B2(net1892),
    .A2(net6913),
    .A1(\shift_reg[177] ));
 sg13g2_nor2_1 _28005_ (.A(net2282),
    .B(net6545),
    .Y(_19544_));
 sg13g2_a21oi_1 _28006_ (.A1(net6545),
    .A2(_19543_),
    .Y(_00360_),
    .B1(_19544_));
 sg13g2_a22oi_1 _28007_ (.Y(_19545_),
    .B1(net6647),
    .B2(net2011),
    .A2(net6912),
    .A1(\shift_reg[178] ));
 sg13g2_nor2_1 _28008_ (.A(net2678),
    .B(net6544),
    .Y(_19546_));
 sg13g2_a21oi_1 _28009_ (.A1(net6543),
    .A2(_19545_),
    .Y(_00361_),
    .B1(_19546_));
 sg13g2_a22oi_1 _28010_ (.Y(_19547_),
    .B1(net6647),
    .B2(\inv_result[171] ),
    .A2(net6913),
    .A1(\shift_reg[179] ));
 sg13g2_nor2_1 _28011_ (.A(net2293),
    .B(net6545),
    .Y(_19548_));
 sg13g2_a21oi_1 _28012_ (.A1(net6545),
    .A2(_19547_),
    .Y(_00362_),
    .B1(_19548_));
 sg13g2_a22oi_1 _28013_ (.Y(_19549_),
    .B1(net6647),
    .B2(net1197),
    .A2(net6912),
    .A1(net3310));
 sg13g2_nor2_1 _28014_ (.A(net3518),
    .B(net6548),
    .Y(_19550_));
 sg13g2_a21oi_1 _28015_ (.A1(net6548),
    .A2(_19549_),
    .Y(_00363_),
    .B1(_19550_));
 sg13g2_a22oi_1 _28016_ (.Y(_19551_),
    .B1(net6647),
    .B2(net1292),
    .A2(net6912),
    .A1(net3498));
 sg13g2_nor2_1 _28017_ (.A(net3548),
    .B(net6550),
    .Y(_19552_));
 sg13g2_a21oi_1 _28018_ (.A1(net6550),
    .A2(_19551_),
    .Y(_00364_),
    .B1(_19552_));
 sg13g2_a22oi_1 _28019_ (.Y(_19553_),
    .B1(net6645),
    .B2(\inv_result[174] ),
    .A2(net6911),
    .A1(\shift_reg[182] ));
 sg13g2_nor2_1 _28020_ (.A(net2233),
    .B(net6543),
    .Y(_19554_));
 sg13g2_a21oi_1 _28021_ (.A1(net6543),
    .A2(_19553_),
    .Y(_00365_),
    .B1(_19554_));
 sg13g2_a22oi_1 _28022_ (.Y(_19555_),
    .B1(net6647),
    .B2(net1887),
    .A2(net6911),
    .A1(net3177));
 sg13g2_nor2_1 _28023_ (.A(net3512),
    .B(net6548),
    .Y(_19556_));
 sg13g2_a21oi_1 _28024_ (.A1(net6548),
    .A2(_19555_),
    .Y(_00366_),
    .B1(_19556_));
 sg13g2_a22oi_1 _28025_ (.Y(_19557_),
    .B1(net6643),
    .B2(net1530),
    .A2(net6910),
    .A1(net2442));
 sg13g2_nor2_1 _28026_ (.A(net2847),
    .B(net6544),
    .Y(_19558_));
 sg13g2_a21oi_1 _28027_ (.A1(net6544),
    .A2(_19557_),
    .Y(_00367_),
    .B1(_19558_));
 sg13g2_a22oi_1 _28028_ (.Y(_19559_),
    .B1(net6643),
    .B2(net2012),
    .A2(net6910),
    .A1(\shift_reg[185] ));
 sg13g2_nor2_1 _28029_ (.A(net2211),
    .B(net6538),
    .Y(_19560_));
 sg13g2_a21oi_1 _28030_ (.A1(net6543),
    .A2(_19559_),
    .Y(_00368_),
    .B1(_19560_));
 sg13g2_a22oi_1 _28031_ (.Y(_19561_),
    .B1(net6643),
    .B2(net1662),
    .A2(net6909),
    .A1(\shift_reg[186] ));
 sg13g2_nor2_1 _28032_ (.A(net2321),
    .B(net6539),
    .Y(_19562_));
 sg13g2_a21oi_1 _28033_ (.A1(net6538),
    .A2(_19561_),
    .Y(_00369_),
    .B1(_19562_));
 sg13g2_a22oi_1 _28034_ (.Y(_19563_),
    .B1(net6643),
    .B2(\inv_result[179] ),
    .A2(net6909),
    .A1(net2293));
 sg13g2_nor2_1 _28035_ (.A(net2351),
    .B(net6543),
    .Y(_19564_));
 sg13g2_a21oi_1 _28036_ (.A1(net6543),
    .A2(_19563_),
    .Y(_00370_),
    .B1(_19564_));
 sg13g2_a22oi_1 _28037_ (.Y(_19565_),
    .B1(net6642),
    .B2(net1882),
    .A2(net6909),
    .A1(\shift_reg[188] ));
 sg13g2_nor2_1 _28038_ (.A(net2604),
    .B(net6543),
    .Y(_19566_));
 sg13g2_a21oi_1 _28039_ (.A1(net6543),
    .A2(_19565_),
    .Y(_00371_),
    .B1(_19566_));
 sg13g2_a22oi_1 _28040_ (.Y(_19567_),
    .B1(net6642),
    .B2(net1710),
    .A2(net6909),
    .A1(\shift_reg[189] ));
 sg13g2_nor2_1 _28041_ (.A(net2535),
    .B(net6541),
    .Y(_19568_));
 sg13g2_a21oi_1 _28042_ (.A1(net6538),
    .A2(_19567_),
    .Y(_00372_),
    .B1(_19568_));
 sg13g2_a22oi_1 _28043_ (.Y(_19569_),
    .B1(net6642),
    .B2(net1247),
    .A2(net6909),
    .A1(net2233));
 sg13g2_nor2_1 _28044_ (.A(net2625),
    .B(net6538),
    .Y(_19570_));
 sg13g2_a21oi_1 _28045_ (.A1(net6538),
    .A2(_19569_),
    .Y(_00373_),
    .B1(_19570_));
 sg13g2_a22oi_1 _28046_ (.Y(_19571_),
    .B1(net6643),
    .B2(net1677),
    .A2(net6909),
    .A1(\shift_reg[191] ));
 sg13g2_nor2_1 _28047_ (.A(net2556),
    .B(net6541),
    .Y(_19572_));
 sg13g2_a21oi_1 _28048_ (.A1(net6538),
    .A2(_19571_),
    .Y(_00374_),
    .B1(_19572_));
 sg13g2_a22oi_1 _28049_ (.Y(_19573_),
    .B1(net6642),
    .B2(net1938),
    .A2(net6909),
    .A1(net2847));
 sg13g2_nor2_1 _28050_ (.A(net2849),
    .B(net6539),
    .Y(_19574_));
 sg13g2_a21oi_1 _28051_ (.A1(net6539),
    .A2(_19573_),
    .Y(_00375_),
    .B1(_19574_));
 sg13g2_a22oi_1 _28052_ (.Y(_19575_),
    .B1(net6642),
    .B2(net1355),
    .A2(net6906),
    .A1(net2211));
 sg13g2_nor2_1 _28053_ (.A(net2784),
    .B(net6539),
    .Y(_19576_));
 sg13g2_a21oi_1 _28054_ (.A1(net6539),
    .A2(_19575_),
    .Y(_00376_),
    .B1(_19576_));
 sg13g2_a22oi_1 _28055_ (.Y(_19577_),
    .B1(net6641),
    .B2(net1853),
    .A2(net6906),
    .A1(net2321));
 sg13g2_nor2_1 _28056_ (.A(net2957),
    .B(net6538),
    .Y(_19578_));
 sg13g2_a21oi_1 _28057_ (.A1(net6538),
    .A2(_19577_),
    .Y(_00377_),
    .B1(_19578_));
 sg13g2_a22oi_1 _28058_ (.Y(_19579_),
    .B1(net6642),
    .B2(net1228),
    .A2(net6909),
    .A1(\shift_reg[195] ));
 sg13g2_nor2_1 _28059_ (.A(net2277),
    .B(net6539),
    .Y(_19580_));
 sg13g2_a21oi_1 _28060_ (.A1(net6539),
    .A2(_19579_),
    .Y(_00378_),
    .B1(_19580_));
 sg13g2_a22oi_1 _28061_ (.Y(_19581_),
    .B1(net6641),
    .B2(net1205),
    .A2(net6906),
    .A1(net2604));
 sg13g2_nor2_1 _28062_ (.A(net3102),
    .B(net6540),
    .Y(_19582_));
 sg13g2_a21oi_1 _28063_ (.A1(net6540),
    .A2(_19581_),
    .Y(_00379_),
    .B1(_19582_));
 sg13g2_a22oi_1 _28064_ (.Y(_19583_),
    .B1(net6642),
    .B2(net1464),
    .A2(net6907),
    .A1(\shift_reg[197] ));
 sg13g2_nor2_1 _28065_ (.A(net2248),
    .B(net6540),
    .Y(_19584_));
 sg13g2_a21oi_1 _28066_ (.A1(net6540),
    .A2(_19583_),
    .Y(_00380_),
    .B1(_19584_));
 sg13g2_a22oi_1 _28067_ (.Y(_19585_),
    .B1(net6641),
    .B2(net2125),
    .A2(net6907),
    .A1(\shift_reg[198] ));
 sg13g2_nor2_1 _28068_ (.A(net2507),
    .B(net6540),
    .Y(_19586_));
 sg13g2_a21oi_1 _28069_ (.A1(net6540),
    .A2(_19585_),
    .Y(_00381_),
    .B1(_19586_));
 sg13g2_a22oi_1 _28070_ (.Y(_19587_),
    .B1(net6642),
    .B2(net1985),
    .A2(net6907),
    .A1(net2556));
 sg13g2_nor2_1 _28071_ (.A(net2755),
    .B(net6540),
    .Y(_19588_));
 sg13g2_a21oi_1 _28072_ (.A1(net6540),
    .A2(_19587_),
    .Y(_00382_),
    .B1(_19588_));
 sg13g2_a22oi_1 _28073_ (.Y(_19589_),
    .B1(net6639),
    .B2(net2285),
    .A2(net6905),
    .A1(net2849));
 sg13g2_nor2_1 _28074_ (.A(net3026),
    .B(net6535),
    .Y(_19590_));
 sg13g2_a21oi_1 _28075_ (.A1(net6533),
    .A2(_19589_),
    .Y(_00383_),
    .B1(_19590_));
 sg13g2_a22oi_1 _28076_ (.Y(_19591_),
    .B1(net6639),
    .B2(net2213),
    .A2(net6905),
    .A1(\shift_reg[201] ));
 sg13g2_nor2_1 _28077_ (.A(net2546),
    .B(net6533),
    .Y(_19592_));
 sg13g2_a21oi_1 _28078_ (.A1(net6533),
    .A2(_19591_),
    .Y(_00384_),
    .B1(_19592_));
 sg13g2_a22oi_1 _28079_ (.Y(_19593_),
    .B1(net6639),
    .B2(net2051),
    .A2(net6904),
    .A1(net2957));
 sg13g2_nor2_1 _28080_ (.A(net3202),
    .B(net6535),
    .Y(_19594_));
 sg13g2_a21oi_1 _28081_ (.A1(net6535),
    .A2(_19593_),
    .Y(_00385_),
    .B1(_19594_));
 sg13g2_a22oi_1 _28082_ (.Y(_19595_),
    .B1(net6641),
    .B2(net1674),
    .A2(net6904),
    .A1(net2277));
 sg13g2_nor2_1 _28083_ (.A(net3024),
    .B(net6533),
    .Y(_19596_));
 sg13g2_a21oi_1 _28084_ (.A1(net6534),
    .A2(_19595_),
    .Y(_00386_),
    .B1(_19596_));
 sg13g2_a22oi_1 _28085_ (.Y(_19597_),
    .B1(net6638),
    .B2(net1859),
    .A2(net6904),
    .A1(\shift_reg[204] ));
 sg13g2_nor2_1 _28086_ (.A(net3002),
    .B(net6534),
    .Y(_19598_));
 sg13g2_a21oi_1 _28087_ (.A1(net6534),
    .A2(_19597_),
    .Y(_00387_),
    .B1(_19598_));
 sg13g2_a22oi_1 _28088_ (.Y(_19599_),
    .B1(net6639),
    .B2(net2001),
    .A2(net6904),
    .A1(net2248));
 sg13g2_nor2_1 _28089_ (.A(net3410),
    .B(net6535),
    .Y(_19600_));
 sg13g2_a21oi_1 _28090_ (.A1(net6535),
    .A2(_19599_),
    .Y(_00388_),
    .B1(_19600_));
 sg13g2_a22oi_1 _28091_ (.Y(_19601_),
    .B1(net6639),
    .B2(net1198),
    .A2(net6905),
    .A1(net2507));
 sg13g2_nor2_1 _28092_ (.A(net2698),
    .B(net6515),
    .Y(_19602_));
 sg13g2_a21oi_1 _28093_ (.A1(net6515),
    .A2(_19601_),
    .Y(_00389_),
    .B1(_19602_));
 sg13g2_a22oi_1 _28094_ (.Y(_19603_),
    .B1(net6638),
    .B2(net2013),
    .A2(net6904),
    .A1(net2755));
 sg13g2_nor2_1 _28095_ (.A(net3115),
    .B(net6534),
    .Y(_19604_));
 sg13g2_a21oi_1 _28096_ (.A1(net6534),
    .A2(_19603_),
    .Y(_00390_),
    .B1(_19604_));
 sg13g2_a22oi_1 _28097_ (.Y(_19605_),
    .B1(net6638),
    .B2(net2187),
    .A2(net6904),
    .A1(net3026));
 sg13g2_nor2_1 _28098_ (.A(net3470),
    .B(net6533),
    .Y(_19606_));
 sg13g2_a21oi_1 _28099_ (.A1(net6533),
    .A2(_19605_),
    .Y(_00391_),
    .B1(_19606_));
 sg13g2_a22oi_1 _28100_ (.Y(_19607_),
    .B1(net6637),
    .B2(\inv_result[201] ),
    .A2(net6895),
    .A1(\shift_reg[209] ));
 sg13g2_nor2_1 _28101_ (.A(net2171),
    .B(net6516),
    .Y(_19608_));
 sg13g2_a21oi_1 _28102_ (.A1(net6516),
    .A2(_19607_),
    .Y(_00392_),
    .B1(_19608_));
 sg13g2_a22oi_1 _28103_ (.Y(_19609_),
    .B1(net6638),
    .B2(net1932),
    .A2(net6905),
    .A1(net3202));
 sg13g2_nor2_1 _28104_ (.A(net3519),
    .B(net6533),
    .Y(_19610_));
 sg13g2_a21oi_1 _28105_ (.A1(net6533),
    .A2(_19609_),
    .Y(_00393_),
    .B1(_19610_));
 sg13g2_a22oi_1 _28106_ (.Y(_19611_),
    .B1(net6638),
    .B2(\inv_result[203] ),
    .A2(net6905),
    .A1(\shift_reg[211] ));
 sg13g2_nor2_1 _28107_ (.A(net2728),
    .B(net6516),
    .Y(_19612_));
 sg13g2_a21oi_1 _28108_ (.A1(net6516),
    .A2(_19611_),
    .Y(_00394_),
    .B1(_19612_));
 sg13g2_a22oi_1 _28109_ (.Y(_19613_),
    .B1(net6638),
    .B2(net2096),
    .A2(net6904),
    .A1(\shift_reg[212] ));
 sg13g2_nor2_1 _28110_ (.A(net2961),
    .B(net6519),
    .Y(_19614_));
 sg13g2_a21oi_1 _28111_ (.A1(net6518),
    .A2(_19613_),
    .Y(_00395_),
    .B1(_19614_));
 sg13g2_a22oi_1 _28112_ (.Y(_19615_),
    .B1(net6638),
    .B2(net1237),
    .A2(net6904),
    .A1(\shift_reg[213] ));
 sg13g2_nor2_1 _28113_ (.A(net3234),
    .B(net6534),
    .Y(_19616_));
 sg13g2_a21oi_1 _28114_ (.A1(net6534),
    .A2(_19615_),
    .Y(_00396_),
    .B1(_19616_));
 sg13g2_a22oi_1 _28115_ (.Y(_19617_),
    .B1(net6637),
    .B2(net2757),
    .A2(net6895),
    .A1(net2698));
 sg13g2_nor2_1 _28116_ (.A(net3484),
    .B(net6515),
    .Y(_19618_));
 sg13g2_a21oi_1 _28117_ (.A1(net6515),
    .A2(_19617_),
    .Y(_00397_),
    .B1(_19618_));
 sg13g2_a22oi_1 _28118_ (.Y(_19619_),
    .B1(net6638),
    .B2(net2518),
    .A2(net6893),
    .A1(net3115));
 sg13g2_nor2_1 _28119_ (.A(net3395),
    .B(net6519),
    .Y(_19620_));
 sg13g2_a21oi_1 _28120_ (.A1(net6518),
    .A2(_19619_),
    .Y(_00398_),
    .B1(_19620_));
 sg13g2_a22oi_1 _28121_ (.Y(_19621_),
    .B1(net6637),
    .B2(net1291),
    .A2(net6894),
    .A1(\shift_reg[216] ));
 sg13g2_nor2_1 _28122_ (.A(net3432),
    .B(net6518),
    .Y(_19622_));
 sg13g2_a21oi_1 _28123_ (.A1(net6518),
    .A2(_19621_),
    .Y(_00399_),
    .B1(_19622_));
 sg13g2_a22oi_1 _28124_ (.Y(_19623_),
    .B1(net6637),
    .B2(net1984),
    .A2(net6895),
    .A1(net2171));
 sg13g2_nor2_1 _28125_ (.A(net3643),
    .B(net6516),
    .Y(_19624_));
 sg13g2_a21oi_1 _28126_ (.A1(net6516),
    .A2(_19623_),
    .Y(_00400_),
    .B1(_19624_));
 sg13g2_a22oi_1 _28127_ (.Y(_19625_),
    .B1(net6637),
    .B2(net1794),
    .A2(net6895),
    .A1(\shift_reg[218] ));
 sg13g2_nor2_1 _28128_ (.A(net3228),
    .B(net6515),
    .Y(_19626_));
 sg13g2_a21oi_1 _28129_ (.A1(net6519),
    .A2(_19625_),
    .Y(_00401_),
    .B1(_19626_));
 sg13g2_a22oi_1 _28130_ (.Y(_19627_),
    .B1(net6637),
    .B2(net1919),
    .A2(net6894),
    .A1(net2728));
 sg13g2_nor2_1 _28131_ (.A(net3076),
    .B(net6518),
    .Y(_19628_));
 sg13g2_a21oi_1 _28132_ (.A1(net6518),
    .A2(_19627_),
    .Y(_00402_),
    .B1(_19628_));
 sg13g2_a22oi_1 _28133_ (.Y(_19629_),
    .B1(net6640),
    .B2(net2078),
    .A2(net6894),
    .A1(net2961));
 sg13g2_nor2_1 _28134_ (.A(net3503),
    .B(net6519),
    .Y(_19630_));
 sg13g2_a21oi_1 _28135_ (.A1(net6518),
    .A2(_19629_),
    .Y(_00403_),
    .B1(_19630_));
 sg13g2_a22oi_1 _28136_ (.Y(_19631_),
    .B1(net6640),
    .B2(net1248),
    .A2(net6894),
    .A1(net3234));
 sg13g2_nor2_1 _28137_ (.A(net3622),
    .B(net6519),
    .Y(_19632_));
 sg13g2_a21oi_1 _28138_ (.A1(net6519),
    .A2(_19631_),
    .Y(_00404_),
    .B1(_19632_));
 sg13g2_o21ai_1 _28139_ (.B1(net6945),
    .Y(_19633_),
    .A1(trng_ready),
    .A2(net7161));
 sg13g2_a21oi_1 _28140_ (.A1(_18299_),
    .A2(net7150),
    .Y(_19634_),
    .B1(_19633_));
 sg13g2_a21oi_1 _28141_ (.A1(\shift_reg[222] ),
    .A2(net6896),
    .Y(_19635_),
    .B1(_19634_));
 sg13g2_nor2_1 _28142_ (.A(net2631),
    .B(net6521),
    .Y(_19636_));
 sg13g2_a21oi_1 _28143_ (.A1(net6521),
    .A2(_19635_),
    .Y(_00405_),
    .B1(_19636_));
 sg13g2_a21oi_1 _28144_ (.A1(net3172),
    .A2(net7155),
    .Y(_19637_),
    .B1(net6893));
 sg13g2_o21ai_1 _28145_ (.B1(_19637_),
    .Y(_19638_),
    .A1(_18265_),
    .A2(net7155));
 sg13g2_o21ai_1 _28146_ (.B1(_19638_),
    .Y(_19639_),
    .A1(\shift_reg[223] ),
    .A2(net6942));
 sg13g2_nor2_1 _28147_ (.A(net3318),
    .B(net6517),
    .Y(_19640_));
 sg13g2_a21oi_1 _28148_ (.A1(net6517),
    .A2(_19639_),
    .Y(_00406_),
    .B1(_19640_));
 sg13g2_o21ai_1 _28149_ (.B1(net6942),
    .Y(_19641_),
    .A1(net1233),
    .A2(net7155));
 sg13g2_a21oi_1 _28150_ (.A1(_18301_),
    .A2(net7154),
    .Y(_19642_),
    .B1(_19641_));
 sg13g2_a21oi_1 _28151_ (.A1(\shift_reg[224] ),
    .A2(net6893),
    .Y(_19643_),
    .B1(_19642_));
 sg13g2_nor2_1 _28152_ (.A(net2519),
    .B(net6514),
    .Y(_19644_));
 sg13g2_a21oi_1 _28153_ (.A1(net6514),
    .A2(_19643_),
    .Y(_00407_),
    .B1(_19644_));
 sg13g2_o21ai_1 _28154_ (.B1(net6942),
    .Y(_19645_),
    .A1(\inv_cycles[1] ),
    .A2(net7155));
 sg13g2_a21oi_1 _28155_ (.A1(_18300_),
    .A2(net7154),
    .Y(_19646_),
    .B1(_19645_));
 sg13g2_a21oi_1 _28156_ (.A1(\shift_reg[225] ),
    .A2(net6892),
    .Y(_19647_),
    .B1(_19646_));
 sg13g2_nor2_1 _28157_ (.A(net2174),
    .B(net6514),
    .Y(_19648_));
 sg13g2_a21oi_1 _28158_ (.A1(net6514),
    .A2(_19647_),
    .Y(_00408_),
    .B1(_19648_));
 sg13g2_o21ai_1 _28159_ (.B1(net6942),
    .Y(_19649_),
    .A1(net2304),
    .A2(net7154));
 sg13g2_a21oi_1 _28160_ (.A1(_18302_),
    .A2(net7154),
    .Y(_19650_),
    .B1(_19649_));
 sg13g2_a21oi_1 _28161_ (.A1(\shift_reg[226] ),
    .A2(net6893),
    .Y(_19651_),
    .B1(_19650_));
 sg13g2_nor2_1 _28162_ (.A(net2742),
    .B(net6517),
    .Y(_19652_));
 sg13g2_a21oi_1 _28163_ (.A1(net6517),
    .A2(_19651_),
    .Y(_00409_),
    .B1(_19652_));
 sg13g2_a21oi_1 _28164_ (.A1(net1224),
    .A2(net7154),
    .Y(_19653_),
    .B1(net6893));
 sg13g2_o21ai_1 _28165_ (.B1(_19653_),
    .Y(_19654_),
    .A1(_18339_),
    .A2(net7154));
 sg13g2_o21ai_1 _28166_ (.B1(_19654_),
    .Y(_19655_),
    .A1(\shift_reg[227] ),
    .A2(net6943));
 sg13g2_nor2_1 _28167_ (.A(net2800),
    .B(net6517),
    .Y(_19656_));
 sg13g2_a21oi_1 _28168_ (.A1(net6517),
    .A2(_19655_),
    .Y(_00410_),
    .B1(_19656_));
 sg13g2_o21ai_1 _28169_ (.B1(net6943),
    .Y(_19657_),
    .A1(net1203),
    .A2(net7154));
 sg13g2_a21oi_1 _28170_ (.A1(_18304_),
    .A2(net7154),
    .Y(_19658_),
    .B1(_19657_));
 sg13g2_a21oi_1 _28171_ (.A1(\shift_reg[228] ),
    .A2(net6891),
    .Y(_19659_),
    .B1(_19658_));
 sg13g2_nor2_1 _28172_ (.A(net2246),
    .B(net6513),
    .Y(_19660_));
 sg13g2_a21oi_1 _28173_ (.A1(net6513),
    .A2(_19659_),
    .Y(_00411_),
    .B1(_19660_));
 sg13g2_o21ai_1 _28174_ (.B1(net6942),
    .Y(_19661_),
    .A1(net1188),
    .A2(net7156));
 sg13g2_a21oi_1 _28175_ (.A1(_18303_),
    .A2(net7156),
    .Y(_19662_),
    .B1(_19661_));
 sg13g2_a21oi_1 _28176_ (.A1(\shift_reg[229] ),
    .A2(net6893),
    .Y(_19663_),
    .B1(_19662_));
 sg13g2_nor2_1 _28177_ (.A(net3262),
    .B(net6520),
    .Y(_19664_));
 sg13g2_a21oi_1 _28178_ (.A1(net6520),
    .A2(_19663_),
    .Y(_00412_),
    .B1(_19664_));
 sg13g2_o21ai_1 _28179_ (.B1(net6942),
    .Y(_19665_),
    .A1(net1878),
    .A2(net7156));
 sg13g2_a21oi_1 _28180_ (.A1(_18306_),
    .A2(net7156),
    .Y(_19666_),
    .B1(_19665_));
 sg13g2_a21oi_1 _28181_ (.A1(\shift_reg[230] ),
    .A2(net6891),
    .Y(_19667_),
    .B1(_19666_));
 sg13g2_nor2_1 _28182_ (.A(net2330),
    .B(net6513),
    .Y(_19668_));
 sg13g2_a21oi_1 _28183_ (.A1(net6513),
    .A2(_19667_),
    .Y(_00413_),
    .B1(_19668_));
 sg13g2_o21ai_1 _28184_ (.B1(net6941),
    .Y(_19669_),
    .A1(net1766),
    .A2(net7150));
 sg13g2_a21oi_1 _28185_ (.A1(_18305_),
    .A2(net7149),
    .Y(_19670_),
    .B1(_19669_));
 sg13g2_a21oi_1 _28186_ (.A1(\shift_reg[231] ),
    .A2(net6891),
    .Y(_19671_),
    .B1(_19670_));
 sg13g2_nor2_1 _28187_ (.A(net1851),
    .B(net6511),
    .Y(_19672_));
 sg13g2_a21oi_1 _28188_ (.A1(net6511),
    .A2(_19671_),
    .Y(_00414_),
    .B1(_19672_));
 sg13g2_o21ai_1 _28189_ (.B1(net6941),
    .Y(_19673_),
    .A1(net1735),
    .A2(net7149));
 sg13g2_a21oi_1 _28190_ (.A1(_18308_),
    .A2(net7149),
    .Y(_19674_),
    .B1(_19673_));
 sg13g2_a21oi_1 _28191_ (.A1(net2519),
    .A2(net6891),
    .Y(_19675_),
    .B1(_19674_));
 sg13g2_nor2_1 _28192_ (.A(net2525),
    .B(net6512),
    .Y(_19676_));
 sg13g2_a21oi_1 _28193_ (.A1(net6512),
    .A2(_19675_),
    .Y(_00415_),
    .B1(_19676_));
 sg13g2_o21ai_1 _28194_ (.B1(net6942),
    .Y(_19677_),
    .A1(net1415),
    .A2(net7156));
 sg13g2_a21oi_1 _28195_ (.A1(_18307_),
    .A2(net7156),
    .Y(_19678_),
    .B1(_19677_));
 sg13g2_a21oi_1 _28196_ (.A1(net2174),
    .A2(net6891),
    .Y(_19679_),
    .B1(_19678_));
 sg13g2_nor2_1 _28197_ (.A(net2549),
    .B(net6511),
    .Y(_19680_));
 sg13g2_a21oi_1 _28198_ (.A1(net6511),
    .A2(_19679_),
    .Y(_00416_),
    .B1(_19680_));
 sg13g2_o21ai_1 _28199_ (.B1(net6941),
    .Y(_19681_),
    .A1(\perf_triple[0] ),
    .A2(net7149));
 sg13g2_a21oi_1 _28200_ (.A1(_18310_),
    .A2(net7149),
    .Y(_19682_),
    .B1(_19681_));
 sg13g2_a21oi_1 _28201_ (.A1(net2742),
    .A2(net6892),
    .Y(_19683_),
    .B1(_19682_));
 sg13g2_nor2_1 _28202_ (.A(net3062),
    .B(net6514),
    .Y(_19684_));
 sg13g2_a21oi_1 _28203_ (.A1(net6514),
    .A2(_19683_),
    .Y(_00417_),
    .B1(_19684_));
 sg13g2_a21oi_1 _28204_ (.A1(net1664),
    .A2(net7149),
    .Y(_19685_),
    .B1(net6892));
 sg13g2_o21ai_1 _28205_ (.B1(_19685_),
    .Y(_19686_),
    .A1(_18340_),
    .A2(net7149));
 sg13g2_o21ai_1 _28206_ (.B1(_19686_),
    .Y(_19687_),
    .A1(\shift_reg[235] ),
    .A2(net6941));
 sg13g2_nor2_1 _28207_ (.A(net2403),
    .B(net6511),
    .Y(_19688_));
 sg13g2_a21oi_1 _28208_ (.A1(net6511),
    .A2(_19687_),
    .Y(_00418_),
    .B1(_19688_));
 sg13g2_o21ai_1 _28209_ (.B1(net6942),
    .Y(_19689_),
    .A1(net1163),
    .A2(net7150));
 sg13g2_a21oi_1 _28210_ (.A1(_18311_),
    .A2(net7156),
    .Y(_19690_),
    .B1(_19689_));
 sg13g2_a21oi_1 _28211_ (.A1(\shift_reg[236] ),
    .A2(net6891),
    .Y(_19691_),
    .B1(_19690_));
 sg13g2_nor2_1 _28212_ (.A(net2138),
    .B(net6512),
    .Y(_19692_));
 sg13g2_a21oi_1 _28213_ (.A1(net6512),
    .A2(_19691_),
    .Y(_00419_),
    .B1(_19692_));
 sg13g2_a21oi_1 _28214_ (.A1(net1505),
    .A2(net7157),
    .Y(_19693_),
    .B1(net6892));
 sg13g2_o21ai_1 _28215_ (.B1(_19693_),
    .Y(_19694_),
    .A1(_18341_),
    .A2(net7149));
 sg13g2_o21ai_1 _28216_ (.B1(_19694_),
    .Y(_19695_),
    .A1(\shift_reg[237] ),
    .A2(net6941));
 sg13g2_nor2_1 _28217_ (.A(net2608),
    .B(net6511),
    .Y(_19696_));
 sg13g2_a21oi_1 _28218_ (.A1(net6511),
    .A2(_19695_),
    .Y(_00420_),
    .B1(_19696_));
 sg13g2_nand2_1 _28219_ (.Y(_19697_),
    .A(_18312_),
    .B(net7157));
 sg13g2_a21oi_1 _28220_ (.A1(_18342_),
    .A2(_18943_),
    .Y(_19698_),
    .B1(net6891));
 sg13g2_a22oi_1 _28221_ (.Y(_19699_),
    .B1(_19697_),
    .B2(_19698_),
    .A2(net6891),
    .A1(net2330));
 sg13g2_nor2_1 _28222_ (.A(net2391),
    .B(net6512),
    .Y(_19700_));
 sg13g2_a21oi_1 _28223_ (.A1(net6512),
    .A2(_19699_),
    .Y(_00421_),
    .B1(_19700_));
 sg13g2_a21oi_1 _28224_ (.A1(net1422),
    .A2(net7157),
    .Y(_19701_),
    .B1(net6892));
 sg13g2_o21ai_1 _28225_ (.B1(_19701_),
    .Y(_19702_),
    .A1(_18343_),
    .A2(net7151));
 sg13g2_o21ai_1 _28226_ (.B1(_19702_),
    .Y(_19703_),
    .A1(net1851),
    .A2(net6941));
 sg13g2_nor2_1 _28227_ (.A(net2270),
    .B(net6513),
    .Y(_19704_));
 sg13g2_a21oi_1 _28228_ (.A1(net6513),
    .A2(_19703_),
    .Y(_00422_),
    .B1(_19704_));
 sg13g2_o21ai_1 _28229_ (.B1(net6940),
    .Y(_19705_),
    .A1(net2421),
    .A2(net7153));
 sg13g2_a21oi_1 _28230_ (.A1(_18313_),
    .A2(net7153),
    .Y(_19706_),
    .B1(_19705_));
 sg13g2_a21oi_1 _28231_ (.A1(net2525),
    .A2(net6897),
    .Y(_19707_),
    .B1(_19706_));
 sg13g2_nor2_1 _28232_ (.A(net2690),
    .B(net6522),
    .Y(_19708_));
 sg13g2_a21oi_1 _28233_ (.A1(net6512),
    .A2(_19707_),
    .Y(_00423_),
    .B1(_19708_));
 sg13g2_a21oi_1 _28234_ (.A1(net2112),
    .A2(net7151),
    .Y(_19709_),
    .B1(net6897));
 sg13g2_o21ai_1 _28235_ (.B1(_19709_),
    .Y(_19710_),
    .A1(_18344_),
    .A2(net7151));
 sg13g2_o21ai_1 _28236_ (.B1(_19710_),
    .Y(_19711_),
    .A1(net2549),
    .A2(net6940));
 sg13g2_nor2_1 _28237_ (.A(net2636),
    .B(net6523),
    .Y(_19712_));
 sg13g2_a21oi_1 _28238_ (.A1(net6513),
    .A2(_19711_),
    .Y(_00424_),
    .B1(_19712_));
 sg13g2_o21ai_1 _28239_ (.B1(net6940),
    .Y(_19713_),
    .A1(\perf_triple[8] ),
    .A2(net7151));
 sg13g2_a21oi_1 _28240_ (.A1(_18314_),
    .A2(net7151),
    .Y(_19714_),
    .B1(_19713_));
 sg13g2_a21oi_1 _28241_ (.A1(\shift_reg[242] ),
    .A2(net6897),
    .Y(_19715_),
    .B1(_19714_));
 sg13g2_nor2_1 _28242_ (.A(net2564),
    .B(net6522),
    .Y(_19716_));
 sg13g2_a21oi_1 _28243_ (.A1(net6522),
    .A2(_19715_),
    .Y(_00425_),
    .B1(_19716_));
 sg13g2_a21oi_1 _28244_ (.A1(\inv_result[235] ),
    .A2(net7153),
    .Y(_19717_),
    .B1(net6899));
 sg13g2_o21ai_1 _28245_ (.B1(_19717_),
    .Y(_19718_),
    .A1(_18345_),
    .A2(net7151));
 sg13g2_o21ai_1 _28246_ (.B1(_19718_),
    .Y(_19719_),
    .A1(net2403),
    .A2(net6940));
 sg13g2_nor2_1 _28247_ (.A(net3020),
    .B(net6523),
    .Y(_19720_));
 sg13g2_a21oi_1 _28248_ (.A1(net6523),
    .A2(_19719_),
    .Y(_00426_),
    .B1(_19720_));
 sg13g2_o21ai_1 _28249_ (.B1(net6941),
    .Y(_19721_),
    .A1(\perf_double[0] ),
    .A2(net7152));
 sg13g2_a21oi_1 _28250_ (.A1(_18316_),
    .A2(net7151),
    .Y(_19722_),
    .B1(_19721_));
 sg13g2_a21oi_1 _28251_ (.A1(net2138),
    .A2(net6897),
    .Y(_19723_),
    .B1(_19722_));
 sg13g2_nor2_1 _28252_ (.A(net2509),
    .B(net6522),
    .Y(_19724_));
 sg13g2_a21oi_1 _28253_ (.A1(net6522),
    .A2(_19723_),
    .Y(_00427_),
    .B1(_19724_));
 sg13g2_nand2_1 _28254_ (.Y(_19725_),
    .A(_18315_),
    .B(net7151));
 sg13g2_a21oi_1 _28255_ (.A1(_18346_),
    .A2(_18943_),
    .Y(_19726_),
    .B1(net6897));
 sg13g2_a22oi_1 _28256_ (.Y(_19727_),
    .B1(_19725_),
    .B2(_19726_),
    .A2(net6897),
    .A1(net2608));
 sg13g2_nor2_1 _28257_ (.A(net2682),
    .B(net6523),
    .Y(_19728_));
 sg13g2_a21oi_1 _28258_ (.A1(net6526),
    .A2(_19727_),
    .Y(_00428_),
    .B1(_19728_));
 sg13g2_o21ai_1 _28259_ (.B1(net6940),
    .Y(_19729_),
    .A1(net1157),
    .A2(net7152));
 sg13g2_a21oi_1 _28260_ (.A1(_18317_),
    .A2(net7152),
    .Y(_19730_),
    .B1(_19729_));
 sg13g2_a21oi_1 _28261_ (.A1(net2391),
    .A2(net6897),
    .Y(_19731_),
    .B1(_19730_));
 sg13g2_nor2_1 _28262_ (.A(net2618),
    .B(net6522),
    .Y(_19732_));
 sg13g2_a21oi_1 _28263_ (.A1(net6522),
    .A2(_19731_),
    .Y(_00429_),
    .B1(_19732_));
 sg13g2_a21oi_1 _28264_ (.A1(net1681),
    .A2(net7153),
    .Y(_19733_),
    .B1(net6899));
 sg13g2_o21ai_1 _28265_ (.B1(_19733_),
    .Y(_19734_),
    .A1(_18347_),
    .A2(net7152));
 sg13g2_o21ai_1 _28266_ (.B1(_19734_),
    .Y(_19735_),
    .A1(net2270),
    .A2(net6940));
 sg13g2_nor2_1 _28267_ (.A(net2584),
    .B(net6523),
    .Y(_19736_));
 sg13g2_a21oi_1 _28268_ (.A1(net6522),
    .A2(_19735_),
    .Y(_00430_),
    .B1(_19736_));
 sg13g2_o21ai_1 _28269_ (.B1(net6940),
    .Y(_19737_),
    .A1(net1235),
    .A2(net7152));
 sg13g2_a21oi_1 _28270_ (.A1(_18318_),
    .A2(net7152),
    .Y(_19738_),
    .B1(_19737_));
 sg13g2_a21oi_1 _28271_ (.A1(\shift_reg[248] ),
    .A2(net6898),
    .Y(_19739_),
    .B1(_19738_));
 sg13g2_nor2_1 _28272_ (.A(net2649),
    .B(net6524),
    .Y(_19740_));
 sg13g2_a21oi_1 _28273_ (.A1(net6524),
    .A2(_19739_),
    .Y(_00431_),
    .B1(_19740_));
 sg13g2_a21oi_1 _28274_ (.A1(net1904),
    .A2(net7158),
    .Y(_19741_),
    .B1(net6897));
 sg13g2_o21ai_1 _28275_ (.B1(_19741_),
    .Y(_19742_),
    .A1(_18348_),
    .A2(net7158));
 sg13g2_o21ai_1 _28276_ (.B1(_19742_),
    .Y(_19743_),
    .A1(\shift_reg[249] ),
    .A2(net6940));
 sg13g2_nor2_1 _28277_ (.A(net2208),
    .B(net6524),
    .Y(_19744_));
 sg13g2_a21oi_1 _28278_ (.A1(net6523),
    .A2(_19743_),
    .Y(_00432_),
    .B1(_19744_));
 sg13g2_o21ai_1 _28279_ (.B1(net6944),
    .Y(_19745_),
    .A1(net1255),
    .A2(net7158));
 sg13g2_a21oi_1 _28280_ (.A1(_18320_),
    .A2(net7158),
    .Y(_19746_),
    .B1(_19745_));
 sg13g2_a21oi_1 _28281_ (.A1(\shift_reg[250] ),
    .A2(net6898),
    .Y(_19747_),
    .B1(_19746_));
 sg13g2_nor2_1 _28282_ (.A(net2156),
    .B(net6524),
    .Y(_19748_));
 sg13g2_a21oi_1 _28283_ (.A1(net6524),
    .A2(_19747_),
    .Y(_00433_),
    .B1(_19748_));
 sg13g2_a21oi_1 _28284_ (.A1(net1278),
    .A2(net7159),
    .Y(_19749_),
    .B1(net6898));
 sg13g2_o21ai_1 _28285_ (.B1(_19749_),
    .Y(_19750_),
    .A1(_18349_),
    .A2(net7158));
 sg13g2_o21ai_1 _28286_ (.B1(_19750_),
    .Y(_19751_),
    .A1(\shift_reg[251] ),
    .A2(net6944));
 sg13g2_nor2_1 _28287_ (.A(net2158),
    .B(net6525),
    .Y(_19752_));
 sg13g2_a21oi_1 _28288_ (.A1(net6525),
    .A2(_19751_),
    .Y(_00434_),
    .B1(_19752_));
 sg13g2_o21ai_1 _28289_ (.B1(net6944),
    .Y(_19753_),
    .A1(net1286),
    .A2(net7159));
 sg13g2_a21oi_1 _28290_ (.A1(_18322_),
    .A2(net7159),
    .Y(_19754_),
    .B1(_19753_));
 sg13g2_a21oi_1 _28291_ (.A1(net2509),
    .A2(net6898),
    .Y(_19755_),
    .B1(_19754_));
 sg13g2_nor2_1 _28292_ (.A(net2799),
    .B(net6524),
    .Y(_19756_));
 sg13g2_a21oi_1 _28293_ (.A1(net6524),
    .A2(_19755_),
    .Y(_00435_),
    .B1(_19756_));
 sg13g2_nand2_1 _28294_ (.Y(_19757_),
    .A(_18321_),
    .B(net7160));
 sg13g2_a21oi_1 _28295_ (.A1(_18350_),
    .A2(_18943_),
    .Y(_19758_),
    .B1(net6899));
 sg13g2_a22oi_1 _28296_ (.Y(_19759_),
    .B1(_19757_),
    .B2(_19758_),
    .A2(net6899),
    .A1(net2682));
 sg13g2_nor2_1 _28297_ (.A(net2982),
    .B(net6526),
    .Y(_19760_));
 sg13g2_a21oi_1 _28298_ (.A1(net6526),
    .A2(_19759_),
    .Y(_00436_),
    .B1(_19760_));
 sg13g2_o21ai_1 _28299_ (.B1(net6944),
    .Y(_19761_),
    .A1(net1187),
    .A2(net7158));
 sg13g2_a21oi_1 _28300_ (.A1(_18324_),
    .A2(net7158),
    .Y(_19762_),
    .B1(_19761_));
 sg13g2_a21oi_1 _28301_ (.A1(\shift_reg[254] ),
    .A2(net6898),
    .Y(_19763_),
    .B1(_19762_));
 sg13g2_nor2_1 _28302_ (.A(net2109),
    .B(net6525),
    .Y(_19764_));
 sg13g2_a21oi_1 _28303_ (.A1(net6524),
    .A2(_19763_),
    .Y(_00437_),
    .B1(_19764_));
 sg13g2_o21ai_1 _28304_ (.B1(net6944),
    .Y(_19765_),
    .A1(\perf_total[1] ),
    .A2(net7159));
 sg13g2_a21oi_1 _28305_ (.A1(_18323_),
    .A2(net7158),
    .Y(_19766_),
    .B1(_19765_));
 sg13g2_a21oi_1 _28306_ (.A1(\shift_reg[255] ),
    .A2(net6898),
    .Y(_19767_),
    .B1(_19766_));
 sg13g2_nor2_1 _28307_ (.A(net2287),
    .B(net6525),
    .Y(_19768_));
 sg13g2_a21oi_1 _28308_ (.A1(net6525),
    .A2(_19767_),
    .Y(_00438_),
    .B1(_19768_));
 sg13g2_nand2_1 _28309_ (.Y(_19769_),
    .A(_18326_),
    .B(net7159));
 sg13g2_a21oi_1 _28310_ (.A1(_18351_),
    .A2(_18943_),
    .Y(_19770_),
    .B1(net6900));
 sg13g2_a22oi_1 _28311_ (.Y(_19771_),
    .B1(_19769_),
    .B2(_19770_),
    .A2(net6901),
    .A1(\shift_reg[256] ));
 sg13g2_nor2_1 _28312_ (.A(net2626),
    .B(net6527),
    .Y(_19772_));
 sg13g2_a21oi_1 _28313_ (.A1(net6527),
    .A2(_19771_),
    .Y(_00439_),
    .B1(_19772_));
 sg13g2_o21ai_1 _28314_ (.B1(net6944),
    .Y(_19773_),
    .A1(net1161),
    .A2(net7160));
 sg13g2_a21oi_1 _28315_ (.A1(_18325_),
    .A2(net7159),
    .Y(_19774_),
    .B1(_19773_));
 sg13g2_a21oi_1 _28316_ (.A1(net2208),
    .A2(net6900),
    .Y(_19775_),
    .B1(_19774_));
 sg13g2_nor2_1 _28317_ (.A(net2619),
    .B(net6528),
    .Y(_19776_));
 sg13g2_a21oi_1 _28318_ (.A1(net6528),
    .A2(_19775_),
    .Y(_00440_),
    .B1(_19776_));
 sg13g2_o21ai_1 _28319_ (.B1(net6945),
    .Y(_19777_),
    .A1(net1193),
    .A2(net7160));
 sg13g2_a21oi_1 _28320_ (.A1(_18328_),
    .A2(net7160),
    .Y(_19778_),
    .B1(_19777_));
 sg13g2_a21oi_1 _28321_ (.A1(net2156),
    .A2(net6900),
    .Y(_19779_),
    .B1(_19778_));
 sg13g2_nor2_1 _28322_ (.A(net2479),
    .B(net6528),
    .Y(_19780_));
 sg13g2_a21oi_1 _28323_ (.A1(net6528),
    .A2(_19779_),
    .Y(_00441_),
    .B1(_19780_));
 sg13g2_nand2_1 _28324_ (.Y(_19781_),
    .A(_18327_),
    .B(net7159));
 sg13g2_a21oi_1 _28325_ (.A1(_18352_),
    .A2(_18943_),
    .Y(_19782_),
    .B1(net6900));
 sg13g2_a22oi_1 _28326_ (.Y(_19783_),
    .B1(_19781_),
    .B2(_19782_),
    .A2(net6900),
    .A1(net2158));
 sg13g2_nor2_1 _28327_ (.A(net2860),
    .B(net6528),
    .Y(_19784_));
 sg13g2_a21oi_1 _28328_ (.A1(net6527),
    .A2(_19783_),
    .Y(_00442_),
    .B1(_19784_));
 sg13g2_o21ai_1 _28329_ (.B1(net6944),
    .Y(_19785_),
    .A1(net1183),
    .A2(net7161));
 sg13g2_a21oi_1 _28330_ (.A1(_18330_),
    .A2(net7160),
    .Y(_19786_),
    .B1(_19785_));
 sg13g2_a21oi_1 _28331_ (.A1(\shift_reg[260] ),
    .A2(net6900),
    .Y(_19787_),
    .B1(_19786_));
 sg13g2_nor2_1 _28332_ (.A(net2574),
    .B(net6527),
    .Y(_19788_));
 sg13g2_a21oi_1 _28333_ (.A1(net6527),
    .A2(_19787_),
    .Y(_00443_),
    .B1(_19788_));
 sg13g2_nand2_1 _28334_ (.Y(_19789_),
    .A(_18329_),
    .B(net7160));
 sg13g2_a21oi_1 _28335_ (.A1(_18353_),
    .A2(_18943_),
    .Y(_19790_),
    .B1(net6902));
 sg13g2_a22oi_1 _28336_ (.Y(_19791_),
    .B1(_19789_),
    .B2(_19790_),
    .A2(net6902),
    .A1(\shift_reg[261] ));
 sg13g2_nor2_1 _28337_ (.A(net2928),
    .B(net6531),
    .Y(_19792_));
 sg13g2_a21oi_1 _28338_ (.A1(net6531),
    .A2(_19791_),
    .Y(_00444_),
    .B1(_19792_));
 sg13g2_o21ai_1 _28339_ (.B1(net6944),
    .Y(_19793_),
    .A1(net2069),
    .A2(net7161));
 sg13g2_a21oi_1 _28340_ (.A1(_18332_),
    .A2(net7160),
    .Y(_19794_),
    .B1(_19793_));
 sg13g2_a21oi_1 _28341_ (.A1(net2109),
    .A2(net6900),
    .Y(_19795_),
    .B1(_19794_));
 sg13g2_nor2_1 _28342_ (.A(net2570),
    .B(net6527),
    .Y(_19796_));
 sg13g2_a21oi_1 _28343_ (.A1(net6528),
    .A2(_19795_),
    .Y(_00445_),
    .B1(_19796_));
 sg13g2_o21ai_1 _28344_ (.B1(net6945),
    .Y(_19797_),
    .A1(\perf_total[9] ),
    .A2(net7161));
 sg13g2_a21oi_1 _28345_ (.A1(_18331_),
    .A2(net7161),
    .Y(_19798_),
    .B1(_19797_));
 sg13g2_a21oi_1 _28346_ (.A1(net2287),
    .A2(net6900),
    .Y(_19799_),
    .B1(_19798_));
 sg13g2_nor2_1 _28347_ (.A(net2430),
    .B(net6527),
    .Y(_19800_));
 sg13g2_a21oi_1 _28348_ (.A1(net6527),
    .A2(_19799_),
    .Y(_00446_),
    .B1(_19800_));
 sg13g2_nor2b_1 _28349_ (.A(_18617_),
    .B_N(_18909_),
    .Y(_19801_));
 sg13g2_a21oi_1 _28350_ (.A1(_18624_),
    .A2(_19801_),
    .Y(_19802_),
    .B1(net1179));
 sg13g2_a21oi_1 _28351_ (.A1(_18617_),
    .A2(_18909_),
    .Y(_19803_),
    .B1(net6901));
 sg13g2_nor2_1 _28352_ (.A(net1180),
    .B(_19803_),
    .Y(_00447_));
 sg13g2_a22oi_1 _28353_ (.Y(_19804_),
    .B1(_19801_),
    .B2(_18898_),
    .A2(_18900_),
    .A1(net1678));
 sg13g2_inv_1 _28354_ (.Y(_00448_),
    .A(net1679));
 sg13g2_mux2_1 _28355_ (.A0(\u_trng.entropy_bit ),
    .A1(net2851),
    .S(net2257),
    .X(_00449_));
 sg13g2_mux2_1 _28356_ (.A0(\trng_data[0] ),
    .A1(net2279),
    .S(net6677),
    .X(_00450_));
 sg13g2_mux2_1 _28357_ (.A0(\trng_data[1] ),
    .A1(net2264),
    .S(net6677),
    .X(_00451_));
 sg13g2_mux2_1 _28358_ (.A0(\trng_data[2] ),
    .A1(net2062),
    .S(net6677),
    .X(_00452_));
 sg13g2_mux2_1 _28359_ (.A0(net2062),
    .A1(net1962),
    .S(net6677),
    .X(_00453_));
 sg13g2_mux2_1 _28360_ (.A0(net1962),
    .A1(net1917),
    .S(net6677),
    .X(_00454_));
 sg13g2_mux2_1 _28361_ (.A0(net1917),
    .A1(\trng_data[6] ),
    .S(net6677),
    .X(_00455_));
 sg13g2_mux2_1 _28362_ (.A0(\trng_data[6] ),
    .A1(net1361),
    .S(_18632_),
    .X(_00456_));
 sg13g2_nor2_1 _28363_ (.A(net1176),
    .B(trng_ready),
    .Y(_19805_));
 sg13g2_xnor2_1 _28364_ (.Y(_00457_),
    .A(net1176),
    .B(trng_ready));
 sg13g2_mux2_1 _28365_ (.A0(net2542),
    .A1(\u_trng.entropy_bit ),
    .S(_19805_),
    .X(_00458_));
 sg13g2_a21oi_1 _28366_ (.A1(_18181_),
    .A2(_18182_),
    .Y(_00459_),
    .B1(net1147));
 sg13g2_nor2b_2 _28367_ (.A(\u_inv.state[1] ),
    .B_N(\u_inv.state[0] ),
    .Y(_19806_));
 sg13g2_nand2b_2 _28368_ (.Y(_19807_),
    .B(\u_inv.state[0] ),
    .A_N(\u_inv.state[1] ));
 sg13g2_nor2_2 _28369_ (.A(_24689_[0]),
    .B(net7081),
    .Y(_19808_));
 sg13g2_nand2_2 _28370_ (.Y(_19809_),
    .A(net6606),
    .B(net7016));
 sg13g2_and2_1 _28371_ (.A(net7444),
    .B(_19809_),
    .X(_19810_));
 sg13g2_nand2_2 _28372_ (.Y(_19811_),
    .A(net7444),
    .B(_19809_));
 sg13g2_nor2_1 _28373_ (.A(net7225),
    .B(\u_inv.delta_reg[9] ),
    .Y(_19812_));
 sg13g2_nand2b_2 _28374_ (.Y(_19813_),
    .B(net7376),
    .A_N(\u_inv.delta_reg[9] ));
 sg13g2_nor2_1 _28375_ (.A(\u_inv.delta_reg[1] ),
    .B(\u_inv.delta_reg[2] ),
    .Y(_19814_));
 sg13g2_nand2_1 _28376_ (.Y(_19815_),
    .A(_18185_),
    .B(_19814_));
 sg13g2_nor3_1 _28377_ (.A(\u_inv.delta_reg[5] ),
    .B(\u_inv.delta_reg[4] ),
    .C(_19815_),
    .Y(_19816_));
 sg13g2_nand2_1 _28378_ (.Y(_19817_),
    .A(_18186_),
    .B(_19816_));
 sg13g2_nor2_1 _28379_ (.A(\u_inv.delta_reg[7] ),
    .B(_19817_),
    .Y(_19818_));
 sg13g2_a21oi_2 _28380_ (.B1(_19813_),
    .Y(_19819_),
    .A2(_19818_),
    .A1(_18187_));
 sg13g2_a21o_1 _28381_ (.A2(_19812_),
    .A1(\u_inv.delta_double[0] ),
    .B1(_19819_),
    .X(_19820_));
 sg13g2_a21oi_1 _28382_ (.A1(\u_inv.delta_double[0] ),
    .A2(_19812_),
    .Y(_19821_),
    .B1(_19819_));
 sg13g2_nand2_1 _28383_ (.Y(_19822_),
    .A(\u_inv.f_next[2] ),
    .B(\u_inv.f_reg[2] ));
 sg13g2_inv_1 _28384_ (.Y(_19823_),
    .A(_19822_));
 sg13g2_or2_1 _28385_ (.X(_19824_),
    .B(\u_inv.f_reg[2] ),
    .A(\u_inv.f_next[2] ));
 sg13g2_and2_1 _28386_ (.A(_19822_),
    .B(_19824_),
    .X(_19825_));
 sg13g2_nor2b_1 _28387_ (.A(\u_inv.f_next[1] ),
    .B_N(\u_inv.f_reg[1] ),
    .Y(_19826_));
 sg13g2_nand2b_1 _28388_ (.Y(_19827_),
    .B(\u_inv.f_next[1] ),
    .A_N(\u_inv.f_reg[1] ));
 sg13g2_nor2b_1 _28389_ (.A(net7315),
    .B_N(\u_inv.f_reg[0] ),
    .Y(_19828_));
 sg13g2_a21oi_1 _28390_ (.A1(_19827_),
    .A2(_19828_),
    .Y(_19829_),
    .B1(_19826_));
 sg13g2_a221oi_1 _28391_ (.B2(_19828_),
    .C1(_19826_),
    .B1(_19827_),
    .A1(_19822_),
    .Y(_19830_),
    .A2(_19824_));
 sg13g2_nor2b_1 _28392_ (.A(_19829_),
    .B_N(_19825_),
    .Y(_19831_));
 sg13g2_nor3_1 _28393_ (.A(net6205),
    .B(_19830_),
    .C(_19831_),
    .Y(_19832_));
 sg13g2_nor2_1 _28394_ (.A(\u_inv.f_next[2] ),
    .B(net7314),
    .Y(_19833_));
 sg13g2_xnor2_1 _28395_ (.Y(_19834_),
    .A(\u_inv.f_next[1] ),
    .B(\u_inv.f_reg[1] ));
 sg13g2_nand2_1 _28396_ (.Y(_19835_),
    .A(net7315),
    .B(\u_inv.f_reg[0] ));
 sg13g2_nand2_1 _28397_ (.Y(_19836_),
    .A(\u_inv.f_next[1] ),
    .B(\u_inv.f_reg[1] ));
 sg13g2_o21ai_1 _28398_ (.B1(_19836_),
    .Y(_19837_),
    .A1(_19834_),
    .A2(_19835_));
 sg13g2_xnor2_1 _28399_ (.Y(_19838_),
    .A(_19825_),
    .B(_19837_));
 sg13g2_a21oi_1 _28400_ (.A1(net7315),
    .A2(_19838_),
    .Y(_19839_),
    .B1(_19833_));
 sg13g2_nand2_1 _28401_ (.Y(_19840_),
    .A(net6205),
    .B(_19839_));
 sg13g2_nor2b_2 _28402_ (.A(_19832_),
    .B_N(_19840_),
    .Y(_19841_));
 sg13g2_nand2b_2 _28403_ (.Y(_19842_),
    .B(_19840_),
    .A_N(_19832_));
 sg13g2_xor2_1 _28404_ (.B(\u_inv.f_reg[255] ),
    .A(\u_inv.f_next[255] ),
    .X(_19843_));
 sg13g2_xnor2_1 _28405_ (.Y(_19844_),
    .A(\u_inv.f_next[255] ),
    .B(\u_inv.f_reg[255] ));
 sg13g2_and2_1 _28406_ (.A(\u_inv.f_next[254] ),
    .B(\u_inv.f_reg[254] ),
    .X(_19845_));
 sg13g2_xor2_1 _28407_ (.B(\u_inv.f_reg[254] ),
    .A(\u_inv.f_next[254] ),
    .X(_19846_));
 sg13g2_xnor2_1 _28408_ (.Y(_19847_),
    .A(\u_inv.f_next[254] ),
    .B(\u_inv.f_reg[254] ));
 sg13g2_nand2_1 _28409_ (.Y(_19848_),
    .A(\u_inv.f_next[253] ),
    .B(\u_inv.f_reg[253] ));
 sg13g2_nand2_1 _28410_ (.Y(_19849_),
    .A(\u_inv.f_next[252] ),
    .B(\u_inv.f_reg[252] ));
 sg13g2_nand2_1 _28411_ (.Y(_19850_),
    .A(_19848_),
    .B(_19849_));
 sg13g2_o21ai_1 _28412_ (.B1(_19850_),
    .Y(_19851_),
    .A1(\u_inv.f_next[253] ),
    .A2(\u_inv.f_reg[253] ));
 sg13g2_xor2_1 _28413_ (.B(\u_inv.f_reg[253] ),
    .A(\u_inv.f_next[253] ),
    .X(_19852_));
 sg13g2_xnor2_1 _28414_ (.Y(_19853_),
    .A(\u_inv.f_next[253] ),
    .B(\u_inv.f_reg[253] ));
 sg13g2_xor2_1 _28415_ (.B(\u_inv.f_reg[252] ),
    .A(\u_inv.f_next[252] ),
    .X(_19854_));
 sg13g2_xnor2_1 _28416_ (.Y(_19855_),
    .A(\u_inv.f_next[252] ),
    .B(\u_inv.f_reg[252] ));
 sg13g2_nor2_1 _28417_ (.A(_19853_),
    .B(_19855_),
    .Y(_19856_));
 sg13g2_xor2_1 _28418_ (.B(\u_inv.f_reg[251] ),
    .A(\u_inv.f_next[251] ),
    .X(_19857_));
 sg13g2_inv_1 _28419_ (.Y(_19858_),
    .A(_19857_));
 sg13g2_nand2_1 _28420_ (.Y(_19859_),
    .A(\u_inv.f_next[250] ),
    .B(\u_inv.f_reg[250] ));
 sg13g2_xnor2_1 _28421_ (.Y(_19860_),
    .A(\u_inv.f_next[250] ),
    .B(\u_inv.f_reg[250] ));
 sg13g2_nor2_1 _28422_ (.A(_19858_),
    .B(_19860_),
    .Y(_19861_));
 sg13g2_and2_1 _28423_ (.A(\u_inv.f_next[248] ),
    .B(\u_inv.f_reg[248] ),
    .X(_19862_));
 sg13g2_a21oi_1 _28424_ (.A1(\u_inv.f_next[249] ),
    .A2(\u_inv.f_reg[249] ),
    .Y(_19863_),
    .B1(_19862_));
 sg13g2_inv_1 _28425_ (.Y(_19864_),
    .A(_19863_));
 sg13g2_o21ai_1 _28426_ (.B1(_19864_),
    .Y(_19865_),
    .A1(\u_inv.f_next[249] ),
    .A2(\u_inv.f_reg[249] ));
 sg13g2_inv_1 _28427_ (.Y(_19866_),
    .A(_19865_));
 sg13g2_a21oi_1 _28428_ (.A1(_17963_),
    .A2(_18253_),
    .Y(_19867_),
    .B1(_19859_));
 sg13g2_a221oi_1 _28429_ (.B2(_19866_),
    .C1(_19867_),
    .B1(_19861_),
    .A1(\u_inv.f_next[251] ),
    .Y(_19868_),
    .A2(\u_inv.f_reg[251] ));
 sg13g2_inv_1 _28430_ (.Y(_19869_),
    .A(_19868_));
 sg13g2_nor2_1 _28431_ (.A(\u_inv.f_next[223] ),
    .B(\u_inv.f_reg[223] ),
    .Y(_19870_));
 sg13g2_xor2_1 _28432_ (.B(\u_inv.f_reg[223] ),
    .A(\u_inv.f_next[223] ),
    .X(_19871_));
 sg13g2_nand2_1 _28433_ (.Y(_19872_),
    .A(\u_inv.f_next[222] ),
    .B(\u_inv.f_reg[222] ));
 sg13g2_xor2_1 _28434_ (.B(\u_inv.f_reg[222] ),
    .A(\u_inv.f_next[222] ),
    .X(_19873_));
 sg13g2_xnor2_1 _28435_ (.Y(_19874_),
    .A(\u_inv.f_next[222] ),
    .B(\u_inv.f_reg[222] ));
 sg13g2_nand2_1 _28436_ (.Y(_19875_),
    .A(_19871_),
    .B(_19873_));
 sg13g2_nor2_1 _28437_ (.A(\u_inv.f_next[221] ),
    .B(\u_inv.f_reg[221] ),
    .Y(_19876_));
 sg13g2_xnor2_1 _28438_ (.Y(_19877_),
    .A(\u_inv.f_next[221] ),
    .B(\u_inv.f_reg[221] ));
 sg13g2_and2_1 _28439_ (.A(\u_inv.f_next[220] ),
    .B(\u_inv.f_reg[220] ),
    .X(_19878_));
 sg13g2_xor2_1 _28440_ (.B(\u_inv.f_reg[220] ),
    .A(\u_inv.f_next[220] ),
    .X(_19879_));
 sg13g2_xnor2_1 _28441_ (.Y(_19880_),
    .A(\u_inv.f_next[220] ),
    .B(\u_inv.f_reg[220] ));
 sg13g2_nand2b_1 _28442_ (.Y(_19881_),
    .B(_19879_),
    .A_N(_19877_));
 sg13g2_or2_1 _28443_ (.X(_19882_),
    .B(_19881_),
    .A(_19875_));
 sg13g2_nand2_1 _28444_ (.Y(_19883_),
    .A(\u_inv.f_next[218] ),
    .B(\u_inv.f_reg[218] ));
 sg13g2_xor2_1 _28445_ (.B(\u_inv.f_reg[218] ),
    .A(\u_inv.f_next[218] ),
    .X(_19884_));
 sg13g2_xnor2_1 _28446_ (.Y(_19885_),
    .A(\u_inv.f_next[218] ),
    .B(\u_inv.f_reg[218] ));
 sg13g2_nand2_1 _28447_ (.Y(_19886_),
    .A(\u_inv.f_next[219] ),
    .B(\u_inv.f_reg[219] ));
 sg13g2_xor2_1 _28448_ (.B(\u_inv.f_reg[219] ),
    .A(\u_inv.f_next[219] ),
    .X(_19887_));
 sg13g2_nand2_1 _28449_ (.Y(_19888_),
    .A(_19884_),
    .B(_19887_));
 sg13g2_and2_1 _28450_ (.A(\u_inv.f_next[216] ),
    .B(\u_inv.f_reg[216] ),
    .X(_19889_));
 sg13g2_a21o_1 _28451_ (.A2(\u_inv.f_reg[217] ),
    .A1(\u_inv.f_next[217] ),
    .B1(_19889_),
    .X(_19890_));
 sg13g2_o21ai_1 _28452_ (.B1(_19890_),
    .Y(_19891_),
    .A1(\u_inv.f_next[217] ),
    .A2(\u_inv.f_reg[217] ));
 sg13g2_a21oi_1 _28453_ (.A1(_17979_),
    .A2(_18249_),
    .Y(_19892_),
    .B1(_19883_));
 sg13g2_o21ai_1 _28454_ (.B1(_19886_),
    .Y(_19893_),
    .A1(_19888_),
    .A2(_19891_));
 sg13g2_nor2_2 _28455_ (.A(_19892_),
    .B(_19893_),
    .Y(_19894_));
 sg13g2_a21oi_1 _28456_ (.A1(\u_inv.f_next[221] ),
    .A2(\u_inv.f_reg[221] ),
    .Y(_19895_),
    .B1(_19878_));
 sg13g2_nor2_1 _28457_ (.A(_19876_),
    .B(_19895_),
    .Y(_19896_));
 sg13g2_nand2b_1 _28458_ (.Y(_19897_),
    .B(_19896_),
    .A_N(_19875_));
 sg13g2_o21ai_1 _28459_ (.B1(_19897_),
    .Y(_19898_),
    .A1(_19870_),
    .A2(_19872_));
 sg13g2_a21oi_1 _28460_ (.A1(\u_inv.f_next[223] ),
    .A2(\u_inv.f_reg[223] ),
    .Y(_19899_),
    .B1(_19898_));
 sg13g2_o21ai_1 _28461_ (.B1(_19899_),
    .Y(_19900_),
    .A1(_19882_),
    .A2(_19894_));
 sg13g2_xor2_1 _28462_ (.B(\u_inv.f_reg[217] ),
    .A(\u_inv.f_next[217] ),
    .X(_19901_));
 sg13g2_xnor2_1 _28463_ (.Y(_19902_),
    .A(\u_inv.f_next[217] ),
    .B(\u_inv.f_reg[217] ));
 sg13g2_xnor2_1 _28464_ (.Y(_19903_),
    .A(\u_inv.f_next[216] ),
    .B(\u_inv.f_reg[216] ));
 sg13g2_nor2_1 _28465_ (.A(_19902_),
    .B(_19903_),
    .Y(_19904_));
 sg13g2_inv_1 _28466_ (.Y(_19905_),
    .A(_19904_));
 sg13g2_nand2b_1 _28467_ (.Y(_19906_),
    .B(_19904_),
    .A_N(_19888_));
 sg13g2_nor2_1 _28468_ (.A(_19882_),
    .B(_19906_),
    .Y(_19907_));
 sg13g2_and2_1 _28469_ (.A(\u_inv.f_next[214] ),
    .B(\u_inv.f_reg[214] ),
    .X(_19908_));
 sg13g2_xor2_1 _28470_ (.B(\u_inv.f_reg[214] ),
    .A(\u_inv.f_next[214] ),
    .X(_19909_));
 sg13g2_xnor2_1 _28471_ (.Y(_19910_),
    .A(\u_inv.f_next[214] ),
    .B(\u_inv.f_reg[214] ));
 sg13g2_nand2_1 _28472_ (.Y(_19911_),
    .A(\u_inv.f_next[215] ),
    .B(\u_inv.f_reg[215] ));
 sg13g2_xnor2_1 _28473_ (.Y(_19912_),
    .A(\u_inv.f_next[215] ),
    .B(\u_inv.f_reg[215] ));
 sg13g2_xor2_1 _28474_ (.B(\u_inv.f_reg[213] ),
    .A(\u_inv.f_next[213] ),
    .X(_19913_));
 sg13g2_xnor2_1 _28475_ (.Y(_19914_),
    .A(\u_inv.f_next[213] ),
    .B(\u_inv.f_reg[213] ));
 sg13g2_nand2_1 _28476_ (.Y(_19915_),
    .A(\u_inv.f_next[212] ),
    .B(\u_inv.f_reg[212] ));
 sg13g2_xor2_1 _28477_ (.B(\u_inv.f_reg[212] ),
    .A(\u_inv.f_next[212] ),
    .X(_19916_));
 sg13g2_xnor2_1 _28478_ (.Y(_19917_),
    .A(\u_inv.f_next[212] ),
    .B(\u_inv.f_reg[212] ));
 sg13g2_nor2_1 _28479_ (.A(_19914_),
    .B(_19917_),
    .Y(_19918_));
 sg13g2_nor4_1 _28480_ (.A(_19910_),
    .B(_19912_),
    .C(_19914_),
    .D(_19917_),
    .Y(_19919_));
 sg13g2_nand2_1 _28481_ (.Y(_19920_),
    .A(\u_inv.f_next[210] ),
    .B(\u_inv.f_reg[210] ));
 sg13g2_xor2_1 _28482_ (.B(\u_inv.f_reg[210] ),
    .A(\u_inv.f_next[210] ),
    .X(_19921_));
 sg13g2_xnor2_1 _28483_ (.Y(_19922_),
    .A(\u_inv.f_next[210] ),
    .B(\u_inv.f_reg[210] ));
 sg13g2_nor2_1 _28484_ (.A(\u_inv.f_next[211] ),
    .B(\u_inv.f_reg[211] ),
    .Y(_19923_));
 sg13g2_xnor2_1 _28485_ (.Y(_19924_),
    .A(\u_inv.f_next[211] ),
    .B(\u_inv.f_reg[211] ));
 sg13g2_nor2_1 _28486_ (.A(_19922_),
    .B(_19924_),
    .Y(_19925_));
 sg13g2_nor2_1 _28487_ (.A(\u_inv.f_next[209] ),
    .B(\u_inv.f_reg[209] ),
    .Y(_19926_));
 sg13g2_a22oi_1 _28488_ (.Y(_19927_),
    .B1(\u_inv.f_reg[209] ),
    .B2(\u_inv.f_next[209] ),
    .A2(\u_inv.f_reg[208] ),
    .A1(\u_inv.f_next[208] ));
 sg13g2_nor2_1 _28489_ (.A(_19926_),
    .B(_19927_),
    .Y(_19928_));
 sg13g2_a22oi_1 _28490_ (.Y(_19929_),
    .B1(_19925_),
    .B2(_19928_),
    .A2(\u_inv.f_reg[211] ),
    .A1(\u_inv.f_next[211] ));
 sg13g2_o21ai_1 _28491_ (.B1(_19929_),
    .Y(_19930_),
    .A1(_19920_),
    .A2(_19923_));
 sg13g2_o21ai_1 _28492_ (.B1(_19908_),
    .Y(_19931_),
    .A1(\u_inv.f_next[215] ),
    .A2(\u_inv.f_reg[215] ));
 sg13g2_a22oi_1 _28493_ (.Y(_19932_),
    .B1(\u_inv.f_reg[213] ),
    .B2(\u_inv.f_next[213] ),
    .A2(\u_inv.f_reg[212] ),
    .A1(\u_inv.f_next[212] ));
 sg13g2_a21o_1 _28494_ (.A2(_18248_),
    .A1(_17983_),
    .B1(_19932_),
    .X(_19933_));
 sg13g2_nor3_1 _28495_ (.A(_19910_),
    .B(_19912_),
    .C(_19933_),
    .Y(_19934_));
 sg13g2_a21oi_1 _28496_ (.A1(_19919_),
    .A2(_19930_),
    .Y(_19935_),
    .B1(_19934_));
 sg13g2_nand3_1 _28497_ (.B(_19931_),
    .C(_19935_),
    .A(_19911_),
    .Y(_19936_));
 sg13g2_inv_2 _28498_ (.Y(_19937_),
    .A(_19936_));
 sg13g2_xnor2_1 _28499_ (.Y(_19938_),
    .A(\u_inv.f_next[209] ),
    .B(\u_inv.f_reg[209] ));
 sg13g2_xor2_1 _28500_ (.B(\u_inv.f_reg[208] ),
    .A(\u_inv.f_next[208] ),
    .X(_19939_));
 sg13g2_xnor2_1 _28501_ (.Y(_19940_),
    .A(\u_inv.f_next[208] ),
    .B(\u_inv.f_reg[208] ));
 sg13g2_nor2_1 _28502_ (.A(_19938_),
    .B(_19940_),
    .Y(_19941_));
 sg13g2_and2_1 _28503_ (.A(_19925_),
    .B(_19941_),
    .X(_19942_));
 sg13g2_inv_1 _28504_ (.Y(_19943_),
    .A(_19942_));
 sg13g2_and2_1 _28505_ (.A(_19919_),
    .B(_19942_),
    .X(_19944_));
 sg13g2_inv_1 _28506_ (.Y(_19945_),
    .A(_19944_));
 sg13g2_and2_1 _28507_ (.A(_19907_),
    .B(_19944_),
    .X(_19946_));
 sg13g2_nand2_1 _28508_ (.Y(_19947_),
    .A(\u_inv.f_next[207] ),
    .B(\u_inv.f_reg[207] ));
 sg13g2_xnor2_1 _28509_ (.Y(_19948_),
    .A(\u_inv.f_next[207] ),
    .B(\u_inv.f_reg[207] ));
 sg13g2_and2_1 _28510_ (.A(\u_inv.f_next[206] ),
    .B(\u_inv.f_reg[206] ),
    .X(_19949_));
 sg13g2_xor2_1 _28511_ (.B(\u_inv.f_reg[206] ),
    .A(\u_inv.f_next[206] ),
    .X(_19950_));
 sg13g2_xnor2_1 _28512_ (.Y(_19951_),
    .A(\u_inv.f_next[206] ),
    .B(\u_inv.f_reg[206] ));
 sg13g2_nor2_1 _28513_ (.A(_19948_),
    .B(_19951_),
    .Y(_19952_));
 sg13g2_nand2_1 _28514_ (.Y(_19953_),
    .A(\u_inv.f_next[204] ),
    .B(\u_inv.f_reg[204] ));
 sg13g2_xor2_1 _28515_ (.B(\u_inv.f_reg[204] ),
    .A(\u_inv.f_next[204] ),
    .X(_19954_));
 sg13g2_xnor2_1 _28516_ (.Y(_19955_),
    .A(\u_inv.f_next[204] ),
    .B(\u_inv.f_reg[204] ));
 sg13g2_xor2_1 _28517_ (.B(\u_inv.f_reg[205] ),
    .A(\u_inv.f_next[205] ),
    .X(_19956_));
 sg13g2_and2_1 _28518_ (.A(_19954_),
    .B(_19956_),
    .X(_19957_));
 sg13g2_and2_1 _28519_ (.A(_19952_),
    .B(_19957_),
    .X(_19958_));
 sg13g2_nand2_1 _28520_ (.Y(_19959_),
    .A(_19952_),
    .B(_19957_));
 sg13g2_nand2_1 _28521_ (.Y(_19960_),
    .A(\u_inv.f_next[202] ),
    .B(\u_inv.f_reg[202] ));
 sg13g2_xnor2_1 _28522_ (.Y(_19961_),
    .A(\u_inv.f_next[202] ),
    .B(\u_inv.f_reg[202] ));
 sg13g2_inv_1 _28523_ (.Y(_19962_),
    .A(_19961_));
 sg13g2_nor2_1 _28524_ (.A(\u_inv.f_next[203] ),
    .B(\u_inv.f_reg[203] ),
    .Y(_19963_));
 sg13g2_xor2_1 _28525_ (.B(\u_inv.f_reg[203] ),
    .A(\u_inv.f_next[203] ),
    .X(_19964_));
 sg13g2_xnor2_1 _28526_ (.Y(_19965_),
    .A(\u_inv.f_next[203] ),
    .B(\u_inv.f_reg[203] ));
 sg13g2_nor2_1 _28527_ (.A(_19961_),
    .B(_19965_),
    .Y(_19966_));
 sg13g2_nand2_1 _28528_ (.Y(_19967_),
    .A(_19962_),
    .B(_19964_));
 sg13g2_and2_1 _28529_ (.A(\u_inv.f_next[200] ),
    .B(\u_inv.f_reg[200] ),
    .X(_19968_));
 sg13g2_a21oi_1 _28530_ (.A1(\u_inv.f_next[201] ),
    .A2(\u_inv.f_reg[201] ),
    .Y(_19969_),
    .B1(_19968_));
 sg13g2_a21oi_1 _28531_ (.A1(_17991_),
    .A2(_18245_),
    .Y(_19970_),
    .B1(_19969_));
 sg13g2_a22oi_1 _28532_ (.Y(_19971_),
    .B1(_19966_),
    .B2(_19970_),
    .A2(\u_inv.f_reg[203] ),
    .A1(\u_inv.f_next[203] ));
 sg13g2_o21ai_1 _28533_ (.B1(_19971_),
    .Y(_19972_),
    .A1(_19960_),
    .A2(_19963_));
 sg13g2_o21ai_1 _28534_ (.B1(_19949_),
    .Y(_19973_),
    .A1(\u_inv.f_next[207] ),
    .A2(\u_inv.f_reg[207] ));
 sg13g2_a21oi_1 _28535_ (.A1(_17988_),
    .A2(_18246_),
    .Y(_19974_),
    .B1(_19953_));
 sg13g2_a21oi_1 _28536_ (.A1(\u_inv.f_next[205] ),
    .A2(\u_inv.f_reg[205] ),
    .Y(_19975_),
    .B1(_19974_));
 sg13g2_inv_1 _28537_ (.Y(_19976_),
    .A(_19975_));
 sg13g2_a22oi_1 _28538_ (.Y(_19977_),
    .B1(_19976_),
    .B2(_19952_),
    .A2(_19972_),
    .A1(_19958_));
 sg13g2_nand2_1 _28539_ (.Y(_19978_),
    .A(\u_inv.f_next[199] ),
    .B(\u_inv.f_reg[199] ));
 sg13g2_xnor2_1 _28540_ (.Y(_19979_),
    .A(\u_inv.f_next[199] ),
    .B(\u_inv.f_reg[199] ));
 sg13g2_and2_1 _28541_ (.A(\u_inv.f_next[198] ),
    .B(\u_inv.f_reg[198] ),
    .X(_19980_));
 sg13g2_xnor2_1 _28542_ (.Y(_19981_),
    .A(\u_inv.f_next[198] ),
    .B(\u_inv.f_reg[198] ));
 sg13g2_inv_2 _28543_ (.Y(_19982_),
    .A(_19981_));
 sg13g2_xor2_1 _28544_ (.B(\u_inv.f_reg[197] ),
    .A(\u_inv.f_next[197] ),
    .X(_19983_));
 sg13g2_xnor2_1 _28545_ (.Y(_19984_),
    .A(\u_inv.f_next[197] ),
    .B(\u_inv.f_reg[197] ));
 sg13g2_xor2_1 _28546_ (.B(\u_inv.f_reg[196] ),
    .A(\u_inv.f_next[196] ),
    .X(_19985_));
 sg13g2_xnor2_1 _28547_ (.Y(_19986_),
    .A(\u_inv.f_next[196] ),
    .B(\u_inv.f_reg[196] ));
 sg13g2_nor2_1 _28548_ (.A(_19984_),
    .B(_19986_),
    .Y(_19987_));
 sg13g2_nand3b_1 _28549_ (.B(_19982_),
    .C(_19987_),
    .Y(_19988_),
    .A_N(_19979_));
 sg13g2_xnor2_1 _28550_ (.Y(_19989_),
    .A(\u_inv.f_next[194] ),
    .B(\u_inv.f_reg[194] ));
 sg13g2_xnor2_1 _28551_ (.Y(_19990_),
    .A(\u_inv.f_next[195] ),
    .B(\u_inv.f_reg[195] ));
 sg13g2_or2_1 _28552_ (.X(_19991_),
    .B(_19990_),
    .A(_19989_));
 sg13g2_a22oi_1 _28553_ (.Y(_19992_),
    .B1(\u_inv.f_reg[193] ),
    .B2(\u_inv.f_next[193] ),
    .A2(\u_inv.f_reg[192] ),
    .A1(\u_inv.f_next[192] ));
 sg13g2_inv_1 _28554_ (.Y(_19993_),
    .A(_19992_));
 sg13g2_o21ai_1 _28555_ (.B1(_19993_),
    .Y(_19994_),
    .A1(\u_inv.f_next[193] ),
    .A2(\u_inv.f_reg[193] ));
 sg13g2_nor2_1 _28556_ (.A(_19991_),
    .B(_19994_),
    .Y(_19995_));
 sg13g2_a22oi_1 _28557_ (.Y(_19996_),
    .B1(\u_inv.f_reg[195] ),
    .B2(\u_inv.f_next[195] ),
    .A2(\u_inv.f_reg[194] ),
    .A1(\u_inv.f_next[194] ));
 sg13g2_a21oi_2 _28558_ (.B1(_19996_),
    .Y(_19997_),
    .A2(_18243_),
    .A1(_17995_));
 sg13g2_nor2_1 _28559_ (.A(_19995_),
    .B(_19997_),
    .Y(_19998_));
 sg13g2_or2_1 _28560_ (.X(_19999_),
    .B(_19998_),
    .A(_19988_));
 sg13g2_o21ai_1 _28561_ (.B1(_19980_),
    .Y(_20000_),
    .A1(\u_inv.f_next[199] ),
    .A2(\u_inv.f_reg[199] ));
 sg13g2_a22oi_1 _28562_ (.Y(_20001_),
    .B1(\u_inv.f_reg[197] ),
    .B2(\u_inv.f_next[197] ),
    .A2(\u_inv.f_reg[196] ),
    .A1(\u_inv.f_next[196] ));
 sg13g2_inv_1 _28563_ (.Y(_20002_),
    .A(_20001_));
 sg13g2_o21ai_1 _28564_ (.B1(_20002_),
    .Y(_20003_),
    .A1(\u_inv.f_next[197] ),
    .A2(\u_inv.f_reg[197] ));
 sg13g2_or3_1 _28565_ (.A(_19979_),
    .B(_19981_),
    .C(_20003_),
    .X(_20004_));
 sg13g2_nand4_1 _28566_ (.B(_19999_),
    .C(_20000_),
    .A(_19978_),
    .Y(_20005_),
    .D(_20004_));
 sg13g2_inv_2 _28567_ (.Y(_20006_),
    .A(_20005_));
 sg13g2_xnor2_1 _28568_ (.Y(_20007_),
    .A(\u_inv.f_next[201] ),
    .B(\u_inv.f_reg[201] ));
 sg13g2_xor2_1 _28569_ (.B(\u_inv.f_reg[200] ),
    .A(\u_inv.f_next[200] ),
    .X(_20008_));
 sg13g2_xnor2_1 _28570_ (.Y(_20009_),
    .A(\u_inv.f_next[200] ),
    .B(\u_inv.f_reg[200] ));
 sg13g2_nand2b_1 _28571_ (.Y(_20010_),
    .B(_20008_),
    .A_N(_20007_));
 sg13g2_nor2_1 _28572_ (.A(_19967_),
    .B(_20010_),
    .Y(_20011_));
 sg13g2_inv_1 _28573_ (.Y(_20012_),
    .A(_20011_));
 sg13g2_nor3_1 _28574_ (.A(_19959_),
    .B(_19967_),
    .C(_20010_),
    .Y(_20013_));
 sg13g2_nand2_1 _28575_ (.Y(_20014_),
    .A(_20005_),
    .B(_20013_));
 sg13g2_nand4_1 _28576_ (.B(_19973_),
    .C(_19977_),
    .A(_19947_),
    .Y(_20015_),
    .D(_20014_));
 sg13g2_inv_2 _28577_ (.Y(_20016_),
    .A(_20015_));
 sg13g2_xor2_1 _28578_ (.B(\u_inv.f_reg[191] ),
    .A(\u_inv.f_next[191] ),
    .X(_20017_));
 sg13g2_xnor2_1 _28579_ (.Y(_20018_),
    .A(\u_inv.f_next[191] ),
    .B(\u_inv.f_reg[191] ));
 sg13g2_and2_1 _28580_ (.A(\u_inv.f_next[190] ),
    .B(\u_inv.f_reg[190] ),
    .X(_20019_));
 sg13g2_nand2_1 _28581_ (.Y(_20020_),
    .A(\u_inv.f_next[190] ),
    .B(\u_inv.f_reg[190] ));
 sg13g2_xor2_1 _28582_ (.B(\u_inv.f_reg[190] ),
    .A(\u_inv.f_next[190] ),
    .X(_20021_));
 sg13g2_inv_1 _28583_ (.Y(_20022_),
    .A(_20021_));
 sg13g2_nand2_1 _28584_ (.Y(_20023_),
    .A(_20017_),
    .B(_20021_));
 sg13g2_nand2_1 _28585_ (.Y(_20024_),
    .A(\u_inv.f_next[189] ),
    .B(\u_inv.f_reg[189] ));
 sg13g2_or2_1 _28586_ (.X(_20025_),
    .B(\u_inv.f_reg[189] ),
    .A(\u_inv.f_next[189] ));
 sg13g2_and2_1 _28587_ (.A(_20024_),
    .B(_20025_),
    .X(_20026_));
 sg13g2_nand2_2 _28588_ (.Y(_20027_),
    .A(_20024_),
    .B(_20025_));
 sg13g2_nand2_1 _28589_ (.Y(_20028_),
    .A(\u_inv.f_next[188] ),
    .B(\u_inv.f_reg[188] ));
 sg13g2_xor2_1 _28590_ (.B(\u_inv.f_reg[188] ),
    .A(\u_inv.f_next[188] ),
    .X(_20029_));
 sg13g2_and2_1 _28591_ (.A(_20026_),
    .B(_20029_),
    .X(_20030_));
 sg13g2_nand2b_1 _28592_ (.Y(_20031_),
    .B(_20030_),
    .A_N(_20023_));
 sg13g2_xor2_1 _28593_ (.B(\u_inv.f_reg[185] ),
    .A(\u_inv.f_next[185] ),
    .X(_20032_));
 sg13g2_xnor2_1 _28594_ (.Y(_20033_),
    .A(\u_inv.f_next[185] ),
    .B(\u_inv.f_reg[185] ));
 sg13g2_nand2_1 _28595_ (.Y(_20034_),
    .A(\u_inv.f_next[184] ),
    .B(\u_inv.f_reg[184] ));
 sg13g2_xnor2_1 _28596_ (.Y(_20035_),
    .A(\u_inv.f_next[184] ),
    .B(\u_inv.f_reg[184] ));
 sg13g2_or2_1 _28597_ (.X(_20036_),
    .B(_20035_),
    .A(_20033_));
 sg13g2_and2_1 _28598_ (.A(\u_inv.f_next[186] ),
    .B(\u_inv.f_reg[186] ),
    .X(_20037_));
 sg13g2_xor2_1 _28599_ (.B(\u_inv.f_reg[186] ),
    .A(\u_inv.f_next[186] ),
    .X(_20038_));
 sg13g2_xnor2_1 _28600_ (.Y(_20039_),
    .A(\u_inv.f_next[186] ),
    .B(\u_inv.f_reg[186] ));
 sg13g2_nand2_1 _28601_ (.Y(_20040_),
    .A(\u_inv.f_next[187] ),
    .B(\u_inv.f_reg[187] ));
 sg13g2_xor2_1 _28602_ (.B(\u_inv.f_reg[187] ),
    .A(\u_inv.f_next[187] ),
    .X(_20041_));
 sg13g2_nand2_1 _28603_ (.Y(_20042_),
    .A(_20038_),
    .B(_20041_));
 sg13g2_nor2_1 _28604_ (.A(_18005_),
    .B(_18238_),
    .Y(_20043_));
 sg13g2_nand2_1 _28605_ (.Y(_20044_),
    .A(_18005_),
    .B(_18238_));
 sg13g2_nor2b_2 _28606_ (.A(_20043_),
    .B_N(_20044_),
    .Y(_20045_));
 sg13g2_and2_1 _28607_ (.A(\u_inv.f_next[182] ),
    .B(\u_inv.f_reg[182] ),
    .X(_20046_));
 sg13g2_xor2_1 _28608_ (.B(\u_inv.f_reg[182] ),
    .A(\u_inv.f_next[182] ),
    .X(_20047_));
 sg13g2_xnor2_1 _28609_ (.Y(_20048_),
    .A(\u_inv.f_next[182] ),
    .B(\u_inv.f_reg[182] ));
 sg13g2_nand2_1 _28610_ (.Y(_20049_),
    .A(_20045_),
    .B(_20047_));
 sg13g2_nand2_1 _28611_ (.Y(_20050_),
    .A(\u_inv.f_next[180] ),
    .B(\u_inv.f_reg[180] ));
 sg13g2_xor2_1 _28612_ (.B(\u_inv.f_reg[180] ),
    .A(\u_inv.f_next[180] ),
    .X(_20051_));
 sg13g2_xnor2_1 _28613_ (.Y(_20052_),
    .A(\u_inv.f_next[180] ),
    .B(\u_inv.f_reg[180] ));
 sg13g2_nand2_1 _28614_ (.Y(_20053_),
    .A(\u_inv.f_next[181] ),
    .B(\u_inv.f_reg[181] ));
 sg13g2_xor2_1 _28615_ (.B(\u_inv.f_reg[181] ),
    .A(\u_inv.f_next[181] ),
    .X(_20054_));
 sg13g2_nand2_1 _28616_ (.Y(_20055_),
    .A(_20051_),
    .B(_20054_));
 sg13g2_nor2_1 _28617_ (.A(_20049_),
    .B(_20055_),
    .Y(_20056_));
 sg13g2_nand2_1 _28618_ (.Y(_20057_),
    .A(\u_inv.f_next[178] ),
    .B(\u_inv.f_reg[178] ));
 sg13g2_xor2_1 _28619_ (.B(\u_inv.f_reg[178] ),
    .A(\u_inv.f_next[178] ),
    .X(_20058_));
 sg13g2_xnor2_1 _28620_ (.Y(_20059_),
    .A(\u_inv.f_next[178] ),
    .B(\u_inv.f_reg[178] ));
 sg13g2_xor2_1 _28621_ (.B(\u_inv.f_reg[179] ),
    .A(\u_inv.f_next[179] ),
    .X(_20060_));
 sg13g2_xnor2_1 _28622_ (.Y(_20061_),
    .A(\u_inv.f_next[179] ),
    .B(\u_inv.f_reg[179] ));
 sg13g2_a22oi_1 _28623_ (.Y(_20062_),
    .B1(\u_inv.f_reg[177] ),
    .B2(\u_inv.f_next[177] ),
    .A2(\u_inv.f_reg[176] ),
    .A1(\u_inv.f_next[176] ));
 sg13g2_a21oi_1 _28624_ (.A1(_18008_),
    .A2(_18236_),
    .Y(_20063_),
    .B1(_20062_));
 sg13g2_nand3_1 _28625_ (.B(_20060_),
    .C(_20063_),
    .A(_20058_),
    .Y(_20064_));
 sg13g2_a21oi_1 _28626_ (.A1(_18007_),
    .A2(_18237_),
    .Y(_20065_),
    .B1(_20057_));
 sg13g2_a21oi_1 _28627_ (.A1(\u_inv.f_next[179] ),
    .A2(\u_inv.f_reg[179] ),
    .Y(_20066_),
    .B1(_20065_));
 sg13g2_nand2_1 _28628_ (.Y(_20067_),
    .A(_20064_),
    .B(_20066_));
 sg13g2_nand2_1 _28629_ (.Y(_20068_),
    .A(_20050_),
    .B(_20053_));
 sg13g2_o21ai_1 _28630_ (.B1(_20068_),
    .Y(_20069_),
    .A1(\u_inv.f_next[181] ),
    .A2(\u_inv.f_reg[181] ));
 sg13g2_a221oi_1 _28631_ (.B2(_20067_),
    .C1(_20043_),
    .B1(_20056_),
    .A1(_20044_),
    .Y(_20070_),
    .A2(_20046_));
 sg13g2_o21ai_1 _28632_ (.B1(_20070_),
    .Y(_20071_),
    .A1(_20049_),
    .A2(_20069_));
 sg13g2_nand2_1 _28633_ (.Y(_20072_),
    .A(_20024_),
    .B(_20028_));
 sg13g2_nand2_1 _28634_ (.Y(_20073_),
    .A(_20025_),
    .B(_20072_));
 sg13g2_a21oi_1 _28635_ (.A1(_17998_),
    .A2(_18241_),
    .Y(_20074_),
    .B1(_20020_));
 sg13g2_a21oi_1 _28636_ (.A1(\u_inv.f_next[191] ),
    .A2(\u_inv.f_reg[191] ),
    .Y(_20075_),
    .B1(_20074_));
 sg13g2_a21oi_1 _28637_ (.A1(_18003_),
    .A2(_18239_),
    .Y(_20076_),
    .B1(_20034_));
 sg13g2_a21oi_1 _28638_ (.A1(\u_inv.f_next[185] ),
    .A2(\u_inv.f_reg[185] ),
    .Y(_20077_),
    .B1(_20076_));
 sg13g2_o21ai_1 _28639_ (.B1(_20037_),
    .Y(_20078_),
    .A1(\u_inv.f_next[187] ),
    .A2(\u_inv.f_reg[187] ));
 sg13g2_o21ai_1 _28640_ (.B1(_20040_),
    .Y(_20079_),
    .A1(_20042_),
    .A2(_20077_));
 sg13g2_nor2b_1 _28641_ (.A(_20079_),
    .B_N(_20078_),
    .Y(_20080_));
 sg13g2_inv_1 _28642_ (.Y(_20081_),
    .A(_20080_));
 sg13g2_nor3_1 _28643_ (.A(_20031_),
    .B(_20036_),
    .C(_20042_),
    .Y(_20082_));
 sg13g2_o21ai_1 _28644_ (.B1(_20075_),
    .Y(_20083_),
    .A1(_20031_),
    .A2(_20080_));
 sg13g2_a21oi_1 _28645_ (.A1(_20071_),
    .A2(_20082_),
    .Y(_20084_),
    .B1(_20083_));
 sg13g2_o21ai_1 _28646_ (.B1(_20084_),
    .Y(_20085_),
    .A1(_20023_),
    .A2(_20073_));
 sg13g2_inv_1 _28647_ (.Y(_20086_),
    .A(_20085_));
 sg13g2_xor2_1 _28648_ (.B(\u_inv.f_reg[175] ),
    .A(\u_inv.f_next[175] ),
    .X(_20087_));
 sg13g2_xnor2_1 _28649_ (.Y(_20088_),
    .A(\u_inv.f_next[175] ),
    .B(\u_inv.f_reg[175] ));
 sg13g2_nand2_1 _28650_ (.Y(_20089_),
    .A(\u_inv.f_next[174] ),
    .B(\u_inv.f_reg[174] ));
 sg13g2_xnor2_1 _28651_ (.Y(_20090_),
    .A(\u_inv.f_next[174] ),
    .B(\u_inv.f_reg[174] ));
 sg13g2_nor2_1 _28652_ (.A(_20088_),
    .B(_20090_),
    .Y(_20091_));
 sg13g2_nand2_1 _28653_ (.Y(_20092_),
    .A(\u_inv.f_next[172] ),
    .B(\u_inv.f_reg[172] ));
 sg13g2_a22oi_1 _28654_ (.Y(_20093_),
    .B1(\u_inv.f_reg[173] ),
    .B2(\u_inv.f_next[173] ),
    .A2(\u_inv.f_reg[172] ),
    .A1(\u_inv.f_next[172] ));
 sg13g2_a21o_1 _28655_ (.A2(_18234_),
    .A1(_18012_),
    .B1(_20093_),
    .X(_20094_));
 sg13g2_xnor2_1 _28656_ (.Y(_20095_),
    .A(\u_inv.f_next[172] ),
    .B(\u_inv.f_reg[172] ));
 sg13g2_inv_1 _28657_ (.Y(_20096_),
    .A(_20095_));
 sg13g2_xor2_1 _28658_ (.B(\u_inv.f_reg[173] ),
    .A(\u_inv.f_next[173] ),
    .X(_20097_));
 sg13g2_nor2b_1 _28659_ (.A(_20095_),
    .B_N(_20097_),
    .Y(_20098_));
 sg13g2_and2_1 _28660_ (.A(\u_inv.f_next[170] ),
    .B(\u_inv.f_reg[170] ),
    .X(_20099_));
 sg13g2_a21oi_1 _28661_ (.A1(\u_inv.f_next[171] ),
    .A2(\u_inv.f_reg[171] ),
    .Y(_20100_),
    .B1(_20099_));
 sg13g2_a21oi_1 _28662_ (.A1(_18013_),
    .A2(_18233_),
    .Y(_20101_),
    .B1(_20100_));
 sg13g2_xor2_1 _28663_ (.B(\u_inv.f_reg[170] ),
    .A(\u_inv.f_next[170] ),
    .X(_20102_));
 sg13g2_nor2_1 _28664_ (.A(_18013_),
    .B(\u_inv.f_reg[171] ),
    .Y(_20103_));
 sg13g2_xnor2_1 _28665_ (.Y(_20104_),
    .A(\u_inv.f_next[171] ),
    .B(\u_inv.f_reg[171] ));
 sg13g2_xor2_1 _28666_ (.B(\u_inv.f_reg[171] ),
    .A(\u_inv.f_next[171] ),
    .X(_20105_));
 sg13g2_and2_1 _28667_ (.A(_20102_),
    .B(_20105_),
    .X(_20106_));
 sg13g2_inv_1 _28668_ (.Y(_20107_),
    .A(_20106_));
 sg13g2_nand2_1 _28669_ (.Y(_20108_),
    .A(\u_inv.f_next[169] ),
    .B(\u_inv.f_reg[169] ));
 sg13g2_xor2_1 _28670_ (.B(\u_inv.f_reg[169] ),
    .A(\u_inv.f_next[169] ),
    .X(_20109_));
 sg13g2_nand2_1 _28671_ (.Y(_20110_),
    .A(\u_inv.f_next[168] ),
    .B(\u_inv.f_reg[168] ));
 sg13g2_xor2_1 _28672_ (.B(\u_inv.f_reg[168] ),
    .A(\u_inv.f_next[168] ),
    .X(_20111_));
 sg13g2_xnor2_1 _28673_ (.Y(_20112_),
    .A(\u_inv.f_next[168] ),
    .B(\u_inv.f_reg[168] ));
 sg13g2_nand2_1 _28674_ (.Y(_20113_),
    .A(_20109_),
    .B(_20111_));
 sg13g2_inv_1 _28675_ (.Y(_20114_),
    .A(_20113_));
 sg13g2_nor2_1 _28676_ (.A(\u_inv.f_next[167] ),
    .B(\u_inv.f_reg[167] ),
    .Y(_20115_));
 sg13g2_xor2_1 _28677_ (.B(\u_inv.f_reg[167] ),
    .A(\u_inv.f_next[167] ),
    .X(_20116_));
 sg13g2_nand2_1 _28678_ (.Y(_20117_),
    .A(\u_inv.f_next[166] ),
    .B(\u_inv.f_reg[166] ));
 sg13g2_xor2_1 _28679_ (.B(\u_inv.f_reg[166] ),
    .A(\u_inv.f_next[166] ),
    .X(_20118_));
 sg13g2_xnor2_1 _28680_ (.Y(_20119_),
    .A(\u_inv.f_next[166] ),
    .B(\u_inv.f_reg[166] ));
 sg13g2_and2_1 _28681_ (.A(_20116_),
    .B(_20118_),
    .X(_20120_));
 sg13g2_nor2_1 _28682_ (.A(\u_inv.f_next[165] ),
    .B(\u_inv.f_reg[165] ),
    .Y(_20121_));
 sg13g2_nand2_1 _28683_ (.Y(_20122_),
    .A(\u_inv.f_next[165] ),
    .B(\u_inv.f_reg[165] ));
 sg13g2_nand2_1 _28684_ (.Y(_20123_),
    .A(\u_inv.f_next[164] ),
    .B(\u_inv.f_reg[164] ));
 sg13g2_o21ai_1 _28685_ (.B1(_20122_),
    .Y(_20124_),
    .A1(_20121_),
    .A2(_20123_));
 sg13g2_a22oi_1 _28686_ (.Y(_20125_),
    .B1(_20120_),
    .B2(_20124_),
    .A2(\u_inv.f_reg[167] ),
    .A1(\u_inv.f_next[167] ));
 sg13g2_o21ai_1 _28687_ (.B1(_20125_),
    .Y(_20126_),
    .A1(_20115_),
    .A2(_20117_));
 sg13g2_xor2_1 _28688_ (.B(\u_inv.f_reg[164] ),
    .A(\u_inv.f_next[164] ),
    .X(_20127_));
 sg13g2_xnor2_1 _28689_ (.Y(_20128_),
    .A(\u_inv.f_next[164] ),
    .B(\u_inv.f_reg[164] ));
 sg13g2_nor2b_2 _28690_ (.A(_20121_),
    .B_N(_20122_),
    .Y(_20129_));
 sg13g2_nand2b_1 _28691_ (.Y(_20130_),
    .B(_20122_),
    .A_N(_20121_));
 sg13g2_nor2_1 _28692_ (.A(_20128_),
    .B(_20130_),
    .Y(_20131_));
 sg13g2_and2_1 _28693_ (.A(_20120_),
    .B(_20131_),
    .X(_20132_));
 sg13g2_inv_1 _28694_ (.Y(_20133_),
    .A(_20132_));
 sg13g2_and2_1 _28695_ (.A(\u_inv.f_next[162] ),
    .B(\u_inv.f_reg[162] ),
    .X(_20134_));
 sg13g2_xor2_1 _28696_ (.B(\u_inv.f_reg[162] ),
    .A(\u_inv.f_next[162] ),
    .X(_20135_));
 sg13g2_nand2_1 _28697_ (.Y(_20136_),
    .A(_18017_),
    .B(_18231_));
 sg13g2_nand2_1 _28698_ (.Y(_20137_),
    .A(\u_inv.f_next[163] ),
    .B(\u_inv.f_reg[163] ));
 sg13g2_and2_1 _28699_ (.A(_20136_),
    .B(_20137_),
    .X(_20138_));
 sg13g2_nand2_1 _28700_ (.Y(_20139_),
    .A(_20135_),
    .B(_20138_));
 sg13g2_nand2_1 _28701_ (.Y(_20140_),
    .A(\u_inv.f_next[160] ),
    .B(\u_inv.f_reg[160] ));
 sg13g2_a21oi_1 _28702_ (.A1(_18019_),
    .A2(_18230_),
    .Y(_20141_),
    .B1(_20140_));
 sg13g2_a21oi_1 _28703_ (.A1(\u_inv.f_next[161] ),
    .A2(\u_inv.f_reg[161] ),
    .Y(_20142_),
    .B1(_20141_));
 sg13g2_o21ai_1 _28704_ (.B1(_20137_),
    .Y(_20143_),
    .A1(_20139_),
    .A2(_20142_));
 sg13g2_a21oi_2 _28705_ (.B1(_20143_),
    .Y(_20144_),
    .A2(_20136_),
    .A1(_20134_));
 sg13g2_inv_1 _28706_ (.Y(_20145_),
    .A(_20144_));
 sg13g2_a21oi_1 _28707_ (.A1(_20132_),
    .A2(_20145_),
    .Y(_20146_),
    .B1(_20126_));
 sg13g2_nand2_1 _28708_ (.Y(_20147_),
    .A(_20108_),
    .B(_20110_));
 sg13g2_o21ai_1 _28709_ (.B1(_20147_),
    .Y(_20148_),
    .A1(\u_inv.f_next[169] ),
    .A2(\u_inv.f_reg[169] ));
 sg13g2_o21ai_1 _28710_ (.B1(_20148_),
    .Y(_20149_),
    .A1(_20113_),
    .A2(_20146_));
 sg13g2_and2_1 _28711_ (.A(_20098_),
    .B(_20106_),
    .X(_20150_));
 sg13g2_a22oi_1 _28712_ (.Y(_20151_),
    .B1(_20149_),
    .B2(_20150_),
    .A2(_20101_),
    .A1(_20098_));
 sg13g2_nand2_1 _28713_ (.Y(_20152_),
    .A(_20094_),
    .B(_20151_));
 sg13g2_a21oi_1 _28714_ (.A1(_18010_),
    .A2(_18235_),
    .Y(_20153_),
    .B1(_20089_));
 sg13g2_a221oi_1 _28715_ (.B2(_20152_),
    .C1(_20153_),
    .B1(_20091_),
    .A1(\u_inv.f_next[175] ),
    .Y(_20154_),
    .A2(\u_inv.f_reg[175] ));
 sg13g2_nor2_1 _28716_ (.A(\u_inv.f_next[159] ),
    .B(\u_inv.f_reg[159] ),
    .Y(_20155_));
 sg13g2_xor2_1 _28717_ (.B(\u_inv.f_reg[159] ),
    .A(\u_inv.f_next[159] ),
    .X(_20156_));
 sg13g2_nand2_1 _28718_ (.Y(_20157_),
    .A(\u_inv.f_next[158] ),
    .B(\u_inv.f_reg[158] ));
 sg13g2_xor2_1 _28719_ (.B(\u_inv.f_reg[158] ),
    .A(\u_inv.f_next[158] ),
    .X(_20158_));
 sg13g2_xnor2_1 _28720_ (.Y(_20159_),
    .A(\u_inv.f_next[158] ),
    .B(\u_inv.f_reg[158] ));
 sg13g2_and2_1 _28721_ (.A(_20156_),
    .B(_20158_),
    .X(_20160_));
 sg13g2_nor2_1 _28722_ (.A(\u_inv.f_next[157] ),
    .B(\u_inv.f_reg[157] ),
    .Y(_20161_));
 sg13g2_xor2_1 _28723_ (.B(\u_inv.f_reg[157] ),
    .A(\u_inv.f_next[157] ),
    .X(_20162_));
 sg13g2_xnor2_1 _28724_ (.Y(_20163_),
    .A(\u_inv.f_next[157] ),
    .B(\u_inv.f_reg[157] ));
 sg13g2_and2_1 _28725_ (.A(\u_inv.f_next[156] ),
    .B(\u_inv.f_reg[156] ),
    .X(_20164_));
 sg13g2_xnor2_1 _28726_ (.Y(_20165_),
    .A(\u_inv.f_next[156] ),
    .B(\u_inv.f_reg[156] ));
 sg13g2_nor2_1 _28727_ (.A(_20163_),
    .B(_20165_),
    .Y(_20166_));
 sg13g2_and2_1 _28728_ (.A(_20160_),
    .B(_20166_),
    .X(_20167_));
 sg13g2_inv_1 _28729_ (.Y(_20168_),
    .A(_20167_));
 sg13g2_xor2_1 _28730_ (.B(\u_inv.f_reg[153] ),
    .A(\u_inv.f_next[153] ),
    .X(_20169_));
 sg13g2_xnor2_1 _28731_ (.Y(_20170_),
    .A(\u_inv.f_next[153] ),
    .B(\u_inv.f_reg[153] ));
 sg13g2_and2_1 _28732_ (.A(\u_inv.f_next[152] ),
    .B(\u_inv.f_reg[152] ),
    .X(_20171_));
 sg13g2_xor2_1 _28733_ (.B(\u_inv.f_reg[152] ),
    .A(\u_inv.f_next[152] ),
    .X(_20172_));
 sg13g2_xnor2_1 _28734_ (.Y(_20173_),
    .A(\u_inv.f_next[152] ),
    .B(\u_inv.f_reg[152] ));
 sg13g2_nand2_1 _28735_ (.Y(_20174_),
    .A(_20169_),
    .B(_20172_));
 sg13g2_nand2_1 _28736_ (.Y(_20175_),
    .A(\u_inv.f_next[154] ),
    .B(\u_inv.f_reg[154] ));
 sg13g2_xor2_1 _28737_ (.B(\u_inv.f_reg[154] ),
    .A(\u_inv.f_next[154] ),
    .X(_20176_));
 sg13g2_nand2_1 _28738_ (.Y(_20177_),
    .A(\u_inv.f_next[155] ),
    .B(\u_inv.f_reg[155] ));
 sg13g2_xor2_1 _28739_ (.B(\u_inv.f_reg[155] ),
    .A(\u_inv.f_next[155] ),
    .X(_20178_));
 sg13g2_nand2_1 _28740_ (.Y(_20179_),
    .A(_20176_),
    .B(_20178_));
 sg13g2_or2_1 _28741_ (.X(_20180_),
    .B(_20179_),
    .A(_20174_));
 sg13g2_nor2_1 _28742_ (.A(_20168_),
    .B(_20180_),
    .Y(_20181_));
 sg13g2_xor2_1 _28743_ (.B(\u_inv.f_reg[149] ),
    .A(\u_inv.f_next[149] ),
    .X(_20182_));
 sg13g2_xnor2_1 _28744_ (.Y(_20183_),
    .A(\u_inv.f_next[149] ),
    .B(\u_inv.f_reg[149] ));
 sg13g2_and2_1 _28745_ (.A(\u_inv.f_next[148] ),
    .B(\u_inv.f_reg[148] ),
    .X(_20184_));
 sg13g2_xor2_1 _28746_ (.B(\u_inv.f_reg[148] ),
    .A(\u_inv.f_next[148] ),
    .X(_20185_));
 sg13g2_xnor2_1 _28747_ (.Y(_20186_),
    .A(\u_inv.f_next[148] ),
    .B(\u_inv.f_reg[148] ));
 sg13g2_nor2_1 _28748_ (.A(_20183_),
    .B(_20186_),
    .Y(_20187_));
 sg13g2_nor2_1 _28749_ (.A(\u_inv.f_next[151] ),
    .B(\u_inv.f_reg[151] ),
    .Y(_20188_));
 sg13g2_xor2_1 _28750_ (.B(\u_inv.f_reg[151] ),
    .A(\u_inv.f_next[151] ),
    .X(_20189_));
 sg13g2_xnor2_1 _28751_ (.Y(_20190_),
    .A(\u_inv.f_next[151] ),
    .B(\u_inv.f_reg[151] ));
 sg13g2_nand2_1 _28752_ (.Y(_20191_),
    .A(\u_inv.f_next[150] ),
    .B(\u_inv.f_reg[150] ));
 sg13g2_xnor2_1 _28753_ (.Y(_20192_),
    .A(\u_inv.f_next[150] ),
    .B(\u_inv.f_reg[150] ));
 sg13g2_nor2_1 _28754_ (.A(_20190_),
    .B(_20192_),
    .Y(_20193_));
 sg13g2_and2_1 _28755_ (.A(_20187_),
    .B(_20193_),
    .X(_20194_));
 sg13g2_xnor2_1 _28756_ (.Y(_20195_),
    .A(\u_inv.f_next[147] ),
    .B(\u_inv.f_reg[147] ));
 sg13g2_xor2_1 _28757_ (.B(\u_inv.f_reg[147] ),
    .A(\u_inv.f_next[147] ),
    .X(_20196_));
 sg13g2_nand2_1 _28758_ (.Y(_20197_),
    .A(\u_inv.f_next[146] ),
    .B(\u_inv.f_reg[146] ));
 sg13g2_xor2_1 _28759_ (.B(\u_inv.f_reg[146] ),
    .A(\u_inv.f_next[146] ),
    .X(_20198_));
 sg13g2_nand2_1 _28760_ (.Y(_20199_),
    .A(_20196_),
    .B(_20198_));
 sg13g2_inv_1 _28761_ (.Y(_20200_),
    .A(_20199_));
 sg13g2_nor2_1 _28762_ (.A(\u_inv.f_next[145] ),
    .B(\u_inv.f_reg[145] ),
    .Y(_20201_));
 sg13g2_nand2_1 _28763_ (.Y(_20202_),
    .A(\u_inv.f_next[145] ),
    .B(\u_inv.f_reg[145] ));
 sg13g2_and2_1 _28764_ (.A(\u_inv.f_next[144] ),
    .B(\u_inv.f_reg[144] ),
    .X(_20203_));
 sg13g2_nand2_1 _28765_ (.Y(_20204_),
    .A(\u_inv.f_next[144] ),
    .B(\u_inv.f_reg[144] ));
 sg13g2_o21ai_1 _28766_ (.B1(_20202_),
    .Y(_20205_),
    .A1(_20201_),
    .A2(_20204_));
 sg13g2_inv_1 _28767_ (.Y(_20206_),
    .A(_20205_));
 sg13g2_a21oi_1 _28768_ (.A1(_18026_),
    .A2(_18227_),
    .Y(_20207_),
    .B1(_20197_));
 sg13g2_a21oi_1 _28769_ (.A1(\u_inv.f_next[147] ),
    .A2(\u_inv.f_reg[147] ),
    .Y(_20208_),
    .B1(_20207_));
 sg13g2_o21ai_1 _28770_ (.B1(_20208_),
    .Y(_20209_),
    .A1(_20199_),
    .A2(_20206_));
 sg13g2_nor2_1 _28771_ (.A(_20188_),
    .B(_20191_),
    .Y(_20210_));
 sg13g2_a21oi_1 _28772_ (.A1(\u_inv.f_next[151] ),
    .A2(\u_inv.f_reg[151] ),
    .Y(_20211_),
    .B1(_20210_));
 sg13g2_a21oi_1 _28773_ (.A1(\u_inv.f_next[149] ),
    .A2(\u_inv.f_reg[149] ),
    .Y(_20212_),
    .B1(_20184_));
 sg13g2_a21oi_1 _28774_ (.A1(_18025_),
    .A2(_18228_),
    .Y(_20213_),
    .B1(_20212_));
 sg13g2_a22oi_1 _28775_ (.Y(_20214_),
    .B1(_20213_),
    .B2(_20193_),
    .A2(_20209_),
    .A1(_20194_));
 sg13g2_nand2_2 _28776_ (.Y(_20215_),
    .A(_20211_),
    .B(_20214_));
 sg13g2_a21oi_1 _28777_ (.A1(\u_inv.f_next[157] ),
    .A2(\u_inv.f_reg[157] ),
    .Y(_20216_),
    .B1(_20164_));
 sg13g2_nor2_1 _28778_ (.A(_20161_),
    .B(_20216_),
    .Y(_20217_));
 sg13g2_nor2_1 _28779_ (.A(_20155_),
    .B(_20157_),
    .Y(_20218_));
 sg13g2_a221oi_1 _28780_ (.B2(_20217_),
    .C1(_20218_),
    .B1(_20160_),
    .A1(\u_inv.f_next[159] ),
    .Y(_20219_),
    .A2(\u_inv.f_reg[159] ));
 sg13g2_a21oi_1 _28781_ (.A1(\u_inv.f_next[153] ),
    .A2(\u_inv.f_reg[153] ),
    .Y(_20220_),
    .B1(_20171_));
 sg13g2_inv_1 _28782_ (.Y(_20221_),
    .A(_20220_));
 sg13g2_o21ai_1 _28783_ (.B1(_20221_),
    .Y(_20222_),
    .A1(\u_inv.f_next[153] ),
    .A2(\u_inv.f_reg[153] ));
 sg13g2_a21oi_1 _28784_ (.A1(_18021_),
    .A2(_18229_),
    .Y(_20223_),
    .B1(_20175_));
 sg13g2_o21ai_1 _28785_ (.B1(_20177_),
    .Y(_20224_),
    .A1(_20179_),
    .A2(_20222_));
 sg13g2_nor2_1 _28786_ (.A(_20223_),
    .B(_20224_),
    .Y(_20225_));
 sg13g2_o21ai_1 _28787_ (.B1(_20219_),
    .Y(_20226_),
    .A1(_20168_),
    .A2(_20225_));
 sg13g2_a21o_2 _28788_ (.A2(_20215_),
    .A1(_20181_),
    .B1(_20226_),
    .X(_20227_));
 sg13g2_nand2_1 _28789_ (.Y(_20228_),
    .A(\u_inv.f_next[127] ),
    .B(\u_inv.f_reg[127] ));
 sg13g2_nor2_1 _28790_ (.A(\u_inv.f_next[127] ),
    .B(\u_inv.f_reg[127] ),
    .Y(_20229_));
 sg13g2_xnor2_1 _28791_ (.Y(_20230_),
    .A(\u_inv.f_next[127] ),
    .B(\u_inv.f_reg[127] ));
 sg13g2_nand2_1 _28792_ (.Y(_20231_),
    .A(\u_inv.f_next[126] ),
    .B(\u_inv.f_reg[126] ));
 sg13g2_xor2_1 _28793_ (.B(\u_inv.f_reg[126] ),
    .A(\u_inv.f_next[126] ),
    .X(_20232_));
 sg13g2_xnor2_1 _28794_ (.Y(_20233_),
    .A(\u_inv.f_next[126] ),
    .B(\u_inv.f_reg[126] ));
 sg13g2_nor2_1 _28795_ (.A(_20230_),
    .B(_20233_),
    .Y(_20234_));
 sg13g2_xor2_1 _28796_ (.B(\u_inv.f_reg[124] ),
    .A(\u_inv.f_next[124] ),
    .X(_20235_));
 sg13g2_xnor2_1 _28797_ (.Y(_20236_),
    .A(\u_inv.f_next[124] ),
    .B(\u_inv.f_reg[124] ));
 sg13g2_xnor2_1 _28798_ (.Y(_20237_),
    .A(\u_inv.f_next[125] ),
    .B(\u_inv.f_reg[125] ));
 sg13g2_nor2_1 _28799_ (.A(_20236_),
    .B(_20237_),
    .Y(_20238_));
 sg13g2_nand2_1 _28800_ (.Y(_20239_),
    .A(_20234_),
    .B(_20238_));
 sg13g2_xor2_1 _28801_ (.B(\u_inv.f_reg[121] ),
    .A(\u_inv.f_next[121] ),
    .X(_20240_));
 sg13g2_and2_1 _28802_ (.A(\u_inv.f_next[120] ),
    .B(\u_inv.f_reg[120] ),
    .X(_20241_));
 sg13g2_xor2_1 _28803_ (.B(\u_inv.f_reg[120] ),
    .A(\u_inv.f_next[120] ),
    .X(_20242_));
 sg13g2_nand2_1 _28804_ (.Y(_20243_),
    .A(_20240_),
    .B(_20242_));
 sg13g2_nand2_1 _28805_ (.Y(_20244_),
    .A(\u_inv.f_next[122] ),
    .B(\u_inv.f_reg[122] ));
 sg13g2_xor2_1 _28806_ (.B(\u_inv.f_reg[122] ),
    .A(\u_inv.f_next[122] ),
    .X(_20245_));
 sg13g2_xnor2_1 _28807_ (.Y(_20246_),
    .A(\u_inv.f_next[122] ),
    .B(\u_inv.f_reg[122] ));
 sg13g2_xor2_1 _28808_ (.B(\u_inv.f_reg[123] ),
    .A(\u_inv.f_next[123] ),
    .X(_20247_));
 sg13g2_nand2_1 _28809_ (.Y(_20248_),
    .A(_20245_),
    .B(_20247_));
 sg13g2_inv_1 _28810_ (.Y(_20249_),
    .A(_20248_));
 sg13g2_nor3_1 _28811_ (.A(_20239_),
    .B(_20243_),
    .C(_20248_),
    .Y(_20250_));
 sg13g2_and2_1 _28812_ (.A(\u_inv.f_next[119] ),
    .B(\u_inv.f_reg[119] ),
    .X(_20251_));
 sg13g2_or2_1 _28813_ (.X(_20252_),
    .B(\u_inv.f_reg[119] ),
    .A(\u_inv.f_next[119] ));
 sg13g2_nor2b_2 _28814_ (.A(_20251_),
    .B_N(_20252_),
    .Y(_20253_));
 sg13g2_and2_1 _28815_ (.A(\u_inv.f_next[118] ),
    .B(\u_inv.f_reg[118] ),
    .X(_20254_));
 sg13g2_xnor2_1 _28816_ (.Y(_20255_),
    .A(\u_inv.f_next[118] ),
    .B(\u_inv.f_reg[118] ));
 sg13g2_inv_1 _28817_ (.Y(_20256_),
    .A(_20255_));
 sg13g2_nand2_1 _28818_ (.Y(_20257_),
    .A(_20253_),
    .B(_20256_));
 sg13g2_xor2_1 _28819_ (.B(\u_inv.f_reg[117] ),
    .A(\u_inv.f_next[117] ),
    .X(_20258_));
 sg13g2_nand2_1 _28820_ (.Y(_20259_),
    .A(\u_inv.f_next[116] ),
    .B(\u_inv.f_reg[116] ));
 sg13g2_nor2_1 _28821_ (.A(\u_inv.f_next[116] ),
    .B(\u_inv.f_reg[116] ),
    .Y(_20260_));
 sg13g2_xor2_1 _28822_ (.B(\u_inv.f_reg[116] ),
    .A(\u_inv.f_next[116] ),
    .X(_20261_));
 sg13g2_and2_1 _28823_ (.A(_20258_),
    .B(_20261_),
    .X(_20262_));
 sg13g2_inv_1 _28824_ (.Y(_20263_),
    .A(_20262_));
 sg13g2_nor2_1 _28825_ (.A(_20257_),
    .B(_20263_),
    .Y(_20264_));
 sg13g2_and2_1 _28826_ (.A(\u_inv.f_next[114] ),
    .B(\u_inv.f_reg[114] ),
    .X(_20265_));
 sg13g2_xor2_1 _28827_ (.B(\u_inv.f_reg[114] ),
    .A(\u_inv.f_next[114] ),
    .X(_20266_));
 sg13g2_nand2_1 _28828_ (.Y(_20267_),
    .A(\u_inv.f_next[115] ),
    .B(\u_inv.f_reg[115] ));
 sg13g2_xor2_1 _28829_ (.B(\u_inv.f_reg[115] ),
    .A(\u_inv.f_next[115] ),
    .X(_20268_));
 sg13g2_xnor2_1 _28830_ (.Y(_20269_),
    .A(\u_inv.f_next[115] ),
    .B(\u_inv.f_reg[115] ));
 sg13g2_and2_1 _28831_ (.A(_20266_),
    .B(_20268_),
    .X(_20270_));
 sg13g2_nand2_1 _28832_ (.Y(_20271_),
    .A(_20266_),
    .B(_20268_));
 sg13g2_a22oi_1 _28833_ (.Y(_20272_),
    .B1(\u_inv.f_reg[113] ),
    .B2(\u_inv.f_next[113] ),
    .A2(\u_inv.f_reg[112] ),
    .A1(\u_inv.f_next[112] ));
 sg13g2_inv_1 _28834_ (.Y(_20273_),
    .A(_20272_));
 sg13g2_o21ai_1 _28835_ (.B1(_20273_),
    .Y(_20274_),
    .A1(\u_inv.f_next[113] ),
    .A2(\u_inv.f_reg[113] ));
 sg13g2_nor2_1 _28836_ (.A(_20271_),
    .B(_20274_),
    .Y(_20275_));
 sg13g2_o21ai_1 _28837_ (.B1(_20265_),
    .Y(_20276_),
    .A1(\u_inv.f_next[115] ),
    .A2(\u_inv.f_reg[115] ));
 sg13g2_nand2_1 _28838_ (.Y(_20277_),
    .A(_20267_),
    .B(_20276_));
 sg13g2_o21ai_1 _28839_ (.B1(_20264_),
    .Y(_20278_),
    .A1(_20275_),
    .A2(_20277_));
 sg13g2_a21o_1 _28840_ (.A2(_20254_),
    .A1(_20252_),
    .B1(_20251_),
    .X(_20279_));
 sg13g2_a21oi_1 _28841_ (.A1(_18041_),
    .A2(_18219_),
    .Y(_20280_),
    .B1(_20259_));
 sg13g2_a21oi_1 _28842_ (.A1(\u_inv.f_next[117] ),
    .A2(\u_inv.f_reg[117] ),
    .Y(_20281_),
    .B1(_20280_));
 sg13g2_o21ai_1 _28843_ (.B1(_20278_),
    .Y(_20282_),
    .A1(_20257_),
    .A2(_20281_));
 sg13g2_nor2_1 _28844_ (.A(_20279_),
    .B(_20282_),
    .Y(_20283_));
 sg13g2_nor2b_1 _28845_ (.A(_20283_),
    .B_N(_20250_),
    .Y(_20284_));
 sg13g2_a22oi_1 _28846_ (.Y(_20285_),
    .B1(\u_inv.f_reg[125] ),
    .B2(\u_inv.f_next[125] ),
    .A2(\u_inv.f_reg[124] ),
    .A1(\u_inv.f_next[124] ));
 sg13g2_a21oi_1 _28847_ (.A1(_18035_),
    .A2(_18223_),
    .Y(_20286_),
    .B1(_20285_));
 sg13g2_and2_1 _28848_ (.A(_20234_),
    .B(_20286_),
    .X(_20287_));
 sg13g2_o21ai_1 _28849_ (.B1(_20228_),
    .Y(_20288_),
    .A1(_20229_),
    .A2(_20231_));
 sg13g2_a21oi_1 _28850_ (.A1(\u_inv.f_next[121] ),
    .A2(\u_inv.f_reg[121] ),
    .Y(_20289_),
    .B1(_20241_));
 sg13g2_a21oi_2 _28851_ (.B1(_20289_),
    .Y(_20290_),
    .A2(_18221_),
    .A1(_18039_));
 sg13g2_nand2_1 _28852_ (.Y(_20291_),
    .A(_20249_),
    .B(_20290_));
 sg13g2_a21oi_1 _28853_ (.A1(_18037_),
    .A2(_18222_),
    .Y(_20292_),
    .B1(_20244_));
 sg13g2_a21oi_1 _28854_ (.A1(\u_inv.f_next[123] ),
    .A2(\u_inv.f_reg[123] ),
    .Y(_20293_),
    .B1(_20292_));
 sg13g2_a21oi_1 _28855_ (.A1(_20291_),
    .A2(_20293_),
    .Y(_20294_),
    .B1(_20239_));
 sg13g2_nor4_2 _28856_ (.A(_20284_),
    .B(_20287_),
    .C(_20288_),
    .Y(_20295_),
    .D(_20294_));
 sg13g2_xnor2_1 _28857_ (.Y(_20296_),
    .A(\u_inv.f_next[47] ),
    .B(\u_inv.f_reg[47] ));
 sg13g2_nand2_1 _28858_ (.Y(_20297_),
    .A(\u_inv.f_next[46] ),
    .B(\u_inv.f_reg[46] ));
 sg13g2_xnor2_1 _28859_ (.Y(_20298_),
    .A(\u_inv.f_next[46] ),
    .B(\u_inv.f_reg[46] ));
 sg13g2_nor2_1 _28860_ (.A(_20296_),
    .B(_20298_),
    .Y(_20299_));
 sg13g2_nand2_1 _28861_ (.Y(_20300_),
    .A(\u_inv.f_next[44] ),
    .B(\u_inv.f_reg[44] ));
 sg13g2_xor2_1 _28862_ (.B(\u_inv.f_reg[44] ),
    .A(\u_inv.f_next[44] ),
    .X(_20301_));
 sg13g2_nor2_1 _28863_ (.A(\u_inv.f_next[45] ),
    .B(\u_inv.f_reg[45] ),
    .Y(_20302_));
 sg13g2_nand2_1 _28864_ (.Y(_20303_),
    .A(\u_inv.f_next[45] ),
    .B(\u_inv.f_reg[45] ));
 sg13g2_nor2b_2 _28865_ (.A(_20302_),
    .B_N(_20303_),
    .Y(_20304_));
 sg13g2_inv_1 _28866_ (.Y(_20305_),
    .A(_20304_));
 sg13g2_and2_1 _28867_ (.A(_20301_),
    .B(_20304_),
    .X(_20306_));
 sg13g2_nand2_1 _28868_ (.Y(_20307_),
    .A(_20299_),
    .B(_20306_));
 sg13g2_nor2b_1 _28869_ (.A(\u_inv.f_reg[43] ),
    .B_N(\u_inv.f_next[43] ),
    .Y(_20308_));
 sg13g2_xnor2_1 _28870_ (.Y(_20309_),
    .A(\u_inv.f_next[43] ),
    .B(\u_inv.f_reg[43] ));
 sg13g2_xor2_1 _28871_ (.B(\u_inv.f_reg[43] ),
    .A(\u_inv.f_next[43] ),
    .X(_20310_));
 sg13g2_nand2_1 _28872_ (.Y(_20311_),
    .A(\u_inv.f_next[42] ),
    .B(\u_inv.f_reg[42] ));
 sg13g2_xor2_1 _28873_ (.B(\u_inv.f_reg[42] ),
    .A(\u_inv.f_next[42] ),
    .X(_20312_));
 sg13g2_xnor2_1 _28874_ (.Y(_20313_),
    .A(\u_inv.f_next[42] ),
    .B(\u_inv.f_reg[42] ));
 sg13g2_nor2_1 _28875_ (.A(_20309_),
    .B(_20313_),
    .Y(_20314_));
 sg13g2_nand2_1 _28876_ (.Y(_20315_),
    .A(_20310_),
    .B(_20312_));
 sg13g2_nor2_1 _28877_ (.A(\u_inv.f_next[41] ),
    .B(\u_inv.f_reg[41] ),
    .Y(_20316_));
 sg13g2_a22oi_1 _28878_ (.Y(_20317_),
    .B1(\u_inv.f_reg[41] ),
    .B2(\u_inv.f_next[41] ),
    .A2(\u_inv.f_reg[40] ),
    .A1(\u_inv.f_next[40] ));
 sg13g2_nor2_1 _28879_ (.A(_20316_),
    .B(_20317_),
    .Y(_20318_));
 sg13g2_nor2_1 _28880_ (.A(\u_inv.f_next[43] ),
    .B(\u_inv.f_reg[43] ),
    .Y(_20319_));
 sg13g2_nand2_1 _28881_ (.Y(_20320_),
    .A(\u_inv.f_next[43] ),
    .B(\u_inv.f_reg[43] ));
 sg13g2_o21ai_1 _28882_ (.B1(_20320_),
    .Y(_20321_),
    .A1(_20311_),
    .A2(_20319_));
 sg13g2_inv_1 _28883_ (.Y(_20322_),
    .A(_20321_));
 sg13g2_a21oi_1 _28884_ (.A1(_20314_),
    .A2(_20318_),
    .Y(_20323_),
    .B1(_20321_));
 sg13g2_a21oi_1 _28885_ (.A1(_18078_),
    .A2(_18203_),
    .Y(_20324_),
    .B1(_20297_));
 sg13g2_o21ai_1 _28886_ (.B1(_20303_),
    .Y(_20325_),
    .A1(_20300_),
    .A2(_20302_));
 sg13g2_a221oi_1 _28887_ (.B2(_20325_),
    .C1(_20324_),
    .B1(_20299_),
    .A1(\u_inv.f_next[47] ),
    .Y(_20326_),
    .A2(\u_inv.f_reg[47] ));
 sg13g2_o21ai_1 _28888_ (.B1(_20326_),
    .Y(_20327_),
    .A1(_20307_),
    .A2(_20323_));
 sg13g2_nand2_1 _28889_ (.Y(_20328_),
    .A(\u_inv.f_next[30] ),
    .B(\u_inv.f_reg[30] ));
 sg13g2_xor2_1 _28890_ (.B(\u_inv.f_reg[30] ),
    .A(\u_inv.f_next[30] ),
    .X(_20329_));
 sg13g2_nand2_1 _28891_ (.Y(_20330_),
    .A(\u_inv.f_next[31] ),
    .B(\u_inv.f_reg[31] ));
 sg13g2_nor2_1 _28892_ (.A(\u_inv.f_next[31] ),
    .B(\u_inv.f_reg[31] ),
    .Y(_20331_));
 sg13g2_xor2_1 _28893_ (.B(\u_inv.f_reg[31] ),
    .A(\u_inv.f_next[31] ),
    .X(_20332_));
 sg13g2_inv_1 _28894_ (.Y(_20333_),
    .A(_20332_));
 sg13g2_and2_1 _28895_ (.A(_20329_),
    .B(_20332_),
    .X(_20334_));
 sg13g2_nor2_1 _28896_ (.A(\u_inv.f_next[29] ),
    .B(\u_inv.f_reg[29] ),
    .Y(_20335_));
 sg13g2_nand2_1 _28897_ (.Y(_20336_),
    .A(\u_inv.f_next[28] ),
    .B(\u_inv.f_reg[28] ));
 sg13g2_nor2_1 _28898_ (.A(_20335_),
    .B(_20336_),
    .Y(_20337_));
 sg13g2_a21oi_1 _28899_ (.A1(\u_inv.f_next[29] ),
    .A2(\u_inv.f_reg[29] ),
    .Y(_20338_),
    .B1(_20337_));
 sg13g2_and2_1 _28900_ (.A(\u_inv.f_next[27] ),
    .B(\u_inv.f_reg[27] ),
    .X(_20339_));
 sg13g2_or2_1 _28901_ (.X(_20340_),
    .B(\u_inv.f_reg[27] ),
    .A(\u_inv.f_next[27] ));
 sg13g2_and2_1 _28902_ (.A(\u_inv.f_next[26] ),
    .B(\u_inv.f_reg[26] ),
    .X(_20341_));
 sg13g2_nand2_1 _28903_ (.Y(_20342_),
    .A(\u_inv.f_next[25] ),
    .B(\u_inv.f_reg[25] ));
 sg13g2_nor2_1 _28904_ (.A(\u_inv.f_next[25] ),
    .B(\u_inv.f_reg[25] ),
    .Y(_20343_));
 sg13g2_nand2_1 _28905_ (.Y(_20344_),
    .A(\u_inv.f_next[24] ),
    .B(\u_inv.f_reg[24] ));
 sg13g2_xor2_1 _28906_ (.B(\u_inv.f_reg[22] ),
    .A(\u_inv.f_next[22] ),
    .X(_20345_));
 sg13g2_inv_1 _28907_ (.Y(_20346_),
    .A(_20345_));
 sg13g2_nor2_1 _28908_ (.A(\u_inv.f_next[23] ),
    .B(\u_inv.f_reg[23] ),
    .Y(_20347_));
 sg13g2_xor2_1 _28909_ (.B(\u_inv.f_reg[23] ),
    .A(\u_inv.f_next[23] ),
    .X(_20348_));
 sg13g2_xnor2_1 _28910_ (.Y(_20349_),
    .A(\u_inv.f_next[23] ),
    .B(\u_inv.f_reg[23] ));
 sg13g2_nor2_1 _28911_ (.A(_20346_),
    .B(_20349_),
    .Y(_20350_));
 sg13g2_nand2_1 _28912_ (.Y(_20351_),
    .A(net7300),
    .B(\u_inv.f_reg[19] ));
 sg13g2_nor2_1 _28913_ (.A(net7300),
    .B(\u_inv.f_reg[19] ),
    .Y(_20352_));
 sg13g2_and2_1 _28914_ (.A(\u_inv.f_next[18] ),
    .B(\u_inv.f_reg[18] ),
    .X(_20353_));
 sg13g2_nand2_1 _28915_ (.Y(_20354_),
    .A(\u_inv.f_next[17] ),
    .B(\u_inv.f_reg[17] ));
 sg13g2_or2_1 _28916_ (.X(_20355_),
    .B(\u_inv.f_reg[17] ),
    .A(\u_inv.f_next[17] ));
 sg13g2_nand2_1 _28917_ (.Y(_20356_),
    .A(\u_inv.f_next[16] ),
    .B(\u_inv.f_reg[16] ));
 sg13g2_nand2_1 _28918_ (.Y(_20357_),
    .A(\u_inv.f_next[15] ),
    .B(\u_inv.f_reg[15] ));
 sg13g2_or2_1 _28919_ (.X(_20358_),
    .B(\u_inv.f_reg[15] ),
    .A(\u_inv.f_next[15] ));
 sg13g2_nand2_1 _28920_ (.Y(_20359_),
    .A(\u_inv.f_next[14] ),
    .B(\u_inv.f_reg[14] ));
 sg13g2_xnor2_1 _28921_ (.Y(_20360_),
    .A(\u_inv.f_next[14] ),
    .B(\u_inv.f_reg[14] ));
 sg13g2_or2_1 _28922_ (.X(_20361_),
    .B(\u_inv.f_reg[13] ),
    .A(\u_inv.f_next[13] ));
 sg13g2_nand2_1 _28923_ (.Y(_20362_),
    .A(\u_inv.f_next[13] ),
    .B(\u_inv.f_reg[13] ));
 sg13g2_nand2_1 _28924_ (.Y(_20363_),
    .A(\u_inv.f_next[12] ),
    .B(\u_inv.f_reg[12] ));
 sg13g2_xor2_1 _28925_ (.B(\u_inv.f_reg[12] ),
    .A(\u_inv.f_next[12] ),
    .X(_20364_));
 sg13g2_inv_1 _28926_ (.Y(_20365_),
    .A(_20364_));
 sg13g2_nor2_1 _28927_ (.A(\u_inv.f_next[11] ),
    .B(\u_inv.f_reg[11] ),
    .Y(_20366_));
 sg13g2_and2_1 _28928_ (.A(\u_inv.f_next[11] ),
    .B(\u_inv.f_reg[11] ),
    .X(_20367_));
 sg13g2_nand2_1 _28929_ (.Y(_20368_),
    .A(\u_inv.f_next[10] ),
    .B(\u_inv.f_reg[10] ));
 sg13g2_xor2_1 _28930_ (.B(\u_inv.f_reg[10] ),
    .A(\u_inv.f_next[10] ),
    .X(_20369_));
 sg13g2_nand2_1 _28931_ (.Y(_20370_),
    .A(_18095_),
    .B(_18195_));
 sg13g2_and2_1 _28932_ (.A(\u_inv.f_next[8] ),
    .B(\u_inv.f_reg[8] ),
    .X(_20371_));
 sg13g2_xor2_1 _28933_ (.B(\u_inv.f_reg[8] ),
    .A(\u_inv.f_next[8] ),
    .X(_20372_));
 sg13g2_nand2_1 _28934_ (.Y(_20373_),
    .A(\u_inv.f_next[7] ),
    .B(\u_inv.f_reg[7] ));
 sg13g2_xnor2_1 _28935_ (.Y(_20374_),
    .A(\u_inv.f_next[7] ),
    .B(\u_inv.f_reg[7] ));
 sg13g2_and2_1 _28936_ (.A(\u_inv.f_next[6] ),
    .B(\u_inv.f_reg[6] ),
    .X(_20375_));
 sg13g2_xor2_1 _28937_ (.B(\u_inv.f_reg[6] ),
    .A(\u_inv.f_next[6] ),
    .X(_20376_));
 sg13g2_nand2_1 _28938_ (.Y(_20377_),
    .A(\u_inv.f_next[5] ),
    .B(\u_inv.f_reg[5] ));
 sg13g2_xnor2_1 _28939_ (.Y(_20378_),
    .A(\u_inv.f_next[5] ),
    .B(\u_inv.f_reg[5] ));
 sg13g2_nor2_1 _28940_ (.A(_18096_),
    .B(_18191_),
    .Y(_20379_));
 sg13g2_xor2_1 _28941_ (.B(\u_inv.f_reg[4] ),
    .A(\u_inv.f_next[4] ),
    .X(_20380_));
 sg13g2_nand2_1 _28942_ (.Y(_20381_),
    .A(\u_inv.f_next[3] ),
    .B(\u_inv.f_reg[3] ));
 sg13g2_xnor2_1 _28943_ (.Y(_20382_),
    .A(\u_inv.f_next[3] ),
    .B(\u_inv.f_reg[3] ));
 sg13g2_a21oi_1 _28944_ (.A1(_19825_),
    .A2(_19837_),
    .Y(_20383_),
    .B1(_19823_));
 sg13g2_o21ai_1 _28945_ (.B1(_20381_),
    .Y(_20384_),
    .A1(_20382_),
    .A2(_20383_));
 sg13g2_a21oi_1 _28946_ (.A1(_20380_),
    .A2(_20384_),
    .Y(_20385_),
    .B1(_20379_));
 sg13g2_o21ai_1 _28947_ (.B1(_20377_),
    .Y(_20386_),
    .A1(_20378_),
    .A2(_20385_));
 sg13g2_a21oi_1 _28948_ (.A1(_20376_),
    .A2(_20386_),
    .Y(_20387_),
    .B1(_20375_));
 sg13g2_o21ai_1 _28949_ (.B1(_20373_),
    .Y(_20388_),
    .A1(_20374_),
    .A2(_20387_));
 sg13g2_a21oi_1 _28950_ (.A1(_20372_),
    .A2(_20388_),
    .Y(_20389_),
    .B1(_20371_));
 sg13g2_a221oi_1 _28951_ (.B2(_20388_),
    .C1(_20371_),
    .B1(_20372_),
    .A1(\u_inv.f_next[9] ),
    .Y(_20390_),
    .A2(\u_inv.f_reg[9] ));
 sg13g2_a21oi_1 _28952_ (.A1(_18095_),
    .A2(_18195_),
    .Y(_20391_),
    .B1(_20390_));
 sg13g2_nand3b_1 _28953_ (.B(_20369_),
    .C(_20370_),
    .Y(_20392_),
    .A_N(_20390_));
 sg13g2_nand2_1 _28954_ (.Y(_20393_),
    .A(_20368_),
    .B(_20392_));
 sg13g2_a21oi_1 _28955_ (.A1(_20368_),
    .A2(_20392_),
    .Y(_20394_),
    .B1(_20366_));
 sg13g2_or2_1 _28956_ (.X(_20395_),
    .B(_20394_),
    .A(_20367_));
 sg13g2_o21ai_1 _28957_ (.B1(_20364_),
    .Y(_20396_),
    .A1(_20367_),
    .A2(_20394_));
 sg13g2_nand2_1 _28958_ (.Y(_20397_),
    .A(_20363_),
    .B(_20396_));
 sg13g2_nand3_1 _28959_ (.B(_20363_),
    .C(_20396_),
    .A(_20362_),
    .Y(_20398_));
 sg13g2_nand2_1 _28960_ (.Y(_20399_),
    .A(_20361_),
    .B(_20398_));
 sg13g2_nand3b_1 _28961_ (.B(_20361_),
    .C(_20398_),
    .Y(_20400_),
    .A_N(_20360_));
 sg13g2_nand2_1 _28962_ (.Y(_20401_),
    .A(_20359_),
    .B(_20400_));
 sg13g2_nand3_1 _28963_ (.B(_20359_),
    .C(_20400_),
    .A(_20357_),
    .Y(_20402_));
 sg13g2_nand2_1 _28964_ (.Y(_20403_),
    .A(_20358_),
    .B(_20402_));
 sg13g2_xnor2_1 _28965_ (.Y(_20404_),
    .A(\u_inv.f_next[16] ),
    .B(\u_inv.f_reg[16] ));
 sg13g2_o21ai_1 _28966_ (.B1(_20356_),
    .Y(_20405_),
    .A1(_20403_),
    .A2(_20404_));
 sg13g2_nand2b_1 _28967_ (.Y(_20406_),
    .B(_20355_),
    .A_N(_20356_));
 sg13g2_nand2_2 _28968_ (.Y(_20407_),
    .A(_20354_),
    .B(_20355_));
 sg13g2_nor2_1 _28969_ (.A(_20404_),
    .B(_20407_),
    .Y(_20408_));
 sg13g2_nand3_1 _28970_ (.B(_20402_),
    .C(_20408_),
    .A(_20358_),
    .Y(_20409_));
 sg13g2_nand3_1 _28971_ (.B(_20406_),
    .C(_20409_),
    .A(_20354_),
    .Y(_20410_));
 sg13g2_xor2_1 _28972_ (.B(\u_inv.f_reg[18] ),
    .A(\u_inv.f_next[18] ),
    .X(_20411_));
 sg13g2_a21oi_1 _28973_ (.A1(_20410_),
    .A2(_20411_),
    .Y(_20412_),
    .B1(_20353_));
 sg13g2_nor2b_1 _28974_ (.A(_20352_),
    .B_N(_20353_),
    .Y(_20413_));
 sg13g2_xor2_1 _28975_ (.B(\u_inv.f_reg[19] ),
    .A(net7300),
    .X(_20414_));
 sg13g2_xnor2_1 _28976_ (.Y(_20415_),
    .A(net7300),
    .B(\u_inv.f_reg[19] ));
 sg13g2_and2_1 _28977_ (.A(_20411_),
    .B(_20414_),
    .X(_20416_));
 sg13g2_a221oi_1 _28978_ (.B2(_20416_),
    .C1(_20413_),
    .B1(_20410_),
    .A1(net7300),
    .Y(_20417_),
    .A2(\u_inv.f_reg[19] ));
 sg13g2_o21ai_1 _28979_ (.B1(_20351_),
    .Y(_20418_),
    .A1(_20352_),
    .A2(_20412_));
 sg13g2_xor2_1 _28980_ (.B(\u_inv.f_reg[21] ),
    .A(\u_inv.f_next[21] ),
    .X(_20419_));
 sg13g2_nor2_1 _28981_ (.A(_18090_),
    .B(_18196_),
    .Y(_20420_));
 sg13g2_xor2_1 _28982_ (.B(\u_inv.f_reg[20] ),
    .A(\u_inv.f_next[20] ),
    .X(_20421_));
 sg13g2_and2_1 _28983_ (.A(_20419_),
    .B(_20421_),
    .X(_20422_));
 sg13g2_nand2_1 _28984_ (.Y(_20423_),
    .A(_20350_),
    .B(_20422_));
 sg13g2_nor3_1 _28985_ (.A(_18089_),
    .B(_18198_),
    .C(_20347_),
    .Y(_20424_));
 sg13g2_a21oi_1 _28986_ (.A1(\u_inv.f_next[21] ),
    .A2(\u_inv.f_reg[21] ),
    .Y(_20425_),
    .B1(_20420_));
 sg13g2_inv_1 _28987_ (.Y(_20426_),
    .A(_20425_));
 sg13g2_o21ai_1 _28988_ (.B1(_20426_),
    .Y(_20427_),
    .A1(\u_inv.f_next[21] ),
    .A2(\u_inv.f_reg[21] ));
 sg13g2_inv_1 _28989_ (.Y(_20428_),
    .A(_20427_));
 sg13g2_a221oi_1 _28990_ (.B2(_20428_),
    .C1(_20424_),
    .B1(_20350_),
    .A1(\u_inv.f_next[23] ),
    .Y(_20429_),
    .A2(\u_inv.f_reg[23] ));
 sg13g2_o21ai_1 _28991_ (.B1(_20429_),
    .Y(_20430_),
    .A1(_20417_),
    .A2(_20423_));
 sg13g2_xor2_1 _28992_ (.B(\u_inv.f_reg[24] ),
    .A(\u_inv.f_next[24] ),
    .X(_20431_));
 sg13g2_nand2_1 _28993_ (.Y(_20432_),
    .A(_20430_),
    .B(_20431_));
 sg13g2_o21ai_1 _28994_ (.B1(_20342_),
    .Y(_20433_),
    .A1(_20343_),
    .A2(_20344_));
 sg13g2_xnor2_1 _28995_ (.Y(_20434_),
    .A(\u_inv.f_next[25] ),
    .B(\u_inv.f_reg[25] ));
 sg13g2_inv_1 _28996_ (.Y(_20435_),
    .A(_20434_));
 sg13g2_and2_1 _28997_ (.A(_20431_),
    .B(_20435_),
    .X(_20436_));
 sg13g2_a21o_2 _28998_ (.A2(_20436_),
    .A1(_20430_),
    .B1(_20433_),
    .X(_20437_));
 sg13g2_xor2_1 _28999_ (.B(\u_inv.f_reg[26] ),
    .A(\u_inv.f_next[26] ),
    .X(_20438_));
 sg13g2_a21oi_1 _29000_ (.A1(_20437_),
    .A2(_20438_),
    .Y(_20439_),
    .B1(_20341_));
 sg13g2_nor2b_2 _29001_ (.A(_20339_),
    .B_N(_20340_),
    .Y(_20440_));
 sg13g2_and2_1 _29002_ (.A(_20438_),
    .B(_20440_),
    .X(_20441_));
 sg13g2_a221oi_1 _29003_ (.B2(_20441_),
    .C1(_20339_),
    .B1(_20437_),
    .A1(_20340_),
    .Y(_20442_),
    .A2(_20341_));
 sg13g2_xor2_1 _29004_ (.B(\u_inv.f_reg[29] ),
    .A(\u_inv.f_next[29] ),
    .X(_20443_));
 sg13g2_xnor2_1 _29005_ (.Y(_20444_),
    .A(\u_inv.f_next[29] ),
    .B(\u_inv.f_reg[29] ));
 sg13g2_nor2_1 _29006_ (.A(\u_inv.f_next[28] ),
    .B(\u_inv.f_reg[28] ),
    .Y(_20445_));
 sg13g2_xor2_1 _29007_ (.B(\u_inv.f_reg[28] ),
    .A(\u_inv.f_next[28] ),
    .X(_20446_));
 sg13g2_nand2_1 _29008_ (.Y(_20447_),
    .A(_20443_),
    .B(_20446_));
 sg13g2_o21ai_1 _29009_ (.B1(_20338_),
    .Y(_20448_),
    .A1(_20442_),
    .A2(_20447_));
 sg13g2_nand3_1 _29010_ (.B(_20443_),
    .C(_20446_),
    .A(_20334_),
    .Y(_20449_));
 sg13g2_nand2b_1 _29011_ (.Y(_20450_),
    .B(_20334_),
    .A_N(_20338_));
 sg13g2_o21ai_1 _29012_ (.B1(_20450_),
    .Y(_20451_),
    .A1(_20442_),
    .A2(_20449_));
 sg13g2_o21ai_1 _29013_ (.B1(_20330_),
    .Y(_20452_),
    .A1(_20328_),
    .A2(_20331_));
 sg13g2_nor2_1 _29014_ (.A(_20451_),
    .B(_20452_),
    .Y(_20453_));
 sg13g2_nand2_1 _29015_ (.Y(_20454_),
    .A(\u_inv.f_next[34] ),
    .B(\u_inv.f_reg[34] ));
 sg13g2_xor2_1 _29016_ (.B(\u_inv.f_reg[34] ),
    .A(\u_inv.f_next[34] ),
    .X(_20455_));
 sg13g2_nand2_1 _29017_ (.Y(_20456_),
    .A(\u_inv.f_next[35] ),
    .B(\u_inv.f_reg[35] ));
 sg13g2_nor2_1 _29018_ (.A(\u_inv.f_next[35] ),
    .B(\u_inv.f_reg[35] ),
    .Y(_20457_));
 sg13g2_xor2_1 _29019_ (.B(\u_inv.f_reg[35] ),
    .A(\u_inv.f_next[35] ),
    .X(_20458_));
 sg13g2_nand2_1 _29020_ (.Y(_20459_),
    .A(_20455_),
    .B(_20458_));
 sg13g2_xor2_1 _29021_ (.B(\u_inv.f_reg[33] ),
    .A(\u_inv.f_next[33] ),
    .X(_20460_));
 sg13g2_xnor2_1 _29022_ (.Y(_20461_),
    .A(\u_inv.f_next[32] ),
    .B(\u_inv.f_reg[32] ));
 sg13g2_inv_1 _29023_ (.Y(_20462_),
    .A(_20461_));
 sg13g2_nand2_1 _29024_ (.Y(_20463_),
    .A(_20460_),
    .B(_20462_));
 sg13g2_nor2_1 _29025_ (.A(_20459_),
    .B(_20463_),
    .Y(_20464_));
 sg13g2_o21ai_1 _29026_ (.B1(_20464_),
    .Y(_20465_),
    .A1(_20451_),
    .A2(_20452_));
 sg13g2_o21ai_1 _29027_ (.B1(_20456_),
    .Y(_20466_),
    .A1(_20454_),
    .A2(_20457_));
 sg13g2_a22oi_1 _29028_ (.Y(_20467_),
    .B1(\u_inv.f_reg[33] ),
    .B2(\u_inv.f_next[33] ),
    .A2(\u_inv.f_reg[32] ),
    .A1(\u_inv.f_next[32] ));
 sg13g2_inv_1 _29029_ (.Y(_20468_),
    .A(_20467_));
 sg13g2_o21ai_1 _29030_ (.B1(_20468_),
    .Y(_20469_),
    .A1(\u_inv.f_next[33] ),
    .A2(\u_inv.f_reg[33] ));
 sg13g2_nor2_1 _29031_ (.A(_20459_),
    .B(_20469_),
    .Y(_20470_));
 sg13g2_nor2_1 _29032_ (.A(_20466_),
    .B(_20470_),
    .Y(_20471_));
 sg13g2_nand2_1 _29033_ (.Y(_20472_),
    .A(_20465_),
    .B(_20471_));
 sg13g2_xnor2_1 _29034_ (.Y(_20473_),
    .A(\u_inv.f_next[39] ),
    .B(\u_inv.f_reg[39] ));
 sg13g2_nand2_1 _29035_ (.Y(_20474_),
    .A(\u_inv.f_next[38] ),
    .B(\u_inv.f_reg[38] ));
 sg13g2_xnor2_1 _29036_ (.Y(_20475_),
    .A(\u_inv.f_next[38] ),
    .B(\u_inv.f_reg[38] ));
 sg13g2_nor2_1 _29037_ (.A(_20473_),
    .B(_20475_),
    .Y(_20476_));
 sg13g2_nand2_1 _29038_ (.Y(_20477_),
    .A(\u_inv.f_next[36] ),
    .B(\u_inv.f_reg[36] ));
 sg13g2_xnor2_1 _29039_ (.Y(_20478_),
    .A(\u_inv.f_next[36] ),
    .B(\u_inv.f_reg[36] ));
 sg13g2_nor2_1 _29040_ (.A(\u_inv.f_next[37] ),
    .B(\u_inv.f_reg[37] ),
    .Y(_20479_));
 sg13g2_nand2_1 _29041_ (.Y(_20480_),
    .A(\u_inv.f_next[37] ),
    .B(\u_inv.f_reg[37] ));
 sg13g2_nor2b_2 _29042_ (.A(_20479_),
    .B_N(_20480_),
    .Y(_20481_));
 sg13g2_nand2b_1 _29043_ (.Y(_20482_),
    .B(_20480_),
    .A_N(_20479_));
 sg13g2_nor2_1 _29044_ (.A(_20478_),
    .B(_20482_),
    .Y(_20483_));
 sg13g2_nand2_1 _29045_ (.Y(_20484_),
    .A(_20476_),
    .B(_20483_));
 sg13g2_a21o_2 _29046_ (.A2(_20471_),
    .A1(_20465_),
    .B1(_20484_),
    .X(_20485_));
 sg13g2_a21oi_1 _29047_ (.A1(_18081_),
    .A2(_18202_),
    .Y(_20486_),
    .B1(_20474_));
 sg13g2_o21ai_1 _29048_ (.B1(_20480_),
    .Y(_20487_),
    .A1(_20477_),
    .A2(_20479_));
 sg13g2_a221oi_1 _29049_ (.B2(_20487_),
    .C1(_20486_),
    .B1(_20476_),
    .A1(\u_inv.f_next[39] ),
    .Y(_20488_),
    .A2(\u_inv.f_reg[39] ));
 sg13g2_nand2_1 _29050_ (.Y(_20489_),
    .A(_20485_),
    .B(_20488_));
 sg13g2_xnor2_1 _29051_ (.Y(_20490_),
    .A(\u_inv.f_next[40] ),
    .B(\u_inv.f_reg[40] ));
 sg13g2_xnor2_1 _29052_ (.Y(_20491_),
    .A(\u_inv.f_next[41] ),
    .B(\u_inv.f_reg[41] ));
 sg13g2_nor2_1 _29053_ (.A(_20490_),
    .B(_20491_),
    .Y(_20492_));
 sg13g2_nor4_1 _29054_ (.A(_20307_),
    .B(_20315_),
    .C(_20490_),
    .D(_20491_),
    .Y(_20493_));
 sg13g2_inv_1 _29055_ (.Y(_20494_),
    .A(_20493_));
 sg13g2_a21oi_2 _29056_ (.B1(_20494_),
    .Y(_20495_),
    .A2(_20488_),
    .A1(_20485_));
 sg13g2_nor2_1 _29057_ (.A(_20327_),
    .B(_20495_),
    .Y(_20496_));
 sg13g2_nor2_1 _29058_ (.A(\u_inv.f_next[49] ),
    .B(\u_inv.f_reg[49] ),
    .Y(_20497_));
 sg13g2_nand2_1 _29059_ (.Y(_20498_),
    .A(\u_inv.f_next[49] ),
    .B(\u_inv.f_reg[49] ));
 sg13g2_nor2b_2 _29060_ (.A(_20497_),
    .B_N(_20498_),
    .Y(_20499_));
 sg13g2_nand2b_1 _29061_ (.Y(_20500_),
    .B(_20498_),
    .A_N(_20497_));
 sg13g2_nand2_1 _29062_ (.Y(_20501_),
    .A(\u_inv.f_next[48] ),
    .B(\u_inv.f_reg[48] ));
 sg13g2_xnor2_1 _29063_ (.Y(_20502_),
    .A(\u_inv.f_next[48] ),
    .B(\u_inv.f_reg[48] ));
 sg13g2_nor3_1 _29064_ (.A(_20496_),
    .B(_20500_),
    .C(_20502_),
    .Y(_20503_));
 sg13g2_nor2_1 _29065_ (.A(\u_inv.f_next[51] ),
    .B(\u_inv.f_reg[51] ),
    .Y(_20504_));
 sg13g2_nand2_1 _29066_ (.Y(_20505_),
    .A(\u_inv.f_next[50] ),
    .B(\u_inv.f_reg[50] ));
 sg13g2_nor2_1 _29067_ (.A(_20504_),
    .B(_20505_),
    .Y(_20506_));
 sg13g2_o21ai_1 _29068_ (.B1(_20498_),
    .Y(_20507_),
    .A1(_20497_),
    .A2(_20501_));
 sg13g2_xnor2_1 _29069_ (.Y(_20508_),
    .A(\u_inv.f_next[50] ),
    .B(\u_inv.f_reg[50] ));
 sg13g2_xnor2_1 _29070_ (.Y(_20509_),
    .A(\u_inv.f_next[51] ),
    .B(\u_inv.f_reg[51] ));
 sg13g2_nor2_1 _29071_ (.A(_20508_),
    .B(_20509_),
    .Y(_20510_));
 sg13g2_or4_1 _29072_ (.A(_20500_),
    .B(_20502_),
    .C(_20508_),
    .D(_20509_),
    .X(_20511_));
 sg13g2_inv_1 _29073_ (.Y(_20512_),
    .A(_20511_));
 sg13g2_o21ai_1 _29074_ (.B1(_20512_),
    .Y(_20513_),
    .A1(_20327_),
    .A2(_20495_));
 sg13g2_a221oi_1 _29075_ (.B2(_20510_),
    .C1(_20506_),
    .B1(_20507_),
    .A1(\u_inv.f_next[51] ),
    .Y(_20514_),
    .A2(\u_inv.f_reg[51] ));
 sg13g2_nand2_1 _29076_ (.Y(_20515_),
    .A(_20513_),
    .B(_20514_));
 sg13g2_nand2_1 _29077_ (.Y(_20516_),
    .A(\u_inv.f_next[54] ),
    .B(\u_inv.f_reg[54] ));
 sg13g2_nor2_1 _29078_ (.A(\u_inv.f_next[54] ),
    .B(\u_inv.f_reg[54] ),
    .Y(_20517_));
 sg13g2_xor2_1 _29079_ (.B(\u_inv.f_reg[54] ),
    .A(\u_inv.f_next[54] ),
    .X(_20518_));
 sg13g2_xor2_1 _29080_ (.B(\u_inv.f_reg[55] ),
    .A(\u_inv.f_next[55] ),
    .X(_20519_));
 sg13g2_and2_1 _29081_ (.A(_20518_),
    .B(_20519_),
    .X(_20520_));
 sg13g2_nor2_1 _29082_ (.A(\u_inv.f_next[53] ),
    .B(\u_inv.f_reg[53] ),
    .Y(_20521_));
 sg13g2_xor2_1 _29083_ (.B(\u_inv.f_reg[53] ),
    .A(\u_inv.f_next[53] ),
    .X(_20522_));
 sg13g2_xnor2_1 _29084_ (.Y(_20523_),
    .A(\u_inv.f_next[53] ),
    .B(\u_inv.f_reg[53] ));
 sg13g2_and2_1 _29085_ (.A(\u_inv.f_next[52] ),
    .B(\u_inv.f_reg[52] ),
    .X(_20524_));
 sg13g2_xor2_1 _29086_ (.B(\u_inv.f_reg[52] ),
    .A(\u_inv.f_next[52] ),
    .X(_20525_));
 sg13g2_xnor2_1 _29087_ (.Y(_20526_),
    .A(\u_inv.f_next[52] ),
    .B(\u_inv.f_reg[52] ));
 sg13g2_nor2_1 _29088_ (.A(_20523_),
    .B(_20526_),
    .Y(_20527_));
 sg13g2_nand2_1 _29089_ (.Y(_20528_),
    .A(_20520_),
    .B(_20527_));
 sg13g2_a21oi_1 _29090_ (.A1(_20513_),
    .A2(_20514_),
    .Y(_20529_),
    .B1(_20528_));
 sg13g2_a21oi_1 _29091_ (.A1(_18074_),
    .A2(_18205_),
    .Y(_20530_),
    .B1(_20516_));
 sg13g2_a21oi_1 _29092_ (.A1(\u_inv.f_next[53] ),
    .A2(\u_inv.f_reg[53] ),
    .Y(_20531_),
    .B1(_20524_));
 sg13g2_nor2_1 _29093_ (.A(_20521_),
    .B(_20531_),
    .Y(_20532_));
 sg13g2_a221oi_1 _29094_ (.B2(_20532_),
    .C1(_20530_),
    .B1(_20520_),
    .A1(\u_inv.f_next[55] ),
    .Y(_20533_),
    .A2(\u_inv.f_reg[55] ));
 sg13g2_inv_1 _29095_ (.Y(_20534_),
    .A(_20533_));
 sg13g2_nand2b_2 _29096_ (.Y(_20535_),
    .B(_20533_),
    .A_N(_20529_));
 sg13g2_xor2_1 _29097_ (.B(\u_inv.f_reg[61] ),
    .A(\u_inv.f_next[61] ),
    .X(_20536_));
 sg13g2_and2_1 _29098_ (.A(\u_inv.f_next[60] ),
    .B(\u_inv.f_reg[60] ),
    .X(_20537_));
 sg13g2_xor2_1 _29099_ (.B(\u_inv.f_reg[60] ),
    .A(\u_inv.f_next[60] ),
    .X(_20538_));
 sg13g2_inv_1 _29100_ (.Y(_20539_),
    .A(_20538_));
 sg13g2_nand2_1 _29101_ (.Y(_20540_),
    .A(\u_inv.f_next[63] ),
    .B(\u_inv.f_reg[63] ));
 sg13g2_nor2_1 _29102_ (.A(\u_inv.f_next[63] ),
    .B(\u_inv.f_reg[63] ),
    .Y(_20541_));
 sg13g2_xor2_1 _29103_ (.B(\u_inv.f_reg[63] ),
    .A(\u_inv.f_next[63] ),
    .X(_20542_));
 sg13g2_nand2_1 _29104_ (.Y(_20543_),
    .A(\u_inv.f_next[62] ),
    .B(\u_inv.f_reg[62] ));
 sg13g2_xor2_1 _29105_ (.B(\u_inv.f_reg[62] ),
    .A(\u_inv.f_next[62] ),
    .X(_20544_));
 sg13g2_nand2_1 _29106_ (.Y(_20545_),
    .A(_20542_),
    .B(_20544_));
 sg13g2_nand4_1 _29107_ (.B(_20538_),
    .C(_20542_),
    .A(_20536_),
    .Y(_20546_),
    .D(_20544_));
 sg13g2_nand2_1 _29108_ (.Y(_20547_),
    .A(\u_inv.f_next[59] ),
    .B(_18206_));
 sg13g2_xor2_1 _29109_ (.B(\u_inv.f_reg[59] ),
    .A(\u_inv.f_next[59] ),
    .X(_20548_));
 sg13g2_nor2b_1 _29110_ (.A(\u_inv.f_reg[58] ),
    .B_N(\u_inv.f_next[58] ),
    .Y(_20549_));
 sg13g2_xnor2_1 _29111_ (.Y(_20550_),
    .A(\u_inv.f_next[58] ),
    .B(\u_inv.f_reg[58] ));
 sg13g2_xor2_1 _29112_ (.B(\u_inv.f_reg[58] ),
    .A(\u_inv.f_next[58] ),
    .X(_20551_));
 sg13g2_nand2_1 _29113_ (.Y(_20552_),
    .A(_20548_),
    .B(_20551_));
 sg13g2_nand2_1 _29114_ (.Y(_20553_),
    .A(\u_inv.f_next[57] ),
    .B(\u_inv.f_reg[57] ));
 sg13g2_nor2_1 _29115_ (.A(\u_inv.f_next[57] ),
    .B(\u_inv.f_reg[57] ),
    .Y(_20554_));
 sg13g2_xor2_1 _29116_ (.B(\u_inv.f_reg[57] ),
    .A(\u_inv.f_next[57] ),
    .X(_20555_));
 sg13g2_xnor2_1 _29117_ (.Y(_20556_),
    .A(\u_inv.f_next[57] ),
    .B(\u_inv.f_reg[57] ));
 sg13g2_nand2_1 _29118_ (.Y(_20557_),
    .A(\u_inv.f_next[56] ),
    .B(\u_inv.f_reg[56] ));
 sg13g2_xor2_1 _29119_ (.B(\u_inv.f_reg[56] ),
    .A(\u_inv.f_next[56] ),
    .X(_20558_));
 sg13g2_xnor2_1 _29120_ (.Y(_20559_),
    .A(\u_inv.f_next[56] ),
    .B(\u_inv.f_reg[56] ));
 sg13g2_nor2_1 _29121_ (.A(_20556_),
    .B(_20559_),
    .Y(_20560_));
 sg13g2_nor4_1 _29122_ (.A(_20546_),
    .B(_20552_),
    .C(_20556_),
    .D(_20559_),
    .Y(_20561_));
 sg13g2_o21ai_1 _29123_ (.B1(_20561_),
    .Y(_20562_),
    .A1(_20529_),
    .A2(_20534_));
 sg13g2_o21ai_1 _29124_ (.B1(_20553_),
    .Y(_20563_),
    .A1(_20554_),
    .A2(_20557_));
 sg13g2_nand2b_1 _29125_ (.Y(_20564_),
    .B(_20563_),
    .A_N(_20552_));
 sg13g2_nand2_1 _29126_ (.Y(_20565_),
    .A(\u_inv.f_next[58] ),
    .B(\u_inv.f_reg[58] ));
 sg13g2_o21ai_1 _29127_ (.B1(_20565_),
    .Y(_20566_),
    .A1(_18072_),
    .A2(_18206_));
 sg13g2_o21ai_1 _29128_ (.B1(_20566_),
    .Y(_20567_),
    .A1(\u_inv.f_next[59] ),
    .A2(\u_inv.f_reg[59] ));
 sg13g2_a21oi_1 _29129_ (.A1(_20564_),
    .A2(_20567_),
    .Y(_20568_),
    .B1(_20546_));
 sg13g2_o21ai_1 _29130_ (.B1(_20540_),
    .Y(_20569_),
    .A1(_20541_),
    .A2(_20543_));
 sg13g2_a21oi_1 _29131_ (.A1(\u_inv.f_next[61] ),
    .A2(\u_inv.f_reg[61] ),
    .Y(_20570_),
    .B1(_20537_));
 sg13g2_inv_1 _29132_ (.Y(_20571_),
    .A(_20570_));
 sg13g2_o21ai_1 _29133_ (.B1(_20571_),
    .Y(_20572_),
    .A1(\u_inv.f_next[61] ),
    .A2(\u_inv.f_reg[61] ));
 sg13g2_nor2_1 _29134_ (.A(_20568_),
    .B(_20569_),
    .Y(_20573_));
 sg13g2_o21ai_1 _29135_ (.B1(_20573_),
    .Y(_20574_),
    .A1(_20545_),
    .A2(_20572_));
 sg13g2_inv_1 _29136_ (.Y(_20575_),
    .A(_20574_));
 sg13g2_and2_1 _29137_ (.A(_20562_),
    .B(_20575_),
    .X(_20576_));
 sg13g2_nand2_1 _29138_ (.Y(_20577_),
    .A(\u_inv.f_next[66] ),
    .B(\u_inv.f_reg[66] ));
 sg13g2_xor2_1 _29139_ (.B(\u_inv.f_reg[66] ),
    .A(\u_inv.f_next[66] ),
    .X(_20578_));
 sg13g2_xnor2_1 _29140_ (.Y(_20579_),
    .A(\u_inv.f_next[66] ),
    .B(\u_inv.f_reg[66] ));
 sg13g2_nand2_1 _29141_ (.Y(_20580_),
    .A(\u_inv.f_next[67] ),
    .B(\u_inv.f_reg[67] ));
 sg13g2_nor2_1 _29142_ (.A(\u_inv.f_next[67] ),
    .B(\u_inv.f_reg[67] ),
    .Y(_20581_));
 sg13g2_xnor2_1 _29143_ (.Y(_20582_),
    .A(\u_inv.f_next[67] ),
    .B(\u_inv.f_reg[67] ));
 sg13g2_nand2_1 _29144_ (.Y(_20583_),
    .A(\u_inv.f_next[65] ),
    .B(\u_inv.f_reg[65] ));
 sg13g2_xnor2_1 _29145_ (.Y(_20584_),
    .A(\u_inv.f_next[65] ),
    .B(\u_inv.f_reg[65] ));
 sg13g2_nand2_1 _29146_ (.Y(_20585_),
    .A(\u_inv.f_next[64] ),
    .B(\u_inv.f_reg[64] ));
 sg13g2_xnor2_1 _29147_ (.Y(_20586_),
    .A(\u_inv.f_next[64] ),
    .B(\u_inv.f_reg[64] ));
 sg13g2_or4_1 _29148_ (.A(_20579_),
    .B(_20582_),
    .C(_20584_),
    .D(_20586_),
    .X(_20587_));
 sg13g2_a21oi_1 _29149_ (.A1(_20562_),
    .A2(_20575_),
    .Y(_20588_),
    .B1(_20587_));
 sg13g2_o21ai_1 _29150_ (.B1(_20580_),
    .Y(_20589_),
    .A1(_20577_),
    .A2(_20581_));
 sg13g2_nand2_1 _29151_ (.Y(_20590_),
    .A(_20583_),
    .B(_20585_));
 sg13g2_o21ai_1 _29152_ (.B1(_20590_),
    .Y(_20591_),
    .A1(\u_inv.f_next[65] ),
    .A2(\u_inv.f_reg[65] ));
 sg13g2_nor3_1 _29153_ (.A(_20579_),
    .B(_20582_),
    .C(_20591_),
    .Y(_20592_));
 sg13g2_nor2_1 _29154_ (.A(_20589_),
    .B(_20592_),
    .Y(_20593_));
 sg13g2_inv_1 _29155_ (.Y(_20594_),
    .A(_20593_));
 sg13g2_nand2b_2 _29156_ (.Y(_20595_),
    .B(_20593_),
    .A_N(_20588_));
 sg13g2_nand2_1 _29157_ (.Y(_20596_),
    .A(\u_inv.f_next[70] ),
    .B(\u_inv.f_reg[70] ));
 sg13g2_xnor2_1 _29158_ (.Y(_20597_),
    .A(\u_inv.f_next[70] ),
    .B(\u_inv.f_reg[70] ));
 sg13g2_nor2_1 _29159_ (.A(\u_inv.f_next[71] ),
    .B(\u_inv.f_reg[71] ),
    .Y(_20598_));
 sg13g2_xor2_1 _29160_ (.B(\u_inv.f_reg[71] ),
    .A(\u_inv.f_next[71] ),
    .X(_20599_));
 sg13g2_xnor2_1 _29161_ (.Y(_20600_),
    .A(\u_inv.f_next[71] ),
    .B(\u_inv.f_reg[71] ));
 sg13g2_nor2_1 _29162_ (.A(_20597_),
    .B(_20600_),
    .Y(_20601_));
 sg13g2_xor2_1 _29163_ (.B(\u_inv.f_reg[69] ),
    .A(\u_inv.f_next[69] ),
    .X(_20602_));
 sg13g2_xnor2_1 _29164_ (.Y(_20603_),
    .A(\u_inv.f_next[69] ),
    .B(\u_inv.f_reg[69] ));
 sg13g2_and2_1 _29165_ (.A(\u_inv.f_next[68] ),
    .B(\u_inv.f_reg[68] ),
    .X(_20604_));
 sg13g2_xor2_1 _29166_ (.B(\u_inv.f_reg[68] ),
    .A(\u_inv.f_next[68] ),
    .X(_20605_));
 sg13g2_and2_1 _29167_ (.A(_20602_),
    .B(_20605_),
    .X(_20606_));
 sg13g2_and2_1 _29168_ (.A(_20601_),
    .B(_20606_),
    .X(_20607_));
 sg13g2_o21ai_1 _29169_ (.B1(_20607_),
    .Y(_20608_),
    .A1(_20588_),
    .A2(_20594_));
 sg13g2_nor2_1 _29170_ (.A(_20596_),
    .B(_20598_),
    .Y(_20609_));
 sg13g2_a21oi_1 _29171_ (.A1(\u_inv.f_next[69] ),
    .A2(\u_inv.f_reg[69] ),
    .Y(_20610_),
    .B1(_20604_));
 sg13g2_a21oi_1 _29172_ (.A1(_18067_),
    .A2(_18208_),
    .Y(_20611_),
    .B1(_20610_));
 sg13g2_a221oi_1 _29173_ (.B2(_20611_),
    .C1(_20609_),
    .B1(_20601_),
    .A1(\u_inv.f_next[71] ),
    .Y(_20612_),
    .A2(\u_inv.f_reg[71] ));
 sg13g2_nand2_1 _29174_ (.Y(_20613_),
    .A(_20608_),
    .B(_20612_));
 sg13g2_nand2_1 _29175_ (.Y(_20614_),
    .A(\u_inv.f_next[79] ),
    .B(\u_inv.f_reg[79] ));
 sg13g2_nor2_1 _29176_ (.A(\u_inv.f_next[79] ),
    .B(\u_inv.f_reg[79] ),
    .Y(_20615_));
 sg13g2_xor2_1 _29177_ (.B(\u_inv.f_reg[79] ),
    .A(\u_inv.f_next[79] ),
    .X(_20616_));
 sg13g2_inv_1 _29178_ (.Y(_20617_),
    .A(_20616_));
 sg13g2_nand2_1 _29179_ (.Y(_20618_),
    .A(\u_inv.f_next[78] ),
    .B(\u_inv.f_reg[78] ));
 sg13g2_nor2_1 _29180_ (.A(\u_inv.f_next[78] ),
    .B(\u_inv.f_reg[78] ),
    .Y(_20619_));
 sg13g2_xor2_1 _29181_ (.B(\u_inv.f_reg[78] ),
    .A(\u_inv.f_next[78] ),
    .X(_20620_));
 sg13g2_and2_1 _29182_ (.A(\u_inv.f_next[76] ),
    .B(\u_inv.f_reg[76] ),
    .X(_20621_));
 sg13g2_xor2_1 _29183_ (.B(\u_inv.f_reg[76] ),
    .A(\u_inv.f_next[76] ),
    .X(_20622_));
 sg13g2_xnor2_1 _29184_ (.Y(_20623_),
    .A(\u_inv.f_next[76] ),
    .B(\u_inv.f_reg[76] ));
 sg13g2_xor2_1 _29185_ (.B(\u_inv.f_reg[77] ),
    .A(\u_inv.f_next[77] ),
    .X(_20624_));
 sg13g2_and2_1 _29186_ (.A(_20622_),
    .B(_20624_),
    .X(_20625_));
 sg13g2_nand3_1 _29187_ (.B(_20620_),
    .C(_20625_),
    .A(_20616_),
    .Y(_20626_));
 sg13g2_nand2_1 _29188_ (.Y(_20627_),
    .A(\u_inv.f_next[75] ),
    .B(\u_inv.f_reg[75] ));
 sg13g2_xor2_1 _29189_ (.B(\u_inv.f_reg[75] ),
    .A(\u_inv.f_next[75] ),
    .X(_20628_));
 sg13g2_xnor2_1 _29190_ (.Y(_20629_),
    .A(\u_inv.f_next[75] ),
    .B(\u_inv.f_reg[75] ));
 sg13g2_nand2_1 _29191_ (.Y(_20630_),
    .A(\u_inv.f_next[74] ),
    .B(\u_inv.f_reg[74] ));
 sg13g2_xor2_1 _29192_ (.B(\u_inv.f_reg[74] ),
    .A(\u_inv.f_next[74] ),
    .X(_20631_));
 sg13g2_xnor2_1 _29193_ (.Y(_20632_),
    .A(\u_inv.f_next[74] ),
    .B(\u_inv.f_reg[74] ));
 sg13g2_nand2_1 _29194_ (.Y(_20633_),
    .A(_20628_),
    .B(_20631_));
 sg13g2_xor2_1 _29195_ (.B(\u_inv.f_reg[73] ),
    .A(\u_inv.f_next[73] ),
    .X(_20634_));
 sg13g2_and2_1 _29196_ (.A(\u_inv.f_next[72] ),
    .B(\u_inv.f_reg[72] ),
    .X(_20635_));
 sg13g2_xor2_1 _29197_ (.B(\u_inv.f_reg[72] ),
    .A(\u_inv.f_next[72] ),
    .X(_20636_));
 sg13g2_nand2_1 _29198_ (.Y(_20637_),
    .A(_20634_),
    .B(_20636_));
 sg13g2_nor3_1 _29199_ (.A(_20626_),
    .B(_20633_),
    .C(_20637_),
    .Y(_20638_));
 sg13g2_inv_1 _29200_ (.Y(_20639_),
    .A(_20638_));
 sg13g2_a21oi_1 _29201_ (.A1(_20608_),
    .A2(_20612_),
    .Y(_20640_),
    .B1(_20639_));
 sg13g2_a21oi_1 _29202_ (.A1(\u_inv.f_next[73] ),
    .A2(\u_inv.f_reg[73] ),
    .Y(_20641_),
    .B1(_20635_));
 sg13g2_a21oi_1 _29203_ (.A1(_18065_),
    .A2(_18209_),
    .Y(_20642_),
    .B1(_20641_));
 sg13g2_nor2b_1 _29204_ (.A(_20633_),
    .B_N(_20642_),
    .Y(_20643_));
 sg13g2_nand2_1 _29205_ (.Y(_20644_),
    .A(_20627_),
    .B(_20630_));
 sg13g2_o21ai_1 _29206_ (.B1(_20644_),
    .Y(_20645_),
    .A1(\u_inv.f_next[75] ),
    .A2(\u_inv.f_reg[75] ));
 sg13g2_nor2b_1 _29207_ (.A(_20643_),
    .B_N(_20645_),
    .Y(_20646_));
 sg13g2_o21ai_1 _29208_ (.B1(_20614_),
    .Y(_20647_),
    .A1(_20615_),
    .A2(_20618_));
 sg13g2_a21oi_1 _29209_ (.A1(\u_inv.f_next[77] ),
    .A2(\u_inv.f_reg[77] ),
    .Y(_20648_),
    .B1(_20621_));
 sg13g2_a21oi_1 _29210_ (.A1(_18064_),
    .A2(_18210_),
    .Y(_20649_),
    .B1(_20648_));
 sg13g2_nand3_1 _29211_ (.B(_20620_),
    .C(_20649_),
    .A(_20616_),
    .Y(_20650_));
 sg13g2_o21ai_1 _29212_ (.B1(_20650_),
    .Y(_20651_),
    .A1(_20626_),
    .A2(_20646_));
 sg13g2_nor2_1 _29213_ (.A(_20647_),
    .B(_20651_),
    .Y(_20652_));
 sg13g2_inv_1 _29214_ (.Y(_20653_),
    .A(_20652_));
 sg13g2_nor2_1 _29215_ (.A(_20640_),
    .B(_20653_),
    .Y(_20654_));
 sg13g2_xor2_1 _29216_ (.B(\u_inv.f_reg[81] ),
    .A(\u_inv.f_next[81] ),
    .X(_20655_));
 sg13g2_xnor2_1 _29217_ (.Y(_20656_),
    .A(\u_inv.f_next[81] ),
    .B(\u_inv.f_reg[81] ));
 sg13g2_nand2_1 _29218_ (.Y(_20657_),
    .A(\u_inv.f_next[80] ),
    .B(\u_inv.f_reg[80] ));
 sg13g2_xnor2_1 _29219_ (.Y(_20658_),
    .A(\u_inv.f_next[80] ),
    .B(\u_inv.f_reg[80] ));
 sg13g2_nor2_1 _29220_ (.A(_20656_),
    .B(_20658_),
    .Y(_20659_));
 sg13g2_o21ai_1 _29221_ (.B1(_20659_),
    .Y(_20660_),
    .A1(_20640_),
    .A2(_20653_));
 sg13g2_a21oi_1 _29222_ (.A1(_18060_),
    .A2(_18211_),
    .Y(_20661_),
    .B1(_20657_));
 sg13g2_a21oi_1 _29223_ (.A1(\u_inv.f_next[81] ),
    .A2(\u_inv.f_reg[81] ),
    .Y(_20662_),
    .B1(_20661_));
 sg13g2_and2_1 _29224_ (.A(_20660_),
    .B(_20662_),
    .X(_20663_));
 sg13g2_nor2_1 _29225_ (.A(\u_inv.f_next[83] ),
    .B(\u_inv.f_reg[83] ),
    .Y(_20664_));
 sg13g2_nand2_1 _29226_ (.Y(_20665_),
    .A(\u_inv.f_next[83] ),
    .B(\u_inv.f_reg[83] ));
 sg13g2_nor2b_2 _29227_ (.A(_20664_),
    .B_N(_20665_),
    .Y(_20666_));
 sg13g2_nand2_2 _29228_ (.Y(_20667_),
    .A(\u_inv.f_next[82] ),
    .B(\u_inv.f_reg[82] ));
 sg13g2_or2_1 _29229_ (.X(_20668_),
    .B(\u_inv.f_reg[82] ),
    .A(\u_inv.f_next[82] ));
 sg13g2_nand2_2 _29230_ (.Y(_20669_),
    .A(_20667_),
    .B(_20668_));
 sg13g2_nand3_1 _29231_ (.B(_20667_),
    .C(_20668_),
    .A(_20666_),
    .Y(_20670_));
 sg13g2_a21oi_1 _29232_ (.A1(_20660_),
    .A2(_20662_),
    .Y(_20671_),
    .B1(_20670_));
 sg13g2_o21ai_1 _29233_ (.B1(_20665_),
    .Y(_20672_),
    .A1(_20664_),
    .A2(_20667_));
 sg13g2_nor2_2 _29234_ (.A(_20671_),
    .B(_20672_),
    .Y(_20673_));
 sg13g2_and2_1 _29235_ (.A(\u_inv.f_next[86] ),
    .B(\u_inv.f_reg[86] ),
    .X(_20674_));
 sg13g2_xor2_1 _29236_ (.B(\u_inv.f_reg[86] ),
    .A(\u_inv.f_next[86] ),
    .X(_20675_));
 sg13g2_xnor2_1 _29237_ (.Y(_20676_),
    .A(\u_inv.f_next[86] ),
    .B(\u_inv.f_reg[86] ));
 sg13g2_and2_1 _29238_ (.A(\u_inv.f_next[87] ),
    .B(\u_inv.f_reg[87] ),
    .X(_20677_));
 sg13g2_or2_1 _29239_ (.X(_20678_),
    .B(\u_inv.f_reg[87] ),
    .A(\u_inv.f_next[87] ));
 sg13g2_nor2b_1 _29240_ (.A(_20677_),
    .B_N(_20678_),
    .Y(_20679_));
 sg13g2_nand2b_2 _29241_ (.Y(_20680_),
    .B(_20678_),
    .A_N(_20677_));
 sg13g2_nand2_1 _29242_ (.Y(_20681_),
    .A(\u_inv.f_next[85] ),
    .B(\u_inv.f_reg[85] ));
 sg13g2_xor2_1 _29243_ (.B(\u_inv.f_reg[85] ),
    .A(\u_inv.f_next[85] ),
    .X(_20682_));
 sg13g2_nand2_1 _29244_ (.Y(_20683_),
    .A(\u_inv.f_next[84] ),
    .B(\u_inv.f_reg[84] ));
 sg13g2_xor2_1 _29245_ (.B(\u_inv.f_reg[84] ),
    .A(\u_inv.f_next[84] ),
    .X(_20684_));
 sg13g2_xnor2_1 _29246_ (.Y(_20685_),
    .A(\u_inv.f_next[84] ),
    .B(\u_inv.f_reg[84] ));
 sg13g2_nand2_1 _29247_ (.Y(_20686_),
    .A(_20682_),
    .B(_20684_));
 sg13g2_nor3_1 _29248_ (.A(_20676_),
    .B(_20680_),
    .C(_20686_),
    .Y(_20687_));
 sg13g2_o21ai_1 _29249_ (.B1(_20687_),
    .Y(_20688_),
    .A1(_20671_),
    .A2(_20672_));
 sg13g2_a21oi_1 _29250_ (.A1(_20674_),
    .A2(_20678_),
    .Y(_20689_),
    .B1(_20677_));
 sg13g2_nand2_1 _29251_ (.Y(_20690_),
    .A(_20681_),
    .B(_20683_));
 sg13g2_o21ai_1 _29252_ (.B1(_20690_),
    .Y(_20691_),
    .A1(\u_inv.f_next[85] ),
    .A2(\u_inv.f_reg[85] ));
 sg13g2_nor3_1 _29253_ (.A(_20676_),
    .B(_20680_),
    .C(_20691_),
    .Y(_20692_));
 sg13g2_nor2b_2 _29254_ (.A(_20692_),
    .B_N(_20689_),
    .Y(_20693_));
 sg13g2_nand2_2 _29255_ (.Y(_20694_),
    .A(_20688_),
    .B(_20693_));
 sg13g2_nand2_1 _29256_ (.Y(_20695_),
    .A(\u_inv.f_next[95] ),
    .B(\u_inv.f_reg[95] ));
 sg13g2_xnor2_1 _29257_ (.Y(_20696_),
    .A(\u_inv.f_next[95] ),
    .B(\u_inv.f_reg[95] ));
 sg13g2_inv_1 _29258_ (.Y(_20697_),
    .A(_20696_));
 sg13g2_and2_1 _29259_ (.A(\u_inv.f_next[94] ),
    .B(\u_inv.f_reg[94] ),
    .X(_20698_));
 sg13g2_xor2_1 _29260_ (.B(\u_inv.f_reg[94] ),
    .A(\u_inv.f_next[94] ),
    .X(_20699_));
 sg13g2_nor2b_1 _29261_ (.A(_20696_),
    .B_N(_20699_),
    .Y(_20700_));
 sg13g2_xor2_1 _29262_ (.B(\u_inv.f_reg[93] ),
    .A(\u_inv.f_next[93] ),
    .X(_20701_));
 sg13g2_and2_1 _29263_ (.A(\u_inv.f_next[92] ),
    .B(\u_inv.f_reg[92] ),
    .X(_20702_));
 sg13g2_xor2_1 _29264_ (.B(\u_inv.f_reg[92] ),
    .A(\u_inv.f_next[92] ),
    .X(_20703_));
 sg13g2_and2_1 _29265_ (.A(_20701_),
    .B(_20703_),
    .X(_20704_));
 sg13g2_nand2_1 _29266_ (.Y(_20705_),
    .A(_20700_),
    .B(_20704_));
 sg13g2_xnor2_1 _29267_ (.Y(_20706_),
    .A(\u_inv.f_next[91] ),
    .B(\u_inv.f_reg[91] ));
 sg13g2_nand2_1 _29268_ (.Y(_20707_),
    .A(\u_inv.f_next[90] ),
    .B(\u_inv.f_reg[90] ));
 sg13g2_xnor2_1 _29269_ (.Y(_20708_),
    .A(\u_inv.f_next[90] ),
    .B(\u_inv.f_reg[90] ));
 sg13g2_or2_1 _29270_ (.X(_20709_),
    .B(_20708_),
    .A(_20706_));
 sg13g2_nand2_1 _29271_ (.Y(_20710_),
    .A(\u_inv.f_next[89] ),
    .B(\u_inv.f_reg[89] ));
 sg13g2_nor2_1 _29272_ (.A(\u_inv.f_next[89] ),
    .B(\u_inv.f_reg[89] ),
    .Y(_20711_));
 sg13g2_xor2_1 _29273_ (.B(\u_inv.f_reg[89] ),
    .A(\u_inv.f_next[89] ),
    .X(_20712_));
 sg13g2_xnor2_1 _29274_ (.Y(_20713_),
    .A(\u_inv.f_next[89] ),
    .B(\u_inv.f_reg[89] ));
 sg13g2_nand2_1 _29275_ (.Y(_20714_),
    .A(\u_inv.f_next[88] ),
    .B(\u_inv.f_reg[88] ));
 sg13g2_xor2_1 _29276_ (.B(\u_inv.f_reg[88] ),
    .A(\u_inv.f_next[88] ),
    .X(_20715_));
 sg13g2_nand2_1 _29277_ (.Y(_20716_),
    .A(_20712_),
    .B(_20715_));
 sg13g2_inv_1 _29278_ (.Y(_20717_),
    .A(_20716_));
 sg13g2_or3_1 _29279_ (.A(_20705_),
    .B(_20709_),
    .C(_20716_),
    .X(_20718_));
 sg13g2_a21oi_2 _29280_ (.B1(_20718_),
    .Y(_20719_),
    .A2(_20693_),
    .A1(_20688_));
 sg13g2_o21ai_1 _29281_ (.B1(_20710_),
    .Y(_20720_),
    .A1(_20711_),
    .A2(_20714_));
 sg13g2_nand2b_1 _29282_ (.Y(_20721_),
    .B(_20720_),
    .A_N(_20709_));
 sg13g2_a21oi_1 _29283_ (.A1(_18053_),
    .A2(_18213_),
    .Y(_20722_),
    .B1(_20707_));
 sg13g2_a21oi_1 _29284_ (.A1(\u_inv.f_next[91] ),
    .A2(\u_inv.f_reg[91] ),
    .Y(_20723_),
    .B1(_20722_));
 sg13g2_a21oi_1 _29285_ (.A1(_20721_),
    .A2(_20723_),
    .Y(_20724_),
    .B1(_20705_));
 sg13g2_o21ai_1 _29286_ (.B1(_20698_),
    .Y(_20725_),
    .A1(\u_inv.f_next[95] ),
    .A2(\u_inv.f_reg[95] ));
 sg13g2_a21oi_1 _29287_ (.A1(\u_inv.f_next[93] ),
    .A2(\u_inv.f_reg[93] ),
    .Y(_20726_),
    .B1(_20702_));
 sg13g2_a21oi_1 _29288_ (.A1(_18052_),
    .A2(_18214_),
    .Y(_20727_),
    .B1(_20726_));
 sg13g2_a21oi_1 _29289_ (.A1(_20700_),
    .A2(_20727_),
    .Y(_20728_),
    .B1(_20724_));
 sg13g2_nand3_1 _29290_ (.B(_20725_),
    .C(_20728_),
    .A(_20695_),
    .Y(_20729_));
 sg13g2_nor2_2 _29291_ (.A(_20719_),
    .B(_20729_),
    .Y(_20730_));
 sg13g2_nand2_1 _29292_ (.Y(_20731_),
    .A(\u_inv.f_next[101] ),
    .B(\u_inv.f_reg[101] ));
 sg13g2_xor2_1 _29293_ (.B(\u_inv.f_reg[101] ),
    .A(\u_inv.f_next[101] ),
    .X(_20732_));
 sg13g2_inv_2 _29294_ (.Y(_20733_),
    .A(_20732_));
 sg13g2_nand2_1 _29295_ (.Y(_20734_),
    .A(\u_inv.f_next[100] ),
    .B(\u_inv.f_reg[100] ));
 sg13g2_xor2_1 _29296_ (.B(\u_inv.f_reg[100] ),
    .A(\u_inv.f_next[100] ),
    .X(_20735_));
 sg13g2_inv_2 _29297_ (.Y(_20736_),
    .A(_20735_));
 sg13g2_nor2_1 _29298_ (.A(_20733_),
    .B(_20736_),
    .Y(_20737_));
 sg13g2_nand2_1 _29299_ (.Y(_20738_),
    .A(\u_inv.f_next[103] ),
    .B(\u_inv.f_reg[103] ));
 sg13g2_nor2_1 _29300_ (.A(\u_inv.f_next[103] ),
    .B(\u_inv.f_reg[103] ),
    .Y(_20739_));
 sg13g2_xor2_1 _29301_ (.B(\u_inv.f_reg[103] ),
    .A(\u_inv.f_next[103] ),
    .X(_20740_));
 sg13g2_xnor2_1 _29302_ (.Y(_20741_),
    .A(\u_inv.f_next[103] ),
    .B(\u_inv.f_reg[103] ));
 sg13g2_nand2_1 _29303_ (.Y(_20742_),
    .A(\u_inv.f_next[102] ),
    .B(\u_inv.f_reg[102] ));
 sg13g2_xor2_1 _29304_ (.B(\u_inv.f_reg[102] ),
    .A(\u_inv.f_next[102] ),
    .X(_20743_));
 sg13g2_inv_1 _29305_ (.Y(_20744_),
    .A(_20743_));
 sg13g2_nand2_1 _29306_ (.Y(_20745_),
    .A(_20740_),
    .B(_20743_));
 sg13g2_nor3_1 _29307_ (.A(_20733_),
    .B(_20736_),
    .C(_20745_),
    .Y(_20746_));
 sg13g2_nor2b_1 _29308_ (.A(\u_inv.f_reg[99] ),
    .B_N(\u_inv.f_next[99] ),
    .Y(_20747_));
 sg13g2_xnor2_1 _29309_ (.Y(_20748_),
    .A(\u_inv.f_next[99] ),
    .B(\u_inv.f_reg[99] ));
 sg13g2_and2_1 _29310_ (.A(\u_inv.f_next[98] ),
    .B(\u_inv.f_reg[98] ),
    .X(_20749_));
 sg13g2_xor2_1 _29311_ (.B(\u_inv.f_reg[98] ),
    .A(\u_inv.f_next[98] ),
    .X(_20750_));
 sg13g2_xnor2_1 _29312_ (.Y(_20751_),
    .A(\u_inv.f_next[98] ),
    .B(\u_inv.f_reg[98] ));
 sg13g2_nor2_1 _29313_ (.A(_20748_),
    .B(_20751_),
    .Y(_20752_));
 sg13g2_nand2_1 _29314_ (.Y(_20753_),
    .A(\u_inv.f_next[97] ),
    .B(\u_inv.f_reg[97] ));
 sg13g2_or2_1 _29315_ (.X(_20754_),
    .B(\u_inv.f_reg[97] ),
    .A(\u_inv.f_next[97] ));
 sg13g2_and2_1 _29316_ (.A(_20753_),
    .B(_20754_),
    .X(_20755_));
 sg13g2_nand2_1 _29317_ (.Y(_20756_),
    .A(_20753_),
    .B(_20754_));
 sg13g2_nand2_1 _29318_ (.Y(_20757_),
    .A(\u_inv.f_next[96] ),
    .B(\u_inv.f_reg[96] ));
 sg13g2_xor2_1 _29319_ (.B(\u_inv.f_reg[96] ),
    .A(\u_inv.f_next[96] ),
    .X(_20758_));
 sg13g2_xnor2_1 _29320_ (.Y(_20759_),
    .A(\u_inv.f_next[96] ),
    .B(\u_inv.f_reg[96] ));
 sg13g2_nand2_1 _29321_ (.Y(_20760_),
    .A(_20755_),
    .B(_20758_));
 sg13g2_nand4_1 _29322_ (.B(_20752_),
    .C(_20755_),
    .A(_20746_),
    .Y(_20761_),
    .D(_20758_));
 sg13g2_inv_1 _29323_ (.Y(_20762_),
    .A(_20761_));
 sg13g2_o21ai_1 _29324_ (.B1(_20762_),
    .Y(_20763_),
    .A1(_20719_),
    .A2(_20729_));
 sg13g2_nand2_1 _29325_ (.Y(_20764_),
    .A(_20753_),
    .B(_20757_));
 sg13g2_nand2_1 _29326_ (.Y(_20765_),
    .A(_20754_),
    .B(_20764_));
 sg13g2_nor3_1 _29327_ (.A(_20748_),
    .B(_20751_),
    .C(_20765_),
    .Y(_20766_));
 sg13g2_nor2_1 _29328_ (.A(\u_inv.f_next[99] ),
    .B(\u_inv.f_reg[99] ),
    .Y(_20767_));
 sg13g2_a21oi_1 _29329_ (.A1(\u_inv.f_next[99] ),
    .A2(\u_inv.f_reg[99] ),
    .Y(_20768_),
    .B1(_20749_));
 sg13g2_nor2_1 _29330_ (.A(_20767_),
    .B(_20768_),
    .Y(_20769_));
 sg13g2_o21ai_1 _29331_ (.B1(_20746_),
    .Y(_20770_),
    .A1(_20766_),
    .A2(_20769_));
 sg13g2_o21ai_1 _29332_ (.B1(_20738_),
    .Y(_20771_),
    .A1(_20739_),
    .A2(_20742_));
 sg13g2_nand2_1 _29333_ (.Y(_20772_),
    .A(_20731_),
    .B(_20734_));
 sg13g2_o21ai_1 _29334_ (.B1(_20772_),
    .Y(_20773_),
    .A1(\u_inv.f_next[101] ),
    .A2(\u_inv.f_reg[101] ));
 sg13g2_o21ai_1 _29335_ (.B1(_20770_),
    .Y(_20774_),
    .A1(_20745_),
    .A2(_20773_));
 sg13g2_nor2_2 _29336_ (.A(_20771_),
    .B(_20774_),
    .Y(_20775_));
 sg13g2_nand2_1 _29337_ (.Y(_20776_),
    .A(_20763_),
    .B(_20775_));
 sg13g2_xor2_1 _29338_ (.B(\u_inv.f_reg[111] ),
    .A(\u_inv.f_next[111] ),
    .X(_20777_));
 sg13g2_xnor2_1 _29339_ (.Y(_20778_),
    .A(\u_inv.f_next[111] ),
    .B(\u_inv.f_reg[111] ));
 sg13g2_nand2_1 _29340_ (.Y(_20779_),
    .A(\u_inv.f_next[110] ),
    .B(\u_inv.f_reg[110] ));
 sg13g2_xor2_1 _29341_ (.B(\u_inv.f_reg[110] ),
    .A(\u_inv.f_next[110] ),
    .X(_20780_));
 sg13g2_and2_1 _29342_ (.A(_20777_),
    .B(_20780_),
    .X(_20781_));
 sg13g2_nor2_1 _29343_ (.A(\u_inv.f_next[109] ),
    .B(\u_inv.f_reg[109] ),
    .Y(_20782_));
 sg13g2_nand2_1 _29344_ (.Y(_20783_),
    .A(\u_inv.f_next[109] ),
    .B(\u_inv.f_reg[109] ));
 sg13g2_nand2b_2 _29345_ (.Y(_20784_),
    .B(_20783_),
    .A_N(_20782_));
 sg13g2_nand2_1 _29346_ (.Y(_20785_),
    .A(\u_inv.f_next[108] ),
    .B(\u_inv.f_reg[108] ));
 sg13g2_xor2_1 _29347_ (.B(\u_inv.f_reg[108] ),
    .A(\u_inv.f_next[108] ),
    .X(_20786_));
 sg13g2_xnor2_1 _29348_ (.Y(_20787_),
    .A(\u_inv.f_next[108] ),
    .B(\u_inv.f_reg[108] ));
 sg13g2_nor2_1 _29349_ (.A(_20784_),
    .B(_20787_),
    .Y(_20788_));
 sg13g2_nand2_1 _29350_ (.Y(_20789_),
    .A(_20781_),
    .B(_20788_));
 sg13g2_nand2_1 _29351_ (.Y(_20790_),
    .A(\u_inv.f_next[106] ),
    .B(\u_inv.f_reg[106] ));
 sg13g2_xor2_1 _29352_ (.B(\u_inv.f_reg[106] ),
    .A(\u_inv.f_next[106] ),
    .X(_20791_));
 sg13g2_xnor2_1 _29353_ (.Y(_20792_),
    .A(\u_inv.f_next[106] ),
    .B(\u_inv.f_reg[106] ));
 sg13g2_xor2_1 _29354_ (.B(\u_inv.f_reg[107] ),
    .A(\u_inv.f_next[107] ),
    .X(_20793_));
 sg13g2_nand2_1 _29355_ (.Y(_20794_),
    .A(_20791_),
    .B(_20793_));
 sg13g2_xor2_1 _29356_ (.B(\u_inv.f_reg[105] ),
    .A(\u_inv.f_next[105] ),
    .X(_20795_));
 sg13g2_and2_1 _29357_ (.A(\u_inv.f_next[104] ),
    .B(\u_inv.f_reg[104] ),
    .X(_20796_));
 sg13g2_xor2_1 _29358_ (.B(\u_inv.f_reg[104] ),
    .A(\u_inv.f_next[104] ),
    .X(_20797_));
 sg13g2_nand2_1 _29359_ (.Y(_20798_),
    .A(_20795_),
    .B(_20797_));
 sg13g2_nor3_1 _29360_ (.A(_20789_),
    .B(_20794_),
    .C(_20798_),
    .Y(_20799_));
 sg13g2_inv_1 _29361_ (.Y(_20800_),
    .A(_20799_));
 sg13g2_a21oi_2 _29362_ (.B1(_20800_),
    .Y(_20801_),
    .A2(_20775_),
    .A1(_20763_));
 sg13g2_a21oi_1 _29363_ (.A1(\u_inv.f_next[105] ),
    .A2(\u_inv.f_reg[105] ),
    .Y(_20802_),
    .B1(_20796_));
 sg13g2_a21oi_1 _29364_ (.A1(_18049_),
    .A2(_18216_),
    .Y(_20803_),
    .B1(_20802_));
 sg13g2_nand2b_1 _29365_ (.Y(_20804_),
    .B(_20803_),
    .A_N(_20794_));
 sg13g2_a22oi_1 _29366_ (.Y(_20805_),
    .B1(\u_inv.f_reg[107] ),
    .B2(\u_inv.f_next[107] ),
    .A2(\u_inv.f_reg[106] ),
    .A1(\u_inv.f_next[106] ));
 sg13g2_a21o_1 _29367_ (.A2(_18217_),
    .A1(_18047_),
    .B1(_20805_),
    .X(_20806_));
 sg13g2_a21oi_1 _29368_ (.A1(_20804_),
    .A2(_20806_),
    .Y(_20807_),
    .B1(_20789_));
 sg13g2_a21oi_1 _29369_ (.A1(_18044_),
    .A2(_18218_),
    .Y(_20808_),
    .B1(_20779_));
 sg13g2_o21ai_1 _29370_ (.B1(_20783_),
    .Y(_20809_),
    .A1(_20782_),
    .A2(_20785_));
 sg13g2_a221oi_1 _29371_ (.B2(_20809_),
    .C1(_20808_),
    .B1(_20781_),
    .A1(\u_inv.f_next[111] ),
    .Y(_20810_),
    .A2(\u_inv.f_reg[111] ));
 sg13g2_nand2b_2 _29372_ (.Y(_20811_),
    .B(_20810_),
    .A_N(_20807_));
 sg13g2_nor2_1 _29373_ (.A(_20801_),
    .B(_20811_),
    .Y(_20812_));
 sg13g2_xnor2_1 _29374_ (.Y(_20813_),
    .A(\u_inv.f_next[113] ),
    .B(\u_inv.f_reg[113] ));
 sg13g2_xnor2_1 _29375_ (.Y(_20814_),
    .A(\u_inv.f_next[112] ),
    .B(\u_inv.f_reg[112] ));
 sg13g2_nor2_1 _29376_ (.A(_20813_),
    .B(_20814_),
    .Y(_20815_));
 sg13g2_and3_1 _29377_ (.X(_20816_),
    .A(_20264_),
    .B(_20270_),
    .C(_20815_));
 sg13g2_nand2_1 _29378_ (.Y(_20817_),
    .A(_20250_),
    .B(_20816_));
 sg13g2_inv_1 _29379_ (.Y(_20818_),
    .A(_20817_));
 sg13g2_o21ai_1 _29380_ (.B1(_20818_),
    .Y(_20819_),
    .A1(_20801_),
    .A2(_20811_));
 sg13g2_nor2_1 _29381_ (.A(\u_inv.f_next[129] ),
    .B(\u_inv.f_reg[129] ),
    .Y(_20820_));
 sg13g2_xor2_1 _29382_ (.B(\u_inv.f_reg[129] ),
    .A(\u_inv.f_next[129] ),
    .X(_20821_));
 sg13g2_xnor2_1 _29383_ (.Y(_20822_),
    .A(\u_inv.f_next[128] ),
    .B(\u_inv.f_reg[128] ));
 sg13g2_inv_1 _29384_ (.Y(_20823_),
    .A(_20822_));
 sg13g2_and2_1 _29385_ (.A(\u_inv.f_next[132] ),
    .B(\u_inv.f_reg[132] ),
    .X(_20824_));
 sg13g2_xor2_1 _29386_ (.B(\u_inv.f_reg[132] ),
    .A(\u_inv.f_next[132] ),
    .X(_20825_));
 sg13g2_nor2_1 _29387_ (.A(\u_inv.f_next[133] ),
    .B(\u_inv.f_reg[133] ),
    .Y(_20826_));
 sg13g2_xor2_1 _29388_ (.B(\u_inv.f_reg[133] ),
    .A(\u_inv.f_next[133] ),
    .X(_20827_));
 sg13g2_xnor2_1 _29389_ (.Y(_20828_),
    .A(\u_inv.f_next[133] ),
    .B(\u_inv.f_reg[133] ));
 sg13g2_and2_1 _29390_ (.A(_20825_),
    .B(_20827_),
    .X(_20829_));
 sg13g2_nand2_1 _29391_ (.Y(_20830_),
    .A(\u_inv.f_next[134] ),
    .B(\u_inv.f_reg[134] ));
 sg13g2_xor2_1 _29392_ (.B(\u_inv.f_reg[134] ),
    .A(\u_inv.f_next[134] ),
    .X(_20831_));
 sg13g2_nor2_1 _29393_ (.A(\u_inv.f_next[135] ),
    .B(\u_inv.f_reg[135] ),
    .Y(_20832_));
 sg13g2_xor2_1 _29394_ (.B(\u_inv.f_reg[135] ),
    .A(\u_inv.f_next[135] ),
    .X(_20833_));
 sg13g2_xnor2_1 _29395_ (.Y(_20834_),
    .A(\u_inv.f_next[135] ),
    .B(\u_inv.f_reg[135] ));
 sg13g2_and2_1 _29396_ (.A(_20831_),
    .B(_20833_),
    .X(_20835_));
 sg13g2_and2_1 _29397_ (.A(_20829_),
    .B(_20835_),
    .X(_20836_));
 sg13g2_nand2_1 _29398_ (.Y(_20837_),
    .A(\u_inv.f_next[130] ),
    .B(\u_inv.f_reg[130] ));
 sg13g2_xnor2_1 _29399_ (.Y(_20838_),
    .A(\u_inv.f_next[130] ),
    .B(\u_inv.f_reg[130] ));
 sg13g2_nand2_1 _29400_ (.Y(_20839_),
    .A(\u_inv.f_next[131] ),
    .B(\u_inv.f_reg[131] ));
 sg13g2_xor2_1 _29401_ (.B(\u_inv.f_reg[131] ),
    .A(\u_inv.f_next[131] ),
    .X(_20840_));
 sg13g2_nor2b_1 _29402_ (.A(_20838_),
    .B_N(_20840_),
    .Y(_20841_));
 sg13g2_inv_1 _29403_ (.Y(_20842_),
    .A(_20841_));
 sg13g2_and4_1 _29404_ (.A(_20821_),
    .B(_20823_),
    .C(_20836_),
    .D(_20841_),
    .X(_20843_));
 sg13g2_inv_1 _29405_ (.Y(_20844_),
    .A(_20843_));
 sg13g2_a21oi_2 _29406_ (.B1(_20844_),
    .Y(_20845_),
    .A2(_20819_),
    .A1(_20295_));
 sg13g2_a22oi_1 _29407_ (.Y(_20846_),
    .B1(\u_inv.f_reg[129] ),
    .B2(\u_inv.f_next[129] ),
    .A2(\u_inv.f_reg[128] ),
    .A1(\u_inv.f_next[128] ));
 sg13g2_nor2_1 _29408_ (.A(_20820_),
    .B(_20846_),
    .Y(_20847_));
 sg13g2_nand2_1 _29409_ (.Y(_20848_),
    .A(_20837_),
    .B(_20839_));
 sg13g2_o21ai_1 _29410_ (.B1(_20848_),
    .Y(_20849_),
    .A1(\u_inv.f_next[131] ),
    .A2(\u_inv.f_reg[131] ));
 sg13g2_a22oi_1 _29411_ (.Y(_20850_),
    .B1(\u_inv.f_reg[135] ),
    .B2(\u_inv.f_next[135] ),
    .A2(\u_inv.f_reg[134] ),
    .A1(\u_inv.f_next[134] ));
 sg13g2_a21oi_1 _29412_ (.A1(\u_inv.f_next[133] ),
    .A2(\u_inv.f_reg[133] ),
    .Y(_20851_),
    .B1(_20824_));
 sg13g2_nor2_1 _29413_ (.A(_20826_),
    .B(_20851_),
    .Y(_20852_));
 sg13g2_nand2_1 _29414_ (.Y(_20853_),
    .A(_20841_),
    .B(_20847_));
 sg13g2_nand2_1 _29415_ (.Y(_20854_),
    .A(_20849_),
    .B(_20853_));
 sg13g2_a22oi_1 _29416_ (.Y(_20855_),
    .B1(_20854_),
    .B2(_20836_),
    .A2(_20852_),
    .A1(_20835_));
 sg13g2_o21ai_1 _29417_ (.B1(_20855_),
    .Y(_20856_),
    .A1(_20832_),
    .A2(_20850_));
 sg13g2_nor2_2 _29418_ (.A(\u_inv.f_next[137] ),
    .B(\u_inv.f_reg[137] ),
    .Y(_20857_));
 sg13g2_nand2_2 _29419_ (.Y(_20858_),
    .A(\u_inv.f_next[137] ),
    .B(\u_inv.f_reg[137] ));
 sg13g2_nor2b_2 _29420_ (.A(_20857_),
    .B_N(_20858_),
    .Y(_20859_));
 sg13g2_nand2b_2 _29421_ (.Y(_20860_),
    .B(_20858_),
    .A_N(_20857_));
 sg13g2_nand2_1 _29422_ (.Y(_20861_),
    .A(\u_inv.f_next[136] ),
    .B(\u_inv.f_reg[136] ));
 sg13g2_xor2_1 _29423_ (.B(\u_inv.f_reg[136] ),
    .A(\u_inv.f_next[136] ),
    .X(_20862_));
 sg13g2_xor2_1 _29424_ (.B(\u_inv.f_reg[141] ),
    .A(\u_inv.f_next[141] ),
    .X(_20863_));
 sg13g2_xnor2_1 _29425_ (.Y(_20864_),
    .A(\u_inv.f_next[141] ),
    .B(\u_inv.f_reg[141] ));
 sg13g2_nand2_1 _29426_ (.Y(_20865_),
    .A(\u_inv.f_next[140] ),
    .B(\u_inv.f_reg[140] ));
 sg13g2_xnor2_1 _29427_ (.Y(_20866_),
    .A(\u_inv.f_next[140] ),
    .B(\u_inv.f_reg[140] ));
 sg13g2_nor2_1 _29428_ (.A(_20864_),
    .B(_20866_),
    .Y(_20867_));
 sg13g2_nand2_1 _29429_ (.Y(_20868_),
    .A(\u_inv.f_next[142] ),
    .B(\u_inv.f_reg[142] ));
 sg13g2_nor2_1 _29430_ (.A(\u_inv.f_next[142] ),
    .B(\u_inv.f_reg[142] ),
    .Y(_20869_));
 sg13g2_xor2_1 _29431_ (.B(\u_inv.f_reg[142] ),
    .A(\u_inv.f_next[142] ),
    .X(_20870_));
 sg13g2_nand2_1 _29432_ (.Y(_20871_),
    .A(\u_inv.f_next[143] ),
    .B(\u_inv.f_reg[143] ));
 sg13g2_nor2_1 _29433_ (.A(\u_inv.f_next[143] ),
    .B(\u_inv.f_reg[143] ),
    .Y(_20872_));
 sg13g2_xor2_1 _29434_ (.B(\u_inv.f_reg[143] ),
    .A(\u_inv.f_next[143] ),
    .X(_20873_));
 sg13g2_xnor2_1 _29435_ (.Y(_20874_),
    .A(\u_inv.f_next[143] ),
    .B(\u_inv.f_reg[143] ));
 sg13g2_nand3_1 _29436_ (.B(_20870_),
    .C(_20873_),
    .A(_20867_),
    .Y(_20875_));
 sg13g2_and2_1 _29437_ (.A(\u_inv.f_next[138] ),
    .B(\u_inv.f_reg[138] ),
    .X(_20876_));
 sg13g2_xor2_1 _29438_ (.B(\u_inv.f_reg[138] ),
    .A(\u_inv.f_next[138] ),
    .X(_20877_));
 sg13g2_xor2_1 _29439_ (.B(\u_inv.f_reg[139] ),
    .A(\u_inv.f_next[139] ),
    .X(_20878_));
 sg13g2_xnor2_1 _29440_ (.Y(_20879_),
    .A(\u_inv.f_next[139] ),
    .B(\u_inv.f_reg[139] ));
 sg13g2_and2_1 _29441_ (.A(_20877_),
    .B(_20878_),
    .X(_20880_));
 sg13g2_nand3_1 _29442_ (.B(_20862_),
    .C(_20880_),
    .A(_20859_),
    .Y(_20881_));
 sg13g2_nor2_1 _29443_ (.A(_20875_),
    .B(_20881_),
    .Y(_20882_));
 sg13g2_o21ai_1 _29444_ (.B1(_20882_),
    .Y(_20883_),
    .A1(_20845_),
    .A2(_20856_));
 sg13g2_a21o_1 _29445_ (.A2(_20861_),
    .A1(_20858_),
    .B1(_20857_),
    .X(_20884_));
 sg13g2_a21oi_1 _29446_ (.A1(_20858_),
    .A2(_20861_),
    .Y(_20885_),
    .B1(_20857_));
 sg13g2_a21oi_1 _29447_ (.A1(\u_inv.f_next[139] ),
    .A2(\u_inv.f_reg[139] ),
    .Y(_20886_),
    .B1(_20876_));
 sg13g2_a21oi_1 _29448_ (.A1(_18030_),
    .A2(_18224_),
    .Y(_20887_),
    .B1(_20886_));
 sg13g2_o21ai_1 _29449_ (.B1(_20871_),
    .Y(_20888_),
    .A1(_20868_),
    .A2(_20872_));
 sg13g2_a22oi_1 _29450_ (.Y(_20889_),
    .B1(\u_inv.f_reg[141] ),
    .B2(\u_inv.f_next[141] ),
    .A2(\u_inv.f_reg[140] ),
    .A1(\u_inv.f_next[140] ));
 sg13g2_a21oi_1 _29451_ (.A1(_18029_),
    .A2(_18225_),
    .Y(_20890_),
    .B1(_20889_));
 sg13g2_nand3_1 _29452_ (.B(_20873_),
    .C(_20890_),
    .A(_20870_),
    .Y(_20891_));
 sg13g2_a21oi_1 _29453_ (.A1(_20880_),
    .A2(_20885_),
    .Y(_20892_),
    .B1(_20887_));
 sg13g2_o21ai_1 _29454_ (.B1(_20891_),
    .Y(_20893_),
    .A1(_20875_),
    .A2(_20892_));
 sg13g2_nor2_2 _29455_ (.A(_20888_),
    .B(_20893_),
    .Y(_20894_));
 sg13g2_nand2_2 _29456_ (.Y(_20895_),
    .A(_20883_),
    .B(_20894_));
 sg13g2_or2_1 _29457_ (.X(_20896_),
    .B(\u_inv.f_reg[144] ),
    .A(\u_inv.f_next[144] ));
 sg13g2_and2_1 _29458_ (.A(_20204_),
    .B(_20896_),
    .X(_20897_));
 sg13g2_nor2b_1 _29459_ (.A(_20201_),
    .B_N(_20202_),
    .Y(_20898_));
 sg13g2_nand2b_2 _29460_ (.Y(_20899_),
    .B(_20202_),
    .A_N(_20201_));
 sg13g2_nand2_1 _29461_ (.Y(_20900_),
    .A(_20897_),
    .B(_20898_));
 sg13g2_and4_1 _29462_ (.A(_20194_),
    .B(_20200_),
    .C(_20897_),
    .D(_20898_),
    .X(_20901_));
 sg13g2_and2_1 _29463_ (.A(_20181_),
    .B(_20901_),
    .X(_20902_));
 sg13g2_inv_1 _29464_ (.Y(_20903_),
    .A(_20902_));
 sg13g2_a21oi_2 _29465_ (.B1(_20903_),
    .Y(_20904_),
    .A2(_20894_),
    .A1(_20883_));
 sg13g2_xor2_1 _29466_ (.B(\u_inv.f_reg[160] ),
    .A(\u_inv.f_next[160] ),
    .X(_20905_));
 sg13g2_xnor2_1 _29467_ (.Y(_20906_),
    .A(\u_inv.f_next[160] ),
    .B(\u_inv.f_reg[160] ));
 sg13g2_xor2_1 _29468_ (.B(\u_inv.f_reg[161] ),
    .A(\u_inv.f_next[161] ),
    .X(_20907_));
 sg13g2_xnor2_1 _29469_ (.Y(_20908_),
    .A(\u_inv.f_next[161] ),
    .B(\u_inv.f_reg[161] ));
 sg13g2_nor3_2 _29470_ (.A(_20139_),
    .B(_20906_),
    .C(_20908_),
    .Y(_20909_));
 sg13g2_nand3_1 _29471_ (.B(_20150_),
    .C(_20909_),
    .A(_20091_),
    .Y(_20910_));
 sg13g2_nor3_1 _29472_ (.A(_20113_),
    .B(_20133_),
    .C(_20910_),
    .Y(_20911_));
 sg13g2_o21ai_1 _29473_ (.B1(_20911_),
    .Y(_20912_),
    .A1(_20227_),
    .A2(_20904_));
 sg13g2_xor2_1 _29474_ (.B(\u_inv.f_reg[177] ),
    .A(\u_inv.f_next[177] ),
    .X(_20913_));
 sg13g2_xnor2_1 _29475_ (.Y(_20914_),
    .A(\u_inv.f_next[177] ),
    .B(\u_inv.f_reg[177] ));
 sg13g2_xor2_1 _29476_ (.B(\u_inv.f_reg[176] ),
    .A(\u_inv.f_next[176] ),
    .X(_20915_));
 sg13g2_xnor2_1 _29477_ (.Y(_20916_),
    .A(\u_inv.f_next[176] ),
    .B(\u_inv.f_reg[176] ));
 sg13g2_nor4_1 _29478_ (.A(_20059_),
    .B(_20061_),
    .C(_20914_),
    .D(_20916_),
    .Y(_20917_));
 sg13g2_inv_1 _29479_ (.Y(_20918_),
    .A(_20917_));
 sg13g2_nand3_1 _29480_ (.B(_20082_),
    .C(_20917_),
    .A(_20056_),
    .Y(_20919_));
 sg13g2_a21oi_2 _29481_ (.B1(_20919_),
    .Y(_20920_),
    .A2(_20912_),
    .A1(_20154_));
 sg13g2_a21o_2 _29482_ (.A2(_20912_),
    .A1(_20154_),
    .B1(_20919_),
    .X(_20921_));
 sg13g2_xor2_1 _29483_ (.B(\u_inv.f_reg[193] ),
    .A(\u_inv.f_next[193] ),
    .X(_20922_));
 sg13g2_xor2_1 _29484_ (.B(\u_inv.f_reg[192] ),
    .A(\u_inv.f_next[192] ),
    .X(_20923_));
 sg13g2_xnor2_1 _29485_ (.Y(_20924_),
    .A(\u_inv.f_next[192] ),
    .B(\u_inv.f_reg[192] ));
 sg13g2_nand2_1 _29486_ (.Y(_20925_),
    .A(_20922_),
    .B(_20923_));
 sg13g2_nor3_2 _29487_ (.A(_19988_),
    .B(_19991_),
    .C(_20925_),
    .Y(_20926_));
 sg13g2_and2_1 _29488_ (.A(_20013_),
    .B(_20926_),
    .X(_20927_));
 sg13g2_o21ai_1 _29489_ (.B1(_20927_),
    .Y(_20928_),
    .A1(_20085_),
    .A2(_20920_));
 sg13g2_nand2_1 _29490_ (.Y(_20929_),
    .A(_20016_),
    .B(_20928_));
 sg13g2_a221oi_1 _29491_ (.B2(_20015_),
    .C1(_19900_),
    .B1(_19946_),
    .A1(_19907_),
    .Y(_20930_),
    .A2(_19936_));
 sg13g2_and4_1 _29492_ (.A(_19946_),
    .B(_19958_),
    .C(_20011_),
    .D(_20926_),
    .X(_20931_));
 sg13g2_o21ai_1 _29493_ (.B1(_20931_),
    .Y(_20932_),
    .A1(_20085_),
    .A2(_20920_));
 sg13g2_nand2_1 _29494_ (.Y(_20933_),
    .A(_20930_),
    .B(_20932_));
 sg13g2_xor2_1 _29495_ (.B(\u_inv.f_reg[229] ),
    .A(\u_inv.f_next[229] ),
    .X(_20934_));
 sg13g2_nand2_1 _29496_ (.Y(_20935_),
    .A(\u_inv.f_next[228] ),
    .B(\u_inv.f_reg[228] ));
 sg13g2_xor2_1 _29497_ (.B(\u_inv.f_reg[228] ),
    .A(\u_inv.f_next[228] ),
    .X(_20936_));
 sg13g2_xnor2_1 _29498_ (.Y(_20937_),
    .A(\u_inv.f_next[228] ),
    .B(\u_inv.f_reg[228] ));
 sg13g2_and2_1 _29499_ (.A(_20934_),
    .B(_20936_),
    .X(_20938_));
 sg13g2_and2_1 _29500_ (.A(\u_inv.f_next[230] ),
    .B(\u_inv.f_reg[230] ),
    .X(_20939_));
 sg13g2_xor2_1 _29501_ (.B(\u_inv.f_reg[230] ),
    .A(\u_inv.f_next[230] ),
    .X(_20940_));
 sg13g2_xnor2_1 _29502_ (.Y(_20941_),
    .A(\u_inv.f_next[230] ),
    .B(\u_inv.f_reg[230] ));
 sg13g2_nand2_1 _29503_ (.Y(_20942_),
    .A(\u_inv.f_next[231] ),
    .B(\u_inv.f_reg[231] ));
 sg13g2_xor2_1 _29504_ (.B(\u_inv.f_reg[231] ),
    .A(\u_inv.f_next[231] ),
    .X(_20943_));
 sg13g2_xnor2_1 _29505_ (.Y(_20944_),
    .A(\u_inv.f_next[231] ),
    .B(\u_inv.f_reg[231] ));
 sg13g2_nand2_1 _29506_ (.Y(_20945_),
    .A(_20940_),
    .B(_20943_));
 sg13g2_and3_1 _29507_ (.X(_20946_),
    .A(_20938_),
    .B(_20940_),
    .C(_20943_));
 sg13g2_nor2_1 _29508_ (.A(\u_inv.f_next[227] ),
    .B(\u_inv.f_reg[227] ),
    .Y(_20947_));
 sg13g2_xor2_1 _29509_ (.B(\u_inv.f_reg[227] ),
    .A(\u_inv.f_next[227] ),
    .X(_20948_));
 sg13g2_nand2_1 _29510_ (.Y(_20949_),
    .A(\u_inv.f_next[226] ),
    .B(\u_inv.f_reg[226] ));
 sg13g2_xor2_1 _29511_ (.B(\u_inv.f_reg[226] ),
    .A(\u_inv.f_next[226] ),
    .X(_20950_));
 sg13g2_and2_1 _29512_ (.A(_20948_),
    .B(_20950_),
    .X(_20951_));
 sg13g2_and2_1 _29513_ (.A(\u_inv.f_next[224] ),
    .B(\u_inv.f_reg[224] ),
    .X(_20952_));
 sg13g2_xor2_1 _29514_ (.B(\u_inv.f_reg[224] ),
    .A(\u_inv.f_next[224] ),
    .X(_20953_));
 sg13g2_xor2_1 _29515_ (.B(\u_inv.f_reg[225] ),
    .A(\u_inv.f_next[225] ),
    .X(_20954_));
 sg13g2_xnor2_1 _29516_ (.Y(_20955_),
    .A(\u_inv.f_next[225] ),
    .B(\u_inv.f_reg[225] ));
 sg13g2_nand2_1 _29517_ (.Y(_20956_),
    .A(_20953_),
    .B(_20954_));
 sg13g2_and3_1 _29518_ (.X(_20957_),
    .A(_20951_),
    .B(_20953_),
    .C(_20954_));
 sg13g2_inv_1 _29519_ (.Y(_20958_),
    .A(_20957_));
 sg13g2_nand2_1 _29520_ (.Y(_20959_),
    .A(_20946_),
    .B(_20957_));
 sg13g2_nand2_2 _29521_ (.Y(_20960_),
    .A(\u_inv.f_next[232] ),
    .B(\u_inv.f_reg[232] ));
 sg13g2_xor2_1 _29522_ (.B(\u_inv.f_reg[232] ),
    .A(\u_inv.f_next[232] ),
    .X(_20961_));
 sg13g2_xnor2_1 _29523_ (.Y(_20962_),
    .A(\u_inv.f_next[232] ),
    .B(\u_inv.f_reg[232] ));
 sg13g2_nand2_1 _29524_ (.Y(_20963_),
    .A(\u_inv.f_next[233] ),
    .B(\u_inv.f_reg[233] ));
 sg13g2_nor2_1 _29525_ (.A(\u_inv.f_next[233] ),
    .B(\u_inv.f_reg[233] ),
    .Y(_20964_));
 sg13g2_xor2_1 _29526_ (.B(\u_inv.f_reg[233] ),
    .A(\u_inv.f_next[233] ),
    .X(_20965_));
 sg13g2_and2_1 _29527_ (.A(_20961_),
    .B(_20965_),
    .X(_20966_));
 sg13g2_nand2_1 _29528_ (.Y(_20967_),
    .A(\u_inv.f_next[234] ),
    .B(\u_inv.f_reg[234] ));
 sg13g2_xor2_1 _29529_ (.B(\u_inv.f_reg[234] ),
    .A(\u_inv.f_next[234] ),
    .X(_20968_));
 sg13g2_xnor2_1 _29530_ (.Y(_20969_),
    .A(\u_inv.f_next[234] ),
    .B(\u_inv.f_reg[234] ));
 sg13g2_xor2_1 _29531_ (.B(\u_inv.f_reg[235] ),
    .A(\u_inv.f_next[235] ),
    .X(_20970_));
 sg13g2_and2_1 _29532_ (.A(_20968_),
    .B(_20970_),
    .X(_20971_));
 sg13g2_nand2_2 _29533_ (.Y(_20972_),
    .A(\u_inv.f_next[237] ),
    .B(\u_inv.f_reg[237] ));
 sg13g2_nor2_1 _29534_ (.A(\u_inv.f_next[237] ),
    .B(\u_inv.f_reg[237] ),
    .Y(_20973_));
 sg13g2_or2_1 _29535_ (.X(_20974_),
    .B(\u_inv.f_reg[237] ),
    .A(\u_inv.f_next[237] ));
 sg13g2_nand2_2 _29536_ (.Y(_20975_),
    .A(_20972_),
    .B(_20974_));
 sg13g2_nand2_1 _29537_ (.Y(_20976_),
    .A(\u_inv.f_next[236] ),
    .B(\u_inv.f_reg[236] ));
 sg13g2_inv_1 _29538_ (.Y(_20977_),
    .A(_20976_));
 sg13g2_xor2_1 _29539_ (.B(\u_inv.f_reg[236] ),
    .A(\u_inv.f_next[236] ),
    .X(_20978_));
 sg13g2_xnor2_1 _29540_ (.Y(_20979_),
    .A(\u_inv.f_next[236] ),
    .B(\u_inv.f_reg[236] ));
 sg13g2_nor2_1 _29541_ (.A(_20975_),
    .B(_20979_),
    .Y(_20980_));
 sg13g2_nor2_1 _29542_ (.A(\u_inv.f_next[239] ),
    .B(\u_inv.f_reg[239] ),
    .Y(_20981_));
 sg13g2_xor2_1 _29543_ (.B(\u_inv.f_reg[239] ),
    .A(\u_inv.f_next[239] ),
    .X(_20982_));
 sg13g2_xnor2_1 _29544_ (.Y(_20983_),
    .A(\u_inv.f_next[239] ),
    .B(\u_inv.f_reg[239] ));
 sg13g2_nand2_1 _29545_ (.Y(_20984_),
    .A(\u_inv.f_next[238] ),
    .B(\u_inv.f_reg[238] ));
 sg13g2_xnor2_1 _29546_ (.Y(_20985_),
    .A(\u_inv.f_next[238] ),
    .B(\u_inv.f_reg[238] ));
 sg13g2_nor2_1 _29547_ (.A(_20983_),
    .B(_20985_),
    .Y(_20986_));
 sg13g2_nand2_1 _29548_ (.Y(_20987_),
    .A(_20980_),
    .B(_20986_));
 sg13g2_nand2_1 _29549_ (.Y(_20988_),
    .A(_20966_),
    .B(_20971_));
 sg13g2_or2_1 _29550_ (.X(_20989_),
    .B(_20988_),
    .A(_20987_));
 sg13g2_or2_1 _29551_ (.X(_20990_),
    .B(_20989_),
    .A(_20959_));
 sg13g2_a21oi_2 _29552_ (.B1(_20990_),
    .Y(_20991_),
    .A2(_20932_),
    .A1(_20930_));
 sg13g2_a21o_2 _29553_ (.A2(_20932_),
    .A1(_20930_),
    .B1(_20990_),
    .X(_20992_));
 sg13g2_a21oi_1 _29554_ (.A1(\u_inv.f_next[225] ),
    .A2(\u_inv.f_reg[225] ),
    .Y(_20993_),
    .B1(_20952_));
 sg13g2_a21oi_1 _29555_ (.A1(_17976_),
    .A2(_18250_),
    .Y(_20994_),
    .B1(_20993_));
 sg13g2_a22oi_1 _29556_ (.Y(_20995_),
    .B1(_20951_),
    .B2(_20994_),
    .A2(\u_inv.f_reg[227] ),
    .A1(\u_inv.f_next[227] ));
 sg13g2_o21ai_1 _29557_ (.B1(_20995_),
    .Y(_20996_),
    .A1(_20947_),
    .A2(_20949_));
 sg13g2_o21ai_1 _29558_ (.B1(_20939_),
    .Y(_20997_),
    .A1(\u_inv.f_next[231] ),
    .A2(\u_inv.f_reg[231] ));
 sg13g2_nand2_1 _29559_ (.Y(_20998_),
    .A(_20942_),
    .B(_20997_));
 sg13g2_a22oi_1 _29560_ (.Y(_20999_),
    .B1(\u_inv.f_reg[229] ),
    .B2(\u_inv.f_next[229] ),
    .A2(\u_inv.f_reg[228] ),
    .A1(\u_inv.f_next[228] ));
 sg13g2_a21o_2 _29561_ (.A2(_18251_),
    .A1(_17974_),
    .B1(_20999_),
    .X(_21000_));
 sg13g2_a21oi_1 _29562_ (.A1(_20946_),
    .A2(_20996_),
    .Y(_21001_),
    .B1(_20998_));
 sg13g2_o21ai_1 _29563_ (.B1(_21001_),
    .Y(_21002_),
    .A1(_20945_),
    .A2(_21000_));
 sg13g2_inv_2 _29564_ (.Y(_21003_),
    .A(_21002_));
 sg13g2_nor2_1 _29565_ (.A(_20989_),
    .B(_21003_),
    .Y(_21004_));
 sg13g2_nand2_1 _29566_ (.Y(_21005_),
    .A(_20960_),
    .B(_20963_));
 sg13g2_o21ai_1 _29567_ (.B1(_20963_),
    .Y(_21006_),
    .A1(_20960_),
    .A2(_20964_));
 sg13g2_nand2b_1 _29568_ (.Y(_21007_),
    .B(_21005_),
    .A_N(_20964_));
 sg13g2_o21ai_1 _29569_ (.B1(_20972_),
    .Y(_21008_),
    .A1(_20973_),
    .A2(_20976_));
 sg13g2_inv_1 _29570_ (.Y(_21009_),
    .A(_21008_));
 sg13g2_nor2_1 _29571_ (.A(_20981_),
    .B(_20984_),
    .Y(_21010_));
 sg13g2_a221oi_1 _29572_ (.B2(_21008_),
    .C1(_21010_),
    .B1(_20986_),
    .A1(\u_inv.f_next[239] ),
    .Y(_21011_),
    .A2(\u_inv.f_reg[239] ));
 sg13g2_a21oi_1 _29573_ (.A1(_17973_),
    .A2(_18252_),
    .Y(_21012_),
    .B1(_20967_));
 sg13g2_a221oi_1 _29574_ (.B2(_21006_),
    .C1(_21012_),
    .B1(_20971_),
    .A1(\u_inv.f_next[235] ),
    .Y(_21013_),
    .A2(\u_inv.f_reg[235] ));
 sg13g2_inv_1 _29575_ (.Y(_21014_),
    .A(_21013_));
 sg13g2_nand2b_1 _29576_ (.Y(_21015_),
    .B(_21014_),
    .A_N(_20987_));
 sg13g2_nand3b_1 _29577_ (.B(_21011_),
    .C(_21015_),
    .Y(_21016_),
    .A_N(_21004_));
 sg13g2_inv_2 _29578_ (.Y(_21017_),
    .A(_21016_));
 sg13g2_nand2_1 _29579_ (.Y(_21018_),
    .A(\u_inv.f_next[240] ),
    .B(\u_inv.f_reg[240] ));
 sg13g2_xor2_1 _29580_ (.B(\u_inv.f_reg[240] ),
    .A(\u_inv.f_next[240] ),
    .X(_21019_));
 sg13g2_xnor2_1 _29581_ (.Y(_21020_),
    .A(\u_inv.f_next[240] ),
    .B(\u_inv.f_reg[240] ));
 sg13g2_nand2_1 _29582_ (.Y(_21021_),
    .A(\u_inv.f_next[241] ),
    .B(\u_inv.f_reg[241] ));
 sg13g2_nor2_1 _29583_ (.A(\u_inv.f_next[241] ),
    .B(\u_inv.f_reg[241] ),
    .Y(_21022_));
 sg13g2_xor2_1 _29584_ (.B(\u_inv.f_reg[241] ),
    .A(\u_inv.f_next[241] ),
    .X(_21023_));
 sg13g2_and2_1 _29585_ (.A(_21019_),
    .B(_21023_),
    .X(_21024_));
 sg13g2_nor2_1 _29586_ (.A(\u_inv.f_next[245] ),
    .B(\u_inv.f_reg[245] ),
    .Y(_21025_));
 sg13g2_or2_1 _29587_ (.X(_21026_),
    .B(\u_inv.f_reg[245] ),
    .A(\u_inv.f_next[245] ));
 sg13g2_nand2_1 _29588_ (.Y(_21027_),
    .A(\u_inv.f_next[245] ),
    .B(\u_inv.f_reg[245] ));
 sg13g2_nand2_2 _29589_ (.Y(_21028_),
    .A(_21026_),
    .B(_21027_));
 sg13g2_nand2_1 _29590_ (.Y(_21029_),
    .A(\u_inv.f_next[244] ),
    .B(\u_inv.f_reg[244] ));
 sg13g2_inv_1 _29591_ (.Y(_21030_),
    .A(_21029_));
 sg13g2_xor2_1 _29592_ (.B(\u_inv.f_reg[244] ),
    .A(\u_inv.f_next[244] ),
    .X(_21031_));
 sg13g2_xnor2_1 _29593_ (.Y(_21032_),
    .A(\u_inv.f_next[244] ),
    .B(\u_inv.f_reg[244] ));
 sg13g2_nand3_1 _29594_ (.B(_21027_),
    .C(_21031_),
    .A(_21026_),
    .Y(_21033_));
 sg13g2_nor2_1 _29595_ (.A(\u_inv.f_next[247] ),
    .B(\u_inv.f_reg[247] ),
    .Y(_21034_));
 sg13g2_xor2_1 _29596_ (.B(\u_inv.f_reg[247] ),
    .A(\u_inv.f_next[247] ),
    .X(_21035_));
 sg13g2_xnor2_1 _29597_ (.Y(_21036_),
    .A(\u_inv.f_next[247] ),
    .B(\u_inv.f_reg[247] ));
 sg13g2_nand2_1 _29598_ (.Y(_21037_),
    .A(\u_inv.f_next[246] ),
    .B(\u_inv.f_reg[246] ));
 sg13g2_xor2_1 _29599_ (.B(\u_inv.f_reg[246] ),
    .A(\u_inv.f_next[246] ),
    .X(_21038_));
 sg13g2_nand2_1 _29600_ (.Y(_21039_),
    .A(_21035_),
    .B(_21038_));
 sg13g2_nor2_1 _29601_ (.A(_21033_),
    .B(_21039_),
    .Y(_21040_));
 sg13g2_and2_1 _29602_ (.A(\u_inv.f_next[242] ),
    .B(\u_inv.f_reg[242] ),
    .X(_21041_));
 sg13g2_xor2_1 _29603_ (.B(\u_inv.f_reg[242] ),
    .A(\u_inv.f_next[242] ),
    .X(_21042_));
 sg13g2_xnor2_1 _29604_ (.Y(_21043_),
    .A(\u_inv.f_next[242] ),
    .B(\u_inv.f_reg[242] ));
 sg13g2_xnor2_1 _29605_ (.Y(_21044_),
    .A(\u_inv.f_next[243] ),
    .B(\u_inv.f_reg[243] ));
 sg13g2_nor2_1 _29606_ (.A(_21043_),
    .B(_21044_),
    .Y(_21045_));
 sg13g2_and2_1 _29607_ (.A(_21024_),
    .B(_21045_),
    .X(_21046_));
 sg13g2_and2_1 _29608_ (.A(_21040_),
    .B(_21046_),
    .X(_21047_));
 sg13g2_inv_1 _29609_ (.Y(_21048_),
    .A(_21047_));
 sg13g2_a21oi_1 _29610_ (.A1(_20992_),
    .A2(_21017_),
    .Y(_21049_),
    .B1(_21048_));
 sg13g2_o21ai_1 _29611_ (.B1(_21047_),
    .Y(_21050_),
    .A1(_20991_),
    .A2(_21016_));
 sg13g2_o21ai_1 _29612_ (.B1(_21021_),
    .Y(_21051_),
    .A1(_21018_),
    .A2(_21022_));
 sg13g2_inv_1 _29613_ (.Y(_21052_),
    .A(_21051_));
 sg13g2_o21ai_1 _29614_ (.B1(_21027_),
    .Y(_21053_),
    .A1(_21025_),
    .A2(_21029_));
 sg13g2_nand2b_1 _29615_ (.Y(_21054_),
    .B(_21053_),
    .A_N(_21039_));
 sg13g2_o21ai_1 _29616_ (.B1(_21054_),
    .Y(_21055_),
    .A1(_21034_),
    .A2(_21037_));
 sg13g2_a21oi_1 _29617_ (.A1(\u_inv.f_next[247] ),
    .A2(\u_inv.f_reg[247] ),
    .Y(_21056_),
    .B1(_21055_));
 sg13g2_o21ai_1 _29618_ (.B1(_21041_),
    .Y(_21057_),
    .A1(\u_inv.f_next[243] ),
    .A2(\u_inv.f_reg[243] ));
 sg13g2_a22oi_1 _29619_ (.Y(_21058_),
    .B1(_21045_),
    .B2(_21051_),
    .A2(\u_inv.f_reg[243] ),
    .A1(\u_inv.f_next[243] ));
 sg13g2_and2_1 _29620_ (.A(_21057_),
    .B(_21058_),
    .X(_21059_));
 sg13g2_nand2b_1 _29621_ (.Y(_21060_),
    .B(_21040_),
    .A_N(_21059_));
 sg13g2_nand2_2 _29622_ (.Y(_21061_),
    .A(_21056_),
    .B(_21060_));
 sg13g2_inv_1 _29623_ (.Y(_21062_),
    .A(_21061_));
 sg13g2_xor2_1 _29624_ (.B(\u_inv.f_reg[248] ),
    .A(\u_inv.f_next[248] ),
    .X(_21063_));
 sg13g2_xnor2_1 _29625_ (.Y(_21064_),
    .A(\u_inv.f_next[248] ),
    .B(\u_inv.f_reg[248] ));
 sg13g2_xnor2_1 _29626_ (.Y(_21065_),
    .A(\u_inv.f_next[249] ),
    .B(\u_inv.f_reg[249] ));
 sg13g2_nor2_1 _29627_ (.A(_21064_),
    .B(_21065_),
    .Y(_21066_));
 sg13g2_nand2_1 _29628_ (.Y(_21067_),
    .A(_19861_),
    .B(_21066_));
 sg13g2_a21oi_1 _29629_ (.A1(_21050_),
    .A2(_21062_),
    .Y(_21068_),
    .B1(_21067_));
 sg13g2_o21ai_1 _29630_ (.B1(_19856_),
    .Y(_21069_),
    .A1(_19869_),
    .A2(_21068_));
 sg13g2_a21oi_1 _29631_ (.A1(_19851_),
    .A2(_21069_),
    .Y(_21070_),
    .B1(_19847_));
 sg13g2_nor3_1 _29632_ (.A(_19844_),
    .B(_19845_),
    .C(_21070_),
    .Y(_21071_));
 sg13g2_o21ai_1 _29633_ (.B1(_19844_),
    .Y(_21072_),
    .A1(_19845_),
    .A2(_21070_));
 sg13g2_nand3b_1 _29634_ (.B(_21072_),
    .C(net7311),
    .Y(_21073_),
    .A_N(_21071_));
 sg13g2_a21oi_1 _29635_ (.A1(_17961_),
    .A2(net7183),
    .Y(_21074_),
    .B1(net6280));
 sg13g2_nor2_1 _29636_ (.A(_17962_),
    .B(\u_inv.f_reg[254] ),
    .Y(_21075_));
 sg13g2_inv_1 _29637_ (.Y(_21076_),
    .A(_21075_));
 sg13g2_nand2b_1 _29638_ (.Y(_21077_),
    .B(\u_inv.f_next[252] ),
    .A_N(\u_inv.f_reg[252] ));
 sg13g2_nand2b_1 _29639_ (.Y(_21078_),
    .B(_19853_),
    .A_N(_21077_));
 sg13g2_nand2b_1 _29640_ (.Y(_21079_),
    .B(\u_inv.f_next[253] ),
    .A_N(\u_inv.f_reg[253] ));
 sg13g2_and2_1 _29641_ (.A(_21078_),
    .B(_21079_),
    .X(_21080_));
 sg13g2_nor2_1 _29642_ (.A(_19852_),
    .B(_19854_),
    .Y(_21081_));
 sg13g2_nand2b_1 _29643_ (.Y(_21082_),
    .B(\u_inv.f_next[250] ),
    .A_N(\u_inv.f_reg[250] ));
 sg13g2_nor2_1 _29644_ (.A(_17965_),
    .B(\u_inv.f_reg[248] ),
    .Y(_21083_));
 sg13g2_nand2_1 _29645_ (.Y(_21084_),
    .A(_21065_),
    .B(_21083_));
 sg13g2_o21ai_1 _29646_ (.B1(_21084_),
    .Y(_21085_),
    .A1(_17964_),
    .A2(\u_inv.f_reg[249] ));
 sg13g2_nand2_1 _29647_ (.Y(_21086_),
    .A(_19860_),
    .B(_21085_));
 sg13g2_a21o_1 _29648_ (.A2(_21086_),
    .A1(_21082_),
    .B1(_19857_),
    .X(_21087_));
 sg13g2_o21ai_1 _29649_ (.B1(_21087_),
    .Y(_21088_),
    .A1(_17963_),
    .A2(\u_inv.f_reg[251] ));
 sg13g2_nor2_1 _29650_ (.A(_20542_),
    .B(_20544_),
    .Y(_21089_));
 sg13g2_nand3b_1 _29651_ (.B(_20539_),
    .C(_21089_),
    .Y(_21090_),
    .A_N(_20536_));
 sg13g2_nand2b_1 _29652_ (.Y(_21091_),
    .B(_20550_),
    .A_N(_20548_));
 sg13g2_nor2_1 _29653_ (.A(_20518_),
    .B(_20519_),
    .Y(_21092_));
 sg13g2_nor3_1 _29654_ (.A(_18075_),
    .B(\u_inv.f_reg[54] ),
    .C(_20519_),
    .Y(_21093_));
 sg13g2_nand2b_1 _29655_ (.Y(_21094_),
    .B(\u_inv.f_next[53] ),
    .A_N(\u_inv.f_reg[53] ));
 sg13g2_nor2b_1 _29656_ (.A(\u_inv.f_reg[51] ),
    .B_N(\u_inv.f_next[51] ),
    .Y(_21095_));
 sg13g2_nor2_1 _29657_ (.A(_18076_),
    .B(\u_inv.f_reg[50] ),
    .Y(_21096_));
 sg13g2_nor2b_1 _29658_ (.A(\u_inv.f_reg[49] ),
    .B_N(\u_inv.f_next[49] ),
    .Y(_21097_));
 sg13g2_nor2_1 _29659_ (.A(_20455_),
    .B(_20458_),
    .Y(_21098_));
 sg13g2_nand2b_1 _29660_ (.Y(_21099_),
    .B(\u_inv.f_next[35] ),
    .A_N(\u_inv.f_reg[35] ));
 sg13g2_nand2b_1 _29661_ (.Y(_21100_),
    .B(\u_inv.f_next[34] ),
    .A_N(\u_inv.f_reg[34] ));
 sg13g2_o21ai_1 _29662_ (.B1(_21099_),
    .Y(_21101_),
    .A1(_20458_),
    .A2(_21100_));
 sg13g2_nand2_1 _29663_ (.Y(_21102_),
    .A(\u_inv.f_next[33] ),
    .B(_18201_));
 sg13g2_nor2_1 _29664_ (.A(_18086_),
    .B(\u_inv.f_reg[31] ),
    .Y(_21103_));
 sg13g2_nand2_1 _29665_ (.Y(_21104_),
    .A(\u_inv.f_next[30] ),
    .B(_18199_));
 sg13g2_nand2b_1 _29666_ (.Y(_21105_),
    .B(\u_inv.f_next[27] ),
    .A_N(\u_inv.f_reg[27] ));
 sg13g2_nor3_1 _29667_ (.A(_18090_),
    .B(\u_inv.f_reg[20] ),
    .C(_20419_),
    .Y(_21106_));
 sg13g2_a21oi_1 _29668_ (.A1(\u_inv.f_next[21] ),
    .A2(_18197_),
    .Y(_21107_),
    .B1(_21106_));
 sg13g2_nand2b_1 _29669_ (.Y(_21108_),
    .B(net7300),
    .A_N(\u_inv.f_reg[19] ));
 sg13g2_nor2b_1 _29670_ (.A(\u_inv.f_reg[17] ),
    .B_N(\u_inv.f_next[17] ),
    .Y(_21109_));
 sg13g2_nor2_1 _29671_ (.A(_18091_),
    .B(\u_inv.f_reg[15] ),
    .Y(_21110_));
 sg13g2_xor2_1 _29672_ (.B(\u_inv.f_reg[13] ),
    .A(\u_inv.f_next[13] ),
    .X(_21111_));
 sg13g2_nor2_1 _29673_ (.A(_20366_),
    .B(_20367_),
    .Y(_21112_));
 sg13g2_xor2_1 _29674_ (.B(\u_inv.f_reg[9] ),
    .A(\u_inv.f_next[9] ),
    .X(_21113_));
 sg13g2_inv_1 _29675_ (.Y(_21114_),
    .A(_21113_));
 sg13g2_nor2_1 _29676_ (.A(_18097_),
    .B(\u_inv.f_reg[2] ),
    .Y(_21115_));
 sg13g2_o21ai_1 _29677_ (.B1(_20382_),
    .Y(_21116_),
    .A1(_19830_),
    .A2(_21115_));
 sg13g2_nand2b_1 _29678_ (.Y(_21117_),
    .B(\u_inv.f_next[3] ),
    .A_N(\u_inv.f_reg[3] ));
 sg13g2_a21oi_1 _29679_ (.A1(_21116_),
    .A2(_21117_),
    .Y(_21118_),
    .B1(_20380_));
 sg13g2_nor2_1 _29680_ (.A(_18096_),
    .B(\u_inv.f_reg[4] ),
    .Y(_21119_));
 sg13g2_o21ai_1 _29681_ (.B1(_20378_),
    .Y(_21120_),
    .A1(_21118_),
    .A2(_21119_));
 sg13g2_nand2b_1 _29682_ (.Y(_21121_),
    .B(\u_inv.f_next[5] ),
    .A_N(\u_inv.f_reg[5] ));
 sg13g2_a21oi_1 _29683_ (.A1(_21120_),
    .A2(_21121_),
    .Y(_21122_),
    .B1(_20376_));
 sg13g2_nor2b_1 _29684_ (.A(\u_inv.f_reg[6] ),
    .B_N(\u_inv.f_next[6] ),
    .Y(_21123_));
 sg13g2_o21ai_1 _29685_ (.B1(_20374_),
    .Y(_21124_),
    .A1(_21122_),
    .A2(_21123_));
 sg13g2_nand2_1 _29686_ (.Y(_21125_),
    .A(\u_inv.f_next[7] ),
    .B(_18193_));
 sg13g2_a21oi_1 _29687_ (.A1(_21124_),
    .A2(_21125_),
    .Y(_21126_),
    .B1(_20372_));
 sg13g2_nor2b_1 _29688_ (.A(\u_inv.f_reg[8] ),
    .B_N(\u_inv.f_next[8] ),
    .Y(_21127_));
 sg13g2_o21ai_1 _29689_ (.B1(_21114_),
    .Y(_21128_),
    .A1(_21126_),
    .A2(_21127_));
 sg13g2_nand2_1 _29690_ (.Y(_21129_),
    .A(\u_inv.f_next[9] ),
    .B(_18195_));
 sg13g2_a21o_1 _29691_ (.A2(_21129_),
    .A1(_21128_),
    .B1(_20369_),
    .X(_21130_));
 sg13g2_nand2b_1 _29692_ (.Y(_21131_),
    .B(\u_inv.f_next[10] ),
    .A_N(\u_inv.f_reg[10] ));
 sg13g2_a21oi_1 _29693_ (.A1(_21130_),
    .A2(_21131_),
    .Y(_21132_),
    .B1(_21112_));
 sg13g2_nor2b_1 _29694_ (.A(\u_inv.f_reg[11] ),
    .B_N(\u_inv.f_next[11] ),
    .Y(_21133_));
 sg13g2_o21ai_1 _29695_ (.B1(_20365_),
    .Y(_21134_),
    .A1(_21132_),
    .A2(_21133_));
 sg13g2_nand2b_1 _29696_ (.Y(_21135_),
    .B(\u_inv.f_next[12] ),
    .A_N(\u_inv.f_reg[12] ));
 sg13g2_a21oi_2 _29697_ (.B1(_21111_),
    .Y(_21136_),
    .A2(_21135_),
    .A1(_21134_));
 sg13g2_nor2_1 _29698_ (.A(_18093_),
    .B(\u_inv.f_reg[13] ),
    .Y(_21137_));
 sg13g2_o21ai_1 _29699_ (.B1(_20360_),
    .Y(_21138_),
    .A1(_21136_),
    .A2(_21137_));
 sg13g2_nand2b_1 _29700_ (.Y(_21139_),
    .B(\u_inv.f_next[14] ),
    .A_N(\u_inv.f_reg[14] ));
 sg13g2_nand2_1 _29701_ (.Y(_21140_),
    .A(_21138_),
    .B(_21139_));
 sg13g2_a22oi_1 _29702_ (.Y(_21141_),
    .B1(_21138_),
    .B2(_21139_),
    .A2(\u_inv.f_reg[15] ),
    .A1(_18091_));
 sg13g2_or2_1 _29703_ (.X(_21142_),
    .B(_21141_),
    .A(_21110_));
 sg13g2_nor2b_1 _29704_ (.A(\u_inv.f_reg[16] ),
    .B_N(\u_inv.f_next[16] ),
    .Y(_21143_));
 sg13g2_a21o_1 _29705_ (.A2(_21142_),
    .A1(_20404_),
    .B1(_21143_),
    .X(_21144_));
 sg13g2_and2_1 _29706_ (.A(_20404_),
    .B(_20407_),
    .X(_21145_));
 sg13g2_o21ai_1 _29707_ (.B1(_21145_),
    .Y(_21146_),
    .A1(_21110_),
    .A2(_21141_));
 sg13g2_a21oi_1 _29708_ (.A1(_20407_),
    .A2(_21143_),
    .Y(_21147_),
    .B1(_21109_));
 sg13g2_and2_1 _29709_ (.A(_21146_),
    .B(_21147_),
    .X(_21148_));
 sg13g2_nand2b_1 _29710_ (.Y(_21149_),
    .B(\u_inv.f_next[18] ),
    .A_N(\u_inv.f_reg[18] ));
 sg13g2_o21ai_1 _29711_ (.B1(_21149_),
    .Y(_21150_),
    .A1(_20411_),
    .A2(_21148_));
 sg13g2_nand2b_1 _29712_ (.Y(_21151_),
    .B(_20415_),
    .A_N(_20411_));
 sg13g2_a21oi_1 _29713_ (.A1(_21146_),
    .A2(_21147_),
    .Y(_21152_),
    .B1(_21151_));
 sg13g2_or2_1 _29714_ (.X(_21153_),
    .B(_21151_),
    .A(_21148_));
 sg13g2_nand2_1 _29715_ (.Y(_21154_),
    .A(_20415_),
    .B(_21150_));
 sg13g2_o21ai_1 _29716_ (.B1(_21108_),
    .Y(_21155_),
    .A1(_20414_),
    .A2(_21149_));
 sg13g2_inv_1 _29717_ (.Y(_21156_),
    .A(_21155_));
 sg13g2_a21oi_1 _29718_ (.A1(_21153_),
    .A2(_21156_),
    .Y(_21157_),
    .B1(_20421_));
 sg13g2_a21oi_1 _29719_ (.A1(\u_inv.f_next[20] ),
    .A2(_18196_),
    .Y(_21158_),
    .B1(_21157_));
 sg13g2_nor2_1 _29720_ (.A(_20419_),
    .B(_21158_),
    .Y(_21159_));
 sg13g2_a21oi_1 _29721_ (.A1(\u_inv.f_next[21] ),
    .A2(_18197_),
    .Y(_21160_),
    .B1(_21159_));
 sg13g2_nor2b_1 _29722_ (.A(\u_inv.f_reg[23] ),
    .B_N(\u_inv.f_next[23] ),
    .Y(_21161_));
 sg13g2_nand2_1 _29723_ (.Y(_21162_),
    .A(\u_inv.f_next[22] ),
    .B(_18198_));
 sg13g2_o21ai_1 _29724_ (.B1(_21162_),
    .Y(_21163_),
    .A1(_20345_),
    .A2(_21107_));
 sg13g2_a21oi_1 _29725_ (.A1(_20349_),
    .A2(_21163_),
    .Y(_21164_),
    .B1(_21161_));
 sg13g2_nor4_1 _29726_ (.A(_20345_),
    .B(_20348_),
    .C(_20419_),
    .D(_20421_),
    .Y(_21165_));
 sg13g2_o21ai_1 _29727_ (.B1(_21165_),
    .Y(_21166_),
    .A1(_21152_),
    .A2(_21155_));
 sg13g2_a21oi_1 _29728_ (.A1(_21164_),
    .A2(_21166_),
    .Y(_21167_),
    .B1(_20431_));
 sg13g2_nor2_1 _29729_ (.A(_18088_),
    .B(\u_inv.f_reg[24] ),
    .Y(_21168_));
 sg13g2_o21ai_1 _29730_ (.B1(_20434_),
    .Y(_21169_),
    .A1(_21167_),
    .A2(_21168_));
 sg13g2_nand2b_1 _29731_ (.Y(_21170_),
    .B(\u_inv.f_next[25] ),
    .A_N(\u_inv.f_reg[25] ));
 sg13g2_and2_1 _29732_ (.A(_21169_),
    .B(_21170_),
    .X(_21171_));
 sg13g2_nand2b_1 _29733_ (.Y(_21172_),
    .B(\u_inv.f_next[26] ),
    .A_N(\u_inv.f_reg[26] ));
 sg13g2_nor2_1 _29734_ (.A(_20438_),
    .B(_20440_),
    .Y(_21173_));
 sg13g2_inv_1 _29735_ (.Y(_21174_),
    .A(_21173_));
 sg13g2_a21oi_1 _29736_ (.A1(_21169_),
    .A2(_21170_),
    .Y(_21175_),
    .B1(_21174_));
 sg13g2_o21ai_1 _29737_ (.B1(_21105_),
    .Y(_21176_),
    .A1(_20440_),
    .A2(_21172_));
 sg13g2_nor2_1 _29738_ (.A(_21175_),
    .B(_21176_),
    .Y(_21177_));
 sg13g2_nor2_1 _29739_ (.A(_20446_),
    .B(_21177_),
    .Y(_21178_));
 sg13g2_nand2_1 _29740_ (.Y(_21179_),
    .A(_20444_),
    .B(_21178_));
 sg13g2_nor2b_1 _29741_ (.A(\u_inv.f_reg[28] ),
    .B_N(\u_inv.f_next[28] ),
    .Y(_21180_));
 sg13g2_nor2b_1 _29742_ (.A(\u_inv.f_reg[29] ),
    .B_N(\u_inv.f_next[29] ),
    .Y(_21181_));
 sg13g2_a21oi_1 _29743_ (.A1(_20444_),
    .A2(_21180_),
    .Y(_21182_),
    .B1(_21181_));
 sg13g2_o21ai_1 _29744_ (.B1(_21104_),
    .Y(_21183_),
    .A1(_20329_),
    .A2(_21182_));
 sg13g2_a21oi_1 _29745_ (.A1(_20333_),
    .A2(_21183_),
    .Y(_21184_),
    .B1(_21103_));
 sg13g2_nor4_1 _29746_ (.A(_20329_),
    .B(_20332_),
    .C(_20443_),
    .D(_20446_),
    .Y(_21185_));
 sg13g2_o21ai_1 _29747_ (.B1(_21185_),
    .Y(_21186_),
    .A1(_21175_),
    .A2(_21176_));
 sg13g2_nand2_1 _29748_ (.Y(_21187_),
    .A(_21184_),
    .B(_21186_));
 sg13g2_nand2_1 _29749_ (.Y(_21188_),
    .A(_20461_),
    .B(_21187_));
 sg13g2_nand2_1 _29750_ (.Y(_21189_),
    .A(\u_inv.f_next[32] ),
    .B(_18200_));
 sg13g2_nand3b_1 _29751_ (.B(_20461_),
    .C(_21098_),
    .Y(_21190_),
    .A_N(_20460_));
 sg13g2_a21oi_1 _29752_ (.A1(_21184_),
    .A2(_21186_),
    .Y(_21191_),
    .B1(_21190_));
 sg13g2_o21ai_1 _29753_ (.B1(_21102_),
    .Y(_21192_),
    .A1(_20460_),
    .A2(_21189_));
 sg13g2_a21oi_1 _29754_ (.A1(_21098_),
    .A2(_21192_),
    .Y(_21193_),
    .B1(_21101_));
 sg13g2_inv_1 _29755_ (.Y(_21194_),
    .A(_21193_));
 sg13g2_nand2b_1 _29756_ (.Y(_21195_),
    .B(_21193_),
    .A_N(_21191_));
 sg13g2_and2_1 _29757_ (.A(_20473_),
    .B(_20475_),
    .X(_21196_));
 sg13g2_nand3_1 _29758_ (.B(_20482_),
    .C(_21196_),
    .A(_20478_),
    .Y(_21197_));
 sg13g2_inv_1 _29759_ (.Y(_21198_),
    .A(_21197_));
 sg13g2_o21ai_1 _29760_ (.B1(_21198_),
    .Y(_21199_),
    .A1(_21191_),
    .A2(_21194_));
 sg13g2_nor2_1 _29761_ (.A(_18081_),
    .B(\u_inv.f_reg[39] ),
    .Y(_21200_));
 sg13g2_nor2_1 _29762_ (.A(_18082_),
    .B(\u_inv.f_reg[38] ),
    .Y(_21201_));
 sg13g2_nand2b_1 _29763_ (.Y(_21202_),
    .B(\u_inv.f_next[36] ),
    .A_N(\u_inv.f_reg[36] ));
 sg13g2_nor2_1 _29764_ (.A(_20481_),
    .B(_21202_),
    .Y(_21203_));
 sg13g2_nor2b_1 _29765_ (.A(\u_inv.f_reg[37] ),
    .B_N(\u_inv.f_next[37] ),
    .Y(_21204_));
 sg13g2_or2_1 _29766_ (.X(_21205_),
    .B(_21204_),
    .A(_21203_));
 sg13g2_a221oi_1 _29767_ (.B2(_21196_),
    .C1(_21200_),
    .B1(_21205_),
    .A1(_20473_),
    .Y(_21206_),
    .A2(_21201_));
 sg13g2_nand2_1 _29768_ (.Y(_21207_),
    .A(_21199_),
    .B(_21206_));
 sg13g2_nand3_1 _29769_ (.B(_20313_),
    .C(_20491_),
    .A(_20309_),
    .Y(_21208_));
 sg13g2_nand2_1 _29770_ (.Y(_21209_),
    .A(_20296_),
    .B(_20298_));
 sg13g2_nand2b_1 _29771_ (.Y(_21210_),
    .B(_20490_),
    .A_N(_20301_));
 sg13g2_nor4_1 _29772_ (.A(_20304_),
    .B(_21208_),
    .C(_21209_),
    .D(_21210_),
    .Y(_21211_));
 sg13g2_inv_1 _29773_ (.Y(_21212_),
    .A(_21211_));
 sg13g2_a21oi_2 _29774_ (.B1(_21212_),
    .Y(_21213_),
    .A2(_21206_),
    .A1(_21199_));
 sg13g2_nor2b_1 _29775_ (.A(\u_inv.f_reg[46] ),
    .B_N(\u_inv.f_next[46] ),
    .Y(_21214_));
 sg13g2_nor2_1 _29776_ (.A(_18078_),
    .B(\u_inv.f_reg[47] ),
    .Y(_21215_));
 sg13g2_a21oi_1 _29777_ (.A1(_20296_),
    .A2(_21214_),
    .Y(_21216_),
    .B1(_21215_));
 sg13g2_nand2b_1 _29778_ (.Y(_21217_),
    .B(\u_inv.f_next[40] ),
    .A_N(\u_inv.f_reg[40] ));
 sg13g2_nand2b_1 _29779_ (.Y(_21218_),
    .B(_20491_),
    .A_N(_21217_));
 sg13g2_nand2b_1 _29780_ (.Y(_21219_),
    .B(\u_inv.f_next[41] ),
    .A_N(\u_inv.f_reg[41] ));
 sg13g2_a21oi_1 _29781_ (.A1(_21218_),
    .A2(_21219_),
    .Y(_21220_),
    .B1(_20312_));
 sg13g2_nand2b_1 _29782_ (.Y(_21221_),
    .B(\u_inv.f_next[42] ),
    .A_N(\u_inv.f_reg[42] ));
 sg13g2_nand2b_1 _29783_ (.Y(_21222_),
    .B(_21221_),
    .A_N(_21220_));
 sg13g2_a21oi_1 _29784_ (.A1(_20309_),
    .A2(_21222_),
    .Y(_21223_),
    .B1(_20308_));
 sg13g2_nand2b_1 _29785_ (.Y(_21224_),
    .B(\u_inv.f_next[44] ),
    .A_N(\u_inv.f_reg[44] ));
 sg13g2_o21ai_1 _29786_ (.B1(_21224_),
    .Y(_21225_),
    .A1(_20301_),
    .A2(_21223_));
 sg13g2_nor2_1 _29787_ (.A(_18079_),
    .B(\u_inv.f_reg[45] ),
    .Y(_21226_));
 sg13g2_a21oi_1 _29788_ (.A1(_20305_),
    .A2(_21225_),
    .Y(_21227_),
    .B1(_21226_));
 sg13g2_o21ai_1 _29789_ (.B1(_21216_),
    .Y(_21228_),
    .A1(_21209_),
    .A2(_21227_));
 sg13g2_nor2_1 _29790_ (.A(_21213_),
    .B(_21228_),
    .Y(_21229_));
 sg13g2_o21ai_1 _29791_ (.B1(_20502_),
    .Y(_21230_),
    .A1(_21213_),
    .A2(_21228_));
 sg13g2_nand2b_1 _29792_ (.Y(_21231_),
    .B(\u_inv.f_next[48] ),
    .A_N(\u_inv.f_reg[48] ));
 sg13g2_and4_1 _29793_ (.A(_20500_),
    .B(_20502_),
    .C(_20508_),
    .D(_20509_),
    .X(_21232_));
 sg13g2_o21ai_1 _29794_ (.B1(_21232_),
    .Y(_21233_),
    .A1(_21213_),
    .A2(_21228_));
 sg13g2_nor2_1 _29795_ (.A(_20499_),
    .B(_21231_),
    .Y(_21234_));
 sg13g2_or2_1 _29796_ (.X(_21235_),
    .B(_21234_),
    .A(_21097_));
 sg13g2_a21o_1 _29797_ (.A2(_21235_),
    .A1(_20508_),
    .B1(_21096_),
    .X(_21236_));
 sg13g2_a21oi_1 _29798_ (.A1(_20509_),
    .A2(_21236_),
    .Y(_21237_),
    .B1(_21095_));
 sg13g2_a21oi_1 _29799_ (.A1(_21233_),
    .A2(_21237_),
    .Y(_21238_),
    .B1(_20525_));
 sg13g2_nand2b_1 _29800_ (.Y(_21239_),
    .B(\u_inv.f_next[52] ),
    .A_N(\u_inv.f_reg[52] ));
 sg13g2_nand3_1 _29801_ (.B(_20526_),
    .C(_21092_),
    .A(_20523_),
    .Y(_21240_));
 sg13g2_a21oi_1 _29802_ (.A1(_21233_),
    .A2(_21237_),
    .Y(_21241_),
    .B1(_21240_));
 sg13g2_o21ai_1 _29803_ (.B1(_21094_),
    .Y(_21242_),
    .A1(_20522_),
    .A2(_21239_));
 sg13g2_a221oi_1 _29804_ (.B2(_21242_),
    .C1(_21093_),
    .B1(_21092_),
    .A1(\u_inv.f_next[55] ),
    .Y(_21243_),
    .A2(_18205_));
 sg13g2_inv_1 _29805_ (.Y(_21244_),
    .A(_21243_));
 sg13g2_nand2b_2 _29806_ (.Y(_21245_),
    .B(_21243_),
    .A_N(_21241_));
 sg13g2_nand3_1 _29807_ (.B(_20559_),
    .C(_21245_),
    .A(_20556_),
    .Y(_21246_));
 sg13g2_or2_1 _29808_ (.X(_21247_),
    .B(_21246_),
    .A(_21091_));
 sg13g2_nor4_1 _29809_ (.A(_20555_),
    .B(_20558_),
    .C(_21090_),
    .D(_21091_),
    .Y(_21248_));
 sg13g2_o21ai_1 _29810_ (.B1(_21248_),
    .Y(_21249_),
    .A1(_21241_),
    .A2(_21244_));
 sg13g2_nand2b_1 _29811_ (.Y(_21250_),
    .B(\u_inv.f_next[62] ),
    .A_N(\u_inv.f_reg[62] ));
 sg13g2_nand2b_1 _29812_ (.Y(_21251_),
    .B(\u_inv.f_next[61] ),
    .A_N(\u_inv.f_reg[61] ));
 sg13g2_nor2b_1 _29813_ (.A(\u_inv.f_reg[60] ),
    .B_N(\u_inv.f_next[60] ),
    .Y(_21252_));
 sg13g2_nand2b_1 _29814_ (.Y(_21253_),
    .B(\u_inv.f_next[56] ),
    .A_N(\u_inv.f_reg[56] ));
 sg13g2_nand2b_1 _29815_ (.Y(_21254_),
    .B(_20556_),
    .A_N(_21253_));
 sg13g2_nand2b_1 _29816_ (.Y(_21255_),
    .B(\u_inv.f_next[57] ),
    .A_N(\u_inv.f_reg[57] ));
 sg13g2_a21oi_1 _29817_ (.A1(_21254_),
    .A2(_21255_),
    .Y(_21256_),
    .B1(_20551_));
 sg13g2_nor2_1 _29818_ (.A(_20549_),
    .B(_21256_),
    .Y(_21257_));
 sg13g2_o21ai_1 _29819_ (.B1(_20547_),
    .Y(_21258_),
    .A1(_20548_),
    .A2(_21257_));
 sg13g2_inv_1 _29820_ (.Y(_21259_),
    .A(_21258_));
 sg13g2_a21oi_1 _29821_ (.A1(_20539_),
    .A2(_21258_),
    .Y(_21260_),
    .B1(_21252_));
 sg13g2_o21ai_1 _29822_ (.B1(_21251_),
    .Y(_21261_),
    .A1(_20536_),
    .A2(_21260_));
 sg13g2_a22oi_1 _29823_ (.Y(_21262_),
    .B1(_21089_),
    .B2(_21261_),
    .A2(_18207_),
    .A1(\u_inv.f_next[63] ));
 sg13g2_o21ai_1 _29824_ (.B1(_21262_),
    .Y(_21263_),
    .A1(_20542_),
    .A2(_21250_));
 sg13g2_inv_1 _29825_ (.Y(_21264_),
    .A(_21263_));
 sg13g2_nand2_1 _29826_ (.Y(_21265_),
    .A(_21249_),
    .B(_21264_));
 sg13g2_nand4_1 _29827_ (.B(_20582_),
    .C(_20584_),
    .A(_20579_),
    .Y(_21266_),
    .D(_20586_));
 sg13g2_a21oi_1 _29828_ (.A1(_21249_),
    .A2(_21264_),
    .Y(_21267_),
    .B1(_21266_));
 sg13g2_nor2b_1 _29829_ (.A(\u_inv.f_reg[64] ),
    .B_N(\u_inv.f_next[64] ),
    .Y(_21268_));
 sg13g2_nor2b_1 _29830_ (.A(\u_inv.f_reg[65] ),
    .B_N(\u_inv.f_next[65] ),
    .Y(_21269_));
 sg13g2_a21oi_1 _29831_ (.A1(_20584_),
    .A2(_21268_),
    .Y(_21270_),
    .B1(_21269_));
 sg13g2_nand2b_1 _29832_ (.Y(_21271_),
    .B(\u_inv.f_next[66] ),
    .A_N(\u_inv.f_reg[66] ));
 sg13g2_o21ai_1 _29833_ (.B1(_21271_),
    .Y(_21272_),
    .A1(_20578_),
    .A2(_21270_));
 sg13g2_nor2_1 _29834_ (.A(_18068_),
    .B(\u_inv.f_reg[67] ),
    .Y(_21273_));
 sg13g2_a21oi_1 _29835_ (.A1(_20582_),
    .A2(_21272_),
    .Y(_21274_),
    .B1(_21273_));
 sg13g2_inv_1 _29836_ (.Y(_21275_),
    .A(_21274_));
 sg13g2_nand2b_2 _29837_ (.Y(_21276_),
    .B(_21274_),
    .A_N(_21267_));
 sg13g2_nor2_1 _29838_ (.A(_20602_),
    .B(_20605_),
    .Y(_21277_));
 sg13g2_and3_1 _29839_ (.X(_21278_),
    .A(_20597_),
    .B(_20600_),
    .C(_21277_));
 sg13g2_o21ai_1 _29840_ (.B1(_21278_),
    .Y(_21279_),
    .A1(_21267_),
    .A2(_21275_));
 sg13g2_nand2b_1 _29841_ (.Y(_21280_),
    .B(\u_inv.f_next[71] ),
    .A_N(\u_inv.f_reg[71] ));
 sg13g2_nor2_1 _29842_ (.A(_18066_),
    .B(\u_inv.f_reg[70] ),
    .Y(_21281_));
 sg13g2_nor2b_1 _29843_ (.A(\u_inv.f_reg[68] ),
    .B_N(\u_inv.f_next[68] ),
    .Y(_21282_));
 sg13g2_nand2_1 _29844_ (.Y(_21283_),
    .A(_20603_),
    .B(_21282_));
 sg13g2_o21ai_1 _29845_ (.B1(_21283_),
    .Y(_21284_),
    .A1(_18067_),
    .A2(\u_inv.f_reg[69] ));
 sg13g2_a21oi_1 _29846_ (.A1(_20597_),
    .A2(_21284_),
    .Y(_21285_),
    .B1(_21281_));
 sg13g2_o21ai_1 _29847_ (.B1(_21280_),
    .Y(_21286_),
    .A1(_20599_),
    .A2(_21285_));
 sg13g2_inv_1 _29848_ (.Y(_21287_),
    .A(_21286_));
 sg13g2_and2_1 _29849_ (.A(_21279_),
    .B(_21287_),
    .X(_21288_));
 sg13g2_or2_1 _29850_ (.X(_21289_),
    .B(_20636_),
    .A(_20634_));
 sg13g2_nor2_1 _29851_ (.A(_20616_),
    .B(_20620_),
    .Y(_21290_));
 sg13g2_nand2_1 _29852_ (.Y(_21291_),
    .A(_20629_),
    .B(_20632_));
 sg13g2_nor3_1 _29853_ (.A(_20622_),
    .B(_20624_),
    .C(_21291_),
    .Y(_21292_));
 sg13g2_nand3b_1 _29854_ (.B(_21290_),
    .C(_21292_),
    .Y(_21293_),
    .A_N(_21289_));
 sg13g2_a21oi_1 _29855_ (.A1(_21279_),
    .A2(_21287_),
    .Y(_21294_),
    .B1(_21293_));
 sg13g2_nand2b_1 _29856_ (.Y(_21295_),
    .B(\u_inv.f_next[72] ),
    .A_N(\u_inv.f_reg[72] ));
 sg13g2_nor2_1 _29857_ (.A(_20634_),
    .B(_21295_),
    .Y(_21296_));
 sg13g2_a21oi_1 _29858_ (.A1(\u_inv.f_next[73] ),
    .A2(_18209_),
    .Y(_21297_),
    .B1(_21296_));
 sg13g2_nor2b_1 _29859_ (.A(\u_inv.f_reg[74] ),
    .B_N(\u_inv.f_next[74] ),
    .Y(_21298_));
 sg13g2_nor2b_1 _29860_ (.A(\u_inv.f_reg[75] ),
    .B_N(\u_inv.f_next[75] ),
    .Y(_21299_));
 sg13g2_a21oi_1 _29861_ (.A1(_20629_),
    .A2(_21298_),
    .Y(_21300_),
    .B1(_21299_));
 sg13g2_o21ai_1 _29862_ (.B1(_21300_),
    .Y(_21301_),
    .A1(_21291_),
    .A2(_21297_));
 sg13g2_nand2_1 _29863_ (.Y(_21302_),
    .A(\u_inv.f_next[77] ),
    .B(_18210_));
 sg13g2_nor2b_1 _29864_ (.A(\u_inv.f_reg[76] ),
    .B_N(\u_inv.f_next[76] ),
    .Y(_21303_));
 sg13g2_a21oi_1 _29865_ (.A1(_20623_),
    .A2(_21301_),
    .Y(_21304_),
    .B1(_21303_));
 sg13g2_o21ai_1 _29866_ (.B1(_21302_),
    .Y(_21305_),
    .A1(_20624_),
    .A2(_21304_));
 sg13g2_nor2_1 _29867_ (.A(_18062_),
    .B(\u_inv.f_reg[79] ),
    .Y(_21306_));
 sg13g2_nor2_1 _29868_ (.A(_18063_),
    .B(\u_inv.f_reg[78] ),
    .Y(_21307_));
 sg13g2_a221oi_1 _29869_ (.B2(_20617_),
    .C1(_21306_),
    .B1(_21307_),
    .A1(_21290_),
    .Y(_21308_),
    .A2(_21305_));
 sg13g2_inv_1 _29870_ (.Y(_21309_),
    .A(_21308_));
 sg13g2_nand2b_1 _29871_ (.Y(_21310_),
    .B(_21308_),
    .A_N(_21294_));
 sg13g2_and2_1 _29872_ (.A(_20656_),
    .B(_20658_),
    .X(_21311_));
 sg13g2_o21ai_1 _29873_ (.B1(_21311_),
    .Y(_21312_),
    .A1(_21294_),
    .A2(_21309_));
 sg13g2_nand2b_1 _29874_ (.Y(_21313_),
    .B(\u_inv.f_next[80] ),
    .A_N(\u_inv.f_reg[80] ));
 sg13g2_nor2_1 _29875_ (.A(_20655_),
    .B(_21313_),
    .Y(_21314_));
 sg13g2_a21oi_1 _29876_ (.A1(\u_inv.f_next[81] ),
    .A2(_18211_),
    .Y(_21315_),
    .B1(_21314_));
 sg13g2_nand2_1 _29877_ (.Y(_21316_),
    .A(_21312_),
    .B(_21315_));
 sg13g2_nand2b_1 _29878_ (.Y(_21317_),
    .B(_20669_),
    .A_N(_20666_));
 sg13g2_a21oi_1 _29879_ (.A1(_21312_),
    .A2(_21315_),
    .Y(_21318_),
    .B1(_21317_));
 sg13g2_nand2b_1 _29880_ (.Y(_21319_),
    .B(\u_inv.f_next[82] ),
    .A_N(\u_inv.f_reg[82] ));
 sg13g2_nand2b_1 _29881_ (.Y(_21320_),
    .B(\u_inv.f_next[83] ),
    .A_N(\u_inv.f_reg[83] ));
 sg13g2_o21ai_1 _29882_ (.B1(_21320_),
    .Y(_21321_),
    .A1(_20666_),
    .A2(_21319_));
 sg13g2_or2_1 _29883_ (.X(_21322_),
    .B(_21321_),
    .A(_21318_));
 sg13g2_nor4_1 _29884_ (.A(_20675_),
    .B(_20679_),
    .C(_20682_),
    .D(_20684_),
    .Y(_21323_));
 sg13g2_o21ai_1 _29885_ (.B1(_21323_),
    .Y(_21324_),
    .A1(_21318_),
    .A2(_21321_));
 sg13g2_nor2_1 _29886_ (.A(_18058_),
    .B(\u_inv.f_reg[84] ),
    .Y(_21325_));
 sg13g2_nor3_1 _29887_ (.A(_18058_),
    .B(\u_inv.f_reg[84] ),
    .C(_20682_),
    .Y(_21326_));
 sg13g2_nor2b_1 _29888_ (.A(\u_inv.f_reg[85] ),
    .B_N(\u_inv.f_next[85] ),
    .Y(_21327_));
 sg13g2_nor2_1 _29889_ (.A(_21326_),
    .B(_21327_),
    .Y(_21328_));
 sg13g2_nand2b_1 _29890_ (.Y(_21329_),
    .B(\u_inv.f_next[86] ),
    .A_N(\u_inv.f_reg[86] ));
 sg13g2_o21ai_1 _29891_ (.B1(_21329_),
    .Y(_21330_),
    .A1(_20675_),
    .A2(_21328_));
 sg13g2_nor2_1 _29892_ (.A(_18056_),
    .B(\u_inv.f_reg[87] ),
    .Y(_21331_));
 sg13g2_a21oi_1 _29893_ (.A1(_20680_),
    .A2(_21330_),
    .Y(_21332_),
    .B1(_21331_));
 sg13g2_and2_1 _29894_ (.A(_21324_),
    .B(_21332_),
    .X(_21333_));
 sg13g2_nor2_1 _29895_ (.A(_20701_),
    .B(_20703_),
    .Y(_21334_));
 sg13g2_and2_1 _29896_ (.A(_20706_),
    .B(_20708_),
    .X(_21335_));
 sg13g2_nor2_1 _29897_ (.A(_20712_),
    .B(_20715_),
    .Y(_21336_));
 sg13g2_nor2_1 _29898_ (.A(_20697_),
    .B(_20699_),
    .Y(_21337_));
 sg13g2_nand4_1 _29899_ (.B(_21335_),
    .C(_21336_),
    .A(_21334_),
    .Y(_21338_),
    .D(_21337_));
 sg13g2_a21o_2 _29900_ (.A2(_21332_),
    .A1(_21324_),
    .B1(_21338_),
    .X(_21339_));
 sg13g2_nand2_1 _29901_ (.Y(_21340_),
    .A(\u_inv.f_next[93] ),
    .B(_18214_));
 sg13g2_nand2b_1 _29902_ (.Y(_21341_),
    .B(\u_inv.f_next[92] ),
    .A_N(\u_inv.f_reg[92] ));
 sg13g2_nor2_1 _29903_ (.A(_18054_),
    .B(\u_inv.f_reg[90] ),
    .Y(_21342_));
 sg13g2_nand3_1 _29904_ (.B(_18212_),
    .C(_20713_),
    .A(\u_inv.f_next[88] ),
    .Y(_21343_));
 sg13g2_o21ai_1 _29905_ (.B1(_21343_),
    .Y(_21344_),
    .A1(_18055_),
    .A2(\u_inv.f_reg[89] ));
 sg13g2_and2_1 _29906_ (.A(_20708_),
    .B(_21344_),
    .X(_21345_));
 sg13g2_o21ai_1 _29907_ (.B1(_20706_),
    .Y(_21346_),
    .A1(_21342_),
    .A2(_21345_));
 sg13g2_o21ai_1 _29908_ (.B1(_21346_),
    .Y(_21347_),
    .A1(_18053_),
    .A2(\u_inv.f_reg[91] ));
 sg13g2_o21ai_1 _29909_ (.B1(_21340_),
    .Y(_21348_),
    .A1(_20701_),
    .A2(_21341_));
 sg13g2_a21o_1 _29910_ (.A2(_21347_),
    .A1(_21334_),
    .B1(_21348_),
    .X(_21349_));
 sg13g2_nor2b_1 _29911_ (.A(\u_inv.f_reg[95] ),
    .B_N(\u_inv.f_next[95] ),
    .Y(_21350_));
 sg13g2_nor2b_2 _29912_ (.A(\u_inv.f_reg[94] ),
    .B_N(\u_inv.f_next[94] ),
    .Y(_21351_));
 sg13g2_a221oi_1 _29913_ (.B2(_20696_),
    .C1(_21350_),
    .B1(_21351_),
    .A1(_21337_),
    .Y(_21352_),
    .A2(_21349_));
 sg13g2_nand2_1 _29914_ (.Y(_21353_),
    .A(_21339_),
    .B(_21352_));
 sg13g2_nor4_1 _29915_ (.A(_20732_),
    .B(_20735_),
    .C(_20740_),
    .D(_20743_),
    .Y(_21354_));
 sg13g2_nand2_1 _29916_ (.Y(_21355_),
    .A(_20748_),
    .B(_20751_));
 sg13g2_nor3_1 _29917_ (.A(_20755_),
    .B(_20758_),
    .C(_21355_),
    .Y(_21356_));
 sg13g2_nand2_1 _29918_ (.Y(_21357_),
    .A(_21354_),
    .B(_21356_));
 sg13g2_a21oi_2 _29919_ (.B1(_21357_),
    .Y(_21358_),
    .A2(_21352_),
    .A1(_21339_));
 sg13g2_a21o_1 _29920_ (.A2(_21352_),
    .A1(_21339_),
    .B1(_21357_),
    .X(_21359_));
 sg13g2_nand2b_1 _29921_ (.Y(_21360_),
    .B(\u_inv.f_next[103] ),
    .A_N(\u_inv.f_reg[103] ));
 sg13g2_nor2_1 _29922_ (.A(_18051_),
    .B(\u_inv.f_reg[102] ),
    .Y(_21361_));
 sg13g2_nand2b_1 _29923_ (.Y(_21362_),
    .B(\u_inv.f_next[96] ),
    .A_N(\u_inv.f_reg[96] ));
 sg13g2_nor2_1 _29924_ (.A(_20755_),
    .B(_21362_),
    .Y(_21363_));
 sg13g2_a21oi_1 _29925_ (.A1(\u_inv.f_next[97] ),
    .A2(_18215_),
    .Y(_21364_),
    .B1(_21363_));
 sg13g2_nor2b_1 _29926_ (.A(\u_inv.f_reg[98] ),
    .B_N(\u_inv.f_next[98] ),
    .Y(_21365_));
 sg13g2_a21oi_1 _29927_ (.A1(_20748_),
    .A2(_21365_),
    .Y(_21366_),
    .B1(_20747_));
 sg13g2_o21ai_1 _29928_ (.B1(_21366_),
    .Y(_21367_),
    .A1(_21355_),
    .A2(_21364_));
 sg13g2_nor2b_1 _29929_ (.A(\u_inv.f_reg[100] ),
    .B_N(\u_inv.f_next[100] ),
    .Y(_21368_));
 sg13g2_a21oi_1 _29930_ (.A1(_20736_),
    .A2(_21367_),
    .Y(_21369_),
    .B1(_21368_));
 sg13g2_nand2b_1 _29931_ (.Y(_21370_),
    .B(\u_inv.f_next[101] ),
    .A_N(\u_inv.f_reg[101] ));
 sg13g2_o21ai_1 _29932_ (.B1(_21370_),
    .Y(_21371_),
    .A1(_20732_),
    .A2(_21369_));
 sg13g2_a21oi_1 _29933_ (.A1(_20744_),
    .A2(_21371_),
    .Y(_21372_),
    .B1(_21361_));
 sg13g2_o21ai_1 _29934_ (.B1(_21360_),
    .Y(_21373_),
    .A1(_20740_),
    .A2(_21372_));
 sg13g2_inv_1 _29935_ (.Y(_21374_),
    .A(_21373_));
 sg13g2_nor2_1 _29936_ (.A(_21358_),
    .B(_21373_),
    .Y(_21375_));
 sg13g2_nor4_1 _29937_ (.A(_20791_),
    .B(_20793_),
    .C(_20795_),
    .D(_20797_),
    .Y(_21376_));
 sg13g2_nor2_1 _29938_ (.A(_20777_),
    .B(_20780_),
    .Y(_21377_));
 sg13g2_and4_1 _29939_ (.A(_20784_),
    .B(_20787_),
    .C(_21376_),
    .D(_21377_),
    .X(_21378_));
 sg13g2_inv_1 _29940_ (.Y(_21379_),
    .A(_21378_));
 sg13g2_a21oi_1 _29941_ (.A1(_21359_),
    .A2(_21374_),
    .Y(_21380_),
    .B1(_21379_));
 sg13g2_o21ai_1 _29942_ (.B1(_21378_),
    .Y(_21381_),
    .A1(_21358_),
    .A2(_21373_));
 sg13g2_nand2b_1 _29943_ (.Y(_21382_),
    .B(\u_inv.f_next[109] ),
    .A_N(\u_inv.f_reg[109] ));
 sg13g2_nor2b_1 _29944_ (.A(\u_inv.f_reg[108] ),
    .B_N(\u_inv.f_next[108] ),
    .Y(_21383_));
 sg13g2_nor2_1 _29945_ (.A(_18048_),
    .B(\u_inv.f_reg[106] ),
    .Y(_21384_));
 sg13g2_inv_1 _29946_ (.Y(_21385_),
    .A(_21384_));
 sg13g2_nand2b_1 _29947_ (.Y(_21386_),
    .B(\u_inv.f_next[104] ),
    .A_N(\u_inv.f_reg[104] ));
 sg13g2_nor2_1 _29948_ (.A(_20795_),
    .B(_21386_),
    .Y(_21387_));
 sg13g2_nor2_1 _29949_ (.A(_18049_),
    .B(\u_inv.f_reg[105] ),
    .Y(_21388_));
 sg13g2_o21ai_1 _29950_ (.B1(_20792_),
    .Y(_21389_),
    .A1(_21387_),
    .A2(_21388_));
 sg13g2_a21oi_1 _29951_ (.A1(_21385_),
    .A2(_21389_),
    .Y(_21390_),
    .B1(_20793_));
 sg13g2_a21oi_1 _29952_ (.A1(\u_inv.f_next[107] ),
    .A2(_18217_),
    .Y(_21391_),
    .B1(_21390_));
 sg13g2_nor2_1 _29953_ (.A(_20786_),
    .B(_21391_),
    .Y(_21392_));
 sg13g2_o21ai_1 _29954_ (.B1(_20784_),
    .Y(_21393_),
    .A1(_21383_),
    .A2(_21392_));
 sg13g2_nand2_1 _29955_ (.Y(_21394_),
    .A(_21382_),
    .B(_21393_));
 sg13g2_nor2_1 _29956_ (.A(_18045_),
    .B(\u_inv.f_reg[110] ),
    .Y(_21395_));
 sg13g2_a22oi_1 _29957_ (.Y(_21396_),
    .B1(_21395_),
    .B2(_20778_),
    .A2(_21394_),
    .A1(_21377_));
 sg13g2_o21ai_1 _29958_ (.B1(_21396_),
    .Y(_21397_),
    .A1(_18044_),
    .A2(\u_inv.f_reg[111] ));
 sg13g2_inv_1 _29959_ (.Y(_21398_),
    .A(_21397_));
 sg13g2_nand2_2 _29960_ (.Y(_21399_),
    .A(_21381_),
    .B(_21398_));
 sg13g2_or4_1 _29961_ (.A(_20240_),
    .B(_20242_),
    .C(_20245_),
    .D(_20247_),
    .X(_21400_));
 sg13g2_nand2_1 _29962_ (.Y(_21401_),
    .A(_20230_),
    .B(_20233_));
 sg13g2_nand4_1 _29963_ (.B(_20233_),
    .C(_20236_),
    .A(_20230_),
    .Y(_21402_),
    .D(_20237_));
 sg13g2_nor2_2 _29964_ (.A(_21400_),
    .B(_21402_),
    .Y(_21403_));
 sg13g2_nor2_1 _29965_ (.A(_20266_),
    .B(_20268_),
    .Y(_21404_));
 sg13g2_nand3_1 _29966_ (.B(_20814_),
    .C(_21404_),
    .A(_20813_),
    .Y(_21405_));
 sg13g2_nand2b_1 _29967_ (.Y(_21406_),
    .B(_20255_),
    .A_N(_20253_));
 sg13g2_nor4_1 _29968_ (.A(_20258_),
    .B(_20261_),
    .C(_21405_),
    .D(_21406_),
    .Y(_21407_));
 sg13g2_nand2_1 _29969_ (.Y(_21408_),
    .A(_21403_),
    .B(_21407_));
 sg13g2_a21oi_2 _29970_ (.B1(_21408_),
    .Y(_21409_),
    .A2(_21398_),
    .A1(_21381_));
 sg13g2_nor2_1 _29971_ (.A(_18041_),
    .B(\u_inv.f_reg[117] ),
    .Y(_21410_));
 sg13g2_nand2_1 _29972_ (.Y(_21411_),
    .A(\u_inv.f_next[117] ),
    .B(_18219_));
 sg13g2_nand2b_1 _29973_ (.Y(_21412_),
    .B(\u_inv.f_next[116] ),
    .A_N(\u_inv.f_reg[116] ));
 sg13g2_nor2b_1 _29974_ (.A(\u_inv.f_reg[115] ),
    .B_N(\u_inv.f_next[115] ),
    .Y(_21413_));
 sg13g2_nor2_1 _29975_ (.A(_18042_),
    .B(\u_inv.f_reg[114] ),
    .Y(_21414_));
 sg13g2_nor2b_1 _29976_ (.A(\u_inv.f_reg[112] ),
    .B_N(\u_inv.f_next[112] ),
    .Y(_21415_));
 sg13g2_nand2_1 _29977_ (.Y(_21416_),
    .A(_20813_),
    .B(_21415_));
 sg13g2_nand2b_1 _29978_ (.Y(_21417_),
    .B(\u_inv.f_next[113] ),
    .A_N(\u_inv.f_reg[113] ));
 sg13g2_nand2_1 _29979_ (.Y(_21418_),
    .A(_21416_),
    .B(_21417_));
 sg13g2_a221oi_1 _29980_ (.B2(_21404_),
    .C1(_21413_),
    .B1(_21418_),
    .A1(_20269_),
    .Y(_21419_),
    .A2(_21414_));
 sg13g2_o21ai_1 _29981_ (.B1(_21412_),
    .Y(_21420_),
    .A1(_20261_),
    .A2(_21419_));
 sg13g2_nand2b_1 _29982_ (.Y(_21421_),
    .B(_21420_),
    .A_N(_20258_));
 sg13g2_a21oi_1 _29983_ (.A1(_21411_),
    .A2(_21421_),
    .Y(_21422_),
    .B1(_21406_));
 sg13g2_nand2b_1 _29984_ (.Y(_21423_),
    .B(\u_inv.f_next[118] ),
    .A_N(\u_inv.f_reg[118] ));
 sg13g2_a21oi_1 _29985_ (.A1(\u_inv.f_next[119] ),
    .A2(_18220_),
    .Y(_21424_),
    .B1(_21422_));
 sg13g2_o21ai_1 _29986_ (.B1(_21424_),
    .Y(_21425_),
    .A1(_20253_),
    .A2(_21423_));
 sg13g2_inv_1 _29987_ (.Y(_21426_),
    .A(_21425_));
 sg13g2_nor2_1 _29988_ (.A(_18036_),
    .B(\u_inv.f_reg[124] ),
    .Y(_21427_));
 sg13g2_nor2_1 _29989_ (.A(_18034_),
    .B(\u_inv.f_reg[126] ),
    .Y(_21428_));
 sg13g2_nand2b_1 _29990_ (.Y(_21429_),
    .B(\u_inv.f_next[127] ),
    .A_N(\u_inv.f_reg[127] ));
 sg13g2_nor2_1 _29991_ (.A(_18035_),
    .B(\u_inv.f_reg[125] ),
    .Y(_21430_));
 sg13g2_a21oi_1 _29992_ (.A1(_20237_),
    .A2(_21427_),
    .Y(_21431_),
    .B1(_21430_));
 sg13g2_o21ai_1 _29993_ (.B1(_21429_),
    .Y(_21432_),
    .A1(_21401_),
    .A2(_21431_));
 sg13g2_nand2b_1 _29994_ (.Y(_21433_),
    .B(\u_inv.f_next[120] ),
    .A_N(\u_inv.f_reg[120] ));
 sg13g2_nand2_1 _29995_ (.Y(_21434_),
    .A(\u_inv.f_next[121] ),
    .B(_18221_));
 sg13g2_o21ai_1 _29996_ (.B1(_21434_),
    .Y(_21435_),
    .A1(_20240_),
    .A2(_21433_));
 sg13g2_nor2_1 _29997_ (.A(_18038_),
    .B(\u_inv.f_reg[122] ),
    .Y(_21436_));
 sg13g2_a21oi_1 _29998_ (.A1(_20246_),
    .A2(_21435_),
    .Y(_21437_),
    .B1(_21436_));
 sg13g2_nand2_1 _29999_ (.Y(_21438_),
    .A(\u_inv.f_next[123] ),
    .B(_18222_));
 sg13g2_o21ai_1 _30000_ (.B1(_21438_),
    .Y(_21439_),
    .A1(_20247_),
    .A2(_21437_));
 sg13g2_inv_1 _30001_ (.Y(_21440_),
    .A(_21439_));
 sg13g2_a221oi_1 _30002_ (.B2(_20230_),
    .C1(_21432_),
    .B1(_21428_),
    .A1(_21403_),
    .Y(_21441_),
    .A2(_21425_));
 sg13g2_o21ai_1 _30003_ (.B1(_21441_),
    .Y(_21442_),
    .A1(_21402_),
    .A2(_21440_));
 sg13g2_or2_1 _30004_ (.X(_21443_),
    .B(_21442_),
    .A(_21409_));
 sg13g2_nor4_2 _30005_ (.A(_20825_),
    .B(_20827_),
    .C(_20831_),
    .Y(_21444_),
    .D(_20833_));
 sg13g2_nand2b_1 _30006_ (.Y(_21445_),
    .B(_20838_),
    .A_N(_20821_));
 sg13g2_nor3_1 _30007_ (.A(_20823_),
    .B(_20840_),
    .C(_21445_),
    .Y(_21446_));
 sg13g2_and2_1 _30008_ (.A(_21444_),
    .B(_21446_),
    .X(_21447_));
 sg13g2_o21ai_1 _30009_ (.B1(_21447_),
    .Y(_21448_),
    .A1(_21409_),
    .A2(_21442_));
 sg13g2_nor2b_1 _30010_ (.A(\u_inv.f_reg[131] ),
    .B_N(\u_inv.f_next[131] ),
    .Y(_21449_));
 sg13g2_nand2b_1 _30011_ (.Y(_21450_),
    .B(\u_inv.f_next[130] ),
    .A_N(\u_inv.f_reg[130] ));
 sg13g2_nand2b_1 _30012_ (.Y(_21451_),
    .B(\u_inv.f_next[128] ),
    .A_N(\u_inv.f_reg[128] ));
 sg13g2_nor2_1 _30013_ (.A(_20821_),
    .B(_21451_),
    .Y(_21452_));
 sg13g2_nor2b_1 _30014_ (.A(\u_inv.f_reg[129] ),
    .B_N(\u_inv.f_next[129] ),
    .Y(_21453_));
 sg13g2_o21ai_1 _30015_ (.B1(_20838_),
    .Y(_21454_),
    .A1(_21452_),
    .A2(_21453_));
 sg13g2_a21oi_1 _30016_ (.A1(_21450_),
    .A2(_21454_),
    .Y(_21455_),
    .B1(_20840_));
 sg13g2_or2_1 _30017_ (.X(_21456_),
    .B(_21455_),
    .A(_21449_));
 sg13g2_inv_1 _30018_ (.Y(_21457_),
    .A(_21456_));
 sg13g2_nor2b_1 _30019_ (.A(\u_inv.f_reg[134] ),
    .B_N(\u_inv.f_next[134] ),
    .Y(_21458_));
 sg13g2_nand2b_1 _30020_ (.Y(_21459_),
    .B(\u_inv.f_next[133] ),
    .A_N(\u_inv.f_reg[133] ));
 sg13g2_nor2b_1 _30021_ (.A(\u_inv.f_reg[132] ),
    .B_N(\u_inv.f_next[132] ),
    .Y(_21460_));
 sg13g2_nand2_1 _30022_ (.Y(_21461_),
    .A(_20828_),
    .B(_21460_));
 sg13g2_a21oi_1 _30023_ (.A1(_21459_),
    .A2(_21461_),
    .Y(_21462_),
    .B1(_20831_));
 sg13g2_o21ai_1 _30024_ (.B1(_20834_),
    .Y(_21463_),
    .A1(_21458_),
    .A2(_21462_));
 sg13g2_o21ai_1 _30025_ (.B1(_21463_),
    .Y(_21464_),
    .A1(_18032_),
    .A2(\u_inv.f_reg[135] ));
 sg13g2_a21oi_2 _30026_ (.B1(_21464_),
    .Y(_21465_),
    .A2(_21456_),
    .A1(_21444_));
 sg13g2_nand2_1 _30027_ (.Y(_21466_),
    .A(_21448_),
    .B(_21465_));
 sg13g2_nand2_1 _30028_ (.Y(_21467_),
    .A(_20864_),
    .B(_20866_));
 sg13g2_nor3_1 _30029_ (.A(_20870_),
    .B(_20873_),
    .C(_21467_),
    .Y(_21468_));
 sg13g2_nor4_1 _30030_ (.A(_20859_),
    .B(_20862_),
    .C(_20877_),
    .D(_20878_),
    .Y(_21469_));
 sg13g2_nand2_1 _30031_ (.Y(_21470_),
    .A(_21468_),
    .B(_21469_));
 sg13g2_a21oi_1 _30032_ (.A1(_21448_),
    .A2(_21465_),
    .Y(_21471_),
    .B1(_21470_));
 sg13g2_a21o_2 _30033_ (.A2(_21465_),
    .A1(_21448_),
    .B1(_21470_),
    .X(_21472_));
 sg13g2_nor2b_1 _30034_ (.A(\u_inv.f_reg[136] ),
    .B_N(\u_inv.f_next[136] ),
    .Y(_21473_));
 sg13g2_nor2b_1 _30035_ (.A(\u_inv.f_reg[138] ),
    .B_N(\u_inv.f_next[138] ),
    .Y(_21474_));
 sg13g2_nand2b_1 _30036_ (.Y(_21475_),
    .B(\u_inv.f_next[137] ),
    .A_N(\u_inv.f_reg[137] ));
 sg13g2_nand2_1 _30037_ (.Y(_21476_),
    .A(_20860_),
    .B(_21473_));
 sg13g2_a21oi_1 _30038_ (.A1(_21475_),
    .A2(_21476_),
    .Y(_21477_),
    .B1(_20877_));
 sg13g2_o21ai_1 _30039_ (.B1(_20879_),
    .Y(_21478_),
    .A1(_21474_),
    .A2(_21477_));
 sg13g2_o21ai_1 _30040_ (.B1(_21478_),
    .Y(_21479_),
    .A1(_18030_),
    .A2(\u_inv.f_reg[139] ));
 sg13g2_nand2b_1 _30041_ (.Y(_21480_),
    .B(\u_inv.f_next[140] ),
    .A_N(\u_inv.f_reg[140] ));
 sg13g2_nor2_1 _30042_ (.A(_20863_),
    .B(_21480_),
    .Y(_21481_));
 sg13g2_a21oi_1 _30043_ (.A1(\u_inv.f_next[141] ),
    .A2(_18225_),
    .Y(_21482_),
    .B1(_21481_));
 sg13g2_nand2_1 _30044_ (.Y(_21483_),
    .A(\u_inv.f_next[142] ),
    .B(_18226_));
 sg13g2_o21ai_1 _30045_ (.B1(_21483_),
    .Y(_21484_),
    .A1(_20870_),
    .A2(_21482_));
 sg13g2_nor2b_1 _30046_ (.A(\u_inv.f_reg[143] ),
    .B_N(\u_inv.f_next[143] ),
    .Y(_21485_));
 sg13g2_a221oi_1 _30047_ (.B2(_20874_),
    .C1(_21485_),
    .B1(_21484_),
    .A1(_21468_),
    .Y(_21486_),
    .A2(_21479_));
 sg13g2_inv_1 _30048_ (.Y(_21487_),
    .A(_21486_));
 sg13g2_or4_1 _30049_ (.A(_20169_),
    .B(_20172_),
    .C(_20176_),
    .D(_20178_),
    .X(_21488_));
 sg13g2_nand2_1 _30050_ (.Y(_21489_),
    .A(_20163_),
    .B(_20165_));
 sg13g2_nor4_2 _30051_ (.A(_20156_),
    .B(_20158_),
    .C(_21488_),
    .Y(_21490_),
    .D(_21489_));
 sg13g2_nand3b_1 _30052_ (.B(_20899_),
    .C(_20195_),
    .Y(_21491_),
    .A_N(_20198_));
 sg13g2_nand2_1 _30053_ (.Y(_21492_),
    .A(_20190_),
    .B(_20192_));
 sg13g2_nor2_1 _30054_ (.A(_20182_),
    .B(_20185_),
    .Y(_21493_));
 sg13g2_nand2_1 _30055_ (.Y(_21494_),
    .A(_20183_),
    .B(_20186_));
 sg13g2_nor4_1 _30056_ (.A(_20897_),
    .B(_21491_),
    .C(_21492_),
    .D(_21494_),
    .Y(_21495_));
 sg13g2_nand2_1 _30057_ (.Y(_21496_),
    .A(_21490_),
    .B(_21495_));
 sg13g2_a21oi_2 _30058_ (.B1(_21496_),
    .Y(_21497_),
    .A2(_21486_),
    .A1(_21472_));
 sg13g2_nor2b_1 _30059_ (.A(\u_inv.f_reg[157] ),
    .B_N(\u_inv.f_next[157] ),
    .Y(_21498_));
 sg13g2_nand2b_1 _30060_ (.Y(_21499_),
    .B(\u_inv.f_next[156] ),
    .A_N(\u_inv.f_reg[156] ));
 sg13g2_nor2b_1 _30061_ (.A(\u_inv.f_reg[154] ),
    .B_N(\u_inv.f_next[154] ),
    .Y(_21500_));
 sg13g2_nor2_1 _30062_ (.A(_18023_),
    .B(\u_inv.f_reg[152] ),
    .Y(_21501_));
 sg13g2_nand2_1 _30063_ (.Y(_21502_),
    .A(_20170_),
    .B(_21501_));
 sg13g2_nand2b_1 _30064_ (.Y(_21503_),
    .B(\u_inv.f_next[153] ),
    .A_N(\u_inv.f_reg[153] ));
 sg13g2_a21oi_1 _30065_ (.A1(_21502_),
    .A2(_21503_),
    .Y(_21504_),
    .B1(_20176_));
 sg13g2_or2_1 _30066_ (.X(_21505_),
    .B(_21504_),
    .A(_21500_));
 sg13g2_nand2b_1 _30067_ (.Y(_21506_),
    .B(_21505_),
    .A_N(_20178_));
 sg13g2_o21ai_1 _30068_ (.B1(_21506_),
    .Y(_21507_),
    .A1(_18021_),
    .A2(\u_inv.f_reg[155] ));
 sg13g2_nand2_1 _30069_ (.Y(_21508_),
    .A(_20165_),
    .B(_21507_));
 sg13g2_nand2_1 _30070_ (.Y(_21509_),
    .A(_21499_),
    .B(_21508_));
 sg13g2_a21oi_1 _30071_ (.A1(_20163_),
    .A2(_21509_),
    .Y(_21510_),
    .B1(_21498_));
 sg13g2_nor3_1 _30072_ (.A(_20156_),
    .B(_20158_),
    .C(_21510_),
    .Y(_21511_));
 sg13g2_nor2_1 _30073_ (.A(_18025_),
    .B(\u_inv.f_reg[149] ),
    .Y(_21512_));
 sg13g2_nor2b_1 _30074_ (.A(\u_inv.f_reg[148] ),
    .B_N(\u_inv.f_next[148] ),
    .Y(_21513_));
 sg13g2_nand2b_1 _30075_ (.Y(_21514_),
    .B(\u_inv.f_next[145] ),
    .A_N(\u_inv.f_reg[145] ));
 sg13g2_nor2_1 _30076_ (.A(_18027_),
    .B(\u_inv.f_reg[144] ),
    .Y(_21515_));
 sg13g2_nand2_1 _30077_ (.Y(_21516_),
    .A(_20899_),
    .B(_21515_));
 sg13g2_nor2b_1 _30078_ (.A(\u_inv.f_reg[146] ),
    .B_N(\u_inv.f_next[146] ),
    .Y(_21517_));
 sg13g2_a21oi_1 _30079_ (.A1(_21514_),
    .A2(_21516_),
    .Y(_21518_),
    .B1(_20198_));
 sg13g2_o21ai_1 _30080_ (.B1(_20195_),
    .Y(_21519_),
    .A1(_21517_),
    .A2(_21518_));
 sg13g2_o21ai_1 _30081_ (.B1(_21519_),
    .Y(_21520_),
    .A1(_18026_),
    .A2(\u_inv.f_reg[147] ));
 sg13g2_a221oi_1 _30082_ (.B2(_21493_),
    .C1(_21512_),
    .B1(_21520_),
    .A1(_20183_),
    .Y(_21521_),
    .A2(_21513_));
 sg13g2_nor2_1 _30083_ (.A(_18024_),
    .B(\u_inv.f_reg[150] ),
    .Y(_21522_));
 sg13g2_nand2b_1 _30084_ (.Y(_21523_),
    .B(\u_inv.f_next[151] ),
    .A_N(\u_inv.f_reg[151] ));
 sg13g2_o21ai_1 _30085_ (.B1(_21523_),
    .Y(_21524_),
    .A1(_21492_),
    .A2(_21521_));
 sg13g2_a21oi_2 _30086_ (.B1(_21524_),
    .Y(_21525_),
    .A2(_21522_),
    .A1(_20190_));
 sg13g2_nor2b_1 _30087_ (.A(_21525_),
    .B_N(_21490_),
    .Y(_21526_));
 sg13g2_nand2b_1 _30088_ (.Y(_21527_),
    .B(\u_inv.f_next[158] ),
    .A_N(\u_inv.f_reg[158] ));
 sg13g2_nand2b_1 _30089_ (.Y(_21528_),
    .B(\u_inv.f_next[159] ),
    .A_N(\u_inv.f_reg[159] ));
 sg13g2_o21ai_1 _30090_ (.B1(_21528_),
    .Y(_21529_),
    .A1(_20156_),
    .A2(_21527_));
 sg13g2_or3_1 _30091_ (.A(_21511_),
    .B(_21526_),
    .C(_21529_),
    .X(_21530_));
 sg13g2_or2_1 _30092_ (.X(_21531_),
    .B(_21530_),
    .A(_21497_));
 sg13g2_nor2_1 _30093_ (.A(_20905_),
    .B(_20907_),
    .Y(_21532_));
 sg13g2_nor4_1 _30094_ (.A(_20135_),
    .B(_20138_),
    .C(_20905_),
    .D(_20907_),
    .Y(_21533_));
 sg13g2_nor2_1 _30095_ (.A(_20116_),
    .B(_20118_),
    .Y(_21534_));
 sg13g2_nand3_1 _30096_ (.B(_20130_),
    .C(_21534_),
    .A(_20128_),
    .Y(_21535_));
 sg13g2_nand2_1 _30097_ (.Y(_21536_),
    .A(_20088_),
    .B(_20090_));
 sg13g2_or3_1 _30098_ (.A(_20096_),
    .B(_20097_),
    .C(_21536_),
    .X(_21537_));
 sg13g2_nor2_1 _30099_ (.A(_20102_),
    .B(_20105_),
    .Y(_21538_));
 sg13g2_nor4_1 _30100_ (.A(_20102_),
    .B(_20105_),
    .C(_20109_),
    .D(_20111_),
    .Y(_21539_));
 sg13g2_nor2b_1 _30101_ (.A(_21537_),
    .B_N(_21539_),
    .Y(_21540_));
 sg13g2_nand2_1 _30102_ (.Y(_21541_),
    .A(_21533_),
    .B(_21540_));
 sg13g2_nor2_1 _30103_ (.A(_21535_),
    .B(_21541_),
    .Y(_21542_));
 sg13g2_o21ai_1 _30104_ (.B1(_21542_),
    .Y(_21543_),
    .A1(_21497_),
    .A2(_21530_));
 sg13g2_nor2_1 _30105_ (.A(_18018_),
    .B(\u_inv.f_reg[162] ),
    .Y(_21544_));
 sg13g2_nor2b_1 _30106_ (.A(\u_inv.f_reg[160] ),
    .B_N(\u_inv.f_next[160] ),
    .Y(_21545_));
 sg13g2_nor2_1 _30107_ (.A(_18019_),
    .B(\u_inv.f_reg[161] ),
    .Y(_21546_));
 sg13g2_a21oi_1 _30108_ (.A1(_20908_),
    .A2(_21545_),
    .Y(_21547_),
    .B1(_21546_));
 sg13g2_nor2_1 _30109_ (.A(_20135_),
    .B(_21547_),
    .Y(_21548_));
 sg13g2_nor2_1 _30110_ (.A(_21544_),
    .B(_21548_),
    .Y(_21549_));
 sg13g2_nor2_1 _30111_ (.A(_20138_),
    .B(_21549_),
    .Y(_21550_));
 sg13g2_a21oi_2 _30112_ (.B1(_21550_),
    .Y(_21551_),
    .A2(_18231_),
    .A1(\u_inv.f_next[163] ));
 sg13g2_nand2b_1 _30113_ (.Y(_21552_),
    .B(\u_inv.f_next[168] ),
    .A_N(\u_inv.f_reg[168] ));
 sg13g2_nand2b_1 _30114_ (.Y(_21553_),
    .B(\u_inv.f_next[169] ),
    .A_N(\u_inv.f_reg[169] ));
 sg13g2_o21ai_1 _30115_ (.B1(_21553_),
    .Y(_21554_),
    .A1(_20109_),
    .A2(_21552_));
 sg13g2_nor2b_1 _30116_ (.A(\u_inv.f_reg[170] ),
    .B_N(\u_inv.f_next[170] ),
    .Y(_21555_));
 sg13g2_a221oi_1 _30117_ (.B2(_20104_),
    .C1(_20103_),
    .B1(_21555_),
    .A1(_21538_),
    .Y(_21556_),
    .A2(_21554_));
 sg13g2_or2_1 _30118_ (.X(_21557_),
    .B(_21556_),
    .A(_21537_));
 sg13g2_nand2b_1 _30119_ (.Y(_21558_),
    .B(\u_inv.f_next[172] ),
    .A_N(\u_inv.f_reg[172] ));
 sg13g2_nor2_1 _30120_ (.A(_20097_),
    .B(_21558_),
    .Y(_21559_));
 sg13g2_a21oi_1 _30121_ (.A1(\u_inv.f_next[173] ),
    .A2(_18234_),
    .Y(_21560_),
    .B1(_21559_));
 sg13g2_inv_1 _30122_ (.Y(_21561_),
    .A(_21560_));
 sg13g2_or2_1 _30123_ (.X(_21562_),
    .B(_21560_),
    .A(_21536_));
 sg13g2_nand2b_1 _30124_ (.Y(_21563_),
    .B(\u_inv.f_next[174] ),
    .A_N(\u_inv.f_reg[174] ));
 sg13g2_nand2b_1 _30125_ (.Y(_21564_),
    .B(_20088_),
    .A_N(_21563_));
 sg13g2_nand2b_1 _30126_ (.Y(_21565_),
    .B(\u_inv.f_next[166] ),
    .A_N(\u_inv.f_reg[166] ));
 sg13g2_nand2b_1 _30127_ (.Y(_21566_),
    .B(\u_inv.f_next[164] ),
    .A_N(\u_inv.f_reg[164] ));
 sg13g2_nor2_1 _30128_ (.A(_18016_),
    .B(\u_inv.f_reg[165] ),
    .Y(_21567_));
 sg13g2_nand2b_1 _30129_ (.Y(_21568_),
    .B(\u_inv.f_next[165] ),
    .A_N(\u_inv.f_reg[165] ));
 sg13g2_o21ai_1 _30130_ (.B1(_21568_),
    .Y(_21569_),
    .A1(_20129_),
    .A2(_21566_));
 sg13g2_a22oi_1 _30131_ (.Y(_21570_),
    .B1(_21534_),
    .B2(_21569_),
    .A2(_18232_),
    .A1(\u_inv.f_next[167] ));
 sg13g2_o21ai_1 _30132_ (.B1(_21570_),
    .Y(_21571_),
    .A1(_20116_),
    .A2(_21565_));
 sg13g2_nor2_1 _30133_ (.A(_21535_),
    .B(_21551_),
    .Y(_21572_));
 sg13g2_o21ai_1 _30134_ (.B1(_21540_),
    .Y(_21573_),
    .A1(_21571_),
    .A2(_21572_));
 sg13g2_nand4_1 _30135_ (.B(_21562_),
    .C(_21564_),
    .A(_21557_),
    .Y(_21574_),
    .D(_21573_));
 sg13g2_a21oi_2 _30136_ (.B1(_21574_),
    .Y(_21575_),
    .A2(_18235_),
    .A1(\u_inv.f_next[175] ));
 sg13g2_nor2_1 _30137_ (.A(_20038_),
    .B(_20041_),
    .Y(_21576_));
 sg13g2_nand3_1 _30138_ (.B(_20035_),
    .C(_21576_),
    .A(_20033_),
    .Y(_21577_));
 sg13g2_inv_1 _30139_ (.Y(_21578_),
    .A(_21577_));
 sg13g2_nand2_1 _30140_ (.Y(_21579_),
    .A(_20018_),
    .B(_20022_));
 sg13g2_nor4_1 _30141_ (.A(_20026_),
    .B(_20029_),
    .C(_21577_),
    .D(_21579_),
    .Y(_21580_));
 sg13g2_nand2b_1 _30142_ (.Y(_21581_),
    .B(_20048_),
    .A_N(_20045_));
 sg13g2_nor3_1 _30143_ (.A(_20051_),
    .B(_20054_),
    .C(_21581_),
    .Y(_21582_));
 sg13g2_nand4_1 _30144_ (.B(_20061_),
    .C(_20914_),
    .A(_20059_),
    .Y(_21583_),
    .D(_20916_));
 sg13g2_nor4_1 _30145_ (.A(_20051_),
    .B(_20054_),
    .C(_21581_),
    .D(_21583_),
    .Y(_21584_));
 sg13g2_inv_1 _30146_ (.Y(_21585_),
    .A(_21584_));
 sg13g2_nand2_1 _30147_ (.Y(_21586_),
    .A(_21580_),
    .B(_21584_));
 sg13g2_a21oi_2 _30148_ (.B1(_21586_),
    .Y(_21587_),
    .A2(_21575_),
    .A1(_21543_));
 sg13g2_nor2b_1 _30149_ (.A(\u_inv.f_reg[178] ),
    .B_N(\u_inv.f_next[178] ),
    .Y(_21588_));
 sg13g2_nor2_1 _30150_ (.A(_18009_),
    .B(\u_inv.f_reg[176] ),
    .Y(_21589_));
 sg13g2_nand2_1 _30151_ (.Y(_21590_),
    .A(_20914_),
    .B(_21589_));
 sg13g2_nand2_1 _30152_ (.Y(_21591_),
    .A(\u_inv.f_next[177] ),
    .B(_18236_));
 sg13g2_a21oi_1 _30153_ (.A1(_21590_),
    .A2(_21591_),
    .Y(_21592_),
    .B1(_20058_));
 sg13g2_o21ai_1 _30154_ (.B1(_20061_),
    .Y(_21593_),
    .A1(_21588_),
    .A2(_21592_));
 sg13g2_o21ai_1 _30155_ (.B1(_21593_),
    .Y(_21594_),
    .A1(_18007_),
    .A2(\u_inv.f_reg[179] ));
 sg13g2_nand2b_1 _30156_ (.Y(_21595_),
    .B(\u_inv.f_next[180] ),
    .A_N(\u_inv.f_reg[180] ));
 sg13g2_nor2b_1 _30157_ (.A(\u_inv.f_reg[181] ),
    .B_N(\u_inv.f_next[181] ),
    .Y(_21596_));
 sg13g2_nand2b_1 _30158_ (.Y(_21597_),
    .B(\u_inv.f_next[182] ),
    .A_N(\u_inv.f_reg[182] ));
 sg13g2_nor2_1 _30159_ (.A(_20054_),
    .B(_21595_),
    .Y(_21598_));
 sg13g2_nor2_1 _30160_ (.A(_21596_),
    .B(_21598_),
    .Y(_21599_));
 sg13g2_nor2_1 _30161_ (.A(_21581_),
    .B(_21599_),
    .Y(_21600_));
 sg13g2_a221oi_1 _30162_ (.B2(_21594_),
    .C1(_21600_),
    .B1(_21582_),
    .A1(\u_inv.f_next[183] ),
    .Y(_21601_),
    .A2(_18238_));
 sg13g2_o21ai_1 _30163_ (.B1(_21601_),
    .Y(_21602_),
    .A1(_20045_),
    .A2(_21597_));
 sg13g2_nor2_1 _30164_ (.A(_18000_),
    .B(\u_inv.f_reg[188] ),
    .Y(_21603_));
 sg13g2_nand2_1 _30165_ (.Y(_21604_),
    .A(_20027_),
    .B(_21603_));
 sg13g2_nand2b_2 _30166_ (.Y(_21605_),
    .B(\u_inv.f_next[189] ),
    .A_N(\u_inv.f_reg[189] ));
 sg13g2_a21oi_1 _30167_ (.A1(_21604_),
    .A2(_21605_),
    .Y(_21606_),
    .B1(_21579_));
 sg13g2_nor2_1 _30168_ (.A(_17999_),
    .B(\u_inv.f_reg[190] ),
    .Y(_21607_));
 sg13g2_nand2_1 _30169_ (.Y(_21608_),
    .A(_20018_),
    .B(_21607_));
 sg13g2_a21oi_1 _30170_ (.A1(\u_inv.f_next[191] ),
    .A2(_18241_),
    .Y(_21609_),
    .B1(_21606_));
 sg13g2_nand2b_1 _30171_ (.Y(_21610_),
    .B(\u_inv.f_next[184] ),
    .A_N(\u_inv.f_reg[184] ));
 sg13g2_nor2_1 _30172_ (.A(_20032_),
    .B(_21610_),
    .Y(_21611_));
 sg13g2_nor2_1 _30173_ (.A(_18003_),
    .B(\u_inv.f_reg[185] ),
    .Y(_21612_));
 sg13g2_o21ai_1 _30174_ (.B1(_20039_),
    .Y(_21613_),
    .A1(_21611_),
    .A2(_21612_));
 sg13g2_nand2b_1 _30175_ (.Y(_21614_),
    .B(\u_inv.f_next[186] ),
    .A_N(\u_inv.f_reg[186] ));
 sg13g2_a21oi_1 _30176_ (.A1(_21613_),
    .A2(_21614_),
    .Y(_21615_),
    .B1(_20041_));
 sg13g2_a21oi_1 _30177_ (.A1(\u_inv.f_next[187] ),
    .A2(_18240_),
    .Y(_21616_),
    .B1(_21615_));
 sg13g2_nor4_1 _30178_ (.A(_20026_),
    .B(_20029_),
    .C(_21579_),
    .D(_21616_),
    .Y(_21617_));
 sg13g2_a21oi_1 _30179_ (.A1(_21580_),
    .A2(_21602_),
    .Y(_21618_),
    .B1(_21617_));
 sg13g2_nand3_1 _30180_ (.B(_21609_),
    .C(_21618_),
    .A(_21608_),
    .Y(_21619_));
 sg13g2_nor2_1 _30181_ (.A(_21587_),
    .B(_21619_),
    .Y(_21620_));
 sg13g2_nor2_1 _30182_ (.A(_19913_),
    .B(_19916_),
    .Y(_21621_));
 sg13g2_and3_1 _30183_ (.X(_21622_),
    .A(_19910_),
    .B(_19912_),
    .C(_21621_));
 sg13g2_nand4_1 _30184_ (.B(_19924_),
    .C(_19938_),
    .A(_19922_),
    .Y(_21623_),
    .D(_19940_));
 sg13g2_inv_1 _30185_ (.Y(_21624_),
    .A(_21623_));
 sg13g2_nand2_1 _30186_ (.Y(_21625_),
    .A(_21622_),
    .B(_21624_));
 sg13g2_nor2_1 _30187_ (.A(_19871_),
    .B(_19873_),
    .Y(_21626_));
 sg13g2_nand2_1 _30188_ (.Y(_21627_),
    .A(_19877_),
    .B(_19880_));
 sg13g2_nand3_1 _30189_ (.B(_19880_),
    .C(_21626_),
    .A(_19877_),
    .Y(_21628_));
 sg13g2_nor2_1 _30190_ (.A(_19884_),
    .B(_19887_),
    .Y(_21629_));
 sg13g2_and3_1 _30191_ (.X(_21630_),
    .A(_19902_),
    .B(_19903_),
    .C(_21629_));
 sg13g2_nor2b_1 _30192_ (.A(_21628_),
    .B_N(_21630_),
    .Y(_21631_));
 sg13g2_nor2b_2 _30193_ (.A(_21625_),
    .B_N(_21631_),
    .Y(_21632_));
 sg13g2_nand2_1 _30194_ (.Y(_21633_),
    .A(_19948_),
    .B(_19951_));
 sg13g2_nor2_1 _30195_ (.A(_19954_),
    .B(_19956_),
    .Y(_21634_));
 sg13g2_nor2b_1 _30196_ (.A(_21633_),
    .B_N(_21634_),
    .Y(_21635_));
 sg13g2_nand2_1 _30197_ (.Y(_21636_),
    .A(_19961_),
    .B(_19965_));
 sg13g2_nor2b_1 _30198_ (.A(_21636_),
    .B_N(_20007_),
    .Y(_21637_));
 sg13g2_nand2_1 _30199_ (.Y(_21638_),
    .A(_20009_),
    .B(_21637_));
 sg13g2_nand3_1 _30200_ (.B(_21635_),
    .C(_21637_),
    .A(_20009_),
    .Y(_21639_));
 sg13g2_nor2_1 _30201_ (.A(_20922_),
    .B(_20923_),
    .Y(_21640_));
 sg13g2_nand3_1 _30202_ (.B(_19990_),
    .C(_21640_),
    .A(_19989_),
    .Y(_21641_));
 sg13g2_inv_1 _30203_ (.Y(_21642_),
    .A(_21641_));
 sg13g2_nand2_1 _30204_ (.Y(_21643_),
    .A(_19979_),
    .B(_19981_));
 sg13g2_nor4_1 _30205_ (.A(_19983_),
    .B(_19985_),
    .C(_21641_),
    .D(_21643_),
    .Y(_21644_));
 sg13g2_nor2b_1 _30206_ (.A(_21639_),
    .B_N(_21644_),
    .Y(_21645_));
 sg13g2_nand2_1 _30207_ (.Y(_21646_),
    .A(_21632_),
    .B(_21645_));
 sg13g2_inv_1 _30208_ (.Y(_21647_),
    .A(_21646_));
 sg13g2_o21ai_1 _30209_ (.B1(_21647_),
    .Y(_21648_),
    .A1(_21587_),
    .A2(_21619_));
 sg13g2_nand2b_2 _30210_ (.Y(_21649_),
    .B(\u_inv.f_next[197] ),
    .A_N(\u_inv.f_reg[197] ));
 sg13g2_nor2_1 _30211_ (.A(_17994_),
    .B(\u_inv.f_reg[196] ),
    .Y(_21650_));
 sg13g2_nor2_1 _30212_ (.A(_17995_),
    .B(\u_inv.f_reg[195] ),
    .Y(_21651_));
 sg13g2_nand2b_1 _30213_ (.Y(_21652_),
    .B(\u_inv.f_next[194] ),
    .A_N(\u_inv.f_reg[194] ));
 sg13g2_nand2_1 _30214_ (.Y(_21653_),
    .A(\u_inv.f_next[192] ),
    .B(_18242_));
 sg13g2_nor2_1 _30215_ (.A(_20922_),
    .B(_21653_),
    .Y(_21654_));
 sg13g2_nor2_1 _30216_ (.A(_17996_),
    .B(\u_inv.f_reg[193] ),
    .Y(_21655_));
 sg13g2_o21ai_1 _30217_ (.B1(_19989_),
    .Y(_21656_),
    .A1(_21654_),
    .A2(_21655_));
 sg13g2_nand2_1 _30218_ (.Y(_21657_),
    .A(_21652_),
    .B(_21656_));
 sg13g2_a21oi_1 _30219_ (.A1(_19990_),
    .A2(_21657_),
    .Y(_21658_),
    .B1(_21651_));
 sg13g2_nor2_1 _30220_ (.A(_19985_),
    .B(_21658_),
    .Y(_21659_));
 sg13g2_o21ai_1 _30221_ (.B1(_19984_),
    .Y(_21660_),
    .A1(_21650_),
    .A2(_21659_));
 sg13g2_a21oi_1 _30222_ (.A1(_21649_),
    .A2(_21660_),
    .Y(_21661_),
    .B1(_21643_));
 sg13g2_nor2_1 _30223_ (.A(_17992_),
    .B(\u_inv.f_reg[198] ),
    .Y(_21662_));
 sg13g2_nor2b_1 _30224_ (.A(\u_inv.f_reg[199] ),
    .B_N(\u_inv.f_next[199] ),
    .Y(_21663_));
 sg13g2_a21oi_1 _30225_ (.A1(_19979_),
    .A2(_21662_),
    .Y(_21664_),
    .B1(_21663_));
 sg13g2_nor2b_2 _30226_ (.A(_21661_),
    .B_N(_21664_),
    .Y(_21665_));
 sg13g2_nor2b_1 _30227_ (.A(\u_inv.f_reg[200] ),
    .B_N(\u_inv.f_next[200] ),
    .Y(_21666_));
 sg13g2_nor2_1 _30228_ (.A(_17989_),
    .B(\u_inv.f_reg[203] ),
    .Y(_21667_));
 sg13g2_nor2_1 _30229_ (.A(_17990_),
    .B(\u_inv.f_reg[202] ),
    .Y(_21668_));
 sg13g2_a21oi_1 _30230_ (.A1(_19965_),
    .A2(_21668_),
    .Y(_21669_),
    .B1(_21667_));
 sg13g2_nor2_1 _30231_ (.A(_17991_),
    .B(\u_inv.f_reg[201] ),
    .Y(_21670_));
 sg13g2_a21oi_1 _30232_ (.A1(_20007_),
    .A2(_21666_),
    .Y(_21671_),
    .B1(_21670_));
 sg13g2_o21ai_1 _30233_ (.B1(_21669_),
    .Y(_21672_),
    .A1(_21636_),
    .A2(_21671_));
 sg13g2_nand2b_1 _30234_ (.Y(_21673_),
    .B(\u_inv.f_next[204] ),
    .A_N(\u_inv.f_reg[204] ));
 sg13g2_nor2_1 _30235_ (.A(_19956_),
    .B(_21673_),
    .Y(_21674_));
 sg13g2_or2_1 _30236_ (.X(_21675_),
    .B(_21673_),
    .A(_19956_));
 sg13g2_a21oi_1 _30237_ (.A1(\u_inv.f_next[205] ),
    .A2(_18246_),
    .Y(_21676_),
    .B1(_21674_));
 sg13g2_nor2_1 _30238_ (.A(_21633_),
    .B(_21676_),
    .Y(_21677_));
 sg13g2_nor2b_1 _30239_ (.A(\u_inv.f_reg[206] ),
    .B_N(\u_inv.f_next[206] ),
    .Y(_21678_));
 sg13g2_a221oi_1 _30240_ (.B2(_19948_),
    .C1(_21677_),
    .B1(_21678_),
    .A1(_21635_),
    .Y(_21679_),
    .A2(_21672_));
 sg13g2_o21ai_1 _30241_ (.B1(_21679_),
    .Y(_21680_),
    .A1(_21639_),
    .A2(_21665_));
 sg13g2_a21oi_2 _30242_ (.B1(_21680_),
    .Y(_21681_),
    .A2(_18247_),
    .A1(\u_inv.f_next[207] ));
 sg13g2_inv_1 _30243_ (.Y(_21682_),
    .A(_21681_));
 sg13g2_nand2_1 _30244_ (.Y(_21683_),
    .A(\u_inv.f_next[219] ),
    .B(_18249_));
 sg13g2_nand2b_1 _30245_ (.Y(_21684_),
    .B(\u_inv.f_next[218] ),
    .A_N(\u_inv.f_reg[218] ));
 sg13g2_nand2b_1 _30246_ (.Y(_21685_),
    .B(\u_inv.f_next[216] ),
    .A_N(\u_inv.f_reg[216] ));
 sg13g2_nor2_1 _30247_ (.A(_19901_),
    .B(_21685_),
    .Y(_21686_));
 sg13g2_nor2_1 _30248_ (.A(_17980_),
    .B(\u_inv.f_reg[217] ),
    .Y(_21687_));
 sg13g2_or2_1 _30249_ (.X(_21688_),
    .B(_21687_),
    .A(_21686_));
 sg13g2_o21ai_1 _30250_ (.B1(_21683_),
    .Y(_21689_),
    .A1(_19887_),
    .A2(_21684_));
 sg13g2_a21oi_2 _30251_ (.B1(_21689_),
    .Y(_21690_),
    .A2(_21688_),
    .A1(_21629_));
 sg13g2_nor2_1 _30252_ (.A(_17978_),
    .B(\u_inv.f_reg[220] ),
    .Y(_21691_));
 sg13g2_and2_1 _30253_ (.A(_19877_),
    .B(_21691_),
    .X(_21692_));
 sg13g2_nand2b_1 _30254_ (.Y(_21693_),
    .B(\u_inv.f_next[221] ),
    .A_N(\u_inv.f_reg[221] ));
 sg13g2_nand2b_1 _30255_ (.Y(_21694_),
    .B(_21693_),
    .A_N(_21692_));
 sg13g2_nand2b_1 _30256_ (.Y(_21695_),
    .B(\u_inv.f_next[223] ),
    .A_N(\u_inv.f_reg[223] ));
 sg13g2_nand2b_1 _30257_ (.Y(_21696_),
    .B(\u_inv.f_next[222] ),
    .A_N(\u_inv.f_reg[222] ));
 sg13g2_o21ai_1 _30258_ (.B1(_21695_),
    .Y(_21697_),
    .A1(_19871_),
    .A2(_21696_));
 sg13g2_a21oi_1 _30259_ (.A1(_21626_),
    .A2(_21694_),
    .Y(_21698_),
    .B1(_21697_));
 sg13g2_o21ai_1 _30260_ (.B1(_21698_),
    .Y(_21699_),
    .A1(_21628_),
    .A2(_21690_));
 sg13g2_nor2_1 _30261_ (.A(_17986_),
    .B(\u_inv.f_reg[208] ),
    .Y(_21700_));
 sg13g2_nand2_1 _30262_ (.Y(_21701_),
    .A(_19938_),
    .B(_21700_));
 sg13g2_nand2b_1 _30263_ (.Y(_21702_),
    .B(\u_inv.f_next[209] ),
    .A_N(\u_inv.f_reg[209] ));
 sg13g2_a21oi_1 _30264_ (.A1(_21701_),
    .A2(_21702_),
    .Y(_21703_),
    .B1(_19921_));
 sg13g2_nor2b_1 _30265_ (.A(\u_inv.f_reg[210] ),
    .B_N(\u_inv.f_next[210] ),
    .Y(_21704_));
 sg13g2_o21ai_1 _30266_ (.B1(_19924_),
    .Y(_21705_),
    .A1(_21703_),
    .A2(_21704_));
 sg13g2_o21ai_1 _30267_ (.B1(_21705_),
    .Y(_21706_),
    .A1(_17985_),
    .A2(\u_inv.f_reg[211] ));
 sg13g2_nand2b_1 _30268_ (.Y(_21707_),
    .B(\u_inv.f_next[212] ),
    .A_N(\u_inv.f_reg[212] ));
 sg13g2_nor2_1 _30269_ (.A(_19913_),
    .B(_21707_),
    .Y(_21708_));
 sg13g2_a21oi_1 _30270_ (.A1(\u_inv.f_next[213] ),
    .A2(_18248_),
    .Y(_21709_),
    .B1(_21708_));
 sg13g2_nor2b_1 _30271_ (.A(\u_inv.f_reg[214] ),
    .B_N(\u_inv.f_next[214] ),
    .Y(_21710_));
 sg13g2_inv_1 _30272_ (.Y(_21711_),
    .A(_21710_));
 sg13g2_o21ai_1 _30273_ (.B1(_21711_),
    .Y(_21712_),
    .A1(_19909_),
    .A2(_21709_));
 sg13g2_a22oi_1 _30274_ (.Y(_21713_),
    .B1(_21712_),
    .B2(_19912_),
    .A2(_21706_),
    .A1(_21622_));
 sg13g2_o21ai_1 _30275_ (.B1(_21713_),
    .Y(_21714_),
    .A1(_17982_),
    .A2(\u_inv.f_reg[215] ));
 sg13g2_a221oi_1 _30276_ (.B2(_21631_),
    .C1(_21699_),
    .B1(_21714_),
    .A1(_21632_),
    .Y(_21715_),
    .A2(_21682_));
 sg13g2_nand2_1 _30277_ (.Y(_21716_),
    .A(_20941_),
    .B(_20944_));
 sg13g2_nor3_1 _30278_ (.A(_20934_),
    .B(_20936_),
    .C(_21716_),
    .Y(_21717_));
 sg13g2_nor2_1 _30279_ (.A(_20948_),
    .B(_20950_),
    .Y(_21718_));
 sg13g2_nor2_1 _30280_ (.A(_20953_),
    .B(_20954_),
    .Y(_21719_));
 sg13g2_inv_1 _30281_ (.Y(_21720_),
    .A(_21719_));
 sg13g2_nand2_1 _30282_ (.Y(_21721_),
    .A(_21718_),
    .B(_21719_));
 sg13g2_nand3_1 _30283_ (.B(_21718_),
    .C(_21719_),
    .A(_21717_),
    .Y(_21722_));
 sg13g2_and2_1 _30284_ (.A(_20983_),
    .B(_20985_),
    .X(_21723_));
 sg13g2_nand3_1 _30285_ (.B(_20979_),
    .C(_21723_),
    .A(_20975_),
    .Y(_21724_));
 sg13g2_nor4_1 _30286_ (.A(_20961_),
    .B(_20965_),
    .C(_20968_),
    .D(_20970_),
    .Y(_21725_));
 sg13g2_nor2b_1 _30287_ (.A(_21724_),
    .B_N(_21725_),
    .Y(_21726_));
 sg13g2_nand2b_1 _30288_ (.Y(_21727_),
    .B(_21726_),
    .A_N(_21722_));
 sg13g2_a21oi_2 _30289_ (.B1(_21727_),
    .Y(_21728_),
    .A2(_21715_),
    .A1(_21648_));
 sg13g2_nand2b_1 _30290_ (.Y(_21729_),
    .B(\u_inv.f_next[227] ),
    .A_N(\u_inv.f_reg[227] ));
 sg13g2_nor2b_1 _30291_ (.A(\u_inv.f_reg[226] ),
    .B_N(\u_inv.f_next[226] ),
    .Y(_21730_));
 sg13g2_nor2b_1 _30292_ (.A(\u_inv.f_reg[224] ),
    .B_N(\u_inv.f_next[224] ),
    .Y(_21731_));
 sg13g2_nand2_1 _30293_ (.Y(_21732_),
    .A(_20955_),
    .B(_21731_));
 sg13g2_o21ai_1 _30294_ (.B1(_21732_),
    .Y(_21733_),
    .A1(_17976_),
    .A2(\u_inv.f_reg[225] ));
 sg13g2_nand2_1 _30295_ (.Y(_21734_),
    .A(_21718_),
    .B(_21733_));
 sg13g2_nand2b_1 _30296_ (.Y(_21735_),
    .B(_21730_),
    .A_N(_20948_));
 sg13g2_nand3_1 _30297_ (.B(_21734_),
    .C(_21735_),
    .A(_21729_),
    .Y(_21736_));
 sg13g2_nor2b_1 _30298_ (.A(\u_inv.f_reg[231] ),
    .B_N(\u_inv.f_next[231] ),
    .Y(_21737_));
 sg13g2_nor2b_1 _30299_ (.A(\u_inv.f_reg[230] ),
    .B_N(\u_inv.f_next[230] ),
    .Y(_21738_));
 sg13g2_nand2b_1 _30300_ (.Y(_21739_),
    .B(\u_inv.f_next[228] ),
    .A_N(\u_inv.f_reg[228] ));
 sg13g2_nor2_1 _30301_ (.A(_20934_),
    .B(_21739_),
    .Y(_21740_));
 sg13g2_a21oi_1 _30302_ (.A1(\u_inv.f_next[229] ),
    .A2(_18251_),
    .Y(_21741_),
    .B1(_21740_));
 sg13g2_a221oi_1 _30303_ (.B2(_20944_),
    .C1(_21737_),
    .B1(_21738_),
    .A1(_21717_),
    .Y(_21742_),
    .A2(_21736_));
 sg13g2_o21ai_1 _30304_ (.B1(_21742_),
    .Y(_21743_),
    .A1(_21716_),
    .A2(_21741_));
 sg13g2_nand2b_1 _30305_ (.Y(_21744_),
    .B(\u_inv.f_next[232] ),
    .A_N(\u_inv.f_reg[232] ));
 sg13g2_nand2b_1 _30306_ (.Y(_21745_),
    .B(\u_inv.f_next[234] ),
    .A_N(\u_inv.f_reg[234] ));
 sg13g2_nor2b_2 _30307_ (.A(\u_inv.f_reg[233] ),
    .B_N(\u_inv.f_next[233] ),
    .Y(_21746_));
 sg13g2_nor2_1 _30308_ (.A(_20965_),
    .B(_21744_),
    .Y(_21747_));
 sg13g2_o21ai_1 _30309_ (.B1(_20969_),
    .Y(_21748_),
    .A1(_21746_),
    .A2(_21747_));
 sg13g2_a21oi_1 _30310_ (.A1(_21745_),
    .A2(_21748_),
    .Y(_21749_),
    .B1(_20970_));
 sg13g2_a21oi_2 _30311_ (.B1(_21749_),
    .Y(_21750_),
    .A2(_18252_),
    .A1(\u_inv.f_next[235] ));
 sg13g2_nor2_1 _30312_ (.A(_17972_),
    .B(\u_inv.f_reg[236] ),
    .Y(_21751_));
 sg13g2_and2_1 _30313_ (.A(_20975_),
    .B(_21751_),
    .X(_21752_));
 sg13g2_nand2b_1 _30314_ (.Y(_21753_),
    .B(\u_inv.f_next[237] ),
    .A_N(\u_inv.f_reg[237] ));
 sg13g2_nand2b_1 _30315_ (.Y(_21754_),
    .B(_21753_),
    .A_N(_21752_));
 sg13g2_nand2b_1 _30316_ (.Y(_21755_),
    .B(\u_inv.f_next[239] ),
    .A_N(\u_inv.f_reg[239] ));
 sg13g2_nand2b_1 _30317_ (.Y(_21756_),
    .B(\u_inv.f_next[238] ),
    .A_N(\u_inv.f_reg[238] ));
 sg13g2_o21ai_1 _30318_ (.B1(_21755_),
    .Y(_21757_),
    .A1(_20982_),
    .A2(_21756_));
 sg13g2_a21oi_1 _30319_ (.A1(_21723_),
    .A2(_21754_),
    .Y(_21758_),
    .B1(_21757_));
 sg13g2_o21ai_1 _30320_ (.B1(_21758_),
    .Y(_21759_),
    .A1(_21724_),
    .A2(_21750_));
 sg13g2_a21o_2 _30321_ (.A2(_21743_),
    .A1(_21726_),
    .B1(_21759_),
    .X(_21760_));
 sg13g2_or2_1 _30322_ (.X(_21761_),
    .B(_21760_),
    .A(_21728_));
 sg13g2_nor2_1 _30323_ (.A(_21035_),
    .B(_21038_),
    .Y(_21762_));
 sg13g2_nand3_1 _30324_ (.B(_21032_),
    .C(_21762_),
    .A(_21028_),
    .Y(_21763_));
 sg13g2_and2_1 _30325_ (.A(_21043_),
    .B(_21044_),
    .X(_21764_));
 sg13g2_nor2_1 _30326_ (.A(_21019_),
    .B(_21023_),
    .Y(_21765_));
 sg13g2_and2_1 _30327_ (.A(_21764_),
    .B(_21765_),
    .X(_21766_));
 sg13g2_nor2b_1 _30328_ (.A(_21763_),
    .B_N(_21766_),
    .Y(_21767_));
 sg13g2_o21ai_1 _30329_ (.B1(_21767_),
    .Y(_21768_),
    .A1(_21728_),
    .A2(_21760_));
 sg13g2_nor2_1 _30330_ (.A(_17968_),
    .B(\u_inv.f_reg[243] ),
    .Y(_21769_));
 sg13g2_nor2_1 _30331_ (.A(_17969_),
    .B(\u_inv.f_reg[242] ),
    .Y(_21770_));
 sg13g2_nand2b_1 _30332_ (.Y(_21771_),
    .B(\u_inv.f_next[240] ),
    .A_N(\u_inv.f_reg[240] ));
 sg13g2_nand2b_1 _30333_ (.Y(_21772_),
    .B(\u_inv.f_next[241] ),
    .A_N(\u_inv.f_reg[241] ));
 sg13g2_o21ai_1 _30334_ (.B1(_21772_),
    .Y(_21773_),
    .A1(_21023_),
    .A2(_21771_));
 sg13g2_inv_1 _30335_ (.Y(_21774_),
    .A(_21773_));
 sg13g2_a221oi_1 _30336_ (.B2(_21764_),
    .C1(_21769_),
    .B1(_21773_),
    .A1(_21044_),
    .Y(_21775_),
    .A2(_21770_));
 sg13g2_nor2_1 _30337_ (.A(_21763_),
    .B(_21775_),
    .Y(_21776_));
 sg13g2_nor2b_1 _30338_ (.A(\u_inv.f_reg[246] ),
    .B_N(\u_inv.f_next[246] ),
    .Y(_21777_));
 sg13g2_nand2b_1 _30339_ (.Y(_21778_),
    .B(\u_inv.f_next[245] ),
    .A_N(\u_inv.f_reg[245] ));
 sg13g2_nor2_1 _30340_ (.A(_17967_),
    .B(\u_inv.f_reg[244] ),
    .Y(_21779_));
 sg13g2_nand2_1 _30341_ (.Y(_21780_),
    .A(_21028_),
    .B(_21779_));
 sg13g2_a21oi_1 _30342_ (.A1(_21778_),
    .A2(_21780_),
    .Y(_21781_),
    .B1(_21038_));
 sg13g2_o21ai_1 _30343_ (.B1(_21036_),
    .Y(_21782_),
    .A1(_21777_),
    .A2(_21781_));
 sg13g2_o21ai_1 _30344_ (.B1(_21782_),
    .Y(_21783_),
    .A1(_17966_),
    .A2(\u_inv.f_reg[247] ));
 sg13g2_or2_1 _30345_ (.X(_21784_),
    .B(_21783_),
    .A(_21776_));
 sg13g2_inv_1 _30346_ (.Y(_21785_),
    .A(_21784_));
 sg13g2_and2_1 _30347_ (.A(_21768_),
    .B(_21785_),
    .X(_21786_));
 sg13g2_and2_1 _30348_ (.A(_21064_),
    .B(_21065_),
    .X(_21787_));
 sg13g2_inv_1 _30349_ (.Y(_21788_),
    .A(_21787_));
 sg13g2_and3_1 _30350_ (.X(_21789_),
    .A(_19858_),
    .B(_19860_),
    .C(_21787_));
 sg13g2_inv_1 _30351_ (.Y(_21790_),
    .A(_21789_));
 sg13g2_a21oi_1 _30352_ (.A1(_21768_),
    .A2(_21785_),
    .Y(_21791_),
    .B1(_21790_));
 sg13g2_o21ai_1 _30353_ (.B1(_21081_),
    .Y(_21792_),
    .A1(_21088_),
    .A2(_21791_));
 sg13g2_a21oi_1 _30354_ (.A1(_21080_),
    .A2(_21792_),
    .Y(_21793_),
    .B1(_19846_));
 sg13g2_o21ai_1 _30355_ (.B1(_19844_),
    .Y(_21794_),
    .A1(_21075_),
    .A2(_21793_));
 sg13g2_nor3_1 _30356_ (.A(_19844_),
    .B(_21075_),
    .C(_21793_),
    .Y(_21795_));
 sg13g2_nor2_1 _30357_ (.A(net6202),
    .B(_21795_),
    .Y(_21796_));
 sg13g2_a22oi_1 _30358_ (.Y(_21797_),
    .B1(_21794_),
    .B2(_21796_),
    .A2(_21074_),
    .A1(_21073_));
 sg13g2_o21ai_1 _30359_ (.B1(_21024_),
    .Y(_21798_),
    .A1(_20991_),
    .A2(_21016_));
 sg13g2_o21ai_1 _30360_ (.B1(_21046_),
    .Y(_21799_),
    .A1(_20991_),
    .A2(_21016_));
 sg13g2_a21oi_1 _30361_ (.A1(_21059_),
    .A2(_21799_),
    .Y(_21800_),
    .B1(_21033_));
 sg13g2_o21ai_1 _30362_ (.B1(_21038_),
    .Y(_21801_),
    .A1(_21053_),
    .A2(_21800_));
 sg13g2_a21oi_1 _30363_ (.A1(_21037_),
    .A2(_21801_),
    .Y(_21802_),
    .B1(_21035_));
 sg13g2_nand3_1 _30364_ (.B(_21037_),
    .C(_21801_),
    .A(_21035_),
    .Y(_21803_));
 sg13g2_nor2_1 _30365_ (.A(net7181),
    .B(_21802_),
    .Y(_21804_));
 sg13g2_a221oi_1 _30366_ (.B2(_21804_),
    .C1(net6280),
    .B1(_21803_),
    .A1(_17966_),
    .Y(_21805_),
    .A2(net7181));
 sg13g2_o21ai_1 _30367_ (.B1(_21766_),
    .Y(_21806_),
    .A1(_21728_),
    .A2(_21760_));
 sg13g2_a21oi_1 _30368_ (.A1(_21775_),
    .A2(_21806_),
    .Y(_21807_),
    .B1(_21031_));
 sg13g2_o21ai_1 _30369_ (.B1(_21028_),
    .Y(_21808_),
    .A1(_21779_),
    .A2(_21807_));
 sg13g2_a21oi_1 _30370_ (.A1(_21778_),
    .A2(_21808_),
    .Y(_21809_),
    .B1(_21038_));
 sg13g2_nor2_1 _30371_ (.A(_21777_),
    .B(_21809_),
    .Y(_21810_));
 sg13g2_xnor2_1 _30372_ (.Y(_21811_),
    .A(_21036_),
    .B(_21810_));
 sg13g2_a21oi_1 _30373_ (.A1(net6281),
    .A2(_21811_),
    .Y(_21812_),
    .B1(_21805_));
 sg13g2_a21o_1 _30374_ (.A2(_21811_),
    .A1(net6280),
    .B1(_21805_),
    .X(_21813_));
 sg13g2_a21o_2 _30375_ (.A2(_20928_),
    .A1(_20016_),
    .B1(_19945_),
    .X(_21814_));
 sg13g2_and2_1 _30376_ (.A(_19937_),
    .B(_21814_),
    .X(_21815_));
 sg13g2_o21ai_1 _30377_ (.B1(_19891_),
    .Y(_21816_),
    .A1(_19905_),
    .A2(_21815_));
 sg13g2_nand2_1 _30378_ (.Y(_21817_),
    .A(_19884_),
    .B(_21816_));
 sg13g2_nand3_1 _30379_ (.B(_19887_),
    .C(_21817_),
    .A(_19883_),
    .Y(_21818_));
 sg13g2_a21o_1 _30380_ (.A2(_21817_),
    .A1(_19883_),
    .B1(_19887_),
    .X(_21819_));
 sg13g2_nand3_1 _30381_ (.B(_21818_),
    .C(_21819_),
    .A(net7306),
    .Y(_21820_));
 sg13g2_a21oi_1 _30382_ (.A1(_17979_),
    .A2(net7178),
    .Y(_21821_),
    .B1(net6277));
 sg13g2_o21ai_1 _30383_ (.B1(_21645_),
    .Y(_21822_),
    .A1(_21587_),
    .A2(_21619_));
 sg13g2_a21oi_1 _30384_ (.A1(_21681_),
    .A2(_21822_),
    .Y(_21823_),
    .B1(_21625_));
 sg13g2_o21ai_1 _30385_ (.B1(_19903_),
    .Y(_21824_),
    .A1(_21714_),
    .A2(_21823_));
 sg13g2_a21oi_1 _30386_ (.A1(_21685_),
    .A2(_21824_),
    .Y(_21825_),
    .B1(_19901_));
 sg13g2_o21ai_1 _30387_ (.B1(_19885_),
    .Y(_21826_),
    .A1(_21687_),
    .A2(_21825_));
 sg13g2_a21oi_1 _30388_ (.A1(_21684_),
    .A2(_21826_),
    .Y(_21827_),
    .B1(_19887_));
 sg13g2_nand3_1 _30389_ (.B(_21684_),
    .C(_21826_),
    .A(_19887_),
    .Y(_21828_));
 sg13g2_nor2_1 _30390_ (.A(net6196),
    .B(_21827_),
    .Y(_21829_));
 sg13g2_a22oi_1 _30391_ (.Y(_21830_),
    .B1(_21828_),
    .B2(_21829_),
    .A2(_21821_),
    .A1(_21820_));
 sg13g2_inv_1 _30392_ (.Y(_21831_),
    .A(_21830_));
 sg13g2_o21ai_1 _30393_ (.B1(_21066_),
    .Y(_21832_),
    .A1(_21049_),
    .A2(_21061_));
 sg13g2_a21o_1 _30394_ (.A2(_21832_),
    .A1(_19865_),
    .B1(_19860_),
    .X(_21833_));
 sg13g2_nand3_1 _30395_ (.B(_19859_),
    .C(_21833_),
    .A(_19857_),
    .Y(_21834_));
 sg13g2_a21o_1 _30396_ (.A2(_21833_),
    .A1(_19859_),
    .B1(_19857_),
    .X(_21835_));
 sg13g2_nand3_1 _30397_ (.B(_21834_),
    .C(_21835_),
    .A(net7312),
    .Y(_21836_));
 sg13g2_a21oi_1 _30398_ (.A1(_17963_),
    .A2(net7181),
    .Y(_21837_),
    .B1(net6280));
 sg13g2_a21oi_1 _30399_ (.A1(_21768_),
    .A2(_21785_),
    .Y(_21838_),
    .B1(_21788_));
 sg13g2_o21ai_1 _30400_ (.B1(_19860_),
    .Y(_21839_),
    .A1(_21085_),
    .A2(_21838_));
 sg13g2_a21oi_1 _30401_ (.A1(_21082_),
    .A2(_21839_),
    .Y(_21840_),
    .B1(_19857_));
 sg13g2_nand3_1 _30402_ (.B(_21082_),
    .C(_21839_),
    .A(_19857_),
    .Y(_21841_));
 sg13g2_nor2_1 _30403_ (.A(net6202),
    .B(_21840_),
    .Y(_21842_));
 sg13g2_a22oi_1 _30404_ (.Y(_21843_),
    .B1(_21841_),
    .B2(_21842_),
    .A2(_21837_),
    .A1(_21836_));
 sg13g2_a21oi_1 _30405_ (.A1(_21648_),
    .A2(_21715_),
    .Y(_21844_),
    .B1(_21722_));
 sg13g2_o21ai_1 _30406_ (.B1(_20962_),
    .Y(_21845_),
    .A1(_21743_),
    .A2(_21844_));
 sg13g2_a21oi_1 _30407_ (.A1(_21744_),
    .A2(_21845_),
    .Y(_21846_),
    .B1(_20965_));
 sg13g2_o21ai_1 _30408_ (.B1(_20969_),
    .Y(_21847_),
    .A1(_21746_),
    .A2(_21846_));
 sg13g2_a21oi_1 _30409_ (.A1(_21745_),
    .A2(_21847_),
    .Y(_21848_),
    .B1(_20970_));
 sg13g2_nand3_1 _30410_ (.B(_21745_),
    .C(_21847_),
    .A(_20970_),
    .Y(_21849_));
 sg13g2_nor2_1 _30411_ (.A(net6199),
    .B(_21848_),
    .Y(_21850_));
 sg13g2_nand2_1 _30412_ (.Y(_21851_),
    .A(_21849_),
    .B(_21850_));
 sg13g2_a21oi_1 _30413_ (.A1(_20930_),
    .A2(_20932_),
    .Y(_21852_),
    .B1(_20959_));
 sg13g2_a21o_1 _30414_ (.A2(_20932_),
    .A1(_20930_),
    .B1(_20959_),
    .X(_21853_));
 sg13g2_o21ai_1 _30415_ (.B1(_20966_),
    .Y(_21854_),
    .A1(_21002_),
    .A2(_21852_));
 sg13g2_a21oi_1 _30416_ (.A1(_21007_),
    .A2(_21854_),
    .Y(_21855_),
    .B1(_20969_));
 sg13g2_a21oi_1 _30417_ (.A1(\u_inv.f_next[234] ),
    .A2(\u_inv.f_reg[234] ),
    .Y(_21856_),
    .B1(_21855_));
 sg13g2_o21ai_1 _30418_ (.B1(net7309),
    .Y(_21857_),
    .A1(_20970_),
    .A2(_21856_));
 sg13g2_a21o_1 _30419_ (.A2(_21856_),
    .A1(_20970_),
    .B1(_21857_),
    .X(_21858_));
 sg13g2_nor2_1 _30420_ (.A(\u_inv.f_next[235] ),
    .B(net7309),
    .Y(_21859_));
 sg13g2_nor2_1 _30421_ (.A(net6279),
    .B(_21859_),
    .Y(_21860_));
 sg13g2_nand2_1 _30422_ (.Y(_21861_),
    .A(net6199),
    .B(_21858_));
 sg13g2_a22oi_1 _30423_ (.Y(_21862_),
    .B1(_21858_),
    .B2(_21860_),
    .A2(_21850_),
    .A1(_21849_));
 sg13g2_o21ai_1 _30424_ (.B1(_21851_),
    .Y(_21863_),
    .A1(_21859_),
    .A2(_21861_));
 sg13g2_a21oi_1 _30425_ (.A1(_21003_),
    .A2(_21853_),
    .Y(_21864_),
    .B1(_20988_));
 sg13g2_a21o_1 _30426_ (.A2(_21853_),
    .A1(_21003_),
    .B1(_20988_),
    .X(_21865_));
 sg13g2_o21ai_1 _30427_ (.B1(_20980_),
    .Y(_21866_),
    .A1(_21014_),
    .A2(_21864_));
 sg13g2_a21o_1 _30428_ (.A2(_21866_),
    .A1(_21009_),
    .B1(_20985_),
    .X(_21867_));
 sg13g2_a21o_1 _30429_ (.A2(_21867_),
    .A1(_20984_),
    .B1(_20982_),
    .X(_21868_));
 sg13g2_nand3_1 _30430_ (.B(_20984_),
    .C(_21867_),
    .A(_20982_),
    .Y(_21869_));
 sg13g2_and3_1 _30431_ (.X(_21870_),
    .A(net7309),
    .B(_21868_),
    .C(_21869_));
 sg13g2_o21ai_1 _30432_ (.B1(net6199),
    .Y(_21871_),
    .A1(\u_inv.f_next[239] ),
    .A2(net7309));
 sg13g2_nor2_1 _30433_ (.A(_21870_),
    .B(_21871_),
    .Y(_21872_));
 sg13g2_o21ai_1 _30434_ (.B1(_21725_),
    .Y(_21873_),
    .A1(_21743_),
    .A2(_21844_));
 sg13g2_a21oi_1 _30435_ (.A1(_21750_),
    .A2(_21873_),
    .Y(_21874_),
    .B1(_20978_));
 sg13g2_a221oi_1 _30436_ (.B2(_21873_),
    .C1(_20978_),
    .B1(_21750_),
    .A1(_20972_),
    .Y(_21875_),
    .A2(_20974_));
 sg13g2_o21ai_1 _30437_ (.B1(_20985_),
    .Y(_21876_),
    .A1(_21754_),
    .A2(_21875_));
 sg13g2_a21o_1 _30438_ (.A2(_21876_),
    .A1(_21756_),
    .B1(_20982_),
    .X(_21877_));
 sg13g2_nand3_1 _30439_ (.B(_21756_),
    .C(_21876_),
    .A(_20982_),
    .Y(_21878_));
 sg13g2_nand3_1 _30440_ (.B(_21877_),
    .C(_21878_),
    .A(net6279),
    .Y(_21879_));
 sg13g2_nor2b_1 _30441_ (.A(_21872_),
    .B_N(_21879_),
    .Y(_21880_));
 sg13g2_o21ai_1 _30442_ (.B1(_21879_),
    .Y(_21881_),
    .A1(_21870_),
    .A2(_21871_));
 sg13g2_nand2_1 _30443_ (.Y(_21882_),
    .A(\u_inv.f_next[256] ),
    .B(net7181));
 sg13g2_nor2_1 _30444_ (.A(\u_inv.f_next[256] ),
    .B(net7254),
    .Y(_21883_));
 sg13g2_xnor2_1 _30445_ (.Y(_21884_),
    .A(\u_inv.f_next[256] ),
    .B(net7254));
 sg13g2_nand2_1 _30446_ (.Y(_21885_),
    .A(_19843_),
    .B(_19846_));
 sg13g2_o21ai_1 _30447_ (.B1(_19845_),
    .Y(_21886_),
    .A1(\u_inv.f_next[255] ),
    .A2(\u_inv.f_reg[255] ));
 sg13g2_o21ai_1 _30448_ (.B1(_21886_),
    .Y(_21887_),
    .A1(_19851_),
    .A2(_21885_));
 sg13g2_a21oi_1 _30449_ (.A1(\u_inv.f_next[255] ),
    .A2(\u_inv.f_reg[255] ),
    .Y(_21888_),
    .B1(_21887_));
 sg13g2_nand3_1 _30450_ (.B(_19846_),
    .C(_19856_),
    .A(_19843_),
    .Y(_21889_));
 sg13g2_nor2_1 _30451_ (.A(_21067_),
    .B(_21889_),
    .Y(_21890_));
 sg13g2_and2_1 _30452_ (.A(_21061_),
    .B(_21890_),
    .X(_21891_));
 sg13g2_o21ai_1 _30453_ (.B1(_21888_),
    .Y(_21892_),
    .A1(_19868_),
    .A2(_21889_));
 sg13g2_nand2_1 _30454_ (.Y(_21893_),
    .A(_21047_),
    .B(_21890_));
 sg13g2_a21oi_1 _30455_ (.A1(_20992_),
    .A2(_21017_),
    .Y(_21894_),
    .B1(_21893_));
 sg13g2_nor3_1 _30456_ (.A(_21891_),
    .B(_21892_),
    .C(_21894_),
    .Y(_21895_));
 sg13g2_o21ai_1 _30457_ (.B1(net7312),
    .Y(_21896_),
    .A1(_21884_),
    .A2(_21895_));
 sg13g2_o21ai_1 _30458_ (.B1(_21882_),
    .Y(_21897_),
    .A1(_21883_),
    .A2(_21896_));
 sg13g2_and2_1 _30459_ (.A(net6202),
    .B(_21897_),
    .X(_21898_));
 sg13g2_nor4_1 _30460_ (.A(_19843_),
    .B(_19846_),
    .C(_19852_),
    .D(_19854_),
    .Y(_21899_));
 sg13g2_nand2_1 _30461_ (.Y(_21900_),
    .A(_21789_),
    .B(_21899_));
 sg13g2_nor2_1 _30462_ (.A(_17961_),
    .B(\u_inv.f_reg[255] ),
    .Y(_21901_));
 sg13g2_o21ai_1 _30463_ (.B1(_21076_),
    .Y(_21902_),
    .A1(_19846_),
    .A2(_21080_));
 sg13g2_a221oi_1 _30464_ (.B2(_19844_),
    .C1(_21901_),
    .B1(_21902_),
    .A1(_21088_),
    .Y(_21903_),
    .A2(_21899_));
 sg13g2_o21ai_1 _30465_ (.B1(_21903_),
    .Y(_21904_),
    .A1(_21786_),
    .A2(_21900_));
 sg13g2_a21oi_1 _30466_ (.A1(_21884_),
    .A2(_21904_),
    .Y(_21905_),
    .B1(net6202));
 sg13g2_nand2b_1 _30467_ (.Y(_21906_),
    .B(net7254),
    .A_N(\u_inv.f_next[256] ));
 sg13g2_a21o_2 _30468_ (.A2(_21906_),
    .A1(_21905_),
    .B1(_21898_),
    .X(_21907_));
 sg13g2_and2_1 _30469_ (.A(_21884_),
    .B(_21895_),
    .X(_21908_));
 sg13g2_o21ai_1 _30470_ (.B1(_21882_),
    .Y(_21909_),
    .A1(_21896_),
    .A2(_21908_));
 sg13g2_or2_1 _30471_ (.X(_21910_),
    .B(_21904_),
    .A(_21884_));
 sg13g2_a22oi_1 _30472_ (.Y(_21911_),
    .B1(_21910_),
    .B2(_21905_),
    .A2(_21909_),
    .A1(net6202));
 sg13g2_o21ai_1 _30473_ (.B1(_21644_),
    .Y(_21912_),
    .A1(_21587_),
    .A2(_21619_));
 sg13g2_a21oi_1 _30474_ (.A1(_21665_),
    .A2(_21912_),
    .Y(_21913_),
    .B1(_20008_));
 sg13g2_a21oi_1 _30475_ (.A1(_21665_),
    .A2(_21912_),
    .Y(_21914_),
    .B1(_21638_));
 sg13g2_o21ai_1 _30476_ (.B1(_19955_),
    .Y(_21915_),
    .A1(_21672_),
    .A2(_21914_));
 sg13g2_o21ai_1 _30477_ (.B1(_21634_),
    .Y(_21916_),
    .A1(_21672_),
    .A2(_21914_));
 sg13g2_a21oi_1 _30478_ (.A1(_21676_),
    .A2(_21916_),
    .Y(_21917_),
    .B1(_19950_));
 sg13g2_o21ai_1 _30479_ (.B1(_19948_),
    .Y(_21918_),
    .A1(_21678_),
    .A2(_21917_));
 sg13g2_nor3_1 _30480_ (.A(_19948_),
    .B(_21678_),
    .C(_21917_),
    .Y(_21919_));
 sg13g2_nor2_1 _30481_ (.A(net6193),
    .B(_21919_),
    .Y(_21920_));
 sg13g2_o21ai_1 _30482_ (.B1(_20926_),
    .Y(_21921_),
    .A1(_20085_),
    .A2(_20920_));
 sg13g2_a21oi_1 _30483_ (.A1(_20006_),
    .A2(_21921_),
    .Y(_21922_),
    .B1(_20009_));
 sg13g2_a21oi_1 _30484_ (.A1(_20006_),
    .A2(_21921_),
    .Y(_21923_),
    .B1(_20010_));
 sg13g2_a21oi_1 _30485_ (.A1(_20006_),
    .A2(_21921_),
    .Y(_21924_),
    .B1(_20012_));
 sg13g2_o21ai_1 _30486_ (.B1(_19957_),
    .Y(_21925_),
    .A1(_19972_),
    .A2(_21924_));
 sg13g2_a21oi_1 _30487_ (.A1(_19975_),
    .A2(_21925_),
    .Y(_21926_),
    .B1(_19951_));
 sg13g2_o21ai_1 _30488_ (.B1(_19948_),
    .Y(_21927_),
    .A1(_19949_),
    .A2(_21926_));
 sg13g2_or3_1 _30489_ (.A(_19948_),
    .B(_19949_),
    .C(_21926_),
    .X(_21928_));
 sg13g2_nand3_1 _30490_ (.B(_21927_),
    .C(_21928_),
    .A(net7303),
    .Y(_21929_));
 sg13g2_a21oi_1 _30491_ (.A1(_17987_),
    .A2(net7179),
    .Y(_21930_),
    .B1(net6275));
 sg13g2_and2_1 _30492_ (.A(_21929_),
    .B(_21930_),
    .X(_21931_));
 sg13g2_a22oi_1 _30493_ (.Y(_21932_),
    .B1(_21929_),
    .B2(_21930_),
    .A2(_21920_),
    .A1(_21918_));
 sg13g2_a21o_1 _30494_ (.A2(_21920_),
    .A1(_21918_),
    .B1(_21931_),
    .X(_21933_));
 sg13g2_a21oi_1 _30495_ (.A1(_21013_),
    .A2(_21865_),
    .Y(_21934_),
    .B1(_20979_));
 sg13g2_nor3_1 _30496_ (.A(_20978_),
    .B(_21014_),
    .C(_21864_),
    .Y(_21935_));
 sg13g2_o21ai_1 _30497_ (.B1(net7309),
    .Y(_21936_),
    .A1(_21934_),
    .A2(_21935_));
 sg13g2_o21ai_1 _30498_ (.B1(_21936_),
    .Y(_21937_),
    .A1(\u_inv.f_next[236] ),
    .A2(net7310));
 sg13g2_nand3_1 _30499_ (.B(_21750_),
    .C(_21873_),
    .A(_20978_),
    .Y(_21938_));
 sg13g2_nand3b_1 _30500_ (.B(_21938_),
    .C(net6279),
    .Y(_21939_),
    .A_N(_21874_));
 sg13g2_o21ai_1 _30501_ (.B1(_21939_),
    .Y(_21940_),
    .A1(net6279),
    .A2(_21937_));
 sg13g2_a21oi_1 _30502_ (.A1(_21052_),
    .A2(_21798_),
    .Y(_21941_),
    .B1(_21043_));
 sg13g2_and3_1 _30503_ (.X(_21942_),
    .A(_21043_),
    .B(_21052_),
    .C(_21798_));
 sg13g2_o21ai_1 _30504_ (.B1(net7310),
    .Y(_21943_),
    .A1(_21941_),
    .A2(_21942_));
 sg13g2_a21oi_1 _30505_ (.A1(_17969_),
    .A2(net7182),
    .Y(_21944_),
    .B1(net6279));
 sg13g2_nand2_1 _30506_ (.Y(_21945_),
    .A(_21943_),
    .B(_21944_));
 sg13g2_nand2_1 _30507_ (.Y(_21946_),
    .A(_21020_),
    .B(_21761_));
 sg13g2_o21ai_1 _30508_ (.B1(_21765_),
    .Y(_21947_),
    .A1(_21728_),
    .A2(_21760_));
 sg13g2_nand3_1 _30509_ (.B(_21774_),
    .C(_21947_),
    .A(_21042_),
    .Y(_21948_));
 sg13g2_a21oi_1 _30510_ (.A1(_21774_),
    .A2(_21947_),
    .Y(_21949_),
    .B1(_21042_));
 sg13g2_nor2_1 _30511_ (.A(net6200),
    .B(_21949_),
    .Y(_21950_));
 sg13g2_nand2_1 _30512_ (.Y(_21951_),
    .A(_21948_),
    .B(_21950_));
 sg13g2_a22oi_1 _30513_ (.Y(_21952_),
    .B1(_21948_),
    .B2(_21950_),
    .A2(_21944_),
    .A1(_21943_));
 sg13g2_nand2_1 _30514_ (.Y(_21953_),
    .A(_21945_),
    .B(_21951_));
 sg13g2_nand3_1 _30515_ (.B(_21676_),
    .C(_21916_),
    .A(_19950_),
    .Y(_21954_));
 sg13g2_nand2_1 _30516_ (.Y(_21955_),
    .A(net6275),
    .B(_21954_));
 sg13g2_nand3_1 _30517_ (.B(_19975_),
    .C(_21925_),
    .A(_19951_),
    .Y(_21956_));
 sg13g2_nand2b_1 _30518_ (.Y(_21957_),
    .B(_21956_),
    .A_N(_21926_));
 sg13g2_o21ai_1 _30519_ (.B1(net6193),
    .Y(_21958_),
    .A1(\u_inv.f_next[206] ),
    .A2(net7303));
 sg13g2_a21o_1 _30520_ (.A2(_21957_),
    .A1(net7303),
    .B1(_21958_),
    .X(_21959_));
 sg13g2_o21ai_1 _30521_ (.B1(_21959_),
    .Y(_21960_),
    .A1(_21917_),
    .A2(_21955_));
 sg13g2_a21oi_1 _30522_ (.A1(_20930_),
    .A2(_20932_),
    .Y(_21961_),
    .B1(_20956_));
 sg13g2_a21oi_1 _30523_ (.A1(_20930_),
    .A2(_20932_),
    .Y(_21962_),
    .B1(_20958_));
 sg13g2_o21ai_1 _30524_ (.B1(_20936_),
    .Y(_21963_),
    .A1(_20996_),
    .A2(_21962_));
 sg13g2_or3_1 _30525_ (.A(_20936_),
    .B(_20996_),
    .C(_21962_),
    .X(_21964_));
 sg13g2_a21o_1 _30526_ (.A2(_21964_),
    .A1(_21963_),
    .B1(net7177),
    .X(_21965_));
 sg13g2_a21oi_1 _30527_ (.A1(_17975_),
    .A2(net7178),
    .Y(_21966_),
    .B1(net6276));
 sg13g2_a21oi_1 _30528_ (.A1(_21648_),
    .A2(_21715_),
    .Y(_21967_),
    .B1(_21721_));
 sg13g2_or3_1 _30529_ (.A(_20937_),
    .B(_21736_),
    .C(_21967_),
    .X(_21968_));
 sg13g2_o21ai_1 _30530_ (.B1(_20937_),
    .Y(_21969_),
    .A1(_21736_),
    .A2(_21967_));
 sg13g2_and2_1 _30531_ (.A(net6276),
    .B(_21969_),
    .X(_21970_));
 sg13g2_a22oi_1 _30532_ (.Y(_21971_),
    .B1(_21968_),
    .B2(_21970_),
    .A2(_21966_),
    .A1(_21965_));
 sg13g2_a21oi_2 _30533_ (.B1(_20918_),
    .Y(_21972_),
    .A2(_20912_),
    .A1(_20154_));
 sg13g2_nor2_1 _30534_ (.A(_20067_),
    .B(_21972_),
    .Y(_21973_));
 sg13g2_a21oi_2 _30535_ (.B1(_20071_),
    .Y(_21974_),
    .A2(_21972_),
    .A1(_20056_));
 sg13g2_nor3_1 _30536_ (.A(_20036_),
    .B(_20042_),
    .C(_21974_),
    .Y(_21975_));
 sg13g2_o21ai_1 _30537_ (.B1(_20029_),
    .Y(_21976_),
    .A1(_20081_),
    .A2(_21975_));
 sg13g2_nand2_1 _30538_ (.Y(_21977_),
    .A(_20028_),
    .B(_21976_));
 sg13g2_o21ai_1 _30539_ (.B1(net7314),
    .Y(_21978_),
    .A1(_20027_),
    .A2(_21977_));
 sg13g2_a21oi_1 _30540_ (.A1(_20027_),
    .A2(_21977_),
    .Y(_21979_),
    .B1(_21978_));
 sg13g2_o21ai_1 _30541_ (.B1(net6205),
    .Y(_21980_),
    .A1(\u_inv.f_next[189] ),
    .A2(net7314));
 sg13g2_a21oi_2 _30542_ (.B1(_21585_),
    .Y(_21981_),
    .A2(_21575_),
    .A1(_21543_));
 sg13g2_nor2_1 _30543_ (.A(_21602_),
    .B(_21981_),
    .Y(_21982_));
 sg13g2_o21ai_1 _30544_ (.B1(_21578_),
    .Y(_21983_),
    .A1(_21602_),
    .A2(_21981_));
 sg13g2_a21oi_1 _30545_ (.A1(_21616_),
    .A2(_21983_),
    .Y(_21984_),
    .B1(_20029_));
 sg13g2_or3_1 _30546_ (.A(_20027_),
    .B(_21603_),
    .C(_21984_),
    .X(_21985_));
 sg13g2_o21ai_1 _30547_ (.B1(_20027_),
    .Y(_21986_),
    .A1(_21603_),
    .A2(_21984_));
 sg13g2_nand3_1 _30548_ (.B(_21985_),
    .C(_21986_),
    .A(net6283),
    .Y(_21987_));
 sg13g2_o21ai_1 _30549_ (.B1(_21987_),
    .Y(_21988_),
    .A1(_21979_),
    .A2(_21980_));
 sg13g2_a21oi_1 _30550_ (.A1(_19937_),
    .A2(_21814_),
    .Y(_21989_),
    .B1(_19903_));
 sg13g2_and3_1 _30551_ (.X(_21990_),
    .A(_19903_),
    .B(_19937_),
    .C(_21814_));
 sg13g2_o21ai_1 _30552_ (.B1(net7303),
    .Y(_21991_),
    .A1(_21989_),
    .A2(_21990_));
 sg13g2_a21oi_1 _30553_ (.A1(_17981_),
    .A2(net7179),
    .Y(_21992_),
    .B1(net6274));
 sg13g2_nand2_1 _30554_ (.Y(_21993_),
    .A(_21991_),
    .B(_21992_));
 sg13g2_nor3_1 _30555_ (.A(_19903_),
    .B(_21714_),
    .C(_21823_),
    .Y(_21994_));
 sg13g2_nor2_1 _30556_ (.A(net6193),
    .B(_21994_),
    .Y(_21995_));
 sg13g2_nand2_1 _30557_ (.Y(_21996_),
    .A(net6275),
    .B(_21824_));
 sg13g2_a22oi_1 _30558_ (.Y(_21997_),
    .B1(_21995_),
    .B2(_21824_),
    .A2(_21992_),
    .A1(_21991_));
 sg13g2_o21ai_1 _30559_ (.B1(_21993_),
    .Y(_21998_),
    .A1(_21994_),
    .A2(_21996_));
 sg13g2_o21ai_1 _30560_ (.B1(_20069_),
    .Y(_21999_),
    .A1(_20055_),
    .A2(_21973_));
 sg13g2_xnor2_1 _30561_ (.Y(_22000_),
    .A(_20047_),
    .B(_21999_));
 sg13g2_o21ai_1 _30562_ (.B1(net6208),
    .Y(_22001_),
    .A1(\u_inv.f_next[182] ),
    .A2(net7317));
 sg13g2_a21oi_1 _30563_ (.A1(net7319),
    .A2(_22000_),
    .Y(_22002_),
    .B1(_22001_));
 sg13g2_a21oi_1 _30564_ (.A1(_21543_),
    .A2(_21575_),
    .Y(_22003_),
    .B1(_21583_));
 sg13g2_o21ai_1 _30565_ (.B1(_20052_),
    .Y(_22004_),
    .A1(_21594_),
    .A2(_22003_));
 sg13g2_a21oi_1 _30566_ (.A1(_21595_),
    .A2(_22004_),
    .Y(_22005_),
    .B1(_20054_));
 sg13g2_nor3_1 _30567_ (.A(_20048_),
    .B(_21596_),
    .C(_22005_),
    .Y(_22006_));
 sg13g2_o21ai_1 _30568_ (.B1(_20048_),
    .Y(_22007_),
    .A1(_21596_),
    .A2(_22005_));
 sg13g2_nor2_1 _30569_ (.A(net6208),
    .B(_22006_),
    .Y(_22008_));
 sg13g2_a21o_2 _30570_ (.A2(_22008_),
    .A1(_22007_),
    .B1(_22002_),
    .X(_22009_));
 sg13g2_a21oi_1 _30571_ (.A1(_20016_),
    .A2(_20928_),
    .Y(_22010_),
    .B1(_19940_));
 sg13g2_a21oi_1 _30572_ (.A1(\u_inv.f_next[208] ),
    .A2(\u_inv.f_reg[208] ),
    .Y(_22011_),
    .B1(_22010_));
 sg13g2_xnor2_1 _30573_ (.Y(_22012_),
    .A(_19938_),
    .B(_22011_));
 sg13g2_o21ai_1 _30574_ (.B1(net6192),
    .Y(_22013_),
    .A1(\u_inv.f_next[209] ),
    .A2(net7302));
 sg13g2_a21oi_1 _30575_ (.A1(net7302),
    .A2(_22012_),
    .Y(_22014_),
    .B1(_22013_));
 sg13g2_a21oi_1 _30576_ (.A1(_21681_),
    .A2(_21822_),
    .Y(_22015_),
    .B1(_19939_));
 sg13g2_nor3_1 _30577_ (.A(_19938_),
    .B(_21700_),
    .C(_22015_),
    .Y(_22016_));
 sg13g2_o21ai_1 _30578_ (.B1(_19938_),
    .Y(_22017_),
    .A1(_21700_),
    .A2(_22015_));
 sg13g2_nor2_1 _30579_ (.A(net6192),
    .B(_22016_),
    .Y(_22018_));
 sg13g2_a21o_2 _30580_ (.A2(_22018_),
    .A1(_22017_),
    .B1(_22014_),
    .X(_22019_));
 sg13g2_o21ai_1 _30581_ (.B1(_21019_),
    .Y(_22020_),
    .A1(_20991_),
    .A2(_21016_));
 sg13g2_nand3_1 _30582_ (.B(_21017_),
    .C(_21020_),
    .A(_20992_),
    .Y(_22021_));
 sg13g2_nand2_1 _30583_ (.Y(_22022_),
    .A(\u_inv.f_next[240] ),
    .B(net7182));
 sg13g2_nand3_1 _30584_ (.B(_22020_),
    .C(_22021_),
    .A(net7310),
    .Y(_22023_));
 sg13g2_xnor2_1 _30585_ (.Y(_22024_),
    .A(_21019_),
    .B(_21761_));
 sg13g2_nand3_1 _30586_ (.B(_22022_),
    .C(_22023_),
    .A(net6199),
    .Y(_22025_));
 sg13g2_o21ai_1 _30587_ (.B1(_22025_),
    .Y(_22026_),
    .A1(net6200),
    .A2(_22024_));
 sg13g2_inv_1 _30588_ (.Y(_22027_),
    .A(_22026_));
 sg13g2_nor3_1 _30589_ (.A(_19968_),
    .B(_20007_),
    .C(_21922_),
    .Y(_22028_));
 sg13g2_o21ai_1 _30590_ (.B1(_20007_),
    .Y(_22029_),
    .A1(_19968_),
    .A2(_21922_));
 sg13g2_nor2_1 _30591_ (.A(net7180),
    .B(_22028_),
    .Y(_22030_));
 sg13g2_o21ai_1 _30592_ (.B1(net6198),
    .Y(_22031_),
    .A1(\u_inv.f_next[201] ),
    .A2(net7308));
 sg13g2_a21o_1 _30593_ (.A2(_22030_),
    .A1(_22029_),
    .B1(_22031_),
    .X(_22032_));
 sg13g2_nor3_1 _30594_ (.A(_20007_),
    .B(_21666_),
    .C(_21913_),
    .Y(_22033_));
 sg13g2_o21ai_1 _30595_ (.B1(_20007_),
    .Y(_22034_),
    .A1(_21666_),
    .A2(_21913_));
 sg13g2_nand3b_1 _30596_ (.B(_22034_),
    .C(net6282),
    .Y(_22035_),
    .A_N(_22033_));
 sg13g2_nand2_1 _30597_ (.Y(_22036_),
    .A(_22032_),
    .B(_22035_));
 sg13g2_o21ai_1 _30598_ (.B1(_21533_),
    .Y(_22037_),
    .A1(_21497_),
    .A2(_21530_));
 sg13g2_a21oi_1 _30599_ (.A1(_21551_),
    .A2(_22037_),
    .Y(_22038_),
    .B1(_21535_));
 sg13g2_o21ai_1 _30600_ (.B1(_21539_),
    .Y(_22039_),
    .A1(_21571_),
    .A2(_22038_));
 sg13g2_a21o_1 _30601_ (.A2(_22039_),
    .A1(_21556_),
    .B1(_20096_),
    .X(_22040_));
 sg13g2_nor2_1 _30602_ (.A(_20097_),
    .B(_22040_),
    .Y(_22041_));
 sg13g2_o21ai_1 _30603_ (.B1(_20090_),
    .Y(_22042_),
    .A1(_21561_),
    .A2(_22041_));
 sg13g2_nor3_1 _30604_ (.A(_20090_),
    .B(_21561_),
    .C(_22041_),
    .Y(_22043_));
 sg13g2_nor2_1 _30605_ (.A(net6214),
    .B(_22043_),
    .Y(_22044_));
 sg13g2_and2_1 _30606_ (.A(_22042_),
    .B(_22044_),
    .X(_22045_));
 sg13g2_o21ai_1 _30607_ (.B1(_20909_),
    .Y(_22046_),
    .A1(_20227_),
    .A2(_20904_));
 sg13g2_nand2_2 _30608_ (.Y(_22047_),
    .A(_20144_),
    .B(_22046_));
 sg13g2_a21oi_1 _30609_ (.A1(_20144_),
    .A2(_22046_),
    .Y(_22048_),
    .B1(_20133_));
 sg13g2_nor2_1 _30610_ (.A(_20126_),
    .B(_22048_),
    .Y(_22049_));
 sg13g2_o21ai_1 _30611_ (.B1(_20114_),
    .Y(_22050_),
    .A1(_20126_),
    .A2(_22048_));
 sg13g2_nand2_1 _30612_ (.Y(_22051_),
    .A(_20148_),
    .B(_22050_));
 sg13g2_a21oi_1 _30613_ (.A1(_20148_),
    .A2(_22050_),
    .Y(_22052_),
    .B1(_20107_));
 sg13g2_nor2_1 _30614_ (.A(_20101_),
    .B(_22052_),
    .Y(_22053_));
 sg13g2_o21ai_1 _30615_ (.B1(_20098_),
    .Y(_22054_),
    .A1(_20101_),
    .A2(_22052_));
 sg13g2_a21o_1 _30616_ (.A2(_22054_),
    .A1(_20094_),
    .B1(_20090_),
    .X(_22055_));
 sg13g2_nand3_1 _30617_ (.B(_20094_),
    .C(_22054_),
    .A(_20090_),
    .Y(_22056_));
 sg13g2_a21o_1 _30618_ (.A2(_22056_),
    .A1(_22055_),
    .B1(net7196),
    .X(_22057_));
 sg13g2_a21oi_1 _30619_ (.A1(_18011_),
    .A2(net7196),
    .Y(_22058_),
    .B1(net6297));
 sg13g2_a22oi_1 _30620_ (.Y(_22059_),
    .B1(_22057_),
    .B2(_22058_),
    .A2(_22044_),
    .A1(_22042_));
 sg13g2_a21o_1 _30621_ (.A2(_22058_),
    .A1(_22057_),
    .B1(_22045_),
    .X(_22060_));
 sg13g2_o21ai_1 _30622_ (.B1(_20961_),
    .Y(_22061_),
    .A1(_21002_),
    .A2(_21852_));
 sg13g2_nand3_1 _30623_ (.B(_21003_),
    .C(_21853_),
    .A(_20962_),
    .Y(_22062_));
 sg13g2_nand2_1 _30624_ (.Y(_22063_),
    .A(\u_inv.f_next[232] ),
    .B(net7177));
 sg13g2_nand3_1 _30625_ (.B(_22061_),
    .C(_22062_),
    .A(net7305),
    .Y(_22064_));
 sg13g2_or3_1 _30626_ (.A(_20962_),
    .B(_21743_),
    .C(_21844_),
    .X(_22065_));
 sg13g2_and2_1 _30627_ (.A(_21845_),
    .B(_22065_),
    .X(_22066_));
 sg13g2_nand3_1 _30628_ (.B(_22063_),
    .C(_22064_),
    .A(net6194),
    .Y(_22067_));
 sg13g2_o21ai_1 _30629_ (.B1(_22067_),
    .Y(_22068_),
    .A1(net6194),
    .A2(_22066_));
 sg13g2_a21oi_1 _30630_ (.A1(_20154_),
    .A2(_20912_),
    .Y(_22069_),
    .B1(_20916_));
 sg13g2_a21oi_1 _30631_ (.A1(_20913_),
    .A2(_22069_),
    .Y(_22070_),
    .B1(_20063_));
 sg13g2_o21ai_1 _30632_ (.B1(_20057_),
    .Y(_22071_),
    .A1(_20059_),
    .A2(_22070_));
 sg13g2_xnor2_1 _30633_ (.Y(_22072_),
    .A(_20060_),
    .B(_22071_));
 sg13g2_o21ai_1 _30634_ (.B1(net6215),
    .Y(_22073_),
    .A1(\u_inv.f_next[179] ),
    .A2(net7326));
 sg13g2_a21oi_1 _30635_ (.A1(net7326),
    .A2(_22072_),
    .Y(_22074_),
    .B1(_22073_));
 sg13g2_a21oi_1 _30636_ (.A1(_21543_),
    .A2(_21575_),
    .Y(_22075_),
    .B1(_20915_));
 sg13g2_o21ai_1 _30637_ (.B1(_20914_),
    .Y(_22076_),
    .A1(_21589_),
    .A2(_22075_));
 sg13g2_a21oi_1 _30638_ (.A1(_21591_),
    .A2(_22076_),
    .Y(_22077_),
    .B1(_20058_));
 sg13g2_nor3_1 _30639_ (.A(_20061_),
    .B(_21588_),
    .C(_22077_),
    .Y(_22078_));
 sg13g2_o21ai_1 _30640_ (.B1(_20061_),
    .Y(_22079_),
    .A1(_21588_),
    .A2(_22077_));
 sg13g2_nor2_1 _30641_ (.A(net6215),
    .B(_22078_),
    .Y(_22080_));
 sg13g2_a21o_2 _30642_ (.A2(_22080_),
    .A1(_22079_),
    .B1(_22074_),
    .X(_22081_));
 sg13g2_inv_4 _30643_ (.A(_22081_),
    .Y(_22082_));
 sg13g2_o21ai_1 _30644_ (.B1(_20950_),
    .Y(_22083_),
    .A1(_20994_),
    .A2(_21961_));
 sg13g2_or3_1 _30645_ (.A(_20950_),
    .B(_20994_),
    .C(_21961_),
    .X(_22084_));
 sg13g2_nand3_1 _30646_ (.B(_22083_),
    .C(_22084_),
    .A(net7304),
    .Y(_22085_));
 sg13g2_a21oi_1 _30647_ (.A1(_21648_),
    .A2(_21715_),
    .Y(_22086_),
    .B1(_20953_));
 sg13g2_a21oi_1 _30648_ (.A1(_21648_),
    .A2(_21715_),
    .Y(_22087_),
    .B1(_21720_));
 sg13g2_nor2_1 _30649_ (.A(_21733_),
    .B(_22087_),
    .Y(_22088_));
 sg13g2_nor2_1 _30650_ (.A(_20950_),
    .B(_22088_),
    .Y(_22089_));
 sg13g2_xnor2_1 _30651_ (.Y(_22090_),
    .A(_20950_),
    .B(_22088_));
 sg13g2_a21oi_1 _30652_ (.A1(\u_inv.f_next[226] ),
    .A2(net7178),
    .Y(_22091_),
    .B1(net6277));
 sg13g2_a22oi_1 _30653_ (.Y(_22092_),
    .B1(_22091_),
    .B2(_22085_),
    .A2(_22090_),
    .A1(net6276));
 sg13g2_inv_1 _30654_ (.Y(_22093_),
    .A(_22092_));
 sg13g2_nand3_1 _30655_ (.B(_21739_),
    .C(_21969_),
    .A(_20934_),
    .Y(_22094_));
 sg13g2_a21o_1 _30656_ (.A2(_21969_),
    .A1(_21739_),
    .B1(_20934_),
    .X(_22095_));
 sg13g2_nand3_1 _30657_ (.B(_22094_),
    .C(_22095_),
    .A(net6277),
    .Y(_22096_));
 sg13g2_and3_1 _30658_ (.X(_22097_),
    .A(_20934_),
    .B(_20935_),
    .C(_21963_));
 sg13g2_a21oi_1 _30659_ (.A1(_20935_),
    .A2(_21963_),
    .Y(_22098_),
    .B1(_20934_));
 sg13g2_nor3_1 _30660_ (.A(net7178),
    .B(_22097_),
    .C(_22098_),
    .Y(_22099_));
 sg13g2_o21ai_1 _30661_ (.B1(net6194),
    .Y(_22100_),
    .A1(\u_inv.f_next[229] ),
    .A2(net7305));
 sg13g2_o21ai_1 _30662_ (.B1(_22096_),
    .Y(_22101_),
    .A1(_22099_),
    .A2(_22100_));
 sg13g2_a21oi_1 _30663_ (.A1(_20131_),
    .A2(_22047_),
    .Y(_22102_),
    .B1(_20124_));
 sg13g2_o21ai_1 _30664_ (.B1(_20117_),
    .Y(_22103_),
    .A1(_20119_),
    .A2(_22102_));
 sg13g2_xnor2_1 _30665_ (.Y(_22104_),
    .A(_20116_),
    .B(_22103_));
 sg13g2_nor2_1 _30666_ (.A(\u_inv.f_next[167] ),
    .B(net7329),
    .Y(_22105_));
 sg13g2_a21oi_1 _30667_ (.A1(net7329),
    .A2(_22104_),
    .Y(_22106_),
    .B1(_22105_));
 sg13g2_a21o_1 _30668_ (.A2(_22037_),
    .A1(_21551_),
    .B1(_20127_),
    .X(_22107_));
 sg13g2_a21oi_1 _30669_ (.A1(_21566_),
    .A2(_22107_),
    .Y(_22108_),
    .B1(_20129_));
 sg13g2_o21ai_1 _30670_ (.B1(_20119_),
    .Y(_22109_),
    .A1(_21567_),
    .A2(_22108_));
 sg13g2_nand3_1 _30671_ (.B(_21565_),
    .C(_22109_),
    .A(_20116_),
    .Y(_22110_));
 sg13g2_a21oi_1 _30672_ (.A1(_21565_),
    .A2(_22109_),
    .Y(_22111_),
    .B1(_20116_));
 sg13g2_nor2_1 _30673_ (.A(net6217),
    .B(_22111_),
    .Y(_22112_));
 sg13g2_a22oi_1 _30674_ (.Y(_22113_),
    .B1(_22110_),
    .B2(_22112_),
    .A2(_22106_),
    .A1(net6217));
 sg13g2_inv_1 _30675_ (.Y(_22114_),
    .A(_22113_));
 sg13g2_a21o_1 _30676_ (.A2(_20921_),
    .A1(_20086_),
    .B1(_20925_),
    .X(_22115_));
 sg13g2_a21oi_1 _30677_ (.A1(_19994_),
    .A2(_22115_),
    .Y(_22116_),
    .B1(_19991_));
 sg13g2_o21ai_1 _30678_ (.B1(_19985_),
    .Y(_22117_),
    .A1(_19997_),
    .A2(_22116_));
 sg13g2_o21ai_1 _30679_ (.B1(_22117_),
    .Y(_22118_),
    .A1(_17994_),
    .A2(_18244_));
 sg13g2_xnor2_1 _30680_ (.Y(_22119_),
    .A(_19983_),
    .B(_22118_));
 sg13g2_o21ai_1 _30681_ (.B1(net6197),
    .Y(_22120_),
    .A1(\u_inv.f_next[197] ),
    .A2(net7307));
 sg13g2_a21oi_1 _30682_ (.A1(net7308),
    .A2(_22119_),
    .Y(_22121_),
    .B1(_22120_));
 sg13g2_o21ai_1 _30683_ (.B1(_21642_),
    .Y(_22122_),
    .A1(_21587_),
    .A2(_21619_));
 sg13g2_nand2_1 _30684_ (.Y(_22123_),
    .A(_21658_),
    .B(_22122_));
 sg13g2_a21oi_1 _30685_ (.A1(_21658_),
    .A2(_22122_),
    .Y(_22124_),
    .B1(_19985_));
 sg13g2_nor3_1 _30686_ (.A(_19984_),
    .B(_21650_),
    .C(_22124_),
    .Y(_22125_));
 sg13g2_o21ai_1 _30687_ (.B1(_19984_),
    .Y(_22126_),
    .A1(_21650_),
    .A2(_22124_));
 sg13g2_nor2_1 _30688_ (.A(net6198),
    .B(_22125_),
    .Y(_22127_));
 sg13g2_a21oi_2 _30689_ (.B1(_22121_),
    .Y(_22128_),
    .A2(_22127_),
    .A1(_22126_));
 sg13g2_a21oi_1 _30690_ (.A1(_19941_),
    .A2(_20929_),
    .Y(_22129_),
    .B1(_19928_));
 sg13g2_a21oi_1 _30691_ (.A1(_20016_),
    .A2(_20928_),
    .Y(_22130_),
    .B1(_19943_));
 sg13g2_nor2_1 _30692_ (.A(_19930_),
    .B(_22130_),
    .Y(_22131_));
 sg13g2_o21ai_1 _30693_ (.B1(_19916_),
    .Y(_22132_),
    .A1(_19930_),
    .A2(_22130_));
 sg13g2_xnor2_1 _30694_ (.Y(_22133_),
    .A(_19917_),
    .B(_22131_));
 sg13g2_nor2_1 _30695_ (.A(\u_inv.f_next[212] ),
    .B(net7301),
    .Y(_22134_));
 sg13g2_a21oi_1 _30696_ (.A1(net7301),
    .A2(_22133_),
    .Y(_22135_),
    .B1(_22134_));
 sg13g2_a21oi_1 _30697_ (.A1(_21681_),
    .A2(_21822_),
    .Y(_22136_),
    .B1(_21623_));
 sg13g2_nor2_1 _30698_ (.A(_21706_),
    .B(_22136_),
    .Y(_22137_));
 sg13g2_nand2_1 _30699_ (.Y(_22138_),
    .A(_19916_),
    .B(_22137_));
 sg13g2_nor2_1 _30700_ (.A(_19916_),
    .B(_22137_),
    .Y(_22139_));
 sg13g2_nor2_1 _30701_ (.A(net6192),
    .B(_22139_),
    .Y(_22140_));
 sg13g2_a22oi_1 _30702_ (.Y(_22141_),
    .B1(_22138_),
    .B2(_22140_),
    .A2(_22135_),
    .A1(net6192));
 sg13g2_nand3_1 _30703_ (.B(_19915_),
    .C(_22132_),
    .A(_19913_),
    .Y(_22142_));
 sg13g2_a21o_1 _30704_ (.A2(_22132_),
    .A1(_19915_),
    .B1(_19913_),
    .X(_22143_));
 sg13g2_nand3_1 _30705_ (.B(_22142_),
    .C(_22143_),
    .A(net7301),
    .Y(_22144_));
 sg13g2_a21oi_1 _30706_ (.A1(_17983_),
    .A2(net7179),
    .Y(_22145_),
    .B1(net6274));
 sg13g2_nand3b_1 _30707_ (.B(_19913_),
    .C(_21707_),
    .Y(_22146_),
    .A_N(_22139_));
 sg13g2_o21ai_1 _30708_ (.B1(_21621_),
    .Y(_22147_),
    .A1(_21706_),
    .A2(_22136_));
 sg13g2_inv_1 _30709_ (.Y(_22148_),
    .A(_22147_));
 sg13g2_nor3_1 _30710_ (.A(net6192),
    .B(_21708_),
    .C(_22148_),
    .Y(_22149_));
 sg13g2_a22oi_1 _30711_ (.Y(_22150_),
    .B1(_22146_),
    .B2(_22149_),
    .A2(_22145_),
    .A1(_22144_));
 sg13g2_nand3_1 _30712_ (.B(_21771_),
    .C(_21946_),
    .A(_21023_),
    .Y(_22151_));
 sg13g2_o21ai_1 _30713_ (.B1(net6280),
    .Y(_22152_),
    .A1(_21023_),
    .A2(_21771_));
 sg13g2_nor2b_1 _30714_ (.A(_22152_),
    .B_N(_21947_),
    .Y(_22153_));
 sg13g2_nand3_1 _30715_ (.B(_21023_),
    .C(_22020_),
    .A(_21018_),
    .Y(_22154_));
 sg13g2_a21o_1 _30716_ (.A2(_22020_),
    .A1(_21018_),
    .B1(_21023_),
    .X(_22155_));
 sg13g2_nand3_1 _30717_ (.B(_22154_),
    .C(_22155_),
    .A(net7310),
    .Y(_22156_));
 sg13g2_a21oi_1 _30718_ (.A1(_17970_),
    .A2(net7182),
    .Y(_22157_),
    .B1(net6280));
 sg13g2_a22oi_1 _30719_ (.Y(_22158_),
    .B1(_22156_),
    .B2(_22157_),
    .A2(_22153_),
    .A1(_22151_));
 sg13g2_a21oi_1 _30720_ (.A1(_20883_),
    .A2(_20894_),
    .Y(_22159_),
    .B1(_20900_));
 sg13g2_nor2_1 _30721_ (.A(_20205_),
    .B(_22159_),
    .Y(_22160_));
 sg13g2_o21ai_1 _30722_ (.B1(_20200_),
    .Y(_22161_),
    .A1(_20205_),
    .A2(_22159_));
 sg13g2_nand2_1 _30723_ (.Y(_22162_),
    .A(_20208_),
    .B(_22161_));
 sg13g2_a21oi_1 _30724_ (.A1(_20187_),
    .A2(_22162_),
    .Y(_22163_),
    .B1(_20213_));
 sg13g2_xnor2_1 _30725_ (.Y(_22164_),
    .A(_20192_),
    .B(_22163_));
 sg13g2_nand2_1 _30726_ (.Y(_22165_),
    .A(net7357),
    .B(_22164_));
 sg13g2_a21oi_1 _30727_ (.A1(_18024_),
    .A2(net7212),
    .Y(_22166_),
    .B1(net6320));
 sg13g2_a21oi_1 _30728_ (.A1(_21472_),
    .A2(_21486_),
    .Y(_22167_),
    .B1(_20897_));
 sg13g2_a221oi_1 _30729_ (.B2(_21486_),
    .C1(_21491_),
    .B1(_21472_),
    .A1(_20204_),
    .Y(_22168_),
    .A2(_20896_));
 sg13g2_o21ai_1 _30730_ (.B1(_20186_),
    .Y(_22169_),
    .A1(_21520_),
    .A2(_22168_));
 sg13g2_nor2b_1 _30731_ (.A(_21513_),
    .B_N(_22169_),
    .Y(_22170_));
 sg13g2_nor2_1 _30732_ (.A(_20182_),
    .B(_22170_),
    .Y(_22171_));
 sg13g2_inv_1 _30733_ (.Y(_22172_),
    .A(_22171_));
 sg13g2_o21ai_1 _30734_ (.B1(_20192_),
    .Y(_22173_),
    .A1(_21512_),
    .A2(_22171_));
 sg13g2_or3_1 _30735_ (.A(_20192_),
    .B(_21512_),
    .C(_22171_),
    .X(_22174_));
 sg13g2_and3_1 _30736_ (.X(_22175_),
    .A(net6320),
    .B(_22173_),
    .C(_22174_));
 sg13g2_a21oi_1 _30737_ (.A1(_22165_),
    .A2(_22166_),
    .Y(_22176_),
    .B1(_22175_));
 sg13g2_a21o_1 _30738_ (.A2(_22166_),
    .A1(_22165_),
    .B1(_22175_),
    .X(_22177_));
 sg13g2_o21ai_1 _30739_ (.B1(_20862_),
    .Y(_22178_),
    .A1(_20845_),
    .A2(_20856_));
 sg13g2_o21ai_1 _30740_ (.B1(_20884_),
    .Y(_22179_),
    .A1(_20860_),
    .A2(_22178_));
 sg13g2_a21oi_1 _30741_ (.A1(_20880_),
    .A2(_22179_),
    .Y(_22180_),
    .B1(_20887_));
 sg13g2_a21o_1 _30742_ (.A2(_22179_),
    .A1(_20880_),
    .B1(_20887_),
    .X(_22181_));
 sg13g2_a21oi_1 _30743_ (.A1(_20867_),
    .A2(_22181_),
    .Y(_22182_),
    .B1(_20890_));
 sg13g2_o21ai_1 _30744_ (.B1(_20868_),
    .Y(_22183_),
    .A1(_20869_),
    .A2(_22182_));
 sg13g2_a21oi_1 _30745_ (.A1(_20874_),
    .A2(_22183_),
    .Y(_22184_),
    .B1(net7211));
 sg13g2_o21ai_1 _30746_ (.B1(_22184_),
    .Y(_22185_),
    .A1(_20874_),
    .A2(_22183_));
 sg13g2_o21ai_1 _30747_ (.B1(net6237),
    .Y(_22186_),
    .A1(\u_inv.f_next[143] ),
    .A2(net7360));
 sg13g2_inv_1 _30748_ (.Y(_22187_),
    .A(_22186_));
 sg13g2_a21o_2 _30749_ (.A2(_21469_),
    .A1(_21466_),
    .B1(_21479_),
    .X(_22188_));
 sg13g2_nand3_1 _30750_ (.B(_20866_),
    .C(_22188_),
    .A(_20864_),
    .Y(_22189_));
 sg13g2_a21oi_1 _30751_ (.A1(_21482_),
    .A2(_22189_),
    .Y(_22190_),
    .B1(_20870_));
 sg13g2_a21oi_1 _30752_ (.A1(\u_inv.f_next[142] ),
    .A2(_18226_),
    .Y(_22191_),
    .B1(_22190_));
 sg13g2_o21ai_1 _30753_ (.B1(net6319),
    .Y(_22192_),
    .A1(_20873_),
    .A2(_22191_));
 sg13g2_a21oi_1 _30754_ (.A1(_20873_),
    .A2(_22191_),
    .Y(_22193_),
    .B1(_22192_));
 sg13g2_a21oi_2 _30755_ (.B1(_22193_),
    .Y(_22194_),
    .A2(_22187_),
    .A1(_22185_));
 sg13g2_a21oi_1 _30756_ (.A1(_20182_),
    .A2(_22170_),
    .Y(_22195_),
    .B1(net6235));
 sg13g2_a21oi_1 _30757_ (.A1(_20208_),
    .A2(_22161_),
    .Y(_22196_),
    .B1(_20186_));
 sg13g2_or3_1 _30758_ (.A(_20183_),
    .B(_20184_),
    .C(_22196_),
    .X(_22197_));
 sg13g2_o21ai_1 _30759_ (.B1(_20183_),
    .Y(_22198_),
    .A1(_20184_),
    .A2(_22196_));
 sg13g2_nand3_1 _30760_ (.B(_22197_),
    .C(_22198_),
    .A(net7357),
    .Y(_22199_));
 sg13g2_a21oi_1 _30761_ (.A1(_18025_),
    .A2(net7212),
    .Y(_22200_),
    .B1(net6320));
 sg13g2_a22oi_1 _30762_ (.Y(_22201_),
    .B1(_22199_),
    .B2(_22200_),
    .A2(_22195_),
    .A1(_22172_));
 sg13g2_inv_1 _30763_ (.Y(_22202_),
    .A(_22201_));
 sg13g2_nor2_1 _30764_ (.A(_20797_),
    .B(_21375_),
    .Y(_22203_));
 sg13g2_o21ai_1 _30765_ (.B1(_21386_),
    .Y(_22204_),
    .A1(_20797_),
    .A2(_21375_));
 sg13g2_nor2b_1 _30766_ (.A(_20795_),
    .B_N(_22204_),
    .Y(_22205_));
 sg13g2_o21ai_1 _30767_ (.B1(_20792_),
    .Y(_22206_),
    .A1(_21388_),
    .A2(_22205_));
 sg13g2_nor2b_1 _30768_ (.A(_21384_),
    .B_N(_22206_),
    .Y(_22207_));
 sg13g2_a21oi_1 _30769_ (.A1(_20793_),
    .A2(_22207_),
    .Y(_22208_),
    .B1(net6251));
 sg13g2_o21ai_1 _30770_ (.B1(_22208_),
    .Y(_22209_),
    .A1(_20793_),
    .A2(_22207_));
 sg13g2_a21oi_1 _30771_ (.A1(_20763_),
    .A2(_20775_),
    .Y(_22210_),
    .B1(_20798_));
 sg13g2_nor2_2 _30772_ (.A(_20803_),
    .B(_22210_),
    .Y(_22211_));
 sg13g2_o21ai_1 _30773_ (.B1(_20790_),
    .Y(_22212_),
    .A1(_20792_),
    .A2(_22211_));
 sg13g2_xnor2_1 _30774_ (.Y(_22213_),
    .A(_20793_),
    .B(_22212_));
 sg13g2_a21oi_1 _30775_ (.A1(net7381),
    .A2(_22213_),
    .Y(_22214_),
    .B1(net6345));
 sg13g2_o21ai_1 _30776_ (.B1(_22214_),
    .Y(_22215_),
    .A1(\u_inv.f_next[107] ),
    .A2(net7381));
 sg13g2_nand2_2 _30777_ (.Y(_22216_),
    .A(_22209_),
    .B(_22215_));
 sg13g2_or3_1 _30778_ (.A(_20845_),
    .B(_20856_),
    .C(_20862_),
    .X(_22217_));
 sg13g2_nand3_1 _30779_ (.B(_22178_),
    .C(_22217_),
    .A(net7360),
    .Y(_22218_));
 sg13g2_a21oi_1 _30780_ (.A1(_21448_),
    .A2(_21465_),
    .Y(_22219_),
    .B1(_20862_));
 sg13g2_xor2_1 _30781_ (.B(_21466_),
    .A(_20862_),
    .X(_22220_));
 sg13g2_a21oi_1 _30782_ (.A1(\u_inv.f_next[136] ),
    .A2(net7211),
    .Y(_22221_),
    .B1(net6323));
 sg13g2_a22oi_1 _30783_ (.Y(_22222_),
    .B1(_22221_),
    .B2(_22218_),
    .A2(_22220_),
    .A1(net6323));
 sg13g2_o21ai_1 _30784_ (.B1(_20815_),
    .Y(_22223_),
    .A1(_20801_),
    .A2(_20811_));
 sg13g2_nand2_2 _30785_ (.Y(_22224_),
    .A(_20274_),
    .B(_22223_));
 sg13g2_a21oi_2 _30786_ (.B1(_20277_),
    .Y(_22225_),
    .A2(_22224_),
    .A1(_20270_));
 sg13g2_o21ai_1 _30787_ (.B1(_20259_),
    .Y(_22226_),
    .A1(_20260_),
    .A2(_22225_));
 sg13g2_xnor2_1 _30788_ (.Y(_22227_),
    .A(_20258_),
    .B(_22226_));
 sg13g2_nand2_1 _30789_ (.Y(_22228_),
    .A(net7380),
    .B(_22227_));
 sg13g2_a21oi_1 _30790_ (.A1(_18041_),
    .A2(net7228),
    .Y(_22229_),
    .B1(net6333));
 sg13g2_nand2b_1 _30791_ (.Y(_22230_),
    .B(_21399_),
    .A_N(_21405_));
 sg13g2_a21o_1 _30792_ (.A2(_22230_),
    .A1(_21419_),
    .B1(_20261_),
    .X(_22231_));
 sg13g2_a21oi_1 _30793_ (.A1(_21412_),
    .A2(_22231_),
    .Y(_22232_),
    .B1(_20258_));
 sg13g2_nand3_1 _30794_ (.B(_21412_),
    .C(_22231_),
    .A(_20258_),
    .Y(_22233_));
 sg13g2_nor2_1 _30795_ (.A(net6251),
    .B(_22232_),
    .Y(_22234_));
 sg13g2_a22oi_1 _30796_ (.Y(_22235_),
    .B1(_22233_),
    .B2(_22234_),
    .A2(_22229_),
    .A1(_22228_));
 sg13g2_inv_2 _30797_ (.Y(_22236_),
    .A(_22235_));
 sg13g2_o21ai_1 _30798_ (.B1(_20816_),
    .Y(_22237_),
    .A1(_20801_),
    .A2(_20811_));
 sg13g2_nand2_1 _30799_ (.Y(_22238_),
    .A(_20283_),
    .B(_22237_));
 sg13g2_a21oi_1 _30800_ (.A1(_20283_),
    .A2(_22237_),
    .Y(_22239_),
    .B1(_20243_));
 sg13g2_nor2_1 _30801_ (.A(_20290_),
    .B(_22239_),
    .Y(_22240_));
 sg13g2_o21ai_1 _30802_ (.B1(_20249_),
    .Y(_22241_),
    .A1(_20290_),
    .A2(_22239_));
 sg13g2_nand2_1 _30803_ (.Y(_22242_),
    .A(_20293_),
    .B(_22241_));
 sg13g2_a21oi_1 _30804_ (.A1(_20293_),
    .A2(_22241_),
    .Y(_22243_),
    .B1(_20236_));
 sg13g2_xnor2_1 _30805_ (.Y(_22244_),
    .A(_20235_),
    .B(_22242_));
 sg13g2_o21ai_1 _30806_ (.B1(net6245),
    .Y(_22245_),
    .A1(\u_inv.f_next[124] ),
    .A2(net7371));
 sg13g2_a21oi_1 _30807_ (.A1(net7371),
    .A2(_22244_),
    .Y(_22246_),
    .B1(_22245_));
 sg13g2_o21ai_1 _30808_ (.B1(_21407_),
    .Y(_22247_),
    .A1(_21380_),
    .A2(_21397_));
 sg13g2_and2_1 _30809_ (.A(_21426_),
    .B(_22247_),
    .X(_22248_));
 sg13g2_or2_1 _30810_ (.X(_22249_),
    .B(_22248_),
    .A(_21400_));
 sg13g2_nand3_1 _30811_ (.B(_21440_),
    .C(_22249_),
    .A(_20235_),
    .Y(_22250_));
 sg13g2_a21oi_1 _30812_ (.A1(_21440_),
    .A2(_22249_),
    .Y(_22251_),
    .B1(_20235_));
 sg13g2_nor2_1 _30813_ (.A(net6245),
    .B(_22251_),
    .Y(_22252_));
 sg13g2_a21oi_1 _30814_ (.A1(_22250_),
    .A2(_22252_),
    .Y(_22253_),
    .B1(_22246_));
 sg13g2_inv_1 _30815_ (.Y(_22254_),
    .A(_22253_));
 sg13g2_xnor2_1 _30816_ (.Y(_22255_),
    .A(_20266_),
    .B(_22224_));
 sg13g2_a21oi_1 _30817_ (.A1(net7380),
    .A2(_22255_),
    .Y(_22256_),
    .B1(net6344));
 sg13g2_o21ai_1 _30818_ (.B1(_22256_),
    .Y(_22257_),
    .A1(\u_inv.f_next[114] ),
    .A2(net7380));
 sg13g2_and2_1 _30819_ (.A(_20814_),
    .B(_21399_),
    .X(_22258_));
 sg13g2_o21ai_1 _30820_ (.B1(_20813_),
    .Y(_22259_),
    .A1(_21415_),
    .A2(_22258_));
 sg13g2_a21oi_1 _30821_ (.A1(_21417_),
    .A2(_22259_),
    .Y(_22260_),
    .B1(_20266_));
 sg13g2_nand3_1 _30822_ (.B(_21417_),
    .C(_22259_),
    .A(_20266_),
    .Y(_22261_));
 sg13g2_nand2_1 _30823_ (.Y(_22262_),
    .A(net6344),
    .B(_22261_));
 sg13g2_o21ai_1 _30824_ (.B1(_22257_),
    .Y(_22263_),
    .A1(_22260_),
    .A2(_22262_));
 sg13g2_a21oi_1 _30825_ (.A1(_20242_),
    .A2(_22238_),
    .Y(_22264_),
    .B1(_20241_));
 sg13g2_o21ai_1 _30826_ (.B1(net7372),
    .Y(_22265_),
    .A1(_20240_),
    .A2(_22264_));
 sg13g2_a21oi_1 _30827_ (.A1(_20240_),
    .A2(_22264_),
    .Y(_22266_),
    .B1(_22265_));
 sg13g2_o21ai_1 _30828_ (.B1(net6246),
    .Y(_22267_),
    .A1(\u_inv.f_next[121] ),
    .A2(net7372));
 sg13g2_a21o_1 _30829_ (.A2(_22247_),
    .A1(_21426_),
    .B1(_20242_),
    .X(_22268_));
 sg13g2_a21oi_1 _30830_ (.A1(_21433_),
    .A2(_22268_),
    .Y(_22269_),
    .B1(_20240_));
 sg13g2_nand3_1 _30831_ (.B(_21433_),
    .C(_22268_),
    .A(_20240_),
    .Y(_22270_));
 sg13g2_nand3b_1 _30832_ (.B(_22270_),
    .C(net6334),
    .Y(_22271_),
    .A_N(_22269_));
 sg13g2_o21ai_1 _30833_ (.B1(_22271_),
    .Y(_22272_),
    .A1(_22266_),
    .A2(_22267_));
 sg13g2_a21oi_2 _30834_ (.B1(_20822_),
    .Y(_22273_),
    .A2(_20819_),
    .A1(_20295_));
 sg13g2_a21oi_1 _30835_ (.A1(\u_inv.f_next[128] ),
    .A2(\u_inv.f_reg[128] ),
    .Y(_22274_),
    .B1(_22273_));
 sg13g2_xor2_1 _30836_ (.B(_22274_),
    .A(_20821_),
    .X(_22275_));
 sg13g2_o21ai_1 _30837_ (.B1(net6243),
    .Y(_22276_),
    .A1(\u_inv.f_next[129] ),
    .A2(net7367));
 sg13g2_a21o_1 _30838_ (.A2(_22275_),
    .A1(net7368),
    .B1(_22276_),
    .X(_22277_));
 sg13g2_nand2_1 _30839_ (.Y(_22278_),
    .A(_20822_),
    .B(_21443_));
 sg13g2_a21oi_1 _30840_ (.A1(_21451_),
    .A2(_22278_),
    .Y(_22279_),
    .B1(_20821_));
 sg13g2_nand3_1 _30841_ (.B(_21451_),
    .C(_22278_),
    .A(_20821_),
    .Y(_22280_));
 sg13g2_nand2_1 _30842_ (.Y(_22281_),
    .A(net6334),
    .B(_22280_));
 sg13g2_o21ai_1 _30843_ (.B1(_22277_),
    .Y(_22282_),
    .A1(_22279_),
    .A2(_22281_));
 sg13g2_o21ai_1 _30844_ (.B1(_21376_),
    .Y(_22283_),
    .A1(_21358_),
    .A2(_21373_));
 sg13g2_a21oi_1 _30845_ (.A1(_21391_),
    .A2(_22283_),
    .Y(_22284_),
    .B1(_20786_));
 sg13g2_o21ai_1 _30846_ (.B1(_20784_),
    .Y(_22285_),
    .A1(_21383_),
    .A2(_22284_));
 sg13g2_a21oi_1 _30847_ (.A1(_21382_),
    .A2(_22285_),
    .Y(_22286_),
    .B1(_20780_));
 sg13g2_o21ai_1 _30848_ (.B1(_20778_),
    .Y(_22287_),
    .A1(_21395_),
    .A2(_22286_));
 sg13g2_or3_1 _30849_ (.A(_20778_),
    .B(_21395_),
    .C(_22286_),
    .X(_22288_));
 sg13g2_nand3_1 _30850_ (.B(_22287_),
    .C(_22288_),
    .A(net6344),
    .Y(_22289_));
 sg13g2_o21ai_1 _30851_ (.B1(_20806_),
    .Y(_22290_),
    .A1(_20794_),
    .A2(_22211_));
 sg13g2_a21oi_1 _30852_ (.A1(_20788_),
    .A2(_22290_),
    .Y(_22291_),
    .B1(_20809_));
 sg13g2_nand2b_1 _30853_ (.Y(_22292_),
    .B(_20780_),
    .A_N(_22291_));
 sg13g2_nand2_1 _30854_ (.Y(_22293_),
    .A(_20779_),
    .B(_22292_));
 sg13g2_o21ai_1 _30855_ (.B1(net7382),
    .Y(_22294_),
    .A1(_20778_),
    .A2(_22293_));
 sg13g2_a21oi_1 _30856_ (.A1(_20778_),
    .A2(_22293_),
    .Y(_22295_),
    .B1(_22294_));
 sg13g2_o21ai_1 _30857_ (.B1(net6252),
    .Y(_22296_),
    .A1(\u_inv.f_next[111] ),
    .A2(net7382));
 sg13g2_o21ai_1 _30858_ (.B1(_22289_),
    .Y(_22297_),
    .A1(_22295_),
    .A2(_22296_));
 sg13g2_xnor2_1 _30859_ (.Y(_22298_),
    .A(_20866_),
    .B(_22180_));
 sg13g2_o21ai_1 _30860_ (.B1(net6233),
    .Y(_22299_),
    .A1(\u_inv.f_next[140] ),
    .A2(net7356));
 sg13g2_a21oi_1 _30861_ (.A1(net7356),
    .A2(_22298_),
    .Y(_22300_),
    .B1(_22299_));
 sg13g2_a21oi_1 _30862_ (.A1(_20866_),
    .A2(_22188_),
    .Y(_22301_),
    .B1(net6237));
 sg13g2_o21ai_1 _30863_ (.B1(_22301_),
    .Y(_22302_),
    .A1(_20866_),
    .A2(_22188_));
 sg13g2_nor2b_2 _30864_ (.A(_22300_),
    .B_N(_22302_),
    .Y(_22303_));
 sg13g2_nand3_1 _30865_ (.B(_20759_),
    .C(_21353_),
    .A(_20756_),
    .Y(_22304_));
 sg13g2_nand2_1 _30866_ (.Y(_22305_),
    .A(_21364_),
    .B(_22304_));
 sg13g2_nand2b_1 _30867_ (.Y(_22306_),
    .B(_22305_),
    .A_N(_21355_));
 sg13g2_a21oi_1 _30868_ (.A1(_21366_),
    .A2(_22306_),
    .Y(_22307_),
    .B1(_20735_));
 sg13g2_o21ai_1 _30869_ (.B1(_20733_),
    .Y(_22308_),
    .A1(_21368_),
    .A2(_22307_));
 sg13g2_a21oi_1 _30870_ (.A1(_21370_),
    .A2(_22308_),
    .Y(_22309_),
    .B1(_20743_));
 sg13g2_o21ai_1 _30871_ (.B1(_20741_),
    .Y(_22310_),
    .A1(_21361_),
    .A2(_22309_));
 sg13g2_nor3_1 _30872_ (.A(_20741_),
    .B(_21361_),
    .C(_22309_),
    .Y(_22311_));
 sg13g2_nand2_1 _30873_ (.Y(_22312_),
    .A(net6348),
    .B(_22310_));
 sg13g2_o21ai_1 _30874_ (.B1(_20765_),
    .Y(_22313_),
    .A1(_20730_),
    .A2(_20760_));
 sg13g2_and2_1 _30875_ (.A(_20752_),
    .B(_22313_),
    .X(_22314_));
 sg13g2_nor2_1 _30876_ (.A(_20769_),
    .B(_22314_),
    .Y(_22315_));
 sg13g2_o21ai_1 _30877_ (.B1(_20737_),
    .Y(_22316_),
    .A1(_20769_),
    .A2(_22314_));
 sg13g2_a21oi_1 _30878_ (.A1(_20773_),
    .A2(_22316_),
    .Y(_22317_),
    .B1(_20744_));
 sg13g2_a21oi_1 _30879_ (.A1(\u_inv.f_next[102] ),
    .A2(\u_inv.f_reg[102] ),
    .Y(_22318_),
    .B1(_22317_));
 sg13g2_xnor2_1 _30880_ (.Y(_22319_),
    .A(_20741_),
    .B(_22318_));
 sg13g2_a21oi_1 _30881_ (.A1(net7387),
    .A2(_22319_),
    .Y(_22320_),
    .B1(net6356));
 sg13g2_o21ai_1 _30882_ (.B1(_22320_),
    .Y(_22321_),
    .A1(\u_inv.f_next[103] ),
    .A2(net7387));
 sg13g2_o21ai_1 _30883_ (.B1(_22321_),
    .Y(_22322_),
    .A1(_22311_),
    .A2(_22312_));
 sg13g2_xnor2_1 _30884_ (.Y(_22323_),
    .A(_20261_),
    .B(_22225_));
 sg13g2_nor2_1 _30885_ (.A(net7228),
    .B(_22323_),
    .Y(_22324_));
 sg13g2_o21ai_1 _30886_ (.B1(net6251),
    .Y(_22325_),
    .A1(\u_inv.f_next[116] ),
    .A2(net7380));
 sg13g2_nand3_1 _30887_ (.B(_21419_),
    .C(_22230_),
    .A(_20261_),
    .Y(_22326_));
 sg13g2_nand3_1 _30888_ (.B(_22231_),
    .C(_22326_),
    .A(net6333),
    .Y(_22327_));
 sg13g2_o21ai_1 _30889_ (.B1(_22327_),
    .Y(_22328_),
    .A1(_22324_),
    .A2(_22325_));
 sg13g2_nor2_1 _30890_ (.A(_20812_),
    .B(_20814_),
    .Y(_22329_));
 sg13g2_a21oi_1 _30891_ (.A1(\u_inv.f_next[112] ),
    .A2(\u_inv.f_reg[112] ),
    .Y(_22330_),
    .B1(_22329_));
 sg13g2_xnor2_1 _30892_ (.Y(_22331_),
    .A(_20813_),
    .B(_22330_));
 sg13g2_o21ai_1 _30893_ (.B1(net6251),
    .Y(_22332_),
    .A1(\u_inv.f_next[113] ),
    .A2(net7380));
 sg13g2_a21oi_1 _30894_ (.A1(net7380),
    .A2(_22331_),
    .Y(_22333_),
    .B1(_22332_));
 sg13g2_nor3_1 _30895_ (.A(_20813_),
    .B(_21415_),
    .C(_22258_),
    .Y(_22334_));
 sg13g2_nor2_1 _30896_ (.A(net6251),
    .B(_22334_),
    .Y(_22335_));
 sg13g2_a21oi_2 _30897_ (.B1(_22333_),
    .Y(_22336_),
    .A2(_22335_),
    .A1(_22259_));
 sg13g2_xnor2_1 _30898_ (.Y(_22337_),
    .A(_20822_),
    .B(_21443_));
 sg13g2_nand3_1 _30899_ (.B(_20819_),
    .C(_20822_),
    .A(_20295_),
    .Y(_22338_));
 sg13g2_nand3b_1 _30900_ (.B(_22338_),
    .C(net7367),
    .Y(_22339_),
    .A_N(_22273_));
 sg13g2_a21oi_1 _30901_ (.A1(\u_inv.f_next[128] ),
    .A2(net7219),
    .Y(_22340_),
    .B1(net6334));
 sg13g2_a22oi_1 _30902_ (.Y(_22341_),
    .B1(_22339_),
    .B2(_22340_),
    .A2(_22337_),
    .A1(net6334));
 sg13g2_nand2_1 _30903_ (.Y(_22342_),
    .A(_20786_),
    .B(_22290_));
 sg13g2_nand2_1 _30904_ (.Y(_22343_),
    .A(_20785_),
    .B(_22342_));
 sg13g2_o21ai_1 _30905_ (.B1(net7381),
    .Y(_22344_),
    .A1(_20784_),
    .A2(_22343_));
 sg13g2_a21oi_1 _30906_ (.A1(_20784_),
    .A2(_22343_),
    .Y(_22345_),
    .B1(_22344_));
 sg13g2_o21ai_1 _30907_ (.B1(net6252),
    .Y(_22346_),
    .A1(\u_inv.f_next[109] ),
    .A2(net7382));
 sg13g2_or3_1 _30908_ (.A(_20784_),
    .B(_21383_),
    .C(_22284_),
    .X(_22347_));
 sg13g2_nand3_1 _30909_ (.B(_22285_),
    .C(_22347_),
    .A(net6345),
    .Y(_22348_));
 sg13g2_o21ai_1 _30910_ (.B1(_22348_),
    .Y(_22349_),
    .A1(_22345_),
    .A2(_22346_));
 sg13g2_xnor2_1 _30911_ (.Y(_22350_),
    .A(_20814_),
    .B(_21399_));
 sg13g2_a21oi_1 _30912_ (.A1(_20812_),
    .A2(_20814_),
    .Y(_22351_),
    .B1(net7227));
 sg13g2_nand2b_1 _30913_ (.Y(_22352_),
    .B(_22351_),
    .A_N(_22329_));
 sg13g2_a21oi_1 _30914_ (.A1(\u_inv.f_next[112] ),
    .A2(net7228),
    .Y(_22353_),
    .B1(net6344));
 sg13g2_a22oi_1 _30915_ (.Y(_22354_),
    .B1(_22352_),
    .B2(_22353_),
    .A2(_22350_),
    .A1(net6344));
 sg13g2_a21oi_1 _30916_ (.A1(_20776_),
    .A2(_20797_),
    .Y(_22355_),
    .B1(_20796_));
 sg13g2_a21oi_1 _30917_ (.A1(_20795_),
    .A2(_22355_),
    .Y(_22356_),
    .B1(net7227));
 sg13g2_o21ai_1 _30918_ (.B1(_22356_),
    .Y(_22357_),
    .A1(_20795_),
    .A2(_22355_));
 sg13g2_a21oi_1 _30919_ (.A1(_18049_),
    .A2(net7227),
    .Y(_22358_),
    .B1(net6344));
 sg13g2_xnor2_1 _30920_ (.Y(_22359_),
    .A(_20795_),
    .B(_22204_));
 sg13g2_a22oi_1 _30921_ (.Y(_22360_),
    .B1(_22359_),
    .B2(net6345),
    .A2(_22358_),
    .A1(_22357_));
 sg13g2_xnor2_1 _30922_ (.Y(_22361_),
    .A(_20786_),
    .B(_22290_));
 sg13g2_nor2_1 _30923_ (.A(\u_inv.f_next[108] ),
    .B(net7381),
    .Y(_22362_));
 sg13g2_a21oi_1 _30924_ (.A1(net7381),
    .A2(_22361_),
    .Y(_22363_),
    .B1(_22362_));
 sg13g2_nand3_1 _30925_ (.B(_21391_),
    .C(_22283_),
    .A(_20786_),
    .Y(_22364_));
 sg13g2_nor2_1 _30926_ (.A(net6251),
    .B(_22284_),
    .Y(_22365_));
 sg13g2_a22oi_1 _30927_ (.Y(_22366_),
    .B1(_22364_),
    .B2(_22365_),
    .A2(_22363_),
    .A1(net6251));
 sg13g2_nand2_2 _30928_ (.Y(_22367_),
    .A(_22360_),
    .B(_22366_));
 sg13g2_xnor2_1 _30929_ (.Y(_22368_),
    .A(_20792_),
    .B(_22211_));
 sg13g2_a21oi_1 _30930_ (.A1(net7381),
    .A2(_22368_),
    .Y(_22369_),
    .B1(net6345));
 sg13g2_o21ai_1 _30931_ (.B1(_22369_),
    .Y(_22370_),
    .A1(\u_inv.f_next[106] ),
    .A2(net7381));
 sg13g2_nor3_1 _30932_ (.A(_20792_),
    .B(_21388_),
    .C(_22205_),
    .Y(_22371_));
 sg13g2_nand2_1 _30933_ (.Y(_22372_),
    .A(net6345),
    .B(_22206_));
 sg13g2_o21ai_1 _30934_ (.B1(_22370_),
    .Y(_22373_),
    .A1(_22371_),
    .A2(_22372_));
 sg13g2_xnor2_1 _30935_ (.Y(_22374_),
    .A(_20242_),
    .B(_22238_));
 sg13g2_o21ai_1 _30936_ (.B1(net6245),
    .Y(_22375_),
    .A1(\u_inv.f_next[120] ),
    .A2(net7371));
 sg13g2_a21oi_1 _30937_ (.A1(net7372),
    .A2(_22374_),
    .Y(_22376_),
    .B1(_22375_));
 sg13g2_a21oi_1 _30938_ (.A1(_20242_),
    .A2(_22248_),
    .Y(_22377_),
    .B1(net6246));
 sg13g2_a21o_2 _30939_ (.A2(_22377_),
    .A1(_22268_),
    .B1(_22376_),
    .X(_22378_));
 sg13g2_a21oi_2 _30940_ (.B1(_20847_),
    .Y(_22379_),
    .A2(_22273_),
    .A1(_20821_));
 sg13g2_o21ai_1 _30941_ (.B1(_20849_),
    .Y(_22380_),
    .A1(_20842_),
    .A2(_22379_));
 sg13g2_xnor2_1 _30942_ (.Y(_22381_),
    .A(_20825_),
    .B(_22380_));
 sg13g2_o21ai_1 _30943_ (.B1(net6241),
    .Y(_22382_),
    .A1(\u_inv.f_next[132] ),
    .A2(net7365));
 sg13g2_a21o_1 _30944_ (.A2(_22381_),
    .A1(net7367),
    .B1(_22382_),
    .X(_22383_));
 sg13g2_o21ai_1 _30945_ (.B1(_21446_),
    .Y(_22384_),
    .A1(_21409_),
    .A2(_21442_));
 sg13g2_and2_1 _30946_ (.A(_21457_),
    .B(_22384_),
    .X(_22385_));
 sg13g2_a21oi_1 _30947_ (.A1(_21457_),
    .A2(_22384_),
    .Y(_22386_),
    .B1(_20825_));
 sg13g2_a21o_1 _30948_ (.A2(_22385_),
    .A1(_20825_),
    .B1(net6242),
    .X(_22387_));
 sg13g2_o21ai_1 _30949_ (.B1(_22383_),
    .Y(_22388_),
    .A1(_22386_),
    .A2(_22387_));
 sg13g2_nand3_1 _30950_ (.B(_21382_),
    .C(_22285_),
    .A(_20780_),
    .Y(_22389_));
 sg13g2_nand2b_1 _30951_ (.Y(_22390_),
    .B(_22389_),
    .A_N(_22286_));
 sg13g2_nand2b_1 _30952_ (.Y(_22391_),
    .B(_22291_),
    .A_N(_20780_));
 sg13g2_nand3_1 _30953_ (.B(_22292_),
    .C(_22391_),
    .A(net7382),
    .Y(_22392_));
 sg13g2_a21oi_1 _30954_ (.A1(\u_inv.f_next[110] ),
    .A2(net7228),
    .Y(_22393_),
    .B1(net6345));
 sg13g2_a22oi_1 _30955_ (.Y(_22394_),
    .B1(_22392_),
    .B2(_22393_),
    .A2(_22390_),
    .A1(net6345));
 sg13g2_nand3_1 _30956_ (.B(_20773_),
    .C(_22316_),
    .A(_20744_),
    .Y(_22395_));
 sg13g2_nand2b_1 _30957_ (.Y(_22396_),
    .B(_22395_),
    .A_N(_22317_));
 sg13g2_nor2_1 _30958_ (.A(\u_inv.f_next[102] ),
    .B(net7387),
    .Y(_22397_));
 sg13g2_a21oi_1 _30959_ (.A1(net7387),
    .A2(_22396_),
    .Y(_22398_),
    .B1(_22397_));
 sg13g2_nand3_1 _30960_ (.B(_21370_),
    .C(_22308_),
    .A(_20743_),
    .Y(_22399_));
 sg13g2_nor2_1 _30961_ (.A(net6255),
    .B(_22309_),
    .Y(_22400_));
 sg13g2_a22oi_1 _30962_ (.Y(_22401_),
    .B1(_22399_),
    .B2(_22400_),
    .A2(_22398_),
    .A1(net6255));
 sg13g2_inv_4 _30963_ (.A(_22401_),
    .Y(_22402_));
 sg13g2_nor3_1 _30964_ (.A(_20733_),
    .B(_21368_),
    .C(_22307_),
    .Y(_22403_));
 sg13g2_nor2_1 _30965_ (.A(net6255),
    .B(_22403_),
    .Y(_22404_));
 sg13g2_o21ai_1 _30966_ (.B1(_20734_),
    .Y(_22405_),
    .A1(_20736_),
    .A2(_22315_));
 sg13g2_xnor2_1 _30967_ (.Y(_22406_),
    .A(_20732_),
    .B(_22405_));
 sg13g2_o21ai_1 _30968_ (.B1(net6255),
    .Y(_22407_),
    .A1(\u_inv.f_next[101] ),
    .A2(net7387));
 sg13g2_a21oi_1 _30969_ (.A1(net7387),
    .A2(_22406_),
    .Y(_22408_),
    .B1(_22407_));
 sg13g2_a21o_2 _30970_ (.A2(_22404_),
    .A1(_22308_),
    .B1(_22408_),
    .X(_22409_));
 sg13g2_a21oi_1 _30971_ (.A1(_20694_),
    .A2(_20717_),
    .Y(_22410_),
    .B1(_20720_));
 sg13g2_o21ai_1 _30972_ (.B1(_20723_),
    .Y(_22411_),
    .A1(_20709_),
    .A2(_22410_));
 sg13g2_a21oi_1 _30973_ (.A1(_20704_),
    .A2(_22411_),
    .Y(_22412_),
    .B1(_20727_));
 sg13g2_nor2b_1 _30974_ (.A(_22412_),
    .B_N(_20699_),
    .Y(_22413_));
 sg13g2_nor2_1 _30975_ (.A(_20698_),
    .B(_22413_),
    .Y(_22414_));
 sg13g2_xnor2_1 _30976_ (.Y(_22415_),
    .A(_20696_),
    .B(_22414_));
 sg13g2_nor2_1 _30977_ (.A(\u_inv.f_next[95] ),
    .B(net7402),
    .Y(_22416_));
 sg13g2_a21oi_1 _30978_ (.A1(net7402),
    .A2(_22415_),
    .Y(_22417_),
    .B1(_22416_));
 sg13g2_nor2b_1 _30979_ (.A(_21333_),
    .B_N(_21336_),
    .Y(_22418_));
 sg13g2_nand2b_1 _30980_ (.Y(_22419_),
    .B(_21336_),
    .A_N(_21333_));
 sg13g2_a21oi_1 _30981_ (.A1(_21335_),
    .A2(_22418_),
    .Y(_22420_),
    .B1(_21347_));
 sg13g2_or2_1 _30982_ (.X(_22421_),
    .B(_22420_),
    .A(_20703_));
 sg13g2_a21o_1 _30983_ (.A2(_22421_),
    .A1(_21341_),
    .B1(_20701_),
    .X(_22422_));
 sg13g2_a21oi_1 _30984_ (.A1(_21340_),
    .A2(_22422_),
    .Y(_22423_),
    .B1(_20699_));
 sg13g2_nor3_1 _30985_ (.A(_20696_),
    .B(_21351_),
    .C(_22423_),
    .Y(_22424_));
 sg13g2_o21ai_1 _30986_ (.B1(_20696_),
    .Y(_22425_),
    .A1(_21351_),
    .A2(_22423_));
 sg13g2_nor2_1 _30987_ (.A(net6265),
    .B(_22424_),
    .Y(_22426_));
 sg13g2_a22oi_1 _30988_ (.Y(_22427_),
    .B1(_22425_),
    .B2(_22426_),
    .A2(_22417_),
    .A1(net6265));
 sg13g2_a21oi_1 _30989_ (.A1(_21364_),
    .A2(_22304_),
    .Y(_22428_),
    .B1(_20750_));
 sg13g2_nor3_1 _30990_ (.A(_20748_),
    .B(_21365_),
    .C(_22428_),
    .Y(_22429_));
 sg13g2_a21oi_1 _30991_ (.A1(_20748_),
    .A2(_21365_),
    .Y(_22430_),
    .B1(net6255));
 sg13g2_nand2_1 _30992_ (.Y(_22431_),
    .A(_22306_),
    .B(_22430_));
 sg13g2_a21oi_1 _30993_ (.A1(_20750_),
    .A2(_22313_),
    .Y(_22432_),
    .B1(_20749_));
 sg13g2_xnor2_1 _30994_ (.Y(_22433_),
    .A(_20748_),
    .B(_22432_));
 sg13g2_a21oi_1 _30995_ (.A1(net7388),
    .A2(_22433_),
    .Y(_22434_),
    .B1(net6348));
 sg13g2_o21ai_1 _30996_ (.B1(_22434_),
    .Y(_22435_),
    .A1(\u_inv.f_next[99] ),
    .A2(net7388));
 sg13g2_o21ai_1 _30997_ (.B1(_22435_),
    .Y(_22436_),
    .A1(_22429_),
    .A2(_22431_));
 sg13g2_a21oi_1 _30998_ (.A1(_20703_),
    .A2(_22411_),
    .Y(_22437_),
    .B1(_20702_));
 sg13g2_o21ai_1 _30999_ (.B1(net7402),
    .Y(_22438_),
    .A1(_20701_),
    .A2(_22437_));
 sg13g2_a21oi_1 _31000_ (.A1(_20701_),
    .A2(_22437_),
    .Y(_22439_),
    .B1(_22438_));
 sg13g2_o21ai_1 _31001_ (.B1(net6265),
    .Y(_22440_),
    .A1(\u_inv.f_next[93] ),
    .A2(net7402));
 sg13g2_nand3_1 _31002_ (.B(_21341_),
    .C(_22421_),
    .A(_20701_),
    .Y(_22441_));
 sg13g2_nand3_1 _31003_ (.B(_22422_),
    .C(_22441_),
    .A(net6359),
    .Y(_22442_));
 sg13g2_o21ai_1 _31004_ (.B1(_22442_),
    .Y(_22443_),
    .A1(_22439_),
    .A2(_22440_));
 sg13g2_xnor2_1 _31005_ (.Y(_22444_),
    .A(_20750_),
    .B(_22313_));
 sg13g2_o21ai_1 _31006_ (.B1(net6255),
    .Y(_22445_),
    .A1(\u_inv.f_next[98] ),
    .A2(net7388));
 sg13g2_a21oi_1 _31007_ (.A1(net7388),
    .A2(_22444_),
    .Y(_22446_),
    .B1(_22445_));
 sg13g2_o21ai_1 _31008_ (.B1(net6348),
    .Y(_22447_),
    .A1(_20751_),
    .A2(_22305_));
 sg13g2_nor2_1 _31009_ (.A(_22428_),
    .B(_22447_),
    .Y(_22448_));
 sg13g2_nor2_2 _31010_ (.A(_22446_),
    .B(_22448_),
    .Y(_22449_));
 sg13g2_a21oi_1 _31011_ (.A1(_20685_),
    .A2(_21322_),
    .Y(_22450_),
    .B1(_21325_));
 sg13g2_nor2_1 _31012_ (.A(_20682_),
    .B(_22450_),
    .Y(_22451_));
 sg13g2_o21ai_1 _31013_ (.B1(_20676_),
    .Y(_22452_),
    .A1(_21327_),
    .A2(_22451_));
 sg13g2_nand2_1 _31014_ (.Y(_22453_),
    .A(_21329_),
    .B(_22452_));
 sg13g2_o21ai_1 _31015_ (.B1(net6360),
    .Y(_22454_),
    .A1(_20680_),
    .A2(_22453_));
 sg13g2_a21oi_1 _31016_ (.A1(_20680_),
    .A2(_22453_),
    .Y(_22455_),
    .B1(_22454_));
 sg13g2_o21ai_1 _31017_ (.B1(_20691_),
    .Y(_22456_),
    .A1(_20673_),
    .A2(_20686_));
 sg13g2_a21oi_1 _31018_ (.A1(_20675_),
    .A2(_22456_),
    .Y(_22457_),
    .B1(_20674_));
 sg13g2_a21oi_1 _31019_ (.A1(_20679_),
    .A2(_22457_),
    .Y(_22458_),
    .B1(net7236));
 sg13g2_o21ai_1 _31020_ (.B1(_22458_),
    .Y(_22459_),
    .A1(_20679_),
    .A2(_22457_));
 sg13g2_a21oi_1 _31021_ (.A1(_18056_),
    .A2(net7236),
    .Y(_22460_),
    .B1(net6360));
 sg13g2_a21oi_1 _31022_ (.A1(_22459_),
    .A2(_22460_),
    .Y(_22461_),
    .B1(_22455_));
 sg13g2_inv_1 _31023_ (.Y(_22462_),
    .A(_22461_));
 sg13g2_o21ai_1 _31024_ (.B1(_20707_),
    .Y(_22463_),
    .A1(_20708_),
    .A2(_22410_));
 sg13g2_a21oi_1 _31025_ (.A1(_20706_),
    .A2(_22463_),
    .Y(_22464_),
    .B1(net7244));
 sg13g2_o21ai_1 _31026_ (.B1(_22464_),
    .Y(_22465_),
    .A1(_20706_),
    .A2(_22463_));
 sg13g2_o21ai_1 _31027_ (.B1(_22465_),
    .Y(_22466_),
    .A1(\u_inv.f_next[91] ),
    .A2(net7403));
 sg13g2_o21ai_1 _31028_ (.B1(_20708_),
    .Y(_22467_),
    .A1(_21344_),
    .A2(_22418_));
 sg13g2_nand2b_1 _31029_ (.Y(_22468_),
    .B(_22467_),
    .A_N(_21342_));
 sg13g2_a21oi_1 _31030_ (.A1(_20706_),
    .A2(_22468_),
    .Y(_22469_),
    .B1(net6265));
 sg13g2_o21ai_1 _31031_ (.B1(_22469_),
    .Y(_22470_),
    .A1(_20706_),
    .A2(_22468_));
 sg13g2_o21ai_1 _31032_ (.B1(_22470_),
    .Y(_22471_),
    .A1(net6359),
    .A2(_22466_));
 sg13g2_xnor2_1 _31033_ (.Y(_22472_),
    .A(_20776_),
    .B(_20797_));
 sg13g2_nor2_1 _31034_ (.A(\u_inv.f_next[104] ),
    .B(net7381),
    .Y(_22473_));
 sg13g2_a21oi_1 _31035_ (.A1(net7382),
    .A2(_22472_),
    .Y(_22474_),
    .B1(_22473_));
 sg13g2_nand2_1 _31036_ (.Y(_22475_),
    .A(_20797_),
    .B(_21375_));
 sg13g2_nor2_1 _31037_ (.A(net6252),
    .B(_22203_),
    .Y(_22476_));
 sg13g2_a22oi_1 _31038_ (.Y(_22477_),
    .B1(_22475_),
    .B2(_22476_),
    .A2(_22474_),
    .A1(net6251));
 sg13g2_inv_2 _31039_ (.Y(_22478_),
    .A(_22477_));
 sg13g2_xnor2_1 _31040_ (.Y(_22479_),
    .A(_20703_),
    .B(_22411_));
 sg13g2_nor2_1 _31041_ (.A(\u_inv.f_next[92] ),
    .B(net7403),
    .Y(_22480_));
 sg13g2_a21oi_1 _31042_ (.A1(net7403),
    .A2(_22479_),
    .Y(_22481_),
    .B1(_22480_));
 sg13g2_nand2_1 _31043_ (.Y(_22482_),
    .A(_20703_),
    .B(_22420_));
 sg13g2_and2_1 _31044_ (.A(net6359),
    .B(_22421_),
    .X(_22483_));
 sg13g2_a22oi_1 _31045_ (.Y(_22484_),
    .B1(_22482_),
    .B2(_22483_),
    .A2(_22481_),
    .A1(net6265));
 sg13g2_a21oi_1 _31046_ (.A1(_20759_),
    .A2(_21353_),
    .Y(_22485_),
    .B1(_20756_));
 sg13g2_nand3b_1 _31047_ (.B(_22304_),
    .C(net6348),
    .Y(_22486_),
    .A_N(_21363_));
 sg13g2_a21oi_1 _31048_ (.A1(_21362_),
    .A2(_22485_),
    .Y(_22487_),
    .B1(_22486_));
 sg13g2_o21ai_1 _31049_ (.B1(_20757_),
    .Y(_22488_),
    .A1(_20730_),
    .A2(_20759_));
 sg13g2_xnor2_1 _31050_ (.Y(_22489_),
    .A(_20755_),
    .B(_22488_));
 sg13g2_o21ai_1 _31051_ (.B1(net6256),
    .Y(_22490_),
    .A1(\u_inv.f_next[97] ),
    .A2(net7388));
 sg13g2_a21oi_1 _31052_ (.A1(net7388),
    .A2(_22489_),
    .Y(_22491_),
    .B1(_22490_));
 sg13g2_nor2_2 _31053_ (.A(_22487_),
    .B(_22491_),
    .Y(_22492_));
 sg13g2_inv_2 _31054_ (.Y(_22493_),
    .A(_22492_));
 sg13g2_a21oi_1 _31055_ (.A1(\u_inv.f_next[88] ),
    .A2(_18212_),
    .Y(_22494_),
    .B1(_20713_));
 sg13g2_o21ai_1 _31056_ (.B1(_22494_),
    .Y(_22495_),
    .A1(_20715_),
    .A2(_21333_));
 sg13g2_nand4_1 _31057_ (.B(_21343_),
    .C(_22419_),
    .A(net6359),
    .Y(_22496_),
    .D(_22495_));
 sg13g2_nand2_1 _31058_ (.Y(_22497_),
    .A(_20694_),
    .B(_20715_));
 sg13g2_nand3_1 _31059_ (.B(_20714_),
    .C(_22497_),
    .A(_20712_),
    .Y(_22498_));
 sg13g2_a21oi_1 _31060_ (.A1(_20714_),
    .A2(_22497_),
    .Y(_22499_),
    .B1(_20712_));
 sg13g2_nand2_1 _31061_ (.Y(_22500_),
    .A(net7402),
    .B(_22498_));
 sg13g2_nor2_1 _31062_ (.A(\u_inv.f_next[89] ),
    .B(net7402),
    .Y(_22501_));
 sg13g2_o21ai_1 _31063_ (.B1(net6265),
    .Y(_22502_),
    .A1(_22499_),
    .A2(_22500_));
 sg13g2_o21ai_1 _31064_ (.B1(_22496_),
    .Y(_22503_),
    .A1(_22501_),
    .A2(_22502_));
 sg13g2_nand2b_1 _31065_ (.Y(_22504_),
    .B(_21276_),
    .A_N(_20605_));
 sg13g2_nand2_1 _31066_ (.Y(_22505_),
    .A(_21276_),
    .B(_21277_));
 sg13g2_nand2b_1 _31067_ (.Y(_22506_),
    .B(_22505_),
    .A_N(_21284_));
 sg13g2_and2_1 _31068_ (.A(_20597_),
    .B(_22506_),
    .X(_22507_));
 sg13g2_nor2_1 _31069_ (.A(_21281_),
    .B(_22507_),
    .Y(_22508_));
 sg13g2_nor2_1 _31070_ (.A(_20599_),
    .B(_22508_),
    .Y(_22509_));
 sg13g2_nand2_1 _31071_ (.Y(_22510_),
    .A(_20599_),
    .B(_22508_));
 sg13g2_nor2_1 _31072_ (.A(net6264),
    .B(_22509_),
    .Y(_22511_));
 sg13g2_nand2_1 _31073_ (.Y(_22512_),
    .A(_22510_),
    .B(_22511_));
 sg13g2_a21oi_1 _31074_ (.A1(_20595_),
    .A2(_20606_),
    .Y(_22513_),
    .B1(_20611_));
 sg13g2_o21ai_1 _31075_ (.B1(_20596_),
    .Y(_22514_),
    .A1(_20597_),
    .A2(_22513_));
 sg13g2_a21oi_1 _31076_ (.A1(_20600_),
    .A2(_22514_),
    .Y(_22515_),
    .B1(net7236));
 sg13g2_o21ai_1 _31077_ (.B1(_22515_),
    .Y(_22516_),
    .A1(_20600_),
    .A2(_22514_));
 sg13g2_nor2_1 _31078_ (.A(\u_inv.f_next[71] ),
    .B(net7397),
    .Y(_22517_));
 sg13g2_nor2_1 _31079_ (.A(net6358),
    .B(_22517_),
    .Y(_22518_));
 sg13g2_nand2_1 _31080_ (.Y(_22519_),
    .A(net6264),
    .B(_22516_));
 sg13g2_a22oi_1 _31081_ (.Y(_22520_),
    .B1(_22516_),
    .B2(_22518_),
    .A2(_22511_),
    .A1(_22510_));
 sg13g2_o21ai_1 _31082_ (.B1(_22512_),
    .Y(_22521_),
    .A1(_22517_),
    .A2(_22519_));
 sg13g2_xnor2_1 _31083_ (.Y(_22522_),
    .A(_20597_),
    .B(_22513_));
 sg13g2_a21oi_1 _31084_ (.A1(net7397),
    .A2(_22522_),
    .Y(_22523_),
    .B1(net6358));
 sg13g2_o21ai_1 _31085_ (.B1(_22523_),
    .Y(_22524_),
    .A1(\u_inv.f_next[70] ),
    .A2(net7397));
 sg13g2_o21ai_1 _31086_ (.B1(net6358),
    .Y(_22525_),
    .A1(_20597_),
    .A2(_22506_));
 sg13g2_o21ai_1 _31087_ (.B1(_22524_),
    .Y(_22526_),
    .A1(_22507_),
    .A2(_22525_));
 sg13g2_a21oi_2 _31088_ (.B1(_20563_),
    .Y(_22527_),
    .A2(_20560_),
    .A1(_20535_));
 sg13g2_o21ai_1 _31089_ (.B1(_20567_),
    .Y(_22528_),
    .A1(_20552_),
    .A2(_22527_));
 sg13g2_nand3_1 _31090_ (.B(_20538_),
    .C(_22528_),
    .A(_20536_),
    .Y(_22529_));
 sg13g2_nand2_1 _31091_ (.Y(_22530_),
    .A(_20572_),
    .B(_22529_));
 sg13g2_nand2_1 _31092_ (.Y(_22531_),
    .A(_20544_),
    .B(_22530_));
 sg13g2_a21oi_1 _31093_ (.A1(_20543_),
    .A2(_22531_),
    .Y(_22532_),
    .B1(_20542_));
 sg13g2_nand3_1 _31094_ (.B(_20543_),
    .C(_22531_),
    .A(_20542_),
    .Y(_22533_));
 sg13g2_nor2_1 _31095_ (.A(net7237),
    .B(_22532_),
    .Y(_22534_));
 sg13g2_a221oi_1 _31096_ (.B2(_22534_),
    .C1(net6361),
    .B1(_22533_),
    .A1(_18070_),
    .Y(_22535_),
    .A2(net7237));
 sg13g2_a21oi_1 _31097_ (.A1(_21247_),
    .A2(_21259_),
    .Y(_22536_),
    .B1(_20538_));
 sg13g2_nor2_1 _31098_ (.A(_21252_),
    .B(_22536_),
    .Y(_22537_));
 sg13g2_or2_1 _31099_ (.X(_22538_),
    .B(_22537_),
    .A(_20536_));
 sg13g2_a21o_1 _31100_ (.A2(_22538_),
    .A1(_21251_),
    .B1(_20544_),
    .X(_22539_));
 sg13g2_nand2_1 _31101_ (.Y(_22540_),
    .A(_21250_),
    .B(_22539_));
 sg13g2_xnor2_1 _31102_ (.Y(_22541_),
    .A(_20542_),
    .B(_22540_));
 sg13g2_a21oi_1 _31103_ (.A1(net6361),
    .A2(_22541_),
    .Y(_22542_),
    .B1(_22535_));
 sg13g2_inv_1 _31104_ (.Y(_22543_),
    .A(_22542_));
 sg13g2_nor2_1 _31105_ (.A(_20603_),
    .B(_21282_),
    .Y(_22544_));
 sg13g2_nand3_1 _31106_ (.B(_21283_),
    .C(_22505_),
    .A(net6358),
    .Y(_22545_));
 sg13g2_a21oi_1 _31107_ (.A1(_22504_),
    .A2(_22544_),
    .Y(_22546_),
    .B1(_22545_));
 sg13g2_a21oi_1 _31108_ (.A1(_20595_),
    .A2(_20605_),
    .Y(_22547_),
    .B1(_20604_));
 sg13g2_xnor2_1 _31109_ (.Y(_22548_),
    .A(_20603_),
    .B(_22547_));
 sg13g2_o21ai_1 _31110_ (.B1(net6264),
    .Y(_22549_),
    .A1(\u_inv.f_next[69] ),
    .A2(net7397));
 sg13g2_a21oi_1 _31111_ (.A1(net7397),
    .A2(_22548_),
    .Y(_22550_),
    .B1(_22549_));
 sg13g2_nor2_1 _31112_ (.A(_22546_),
    .B(_22550_),
    .Y(_22551_));
 sg13g2_inv_1 _31113_ (.Y(_22552_),
    .A(_22551_));
 sg13g2_xnor2_1 _31114_ (.Y(_22553_),
    .A(_20544_),
    .B(_22530_));
 sg13g2_o21ai_1 _31115_ (.B1(net6260),
    .Y(_22554_),
    .A1(\u_inv.f_next[62] ),
    .A2(net7395));
 sg13g2_a21oi_1 _31116_ (.A1(net7395),
    .A2(_22553_),
    .Y(_22555_),
    .B1(_22554_));
 sg13g2_nand3_1 _31117_ (.B(_21251_),
    .C(_22538_),
    .A(_20544_),
    .Y(_22556_));
 sg13g2_nand3_1 _31118_ (.B(_22539_),
    .C(_22556_),
    .A(net6361),
    .Y(_22557_));
 sg13g2_nand2b_2 _31119_ (.Y(_22558_),
    .B(_22557_),
    .A_N(_22555_));
 sg13g2_o21ai_1 _31120_ (.B1(_20585_),
    .Y(_22559_),
    .A1(_20576_),
    .A2(_20586_));
 sg13g2_xor2_1 _31121_ (.B(_22559_),
    .A(_20584_),
    .X(_22560_));
 sg13g2_o21ai_1 _31122_ (.B1(net6260),
    .Y(_22561_),
    .A1(\u_inv.f_next[65] ),
    .A2(net7396));
 sg13g2_a21o_1 _31123_ (.A2(_22560_),
    .A1(net7396),
    .B1(_22561_),
    .X(_22562_));
 sg13g2_a21o_1 _31124_ (.A2(_21265_),
    .A1(_20586_),
    .B1(_21268_),
    .X(_22563_));
 sg13g2_xnor2_1 _31125_ (.Y(_22564_),
    .A(_20584_),
    .B(_22563_));
 sg13g2_o21ai_1 _31126_ (.B1(_22562_),
    .Y(_22565_),
    .A1(net6260),
    .A2(_22564_));
 sg13g2_xnor2_1 _31127_ (.Y(_22566_),
    .A(_20595_),
    .B(_20605_));
 sg13g2_o21ai_1 _31128_ (.B1(net6264),
    .Y(_22567_),
    .A1(\u_inv.f_next[68] ),
    .A2(net7397));
 sg13g2_a21oi_1 _31129_ (.A1(net7397),
    .A2(_22566_),
    .Y(_22568_),
    .B1(_22567_));
 sg13g2_xnor2_1 _31130_ (.Y(_22569_),
    .A(_20605_),
    .B(_21276_));
 sg13g2_a21oi_2 _31131_ (.B1(_22568_),
    .Y(_22570_),
    .A2(_22569_),
    .A1(net6358));
 sg13g2_nor2b_1 _31132_ (.A(_21238_),
    .B_N(_21239_),
    .Y(_22571_));
 sg13g2_or2_1 _31133_ (.X(_22572_),
    .B(_22571_),
    .A(_20522_));
 sg13g2_a21oi_1 _31134_ (.A1(_21094_),
    .A2(_22572_),
    .Y(_22573_),
    .B1(_20518_));
 sg13g2_a21oi_1 _31135_ (.A1(\u_inv.f_next[54] ),
    .A2(_18204_),
    .Y(_22574_),
    .B1(_22573_));
 sg13g2_o21ai_1 _31136_ (.B1(net6348),
    .Y(_22575_),
    .A1(_20519_),
    .A2(_22574_));
 sg13g2_a21oi_1 _31137_ (.A1(_20519_),
    .A2(_22574_),
    .Y(_22576_),
    .B1(_22575_));
 sg13g2_a21oi_1 _31138_ (.A1(_20515_),
    .A2(_20527_),
    .Y(_22577_),
    .B1(_20532_));
 sg13g2_o21ai_1 _31139_ (.B1(_20516_),
    .Y(_22578_),
    .A1(_20517_),
    .A2(_22577_));
 sg13g2_xnor2_1 _31140_ (.Y(_22579_),
    .A(_20519_),
    .B(_22578_));
 sg13g2_nand2_1 _31141_ (.Y(_22580_),
    .A(net7384),
    .B(_22579_));
 sg13g2_a21oi_1 _31142_ (.A1(_18074_),
    .A2(net7229),
    .Y(_22581_),
    .B1(net6347));
 sg13g2_a21oi_1 _31143_ (.A1(_22580_),
    .A2(_22581_),
    .Y(_22582_),
    .B1(_22576_));
 sg13g2_a21o_1 _31144_ (.A2(_22581_),
    .A1(_22580_),
    .B1(_22576_),
    .X(_22583_));
 sg13g2_o21ai_1 _31145_ (.B1(net7395),
    .Y(_22584_),
    .A1(_20550_),
    .A2(_22527_));
 sg13g2_a21o_1 _31146_ (.A2(_22527_),
    .A1(_20550_),
    .B1(_22584_),
    .X(_22585_));
 sg13g2_and2_1 _31147_ (.A(_21246_),
    .B(_21254_),
    .X(_22586_));
 sg13g2_nand2_1 _31148_ (.Y(_22587_),
    .A(_21255_),
    .B(_22586_));
 sg13g2_xnor2_1 _31149_ (.Y(_22588_),
    .A(_20550_),
    .B(_22587_));
 sg13g2_a21oi_1 _31150_ (.A1(\u_inv.f_next[58] ),
    .A2(net7237),
    .Y(_22589_),
    .B1(net6347));
 sg13g2_a22oi_1 _31151_ (.Y(_22590_),
    .B1(_22589_),
    .B2(_22585_),
    .A2(_22588_),
    .A1(net6347));
 sg13g2_xnor2_1 _31152_ (.Y(_22591_),
    .A(_20538_),
    .B(_22528_));
 sg13g2_o21ai_1 _31153_ (.B1(net6260),
    .Y(_22592_),
    .A1(\u_inv.f_next[60] ),
    .A2(net7395));
 sg13g2_a21oi_1 _31154_ (.A1(net7395),
    .A2(_22591_),
    .Y(_22593_),
    .B1(_22592_));
 sg13g2_nand3_1 _31155_ (.B(_21247_),
    .C(_21259_),
    .A(_20538_),
    .Y(_22594_));
 sg13g2_nor2_1 _31156_ (.A(net6260),
    .B(_22536_),
    .Y(_22595_));
 sg13g2_a21o_2 _31157_ (.A2(_22595_),
    .A1(_22594_),
    .B1(_22593_),
    .X(_22596_));
 sg13g2_xor2_1 _31158_ (.B(_21265_),
    .A(_20586_),
    .X(_22597_));
 sg13g2_a21oi_1 _31159_ (.A1(_20576_),
    .A2(_20586_),
    .Y(_22598_),
    .B1(net7237));
 sg13g2_o21ai_1 _31160_ (.B1(_22598_),
    .Y(_22599_),
    .A1(_20576_),
    .A2(_20586_));
 sg13g2_nand2_1 _31161_ (.Y(_22600_),
    .A(\u_inv.f_next[64] ),
    .B(net7237));
 sg13g2_nand3_1 _31162_ (.B(_22599_),
    .C(_22600_),
    .A(net6261),
    .Y(_22601_));
 sg13g2_o21ai_1 _31163_ (.B1(_22601_),
    .Y(_22602_),
    .A1(net6261),
    .A2(_22597_));
 sg13g2_nor2_1 _31164_ (.A(_20503_),
    .B(_20507_),
    .Y(_22603_));
 sg13g2_o21ai_1 _31165_ (.B1(_20505_),
    .Y(_22604_),
    .A1(_20508_),
    .A2(_22603_));
 sg13g2_o21ai_1 _31166_ (.B1(net7386),
    .Y(_22605_),
    .A1(_20509_),
    .A2(_22604_));
 sg13g2_a21o_1 _31167_ (.A2(_22604_),
    .A1(_20509_),
    .B1(_22605_),
    .X(_22606_));
 sg13g2_o21ai_1 _31168_ (.B1(_22606_),
    .Y(_22607_),
    .A1(\u_inv.f_next[51] ),
    .A2(net7386));
 sg13g2_a21oi_1 _31169_ (.A1(_21230_),
    .A2(_21231_),
    .Y(_22608_),
    .B1(_20499_));
 sg13g2_or2_1 _31170_ (.X(_22609_),
    .B(_22608_),
    .A(_21097_));
 sg13g2_nand2_1 _31171_ (.Y(_22610_),
    .A(_20508_),
    .B(_22609_));
 sg13g2_nand2b_1 _31172_ (.Y(_22611_),
    .B(_22610_),
    .A_N(_21096_));
 sg13g2_a21oi_1 _31173_ (.A1(_20509_),
    .A2(_22611_),
    .Y(_22612_),
    .B1(net6253));
 sg13g2_o21ai_1 _31174_ (.B1(_22612_),
    .Y(_22613_),
    .A1(_20509_),
    .A2(_22611_));
 sg13g2_o21ai_1 _31175_ (.B1(_22613_),
    .Y(_22614_),
    .A1(net6347),
    .A2(_22607_));
 sg13g2_nand2_1 _31176_ (.Y(_22615_),
    .A(_20535_),
    .B(_20558_));
 sg13g2_xnor2_1 _31177_ (.Y(_22616_),
    .A(_20535_),
    .B(_20558_));
 sg13g2_o21ai_1 _31178_ (.B1(net6253),
    .Y(_22617_),
    .A1(\u_inv.f_next[56] ),
    .A2(net7385));
 sg13g2_a21oi_1 _31179_ (.A1(net7385),
    .A2(_22616_),
    .Y(_22618_),
    .B1(_22617_));
 sg13g2_xnor2_1 _31180_ (.Y(_22619_),
    .A(_20558_),
    .B(_21245_));
 sg13g2_a21oi_2 _31181_ (.B1(_22618_),
    .Y(_22620_),
    .A2(_22619_),
    .A1(net6347));
 sg13g2_a21oi_2 _31182_ (.B1(_20318_),
    .Y(_22621_),
    .A2(_20492_),
    .A1(_20489_));
 sg13g2_o21ai_1 _31183_ (.B1(_20311_),
    .Y(_22622_),
    .A1(_20313_),
    .A2(_22621_));
 sg13g2_o21ai_1 _31184_ (.B1(net7379),
    .Y(_22623_),
    .A1(_20309_),
    .A2(_22622_));
 sg13g2_a21oi_1 _31185_ (.A1(_20309_),
    .A2(_22622_),
    .Y(_22624_),
    .B1(_22623_));
 sg13g2_o21ai_1 _31186_ (.B1(net6250),
    .Y(_22625_),
    .A1(\u_inv.f_next[43] ),
    .A2(net7378));
 sg13g2_nand2_1 _31187_ (.Y(_22626_),
    .A(_20490_),
    .B(_21207_));
 sg13g2_nand2_1 _31188_ (.Y(_22627_),
    .A(_21217_),
    .B(_22626_));
 sg13g2_nand2_1 _31189_ (.Y(_22628_),
    .A(_20491_),
    .B(_22627_));
 sg13g2_and2_1 _31190_ (.A(_21219_),
    .B(_22628_),
    .X(_22629_));
 sg13g2_or2_1 _31191_ (.X(_22630_),
    .B(_22629_),
    .A(_20312_));
 sg13g2_a21o_1 _31192_ (.A2(_22630_),
    .A1(_21221_),
    .B1(_20310_),
    .X(_22631_));
 sg13g2_nand3_1 _31193_ (.B(_21221_),
    .C(_22630_),
    .A(_20310_),
    .Y(_22632_));
 sg13g2_nand3_1 _31194_ (.B(_22631_),
    .C(_22632_),
    .A(net6343),
    .Y(_22633_));
 sg13g2_o21ai_1 _31195_ (.B1(_22633_),
    .Y(_22634_),
    .A1(_22624_),
    .A2(_22625_));
 sg13g2_inv_2 _31196_ (.Y(_22635_),
    .A(_22634_));
 sg13g2_xnor2_1 _31197_ (.Y(_22636_),
    .A(_20508_),
    .B(_22603_));
 sg13g2_nor2_1 _31198_ (.A(\u_inv.f_next[50] ),
    .B(net7386),
    .Y(_22637_));
 sg13g2_a21oi_1 _31199_ (.A1(net7386),
    .A2(_22636_),
    .Y(_22638_),
    .B1(_22637_));
 sg13g2_nor2_1 _31200_ (.A(_20508_),
    .B(_22609_),
    .Y(_22639_));
 sg13g2_nor2_1 _31201_ (.A(net6253),
    .B(_22639_),
    .Y(_22640_));
 sg13g2_a22oi_1 _31202_ (.Y(_22641_),
    .B1(_22640_),
    .B2(_22610_),
    .A2(_22638_),
    .A1(net6253));
 sg13g2_inv_1 _31203_ (.Y(_22642_),
    .A(_22641_));
 sg13g2_xnor2_1 _31204_ (.Y(_22643_),
    .A(_20313_),
    .B(_22621_));
 sg13g2_o21ai_1 _31205_ (.B1(net6250),
    .Y(_22644_),
    .A1(\u_inv.f_next[42] ),
    .A2(net7378));
 sg13g2_a21oi_1 _31206_ (.A1(net7378),
    .A2(_22643_),
    .Y(_22645_),
    .B1(_22644_));
 sg13g2_a21oi_1 _31207_ (.A1(_20312_),
    .A2(_22629_),
    .Y(_22646_),
    .B1(net6250));
 sg13g2_a21o_2 _31208_ (.A2(_22646_),
    .A1(_22630_),
    .B1(_22645_),
    .X(_22647_));
 sg13g2_o21ai_1 _31209_ (.B1(_20501_),
    .Y(_22648_),
    .A1(_20496_),
    .A2(_20502_));
 sg13g2_xnor2_1 _31210_ (.Y(_22649_),
    .A(_20499_),
    .B(_22648_));
 sg13g2_o21ai_1 _31211_ (.B1(net6253),
    .Y(_22650_),
    .A1(\u_inv.f_next[49] ),
    .A2(net7386));
 sg13g2_a21oi_1 _31212_ (.A1(net7386),
    .A2(_22649_),
    .Y(_22651_),
    .B1(_22650_));
 sg13g2_nand3_1 _31213_ (.B(_21230_),
    .C(_21231_),
    .A(_20499_),
    .Y(_22652_));
 sg13g2_nor2_1 _31214_ (.A(net6253),
    .B(_22608_),
    .Y(_22653_));
 sg13g2_a21o_2 _31215_ (.A2(_22653_),
    .A1(_22652_),
    .B1(_22651_),
    .X(_22654_));
 sg13g2_a21oi_1 _31216_ (.A1(_20472_),
    .A2(_20483_),
    .Y(_22655_),
    .B1(_20487_));
 sg13g2_o21ai_1 _31217_ (.B1(_20474_),
    .Y(_22656_),
    .A1(_20475_),
    .A2(_22655_));
 sg13g2_a21oi_1 _31218_ (.A1(_20473_),
    .A2(_22656_),
    .Y(_22657_),
    .B1(net7227));
 sg13g2_o21ai_1 _31219_ (.B1(_22657_),
    .Y(_22658_),
    .A1(_20473_),
    .A2(_22656_));
 sg13g2_o21ai_1 _31220_ (.B1(_22658_),
    .Y(_22659_),
    .A1(\u_inv.f_next[39] ),
    .A2(net7378));
 sg13g2_nand2_1 _31221_ (.Y(_22660_),
    .A(_20478_),
    .B(_21195_));
 sg13g2_a21oi_1 _31222_ (.A1(_21202_),
    .A2(_22660_),
    .Y(_22661_),
    .B1(_20481_));
 sg13g2_o21ai_1 _31223_ (.B1(_20475_),
    .Y(_22662_),
    .A1(_21204_),
    .A2(_22661_));
 sg13g2_nand2b_1 _31224_ (.Y(_22663_),
    .B(_22662_),
    .A_N(_21201_));
 sg13g2_a21oi_1 _31225_ (.A1(_20473_),
    .A2(_22663_),
    .Y(_22664_),
    .B1(net6250));
 sg13g2_o21ai_1 _31226_ (.B1(_22664_),
    .Y(_22665_),
    .A1(_20473_),
    .A2(_22663_));
 sg13g2_o21ai_1 _31227_ (.B1(_22665_),
    .Y(_22666_),
    .A1(net6332),
    .A2(_22659_));
 sg13g2_and2_1 _31228_ (.A(_20557_),
    .B(_22615_),
    .X(_22667_));
 sg13g2_o21ai_1 _31229_ (.B1(net7385),
    .Y(_22668_),
    .A1(_20555_),
    .A2(_22667_));
 sg13g2_a21oi_1 _31230_ (.A1(_20555_),
    .A2(_22667_),
    .Y(_22669_),
    .B1(_22668_));
 sg13g2_o21ai_1 _31231_ (.B1(net6254),
    .Y(_22670_),
    .A1(\u_inv.f_next[57] ),
    .A2(net7385));
 sg13g2_a21oi_1 _31232_ (.A1(_20559_),
    .A2(_21245_),
    .Y(_22671_),
    .B1(_20556_));
 sg13g2_nand2_1 _31233_ (.Y(_22672_),
    .A(_21253_),
    .B(_22671_));
 sg13g2_nand3_1 _31234_ (.B(_22586_),
    .C(_22672_),
    .A(net6347),
    .Y(_22673_));
 sg13g2_o21ai_1 _31235_ (.B1(_22673_),
    .Y(_22674_),
    .A1(_22669_),
    .A2(_22670_));
 sg13g2_o21ai_1 _31236_ (.B1(_20322_),
    .Y(_22675_),
    .A1(_20315_),
    .A2(_22621_));
 sg13g2_a21oi_1 _31237_ (.A1(_20306_),
    .A2(_22675_),
    .Y(_22676_),
    .B1(_20325_));
 sg13g2_xnor2_1 _31238_ (.Y(_22677_),
    .A(_20298_),
    .B(_22676_));
 sg13g2_nor2_1 _31239_ (.A(\u_inv.f_next[46] ),
    .B(net7379),
    .Y(_22678_));
 sg13g2_a21oi_1 _31240_ (.A1(net7378),
    .A2(_22677_),
    .Y(_22679_),
    .B1(_22678_));
 sg13g2_o21ai_1 _31241_ (.B1(_21223_),
    .Y(_22680_),
    .A1(_21208_),
    .A2(_22626_));
 sg13g2_nand2b_1 _31242_ (.Y(_22681_),
    .B(_22680_),
    .A_N(_20301_));
 sg13g2_and2_1 _31243_ (.A(_21224_),
    .B(_22681_),
    .X(_22682_));
 sg13g2_nor2_1 _31244_ (.A(_20304_),
    .B(_22682_),
    .Y(_22683_));
 sg13g2_or3_1 _31245_ (.A(_20298_),
    .B(_21226_),
    .C(_22683_),
    .X(_22684_));
 sg13g2_o21ai_1 _31246_ (.B1(_20298_),
    .Y(_22685_),
    .A1(_21226_),
    .A2(_22683_));
 sg13g2_and2_1 _31247_ (.A(net6343),
    .B(_22685_),
    .X(_22686_));
 sg13g2_a22oi_1 _31248_ (.Y(_22687_),
    .B1(_22684_),
    .B2(_22686_),
    .A2(_22679_),
    .A1(net6250));
 sg13g2_inv_1 _31249_ (.Y(_22688_),
    .A(_22687_));
 sg13g2_a21oi_1 _31250_ (.A1(_20515_),
    .A2(_20525_),
    .Y(_22689_),
    .B1(_20524_));
 sg13g2_xnor2_1 _31251_ (.Y(_22690_),
    .A(_20523_),
    .B(_22689_));
 sg13g2_o21ai_1 _31252_ (.B1(net6254),
    .Y(_22691_),
    .A1(\u_inv.f_next[53] ),
    .A2(net7384));
 sg13g2_a21oi_1 _31253_ (.A1(net7384),
    .A2(_22690_),
    .Y(_22692_),
    .B1(_22691_));
 sg13g2_a21oi_1 _31254_ (.A1(_20522_),
    .A2(_22571_),
    .Y(_22693_),
    .B1(net6254));
 sg13g2_a21oi_1 _31255_ (.A1(_22572_),
    .A2(_22693_),
    .Y(_22694_),
    .B1(_22692_));
 sg13g2_inv_1 _31256_ (.Y(_22695_),
    .A(_22694_));
 sg13g2_xnor2_1 _31257_ (.Y(_22696_),
    .A(_20515_),
    .B(_20525_));
 sg13g2_nor2_1 _31258_ (.A(\u_inv.f_next[52] ),
    .B(net7384),
    .Y(_22697_));
 sg13g2_a21oi_1 _31259_ (.A1(net7384),
    .A2(_22696_),
    .Y(_22698_),
    .B1(_22697_));
 sg13g2_nand3_1 _31260_ (.B(_21233_),
    .C(_21237_),
    .A(_20525_),
    .Y(_22699_));
 sg13g2_nor2_1 _31261_ (.A(net6254),
    .B(_21238_),
    .Y(_22700_));
 sg13g2_a22oi_1 _31262_ (.Y(_22701_),
    .B1(_22699_),
    .B2(_22700_),
    .A2(_22698_),
    .A1(net6253));
 sg13g2_nand2_1 _31263_ (.Y(_22702_),
    .A(_20301_),
    .B(_22675_));
 sg13g2_nand3_1 _31264_ (.B(_20304_),
    .C(_22702_),
    .A(_20300_),
    .Y(_22703_));
 sg13g2_a21o_1 _31265_ (.A2(_22702_),
    .A1(_20300_),
    .B1(_20304_),
    .X(_22704_));
 sg13g2_nand3_1 _31266_ (.B(_22703_),
    .C(_22704_),
    .A(net7379),
    .Y(_22705_));
 sg13g2_a21oi_1 _31267_ (.A1(_18079_),
    .A2(net7227),
    .Y(_22706_),
    .B1(net6343));
 sg13g2_nand2_1 _31268_ (.Y(_22707_),
    .A(_20304_),
    .B(_22682_));
 sg13g2_nor2_1 _31269_ (.A(net6250),
    .B(_22683_),
    .Y(_22708_));
 sg13g2_a22oi_1 _31270_ (.Y(_22709_),
    .B1(_22707_),
    .B2(_22708_),
    .A2(_22706_),
    .A1(_22705_));
 sg13g2_inv_1 _31271_ (.Y(_22710_),
    .A(_22709_));
 sg13g2_a21oi_1 _31272_ (.A1(_20485_),
    .A2(_20488_),
    .Y(_22711_),
    .B1(_20490_));
 sg13g2_a21oi_1 _31273_ (.A1(\u_inv.f_next[40] ),
    .A2(\u_inv.f_reg[40] ),
    .Y(_22712_),
    .B1(_22711_));
 sg13g2_xnor2_1 _31274_ (.Y(_22713_),
    .A(_20491_),
    .B(_22712_));
 sg13g2_nand2_1 _31275_ (.Y(_22714_),
    .A(net7378),
    .B(_22713_));
 sg13g2_o21ai_1 _31276_ (.B1(_22714_),
    .Y(_22715_),
    .A1(\u_inv.f_next[41] ),
    .A2(net7378));
 sg13g2_o21ai_1 _31277_ (.B1(net6343),
    .Y(_22716_),
    .A1(_20491_),
    .A2(_22627_));
 sg13g2_nand2b_1 _31278_ (.Y(_22717_),
    .B(_22628_),
    .A_N(_22716_));
 sg13g2_o21ai_1 _31279_ (.B1(_22717_),
    .Y(_22718_),
    .A1(net6343),
    .A2(_22715_));
 sg13g2_xnor2_1 _31280_ (.Y(_22719_),
    .A(_20496_),
    .B(_20502_));
 sg13g2_o21ai_1 _31281_ (.B1(net6253),
    .Y(_22720_),
    .A1(\u_inv.f_next[48] ),
    .A2(net7386));
 sg13g2_a21oi_1 _31282_ (.A1(net7386),
    .A2(_22719_),
    .Y(_22721_),
    .B1(_22720_));
 sg13g2_xnor2_1 _31283_ (.Y(_22722_),
    .A(_20502_),
    .B(_21229_));
 sg13g2_a21oi_2 _31284_ (.B1(_22721_),
    .Y(_22723_),
    .A2(_22722_),
    .A1(net6343));
 sg13g2_nand2b_1 _31285_ (.Y(_22724_),
    .B(_22723_),
    .A_N(_22718_));
 sg13g2_xnor2_1 _31286_ (.Y(_22725_),
    .A(_20475_),
    .B(_22655_));
 sg13g2_a21oi_1 _31287_ (.A1(net7370),
    .A2(_22725_),
    .Y(_22726_),
    .B1(net6332));
 sg13g2_o21ai_1 _31288_ (.B1(_22726_),
    .Y(_22727_),
    .A1(\u_inv.f_next[38] ),
    .A2(net7370));
 sg13g2_nor3_1 _31289_ (.A(_20475_),
    .B(_21204_),
    .C(_22661_),
    .Y(_22728_));
 sg13g2_nand2_1 _31290_ (.Y(_22729_),
    .A(net6332),
    .B(_22662_));
 sg13g2_o21ai_1 _31291_ (.B1(_22727_),
    .Y(_22730_),
    .A1(_22728_),
    .A2(_22729_));
 sg13g2_xnor2_1 _31292_ (.Y(_22731_),
    .A(_20301_),
    .B(_22680_));
 sg13g2_xnor2_1 _31293_ (.Y(_22732_),
    .A(_20301_),
    .B(_22675_));
 sg13g2_o21ai_1 _31294_ (.B1(net6252),
    .Y(_22733_),
    .A1(\u_inv.f_next[44] ),
    .A2(net7379));
 sg13g2_a21oi_1 _31295_ (.A1(net7379),
    .A2(_22732_),
    .Y(_22734_),
    .B1(_22733_));
 sg13g2_a21oi_2 _31296_ (.B1(_22734_),
    .Y(_22735_),
    .A2(_22731_),
    .A1(net6343));
 sg13g2_inv_1 _31297_ (.Y(_22736_),
    .A(_22735_));
 sg13g2_xnor2_1 _31298_ (.Y(_22737_),
    .A(_20489_),
    .B(_20490_));
 sg13g2_nor2_1 _31299_ (.A(net7227),
    .B(_22737_),
    .Y(_22738_));
 sg13g2_o21ai_1 _31300_ (.B1(net6250),
    .Y(_22739_),
    .A1(\u_inv.f_next[40] ),
    .A2(net7378));
 sg13g2_o21ai_1 _31301_ (.B1(net6343),
    .Y(_22740_),
    .A1(_20490_),
    .A2(_21207_));
 sg13g2_nand2b_1 _31302_ (.Y(_22741_),
    .B(_22626_),
    .A_N(_22740_));
 sg13g2_o21ai_1 _31303_ (.B1(_22741_),
    .Y(_22742_),
    .A1(_22738_),
    .A2(_22739_));
 sg13g2_nand2b_1 _31304_ (.Y(_22743_),
    .B(_20472_),
    .A_N(_20478_));
 sg13g2_nand3_1 _31305_ (.B(_20481_),
    .C(_22743_),
    .A(_20477_),
    .Y(_22744_));
 sg13g2_a21o_1 _31306_ (.A2(_22743_),
    .A1(_20477_),
    .B1(_20481_),
    .X(_22745_));
 sg13g2_nand3_1 _31307_ (.B(_22744_),
    .C(_22745_),
    .A(net7370),
    .Y(_22746_));
 sg13g2_o21ai_1 _31308_ (.B1(net6244),
    .Y(_22747_),
    .A1(\u_inv.f_next[37] ),
    .A2(net7370));
 sg13g2_nand2b_1 _31309_ (.Y(_22748_),
    .B(_22746_),
    .A_N(_22747_));
 sg13g2_nand3_1 _31310_ (.B(_21202_),
    .C(_22660_),
    .A(_20481_),
    .Y(_22749_));
 sg13g2_nand2_1 _31311_ (.Y(_22750_),
    .A(net6333),
    .B(_22749_));
 sg13g2_o21ai_1 _31312_ (.B1(_22748_),
    .Y(_22751_),
    .A1(_22661_),
    .A2(_22750_));
 sg13g2_nand3_1 _31313_ (.B(_20471_),
    .C(_20478_),
    .A(_20465_),
    .Y(_22752_));
 sg13g2_a21oi_1 _31314_ (.A1(_22743_),
    .A2(_22752_),
    .Y(_22753_),
    .B1(net7220));
 sg13g2_o21ai_1 _31315_ (.B1(net6244),
    .Y(_22754_),
    .A1(\u_inv.f_next[36] ),
    .A2(net7370));
 sg13g2_o21ai_1 _31316_ (.B1(net6333),
    .Y(_22755_),
    .A1(_20478_),
    .A2(_21195_));
 sg13g2_nand2b_1 _31317_ (.Y(_22756_),
    .B(_22660_),
    .A_N(_22755_));
 sg13g2_o21ai_1 _31318_ (.B1(_22756_),
    .Y(_22757_),
    .A1(_22753_),
    .A2(_22754_));
 sg13g2_nor2_1 _31319_ (.A(_20453_),
    .B(_20461_),
    .Y(_22758_));
 sg13g2_a21oi_1 _31320_ (.A1(\u_inv.f_next[32] ),
    .A2(\u_inv.f_reg[32] ),
    .Y(_22759_),
    .B1(_22758_));
 sg13g2_xor2_1 _31321_ (.B(_22759_),
    .A(_20460_),
    .X(_22760_));
 sg13g2_o21ai_1 _31322_ (.B1(net6244),
    .Y(_22761_),
    .A1(\u_inv.f_next[33] ),
    .A2(net7369));
 sg13g2_a21o_1 _31323_ (.A2(_22760_),
    .A1(net7369),
    .B1(_22761_),
    .X(_22762_));
 sg13g2_nand3_1 _31324_ (.B(_21188_),
    .C(_21189_),
    .A(_20460_),
    .Y(_22763_));
 sg13g2_a21oi_1 _31325_ (.A1(_21188_),
    .A2(_21189_),
    .Y(_22764_),
    .B1(_20460_));
 sg13g2_nand2_1 _31326_ (.Y(_22765_),
    .A(net6332),
    .B(_22763_));
 sg13g2_o21ai_1 _31327_ (.B1(_22762_),
    .Y(_22766_),
    .A1(_22764_),
    .A2(_22765_));
 sg13g2_nand2_1 _31328_ (.Y(_22767_),
    .A(_20329_),
    .B(_20448_));
 sg13g2_and2_1 _31329_ (.A(_20328_),
    .B(_22767_),
    .X(_22768_));
 sg13g2_xnor2_1 _31330_ (.Y(_22769_),
    .A(_20333_),
    .B(_22768_));
 sg13g2_nor2_1 _31331_ (.A(\u_inv.f_next[31] ),
    .B(net7366),
    .Y(_22770_));
 sg13g2_a21oi_1 _31332_ (.A1(net7366),
    .A2(_22769_),
    .Y(_22771_),
    .B1(_22770_));
 sg13g2_nor2_1 _31333_ (.A(_21178_),
    .B(_21180_),
    .Y(_22772_));
 sg13g2_a21oi_1 _31334_ (.A1(_21179_),
    .A2(_21182_),
    .Y(_22773_),
    .B1(_20329_));
 sg13g2_a21oi_1 _31335_ (.A1(\u_inv.f_next[30] ),
    .A2(_18199_),
    .Y(_22774_),
    .B1(_22773_));
 sg13g2_nand2_1 _31336_ (.Y(_22775_),
    .A(_20332_),
    .B(_22774_));
 sg13g2_nor2_1 _31337_ (.A(_20332_),
    .B(_22774_),
    .Y(_22776_));
 sg13g2_nor2_1 _31338_ (.A(net6242),
    .B(_22776_),
    .Y(_22777_));
 sg13g2_a22oi_1 _31339_ (.Y(_22778_),
    .B1(_22775_),
    .B2(_22777_),
    .A2(_22771_),
    .A1(net6242));
 sg13g2_inv_2 _31340_ (.Y(_22779_),
    .A(_22778_));
 sg13g2_xnor2_1 _31341_ (.Y(_22780_),
    .A(_20462_),
    .B(_21187_));
 sg13g2_a21o_1 _31342_ (.A2(_20461_),
    .A1(_20453_),
    .B1(net7220),
    .X(_22781_));
 sg13g2_a21oi_1 _31343_ (.A1(\u_inv.f_next[32] ),
    .A2(net7220),
    .Y(_22782_),
    .B1(net6332));
 sg13g2_o21ai_1 _31344_ (.B1(_22782_),
    .Y(_22783_),
    .A1(_22758_),
    .A2(_22781_));
 sg13g2_o21ai_1 _31345_ (.B1(_22783_),
    .Y(_22784_),
    .A1(net6244),
    .A2(_22780_));
 sg13g2_xnor2_1 _31346_ (.Y(_22785_),
    .A(_20329_),
    .B(_20448_));
 sg13g2_nor2_1 _31347_ (.A(\u_inv.f_next[30] ),
    .B(net7366),
    .Y(_22786_));
 sg13g2_a21oi_1 _31348_ (.A1(net7366),
    .A2(_22785_),
    .Y(_22787_),
    .B1(_22786_));
 sg13g2_nand3_1 _31349_ (.B(_21179_),
    .C(_21182_),
    .A(_20329_),
    .Y(_22788_));
 sg13g2_nor2_1 _31350_ (.A(net6241),
    .B(_22773_),
    .Y(_22789_));
 sg13g2_a22oi_1 _31351_ (.Y(_22790_),
    .B1(_22788_),
    .B2(_22789_),
    .A2(_22787_),
    .A1(net6242));
 sg13g2_o21ai_1 _31352_ (.B1(_20336_),
    .Y(_22791_),
    .A1(_20442_),
    .A2(_20445_));
 sg13g2_o21ai_1 _31353_ (.B1(net7365),
    .Y(_22792_),
    .A1(_20444_),
    .A2(_22791_));
 sg13g2_a21oi_1 _31354_ (.A1(_20444_),
    .A2(_22791_),
    .Y(_22793_),
    .B1(_22792_));
 sg13g2_o21ai_1 _31355_ (.B1(net6241),
    .Y(_22794_),
    .A1(\u_inv.f_next[29] ),
    .A2(net7365));
 sg13g2_xnor2_1 _31356_ (.Y(_22795_),
    .A(_20444_),
    .B(_22772_));
 sg13g2_nand2_1 _31357_ (.Y(_22796_),
    .A(net6331),
    .B(_22795_));
 sg13g2_o21ai_1 _31358_ (.B1(_22796_),
    .Y(_22797_),
    .A1(_22793_),
    .A2(_22794_));
 sg13g2_a21oi_1 _31359_ (.A1(_20446_),
    .A2(_21177_),
    .Y(_22798_),
    .B1(net6241));
 sg13g2_nor2b_1 _31360_ (.A(_21178_),
    .B_N(_22798_),
    .Y(_22799_));
 sg13g2_xor2_1 _31361_ (.B(_20446_),
    .A(_20442_),
    .X(_22800_));
 sg13g2_o21ai_1 _31362_ (.B1(net6241),
    .Y(_22801_),
    .A1(\u_inv.f_next[28] ),
    .A2(net7365));
 sg13g2_a21oi_1 _31363_ (.A1(net7365),
    .A2(_22800_),
    .Y(_22802_),
    .B1(_22801_));
 sg13g2_or2_1 _31364_ (.X(_22803_),
    .B(_22802_),
    .A(_22799_));
 sg13g2_xor2_1 _31365_ (.B(_20440_),
    .A(_20439_),
    .X(_22804_));
 sg13g2_o21ai_1 _31366_ (.B1(net6236),
    .Y(_22805_),
    .A1(\u_inv.f_next[27] ),
    .A2(net7358));
 sg13g2_a21oi_1 _31367_ (.A1(net7358),
    .A2(_22804_),
    .Y(_22806_),
    .B1(_22805_));
 sg13g2_o21ai_1 _31368_ (.B1(_20440_),
    .Y(_22807_),
    .A1(_20438_),
    .A2(_21171_));
 sg13g2_nand2b_1 _31369_ (.Y(_22808_),
    .B(_21172_),
    .A_N(_22807_));
 sg13g2_o21ai_1 _31370_ (.B1(net6321),
    .Y(_22809_),
    .A1(_20440_),
    .A2(_21172_));
 sg13g2_nor2_1 _31371_ (.A(_21175_),
    .B(_22809_),
    .Y(_22810_));
 sg13g2_a21o_2 _31372_ (.A2(_22810_),
    .A1(_22808_),
    .B1(_22806_),
    .X(_22811_));
 sg13g2_xnor2_1 _31373_ (.Y(_22812_),
    .A(_20438_),
    .B(_21171_));
 sg13g2_a21oi_1 _31374_ (.A1(_20437_),
    .A2(_20438_),
    .Y(_22813_),
    .B1(net7212));
 sg13g2_o21ai_1 _31375_ (.B1(_22813_),
    .Y(_22814_),
    .A1(_20437_),
    .A2(_20438_));
 sg13g2_a21oi_1 _31376_ (.A1(\u_inv.f_next[26] ),
    .A2(net7212),
    .Y(_22815_),
    .B1(net6321));
 sg13g2_a22oi_1 _31377_ (.Y(_22816_),
    .B1(_22814_),
    .B2(_22815_),
    .A2(_22812_),
    .A1(net6321));
 sg13g2_nand3_1 _31378_ (.B(_20432_),
    .C(_20435_),
    .A(_20344_),
    .Y(_22817_));
 sg13g2_a21oi_1 _31379_ (.A1(_20344_),
    .A2(_20432_),
    .Y(_22818_),
    .B1(_20435_));
 sg13g2_nor2_1 _31380_ (.A(net7213),
    .B(_22818_),
    .Y(_22819_));
 sg13g2_a221oi_1 _31381_ (.B2(_22819_),
    .C1(net6318),
    .B1(_22817_),
    .A1(_18087_),
    .Y(_22820_),
    .A2(net7213));
 sg13g2_or3_1 _31382_ (.A(_20434_),
    .B(_21167_),
    .C(_21168_),
    .X(_22821_));
 sg13g2_nand3_1 _31383_ (.B(_21169_),
    .C(_22821_),
    .A(net6318),
    .Y(_22822_));
 sg13g2_nand2b_2 _31384_ (.Y(_22823_),
    .B(_22822_),
    .A_N(_22820_));
 sg13g2_a21oi_1 _31385_ (.A1(_20418_),
    .A2(_20422_),
    .Y(_22824_),
    .B1(_20428_));
 sg13g2_nor2_1 _31386_ (.A(_20346_),
    .B(_22824_),
    .Y(_22825_));
 sg13g2_a21oi_1 _31387_ (.A1(\u_inv.f_next[22] ),
    .A2(\u_inv.f_reg[22] ),
    .Y(_22826_),
    .B1(_22825_));
 sg13g2_o21ai_1 _31388_ (.B1(net7353),
    .Y(_22827_),
    .A1(_20348_),
    .A2(_22826_));
 sg13g2_a21oi_1 _31389_ (.A1(_20348_),
    .A2(_22826_),
    .Y(_22828_),
    .B1(_22827_));
 sg13g2_o21ai_1 _31390_ (.B1(net6232),
    .Y(_22829_),
    .A1(\u_inv.f_next[23] ),
    .A2(net7353));
 sg13g2_nor2_1 _31391_ (.A(_20345_),
    .B(_21160_),
    .Y(_22830_));
 sg13g2_a21oi_1 _31392_ (.A1(\u_inv.f_next[22] ),
    .A2(_18198_),
    .Y(_22831_),
    .B1(_22830_));
 sg13g2_a21oi_1 _31393_ (.A1(_20348_),
    .A2(_22831_),
    .Y(_22832_),
    .B1(net6232));
 sg13g2_o21ai_1 _31394_ (.B1(_22832_),
    .Y(_22833_),
    .A1(_20348_),
    .A2(_22831_));
 sg13g2_o21ai_1 _31395_ (.B1(_22833_),
    .Y(_22834_),
    .A1(_22828_),
    .A2(_22829_));
 sg13g2_nand3_1 _31396_ (.B(_21164_),
    .C(_21166_),
    .A(_20431_),
    .Y(_22835_));
 sg13g2_nor2_1 _31397_ (.A(net6232),
    .B(_21167_),
    .Y(_22836_));
 sg13g2_xnor2_1 _31398_ (.Y(_22837_),
    .A(_20430_),
    .B(_20431_));
 sg13g2_nor2_1 _31399_ (.A(\u_inv.f_next[24] ),
    .B(net7353),
    .Y(_22838_));
 sg13g2_a21oi_1 _31400_ (.A1(net7353),
    .A2(_22837_),
    .Y(_22839_),
    .B1(_22838_));
 sg13g2_a22oi_1 _31401_ (.Y(_22840_),
    .B1(_22839_),
    .B2(net6232),
    .A2(_22836_),
    .A1(_22835_));
 sg13g2_nand2_1 _31402_ (.Y(_22841_),
    .A(_20345_),
    .B(_21160_));
 sg13g2_nor2_1 _31403_ (.A(net6225),
    .B(_22830_),
    .Y(_22842_));
 sg13g2_xnor2_1 _31404_ (.Y(_22843_),
    .A(_20346_),
    .B(_22824_));
 sg13g2_nor2_1 _31405_ (.A(\u_inv.f_next[22] ),
    .B(net7343),
    .Y(_22844_));
 sg13g2_a21oi_1 _31406_ (.A1(net7343),
    .A2(_22843_),
    .Y(_22845_),
    .B1(_22844_));
 sg13g2_a22oi_1 _31407_ (.Y(_22846_),
    .B1(_22845_),
    .B2(net6225),
    .A2(_22842_),
    .A1(_22841_));
 sg13g2_inv_1 _31408_ (.Y(_22847_),
    .A(_22846_));
 sg13g2_nand3_1 _31409_ (.B(_21153_),
    .C(_21156_),
    .A(_20421_),
    .Y(_22848_));
 sg13g2_nor2_1 _31410_ (.A(net6225),
    .B(_21157_),
    .Y(_22849_));
 sg13g2_xor2_1 _31411_ (.B(_20421_),
    .A(_20417_),
    .X(_22850_));
 sg13g2_o21ai_1 _31412_ (.B1(net6225),
    .Y(_22851_),
    .A1(\u_inv.f_next[20] ),
    .A2(net7343));
 sg13g2_a21oi_1 _31413_ (.A1(net7343),
    .A2(_22850_),
    .Y(_22852_),
    .B1(_22851_));
 sg13g2_a21o_2 _31414_ (.A2(_22849_),
    .A1(_22848_),
    .B1(_22852_),
    .X(_22853_));
 sg13g2_o21ai_1 _31415_ (.B1(net7343),
    .Y(_22854_),
    .A1(_20412_),
    .A2(_20414_));
 sg13g2_a21oi_1 _31416_ (.A1(_20412_),
    .A2(_20414_),
    .Y(_22855_),
    .B1(_22854_));
 sg13g2_o21ai_1 _31417_ (.B1(net6225),
    .Y(_22856_),
    .A1(net7300),
    .A2(net7343));
 sg13g2_or2_1 _31418_ (.X(_22857_),
    .B(_21150_),
    .A(_20415_));
 sg13g2_nand3_1 _31419_ (.B(_21154_),
    .C(_22857_),
    .A(net6309),
    .Y(_22858_));
 sg13g2_o21ai_1 _31420_ (.B1(_22858_),
    .Y(_22859_),
    .A1(_22855_),
    .A2(_22856_));
 sg13g2_xnor2_1 _31421_ (.Y(_22860_),
    .A(_20411_),
    .B(_21148_));
 sg13g2_xor2_1 _31422_ (.B(_20411_),
    .A(_20410_),
    .X(_22861_));
 sg13g2_nand2_1 _31423_ (.Y(_22862_),
    .A(net7343),
    .B(_22861_));
 sg13g2_a21oi_1 _31424_ (.A1(\u_inv.f_next[18] ),
    .A2(net7203),
    .Y(_22863_),
    .B1(net6309));
 sg13g2_a22oi_1 _31425_ (.Y(_22864_),
    .B1(_22862_),
    .B2(_22863_),
    .A2(_22860_),
    .A1(net6309));
 sg13g2_xor2_1 _31426_ (.B(_20407_),
    .A(_20405_),
    .X(_22865_));
 sg13g2_o21ai_1 _31427_ (.B1(net6223),
    .Y(_22866_),
    .A1(\u_inv.f_next[17] ),
    .A2(net7339));
 sg13g2_a21oi_1 _31428_ (.A1(net7339),
    .A2(_22865_),
    .Y(_22867_),
    .B1(_22866_));
 sg13g2_a21oi_1 _31429_ (.A1(_20407_),
    .A2(_21144_),
    .Y(_22868_),
    .B1(net6223));
 sg13g2_o21ai_1 _31430_ (.B1(_22868_),
    .Y(_22869_),
    .A1(_20407_),
    .A2(_21144_));
 sg13g2_nand2b_2 _31431_ (.Y(_22870_),
    .B(_22869_),
    .A_N(_22867_));
 sg13g2_xnor2_1 _31432_ (.Y(_22871_),
    .A(_20404_),
    .B(_21142_));
 sg13g2_xnor2_1 _31433_ (.Y(_22872_),
    .A(_20403_),
    .B(_20404_));
 sg13g2_o21ai_1 _31434_ (.B1(net6223),
    .Y(_22873_),
    .A1(\u_inv.f_next[16] ),
    .A2(net7339));
 sg13g2_a21o_1 _31435_ (.A2(_22872_),
    .A1(net7339),
    .B1(_22873_),
    .X(_22874_));
 sg13g2_o21ai_1 _31436_ (.B1(_22874_),
    .Y(_22875_),
    .A1(net6223),
    .A2(_22871_));
 sg13g2_nand2_2 _31437_ (.Y(_22876_),
    .A(_20357_),
    .B(_20358_));
 sg13g2_a21oi_1 _31438_ (.A1(_20401_),
    .A2(_22876_),
    .Y(_22877_),
    .B1(net7197));
 sg13g2_o21ai_1 _31439_ (.B1(_22877_),
    .Y(_22878_),
    .A1(_20401_),
    .A2(_22876_));
 sg13g2_o21ai_1 _31440_ (.B1(_22878_),
    .Y(_22879_),
    .A1(\u_inv.f_next[15] ),
    .A2(net7329));
 sg13g2_a21oi_1 _31441_ (.A1(_21140_),
    .A2(_22876_),
    .Y(_22880_),
    .B1(net6218));
 sg13g2_o21ai_1 _31442_ (.B1(_22880_),
    .Y(_22881_),
    .A1(_21140_),
    .A2(_22876_));
 sg13g2_o21ai_1 _31443_ (.B1(_22881_),
    .Y(_22882_),
    .A1(net6298),
    .A2(_22879_));
 sg13g2_nor3_1 _31444_ (.A(_20360_),
    .B(_21136_),
    .C(_21137_),
    .Y(_22883_));
 sg13g2_nand2_1 _31445_ (.Y(_22884_),
    .A(net6298),
    .B(_21138_));
 sg13g2_xnor2_1 _31446_ (.Y(_22885_),
    .A(_20360_),
    .B(_20399_));
 sg13g2_o21ai_1 _31447_ (.B1(net6217),
    .Y(_22886_),
    .A1(\u_inv.f_next[14] ),
    .A2(net7328));
 sg13g2_a21o_1 _31448_ (.A2(_22885_),
    .A1(net7328),
    .B1(_22886_),
    .X(_22887_));
 sg13g2_o21ai_1 _31449_ (.B1(_22887_),
    .Y(_22888_),
    .A1(_22883_),
    .A2(_22884_));
 sg13g2_xnor2_1 _31450_ (.Y(_22889_),
    .A(_20397_),
    .B(_21111_));
 sg13g2_o21ai_1 _31451_ (.B1(net6213),
    .Y(_22890_),
    .A1(\u_inv.f_next[13] ),
    .A2(net7325));
 sg13g2_a21oi_1 _31452_ (.A1(net7325),
    .A2(_22889_),
    .Y(_22891_),
    .B1(_22890_));
 sg13g2_nand3_1 _31453_ (.B(_21134_),
    .C(_21135_),
    .A(_21111_),
    .Y(_22892_));
 sg13g2_nor2_1 _31454_ (.A(net6213),
    .B(_21136_),
    .Y(_22893_));
 sg13g2_a21o_2 _31455_ (.A2(_22893_),
    .A1(_22892_),
    .B1(_22891_),
    .X(_22894_));
 sg13g2_nor3_1 _31456_ (.A(_20365_),
    .B(_21132_),
    .C(_21133_),
    .Y(_22895_));
 sg13g2_nor2_1 _31457_ (.A(net6213),
    .B(_22895_),
    .Y(_22896_));
 sg13g2_xnor2_1 _31458_ (.Y(_22897_),
    .A(_20364_),
    .B(_20395_));
 sg13g2_nor2_1 _31459_ (.A(\u_inv.f_next[12] ),
    .B(net7325),
    .Y(_22898_));
 sg13g2_a21oi_1 _31460_ (.A1(net7325),
    .A2(_22897_),
    .Y(_22899_),
    .B1(_22898_));
 sg13g2_a22oi_1 _31461_ (.Y(_22900_),
    .B1(_22899_),
    .B2(net6213),
    .A2(_22896_),
    .A1(_21134_));
 sg13g2_inv_1 _31462_ (.Y(_22901_),
    .A(_22900_));
 sg13g2_xnor2_1 _31463_ (.Y(_22902_),
    .A(_20393_),
    .B(_21112_));
 sg13g2_o21ai_1 _31464_ (.B1(net6215),
    .Y(_22903_),
    .A1(\u_inv.f_next[11] ),
    .A2(net7324));
 sg13g2_a21oi_1 _31465_ (.A1(net7324),
    .A2(_22902_),
    .Y(_22904_),
    .B1(_22903_));
 sg13g2_nand3_1 _31466_ (.B(_21130_),
    .C(_21131_),
    .A(_21112_),
    .Y(_22905_));
 sg13g2_nor2_1 _31467_ (.A(net6215),
    .B(_21132_),
    .Y(_22906_));
 sg13g2_a21oi_2 _31468_ (.B1(_22904_),
    .Y(_22907_),
    .A2(_22906_),
    .A1(_22905_));
 sg13g2_nand3_1 _31469_ (.B(_21128_),
    .C(_21129_),
    .A(_20369_),
    .Y(_22908_));
 sg13g2_and2_1 _31470_ (.A(net6297),
    .B(_22908_),
    .X(_22909_));
 sg13g2_xnor2_1 _31471_ (.Y(_22910_),
    .A(_20369_),
    .B(_20391_));
 sg13g2_nor2_1 _31472_ (.A(\u_inv.f_next[10] ),
    .B(net7324),
    .Y(_22911_));
 sg13g2_a21oi_1 _31473_ (.A1(net7324),
    .A2(_22910_),
    .Y(_22912_),
    .B1(_22911_));
 sg13g2_a22oi_1 _31474_ (.Y(_22913_),
    .B1(_22912_),
    .B2(net6215),
    .A2(_22909_),
    .A1(_21130_));
 sg13g2_xnor2_1 _31475_ (.Y(_22914_),
    .A(_20389_),
    .B(_21114_));
 sg13g2_o21ai_1 _31476_ (.B1(net6215),
    .Y(_22915_),
    .A1(\u_inv.f_next[9] ),
    .A2(net7317));
 sg13g2_a21o_1 _31477_ (.A2(_22914_),
    .A1(net7317),
    .B1(_22915_),
    .X(_22916_));
 sg13g2_nor3_1 _31478_ (.A(_21114_),
    .B(_21126_),
    .C(_21127_),
    .Y(_22917_));
 sg13g2_nand2_1 _31479_ (.Y(_22918_),
    .A(net6287),
    .B(_21128_));
 sg13g2_o21ai_1 _31480_ (.B1(_22916_),
    .Y(_22919_),
    .A1(_22917_),
    .A2(_22918_));
 sg13g2_nand3_1 _31481_ (.B(_21124_),
    .C(_21125_),
    .A(_20372_),
    .Y(_22920_));
 sg13g2_nand2_1 _31482_ (.Y(_22921_),
    .A(net6287),
    .B(_22920_));
 sg13g2_xnor2_1 _31483_ (.Y(_22922_),
    .A(_20372_),
    .B(_20388_));
 sg13g2_o21ai_1 _31484_ (.B1(net6208),
    .Y(_22923_),
    .A1(\u_inv.f_next[8] ),
    .A2(net7317));
 sg13g2_a21o_1 _31485_ (.A2(_22922_),
    .A1(net7317),
    .B1(_22923_),
    .X(_22924_));
 sg13g2_o21ai_1 _31486_ (.B1(_22924_),
    .Y(_22925_),
    .A1(_21126_),
    .A2(_22921_));
 sg13g2_or3_1 _31487_ (.A(_20374_),
    .B(_21122_),
    .C(_21123_),
    .X(_22926_));
 sg13g2_nand2_1 _31488_ (.Y(_22927_),
    .A(_21124_),
    .B(_22926_));
 sg13g2_o21ai_1 _31489_ (.B1(net7318),
    .Y(_22928_),
    .A1(_20374_),
    .A2(_20387_));
 sg13g2_a21o_1 _31490_ (.A2(_20387_),
    .A1(_20374_),
    .B1(_22928_),
    .X(_22929_));
 sg13g2_a21oi_1 _31491_ (.A1(\u_inv.f_next[7] ),
    .A2(net7186),
    .Y(_22930_),
    .B1(net6286));
 sg13g2_a22oi_1 _31492_ (.Y(_22931_),
    .B1(_22929_),
    .B2(_22930_),
    .A2(_22927_),
    .A1(net6286));
 sg13g2_nand3_1 _31493_ (.B(_21120_),
    .C(_21121_),
    .A(_20376_),
    .Y(_22932_));
 sg13g2_nand2b_1 _31494_ (.Y(_22933_),
    .B(_22932_),
    .A_N(_21122_));
 sg13g2_a21oi_1 _31495_ (.A1(_20376_),
    .A2(_20386_),
    .Y(_22934_),
    .B1(net7186));
 sg13g2_o21ai_1 _31496_ (.B1(_22934_),
    .Y(_22935_),
    .A1(_20376_),
    .A2(_20386_));
 sg13g2_a21oi_1 _31497_ (.A1(\u_inv.f_next[6] ),
    .A2(net7186),
    .Y(_22936_),
    .B1(net6286));
 sg13g2_a22oi_1 _31498_ (.Y(_22937_),
    .B1(_22935_),
    .B2(_22936_),
    .A2(_22933_),
    .A1(net6286));
 sg13g2_or3_1 _31499_ (.A(_20378_),
    .B(_21118_),
    .C(_21119_),
    .X(_22938_));
 sg13g2_nand3_1 _31500_ (.B(_21120_),
    .C(_22938_),
    .A(net6286),
    .Y(_22939_));
 sg13g2_xor2_1 _31501_ (.B(_20385_),
    .A(_20378_),
    .X(_22940_));
 sg13g2_nor2_1 _31502_ (.A(net7186),
    .B(_22940_),
    .Y(_22941_));
 sg13g2_o21ai_1 _31503_ (.B1(net6207),
    .Y(_22942_),
    .A1(\u_inv.f_next[5] ),
    .A2(net7318));
 sg13g2_o21ai_1 _31504_ (.B1(_22939_),
    .Y(_22943_),
    .A1(_22941_),
    .A2(_22942_));
 sg13g2_nand3_1 _31505_ (.B(_21116_),
    .C(_21117_),
    .A(_20380_),
    .Y(_22944_));
 sg13g2_nand2b_1 _31506_ (.Y(_22945_),
    .B(_22944_),
    .A_N(_21118_));
 sg13g2_xor2_1 _31507_ (.B(_20384_),
    .A(_20380_),
    .X(_22946_));
 sg13g2_nand2_1 _31508_ (.Y(_22947_),
    .A(net7314),
    .B(_22946_));
 sg13g2_a21oi_1 _31509_ (.A1(\u_inv.f_next[4] ),
    .A2(net7185),
    .Y(_22948_),
    .B1(net6283));
 sg13g2_a22oi_1 _31510_ (.Y(_22949_),
    .B1(_22947_),
    .B2(_22948_),
    .A2(_22945_),
    .A1(net6283));
 sg13g2_nand2_1 _31511_ (.Y(_22950_),
    .A(\u_inv.f_reg[0] ),
    .B(net6284));
 sg13g2_a21oi_1 _31512_ (.A1(_18183_),
    .A2(_19834_),
    .Y(_22951_),
    .B1(net7184));
 sg13g2_o21ai_1 _31513_ (.B1(_22951_),
    .Y(_22952_),
    .A1(_19834_),
    .A2(_19835_));
 sg13g2_o21ai_1 _31514_ (.B1(_22952_),
    .Y(_22953_),
    .A1(_18098_),
    .A2(net7315));
 sg13g2_xor2_1 _31515_ (.B(_22953_),
    .A(_22950_),
    .X(_22954_));
 sg13g2_or3_1 _31516_ (.A(_19830_),
    .B(_20382_),
    .C(_21115_),
    .X(_22955_));
 sg13g2_nand2_1 _31517_ (.Y(_22956_),
    .A(_21116_),
    .B(_22955_));
 sg13g2_xor2_1 _31518_ (.B(_20383_),
    .A(_20382_),
    .X(_22957_));
 sg13g2_nand2_1 _31519_ (.Y(_22958_),
    .A(net7314),
    .B(_22957_));
 sg13g2_a21oi_1 _31520_ (.A1(\u_inv.f_next[3] ),
    .A2(net7184),
    .Y(_22959_),
    .B1(net6283));
 sg13g2_a22oi_1 _31521_ (.Y(_22960_),
    .B1(_22958_),
    .B2(_22959_),
    .A2(_22956_),
    .A1(net6283));
 sg13g2_nand3b_1 _31522_ (.B(_19841_),
    .C(_22954_),
    .Y(_22961_),
    .A_N(_22960_));
 sg13g2_or4_1 _31523_ (.A(_22937_),
    .B(_22943_),
    .C(_22949_),
    .D(_22961_),
    .X(_22962_));
 sg13g2_nor4_1 _31524_ (.A(_22919_),
    .B(_22925_),
    .C(_22931_),
    .D(_22962_),
    .Y(_22963_));
 sg13g2_nand4_1 _31525_ (.B(_22907_),
    .C(_22913_),
    .A(_22900_),
    .Y(_22964_),
    .D(_22963_));
 sg13g2_or4_1 _31526_ (.A(_22882_),
    .B(_22888_),
    .C(_22894_),
    .D(_22964_),
    .X(_22965_));
 sg13g2_or4_1 _31527_ (.A(_22864_),
    .B(_22870_),
    .C(_22875_),
    .D(_22965_),
    .X(_22966_));
 sg13g2_nor3_1 _31528_ (.A(_22853_),
    .B(_22859_),
    .C(_22966_),
    .Y(_22967_));
 sg13g2_a21oi_1 _31529_ (.A1(_20418_),
    .A2(_20421_),
    .Y(_22968_),
    .B1(_20420_));
 sg13g2_xor2_1 _31530_ (.B(_22968_),
    .A(_20419_),
    .X(_22969_));
 sg13g2_o21ai_1 _31531_ (.B1(net6225),
    .Y(_22970_),
    .A1(\u_inv.f_next[21] ),
    .A2(net7345));
 sg13g2_a21oi_1 _31532_ (.A1(net7345),
    .A2(_22969_),
    .Y(_22971_),
    .B1(_22970_));
 sg13g2_o21ai_1 _31533_ (.B1(net6309),
    .Y(_22972_),
    .A1(_20419_),
    .A2(_21158_));
 sg13g2_a21oi_1 _31534_ (.A1(_20419_),
    .A2(_21158_),
    .Y(_22973_),
    .B1(_22972_));
 sg13g2_nor2_2 _31535_ (.A(_22971_),
    .B(_22973_),
    .Y(_22974_));
 sg13g2_nand4_1 _31536_ (.B(_22846_),
    .C(_22967_),
    .A(_22840_),
    .Y(_22975_),
    .D(_22974_));
 sg13g2_or4_1 _31537_ (.A(_22816_),
    .B(_22823_),
    .C(_22834_),
    .D(_22975_),
    .X(_22976_));
 sg13g2_nor4_1 _31538_ (.A(_22797_),
    .B(_22803_),
    .C(_22811_),
    .D(_22976_),
    .Y(_22977_));
 sg13g2_nand4_1 _31539_ (.B(_22784_),
    .C(_22790_),
    .A(_22778_),
    .Y(_22978_),
    .D(_22977_));
 sg13g2_nor3_1 _31540_ (.A(_22757_),
    .B(_22766_),
    .C(_22978_),
    .Y(_22979_));
 sg13g2_a21oi_1 _31541_ (.A1(\u_inv.f_next[33] ),
    .A2(_18201_),
    .Y(_22980_),
    .B1(_22764_));
 sg13g2_or2_1 _31542_ (.X(_22981_),
    .B(_22980_),
    .A(_20455_));
 sg13g2_a21oi_1 _31543_ (.A1(_20455_),
    .A2(_22980_),
    .Y(_22982_),
    .B1(net6244));
 sg13g2_o21ai_1 _31544_ (.B1(_20469_),
    .Y(_22983_),
    .A1(_20453_),
    .A2(_20463_));
 sg13g2_nand2_1 _31545_ (.Y(_22984_),
    .A(_20455_),
    .B(_22983_));
 sg13g2_xnor2_1 _31546_ (.Y(_22985_),
    .A(_20455_),
    .B(_22983_));
 sg13g2_o21ai_1 _31547_ (.B1(net6244),
    .Y(_22986_),
    .A1(\u_inv.f_next[34] ),
    .A2(net7369));
 sg13g2_a21oi_1 _31548_ (.A1(net7369),
    .A2(_22985_),
    .Y(_22987_),
    .B1(_22986_));
 sg13g2_a21o_2 _31549_ (.A2(_22982_),
    .A1(_22981_),
    .B1(_22987_),
    .X(_22988_));
 sg13g2_nor3_1 _31550_ (.A(_22742_),
    .B(_22751_),
    .C(_22988_),
    .Y(_22989_));
 sg13g2_a21o_1 _31551_ (.A2(_22984_),
    .A1(_20454_),
    .B1(_20458_),
    .X(_22990_));
 sg13g2_nand3_1 _31552_ (.B(_20458_),
    .C(_22984_),
    .A(_20454_),
    .Y(_22991_));
 sg13g2_nand3_1 _31553_ (.B(_22990_),
    .C(_22991_),
    .A(net7369),
    .Y(_22992_));
 sg13g2_o21ai_1 _31554_ (.B1(_22992_),
    .Y(_22993_),
    .A1(\u_inv.f_next[35] ),
    .A2(net7370));
 sg13g2_and3_1 _31555_ (.X(_22994_),
    .A(_20458_),
    .B(_21100_),
    .C(_22981_));
 sg13g2_a21oi_1 _31556_ (.A1(_21100_),
    .A2(_22981_),
    .Y(_22995_),
    .B1(_20458_));
 sg13g2_or3_1 _31557_ (.A(net6246),
    .B(_22994_),
    .C(_22995_),
    .X(_22996_));
 sg13g2_o21ai_1 _31558_ (.B1(_22996_),
    .Y(_22997_),
    .A1(net6332),
    .A2(_22993_));
 sg13g2_o21ai_1 _31559_ (.B1(_20297_),
    .Y(_22998_),
    .A1(_20298_),
    .A2(_22676_));
 sg13g2_a21oi_1 _31560_ (.A1(_20296_),
    .A2(_22998_),
    .Y(_22999_),
    .B1(net7227));
 sg13g2_o21ai_1 _31561_ (.B1(_22999_),
    .Y(_23000_),
    .A1(_20296_),
    .A2(_22998_));
 sg13g2_a21oi_1 _31562_ (.A1(_18078_),
    .A2(net7227),
    .Y(_23001_),
    .B1(net6346));
 sg13g2_nand2_1 _31563_ (.Y(_23002_),
    .A(_23000_),
    .B(_23001_));
 sg13g2_nand2b_1 _31564_ (.Y(_23003_),
    .B(_22685_),
    .A_N(_21214_));
 sg13g2_xnor2_1 _31565_ (.Y(_23004_),
    .A(_20296_),
    .B(_23003_));
 sg13g2_o21ai_1 _31566_ (.B1(_23002_),
    .Y(_23005_),
    .A1(net6250),
    .A2(_23004_));
 sg13g2_xor2_1 _31567_ (.B(_22577_),
    .A(_20518_),
    .X(_23006_));
 sg13g2_o21ai_1 _31568_ (.B1(net6254),
    .Y(_23007_),
    .A1(\u_inv.f_next[54] ),
    .A2(net7384));
 sg13g2_a21o_1 _31569_ (.A2(_23006_),
    .A1(net7384),
    .B1(_23007_),
    .X(_23008_));
 sg13g2_nand3_1 _31570_ (.B(_21094_),
    .C(_22572_),
    .A(_20518_),
    .Y(_23009_));
 sg13g2_nand2_1 _31571_ (.Y(_23010_),
    .A(net6347),
    .B(_23009_));
 sg13g2_o21ai_1 _31572_ (.B1(_23008_),
    .Y(_23011_),
    .A1(_22573_),
    .A2(_23010_));
 sg13g2_a21oi_1 _31573_ (.A1(_20538_),
    .A2(_22528_),
    .Y(_23012_),
    .B1(_20537_));
 sg13g2_or2_1 _31574_ (.X(_23013_),
    .B(_23012_),
    .A(_20536_));
 sg13g2_a21oi_1 _31575_ (.A1(_20536_),
    .A2(_23012_),
    .Y(_23014_),
    .B1(net7237));
 sg13g2_a221oi_1 _31576_ (.B2(_23014_),
    .C1(net6361),
    .B1(_23013_),
    .A1(_18071_),
    .Y(_23015_),
    .A2(net7237));
 sg13g2_a21oi_1 _31577_ (.A1(_20536_),
    .A2(_22537_),
    .Y(_23016_),
    .B1(net6260));
 sg13g2_a21oi_2 _31578_ (.B1(_23015_),
    .Y(_23017_),
    .A2(_23016_),
    .A1(_22538_));
 sg13g2_a21oi_1 _31579_ (.A1(_20550_),
    .A2(_22587_),
    .Y(_23018_),
    .B1(_20549_));
 sg13g2_a21oi_1 _31580_ (.A1(_20548_),
    .A2(_23018_),
    .Y(_23019_),
    .B1(net6254));
 sg13g2_o21ai_1 _31581_ (.B1(_23019_),
    .Y(_23020_),
    .A1(_20548_),
    .A2(_23018_));
 sg13g2_o21ai_1 _31582_ (.B1(_20565_),
    .Y(_23021_),
    .A1(_20550_),
    .A2(_22527_));
 sg13g2_xnor2_1 _31583_ (.Y(_23022_),
    .A(_20548_),
    .B(_23021_));
 sg13g2_a21oi_1 _31584_ (.A1(net7384),
    .A2(_23022_),
    .Y(_23023_),
    .B1(net6347));
 sg13g2_o21ai_1 _31585_ (.B1(_23023_),
    .Y(_23024_),
    .A1(\u_inv.f_next[59] ),
    .A2(net7385));
 sg13g2_nand2_2 _31586_ (.Y(_23025_),
    .A(_23020_),
    .B(_23024_));
 sg13g2_a21oi_1 _31587_ (.A1(_20608_),
    .A2(_20612_),
    .Y(_23026_),
    .B1(_20637_));
 sg13g2_nor2_2 _31588_ (.A(_20642_),
    .B(_23026_),
    .Y(_23027_));
 sg13g2_xnor2_1 _31589_ (.Y(_23028_),
    .A(_20632_),
    .B(_23027_));
 sg13g2_nor2_1 _31590_ (.A(\u_inv.f_next[74] ),
    .B(net7400),
    .Y(_23029_));
 sg13g2_a21oi_1 _31591_ (.A1(net7400),
    .A2(_23028_),
    .Y(_23030_),
    .B1(_23029_));
 sg13g2_a21o_1 _31592_ (.A2(_21287_),
    .A1(_21279_),
    .B1(_21289_),
    .X(_23031_));
 sg13g2_nand3_1 _31593_ (.B(_21297_),
    .C(_23031_),
    .A(_20631_),
    .Y(_23032_));
 sg13g2_a21oi_1 _31594_ (.A1(_21297_),
    .A2(_23031_),
    .Y(_23033_),
    .B1(_20631_));
 sg13g2_nor2_1 _31595_ (.A(net6262),
    .B(_23033_),
    .Y(_23034_));
 sg13g2_a22oi_1 _31596_ (.Y(_23035_),
    .B1(_23032_),
    .B2(_23034_),
    .A2(_23030_),
    .A1(net6262));
 sg13g2_xnor2_1 _31597_ (.Y(_23036_),
    .A(_20613_),
    .B(_20636_));
 sg13g2_or2_1 _31598_ (.X(_23037_),
    .B(net7400),
    .A(\u_inv.f_next[72] ));
 sg13g2_a21oi_1 _31599_ (.A1(net7400),
    .A2(_23036_),
    .Y(_23038_),
    .B1(net6357));
 sg13g2_xor2_1 _31600_ (.B(_21288_),
    .A(_20636_),
    .X(_23039_));
 sg13g2_a22oi_1 _31601_ (.Y(_23040_),
    .B1(_23039_),
    .B2(net6357),
    .A2(_23038_),
    .A1(_23037_));
 sg13g2_inv_1 _31602_ (.Y(_23041_),
    .A(_23040_));
 sg13g2_and2_1 _31603_ (.A(_20634_),
    .B(_21295_),
    .X(_23042_));
 sg13g2_o21ai_1 _31604_ (.B1(_23042_),
    .Y(_23043_),
    .A1(_20636_),
    .A2(_21288_));
 sg13g2_nor2_1 _31605_ (.A(net6262),
    .B(_21296_),
    .Y(_23044_));
 sg13g2_and2_1 _31606_ (.A(_23031_),
    .B(_23044_),
    .X(_23045_));
 sg13g2_a21oi_1 _31607_ (.A1(_20613_),
    .A2(_20636_),
    .Y(_23046_),
    .B1(_20635_));
 sg13g2_xor2_1 _31608_ (.B(_23046_),
    .A(_20634_),
    .X(_23047_));
 sg13g2_o21ai_1 _31609_ (.B1(net6262),
    .Y(_23048_),
    .A1(\u_inv.f_next[73] ),
    .A2(net7400));
 sg13g2_a21oi_1 _31610_ (.A1(net7400),
    .A2(_23047_),
    .Y(_23049_),
    .B1(_23048_));
 sg13g2_a21o_2 _31611_ (.A2(_23045_),
    .A1(_23043_),
    .B1(_23049_),
    .X(_23050_));
 sg13g2_or3_1 _31612_ (.A(_20576_),
    .B(_20584_),
    .C(_20586_),
    .X(_23051_));
 sg13g2_a21o_1 _31613_ (.A2(_23051_),
    .A1(_20591_),
    .B1(_20579_),
    .X(_23052_));
 sg13g2_nand3_1 _31614_ (.B(_20591_),
    .C(_23051_),
    .A(_20579_),
    .Y(_23053_));
 sg13g2_nand3_1 _31615_ (.B(_23052_),
    .C(_23053_),
    .A(net7396),
    .Y(_23054_));
 sg13g2_o21ai_1 _31616_ (.B1(_23054_),
    .Y(_23055_),
    .A1(_18069_),
    .A2(net7395));
 sg13g2_a21oi_1 _31617_ (.A1(_20584_),
    .A2(_22563_),
    .Y(_23056_),
    .B1(_21269_));
 sg13g2_o21ai_1 _31618_ (.B1(net6361),
    .Y(_23057_),
    .A1(_20578_),
    .A2(_23056_));
 sg13g2_a21oi_1 _31619_ (.A1(_20578_),
    .A2(_23056_),
    .Y(_23058_),
    .B1(_23057_));
 sg13g2_a21oi_1 _31620_ (.A1(net6260),
    .A2(_23055_),
    .Y(_23059_),
    .B1(_23058_));
 sg13g2_a21o_1 _31621_ (.A2(_23055_),
    .A1(net6261),
    .B1(_23058_),
    .X(_23060_));
 sg13g2_o21ai_1 _31622_ (.B1(_20630_),
    .Y(_23061_),
    .A1(_20632_),
    .A2(_23027_));
 sg13g2_xnor2_1 _31623_ (.Y(_23062_),
    .A(_20628_),
    .B(_23061_));
 sg13g2_o21ai_1 _31624_ (.B1(net6262),
    .Y(_23063_),
    .A1(\u_inv.f_next[75] ),
    .A2(net7400));
 sg13g2_a21oi_1 _31625_ (.A1(net7400),
    .A2(_23062_),
    .Y(_23064_),
    .B1(_23063_));
 sg13g2_nor3_1 _31626_ (.A(_20629_),
    .B(_21298_),
    .C(_23033_),
    .Y(_23065_));
 sg13g2_o21ai_1 _31627_ (.B1(_20629_),
    .Y(_23066_),
    .A1(_21298_),
    .A2(_23033_));
 sg13g2_nor2_1 _31628_ (.A(net6262),
    .B(_23065_),
    .Y(_23067_));
 sg13g2_a21o_2 _31629_ (.A2(_23067_),
    .A1(_23066_),
    .B1(_23064_),
    .X(_23068_));
 sg13g2_nand2_1 _31630_ (.Y(_23069_),
    .A(_20655_),
    .B(_21313_));
 sg13g2_a21oi_1 _31631_ (.A1(_20658_),
    .A2(_21310_),
    .Y(_23070_),
    .B1(_23069_));
 sg13g2_nand3b_1 _31632_ (.B(net6357),
    .C(_21312_),
    .Y(_23071_),
    .A_N(_21314_));
 sg13g2_or2_1 _31633_ (.X(_23072_),
    .B(_20658_),
    .A(_20654_));
 sg13g2_a21o_1 _31634_ (.A2(_23072_),
    .A1(_20657_),
    .B1(_20655_),
    .X(_23073_));
 sg13g2_nand3_1 _31635_ (.B(_20657_),
    .C(_23072_),
    .A(_20655_),
    .Y(_23074_));
 sg13g2_nand3_1 _31636_ (.B(_23073_),
    .C(_23074_),
    .A(net7398),
    .Y(_23075_));
 sg13g2_o21ai_1 _31637_ (.B1(net6264),
    .Y(_23076_),
    .A1(\u_inv.f_next[81] ),
    .A2(net7397));
 sg13g2_nand2b_1 _31638_ (.Y(_23077_),
    .B(_23075_),
    .A_N(_23076_));
 sg13g2_o21ai_1 _31639_ (.B1(_23077_),
    .Y(_23078_),
    .A1(_23070_),
    .A2(_23071_));
 sg13g2_nand2_1 _31640_ (.Y(_23079_),
    .A(_20577_),
    .B(_23052_));
 sg13g2_o21ai_1 _31641_ (.B1(net7395),
    .Y(_23080_),
    .A1(_20582_),
    .A2(_23079_));
 sg13g2_a21oi_1 _31642_ (.A1(_20582_),
    .A2(_23079_),
    .Y(_23081_),
    .B1(_23080_));
 sg13g2_o21ai_1 _31643_ (.B1(net6260),
    .Y(_23082_),
    .A1(\u_inv.f_next[67] ),
    .A2(net7395));
 sg13g2_o21ai_1 _31644_ (.B1(_21271_),
    .Y(_23083_),
    .A1(_20578_),
    .A2(_23056_));
 sg13g2_o21ai_1 _31645_ (.B1(net6361),
    .Y(_23084_),
    .A1(_20582_),
    .A2(_23083_));
 sg13g2_a21o_1 _31646_ (.A2(_23083_),
    .A1(_20582_),
    .B1(_23084_),
    .X(_23085_));
 sg13g2_o21ai_1 _31647_ (.B1(_23085_),
    .Y(_23086_),
    .A1(_23081_),
    .A2(_23082_));
 sg13g2_nand2_1 _31648_ (.Y(_23087_),
    .A(_20654_),
    .B(_20658_));
 sg13g2_nand3_1 _31649_ (.B(_23072_),
    .C(_23087_),
    .A(net7398),
    .Y(_23088_));
 sg13g2_o21ai_1 _31650_ (.B1(_23088_),
    .Y(_23089_),
    .A1(_18061_),
    .A2(net7401));
 sg13g2_xor2_1 _31651_ (.B(_21310_),
    .A(_20658_),
    .X(_23090_));
 sg13g2_mux2_1 _31652_ (.A0(_23089_),
    .A1(_23090_),
    .S(net6358),
    .X(_23091_));
 sg13g2_nor2_1 _31653_ (.A(_20663_),
    .B(_20669_),
    .Y(_23092_));
 sg13g2_xnor2_1 _31654_ (.Y(_23093_),
    .A(_20663_),
    .B(_20669_));
 sg13g2_o21ai_1 _31655_ (.B1(net6263),
    .Y(_23094_),
    .A1(\u_inv.f_next[82] ),
    .A2(net7398));
 sg13g2_a21o_1 _31656_ (.A2(_23093_),
    .A1(net7398),
    .B1(_23094_),
    .X(_23095_));
 sg13g2_xnor2_1 _31657_ (.Y(_23096_),
    .A(_20669_),
    .B(_21316_));
 sg13g2_o21ai_1 _31658_ (.B1(_23095_),
    .Y(_23097_),
    .A1(net6263),
    .A2(_23096_));
 sg13g2_nand2_1 _31659_ (.Y(_23098_),
    .A(_20666_),
    .B(_21319_));
 sg13g2_a21oi_1 _31660_ (.A1(_20669_),
    .A2(_21316_),
    .Y(_23099_),
    .B1(_23098_));
 sg13g2_o21ai_1 _31661_ (.B1(net6357),
    .Y(_23100_),
    .A1(_20666_),
    .A2(_21319_));
 sg13g2_or2_1 _31662_ (.X(_23101_),
    .B(_23100_),
    .A(_21318_));
 sg13g2_a21oi_1 _31663_ (.A1(\u_inv.f_next[82] ),
    .A2(\u_inv.f_reg[82] ),
    .Y(_23102_),
    .B1(_23092_));
 sg13g2_a21oi_1 _31664_ (.A1(_20666_),
    .A2(_23102_),
    .Y(_23103_),
    .B1(net7236));
 sg13g2_o21ai_1 _31665_ (.B1(_23103_),
    .Y(_23104_),
    .A1(_20666_),
    .A2(_23102_));
 sg13g2_o21ai_1 _31666_ (.B1(net6265),
    .Y(_23105_),
    .A1(\u_inv.f_next[83] ),
    .A2(net7402));
 sg13g2_nand2b_1 _31667_ (.Y(_23106_),
    .B(_23104_),
    .A_N(_23105_));
 sg13g2_o21ai_1 _31668_ (.B1(_23106_),
    .Y(_23107_),
    .A1(_23099_),
    .A2(_23101_));
 sg13g2_nand2b_1 _31669_ (.Y(_23108_),
    .B(_23066_),
    .A_N(_21299_));
 sg13g2_xnor2_1 _31670_ (.Y(_23109_),
    .A(_20623_),
    .B(_23108_));
 sg13g2_o21ai_1 _31671_ (.B1(_20645_),
    .Y(_23110_),
    .A1(_20633_),
    .A2(_23027_));
 sg13g2_a21oi_1 _31672_ (.A1(_20622_),
    .A2(_23110_),
    .Y(_23111_),
    .B1(net7236));
 sg13g2_o21ai_1 _31673_ (.B1(_23111_),
    .Y(_23112_),
    .A1(_20622_),
    .A2(_23110_));
 sg13g2_a21oi_1 _31674_ (.A1(\u_inv.f_next[76] ),
    .A2(net7236),
    .Y(_23113_),
    .B1(net6357));
 sg13g2_a22oi_1 _31675_ (.Y(_23114_),
    .B1(_23112_),
    .B2(_23113_),
    .A2(_23109_),
    .A1(net6357));
 sg13g2_xnor2_1 _31676_ (.Y(_23115_),
    .A(_20673_),
    .B(_20685_));
 sg13g2_a21oi_1 _31677_ (.A1(net7398),
    .A2(_23115_),
    .Y(_23116_),
    .B1(net6357));
 sg13g2_o21ai_1 _31678_ (.B1(_23116_),
    .Y(_23117_),
    .A1(\u_inv.f_next[84] ),
    .A2(net7398));
 sg13g2_xnor2_1 _31679_ (.Y(_23118_),
    .A(_20685_),
    .B(_21322_));
 sg13g2_o21ai_1 _31680_ (.B1(_23117_),
    .Y(_23119_),
    .A1(net6263),
    .A2(_23118_));
 sg13g2_nand4_1 _31681_ (.B(_23017_),
    .C(_23040_),
    .A(_22551_),
    .Y(_23120_),
    .D(_23059_));
 sg13g2_or4_1 _31682_ (.A(_23050_),
    .B(_23086_),
    .C(_23091_),
    .D(_23120_),
    .X(_23121_));
 sg13g2_nor4_1 _31683_ (.A(_23068_),
    .B(_23078_),
    .C(_23097_),
    .D(_23121_),
    .Y(_23122_));
 sg13g2_nor3_1 _31684_ (.A(_22724_),
    .B(_22730_),
    .C(_22997_),
    .Y(_23123_));
 sg13g2_nand3_1 _31685_ (.B(_22989_),
    .C(_23123_),
    .A(_22979_),
    .Y(_23124_));
 sg13g2_nand3b_1 _31686_ (.B(_22701_),
    .C(_22735_),
    .Y(_23125_),
    .A_N(_22666_));
 sg13g2_nor4_1 _31687_ (.A(_22647_),
    .B(_22654_),
    .C(_23124_),
    .D(_23125_),
    .Y(_23126_));
 sg13g2_nand4_1 _31688_ (.B(_22641_),
    .C(_22687_),
    .A(_22620_),
    .Y(_23127_),
    .D(_23126_));
 sg13g2_nand4_1 _31689_ (.B(_22635_),
    .C(_22694_),
    .A(_22602_),
    .Y(_23128_),
    .D(_22709_));
 sg13g2_nor4_1 _31690_ (.A(_22590_),
    .B(_22614_),
    .C(_22674_),
    .D(_23011_),
    .Y(_23129_));
 sg13g2_nand2b_1 _31691_ (.Y(_23130_),
    .B(_23129_),
    .A_N(_22565_));
 sg13g2_nor4_1 _31692_ (.A(_23005_),
    .B(_23127_),
    .C(_23128_),
    .D(_23130_),
    .Y(_23131_));
 sg13g2_nor2_1 _31693_ (.A(_22596_),
    .B(_23025_),
    .Y(_23132_));
 sg13g2_nand4_1 _31694_ (.B(_22582_),
    .C(_23131_),
    .A(_22570_),
    .Y(_23133_),
    .D(_23132_));
 sg13g2_nor3_1 _31695_ (.A(_22526_),
    .B(_22558_),
    .C(_23133_),
    .Y(_23134_));
 sg13g2_and4_1 _31696_ (.A(_22520_),
    .B(_22542_),
    .C(_23035_),
    .D(_23134_),
    .X(_23135_));
 sg13g2_nand3b_1 _31697_ (.B(_23122_),
    .C(_23135_),
    .Y(_23136_),
    .A_N(_23114_));
 sg13g2_nor2_1 _31698_ (.A(_20694_),
    .B(_20715_),
    .Y(_23137_));
 sg13g2_nor2_1 _31699_ (.A(net7236),
    .B(_23137_),
    .Y(_23138_));
 sg13g2_xnor2_1 _31700_ (.Y(_23139_),
    .A(_20715_),
    .B(_21333_));
 sg13g2_a221oi_1 _31701_ (.B2(_23138_),
    .C1(net6359),
    .B1(_22497_),
    .A1(\u_inv.f_next[88] ),
    .Y(_23140_),
    .A2(net7244));
 sg13g2_a21oi_2 _31702_ (.B1(_23140_),
    .Y(_23141_),
    .A2(_23139_),
    .A1(net6359));
 sg13g2_o21ai_1 _31703_ (.B1(_20683_),
    .Y(_23142_),
    .A1(_20673_),
    .A2(_20685_));
 sg13g2_o21ai_1 _31704_ (.B1(net7404),
    .Y(_23143_),
    .A1(_20682_),
    .A2(_23142_));
 sg13g2_a21oi_1 _31705_ (.A1(_20682_),
    .A2(_23142_),
    .Y(_23144_),
    .B1(_23143_));
 sg13g2_nor2b_1 _31706_ (.A(net7404),
    .B_N(\u_inv.f_next[85] ),
    .Y(_23145_));
 sg13g2_o21ai_1 _31707_ (.B1(net6266),
    .Y(_23146_),
    .A1(_23144_),
    .A2(_23145_));
 sg13g2_xnor2_1 _31708_ (.Y(_23147_),
    .A(_20682_),
    .B(_22450_));
 sg13g2_o21ai_1 _31709_ (.B1(_23146_),
    .Y(_23148_),
    .A1(net6266),
    .A2(_23147_));
 sg13g2_a21oi_1 _31710_ (.A1(_20622_),
    .A2(_23110_),
    .Y(_23149_),
    .B1(_20621_));
 sg13g2_xor2_1 _31711_ (.B(_23149_),
    .A(_20624_),
    .X(_23150_));
 sg13g2_o21ai_1 _31712_ (.B1(net6262),
    .Y(_23151_),
    .A1(\u_inv.f_next[77] ),
    .A2(net7399));
 sg13g2_a21oi_1 _31713_ (.A1(net7399),
    .A2(_23150_),
    .Y(_23152_),
    .B1(_23151_));
 sg13g2_a21oi_1 _31714_ (.A1(_20623_),
    .A2(_23108_),
    .Y(_23153_),
    .B1(_21303_));
 sg13g2_or2_1 _31715_ (.X(_23154_),
    .B(_23153_),
    .A(_20624_));
 sg13g2_a21oi_1 _31716_ (.A1(_20624_),
    .A2(_23153_),
    .Y(_23155_),
    .B1(net6262));
 sg13g2_a21o_2 _31717_ (.A2(_23155_),
    .A1(_23154_),
    .B1(_23152_),
    .X(_23156_));
 sg13g2_or4_1 _31718_ (.A(_23107_),
    .B(_23119_),
    .C(_23136_),
    .D(_23156_),
    .X(_23157_));
 sg13g2_nor4_1 _31719_ (.A(_22503_),
    .B(_23141_),
    .C(_23148_),
    .D(_23157_),
    .Y(_23158_));
 sg13g2_a21oi_1 _31720_ (.A1(_20625_),
    .A2(_23110_),
    .Y(_23159_),
    .B1(_20649_));
 sg13g2_o21ai_1 _31721_ (.B1(_20618_),
    .Y(_23160_),
    .A1(_20619_),
    .A2(_23159_));
 sg13g2_xnor2_1 _31722_ (.Y(_23161_),
    .A(_20616_),
    .B(_23160_));
 sg13g2_o21ai_1 _31723_ (.B1(net6263),
    .Y(_23162_),
    .A1(\u_inv.f_next[79] ),
    .A2(net7398));
 sg13g2_a21oi_1 _31724_ (.A1(net7398),
    .A2(_23161_),
    .Y(_23163_),
    .B1(_23162_));
 sg13g2_and2_1 _31725_ (.A(_21302_),
    .B(_23154_),
    .X(_23164_));
 sg13g2_nor2_1 _31726_ (.A(_20620_),
    .B(_23164_),
    .Y(_23165_));
 sg13g2_nor2_1 _31727_ (.A(_21307_),
    .B(_23165_),
    .Y(_23166_));
 sg13g2_o21ai_1 _31728_ (.B1(net6358),
    .Y(_23167_),
    .A1(_20616_),
    .A2(_23166_));
 sg13g2_a21oi_1 _31729_ (.A1(_20616_),
    .A2(_23166_),
    .Y(_23168_),
    .B1(_23167_));
 sg13g2_nor2_2 _31730_ (.A(_23163_),
    .B(_23168_),
    .Y(_23169_));
 sg13g2_xor2_1 _31731_ (.B(_23159_),
    .A(_20620_),
    .X(_23170_));
 sg13g2_a21oi_1 _31732_ (.A1(net7399),
    .A2(_23170_),
    .Y(_23171_),
    .B1(net6357));
 sg13g2_o21ai_1 _31733_ (.B1(_23171_),
    .Y(_23172_),
    .A1(\u_inv.f_next[78] ),
    .A2(net7399));
 sg13g2_and2_1 _31734_ (.A(_20620_),
    .B(_23164_),
    .X(_23173_));
 sg13g2_o21ai_1 _31735_ (.B1(net6361),
    .Y(_23174_),
    .A1(_20620_),
    .A2(_23164_));
 sg13g2_o21ai_1 _31736_ (.B1(_23172_),
    .Y(_23175_),
    .A1(_23173_),
    .A2(_23174_));
 sg13g2_xnor2_1 _31737_ (.Y(_23176_),
    .A(_20708_),
    .B(_22410_));
 sg13g2_nor2_1 _31738_ (.A(\u_inv.f_next[90] ),
    .B(net7403),
    .Y(_23177_));
 sg13g2_a21oi_1 _31739_ (.A1(net7403),
    .A2(_23176_),
    .Y(_23178_),
    .B1(_23177_));
 sg13g2_or3_1 _31740_ (.A(_20708_),
    .B(_21344_),
    .C(_22418_),
    .X(_23179_));
 sg13g2_and2_1 _31741_ (.A(net6360),
    .B(_22467_),
    .X(_23180_));
 sg13g2_a22oi_1 _31742_ (.Y(_23181_),
    .B1(_23179_),
    .B2(_23180_),
    .A2(_23178_),
    .A1(net6266));
 sg13g2_inv_1 _31743_ (.Y(_23182_),
    .A(_23181_));
 sg13g2_xnor2_1 _31744_ (.Y(_23183_),
    .A(_20675_),
    .B(_22456_));
 sg13g2_a21oi_1 _31745_ (.A1(net7404),
    .A2(_23183_),
    .Y(_23184_),
    .B1(net6360));
 sg13g2_o21ai_1 _31746_ (.B1(_23184_),
    .Y(_23185_),
    .A1(\u_inv.f_next[86] ),
    .A2(net7404));
 sg13g2_nor3_1 _31747_ (.A(_20676_),
    .B(_21327_),
    .C(_22451_),
    .Y(_23186_));
 sg13g2_nand2_1 _31748_ (.Y(_23187_),
    .A(net6360),
    .B(_22452_));
 sg13g2_o21ai_1 _31749_ (.B1(_23185_),
    .Y(_23188_),
    .A1(_23186_),
    .A2(_23187_));
 sg13g2_xnor2_1 _31750_ (.Y(_23189_),
    .A(_20759_),
    .B(_21353_));
 sg13g2_o21ai_1 _31751_ (.B1(net7388),
    .Y(_23190_),
    .A1(_20730_),
    .A2(_20759_));
 sg13g2_a21o_1 _31752_ (.A2(_20759_),
    .A1(_20730_),
    .B1(_23190_),
    .X(_23191_));
 sg13g2_a21oi_1 _31753_ (.A1(\u_inv.f_next[96] ),
    .A2(net7229),
    .Y(_23192_),
    .B1(net6348));
 sg13g2_a22oi_1 _31754_ (.Y(_23193_),
    .B1(_23191_),
    .B2(_23192_),
    .A2(_23189_),
    .A1(net6348));
 sg13g2_xnor2_1 _31755_ (.Y(_23194_),
    .A(_20736_),
    .B(_22315_));
 sg13g2_nor2_1 _31756_ (.A(\u_inv.f_next[100] ),
    .B(net7387),
    .Y(_23195_));
 sg13g2_a21oi_1 _31757_ (.A1(net7387),
    .A2(_23194_),
    .Y(_23196_),
    .B1(_23195_));
 sg13g2_nand3_1 _31758_ (.B(_21366_),
    .C(_22306_),
    .A(_20735_),
    .Y(_23197_));
 sg13g2_nor2_1 _31759_ (.A(net6255),
    .B(_22307_),
    .Y(_23198_));
 sg13g2_a22oi_1 _31760_ (.Y(_23199_),
    .B1(_23197_),
    .B2(_23198_),
    .A2(_23196_),
    .A1(net6255));
 sg13g2_nand2b_1 _31761_ (.Y(_23200_),
    .B(_22412_),
    .A_N(_20699_));
 sg13g2_nand3b_1 _31762_ (.B(_23200_),
    .C(net7402),
    .Y(_23201_),
    .A_N(_22413_));
 sg13g2_nand3_1 _31763_ (.B(_21340_),
    .C(_22422_),
    .A(_20699_),
    .Y(_23202_));
 sg13g2_nand2b_1 _31764_ (.Y(_23203_),
    .B(_23202_),
    .A_N(_22423_));
 sg13g2_a21oi_1 _31765_ (.A1(\u_inv.f_next[94] ),
    .A2(net7244),
    .Y(_23204_),
    .B1(net6359));
 sg13g2_a22oi_1 _31766_ (.Y(_23205_),
    .B1(_23204_),
    .B2(_23201_),
    .A2(_23203_),
    .A1(net6359));
 sg13g2_o21ai_1 _31767_ (.B1(_20245_),
    .Y(_23206_),
    .A1(_20290_),
    .A2(_22239_));
 sg13g2_a21oi_1 _31768_ (.A1(_20246_),
    .A2(_22240_),
    .Y(_23207_),
    .B1(net7219));
 sg13g2_a21oi_1 _31769_ (.A1(\u_inv.f_next[121] ),
    .A2(_18221_),
    .Y(_23208_),
    .B1(_22269_));
 sg13g2_nor2_1 _31770_ (.A(_20245_),
    .B(_23208_),
    .Y(_23209_));
 sg13g2_xnor2_1 _31771_ (.Y(_23210_),
    .A(_20245_),
    .B(_23208_));
 sg13g2_a221oi_1 _31772_ (.B2(_23207_),
    .C1(net6334),
    .B1(_23206_),
    .A1(\u_inv.f_next[122] ),
    .Y(_23211_),
    .A2(net7220));
 sg13g2_a21oi_2 _31773_ (.B1(_23211_),
    .Y(_23212_),
    .A2(_23210_),
    .A1(net6334));
 sg13g2_a21oi_1 _31774_ (.A1(\u_inv.f_next[124] ),
    .A2(\u_inv.f_reg[124] ),
    .Y(_23213_),
    .B1(_22243_));
 sg13g2_xnor2_1 _31775_ (.Y(_23214_),
    .A(_20237_),
    .B(_23213_));
 sg13g2_o21ai_1 _31776_ (.B1(net6245),
    .Y(_23215_),
    .A1(\u_inv.f_next[125] ),
    .A2(net7371));
 sg13g2_a21oi_1 _31777_ (.A1(net7371),
    .A2(_23214_),
    .Y(_23216_),
    .B1(_23215_));
 sg13g2_nor3_1 _31778_ (.A(_20237_),
    .B(_21427_),
    .C(_22251_),
    .Y(_23217_));
 sg13g2_o21ai_1 _31779_ (.B1(_20237_),
    .Y(_23218_),
    .A1(_21427_),
    .A2(_22251_));
 sg13g2_nor2_1 _31780_ (.A(net6245),
    .B(_23217_),
    .Y(_23219_));
 sg13g2_a21o_2 _31781_ (.A2(_23219_),
    .A1(_23218_),
    .B1(_23216_),
    .X(_23220_));
 sg13g2_nand3_1 _31782_ (.B(_21472_),
    .C(_21486_),
    .A(_20897_),
    .Y(_23221_));
 sg13g2_nand2b_1 _31783_ (.Y(_23222_),
    .B(_23221_),
    .A_N(_22167_));
 sg13g2_a21oi_1 _31784_ (.A1(_20895_),
    .A2(_20897_),
    .Y(_23223_),
    .B1(net7212));
 sg13g2_o21ai_1 _31785_ (.B1(_23223_),
    .Y(_23224_),
    .A1(_20895_),
    .A2(_20897_));
 sg13g2_a21oi_1 _31786_ (.A1(\u_inv.f_next[144] ),
    .A2(net7212),
    .Y(_23225_),
    .B1(net6320));
 sg13g2_a22oi_1 _31787_ (.Y(_23226_),
    .B1(_23224_),
    .B2(_23225_),
    .A2(_23222_),
    .A1(net6321));
 sg13g2_a21oi_1 _31788_ (.A1(_20825_),
    .A2(_22380_),
    .Y(_23227_),
    .B1(_20824_));
 sg13g2_o21ai_1 _31789_ (.B1(net7365),
    .Y(_23228_),
    .A1(_20827_),
    .A2(_23227_));
 sg13g2_a21oi_1 _31790_ (.A1(_20827_),
    .A2(_23227_),
    .Y(_23229_),
    .B1(_23228_));
 sg13g2_o21ai_1 _31791_ (.B1(net6241),
    .Y(_23230_),
    .A1(\u_inv.f_next[133] ),
    .A2(net7365));
 sg13g2_o21ai_1 _31792_ (.B1(_20828_),
    .Y(_23231_),
    .A1(_21460_),
    .A2(_22386_));
 sg13g2_or3_1 _31793_ (.A(_20828_),
    .B(_21460_),
    .C(_22386_),
    .X(_23232_));
 sg13g2_nand3_1 _31794_ (.B(_23231_),
    .C(_23232_),
    .A(net6331),
    .Y(_23233_));
 sg13g2_o21ai_1 _31795_ (.B1(_23233_),
    .Y(_23234_),
    .A1(_23229_),
    .A2(_23230_));
 sg13g2_a21o_1 _31796_ (.A2(_22178_),
    .A1(_20861_),
    .B1(_20859_),
    .X(_23235_));
 sg13g2_nand3_1 _31797_ (.B(_20861_),
    .C(_22178_),
    .A(_20859_),
    .Y(_23236_));
 sg13g2_nand3_1 _31798_ (.B(_23235_),
    .C(_23236_),
    .A(net7360),
    .Y(_23237_));
 sg13g2_a21oi_1 _31799_ (.A1(_18031_),
    .A2(net7211),
    .Y(_23238_),
    .B1(net6323));
 sg13g2_o21ai_1 _31800_ (.B1(_20860_),
    .Y(_23239_),
    .A1(_21473_),
    .A2(_22219_));
 sg13g2_nor3_1 _31801_ (.A(_20860_),
    .B(_21473_),
    .C(_22219_),
    .Y(_23240_));
 sg13g2_nor2_1 _31802_ (.A(net6237),
    .B(_23240_),
    .Y(_23241_));
 sg13g2_a22oi_1 _31803_ (.Y(_23242_),
    .B1(_23239_),
    .B2(_23241_),
    .A2(_23238_),
    .A1(_23237_));
 sg13g2_inv_2 _31804_ (.Y(_23243_),
    .A(_23242_));
 sg13g2_xnor2_1 _31805_ (.Y(_23244_),
    .A(_20838_),
    .B(_22379_));
 sg13g2_nor2_1 _31806_ (.A(\u_inv.f_next[130] ),
    .B(net7368),
    .Y(_23245_));
 sg13g2_a21oi_1 _31807_ (.A1(net7368),
    .A2(_23244_),
    .Y(_23246_),
    .B1(_23245_));
 sg13g2_nor3_1 _31808_ (.A(_20838_),
    .B(_21453_),
    .C(_22279_),
    .Y(_23247_));
 sg13g2_o21ai_1 _31809_ (.B1(_20838_),
    .Y(_23248_),
    .A1(_21453_),
    .A2(_22279_));
 sg13g2_nor2_1 _31810_ (.A(net6243),
    .B(_23247_),
    .Y(_23249_));
 sg13g2_a22oi_1 _31811_ (.Y(_23250_),
    .B1(_23248_),
    .B2(_23249_),
    .A2(_23246_),
    .A1(net6243));
 sg13g2_inv_2 _31812_ (.Y(_23251_),
    .A(_23250_));
 sg13g2_o21ai_1 _31813_ (.B1(_20281_),
    .Y(_23252_),
    .A1(_20263_),
    .A2(_22225_));
 sg13g2_xnor2_1 _31814_ (.Y(_23253_),
    .A(_20256_),
    .B(_23252_));
 sg13g2_a21oi_1 _31815_ (.A1(net7380),
    .A2(_23253_),
    .Y(_23254_),
    .B1(net6333));
 sg13g2_o21ai_1 _31816_ (.B1(_23254_),
    .Y(_23255_),
    .A1(\u_inv.f_next[118] ),
    .A2(net7380));
 sg13g2_o21ai_1 _31817_ (.B1(_20255_),
    .Y(_23256_),
    .A1(_21410_),
    .A2(_22232_));
 sg13g2_nor3_1 _31818_ (.A(_20255_),
    .B(_21410_),
    .C(_22232_),
    .Y(_23257_));
 sg13g2_nand2_1 _31819_ (.Y(_23258_),
    .A(net6333),
    .B(_23256_));
 sg13g2_o21ai_1 _31820_ (.B1(_23255_),
    .Y(_23259_),
    .A1(_23257_),
    .A2(_23258_));
 sg13g2_a21oi_1 _31821_ (.A1(_20266_),
    .A2(_22224_),
    .Y(_23260_),
    .B1(_20265_));
 sg13g2_a21oi_1 _31822_ (.A1(_20268_),
    .A2(_23260_),
    .Y(_23261_),
    .B1(net7228));
 sg13g2_o21ai_1 _31823_ (.B1(_23261_),
    .Y(_23262_),
    .A1(_20268_),
    .A2(_23260_));
 sg13g2_o21ai_1 _31824_ (.B1(_23262_),
    .Y(_23263_),
    .A1(\u_inv.f_next[115] ),
    .A2(net7383));
 sg13g2_o21ai_1 _31825_ (.B1(_20269_),
    .Y(_23264_),
    .A1(_21414_),
    .A2(_22260_));
 sg13g2_or3_1 _31826_ (.A(_20269_),
    .B(_21414_),
    .C(_22260_),
    .X(_23265_));
 sg13g2_nand3_1 _31827_ (.B(_23264_),
    .C(_23265_),
    .A(net6344),
    .Y(_23266_));
 sg13g2_o21ai_1 _31828_ (.B1(_23266_),
    .Y(_23267_),
    .A1(net6344),
    .A2(_23263_));
 sg13g2_xor2_1 _31829_ (.B(_22182_),
    .A(_20870_),
    .X(_23268_));
 sg13g2_o21ai_1 _31830_ (.B1(net6233),
    .Y(_23269_),
    .A1(\u_inv.f_next[142] ),
    .A2(net7356));
 sg13g2_a21oi_1 _31831_ (.A1(net7356),
    .A2(_23268_),
    .Y(_23270_),
    .B1(_23269_));
 sg13g2_and3_1 _31832_ (.X(_23271_),
    .A(_20870_),
    .B(_21482_),
    .C(_22189_));
 sg13g2_nor3_1 _31833_ (.A(net6233),
    .B(_22190_),
    .C(_23271_),
    .Y(_23272_));
 sg13g2_nor2_2 _31834_ (.A(_23270_),
    .B(_23272_),
    .Y(_23273_));
 sg13g2_xnor2_1 _31835_ (.Y(_23274_),
    .A(_20185_),
    .B(_22162_));
 sg13g2_o21ai_1 _31836_ (.B1(net6235),
    .Y(_23275_),
    .A1(\u_inv.f_next[148] ),
    .A2(net7357));
 sg13g2_a21o_1 _31837_ (.A2(_23274_),
    .A1(net7358),
    .B1(_23275_),
    .X(_23276_));
 sg13g2_nor3_1 _31838_ (.A(_20186_),
    .B(_21520_),
    .C(_22168_),
    .Y(_23277_));
 sg13g2_nand2_1 _31839_ (.Y(_23278_),
    .A(net6320),
    .B(_22169_));
 sg13g2_o21ai_1 _31840_ (.B1(_23276_),
    .Y(_23279_),
    .A1(_23277_),
    .A2(_23278_));
 sg13g2_nand2_1 _31841_ (.Y(_23280_),
    .A(_20127_),
    .B(_22047_));
 sg13g2_xnor2_1 _31842_ (.Y(_23281_),
    .A(_20127_),
    .B(_22047_));
 sg13g2_o21ai_1 _31843_ (.B1(net6217),
    .Y(_23282_),
    .A1(\u_inv.f_next[164] ),
    .A2(net7328));
 sg13g2_a21oi_1 _31844_ (.A1(net7328),
    .A2(_23281_),
    .Y(_23283_),
    .B1(_23282_));
 sg13g2_nand3_1 _31845_ (.B(_21551_),
    .C(_22037_),
    .A(_20127_),
    .Y(_23284_));
 sg13g2_and2_1 _31846_ (.A(_22107_),
    .B(_23284_),
    .X(_23285_));
 sg13g2_a21oi_2 _31847_ (.B1(_23283_),
    .Y(_23286_),
    .A2(_23285_),
    .A1(net6298));
 sg13g2_nand3_1 _31848_ (.B(_21543_),
    .C(_21575_),
    .A(_20915_),
    .Y(_23287_));
 sg13g2_nand2b_1 _31849_ (.Y(_23288_),
    .B(_23287_),
    .A_N(_22075_));
 sg13g2_nand3_1 _31850_ (.B(_20912_),
    .C(_20916_),
    .A(_20154_),
    .Y(_23289_));
 sg13g2_nand3b_1 _31851_ (.B(_23289_),
    .C(net7324),
    .Y(_23290_),
    .A_N(_22069_));
 sg13g2_a21oi_1 _31852_ (.A1(\u_inv.f_next[176] ),
    .A2(net7196),
    .Y(_23291_),
    .B1(net6297));
 sg13g2_a22oi_1 _31853_ (.Y(_23292_),
    .B1(_23290_),
    .B2(_23291_),
    .A2(_23288_),
    .A1(net6297));
 sg13g2_a21o_1 _31854_ (.A2(_23231_),
    .A1(_21459_),
    .B1(_20831_),
    .X(_23293_));
 sg13g2_nand2b_1 _31855_ (.Y(_23294_),
    .B(_23293_),
    .A_N(_21458_));
 sg13g2_a21oi_1 _31856_ (.A1(_20834_),
    .A2(_23294_),
    .Y(_23295_),
    .B1(net6241));
 sg13g2_o21ai_1 _31857_ (.B1(_23295_),
    .Y(_23296_),
    .A1(_20834_),
    .A2(_23294_));
 sg13g2_a21oi_1 _31858_ (.A1(_20829_),
    .A2(_22380_),
    .Y(_23297_),
    .B1(_20852_));
 sg13g2_nand2b_1 _31859_ (.Y(_23298_),
    .B(_20831_),
    .A_N(_23297_));
 sg13g2_a21oi_1 _31860_ (.A1(_20830_),
    .A2(_23298_),
    .Y(_23299_),
    .B1(_20833_));
 sg13g2_and3_1 _31861_ (.X(_23300_),
    .A(_20830_),
    .B(_20833_),
    .C(_23298_));
 sg13g2_nor3_1 _31862_ (.A(net7219),
    .B(_23299_),
    .C(_23300_),
    .Y(_23301_));
 sg13g2_o21ai_1 _31863_ (.B1(net6241),
    .Y(_23302_),
    .A1(\u_inv.f_next[135] ),
    .A2(net7365));
 sg13g2_o21ai_1 _31864_ (.B1(_23296_),
    .Y(_23303_),
    .A1(_23301_),
    .A2(_23302_));
 sg13g2_a21oi_1 _31865_ (.A1(_21475_),
    .A2(_23239_),
    .Y(_23304_),
    .B1(_20877_));
 sg13g2_o21ai_1 _31866_ (.B1(_20879_),
    .Y(_23305_),
    .A1(_21474_),
    .A2(_23304_));
 sg13g2_nor3_1 _31867_ (.A(_20879_),
    .B(_21474_),
    .C(_23304_),
    .Y(_23306_));
 sg13g2_nor2_1 _31868_ (.A(net6237),
    .B(_23306_),
    .Y(_23307_));
 sg13g2_a21oi_1 _31869_ (.A1(_20877_),
    .A2(_22179_),
    .Y(_23308_),
    .B1(_20876_));
 sg13g2_xnor2_1 _31870_ (.Y(_23309_),
    .A(_20879_),
    .B(_23308_));
 sg13g2_o21ai_1 _31871_ (.B1(net6237),
    .Y(_23310_),
    .A1(\u_inv.f_next[139] ),
    .A2(net7360));
 sg13g2_a21oi_1 _31872_ (.A1(net7360),
    .A2(_23309_),
    .Y(_23311_),
    .B1(_23310_));
 sg13g2_a21o_2 _31873_ (.A2(_23307_),
    .A1(_23305_),
    .B1(_23311_),
    .X(_23312_));
 sg13g2_nor2_1 _31874_ (.A(_21436_),
    .B(_23209_),
    .Y(_23313_));
 sg13g2_a21oi_1 _31875_ (.A1(_20247_),
    .A2(_23313_),
    .Y(_23314_),
    .B1(net6245));
 sg13g2_o21ai_1 _31876_ (.B1(_23314_),
    .Y(_23315_),
    .A1(_20247_),
    .A2(_23313_));
 sg13g2_and3_1 _31877_ (.X(_23316_),
    .A(_20244_),
    .B(_20247_),
    .C(_23206_));
 sg13g2_a21oi_1 _31878_ (.A1(_20244_),
    .A2(_23206_),
    .Y(_23317_),
    .B1(_20247_));
 sg13g2_nor3_1 _31879_ (.A(net7220),
    .B(_23316_),
    .C(_23317_),
    .Y(_23318_));
 sg13g2_o21ai_1 _31880_ (.B1(net6245),
    .Y(_23319_),
    .A1(\u_inv.f_next[123] ),
    .A2(net7371));
 sg13g2_o21ai_1 _31881_ (.B1(_23315_),
    .Y(_23320_),
    .A1(_23318_),
    .A2(_23319_));
 sg13g2_nand3_1 _31882_ (.B(_21423_),
    .C(_23256_),
    .A(_20253_),
    .Y(_23321_));
 sg13g2_a21o_1 _31883_ (.A2(_23256_),
    .A1(_21423_),
    .B1(_20253_),
    .X(_23322_));
 sg13g2_nand3_1 _31884_ (.B(_23321_),
    .C(_23322_),
    .A(net6333),
    .Y(_23323_));
 sg13g2_a21oi_1 _31885_ (.A1(_20256_),
    .A2(_23252_),
    .Y(_23324_),
    .B1(_20254_));
 sg13g2_o21ai_1 _31886_ (.B1(net7371),
    .Y(_23325_),
    .A1(_20253_),
    .A2(_23324_));
 sg13g2_a21oi_1 _31887_ (.A1(_20253_),
    .A2(_23324_),
    .Y(_23326_),
    .B1(_23325_));
 sg13g2_o21ai_1 _31888_ (.B1(net6245),
    .Y(_23327_),
    .A1(\u_inv.f_next[119] ),
    .A2(net7371));
 sg13g2_o21ai_1 _31889_ (.B1(_23323_),
    .Y(_23328_),
    .A1(_23326_),
    .A2(_23327_));
 sg13g2_xnor2_1 _31890_ (.Y(_23329_),
    .A(_20906_),
    .B(_21531_));
 sg13g2_nor3_1 _31891_ (.A(_20227_),
    .B(_20904_),
    .C(_20905_),
    .Y(_23330_));
 sg13g2_o21ai_1 _31892_ (.B1(_20905_),
    .Y(_23331_),
    .A1(_20227_),
    .A2(_20904_));
 sg13g2_nand3b_1 _31893_ (.B(_23331_),
    .C(net7339),
    .Y(_23332_),
    .A_N(_23330_));
 sg13g2_a21oi_1 _31894_ (.A1(\u_inv.f_next[160] ),
    .A2(net7204),
    .Y(_23333_),
    .B1(net6307));
 sg13g2_a22oi_1 _31895_ (.Y(_23334_),
    .B1(_23332_),
    .B2(_23333_),
    .A2(_23329_),
    .A1(net6307));
 sg13g2_a21oi_1 _31896_ (.A1(_20895_),
    .A2(_20897_),
    .Y(_23335_),
    .B1(_20203_));
 sg13g2_xnor2_1 _31897_ (.Y(_23336_),
    .A(_20899_),
    .B(_23335_));
 sg13g2_o21ai_1 _31898_ (.B1(net6236),
    .Y(_23337_),
    .A1(\u_inv.f_next[145] ),
    .A2(net7359));
 sg13g2_a21oi_1 _31899_ (.A1(net7358),
    .A2(_23336_),
    .Y(_23338_),
    .B1(_23337_));
 sg13g2_nor3_1 _31900_ (.A(_20899_),
    .B(_21515_),
    .C(_22167_),
    .Y(_23339_));
 sg13g2_o21ai_1 _31901_ (.B1(_20899_),
    .Y(_23340_),
    .A1(_21515_),
    .A2(_22167_));
 sg13g2_nor2_1 _31902_ (.A(net6236),
    .B(_23339_),
    .Y(_23341_));
 sg13g2_a21o_2 _31903_ (.A2(_23341_),
    .A1(_23340_),
    .B1(_23338_),
    .X(_23342_));
 sg13g2_inv_1 _31904_ (.Y(_23343_),
    .A(_23342_));
 sg13g2_a21oi_1 _31905_ (.A1(_20866_),
    .A2(_22188_),
    .Y(_23344_),
    .B1(_20864_));
 sg13g2_nand2_1 _31906_ (.Y(_23345_),
    .A(_21480_),
    .B(_23344_));
 sg13g2_nor2_1 _31907_ (.A(net6234),
    .B(_21481_),
    .Y(_23346_));
 sg13g2_and2_1 _31908_ (.A(_22189_),
    .B(_23346_),
    .X(_23347_));
 sg13g2_o21ai_1 _31909_ (.B1(_20865_),
    .Y(_23348_),
    .A1(_20866_),
    .A2(_22180_));
 sg13g2_xnor2_1 _31910_ (.Y(_23349_),
    .A(_20863_),
    .B(_23348_));
 sg13g2_o21ai_1 _31911_ (.B1(net6233),
    .Y(_23350_),
    .A1(\u_inv.f_next[141] ),
    .A2(net7356));
 sg13g2_a21oi_1 _31912_ (.A1(net7356),
    .A2(_23349_),
    .Y(_23351_),
    .B1(_23350_));
 sg13g2_a21oi_1 _31913_ (.A1(_23345_),
    .A2(_23347_),
    .Y(_23352_),
    .B1(_23351_));
 sg13g2_inv_1 _31914_ (.Y(_23353_),
    .A(_23352_));
 sg13g2_a21oi_1 _31915_ (.A1(_20906_),
    .A2(_21531_),
    .Y(_23354_),
    .B1(_20908_));
 sg13g2_nand2b_1 _31916_ (.Y(_23355_),
    .B(_23354_),
    .A_N(_21545_));
 sg13g2_o21ai_1 _31917_ (.B1(_21532_),
    .Y(_23356_),
    .A1(_21497_),
    .A2(_21530_));
 sg13g2_a221oi_1 _31918_ (.B2(_20908_),
    .C1(net6223),
    .B1(_21545_),
    .A1(_21531_),
    .Y(_23357_),
    .A2(_21532_));
 sg13g2_nand2_1 _31919_ (.Y(_23358_),
    .A(_20140_),
    .B(_23331_));
 sg13g2_xnor2_1 _31920_ (.Y(_23359_),
    .A(_20907_),
    .B(_23358_));
 sg13g2_o21ai_1 _31921_ (.B1(net6223),
    .Y(_23360_),
    .A1(\u_inv.f_next[161] ),
    .A2(net7339));
 sg13g2_a21oi_1 _31922_ (.A1(net7340),
    .A2(_23359_),
    .Y(_23361_),
    .B1(_23360_));
 sg13g2_a21oi_2 _31923_ (.B1(_23361_),
    .Y(_23362_),
    .A2(_23357_),
    .A1(_23355_));
 sg13g2_a21oi_1 _31924_ (.A1(_20238_),
    .A2(_22242_),
    .Y(_23363_),
    .B1(_20286_));
 sg13g2_xnor2_1 _31925_ (.Y(_23364_),
    .A(_20233_),
    .B(_23363_));
 sg13g2_a21oi_1 _31926_ (.A1(net7369),
    .A2(_23364_),
    .Y(_23365_),
    .B1(net6332));
 sg13g2_o21ai_1 _31927_ (.B1(_23365_),
    .Y(_23366_),
    .A1(\u_inv.f_next[126] ),
    .A2(net7370));
 sg13g2_nor2b_1 _31928_ (.A(_21430_),
    .B_N(_23218_),
    .Y(_23367_));
 sg13g2_nor2_1 _31929_ (.A(_20232_),
    .B(_23367_),
    .Y(_23368_));
 sg13g2_a21o_1 _31930_ (.A2(_23367_),
    .A1(_20232_),
    .B1(net6244),
    .X(_23369_));
 sg13g2_o21ai_1 _31931_ (.B1(_23366_),
    .Y(_23370_),
    .A1(_23368_),
    .A2(_23369_));
 sg13g2_a21oi_2 _31932_ (.B1(_20215_),
    .Y(_23371_),
    .A2(_20901_),
    .A1(_20895_));
 sg13g2_nor2_1 _31933_ (.A(_20173_),
    .B(_23371_),
    .Y(_23372_));
 sg13g2_xnor2_1 _31934_ (.Y(_23373_),
    .A(_20173_),
    .B(_23371_));
 sg13g2_o21ai_1 _31935_ (.B1(net6235),
    .Y(_23374_),
    .A1(\u_inv.f_next[152] ),
    .A2(net7357));
 sg13g2_a21oi_1 _31936_ (.A1(net7357),
    .A2(_23373_),
    .Y(_23375_),
    .B1(_23374_));
 sg13g2_o21ai_1 _31937_ (.B1(_21495_),
    .Y(_23376_),
    .A1(_21471_),
    .A2(_21487_));
 sg13g2_a21oi_1 _31938_ (.A1(_21525_),
    .A2(_23376_),
    .Y(_23377_),
    .B1(_20172_));
 sg13g2_and3_1 _31939_ (.X(_23378_),
    .A(_20172_),
    .B(_21525_),
    .C(_23376_));
 sg13g2_nor3_1 _31940_ (.A(net6235),
    .B(_23377_),
    .C(_23378_),
    .Y(_23379_));
 sg13g2_nor2_1 _31941_ (.A(_23375_),
    .B(_23379_),
    .Y(_23380_));
 sg13g2_inv_4 _31942_ (.A(_23380_),
    .Y(_23381_));
 sg13g2_o21ai_1 _31943_ (.B1(_20142_),
    .Y(_23382_),
    .A1(_20908_),
    .A2(_23331_));
 sg13g2_xnor2_1 _31944_ (.Y(_23383_),
    .A(_20135_),
    .B(_23382_));
 sg13g2_o21ai_1 _31945_ (.B1(net6223),
    .Y(_23384_),
    .A1(\u_inv.f_next[162] ),
    .A2(net7339));
 sg13g2_a21oi_1 _31946_ (.A1(net7340),
    .A2(_23383_),
    .Y(_23385_),
    .B1(_23384_));
 sg13g2_nand3_1 _31947_ (.B(_21547_),
    .C(_23356_),
    .A(_20135_),
    .Y(_23386_));
 sg13g2_a21oi_1 _31948_ (.A1(_21547_),
    .A2(_23356_),
    .Y(_23387_),
    .B1(_20135_));
 sg13g2_nor2_1 _31949_ (.A(net6224),
    .B(_23387_),
    .Y(_23388_));
 sg13g2_a21o_2 _31950_ (.A2(_23388_),
    .A1(_23386_),
    .B1(_23385_),
    .X(_23389_));
 sg13g2_a21oi_1 _31951_ (.A1(_21450_),
    .A2(_23248_),
    .Y(_23390_),
    .B1(_20840_));
 sg13g2_nand3_1 _31952_ (.B(_21450_),
    .C(_23248_),
    .A(_20840_),
    .Y(_23391_));
 sg13g2_nor2_1 _31953_ (.A(net6243),
    .B(_23390_),
    .Y(_23392_));
 sg13g2_o21ai_1 _31954_ (.B1(_20837_),
    .Y(_23393_),
    .A1(_20838_),
    .A2(_22379_));
 sg13g2_xnor2_1 _31955_ (.Y(_23394_),
    .A(_20840_),
    .B(_23393_));
 sg13g2_o21ai_1 _31956_ (.B1(net6242),
    .Y(_23395_),
    .A1(\u_inv.f_next[131] ),
    .A2(net7367));
 sg13g2_a21oi_1 _31957_ (.A1(net7367),
    .A2(_23394_),
    .Y(_23396_),
    .B1(_23395_));
 sg13g2_a21oi_2 _31958_ (.B1(_23396_),
    .Y(_23397_),
    .A2(_23392_),
    .A1(_23391_));
 sg13g2_nand2b_1 _31959_ (.Y(_23398_),
    .B(_23297_),
    .A_N(_20831_));
 sg13g2_nand3_1 _31960_ (.B(_23298_),
    .C(_23398_),
    .A(net7366),
    .Y(_23399_));
 sg13g2_nand3_1 _31961_ (.B(_21459_),
    .C(_23231_),
    .A(_20831_),
    .Y(_23400_));
 sg13g2_nand2_1 _31962_ (.Y(_23401_),
    .A(_23293_),
    .B(_23400_));
 sg13g2_a21oi_1 _31963_ (.A1(\u_inv.f_next[134] ),
    .A2(net7219),
    .Y(_23402_),
    .B1(net6331));
 sg13g2_a22oi_1 _31964_ (.Y(_23403_),
    .B1(_23402_),
    .B2(_23399_),
    .A2(_23401_),
    .A1(net6331));
 sg13g2_xnor2_1 _31965_ (.Y(_23404_),
    .A(_20877_),
    .B(_22179_));
 sg13g2_a21oi_1 _31966_ (.A1(net7360),
    .A2(_23404_),
    .Y(_23405_),
    .B1(net6323));
 sg13g2_o21ai_1 _31967_ (.B1(_23405_),
    .Y(_23406_),
    .A1(\u_inv.f_next[138] ),
    .A2(net7360));
 sg13g2_nand3_1 _31968_ (.B(_21475_),
    .C(_23239_),
    .A(_20877_),
    .Y(_23407_));
 sg13g2_nand2_1 _31969_ (.Y(_23408_),
    .A(net6323),
    .B(_23407_));
 sg13g2_o21ai_1 _31970_ (.B1(_23406_),
    .Y(_23409_),
    .A1(_23304_),
    .A2(_23408_));
 sg13g2_nor2_1 _31971_ (.A(_23403_),
    .B(_23409_),
    .Y(_23410_));
 sg13g2_nand3_1 _31972_ (.B(_20129_),
    .C(_23280_),
    .A(_20123_),
    .Y(_23411_));
 sg13g2_a21o_1 _31973_ (.A2(_23280_),
    .A1(_20123_),
    .B1(_20129_),
    .X(_23412_));
 sg13g2_nand3_1 _31974_ (.B(_23411_),
    .C(_23412_),
    .A(net7329),
    .Y(_23413_));
 sg13g2_a21oi_1 _31975_ (.A1(_18016_),
    .A2(net7197),
    .Y(_23414_),
    .B1(net6298));
 sg13g2_nand3_1 _31976_ (.B(_21566_),
    .C(_22107_),
    .A(_20129_),
    .Y(_23415_));
 sg13g2_nor2_1 _31977_ (.A(net6217),
    .B(_22108_),
    .Y(_23416_));
 sg13g2_a22oi_1 _31978_ (.Y(_23417_),
    .B1(_23415_),
    .B2(_23416_),
    .A2(_23414_),
    .A1(_23413_));
 sg13g2_inv_2 _31979_ (.Y(_23418_),
    .A(_23417_));
 sg13g2_o21ai_1 _31980_ (.B1(_20222_),
    .Y(_23419_),
    .A1(_20174_),
    .A2(_23371_));
 sg13g2_nand2_1 _31981_ (.Y(_23420_),
    .A(_20176_),
    .B(_23419_));
 sg13g2_xnor2_1 _31982_ (.Y(_23421_),
    .A(_20176_),
    .B(_23419_));
 sg13g2_nor2_1 _31983_ (.A(\u_inv.f_next[154] ),
    .B(net7354),
    .Y(_23422_));
 sg13g2_a21oi_1 _31984_ (.A1(net7357),
    .A2(_23421_),
    .Y(_23423_),
    .B1(_23422_));
 sg13g2_o21ai_1 _31985_ (.B1(_20170_),
    .Y(_23424_),
    .A1(_21501_),
    .A2(_23377_));
 sg13g2_a21oi_1 _31986_ (.A1(_21503_),
    .A2(_23424_),
    .Y(_23425_),
    .B1(_20176_));
 sg13g2_nand3_1 _31987_ (.B(_21503_),
    .C(_23424_),
    .A(_20176_),
    .Y(_23426_));
 sg13g2_nor2_1 _31988_ (.A(net6235),
    .B(_23425_),
    .Y(_23427_));
 sg13g2_a22oi_1 _31989_ (.Y(_23428_),
    .B1(_23426_),
    .B2(_23427_),
    .A2(_23423_),
    .A1(net6235));
 sg13g2_inv_1 _31990_ (.Y(_23429_),
    .A(_23428_));
 sg13g2_a21oi_1 _31991_ (.A1(\u_inv.f_next[176] ),
    .A2(\u_inv.f_reg[176] ),
    .Y(_23430_),
    .B1(_22069_));
 sg13g2_xnor2_1 _31992_ (.Y(_23431_),
    .A(_20914_),
    .B(_23430_));
 sg13g2_o21ai_1 _31993_ (.B1(net6215),
    .Y(_23432_),
    .A1(\u_inv.f_next[177] ),
    .A2(net7324));
 sg13g2_a21oi_1 _31994_ (.A1(net7324),
    .A2(_23431_),
    .Y(_23433_),
    .B1(_23432_));
 sg13g2_nor3_1 _31995_ (.A(_20914_),
    .B(_21589_),
    .C(_22075_),
    .Y(_23434_));
 sg13g2_nor2_1 _31996_ (.A(net6215),
    .B(_23434_),
    .Y(_23435_));
 sg13g2_a21oi_2 _31997_ (.B1(_23433_),
    .Y(_23436_),
    .A2(_23435_),
    .A1(_22076_));
 sg13g2_inv_1 _31998_ (.Y(_23437_),
    .A(_23436_));
 sg13g2_o21ai_1 _31999_ (.B1(_20225_),
    .Y(_23438_),
    .A1(_20180_),
    .A2(_23371_));
 sg13g2_nor2b_1 _32000_ (.A(_20165_),
    .B_N(_23438_),
    .Y(_23439_));
 sg13g2_or2_1 _32001_ (.X(_23440_),
    .B(_23439_),
    .A(_20164_));
 sg13g2_o21ai_1 _32002_ (.B1(net7354),
    .Y(_23441_),
    .A1(_20163_),
    .A2(_23440_));
 sg13g2_a21oi_1 _32003_ (.A1(_20163_),
    .A2(_23440_),
    .Y(_23442_),
    .B1(_23441_));
 sg13g2_o21ai_1 _32004_ (.B1(net6232),
    .Y(_23443_),
    .A1(\u_inv.f_next[157] ),
    .A2(net7353));
 sg13g2_a21oi_1 _32005_ (.A1(_21525_),
    .A2(_23376_),
    .Y(_23444_),
    .B1(_21488_));
 sg13g2_o21ai_1 _32006_ (.B1(_20165_),
    .Y(_23445_),
    .A1(_21507_),
    .A2(_23444_));
 sg13g2_nand3_1 _32007_ (.B(_21499_),
    .C(_23445_),
    .A(_20162_),
    .Y(_23446_));
 sg13g2_a21oi_1 _32008_ (.A1(_21499_),
    .A2(_23445_),
    .Y(_23447_),
    .B1(_20162_));
 sg13g2_nand3b_1 _32009_ (.B(net6318),
    .C(_23446_),
    .Y(_23448_),
    .A_N(_23447_));
 sg13g2_o21ai_1 _32010_ (.B1(_23448_),
    .Y(_23449_),
    .A1(_23442_),
    .A2(_23443_));
 sg13g2_nor2_1 _32011_ (.A(_21544_),
    .B(_23387_),
    .Y(_23450_));
 sg13g2_a21oi_1 _32012_ (.A1(_20138_),
    .A2(_23450_),
    .Y(_23451_),
    .B1(net6223));
 sg13g2_o21ai_1 _32013_ (.B1(_23451_),
    .Y(_23452_),
    .A1(_20138_),
    .A2(_23450_));
 sg13g2_a21oi_1 _32014_ (.A1(_20135_),
    .A2(_23382_),
    .Y(_23453_),
    .B1(_20134_));
 sg13g2_o21ai_1 _32015_ (.B1(net7340),
    .Y(_23454_),
    .A1(_20138_),
    .A2(_23453_));
 sg13g2_a21oi_1 _32016_ (.A1(_20138_),
    .A2(_23453_),
    .Y(_23455_),
    .B1(_23454_));
 sg13g2_o21ai_1 _32017_ (.B1(net6224),
    .Y(_23456_),
    .A1(\u_inv.f_next[163] ),
    .A2(net7340));
 sg13g2_o21ai_1 _32018_ (.B1(_23452_),
    .Y(_23457_),
    .A1(_23455_),
    .A2(_23456_));
 sg13g2_or3_1 _32019_ (.A(_20170_),
    .B(_20171_),
    .C(_23372_),
    .X(_23458_));
 sg13g2_o21ai_1 _32020_ (.B1(_20170_),
    .Y(_23459_),
    .A1(_20171_),
    .A2(_23372_));
 sg13g2_nand3_1 _32021_ (.B(_23458_),
    .C(_23459_),
    .A(net7357),
    .Y(_23460_));
 sg13g2_a21oi_1 _32022_ (.A1(_18022_),
    .A2(net7212),
    .Y(_23461_),
    .B1(net6320));
 sg13g2_and2_1 _32023_ (.A(_23460_),
    .B(_23461_),
    .X(_23462_));
 sg13g2_nor3_1 _32024_ (.A(_20170_),
    .B(_21501_),
    .C(_23377_),
    .Y(_23463_));
 sg13g2_nor2_1 _32025_ (.A(net6235),
    .B(_23463_),
    .Y(_23464_));
 sg13g2_a22oi_1 _32026_ (.Y(_23465_),
    .B1(_23464_),
    .B2(_23424_),
    .A2(_23461_),
    .A1(_23460_));
 sg13g2_a21o_2 _32027_ (.A2(_23464_),
    .A1(_23424_),
    .B1(_23462_),
    .X(_23466_));
 sg13g2_o21ai_1 _32028_ (.B1(_20231_),
    .Y(_23467_),
    .A1(_20233_),
    .A2(_23363_));
 sg13g2_o21ai_1 _32029_ (.B1(net7369),
    .Y(_23468_),
    .A1(_20230_),
    .A2(_23467_));
 sg13g2_a21oi_1 _32030_ (.A1(_20230_),
    .A2(_23467_),
    .Y(_23469_),
    .B1(_23468_));
 sg13g2_o21ai_1 _32031_ (.B1(net6244),
    .Y(_23470_),
    .A1(\u_inv.f_next[127] ),
    .A2(net7369));
 sg13g2_nor2_1 _32032_ (.A(_23469_),
    .B(_23470_),
    .Y(_23471_));
 sg13g2_nor2_1 _32033_ (.A(_21428_),
    .B(_23368_),
    .Y(_23472_));
 sg13g2_xnor2_1 _32034_ (.Y(_23473_),
    .A(_20230_),
    .B(_23472_));
 sg13g2_a21oi_2 _32035_ (.B1(_23471_),
    .Y(_23474_),
    .A2(_23473_),
    .A1(net6332));
 sg13g2_xor2_1 _32036_ (.B(_23438_),
    .A(_20165_),
    .X(_23475_));
 sg13g2_nor2_1 _32037_ (.A(\u_inv.f_next[156] ),
    .B(net7354),
    .Y(_23476_));
 sg13g2_a21oi_1 _32038_ (.A1(net7354),
    .A2(_23475_),
    .Y(_23477_),
    .B1(_23476_));
 sg13g2_or3_1 _32039_ (.A(_20165_),
    .B(_21507_),
    .C(_23444_),
    .X(_23478_));
 sg13g2_and2_1 _32040_ (.A(net6318),
    .B(_23445_),
    .X(_23479_));
 sg13g2_a22oi_1 _32041_ (.Y(_23480_),
    .B1(_23478_),
    .B2(_23479_),
    .A2(_23477_),
    .A1(net6232));
 sg13g2_o21ai_1 _32042_ (.B1(_20198_),
    .Y(_23481_),
    .A1(_20205_),
    .A2(_22159_));
 sg13g2_xor2_1 _32043_ (.B(_22160_),
    .A(_20198_),
    .X(_23482_));
 sg13g2_nor2_1 _32044_ (.A(\u_inv.f_next[146] ),
    .B(net7358),
    .Y(_23483_));
 sg13g2_a21oi_1 _32045_ (.A1(net7358),
    .A2(_23482_),
    .Y(_23484_),
    .B1(_23483_));
 sg13g2_nand3_1 _32046_ (.B(_21514_),
    .C(_23340_),
    .A(_20198_),
    .Y(_23485_));
 sg13g2_a21oi_1 _32047_ (.A1(_21514_),
    .A2(_23340_),
    .Y(_23486_),
    .B1(_20198_));
 sg13g2_nor2_1 _32048_ (.A(net6236),
    .B(_23486_),
    .Y(_23487_));
 sg13g2_a22oi_1 _32049_ (.Y(_23488_),
    .B1(_23485_),
    .B2(_23487_),
    .A2(_23484_),
    .A1(net6236));
 sg13g2_o21ai_1 _32050_ (.B1(_20924_),
    .Y(_23489_),
    .A1(_21587_),
    .A2(_21619_));
 sg13g2_xnor2_1 _32051_ (.Y(_23490_),
    .A(_20923_),
    .B(_21620_));
 sg13g2_o21ai_1 _32052_ (.B1(_20923_),
    .Y(_23491_),
    .A1(_20085_),
    .A2(_20920_));
 sg13g2_nor3_1 _32053_ (.A(_20085_),
    .B(_20920_),
    .C(_20923_),
    .Y(_23492_));
 sg13g2_nor2_1 _32054_ (.A(net7184),
    .B(_23492_),
    .Y(_23493_));
 sg13g2_a221oi_1 _32055_ (.B2(_23493_),
    .C1(net6284),
    .B1(_23491_),
    .A1(\u_inv.f_next[192] ),
    .Y(_23494_),
    .A2(net7184));
 sg13g2_a21o_2 _32056_ (.A2(_23490_),
    .A1(net6284),
    .B1(_23494_),
    .X(_23495_));
 sg13g2_nor2_1 _32057_ (.A(_21517_),
    .B(_23486_),
    .Y(_23496_));
 sg13g2_a21oi_1 _32058_ (.A1(_20196_),
    .A2(_23496_),
    .Y(_23497_),
    .B1(net6236));
 sg13g2_o21ai_1 _32059_ (.B1(_23497_),
    .Y(_23498_),
    .A1(_20196_),
    .A2(_23496_));
 sg13g2_nand2_1 _32060_ (.Y(_23499_),
    .A(_20197_),
    .B(_23481_));
 sg13g2_xnor2_1 _32061_ (.Y(_23500_),
    .A(_20196_),
    .B(_23499_));
 sg13g2_a21oi_1 _32062_ (.A1(net7358),
    .A2(_23500_),
    .Y(_23501_),
    .B1(net6321));
 sg13g2_o21ai_1 _32063_ (.B1(_23501_),
    .Y(_23502_),
    .A1(\u_inv.f_next[147] ),
    .A2(net7358));
 sg13g2_nand2_2 _32064_ (.Y(_23503_),
    .A(_23498_),
    .B(_23502_));
 sg13g2_nor2b_1 _32065_ (.A(_21522_),
    .B_N(_22173_),
    .Y(_23504_));
 sg13g2_o21ai_1 _32066_ (.B1(net6320),
    .Y(_23505_),
    .A1(_20189_),
    .A2(_23504_));
 sg13g2_a21oi_1 _32067_ (.A1(_20189_),
    .A2(_23504_),
    .Y(_23506_),
    .B1(_23505_));
 sg13g2_o21ai_1 _32068_ (.B1(_20191_),
    .Y(_23507_),
    .A1(_20192_),
    .A2(_22163_));
 sg13g2_o21ai_1 _32069_ (.B1(net7359),
    .Y(_23508_),
    .A1(_20190_),
    .A2(_23507_));
 sg13g2_a21oi_1 _32070_ (.A1(_20190_),
    .A2(_23507_),
    .Y(_23509_),
    .B1(_23508_));
 sg13g2_o21ai_1 _32071_ (.B1(net6235),
    .Y(_23510_),
    .A1(\u_inv.f_next[151] ),
    .A2(net7359));
 sg13g2_nor2_1 _32072_ (.A(_23509_),
    .B(_23510_),
    .Y(_23511_));
 sg13g2_nor2_2 _32073_ (.A(_23506_),
    .B(_23511_),
    .Y(_23512_));
 sg13g2_nand3_1 _32074_ (.B(_21558_),
    .C(_22040_),
    .A(_20097_),
    .Y(_23513_));
 sg13g2_nor3_1 _32075_ (.A(net6213),
    .B(_21559_),
    .C(_22041_),
    .Y(_23514_));
 sg13g2_o21ai_1 _32076_ (.B1(_20092_),
    .Y(_23515_),
    .A1(_20095_),
    .A2(_22053_));
 sg13g2_xnor2_1 _32077_ (.Y(_23516_),
    .A(_20097_),
    .B(_23515_));
 sg13g2_o21ai_1 _32078_ (.B1(net6213),
    .Y(_23517_),
    .A1(\u_inv.f_next[173] ),
    .A2(net7325));
 sg13g2_a21oi_1 _32079_ (.A1(net7325),
    .A2(_23516_),
    .Y(_23518_),
    .B1(_23517_));
 sg13g2_a21o_2 _32080_ (.A2(_23514_),
    .A1(_23513_),
    .B1(_23518_),
    .X(_23519_));
 sg13g2_nand3_1 _32081_ (.B(_21673_),
    .C(_21915_),
    .A(_19956_),
    .Y(_23520_));
 sg13g2_and4_1 _32082_ (.A(net6275),
    .B(_21675_),
    .C(_21916_),
    .D(_23520_),
    .X(_23521_));
 sg13g2_o21ai_1 _32083_ (.B1(_19954_),
    .Y(_23522_),
    .A1(_19972_),
    .A2(_21924_));
 sg13g2_a21o_1 _32084_ (.A2(_23522_),
    .A1(_19953_),
    .B1(_19956_),
    .X(_23523_));
 sg13g2_nand3_1 _32085_ (.B(_19956_),
    .C(_23522_),
    .A(_19953_),
    .Y(_23524_));
 sg13g2_nand3_1 _32086_ (.B(_23523_),
    .C(_23524_),
    .A(net7303),
    .Y(_23525_));
 sg13g2_a21oi_1 _32087_ (.A1(_17988_),
    .A2(net7179),
    .Y(_23526_),
    .B1(net6275));
 sg13g2_a21o_2 _32088_ (.A2(_23526_),
    .A1(_23525_),
    .B1(_23521_),
    .X(_23527_));
 sg13g2_or3_1 _32089_ (.A(_19954_),
    .B(_19972_),
    .C(_21924_),
    .X(_23528_));
 sg13g2_nand2_1 _32090_ (.Y(_23529_),
    .A(_23522_),
    .B(_23528_));
 sg13g2_o21ai_1 _32091_ (.B1(net6193),
    .Y(_23530_),
    .A1(\u_inv.f_next[204] ),
    .A2(net7303));
 sg13g2_a21oi_1 _32092_ (.A1(net7308),
    .A2(_23529_),
    .Y(_23531_),
    .B1(_23530_));
 sg13g2_nor3_1 _32093_ (.A(_19955_),
    .B(_21672_),
    .C(_21914_),
    .Y(_23532_));
 sg13g2_nand3b_1 _32094_ (.B(net6275),
    .C(_21915_),
    .Y(_23533_),
    .A_N(_23532_));
 sg13g2_nor2b_2 _32095_ (.A(_23531_),
    .B_N(_23533_),
    .Y(_23534_));
 sg13g2_a21oi_1 _32096_ (.A1(_19994_),
    .A2(_22115_),
    .Y(_23535_),
    .B1(_19989_));
 sg13g2_nand3_1 _32097_ (.B(_19994_),
    .C(_22115_),
    .A(_19989_),
    .Y(_23536_));
 sg13g2_nand2b_1 _32098_ (.Y(_23537_),
    .B(_23536_),
    .A_N(_23535_));
 sg13g2_o21ai_1 _32099_ (.B1(net6197),
    .Y(_23538_),
    .A1(\u_inv.f_next[194] ),
    .A2(net7307));
 sg13g2_a21oi_1 _32100_ (.A1(net7307),
    .A2(_23537_),
    .Y(_23539_),
    .B1(_23538_));
 sg13g2_a21oi_1 _32101_ (.A1(_21653_),
    .A2(_23489_),
    .Y(_23540_),
    .B1(_20922_));
 sg13g2_nor3_1 _32102_ (.A(_19989_),
    .B(_21655_),
    .C(_23540_),
    .Y(_23541_));
 sg13g2_o21ai_1 _32103_ (.B1(_19989_),
    .Y(_23542_),
    .A1(_21655_),
    .A2(_23540_));
 sg13g2_nor2_1 _32104_ (.A(net6197),
    .B(_23541_),
    .Y(_23543_));
 sg13g2_a21o_2 _32105_ (.A2(_23543_),
    .A1(_23542_),
    .B1(_23539_),
    .X(_23544_));
 sg13g2_o21ai_1 _32106_ (.B1(_20077_),
    .Y(_23545_),
    .A1(_20036_),
    .A2(_21974_));
 sg13g2_xnor2_1 _32107_ (.Y(_23546_),
    .A(_20038_),
    .B(_23545_));
 sg13g2_o21ai_1 _32108_ (.B1(net6207),
    .Y(_23547_),
    .A1(\u_inv.f_next[186] ),
    .A2(net7318));
 sg13g2_a21oi_1 _32109_ (.A1(net7318),
    .A2(_23546_),
    .Y(_23548_),
    .B1(_23547_));
 sg13g2_o21ai_1 _32110_ (.B1(_20035_),
    .Y(_23549_),
    .A1(_21602_),
    .A2(_21981_));
 sg13g2_a21oi_1 _32111_ (.A1(_21610_),
    .A2(_23549_),
    .Y(_23550_),
    .B1(_20032_));
 sg13g2_o21ai_1 _32112_ (.B1(_20039_),
    .Y(_23551_),
    .A1(_21612_),
    .A2(_23550_));
 sg13g2_nor3_1 _32113_ (.A(_20039_),
    .B(_21612_),
    .C(_23550_),
    .Y(_23552_));
 sg13g2_nor2_1 _32114_ (.A(net6207),
    .B(_23552_),
    .Y(_23553_));
 sg13g2_a21o_2 _32115_ (.A2(_23553_),
    .A1(_23551_),
    .B1(_23548_),
    .X(_23554_));
 sg13g2_a21oi_1 _32116_ (.A1(_20166_),
    .A2(_23438_),
    .Y(_23555_),
    .B1(_20217_));
 sg13g2_o21ai_1 _32117_ (.B1(_20157_),
    .Y(_23556_),
    .A1(_20159_),
    .A2(_23555_));
 sg13g2_xnor2_1 _32118_ (.Y(_23557_),
    .A(_20156_),
    .B(_23556_));
 sg13g2_o21ai_1 _32119_ (.B1(net6232),
    .Y(_23558_),
    .A1(\u_inv.f_next[159] ),
    .A2(net7353));
 sg13g2_a21oi_1 _32120_ (.A1(net7353),
    .A2(_23557_),
    .Y(_23559_),
    .B1(_23558_));
 sg13g2_o21ai_1 _32121_ (.B1(_20159_),
    .Y(_23560_),
    .A1(_21498_),
    .A2(_23447_));
 sg13g2_and2_1 _32122_ (.A(_21527_),
    .B(_23560_),
    .X(_23561_));
 sg13g2_a21oi_1 _32123_ (.A1(_20156_),
    .A2(_23561_),
    .Y(_23562_),
    .B1(net6232));
 sg13g2_o21ai_1 _32124_ (.B1(_23562_),
    .Y(_23563_),
    .A1(_20156_),
    .A2(_23561_));
 sg13g2_nand2b_2 _32125_ (.Y(_23564_),
    .B(_23563_),
    .A_N(_23559_));
 sg13g2_xnor2_1 _32126_ (.Y(_23565_),
    .A(_20102_),
    .B(_22051_));
 sg13g2_nor2_1 _32127_ (.A(\u_inv.f_next[170] ),
    .B(net7326),
    .Y(_23566_));
 sg13g2_a21oi_1 _32128_ (.A1(net7328),
    .A2(_23565_),
    .Y(_23567_),
    .B1(_23566_));
 sg13g2_o21ai_1 _32129_ (.B1(_20112_),
    .Y(_23568_),
    .A1(_21571_),
    .A2(_22038_));
 sg13g2_a21o_1 _32130_ (.A2(_23568_),
    .A1(_21552_),
    .B1(_20109_),
    .X(_23569_));
 sg13g2_a21oi_1 _32131_ (.A1(_21553_),
    .A2(_23569_),
    .Y(_23570_),
    .B1(_20102_));
 sg13g2_nand3_1 _32132_ (.B(_21553_),
    .C(_23569_),
    .A(_20102_),
    .Y(_23571_));
 sg13g2_nor2_1 _32133_ (.A(net6214),
    .B(_23570_),
    .Y(_23572_));
 sg13g2_a22oi_1 _32134_ (.Y(_23573_),
    .B1(_23571_),
    .B2(_23572_),
    .A2(_23567_),
    .A1(net6214));
 sg13g2_inv_1 _32135_ (.Y(_23574_),
    .A(_23573_));
 sg13g2_nand3_1 _32136_ (.B(_21616_),
    .C(_21983_),
    .A(_20029_),
    .Y(_23575_));
 sg13g2_nand2b_1 _32137_ (.Y(_23576_),
    .B(_23575_),
    .A_N(_21984_));
 sg13g2_nor3_1 _32138_ (.A(_20029_),
    .B(_20081_),
    .C(_21975_),
    .Y(_23577_));
 sg13g2_nand3b_1 _32139_ (.B(net7314),
    .C(_21976_),
    .Y(_23578_),
    .A_N(_23577_));
 sg13g2_a21oi_1 _32140_ (.A1(\u_inv.f_next[188] ),
    .A2(net7184),
    .Y(_23579_),
    .B1(net6283));
 sg13g2_a22oi_1 _32141_ (.Y(_23580_),
    .B1(_23578_),
    .B2(_23579_),
    .A2(_23576_),
    .A1(net6283));
 sg13g2_nand3_1 _32142_ (.B(_21610_),
    .C(_23549_),
    .A(_20032_),
    .Y(_23581_));
 sg13g2_nor2_1 _32143_ (.A(net6207),
    .B(_23550_),
    .Y(_23582_));
 sg13g2_o21ai_1 _32144_ (.B1(_20034_),
    .Y(_23583_),
    .A1(_20035_),
    .A2(_21974_));
 sg13g2_xnor2_1 _32145_ (.Y(_23584_),
    .A(_20032_),
    .B(_23583_));
 sg13g2_o21ai_1 _32146_ (.B1(net6207),
    .Y(_23585_),
    .A1(\u_inv.f_next[185] ),
    .A2(net7318));
 sg13g2_a21oi_1 _32147_ (.A1(net7318),
    .A2(_23584_),
    .Y(_23586_),
    .B1(_23585_));
 sg13g2_a21o_2 _32148_ (.A2(_23582_),
    .A1(_23581_),
    .B1(_23586_),
    .X(_23587_));
 sg13g2_nand3_1 _32149_ (.B(_21648_),
    .C(_21715_),
    .A(_20953_),
    .Y(_23588_));
 sg13g2_nor2b_1 _32150_ (.A(_22086_),
    .B_N(_23588_),
    .Y(_23589_));
 sg13g2_and2_1 _32151_ (.A(_20933_),
    .B(_20953_),
    .X(_23590_));
 sg13g2_o21ai_1 _32152_ (.B1(net7304),
    .Y(_23591_),
    .A1(_20933_),
    .A2(_20953_));
 sg13g2_nand2_1 _32153_ (.Y(_23592_),
    .A(\u_inv.f_next[224] ),
    .B(net7177));
 sg13g2_o21ai_1 _32154_ (.B1(_23592_),
    .Y(_23593_),
    .A1(_23590_),
    .A2(_23591_));
 sg13g2_mux2_1 _32155_ (.A0(_23589_),
    .A1(_23593_),
    .S(net6195),
    .X(_23594_));
 sg13g2_nand3_1 _32156_ (.B(_20009_),
    .C(_21921_),
    .A(_20006_),
    .Y(_23595_));
 sg13g2_nand2b_1 _32157_ (.Y(_23596_),
    .B(_23595_),
    .A_N(_21922_));
 sg13g2_o21ai_1 _32158_ (.B1(net6198),
    .Y(_23597_),
    .A1(\u_inv.f_next[200] ),
    .A2(net7308));
 sg13g2_a21oi_1 _32159_ (.A1(net7308),
    .A2(_23596_),
    .Y(_23598_),
    .B1(_23597_));
 sg13g2_nand3_1 _32160_ (.B(_21665_),
    .C(_21912_),
    .A(_20008_),
    .Y(_23599_));
 sg13g2_nor2_1 _32161_ (.A(net6198),
    .B(_21913_),
    .Y(_23600_));
 sg13g2_a21o_2 _32162_ (.A2(_23600_),
    .A1(_23599_),
    .B1(_23598_),
    .X(_23601_));
 sg13g2_nand3_1 _32163_ (.B(_21552_),
    .C(_23568_),
    .A(_20109_),
    .Y(_23602_));
 sg13g2_nand3_1 _32164_ (.B(_23569_),
    .C(_23602_),
    .A(net6298),
    .Y(_23603_));
 sg13g2_o21ai_1 _32165_ (.B1(_20111_),
    .Y(_23604_),
    .A1(_20126_),
    .A2(_22048_));
 sg13g2_a21oi_1 _32166_ (.A1(_20110_),
    .A2(_23604_),
    .Y(_23605_),
    .B1(_20109_));
 sg13g2_and3_1 _32167_ (.X(_23606_),
    .A(_20109_),
    .B(_20110_),
    .C(_23604_));
 sg13g2_nor3_1 _32168_ (.A(net7197),
    .B(_23605_),
    .C(_23606_),
    .Y(_23607_));
 sg13g2_o21ai_1 _32169_ (.B1(net6217),
    .Y(_23608_),
    .A1(\u_inv.f_next[169] ),
    .A2(net7328));
 sg13g2_o21ai_1 _32170_ (.B1(_23603_),
    .Y(_23609_),
    .A1(_23607_),
    .A2(_23608_));
 sg13g2_xnor2_1 _32171_ (.Y(_23610_),
    .A(_20035_),
    .B(_21974_));
 sg13g2_o21ai_1 _32172_ (.B1(net6207),
    .Y(_23611_),
    .A1(\u_inv.f_next[184] ),
    .A2(net7318));
 sg13g2_a21oi_1 _32173_ (.A1(net7318),
    .A2(_23610_),
    .Y(_23612_),
    .B1(_23611_));
 sg13g2_xnor2_1 _32174_ (.Y(_23613_),
    .A(_20035_),
    .B(_21982_));
 sg13g2_a21oi_2 _32175_ (.B1(_23612_),
    .Y(_23614_),
    .A2(_23613_),
    .A1(net6286));
 sg13g2_xnor2_1 _32176_ (.Y(_23615_),
    .A(_20112_),
    .B(_22049_));
 sg13g2_o21ai_1 _32177_ (.B1(net6217),
    .Y(_23616_),
    .A1(\u_inv.f_next[168] ),
    .A2(net7328));
 sg13g2_a21oi_1 _32178_ (.A1(net7328),
    .A2(_23615_),
    .Y(_23617_),
    .B1(_23616_));
 sg13g2_or3_1 _32179_ (.A(_20112_),
    .B(_21571_),
    .C(_22038_),
    .X(_23618_));
 sg13g2_and2_1 _32180_ (.A(net6298),
    .B(_23568_),
    .X(_23619_));
 sg13g2_a21oi_2 _32181_ (.B1(_23617_),
    .Y(_23620_),
    .A2(_23619_),
    .A1(_23618_));
 sg13g2_or3_1 _32182_ (.A(_20052_),
    .B(_21594_),
    .C(_22003_),
    .X(_23621_));
 sg13g2_and2_1 _32183_ (.A(net6287),
    .B(_22004_),
    .X(_23622_));
 sg13g2_o21ai_1 _32184_ (.B1(_20051_),
    .Y(_23623_),
    .A1(_20067_),
    .A2(_21972_));
 sg13g2_xnor2_1 _32185_ (.Y(_23624_),
    .A(_20052_),
    .B(_21973_));
 sg13g2_nor2_1 _32186_ (.A(\u_inv.f_next[180] ),
    .B(net7317),
    .Y(_23625_));
 sg13g2_a21oi_1 _32187_ (.A1(net7317),
    .A2(_23624_),
    .Y(_23626_),
    .B1(_23625_));
 sg13g2_a22oi_1 _32188_ (.Y(_23627_),
    .B1(_23626_),
    .B2(net6207),
    .A2(_23622_),
    .A1(_23621_));
 sg13g2_xnor2_1 _32189_ (.Y(_23628_),
    .A(_20159_),
    .B(_23555_));
 sg13g2_a21oi_1 _32190_ (.A1(net7354),
    .A2(_23628_),
    .Y(_23629_),
    .B1(net6318));
 sg13g2_o21ai_1 _32191_ (.B1(_23629_),
    .Y(_23630_),
    .A1(\u_inv.f_next[158] ),
    .A2(net7353));
 sg13g2_nor3_1 _32192_ (.A(_20159_),
    .B(_21498_),
    .C(_23447_),
    .Y(_23631_));
 sg13g2_nand2_1 _32193_ (.Y(_23632_),
    .A(net6318),
    .B(_23560_));
 sg13g2_o21ai_1 _32194_ (.B1(_23630_),
    .Y(_23633_),
    .A1(_23631_),
    .A2(_23632_));
 sg13g2_xnor2_1 _32195_ (.Y(_23634_),
    .A(_20059_),
    .B(_22070_));
 sg13g2_a21oi_1 _32196_ (.A1(net7326),
    .A2(_23634_),
    .Y(_23635_),
    .B1(net6297));
 sg13g2_o21ai_1 _32197_ (.B1(_23635_),
    .Y(_23636_),
    .A1(\u_inv.f_next[178] ),
    .A2(net7324));
 sg13g2_nand3_1 _32198_ (.B(_21591_),
    .C(_22076_),
    .A(_20058_),
    .Y(_23637_));
 sg13g2_nand2_1 _32199_ (.Y(_23638_),
    .A(net6297),
    .B(_23637_));
 sg13g2_o21ai_1 _32200_ (.B1(_23636_),
    .Y(_23639_),
    .A1(_22077_),
    .A2(_23638_));
 sg13g2_xnor2_1 _32201_ (.Y(_23640_),
    .A(_20118_),
    .B(_22102_));
 sg13g2_nor2_1 _32202_ (.A(\u_inv.f_next[166] ),
    .B(net7329),
    .Y(_23641_));
 sg13g2_o21ai_1 _32203_ (.B1(net6217),
    .Y(_23642_),
    .A1(net7197),
    .A2(_23640_));
 sg13g2_nand3b_1 _32204_ (.B(_20118_),
    .C(_21568_),
    .Y(_23643_),
    .A_N(_22108_));
 sg13g2_nand3_1 _32205_ (.B(_22109_),
    .C(_23643_),
    .A(net6298),
    .Y(_23644_));
 sg13g2_o21ai_1 _32206_ (.B1(_23644_),
    .Y(_23645_),
    .A1(_23641_),
    .A2(_23642_));
 sg13g2_nor3_1 _32207_ (.A(_20955_),
    .B(_21731_),
    .C(_22086_),
    .Y(_23646_));
 sg13g2_nand2_1 _32208_ (.Y(_23647_),
    .A(net6276),
    .B(_21732_));
 sg13g2_nor3_1 _32209_ (.A(_22087_),
    .B(_23646_),
    .C(_23647_),
    .Y(_23648_));
 sg13g2_a21oi_1 _32210_ (.A1(_20933_),
    .A2(_20953_),
    .Y(_23649_),
    .B1(_20952_));
 sg13g2_xnor2_1 _32211_ (.Y(_23650_),
    .A(_20955_),
    .B(_23649_));
 sg13g2_o21ai_1 _32212_ (.B1(net6195),
    .Y(_01901_),
    .A1(\u_inv.f_next[225] ),
    .A2(net7304));
 sg13g2_a21oi_1 _32213_ (.A1(net7304),
    .A2(_23650_),
    .Y(_01902_),
    .B1(_01901_));
 sg13g2_nor2_2 _32214_ (.A(_23648_),
    .B(_01902_),
    .Y(_01903_));
 sg13g2_inv_1 _32215_ (.Y(_01904_),
    .A(_01903_));
 sg13g2_and2_1 _32216_ (.A(_20175_),
    .B(_23420_),
    .X(_01905_));
 sg13g2_o21ai_1 _32217_ (.B1(net7357),
    .Y(_01906_),
    .A1(_20178_),
    .A2(_01905_));
 sg13g2_a21oi_1 _32218_ (.A1(_20178_),
    .A2(_01905_),
    .Y(_01907_),
    .B1(_01906_));
 sg13g2_o21ai_1 _32219_ (.B1(net6234),
    .Y(_01908_),
    .A1(\u_inv.f_next[155] ),
    .A2(net7354));
 sg13g2_nor2_1 _32220_ (.A(_21500_),
    .B(_23425_),
    .Y(_01909_));
 sg13g2_o21ai_1 _32221_ (.B1(net6320),
    .Y(_01910_),
    .A1(_20178_),
    .A2(_01909_));
 sg13g2_a21o_1 _32222_ (.A2(_01909_),
    .A1(_20178_),
    .B1(_01910_),
    .X(_01911_));
 sg13g2_o21ai_1 _32223_ (.B1(_01911_),
    .Y(_01912_),
    .A1(_01907_),
    .A2(_01908_));
 sg13g2_o21ai_1 _32224_ (.B1(_23491_),
    .Y(_01913_),
    .A1(_17997_),
    .A2(_18242_));
 sg13g2_xnor2_1 _32225_ (.Y(_01914_),
    .A(_20922_),
    .B(_01913_));
 sg13g2_o21ai_1 _32226_ (.B1(net6205),
    .Y(_01915_),
    .A1(\u_inv.f_next[193] ),
    .A2(net7315));
 sg13g2_a21o_1 _32227_ (.A2(_01914_),
    .A1(net7315),
    .B1(_01915_),
    .X(_01916_));
 sg13g2_nand3_1 _32228_ (.B(_21653_),
    .C(_23489_),
    .A(_20922_),
    .Y(_01917_));
 sg13g2_nand2_1 _32229_ (.Y(_01918_),
    .A(net6278),
    .B(_01917_));
 sg13g2_o21ai_1 _32230_ (.B1(_01916_),
    .Y(_01919_),
    .A1(_23540_),
    .A2(_01918_));
 sg13g2_nand3_1 _32231_ (.B(_21681_),
    .C(_21822_),
    .A(_19939_),
    .Y(_01920_));
 sg13g2_nand2b_1 _32232_ (.Y(_01921_),
    .B(_01920_),
    .A_N(_22015_));
 sg13g2_nor2_1 _32233_ (.A(net7179),
    .B(_22010_),
    .Y(_01922_));
 sg13g2_o21ai_1 _32234_ (.B1(_01922_),
    .Y(_01923_),
    .A1(_19939_),
    .A2(_20929_));
 sg13g2_a21oi_1 _32235_ (.A1(\u_inv.f_next[208] ),
    .A2(net7179),
    .Y(_01924_),
    .B1(net6274));
 sg13g2_a22oi_1 _32236_ (.Y(_01925_),
    .B1(_01923_),
    .B2(_01924_),
    .A2(_01921_),
    .A1(net6274));
 sg13g2_or3_1 _32237_ (.A(_19985_),
    .B(_19997_),
    .C(_22116_),
    .X(_01926_));
 sg13g2_a21oi_1 _32238_ (.A1(_22117_),
    .A2(_01926_),
    .Y(_01927_),
    .B1(net7180));
 sg13g2_o21ai_1 _32239_ (.B1(net6198),
    .Y(_01928_),
    .A1(\u_inv.f_next[196] ),
    .A2(net7307));
 sg13g2_nor2_1 _32240_ (.A(net6197),
    .B(_22124_),
    .Y(_01929_));
 sg13g2_o21ai_1 _32241_ (.B1(_01929_),
    .Y(_01930_),
    .A1(_19986_),
    .A2(_22123_));
 sg13g2_o21ai_1 _32242_ (.B1(_01930_),
    .Y(_01931_),
    .A1(_01927_),
    .A2(_01928_));
 sg13g2_xnor2_1 _32243_ (.Y(_01932_),
    .A(_20095_),
    .B(_22053_));
 sg13g2_o21ai_1 _32244_ (.B1(net6213),
    .Y(_01933_),
    .A1(\u_inv.f_next[172] ),
    .A2(net7325));
 sg13g2_a21oi_1 _32245_ (.A1(net7325),
    .A2(_01932_),
    .Y(_01934_),
    .B1(_01933_));
 sg13g2_nand3_1 _32246_ (.B(_21556_),
    .C(_22039_),
    .A(_20096_),
    .Y(_01935_));
 sg13g2_and2_1 _32247_ (.A(net6297),
    .B(_01935_),
    .X(_01936_));
 sg13g2_a21o_2 _32248_ (.A2(_01936_),
    .A1(_22040_),
    .B1(_01934_),
    .X(_01937_));
 sg13g2_a21oi_1 _32249_ (.A1(_20050_),
    .A2(_23623_),
    .Y(_01938_),
    .B1(_20054_));
 sg13g2_and3_1 _32250_ (.X(_01939_),
    .A(_20050_),
    .B(_20054_),
    .C(_23623_));
 sg13g2_nor3_1 _32251_ (.A(net7186),
    .B(_01938_),
    .C(_01939_),
    .Y(_01940_));
 sg13g2_o21ai_1 _32252_ (.B1(net6207),
    .Y(_01941_),
    .A1(\u_inv.f_next[181] ),
    .A2(net7317));
 sg13g2_nand3_1 _32253_ (.B(_21595_),
    .C(_22004_),
    .A(_20054_),
    .Y(_01942_));
 sg13g2_nand3b_1 _32254_ (.B(_01942_),
    .C(net6287),
    .Y(_01943_),
    .A_N(_22005_));
 sg13g2_o21ai_1 _32255_ (.B1(_01943_),
    .Y(_01944_),
    .A1(_01940_),
    .A2(_01941_));
 sg13g2_nand3_1 _32256_ (.B(_21009_),
    .C(_21866_),
    .A(_20985_),
    .Y(_01945_));
 sg13g2_a21o_1 _32257_ (.A2(_01945_),
    .A1(_21867_),
    .B1(net7182),
    .X(_01946_));
 sg13g2_a21oi_1 _32258_ (.A1(_17971_),
    .A2(net7182),
    .Y(_01947_),
    .B1(net6279));
 sg13g2_nor3_1 _32259_ (.A(_20985_),
    .B(_21754_),
    .C(_21875_),
    .Y(_01948_));
 sg13g2_nor2_1 _32260_ (.A(net6199),
    .B(_01948_),
    .Y(_01949_));
 sg13g2_a22oi_1 _32261_ (.Y(_01950_),
    .B1(_01949_),
    .B2(_21876_),
    .A2(_01947_),
    .A1(_01946_));
 sg13g2_o21ai_1 _32262_ (.B1(_21044_),
    .Y(_01951_),
    .A1(_21770_),
    .A2(_21949_));
 sg13g2_or3_1 _32263_ (.A(_21044_),
    .B(_21770_),
    .C(_21949_),
    .X(_01952_));
 sg13g2_nand3_1 _32264_ (.B(_01951_),
    .C(_01952_),
    .A(net6279),
    .Y(_01953_));
 sg13g2_nor2_1 _32265_ (.A(_21041_),
    .B(_21941_),
    .Y(_01954_));
 sg13g2_xor2_1 _32266_ (.B(_01954_),
    .A(_21044_),
    .X(_01955_));
 sg13g2_a21oi_1 _32267_ (.A1(_17968_),
    .A2(net7182),
    .Y(_01956_),
    .B1(net6279));
 sg13g2_o21ai_1 _32268_ (.B1(_01956_),
    .Y(_01957_),
    .A1(net7182),
    .A2(_01955_));
 sg13g2_nand2_1 _32269_ (.Y(_01958_),
    .A(_01953_),
    .B(_01957_));
 sg13g2_a21o_1 _32270_ (.A2(_21814_),
    .A1(_19937_),
    .B1(_19906_),
    .X(_01959_));
 sg13g2_a21oi_1 _32271_ (.A1(_19894_),
    .A2(_01959_),
    .Y(_01960_),
    .B1(_19881_));
 sg13g2_o21ai_1 _32272_ (.B1(_19873_),
    .Y(_01961_),
    .A1(_19896_),
    .A2(_01960_));
 sg13g2_nand3_1 _32273_ (.B(_19872_),
    .C(_01961_),
    .A(_19871_),
    .Y(_01962_));
 sg13g2_a21o_1 _32274_ (.A2(_01961_),
    .A1(_19872_),
    .B1(_19871_),
    .X(_01963_));
 sg13g2_nand3_1 _32275_ (.B(_01962_),
    .C(_01963_),
    .A(net7304),
    .Y(_01964_));
 sg13g2_a21oi_1 _32276_ (.A1(_17977_),
    .A2(net7177),
    .Y(_01965_),
    .B1(net6276));
 sg13g2_o21ai_1 _32277_ (.B1(_21630_),
    .Y(_01966_),
    .A1(_21714_),
    .A2(_21823_));
 sg13g2_a21oi_1 _32278_ (.A1(_21690_),
    .A2(_01966_),
    .Y(_01967_),
    .B1(_21627_));
 sg13g2_o21ai_1 _32279_ (.B1(_19874_),
    .Y(_01968_),
    .A1(_21694_),
    .A2(_01967_));
 sg13g2_a21oi_1 _32280_ (.A1(_21696_),
    .A2(_01968_),
    .Y(_01969_),
    .B1(_19871_));
 sg13g2_nand3_1 _32281_ (.B(_21696_),
    .C(_01968_),
    .A(_19871_),
    .Y(_01970_));
 sg13g2_nor2_1 _32282_ (.A(net6195),
    .B(_01969_),
    .Y(_01971_));
 sg13g2_a22oi_1 _32283_ (.Y(_01972_),
    .B1(_01970_),
    .B2(_01971_),
    .A2(_01965_),
    .A1(_01964_));
 sg13g2_o21ai_1 _32284_ (.B1(_19920_),
    .Y(_01973_),
    .A1(_19922_),
    .A2(_22129_));
 sg13g2_and2_1 _32285_ (.A(_19924_),
    .B(_01973_),
    .X(_01974_));
 sg13g2_o21ai_1 _32286_ (.B1(net7301),
    .Y(_01975_),
    .A1(_19924_),
    .A2(_01973_));
 sg13g2_a21oi_1 _32287_ (.A1(_17985_),
    .A2(net7179),
    .Y(_01976_),
    .B1(net6274));
 sg13g2_o21ai_1 _32288_ (.B1(_01976_),
    .Y(_01977_),
    .A1(_01974_),
    .A2(_01975_));
 sg13g2_a21oi_1 _32289_ (.A1(_21702_),
    .A2(_22017_),
    .Y(_01978_),
    .B1(_19921_));
 sg13g2_nor2_1 _32290_ (.A(_21704_),
    .B(_01978_),
    .Y(_01979_));
 sg13g2_xor2_1 _32291_ (.B(_01979_),
    .A(_19924_),
    .X(_01980_));
 sg13g2_o21ai_1 _32292_ (.B1(_01977_),
    .Y(_01981_),
    .A1(net6192),
    .A2(_01980_));
 sg13g2_xnor2_1 _32293_ (.Y(_01982_),
    .A(_19884_),
    .B(_21816_));
 sg13g2_o21ai_1 _32294_ (.B1(net6196),
    .Y(_01983_),
    .A1(\u_inv.f_next[218] ),
    .A2(net7306));
 sg13g2_a21oi_1 _32295_ (.A1(net7306),
    .A2(_01982_),
    .Y(_01984_),
    .B1(_01983_));
 sg13g2_nor3_1 _32296_ (.A(_19885_),
    .B(_21687_),
    .C(_21825_),
    .Y(_01985_));
 sg13g2_nor2_1 _32297_ (.A(net6196),
    .B(_01985_),
    .Y(_01986_));
 sg13g2_a21o_2 _32298_ (.A2(_01986_),
    .A1(_21826_),
    .B1(_01984_),
    .X(_01987_));
 sg13g2_o21ai_1 _32299_ (.B1(_19918_),
    .Y(_01988_),
    .A1(_19930_),
    .A2(_22130_));
 sg13g2_a21oi_1 _32300_ (.A1(_19933_),
    .A2(_01988_),
    .Y(_01989_),
    .B1(_19910_));
 sg13g2_o21ai_1 _32301_ (.B1(_19912_),
    .Y(_01990_),
    .A1(_19908_),
    .A2(_01989_));
 sg13g2_or3_1 _32302_ (.A(_19908_),
    .B(_19912_),
    .C(_01989_),
    .X(_01991_));
 sg13g2_and3_1 _32303_ (.X(_01992_),
    .A(net7301),
    .B(_01990_),
    .C(_01991_));
 sg13g2_o21ai_1 _32304_ (.B1(net6192),
    .Y(_01993_),
    .A1(\u_inv.f_next[215] ),
    .A2(net7301));
 sg13g2_a21oi_1 _32305_ (.A1(_21709_),
    .A2(_22147_),
    .Y(_01994_),
    .B1(_19909_));
 sg13g2_or3_1 _32306_ (.A(_19912_),
    .B(_21710_),
    .C(_01994_),
    .X(_01995_));
 sg13g2_o21ai_1 _32307_ (.B1(_19912_),
    .Y(_01996_),
    .A1(_21710_),
    .A2(_01994_));
 sg13g2_nand3_1 _32308_ (.B(_01995_),
    .C(_01996_),
    .A(net6274),
    .Y(_01997_));
 sg13g2_o21ai_1 _32309_ (.B1(_01997_),
    .Y(_01998_),
    .A1(_01992_),
    .A2(_01993_));
 sg13g2_nor3_1 _32310_ (.A(_21038_),
    .B(_21053_),
    .C(_21800_),
    .Y(_01999_));
 sg13g2_nand2_1 _32311_ (.Y(_02000_),
    .A(net7311),
    .B(_21801_));
 sg13g2_nand2_1 _32312_ (.Y(_02001_),
    .A(\u_inv.f_next[246] ),
    .B(net7181));
 sg13g2_o21ai_1 _32313_ (.B1(_02001_),
    .Y(_02002_),
    .A1(_01999_),
    .A2(_02000_));
 sg13g2_nand3_1 _32314_ (.B(_21778_),
    .C(_21808_),
    .A(_21038_),
    .Y(_02003_));
 sg13g2_nor2_1 _32315_ (.A(net6201),
    .B(_21809_),
    .Y(_02004_));
 sg13g2_a22oi_1 _32316_ (.Y(_02005_),
    .B1(_02003_),
    .B2(_02004_),
    .A2(_02002_),
    .A1(net6201));
 sg13g2_and3_1 _32317_ (.X(_02006_),
    .A(_19847_),
    .B(_19851_),
    .C(_21069_));
 sg13g2_o21ai_1 _32318_ (.B1(net7312),
    .Y(_02007_),
    .A1(_21070_),
    .A2(_02006_));
 sg13g2_a21oi_1 _32319_ (.A1(_17962_),
    .A2(net7181),
    .Y(_02008_),
    .B1(net6281));
 sg13g2_nand3_1 _32320_ (.B(_21080_),
    .C(_21792_),
    .A(_19846_),
    .Y(_02009_));
 sg13g2_nor2_1 _32321_ (.A(net6203),
    .B(_21793_),
    .Y(_02010_));
 sg13g2_a22oi_1 _32322_ (.Y(_02011_),
    .B1(_02009_),
    .B2(_02010_),
    .A2(_02008_),
    .A1(_02007_));
 sg13g2_nand3_1 _32323_ (.B(_21007_),
    .C(_21854_),
    .A(_20969_),
    .Y(_02012_));
 sg13g2_nand2b_1 _32324_ (.Y(_02013_),
    .B(_02012_),
    .A_N(_21855_));
 sg13g2_o21ai_1 _32325_ (.B1(net6199),
    .Y(_02014_),
    .A1(\u_inv.f_next[234] ),
    .A2(net7309));
 sg13g2_a21oi_1 _32326_ (.A1(net7309),
    .A2(_02013_),
    .Y(_02015_),
    .B1(_02014_));
 sg13g2_nor3_1 _32327_ (.A(_20969_),
    .B(_21746_),
    .C(_21846_),
    .Y(_02016_));
 sg13g2_nor2_1 _32328_ (.A(net6194),
    .B(_02016_),
    .Y(_02017_));
 sg13g2_a21o_2 _32329_ (.A2(_02017_),
    .A1(_21847_),
    .B1(_02015_),
    .X(_02018_));
 sg13g2_nand3_1 _32330_ (.B(_20949_),
    .C(_22083_),
    .A(_20948_),
    .Y(_02019_));
 sg13g2_a21oi_1 _32331_ (.A1(_20949_),
    .A2(_22083_),
    .Y(_02020_),
    .B1(_20948_));
 sg13g2_nor2_1 _32332_ (.A(net7177),
    .B(_02020_),
    .Y(_02021_));
 sg13g2_o21ai_1 _32333_ (.B1(net6194),
    .Y(_02022_),
    .A1(\u_inv.f_next[227] ),
    .A2(net7305));
 sg13g2_a21o_1 _32334_ (.A2(_02021_),
    .A1(_02019_),
    .B1(_02022_),
    .X(_02023_));
 sg13g2_or2_1 _32335_ (.X(_02024_),
    .B(_22089_),
    .A(_21730_));
 sg13g2_xor2_1 _32336_ (.B(_02024_),
    .A(_20948_),
    .X(_02025_));
 sg13g2_o21ai_1 _32337_ (.B1(_02023_),
    .Y(_02026_),
    .A1(net6195),
    .A2(_02025_));
 sg13g2_o21ai_1 _32338_ (.B1(_20938_),
    .Y(_02027_),
    .A1(_20996_),
    .A2(_21962_));
 sg13g2_a21oi_1 _32339_ (.A1(_21000_),
    .A2(_02027_),
    .Y(_02028_),
    .B1(_20941_));
 sg13g2_nand3_1 _32340_ (.B(_21000_),
    .C(_02027_),
    .A(_20941_),
    .Y(_02029_));
 sg13g2_nand2b_1 _32341_ (.Y(_02030_),
    .B(_02029_),
    .A_N(_02028_));
 sg13g2_o21ai_1 _32342_ (.B1(net6196),
    .Y(_02031_),
    .A1(\u_inv.f_next[230] ),
    .A2(net7305));
 sg13g2_a21oi_1 _32343_ (.A1(net7306),
    .A2(_02030_),
    .Y(_02032_),
    .B1(_02031_));
 sg13g2_o21ai_1 _32344_ (.B1(_21741_),
    .Y(_02033_),
    .A1(_20934_),
    .A2(_21969_));
 sg13g2_a21oi_1 _32345_ (.A1(_20941_),
    .A2(_02033_),
    .Y(_02034_),
    .B1(net6196));
 sg13g2_o21ai_1 _32346_ (.B1(_02034_),
    .Y(_02035_),
    .A1(_20941_),
    .A2(_02033_));
 sg13g2_nand2b_2 _32347_ (.Y(_02036_),
    .B(_02035_),
    .A_N(_02032_));
 sg13g2_and3_1 _32348_ (.X(_02037_),
    .A(_20087_),
    .B(_20089_),
    .C(_22055_));
 sg13g2_a21oi_1 _32349_ (.A1(_20089_),
    .A2(_22055_),
    .Y(_02038_),
    .B1(_20087_));
 sg13g2_nor3_1 _32350_ (.A(net7196),
    .B(_02037_),
    .C(_02038_),
    .Y(_02039_));
 sg13g2_o21ai_1 _32351_ (.B1(net6214),
    .Y(_02040_),
    .A1(\u_inv.f_next[175] ),
    .A2(net7326));
 sg13g2_nand3_1 _32352_ (.B(_21563_),
    .C(_22042_),
    .A(_20087_),
    .Y(_02041_));
 sg13g2_a21o_1 _32353_ (.A2(_22042_),
    .A1(_21563_),
    .B1(_20087_),
    .X(_02042_));
 sg13g2_nand3_1 _32354_ (.B(_02041_),
    .C(_02042_),
    .A(net6297),
    .Y(_02043_));
 sg13g2_o21ai_1 _32355_ (.B1(_02043_),
    .Y(_02044_),
    .A1(_02039_),
    .A2(_02040_));
 sg13g2_o21ai_1 _32356_ (.B1(_19854_),
    .Y(_02045_),
    .A1(_19869_),
    .A2(_21068_));
 sg13g2_and3_1 _32357_ (.X(_02046_),
    .A(_19849_),
    .B(_19852_),
    .C(_02045_));
 sg13g2_a21oi_1 _32358_ (.A1(_19849_),
    .A2(_02045_),
    .Y(_02047_),
    .B1(_19852_));
 sg13g2_nor3_1 _32359_ (.A(net7183),
    .B(_02046_),
    .C(_02047_),
    .Y(_02048_));
 sg13g2_o21ai_1 _32360_ (.B1(net6203),
    .Y(_02049_),
    .A1(\u_inv.f_next[253] ),
    .A2(net7312));
 sg13g2_o21ai_1 _32361_ (.B1(_19855_),
    .Y(_02050_),
    .A1(_21088_),
    .A2(_21791_));
 sg13g2_inv_1 _32362_ (.Y(_02051_),
    .A(_02050_));
 sg13g2_nand3_1 _32363_ (.B(_21077_),
    .C(_02050_),
    .A(_19852_),
    .Y(_02052_));
 sg13g2_nand4_1 _32364_ (.B(_21078_),
    .C(_21792_),
    .A(net6281),
    .Y(_02053_),
    .D(_02052_));
 sg13g2_o21ai_1 _32365_ (.B1(_02053_),
    .Y(_02054_),
    .A1(_02048_),
    .A2(_02049_));
 sg13g2_nor3_1 _32366_ (.A(_20975_),
    .B(_20977_),
    .C(_21934_),
    .Y(_02055_));
 sg13g2_o21ai_1 _32367_ (.B1(_20975_),
    .Y(_02056_),
    .A1(_20977_),
    .A2(_21934_));
 sg13g2_nand3b_1 _32368_ (.B(_02056_),
    .C(net7310),
    .Y(_02057_),
    .A_N(_02055_));
 sg13g2_o21ai_1 _32369_ (.B1(net6199),
    .Y(_02058_),
    .A1(\u_inv.f_next[237] ),
    .A2(net7309));
 sg13g2_inv_1 _32370_ (.Y(_02059_),
    .A(_02058_));
 sg13g2_nor3_1 _32371_ (.A(_20975_),
    .B(_21751_),
    .C(_21874_),
    .Y(_02060_));
 sg13g2_nor4_1 _32372_ (.A(net6199),
    .B(_21752_),
    .C(_21875_),
    .D(_02060_),
    .Y(_02061_));
 sg13g2_a21oi_2 _32373_ (.B1(_02061_),
    .Y(_02062_),
    .A2(_02059_),
    .A1(_02057_));
 sg13g2_a21o_1 _32374_ (.A2(_02059_),
    .A1(_02057_),
    .B1(_02061_),
    .X(_02063_));
 sg13g2_a21oi_1 _32375_ (.A1(_21050_),
    .A2(_21062_),
    .Y(_02064_),
    .B1(_21064_));
 sg13g2_nor3_1 _32376_ (.A(_21049_),
    .B(_21061_),
    .C(_21063_),
    .Y(_02065_));
 sg13g2_o21ai_1 _32377_ (.B1(net7311),
    .Y(_02066_),
    .A1(_02064_),
    .A2(_02065_));
 sg13g2_nand2_1 _32378_ (.Y(_02067_),
    .A(_17965_),
    .B(net7181));
 sg13g2_nand3_1 _32379_ (.B(_02066_),
    .C(_02067_),
    .A(net6201),
    .Y(_02068_));
 sg13g2_a21oi_1 _32380_ (.A1(_21063_),
    .A2(_21786_),
    .Y(_02069_),
    .B1(net6201));
 sg13g2_o21ai_1 _32381_ (.B1(_02069_),
    .Y(_02070_),
    .A1(_21063_),
    .A2(_21786_));
 sg13g2_nand2_1 _32382_ (.Y(_02071_),
    .A(_02068_),
    .B(_02070_));
 sg13g2_a21oi_1 _32383_ (.A1(_20047_),
    .A2(_21999_),
    .Y(_02072_),
    .B1(_20046_));
 sg13g2_a21oi_1 _32384_ (.A1(_20045_),
    .A2(_02072_),
    .Y(_02073_),
    .B1(net7186));
 sg13g2_o21ai_1 _32385_ (.B1(_02073_),
    .Y(_02074_),
    .A1(_20045_),
    .A2(_02072_));
 sg13g2_a21oi_1 _32386_ (.A1(_18005_),
    .A2(net7186),
    .Y(_02075_),
    .B1(net6286));
 sg13g2_a21o_1 _32387_ (.A2(_22007_),
    .A1(_21597_),
    .B1(_20045_),
    .X(_02076_));
 sg13g2_nand3_1 _32388_ (.B(_21597_),
    .C(_22007_),
    .A(_20045_),
    .Y(_02077_));
 sg13g2_and2_1 _32389_ (.A(net6286),
    .B(_02077_),
    .X(_02078_));
 sg13g2_and2_1 _32390_ (.A(_02076_),
    .B(_02078_),
    .X(_02079_));
 sg13g2_a22oi_1 _32391_ (.Y(_02080_),
    .B1(_02076_),
    .B2(_02078_),
    .A2(_02075_),
    .A1(_02074_));
 sg13g2_a21o_1 _32392_ (.A2(_02075_),
    .A1(_02074_),
    .B1(_02079_),
    .X(_02081_));
 sg13g2_nand3_1 _32393_ (.B(_21744_),
    .C(_21845_),
    .A(_20965_),
    .Y(_02082_));
 sg13g2_nand3b_1 _32394_ (.B(_02082_),
    .C(net6276),
    .Y(_02083_),
    .A_N(_21846_));
 sg13g2_and3_1 _32395_ (.X(_02084_),
    .A(_20960_),
    .B(_20965_),
    .C(_22061_));
 sg13g2_a21oi_1 _32396_ (.A1(_20960_),
    .A2(_22061_),
    .Y(_02085_),
    .B1(_20965_));
 sg13g2_nor3_1 _32397_ (.A(net7177),
    .B(_02084_),
    .C(_02085_),
    .Y(_02086_));
 sg13g2_o21ai_1 _32398_ (.B1(net6194),
    .Y(_02087_),
    .A1(\u_inv.f_next[233] ),
    .A2(net7305));
 sg13g2_o21ai_1 _32399_ (.B1(_02083_),
    .Y(_02088_),
    .A1(_02086_),
    .A2(_02087_));
 sg13g2_o21ai_1 _32400_ (.B1(_21065_),
    .Y(_02089_),
    .A1(_19862_),
    .A2(_02064_));
 sg13g2_or3_1 _32401_ (.A(_19862_),
    .B(_21065_),
    .C(_02064_),
    .X(_02090_));
 sg13g2_and3_1 _32402_ (.X(_02091_),
    .A(net7311),
    .B(_02089_),
    .C(_02090_));
 sg13g2_o21ai_1 _32403_ (.B1(net6202),
    .Y(_02092_),
    .A1(\u_inv.f_next[249] ),
    .A2(net7311));
 sg13g2_nor2_1 _32404_ (.A(_21065_),
    .B(_21083_),
    .Y(_02093_));
 sg13g2_o21ai_1 _32405_ (.B1(_02093_),
    .Y(_02094_),
    .A1(_21063_),
    .A2(_21786_));
 sg13g2_nor2_1 _32406_ (.A(net6202),
    .B(_21838_),
    .Y(_02095_));
 sg13g2_nand3_1 _32407_ (.B(_02094_),
    .C(_02095_),
    .A(_21084_),
    .Y(_02096_));
 sg13g2_o21ai_1 _32408_ (.B1(_02096_),
    .Y(_02097_),
    .A1(_02091_),
    .A2(_02092_));
 sg13g2_a21oi_1 _32409_ (.A1(_21059_),
    .A2(_21799_),
    .Y(_02098_),
    .B1(_21032_));
 sg13g2_nand3_1 _32410_ (.B(_21059_),
    .C(_21799_),
    .A(_21032_),
    .Y(_02099_));
 sg13g2_nand2b_1 _32411_ (.Y(_02100_),
    .B(_02099_),
    .A_N(_02098_));
 sg13g2_o21ai_1 _32412_ (.B1(net6201),
    .Y(_02101_),
    .A1(\u_inv.f_next[244] ),
    .A2(net7311));
 sg13g2_a21oi_1 _32413_ (.A1(net7310),
    .A2(_02100_),
    .Y(_02102_),
    .B1(_02101_));
 sg13g2_nand3_1 _32414_ (.B(_21775_),
    .C(_21806_),
    .A(_21031_),
    .Y(_02103_));
 sg13g2_nor2_1 _32415_ (.A(net6200),
    .B(_21807_),
    .Y(_02104_));
 sg13g2_a21o_2 _32416_ (.A2(_02104_),
    .A1(_02103_),
    .B1(_02102_),
    .X(_02105_));
 sg13g2_a21oi_1 _32417_ (.A1(\u_inv.f_next[194] ),
    .A2(\u_inv.f_reg[194] ),
    .Y(_02106_),
    .B1(_23535_));
 sg13g2_xnor2_1 _32418_ (.Y(_02107_),
    .A(_19990_),
    .B(_02106_));
 sg13g2_nand2_1 _32419_ (.Y(_02108_),
    .A(net7307),
    .B(_02107_));
 sg13g2_a21oi_1 _32420_ (.A1(_17995_),
    .A2(net7180),
    .Y(_02109_),
    .B1(net6278));
 sg13g2_nand2_1 _32421_ (.Y(_02110_),
    .A(_21652_),
    .B(_23542_));
 sg13g2_or2_1 _32422_ (.X(_02111_),
    .B(_02110_),
    .A(_19990_));
 sg13g2_a21oi_1 _32423_ (.A1(_19990_),
    .A2(_02110_),
    .Y(_02112_),
    .B1(net6197));
 sg13g2_and2_1 _32424_ (.A(_02111_),
    .B(_02112_),
    .X(_02113_));
 sg13g2_a22oi_1 _32425_ (.Y(_02114_),
    .B1(_02111_),
    .B2(_02112_),
    .A2(_02109_),
    .A1(_02108_));
 sg13g2_a21o_1 _32426_ (.A2(_02109_),
    .A1(_02108_),
    .B1(_02113_),
    .X(_02115_));
 sg13g2_o21ai_1 _32427_ (.B1(_20030_),
    .Y(_02116_),
    .A1(_20081_),
    .A2(_21975_));
 sg13g2_a21oi_1 _32428_ (.A1(_20073_),
    .A2(_02116_),
    .Y(_02117_),
    .B1(_20022_));
 sg13g2_and3_1 _32429_ (.X(_02118_),
    .A(_20022_),
    .B(_20073_),
    .C(_02116_));
 sg13g2_o21ai_1 _32430_ (.B1(net7314),
    .Y(_02119_),
    .A1(_02117_),
    .A2(_02118_));
 sg13g2_a21oi_1 _32431_ (.A1(_17999_),
    .A2(net7184),
    .Y(_02120_),
    .B1(net6284));
 sg13g2_nand2_1 _32432_ (.Y(_02121_),
    .A(_02119_),
    .B(_02120_));
 sg13g2_a21oi_2 _32433_ (.B1(_20021_),
    .Y(_02122_),
    .A2(_21986_),
    .A1(_21605_));
 sg13g2_nand3_1 _32434_ (.B(_21605_),
    .C(_21986_),
    .A(_20021_),
    .Y(_02123_));
 sg13g2_nand2_1 _32435_ (.Y(_02124_),
    .A(net6284),
    .B(_02123_));
 sg13g2_nor2_1 _32436_ (.A(net6205),
    .B(_02122_),
    .Y(_02125_));
 sg13g2_a22oi_1 _32437_ (.Y(_02126_),
    .B1(_02123_),
    .B2(_02125_),
    .A2(_02120_),
    .A1(_02119_));
 sg13g2_o21ai_1 _32438_ (.B1(_02121_),
    .Y(_02127_),
    .A1(_02122_),
    .A2(_02124_));
 sg13g2_o21ai_1 _32439_ (.B1(_19987_),
    .Y(_02128_),
    .A1(_19997_),
    .A2(_22116_));
 sg13g2_a21oi_1 _32440_ (.A1(_20003_),
    .A2(_02128_),
    .Y(_02129_),
    .B1(_19981_));
 sg13g2_and3_1 _32441_ (.X(_02130_),
    .A(_19981_),
    .B(_20003_),
    .C(_02128_));
 sg13g2_o21ai_1 _32442_ (.B1(net7307),
    .Y(_02131_),
    .A1(_02129_),
    .A2(_02130_));
 sg13g2_a21oi_1 _32443_ (.A1(_17992_),
    .A2(net7180),
    .Y(_02132_),
    .B1(net6278));
 sg13g2_nand2_1 _32444_ (.Y(_02133_),
    .A(_02131_),
    .B(_02132_));
 sg13g2_a21oi_2 _32445_ (.B1(_19982_),
    .Y(_02134_),
    .A2(_22126_),
    .A1(_21649_));
 sg13g2_nand3_1 _32446_ (.B(_21649_),
    .C(_22126_),
    .A(_19982_),
    .Y(_02135_));
 sg13g2_nand2_1 _32447_ (.Y(_02136_),
    .A(net6278),
    .B(_02135_));
 sg13g2_nor2_1 _32448_ (.A(net6197),
    .B(_02134_),
    .Y(_02137_));
 sg13g2_a22oi_1 _32449_ (.Y(_02138_),
    .B1(_02135_),
    .B2(_02137_),
    .A2(_02132_),
    .A1(_02131_));
 sg13g2_o21ai_1 _32450_ (.B1(_02133_),
    .Y(_02139_),
    .A1(_02134_),
    .A2(_02136_));
 sg13g2_nand3_1 _32451_ (.B(_21685_),
    .C(_21824_),
    .A(_19901_),
    .Y(_02140_));
 sg13g2_nor2_1 _32452_ (.A(net6193),
    .B(_21825_),
    .Y(_02141_));
 sg13g2_or3_1 _32453_ (.A(_19889_),
    .B(_19902_),
    .C(_21989_),
    .X(_02142_));
 sg13g2_o21ai_1 _32454_ (.B1(_19902_),
    .Y(_02143_),
    .A1(_19889_),
    .A2(_21989_));
 sg13g2_nand3_1 _32455_ (.B(_02142_),
    .C(_02143_),
    .A(net7303),
    .Y(_02144_));
 sg13g2_a21oi_1 _32456_ (.A1(_17980_),
    .A2(net7179),
    .Y(_02145_),
    .B1(net6275));
 sg13g2_a22oi_1 _32457_ (.Y(_02146_),
    .B1(_02144_),
    .B2(_02145_),
    .A2(_02141_),
    .A1(_02140_));
 sg13g2_a21oi_1 _32458_ (.A1(_21690_),
    .A2(_01966_),
    .Y(_02147_),
    .B1(_19879_));
 sg13g2_nor3_1 _32459_ (.A(_19877_),
    .B(_21691_),
    .C(_02147_),
    .Y(_02148_));
 sg13g2_or4_1 _32460_ (.A(net6195),
    .B(_21692_),
    .C(_01967_),
    .D(_02148_),
    .X(_02149_));
 sg13g2_a21oi_1 _32461_ (.A1(_19894_),
    .A2(_01959_),
    .Y(_02150_),
    .B1(_19880_));
 sg13g2_or3_1 _32462_ (.A(_19877_),
    .B(_19878_),
    .C(_02150_),
    .X(_02151_));
 sg13g2_o21ai_1 _32463_ (.B1(_19877_),
    .Y(_02152_),
    .A1(_19878_),
    .A2(_02150_));
 sg13g2_and3_1 _32464_ (.X(_02153_),
    .A(net7304),
    .B(_02151_),
    .C(_02152_));
 sg13g2_o21ai_1 _32465_ (.B1(net6195),
    .Y(_02154_),
    .A1(\u_inv.f_next[221] ),
    .A2(net7304));
 sg13g2_o21ai_1 _32466_ (.B1(_02149_),
    .Y(_02155_),
    .A1(_02153_),
    .A2(_02154_));
 sg13g2_nand3_1 _32467_ (.B(_19894_),
    .C(_01959_),
    .A(_19880_),
    .Y(_02156_));
 sg13g2_nand2_1 _32468_ (.Y(_02157_),
    .A(\u_inv.f_next[220] ),
    .B(net7177));
 sg13g2_nand3b_1 _32469_ (.B(_02156_),
    .C(net7305),
    .Y(_02158_),
    .A_N(_02150_));
 sg13g2_a21oi_1 _32470_ (.A1(_02157_),
    .A2(_02158_),
    .Y(_02159_),
    .B1(net6276));
 sg13g2_nand3_1 _32471_ (.B(_21690_),
    .C(_01966_),
    .A(_19879_),
    .Y(_02160_));
 sg13g2_nor2_1 _32472_ (.A(net6195),
    .B(_02147_),
    .Y(_02161_));
 sg13g2_a21o_2 _32473_ (.A2(_02161_),
    .A1(_02160_),
    .B1(_02159_),
    .X(_02162_));
 sg13g2_nand2b_1 _32474_ (.Y(_02163_),
    .B(_22034_),
    .A_N(_21670_));
 sg13g2_xnor2_1 _32475_ (.Y(_02164_),
    .A(_19961_),
    .B(_02163_));
 sg13g2_nor3_1 _32476_ (.A(_19962_),
    .B(_19970_),
    .C(_21923_),
    .Y(_02165_));
 sg13g2_o21ai_1 _32477_ (.B1(_19962_),
    .Y(_02166_),
    .A1(_19970_),
    .A2(_21923_));
 sg13g2_nor2_1 _32478_ (.A(net7195),
    .B(_02165_),
    .Y(_02167_));
 sg13g2_a221oi_1 _32479_ (.B2(_02167_),
    .C1(net6278),
    .B1(_02166_),
    .A1(\u_inv.f_next[202] ),
    .Y(_02168_),
    .A2(net7180));
 sg13g2_a21o_2 _32480_ (.A2(_02164_),
    .A1(net6282),
    .B1(_02168_),
    .X(_02169_));
 sg13g2_a21oi_1 _32481_ (.A1(_20102_),
    .A2(_22051_),
    .Y(_02170_),
    .B1(_20099_));
 sg13g2_a21oi_1 _32482_ (.A1(_20105_),
    .A2(_02170_),
    .Y(_02171_),
    .B1(net7196));
 sg13g2_o21ai_1 _32483_ (.B1(_02171_),
    .Y(_02172_),
    .A1(_20105_),
    .A2(_02170_));
 sg13g2_a21oi_1 _32484_ (.A1(_18013_),
    .A2(net7196),
    .Y(_02173_),
    .B1(net6300));
 sg13g2_nor3_1 _32485_ (.A(_20104_),
    .B(_21555_),
    .C(_23570_),
    .Y(_02174_));
 sg13g2_o21ai_1 _32486_ (.B1(_20104_),
    .Y(_02175_),
    .A1(_21555_),
    .A2(_23570_));
 sg13g2_nor2_1 _32487_ (.A(net6213),
    .B(_02174_),
    .Y(_02176_));
 sg13g2_a22oi_1 _32488_ (.Y(_02177_),
    .B1(_02175_),
    .B2(_02176_),
    .A2(_02173_),
    .A1(_02172_));
 sg13g2_nand3_1 _32489_ (.B(_21614_),
    .C(_23551_),
    .A(_20041_),
    .Y(_02178_));
 sg13g2_a21oi_1 _32490_ (.A1(_21614_),
    .A2(_23551_),
    .Y(_02179_),
    .B1(_20041_));
 sg13g2_nor2_1 _32491_ (.A(net6205),
    .B(_02179_),
    .Y(_02180_));
 sg13g2_a21oi_1 _32492_ (.A1(_20038_),
    .A2(_23545_),
    .Y(_02181_),
    .B1(_20037_));
 sg13g2_or2_1 _32493_ (.X(_02182_),
    .B(_02181_),
    .A(_20041_));
 sg13g2_a21oi_1 _32494_ (.A1(_20041_),
    .A2(_02181_),
    .Y(_02183_),
    .B1(net7186));
 sg13g2_nand2_1 _32495_ (.Y(_02184_),
    .A(_18001_),
    .B(net7184));
 sg13g2_a21oi_1 _32496_ (.A1(_02182_),
    .A2(_02183_),
    .Y(_02185_),
    .B1(net6283));
 sg13g2_a22oi_1 _32497_ (.Y(_02186_),
    .B1(_02184_),
    .B2(_02185_),
    .A2(_02180_),
    .A1(_02178_));
 sg13g2_and3_1 _32498_ (.X(_02187_),
    .A(_19910_),
    .B(_19933_),
    .C(_01988_));
 sg13g2_o21ai_1 _32499_ (.B1(net7301),
    .Y(_02188_),
    .A1(_01989_),
    .A2(_02187_));
 sg13g2_o21ai_1 _32500_ (.B1(_02188_),
    .Y(_02189_),
    .A1(\u_inv.f_next[214] ),
    .A2(net7301));
 sg13g2_nand3_1 _32501_ (.B(_21709_),
    .C(_22147_),
    .A(_19909_),
    .Y(_02190_));
 sg13g2_nand3b_1 _32502_ (.B(_02190_),
    .C(net6274),
    .Y(_02191_),
    .A_N(_01994_));
 sg13g2_o21ai_1 _32503_ (.B1(_02191_),
    .Y(_02192_),
    .A1(net6274),
    .A2(_02189_));
 sg13g2_xnor2_1 _32504_ (.Y(_02193_),
    .A(_19921_),
    .B(_22129_));
 sg13g2_mux2_1 _32505_ (.A0(\u_inv.f_next[210] ),
    .A1(_02193_),
    .S(net7302),
    .X(_02194_));
 sg13g2_nand3_1 _32506_ (.B(_21702_),
    .C(_22017_),
    .A(_19921_),
    .Y(_02195_));
 sg13g2_nor2_1 _32507_ (.A(net6192),
    .B(_01978_),
    .Y(_02196_));
 sg13g2_and2_1 _32508_ (.A(_02195_),
    .B(_02196_),
    .X(_02197_));
 sg13g2_a22oi_1 _32509_ (.Y(_02198_),
    .B1(_02195_),
    .B2(_02196_),
    .A2(_02194_),
    .A1(net6193));
 sg13g2_a21o_1 _32510_ (.A2(_02194_),
    .A1(net6193),
    .B1(_02197_),
    .X(_02199_));
 sg13g2_o21ai_1 _32511_ (.B1(_21028_),
    .Y(_02200_),
    .A1(_21030_),
    .A2(_02098_));
 sg13g2_nor3_1 _32512_ (.A(_21028_),
    .B(_21030_),
    .C(_02098_),
    .Y(_02201_));
 sg13g2_nand3b_1 _32513_ (.B(net7311),
    .C(_02200_),
    .Y(_02202_),
    .A_N(_02201_));
 sg13g2_o21ai_1 _32514_ (.B1(net6201),
    .Y(_02203_),
    .A1(\u_inv.f_next[245] ),
    .A2(net7311));
 sg13g2_inv_1 _32515_ (.Y(_02204_),
    .A(_02203_));
 sg13g2_nor3_1 _32516_ (.A(_21028_),
    .B(_21779_),
    .C(_21807_),
    .Y(_02205_));
 sg13g2_nor2_1 _32517_ (.A(net6201),
    .B(_02205_),
    .Y(_02206_));
 sg13g2_a22oi_1 _32518_ (.Y(_02207_),
    .B1(_02206_),
    .B2(_21808_),
    .A2(_02204_),
    .A1(_02202_));
 sg13g2_inv_1 _32519_ (.Y(_02208_),
    .A(_02207_));
 sg13g2_nor3_1 _32520_ (.A(_19979_),
    .B(_21662_),
    .C(_02134_),
    .Y(_02209_));
 sg13g2_o21ai_1 _32521_ (.B1(_19979_),
    .Y(_02210_),
    .A1(_21662_),
    .A2(_02134_));
 sg13g2_nor2_1 _32522_ (.A(net6197),
    .B(_02209_),
    .Y(_02211_));
 sg13g2_nor2_1 _32523_ (.A(_19980_),
    .B(_02129_),
    .Y(_02212_));
 sg13g2_xnor2_1 _32524_ (.Y(_02213_),
    .A(_19979_),
    .B(_02212_));
 sg13g2_o21ai_1 _32525_ (.B1(net6197),
    .Y(_02214_),
    .A1(\u_inv.f_next[199] ),
    .A2(net7307));
 sg13g2_a21oi_1 _32526_ (.A1(net7307),
    .A2(_02213_),
    .Y(_02215_),
    .B1(_02214_));
 sg13g2_a21o_2 _32527_ (.A2(_02211_),
    .A1(_02210_),
    .B1(_02215_),
    .X(_02216_));
 sg13g2_or3_1 _32528_ (.A(_19873_),
    .B(_19896_),
    .C(_01960_),
    .X(_02217_));
 sg13g2_a21oi_1 _32529_ (.A1(_01961_),
    .A2(_02217_),
    .Y(_02218_),
    .B1(net7177));
 sg13g2_o21ai_1 _32530_ (.B1(net6195),
    .Y(_02219_),
    .A1(\u_inv.f_next[222] ),
    .A2(net7304));
 sg13g2_nor3_1 _32531_ (.A(_19874_),
    .B(_21694_),
    .C(_01967_),
    .Y(_02220_));
 sg13g2_nand3b_1 _32532_ (.B(net6276),
    .C(_01968_),
    .Y(_02221_),
    .A_N(_02220_));
 sg13g2_o21ai_1 _32533_ (.B1(_02221_),
    .Y(_02222_),
    .A1(_02218_),
    .A2(_02219_));
 sg13g2_or3_1 _32534_ (.A(_19854_),
    .B(_19869_),
    .C(_21068_),
    .X(_02223_));
 sg13g2_a21oi_1 _32535_ (.A1(_02045_),
    .A2(_02223_),
    .Y(_02224_),
    .B1(net7183));
 sg13g2_o21ai_1 _32536_ (.B1(net6203),
    .Y(_02225_),
    .A1(\u_inv.f_next[252] ),
    .A2(net7312));
 sg13g2_nor2_1 _32537_ (.A(_02224_),
    .B(_02225_),
    .Y(_02226_));
 sg13g2_nor3_1 _32538_ (.A(_19855_),
    .B(_21088_),
    .C(_21791_),
    .Y(_02227_));
 sg13g2_nor3_1 _32539_ (.A(net6203),
    .B(_02051_),
    .C(_02227_),
    .Y(_02228_));
 sg13g2_nor2_1 _32540_ (.A(_02226_),
    .B(_02228_),
    .Y(_02229_));
 sg13g2_o21ai_1 _32541_ (.B1(_20018_),
    .Y(_02230_),
    .A1(_21607_),
    .A2(_02122_));
 sg13g2_nor3_1 _32542_ (.A(_20018_),
    .B(_21607_),
    .C(_02122_),
    .Y(_02231_));
 sg13g2_nand3b_1 _32543_ (.B(net6284),
    .C(_02230_),
    .Y(_02232_),
    .A_N(_02231_));
 sg13g2_o21ai_1 _32544_ (.B1(_20018_),
    .Y(_02233_),
    .A1(_20019_),
    .A2(_02117_));
 sg13g2_nand3b_1 _32545_ (.B(_20017_),
    .C(_20020_),
    .Y(_02234_),
    .A_N(_02117_));
 sg13g2_and3_1 _32546_ (.X(_02235_),
    .A(net7314),
    .B(_02233_),
    .C(_02234_));
 sg13g2_o21ai_1 _32547_ (.B1(net6205),
    .Y(_02236_),
    .A1(\u_inv.f_next[191] ),
    .A2(net7315));
 sg13g2_o21ai_1 _32548_ (.B1(_02232_),
    .Y(_02237_),
    .A1(_02235_),
    .A2(_02236_));
 sg13g2_nand3_1 _32549_ (.B(_19865_),
    .C(_21832_),
    .A(_19860_),
    .Y(_02238_));
 sg13g2_a21oi_1 _32550_ (.A1(_21833_),
    .A2(_02238_),
    .Y(_02239_),
    .B1(net7181));
 sg13g2_o21ai_1 _32551_ (.B1(net6201),
    .Y(_02240_),
    .A1(\u_inv.f_next[250] ),
    .A2(net7312));
 sg13g2_nor2_1 _32552_ (.A(_02239_),
    .B(_02240_),
    .Y(_02241_));
 sg13g2_or3_1 _32553_ (.A(_19860_),
    .B(_21085_),
    .C(_21838_),
    .X(_02242_));
 sg13g2_nand3_1 _32554_ (.B(_21839_),
    .C(_02242_),
    .A(net6280),
    .Y(_02243_));
 sg13g2_nor2b_2 _32555_ (.A(_02241_),
    .B_N(_02243_),
    .Y(_02244_));
 sg13g2_o21ai_1 _32556_ (.B1(_02243_),
    .Y(_02245_),
    .A1(_02239_),
    .A2(_02240_));
 sg13g2_a21oi_1 _32557_ (.A1(_20941_),
    .A2(_02033_),
    .Y(_02246_),
    .B1(_21738_));
 sg13g2_a21oi_1 _32558_ (.A1(_20943_),
    .A2(_02246_),
    .Y(_02247_),
    .B1(net6194));
 sg13g2_o21ai_1 _32559_ (.B1(_02247_),
    .Y(_02248_),
    .A1(_20943_),
    .A2(_02246_));
 sg13g2_o21ai_1 _32560_ (.B1(_20944_),
    .Y(_02249_),
    .A1(_20939_),
    .A2(_02028_));
 sg13g2_nor3_1 _32561_ (.A(_20939_),
    .B(_20944_),
    .C(_02028_),
    .Y(_02250_));
 sg13g2_nand2_1 _32562_ (.Y(_02251_),
    .A(net7306),
    .B(_02249_));
 sg13g2_nor2_1 _32563_ (.A(\u_inv.f_next[231] ),
    .B(net7305),
    .Y(_02252_));
 sg13g2_o21ai_1 _32564_ (.B1(net6194),
    .Y(_02253_),
    .A1(_02250_),
    .A2(_02251_));
 sg13g2_o21ai_1 _32565_ (.B1(_02248_),
    .Y(_02254_),
    .A1(_02252_),
    .A2(_02253_));
 sg13g2_nand3_1 _32566_ (.B(_19964_),
    .C(_02166_),
    .A(_19960_),
    .Y(_02255_));
 sg13g2_a21oi_1 _32567_ (.A1(_19960_),
    .A2(_02166_),
    .Y(_02256_),
    .B1(_19964_));
 sg13g2_nand2_1 _32568_ (.Y(_02257_),
    .A(net7308),
    .B(_02255_));
 sg13g2_a21oi_1 _32569_ (.A1(_17989_),
    .A2(net7180),
    .Y(_02258_),
    .B1(net6282));
 sg13g2_o21ai_1 _32570_ (.B1(_02258_),
    .Y(_02259_),
    .A1(_02256_),
    .A2(_02257_));
 sg13g2_a21oi_1 _32571_ (.A1(_19961_),
    .A2(_02163_),
    .Y(_02260_),
    .B1(_21668_));
 sg13g2_xnor2_1 _32572_ (.Y(_02261_),
    .A(_19964_),
    .B(_02260_));
 sg13g2_o21ai_1 _32573_ (.B1(_02259_),
    .Y(_02262_),
    .A1(net6198),
    .A2(_02261_));
 sg13g2_nand4_1 _32574_ (.B(_02080_),
    .C(_02126_),
    .A(_21952_),
    .Y(_02263_),
    .D(_02198_));
 sg13g2_nand3b_1 _32575_ (.B(_02070_),
    .C(_02068_),
    .Y(_02264_),
    .A_N(_02088_));
 sg13g2_or4_1 _32576_ (.A(_21940_),
    .B(_02105_),
    .C(_02263_),
    .D(_02264_),
    .X(_02265_));
 sg13g2_nand2_1 _32577_ (.Y(_02266_),
    .A(_23512_),
    .B(_01903_));
 sg13g2_or2_1 _32578_ (.X(_02267_),
    .B(_01944_),
    .A(_01925_));
 sg13g2_nor4_2 _32579_ (.A(_22216_),
    .B(_22236_),
    .C(_22263_),
    .Y(_02268_),
    .D(_22282_));
 sg13g2_nand2b_2 _32580_ (.Y(_02269_),
    .B(_22427_),
    .A_N(_22272_));
 sg13g2_nor3_2 _32581_ (.A(_22222_),
    .B(_22402_),
    .C(_02269_),
    .Y(_02270_));
 sg13g2_nand4_1 _32582_ (.B(_23352_),
    .C(_02268_),
    .A(_23273_),
    .Y(_02271_),
    .D(_02270_));
 sg13g2_or4_1 _32583_ (.A(_22202_),
    .B(_23389_),
    .C(_23457_),
    .D(_02271_),
    .X(_02272_));
 sg13g2_nor4_1 _32584_ (.A(_22328_),
    .B(_22349_),
    .C(_22378_),
    .D(_22394_),
    .Y(_02273_));
 sg13g2_nor3_1 _32585_ (.A(_22373_),
    .B(_22409_),
    .C(_23205_),
    .Y(_02274_));
 sg13g2_nor3_1 _32586_ (.A(_22471_),
    .B(_22493_),
    .C(_23182_),
    .Y(_02275_));
 sg13g2_nand4_1 _32587_ (.B(_23169_),
    .C(_23199_),
    .A(_22449_),
    .Y(_02276_),
    .D(_02275_));
 sg13g2_nor3_1 _32588_ (.A(_23175_),
    .B(_23188_),
    .C(_23193_),
    .Y(_02277_));
 sg13g2_nand4_1 _32589_ (.B(_22484_),
    .C(_23158_),
    .A(_22461_),
    .Y(_02278_),
    .D(_02277_));
 sg13g2_nor4_1 _32590_ (.A(_22436_),
    .B(_22478_),
    .C(_02276_),
    .D(_02278_),
    .Y(_02279_));
 sg13g2_nor2_1 _32591_ (.A(_22354_),
    .B(_22443_),
    .Y(_02280_));
 sg13g2_nand4_1 _32592_ (.B(_02274_),
    .C(_02279_),
    .A(_22336_),
    .Y(_02281_),
    .D(_02280_));
 sg13g2_nor4_1 _32593_ (.A(_22341_),
    .B(_22367_),
    .C(_22388_),
    .D(_02281_),
    .Y(_02282_));
 sg13g2_and3_2 _32594_ (.X(_02283_),
    .A(_22253_),
    .B(_02273_),
    .C(_02282_));
 sg13g2_nor2b_1 _32595_ (.A(_23279_),
    .B_N(_23362_),
    .Y(_02284_));
 sg13g2_nand4_1 _32596_ (.B(_22194_),
    .C(_02283_),
    .A(_22176_),
    .Y(_02285_),
    .D(_02284_));
 sg13g2_or4_1 _32597_ (.A(_23320_),
    .B(_23328_),
    .C(_23370_),
    .D(_23381_),
    .X(_02286_));
 sg13g2_nor3_2 _32598_ (.A(_22297_),
    .B(_23251_),
    .C(_23267_),
    .Y(_02287_));
 sg13g2_nor4_1 _32599_ (.A(_22322_),
    .B(_23226_),
    .C(_23243_),
    .D(_23259_),
    .Y(_02288_));
 sg13g2_nor4_1 _32600_ (.A(_23212_),
    .B(_23220_),
    .C(_23234_),
    .D(_23334_),
    .Y(_02289_));
 sg13g2_nand4_1 _32601_ (.B(_02287_),
    .C(_02288_),
    .A(_22303_),
    .Y(_02290_),
    .D(_02289_));
 sg13g2_nand4_1 _32602_ (.B(_23343_),
    .C(_23397_),
    .A(_23286_),
    .Y(_02291_),
    .D(_23410_));
 sg13g2_nor2_1 _32603_ (.A(_23292_),
    .B(_23312_),
    .Y(_02292_));
 sg13g2_nand3b_1 _32604_ (.B(_23465_),
    .C(_02292_),
    .Y(_02293_),
    .A_N(_23303_));
 sg13g2_or4_1 _32605_ (.A(_02286_),
    .B(_02290_),
    .C(_02291_),
    .D(_02293_),
    .X(_02294_));
 sg13g2_nand4_1 _32606_ (.B(_23436_),
    .C(_23620_),
    .A(_23417_),
    .Y(_02295_),
    .D(_23627_));
 sg13g2_or4_1 _32607_ (.A(_02272_),
    .B(_02285_),
    .C(_02294_),
    .D(_02295_),
    .X(_02296_));
 sg13g2_nand4_1 _32608_ (.B(_23480_),
    .C(_23488_),
    .A(_23474_),
    .Y(_02297_),
    .D(_23614_));
 sg13g2_nand2_1 _32609_ (.Y(_02298_),
    .A(_23428_),
    .B(_23495_));
 sg13g2_or4_1 _32610_ (.A(_23449_),
    .B(_23503_),
    .C(_02297_),
    .D(_02298_),
    .X(_02299_));
 sg13g2_or4_1 _32611_ (.A(_01937_),
    .B(_02267_),
    .C(_02296_),
    .D(_02299_),
    .X(_02300_));
 sg13g2_or4_1 _32612_ (.A(_21960_),
    .B(_23519_),
    .C(_02266_),
    .D(_02300_),
    .X(_02301_));
 sg13g2_nand4_1 _32613_ (.B(_22068_),
    .C(_22082_),
    .A(_22026_),
    .Y(_02302_),
    .D(_22113_));
 sg13g2_nor3_2 _32614_ (.A(_23645_),
    .B(_01912_),
    .C(_01919_),
    .Y(_02303_));
 sg13g2_nand2_1 _32615_ (.Y(_02304_),
    .A(_22141_),
    .B(_02303_));
 sg13g2_or4_1 _32616_ (.A(_22019_),
    .B(_23564_),
    .C(_02302_),
    .D(_02304_),
    .X(_02305_));
 sg13g2_nand3_1 _32617_ (.B(_23534_),
    .C(_02146_),
    .A(_22128_),
    .Y(_02306_));
 sg13g2_nor4_2 _32618_ (.A(_02265_),
    .B(_02301_),
    .C(_02305_),
    .Y(_02307_),
    .D(_02306_));
 sg13g2_or2_1 _32619_ (.X(_02308_),
    .B(_02222_),
    .A(_02018_));
 sg13g2_nor4_1 _32620_ (.A(_21907_),
    .B(_02054_),
    .C(_02216_),
    .D(_02308_),
    .Y(_02309_));
 sg13g2_nand4_1 _32621_ (.B(_02114_),
    .C(_02138_),
    .A(_22150_),
    .Y(_02310_),
    .D(_02177_));
 sg13g2_nand2_2 _32622_ (.Y(_02311_),
    .A(_02169_),
    .B(_02186_));
 sg13g2_or4_1 _32623_ (.A(_02097_),
    .B(_02155_),
    .C(_02310_),
    .D(_02311_),
    .X(_02312_));
 sg13g2_nand2_1 _32624_ (.Y(_02313_),
    .A(_22059_),
    .B(_22093_));
 sg13g2_nor4_2 _32625_ (.A(_23601_),
    .B(_23609_),
    .C(_23633_),
    .Y(_02314_),
    .D(_23639_));
 sg13g2_nor4_1 _32626_ (.A(_23580_),
    .B(_23587_),
    .C(_23594_),
    .D(_01931_),
    .Y(_02315_));
 sg13g2_nand3b_1 _32627_ (.B(_02314_),
    .C(_02315_),
    .Y(_02316_),
    .A_N(_23527_));
 sg13g2_or4_1 _32628_ (.A(_22101_),
    .B(_02036_),
    .C(_02313_),
    .D(_02316_),
    .X(_02317_));
 sg13g2_and4_1 _32629_ (.A(_21971_),
    .B(_21997_),
    .C(_22032_),
    .D(_22035_),
    .X(_02318_));
 sg13g2_nor2_2 _32630_ (.A(_22009_),
    .B(_23544_),
    .Y(_02319_));
 sg13g2_nor2b_2 _32631_ (.A(_23554_),
    .B_N(_23573_),
    .Y(_02320_));
 sg13g2_nand4_1 _32632_ (.B(_02318_),
    .C(_02319_),
    .A(_22158_),
    .Y(_02321_),
    .D(_02320_));
 sg13g2_or4_1 _32633_ (.A(_21988_),
    .B(_02162_),
    .C(_02192_),
    .D(_02321_),
    .X(_02322_));
 sg13g2_nand4_1 _32634_ (.B(_01953_),
    .C(_01957_),
    .A(_21911_),
    .Y(_02323_),
    .D(_02207_));
 sg13g2_nor4_1 _32635_ (.A(_02312_),
    .B(_02317_),
    .C(_02322_),
    .D(_02323_),
    .Y(_02324_));
 sg13g2_or2_1 _32636_ (.X(_02325_),
    .B(_02044_),
    .A(_02026_));
 sg13g2_nand3_1 _32637_ (.B(_01950_),
    .C(_02062_),
    .A(_21932_),
    .Y(_02326_));
 sg13g2_nor4_1 _32638_ (.A(_21881_),
    .B(_02254_),
    .C(_02325_),
    .D(_02326_),
    .Y(_02327_));
 sg13g2_and4_1 _32639_ (.A(_02307_),
    .B(_02309_),
    .C(_02324_),
    .D(_02327_),
    .X(_02328_));
 sg13g2_and4_1 _32640_ (.A(_21843_),
    .B(_21862_),
    .C(_01972_),
    .D(_02011_),
    .X(_02329_));
 sg13g2_nor4_2 _32641_ (.A(_01981_),
    .B(_02237_),
    .C(_02245_),
    .Y(_02330_),
    .D(_02262_));
 sg13g2_nor4_1 _32642_ (.A(_01987_),
    .B(_01998_),
    .C(_02226_),
    .D(_02228_),
    .Y(_02331_));
 sg13g2_and4_1 _32643_ (.A(_21830_),
    .B(_02005_),
    .C(_02330_),
    .D(_02331_),
    .X(_02332_));
 sg13g2_and4_1 _32644_ (.A(_21797_),
    .B(_21812_),
    .C(_02329_),
    .D(_02332_),
    .X(_02333_));
 sg13g2_nand2_2 _32645_ (.Y(_02334_),
    .A(net5319),
    .B(net5315));
 sg13g2_nand2_2 _32646_ (.Y(_02335_),
    .A(\u_inv.counter[9] ),
    .B(\u_inv.counter[8] ));
 sg13g2_nand2_2 _32647_ (.Y(_02336_),
    .A(_22954_),
    .B(_02335_));
 sg13g2_nand4_1 _32648_ (.B(\u_inv.counter[7] ),
    .C(net7248),
    .A(\u_inv.counter[9] ),
    .Y(_02337_),
    .D(\u_inv.counter[5] ));
 sg13g2_o21ai_1 _32649_ (.B1(\u_inv.counter[2] ),
    .Y(_02338_),
    .A1(\u_inv.counter[1] ),
    .A2(net7250));
 sg13g2_nor2_1 _32650_ (.A(\u_inv.counter[4] ),
    .B(\u_inv.counter[3] ),
    .Y(_02339_));
 sg13g2_a21oi_2 _32651_ (.B1(_02337_),
    .Y(_02340_),
    .A2(_02339_),
    .A1(_02338_));
 sg13g2_nor2_2 _32652_ (.A(_02336_),
    .B(_02340_),
    .Y(_02341_));
 sg13g2_or2_1 _32653_ (.X(_02342_),
    .B(_02340_),
    .A(_02336_));
 sg13g2_a21oi_2 _32654_ (.B1(net5990),
    .Y(_02343_),
    .A2(net5317),
    .A1(net5321));
 sg13g2_nand2_2 _32655_ (.Y(_02344_),
    .A(net5277),
    .B(net6008));
 sg13g2_a21oi_2 _32656_ (.B1(net7023),
    .Y(_02345_),
    .A2(net5315),
    .A1(net5319));
 sg13g2_nor2_2 _32657_ (.A(net7019),
    .B(net5155),
    .Y(_02346_));
 sg13g2_and2_1 _32658_ (.A(net7493),
    .B(net7110),
    .X(_02347_));
 sg13g2_nand2_1 _32659_ (.Y(_02348_),
    .A(net7501),
    .B(net7115));
 sg13g2_nor2_1 _32660_ (.A(net1306),
    .B(net6389),
    .Y(_02349_));
 sg13g2_a22oi_1 _32661_ (.Y(_02350_),
    .B1(_02349_),
    .B2(net7019),
    .A2(net6866),
    .A1(_22954_));
 sg13g2_nor3_1 _32662_ (.A(\u_inv.counter[4] ),
    .B(\u_inv.counter[3] ),
    .C(\u_inv.counter[2] ),
    .Y(_02351_));
 sg13g2_nor2_2 _32663_ (.A(_02337_),
    .B(_02351_),
    .Y(_02352_));
 sg13g2_nor2_2 _32664_ (.A(_02336_),
    .B(_02352_),
    .Y(_02353_));
 sg13g2_nor3_1 _32665_ (.A(_19842_),
    .B(_02336_),
    .C(_02352_),
    .Y(_02354_));
 sg13g2_nand2_2 _32666_ (.Y(_02355_),
    .A(_19841_),
    .B(_02353_));
 sg13g2_a21oi_1 _32667_ (.A1(net5319),
    .A2(net5315),
    .Y(_02356_),
    .B1(net5920));
 sg13g2_nand2_2 _32668_ (.Y(_02357_),
    .A(net5245),
    .B(net5938));
 sg13g2_and2_1 _32669_ (.A(net5235),
    .B(net5937),
    .X(_02358_));
 sg13g2_nand2_1 _32670_ (.Y(_02359_),
    .A(net5237),
    .B(net5943));
 sg13g2_a221oi_1 _32671_ (.B2(_22960_),
    .C1(_02350_),
    .B1(net5130),
    .A1(_19842_),
    .Y(_02360_),
    .A2(_02346_));
 sg13g2_a21oi_1 _32672_ (.A1(net7184),
    .A2(net6389),
    .Y(_00460_),
    .B1(_02360_));
 sg13g2_nor2_1 _32673_ (.A(net5987),
    .B(net5954),
    .Y(_02361_));
 sg13g2_nand2_2 _32674_ (.Y(_02362_),
    .A(net6003),
    .B(net5918));
 sg13g2_a21oi_2 _32675_ (.B1(net5880),
    .Y(_02363_),
    .A2(net5315),
    .A1(net5319));
 sg13g2_nand2_2 _32676_ (.Y(_02364_),
    .A(net5278),
    .B(net5902));
 sg13g2_a21oi_1 _32677_ (.A1(_22949_),
    .A2(net5941),
    .Y(_02365_),
    .B1(net7017));
 sg13g2_a22oi_1 _32678_ (.Y(_02366_),
    .B1(net5202),
    .B2(_22960_),
    .A2(net5157),
    .A1(_19842_));
 sg13g2_o21ai_1 _32679_ (.B1(net6481),
    .Y(_02367_),
    .A1(net1924),
    .A2(net7088));
 sg13g2_a21o_1 _32680_ (.A2(_02366_),
    .A1(_02365_),
    .B1(_02367_),
    .X(_02368_));
 sg13g2_o21ai_1 _32681_ (.B1(_02368_),
    .Y(_00461_),
    .A1(_18098_),
    .A2(net6481));
 sg13g2_nor2_1 _32682_ (.A(net7039),
    .B(net5242),
    .Y(_02369_));
 sg13g2_nand2_2 _32683_ (.Y(_02370_),
    .A(net7111),
    .B(net5159));
 sg13g2_a22oi_1 _32684_ (.Y(_02371_),
    .B1(net5886),
    .B2(_22949_),
    .A2(net5941),
    .A1(_22943_));
 sg13g2_nand2b_1 _32685_ (.Y(_02372_),
    .B(net5236),
    .A_N(_02371_));
 sg13g2_a221oi_1 _32686_ (.B2(net5111),
    .C1(net6388),
    .B1(_22960_),
    .A1(net1537),
    .Y(_02373_),
    .A2(net7017));
 sg13g2_a22oi_1 _32687_ (.Y(_00462_),
    .B1(_02372_),
    .B2(_02373_),
    .A2(net6388),
    .A1(_18097_));
 sg13g2_nor2_2 _32688_ (.A(net5241),
    .B(net6842),
    .Y(_02374_));
 sg13g2_nand2_2 _32689_ (.Y(_02375_),
    .A(net5162),
    .B(net6881));
 sg13g2_and2_1 _32690_ (.A(net5235),
    .B(net5884),
    .X(_02376_));
 sg13g2_nand2_2 _32691_ (.Y(_02377_),
    .A(net5237),
    .B(net5898));
 sg13g2_and2_1 _32692_ (.A(net1648),
    .B(net7021),
    .X(_02378_));
 sg13g2_a221oi_1 _32693_ (.B2(_22943_),
    .C1(_02378_),
    .B1(net5079),
    .A1(_22937_),
    .Y(_02379_),
    .A2(net5134));
 sg13g2_a22oi_1 _32694_ (.Y(_02380_),
    .B1(_22949_),
    .B2(net5095),
    .A2(net6388),
    .A1(net3690));
 sg13g2_o21ai_1 _32695_ (.B1(_02380_),
    .Y(_00463_),
    .A1(net6388),
    .A2(_02379_));
 sg13g2_nand2b_1 _32696_ (.Y(_02381_),
    .B(net6482),
    .A_N(net1295));
 sg13g2_a22oi_1 _32697_ (.Y(_02382_),
    .B1(_02381_),
    .B2(net6837),
    .A2(net5079),
    .A1(_22937_));
 sg13g2_a22oi_1 _32698_ (.Y(_02383_),
    .B1(net5111),
    .B2(_22943_),
    .A2(net5134),
    .A1(_22931_));
 sg13g2_a22oi_1 _32699_ (.Y(_00464_),
    .B1(_02382_),
    .B2(_02383_),
    .A2(net6391),
    .A1(_18096_));
 sg13g2_nand2_1 _32700_ (.Y(_02384_),
    .A(net2327),
    .B(net6392));
 sg13g2_a22oi_1 _32701_ (.Y(_02385_),
    .B1(net5886),
    .B2(_22931_),
    .A2(net5970),
    .A1(_22937_));
 sg13g2_nand2_1 _32702_ (.Y(_02386_),
    .A(net7089),
    .B(_02385_));
 sg13g2_a21oi_1 _32703_ (.A1(_22925_),
    .A2(net5941),
    .Y(_02387_),
    .B1(_02386_));
 sg13g2_o21ai_1 _32704_ (.B1(net6482),
    .Y(_02388_),
    .A1(net1888),
    .A2(net7089));
 sg13g2_o21ai_1 _32705_ (.B1(_02384_),
    .Y(_00465_),
    .A1(_02387_),
    .A2(_02388_));
 sg13g2_nor2_1 _32706_ (.A(net2774),
    .B(net6482),
    .Y(_02389_));
 sg13g2_a22oi_1 _32707_ (.Y(_02390_),
    .B1(net5886),
    .B2(_22925_),
    .A2(net5971),
    .A1(_22931_));
 sg13g2_nor2_1 _32708_ (.A(net7020),
    .B(_02390_),
    .Y(_02391_));
 sg13g2_a221oi_1 _32709_ (.B2(net5135),
    .C1(_02391_),
    .B1(_22919_),
    .A1(net1567),
    .Y(_02392_),
    .A2(net7020));
 sg13g2_a21oi_1 _32710_ (.A1(net6482),
    .A2(_02392_),
    .Y(_00466_),
    .B1(_02389_));
 sg13g2_nand2_1 _32711_ (.Y(_02393_),
    .A(_22925_),
    .B(net5095));
 sg13g2_a221oi_1 _32712_ (.B2(net5080),
    .C1(net6399),
    .B1(_22919_),
    .A1(net1760),
    .Y(_02394_),
    .A2(net7024));
 sg13g2_o21ai_1 _32713_ (.B1(_02394_),
    .Y(_02395_),
    .A1(_22913_),
    .A2(net5124));
 sg13g2_o21ai_1 _32714_ (.B1(_02395_),
    .Y(_02396_),
    .A1(net2132),
    .A2(net6482));
 sg13g2_nand2_1 _32715_ (.Y(_00467_),
    .A(_02393_),
    .B(_02396_));
 sg13g2_nor2_1 _32716_ (.A(_22913_),
    .B(net5070),
    .Y(_02397_));
 sg13g2_nand2_1 _32717_ (.Y(_02398_),
    .A(net1293),
    .B(net7025));
 sg13g2_o21ai_1 _32718_ (.B1(_02398_),
    .Y(_02399_),
    .A1(_22907_),
    .A2(net5125));
 sg13g2_o21ai_1 _32719_ (.B1(net6485),
    .Y(_02400_),
    .A1(_02397_),
    .A2(_02399_));
 sg13g2_a22oi_1 _32720_ (.Y(_02401_),
    .B1(_22919_),
    .B2(net5095),
    .A2(net6392),
    .A1(net3644));
 sg13g2_nand2_1 _32721_ (.Y(_00468_),
    .A(_02400_),
    .B(_02401_));
 sg13g2_a221oi_1 _32722_ (.B2(net5137),
    .C1(net6400),
    .B1(_22901_),
    .A1(net1391),
    .Y(_02402_),
    .A2(net7025));
 sg13g2_o21ai_1 _32723_ (.B1(_02402_),
    .Y(_02403_),
    .A1(_22907_),
    .A2(net5070));
 sg13g2_o21ai_1 _32724_ (.B1(_02403_),
    .Y(_02404_),
    .A1(net3740),
    .A2(net6485));
 sg13g2_o21ai_1 _32725_ (.B1(_02404_),
    .Y(_00469_),
    .A1(_22913_),
    .A2(net5066));
 sg13g2_nor2_1 _32726_ (.A(net3141),
    .B(net6485),
    .Y(_02405_));
 sg13g2_nand2b_1 _32727_ (.Y(_02406_),
    .B(net5977),
    .A_N(_22907_));
 sg13g2_o21ai_1 _32728_ (.B1(_02406_),
    .Y(_02407_),
    .A1(_22900_),
    .A2(net5880));
 sg13g2_and2_1 _32729_ (.A(net7095),
    .B(_02407_),
    .X(_02408_));
 sg13g2_a221oi_1 _32730_ (.B2(net5137),
    .C1(_02408_),
    .B1(_22894_),
    .A1(net1331),
    .Y(_02409_),
    .A2(net7025));
 sg13g2_a21oi_1 _32731_ (.A1(net6485),
    .A2(_02409_),
    .Y(_00470_),
    .B1(_02405_));
 sg13g2_nand2_1 _32732_ (.Y(_02410_),
    .A(net1684),
    .B(net6400));
 sg13g2_o21ai_1 _32733_ (.B1(net7095),
    .Y(_02411_),
    .A1(_22900_),
    .A2(net6004));
 sg13g2_a221oi_1 _32734_ (.B2(_22894_),
    .C1(_02411_),
    .B1(net5892),
    .A1(_22888_),
    .Y(_02412_),
    .A2(net5943));
 sg13g2_o21ai_1 _32735_ (.B1(net6486),
    .Y(_02413_),
    .A1(net1448),
    .A2(net7095));
 sg13g2_o21ai_1 _32736_ (.B1(_02410_),
    .Y(_00471_),
    .A1(_02412_),
    .A2(_02413_));
 sg13g2_nand2b_1 _32737_ (.Y(_02414_),
    .B(net6486),
    .A_N(net1274));
 sg13g2_a22oi_1 _32738_ (.Y(_02415_),
    .B1(net5080),
    .B2(_22888_),
    .A2(net5137),
    .A1(_22882_));
 sg13g2_a22oi_1 _32739_ (.Y(_02416_),
    .B1(_02414_),
    .B2(net6842),
    .A2(net5112),
    .A1(_22894_));
 sg13g2_a22oi_1 _32740_ (.Y(_00472_),
    .B1(_02415_),
    .B2(_02416_),
    .A2(net6400),
    .A1(_18094_));
 sg13g2_a22oi_1 _32741_ (.Y(_02417_),
    .B1(net5112),
    .B2(_22888_),
    .A2(net5137),
    .A1(_22875_));
 sg13g2_a221oi_1 _32742_ (.B2(net5091),
    .C1(net6402),
    .B1(_22882_),
    .A1(net1694),
    .Y(_02418_),
    .A2(net7029));
 sg13g2_a22oi_1 _32743_ (.Y(_00473_),
    .B1(_02417_),
    .B2(_02418_),
    .A2(net6402),
    .A1(_18093_));
 sg13g2_nand2b_1 _32744_ (.Y(_02419_),
    .B(net6487),
    .A_N(net1302));
 sg13g2_a22oi_1 _32745_ (.Y(_02420_),
    .B1(_02419_),
    .B2(net6844),
    .A2(net5091),
    .A1(_22875_));
 sg13g2_a22oi_1 _32746_ (.Y(_02421_),
    .B1(net5112),
    .B2(_22882_),
    .A2(net5138),
    .A1(_22870_));
 sg13g2_a22oi_1 _32747_ (.Y(_00474_),
    .B1(_02420_),
    .B2(_02421_),
    .A2(net6402),
    .A1(_18092_));
 sg13g2_nand2_1 _32748_ (.Y(_02422_),
    .A(net2124),
    .B(net6403));
 sg13g2_a21o_1 _32749_ (.A2(net5946),
    .A1(_22864_),
    .B1(net7031),
    .X(_02423_));
 sg13g2_a221oi_1 _32750_ (.B2(_22870_),
    .C1(_02423_),
    .B1(net5203),
    .A1(_22875_),
    .Y(_02424_),
    .A2(net5158));
 sg13g2_o21ai_1 _32751_ (.B1(net6490),
    .Y(_02425_),
    .A1(net1612),
    .A2(net7096));
 sg13g2_o21ai_1 _32752_ (.B1(_02422_),
    .Y(_00475_),
    .A1(_02424_),
    .A2(_02425_));
 sg13g2_nand2_1 _32753_ (.Y(_02426_),
    .A(net2635),
    .B(net6411));
 sg13g2_a22oi_1 _32754_ (.Y(_02427_),
    .B1(net5896),
    .B2(_22864_),
    .A2(net5980),
    .A1(_22870_));
 sg13g2_nand2_1 _32755_ (.Y(_02428_),
    .A(net7104),
    .B(_02427_));
 sg13g2_a21oi_1 _32756_ (.A1(_22859_),
    .A2(net5947),
    .Y(_02429_),
    .B1(_02428_));
 sg13g2_o21ai_1 _32757_ (.B1(net6488),
    .Y(_02430_),
    .A1(net1870),
    .A2(net7104));
 sg13g2_o21ai_1 _32758_ (.B1(_02426_),
    .Y(_00476_),
    .A1(_02429_),
    .A2(_02430_));
 sg13g2_nor2_1 _32759_ (.A(net2845),
    .B(net6488),
    .Y(_02431_));
 sg13g2_a22oi_1 _32760_ (.Y(_02432_),
    .B1(net5947),
    .B2(_22853_),
    .A2(net5981),
    .A1(_22864_));
 sg13g2_nor2_1 _32761_ (.A(net7032),
    .B(_02432_),
    .Y(_02433_));
 sg13g2_a221oi_1 _32762_ (.B2(net5091),
    .C1(_02433_),
    .B1(_22859_),
    .A1(net1452),
    .Y(_02434_),
    .A2(net7032));
 sg13g2_a21oi_1 _32763_ (.A1(net6488),
    .A2(_02434_),
    .Y(_00477_),
    .B1(_02431_));
 sg13g2_a22oi_1 _32764_ (.Y(_02435_),
    .B1(net5897),
    .B2(_22853_),
    .A2(net5981),
    .A1(_22859_));
 sg13g2_nor2_1 _32765_ (.A(net7033),
    .B(_02435_),
    .Y(_02436_));
 sg13g2_a21oi_1 _32766_ (.A1(net1369),
    .A2(net7033),
    .Y(_02437_),
    .B1(_02436_));
 sg13g2_o21ai_1 _32767_ (.B1(_02437_),
    .Y(_02438_),
    .A1(_22974_),
    .A2(net5125));
 sg13g2_mux2_1 _32768_ (.A0(net3520),
    .A1(_02438_),
    .S(net6488),
    .X(_00478_));
 sg13g2_nor2_1 _32769_ (.A(_22974_),
    .B(net5070),
    .Y(_02439_));
 sg13g2_a221oi_1 _32770_ (.B2(net5139),
    .C1(_02439_),
    .B1(_22847_),
    .A1(net2053),
    .Y(_02440_),
    .A2(net7033));
 sg13g2_a22oi_1 _32771_ (.Y(_02441_),
    .B1(_22853_),
    .B2(net5098),
    .A2(net6413),
    .A1(net3482));
 sg13g2_o21ai_1 _32772_ (.B1(_02441_),
    .Y(_00479_),
    .A1(net6413),
    .A2(_02440_));
 sg13g2_a221oi_1 _32773_ (.B2(_22847_),
    .C1(net7033),
    .B1(net5205),
    .A1(_22834_),
    .Y(_02442_),
    .A2(net5948));
 sg13g2_o21ai_1 _32774_ (.B1(_02442_),
    .Y(_02443_),
    .A1(_22974_),
    .A2(net5241));
 sg13g2_o21ai_1 _32775_ (.B1(net6489),
    .Y(_02444_),
    .A1(net1375),
    .A2(net7105));
 sg13g2_nand2b_1 _32776_ (.Y(_02445_),
    .B(_02443_),
    .A_N(_02444_));
 sg13g2_o21ai_1 _32777_ (.B1(_02445_),
    .Y(_00480_),
    .A1(_18090_),
    .A2(net6489));
 sg13g2_nand2_1 _32778_ (.Y(_02446_),
    .A(net2780),
    .B(net6413));
 sg13g2_o21ai_1 _32779_ (.B1(net7105),
    .Y(_02447_),
    .A1(_22840_),
    .A2(net5924));
 sg13g2_a221oi_1 _32780_ (.B2(_22834_),
    .C1(_02447_),
    .B1(net5205),
    .A1(_22847_),
    .Y(_02448_),
    .A2(net5158));
 sg13g2_o21ai_1 _32781_ (.B1(net6489),
    .Y(_02449_),
    .A1(net1692),
    .A2(net7105));
 sg13g2_o21ai_1 _32782_ (.B1(_02446_),
    .Y(_00481_),
    .A1(_02448_),
    .A2(_02449_));
 sg13g2_nor2_1 _32783_ (.A(_22840_),
    .B(net5071),
    .Y(_02450_));
 sg13g2_a221oi_1 _32784_ (.B2(net5113),
    .C1(net6420),
    .B1(_22834_),
    .A1(net1509),
    .Y(_02451_),
    .A2(net7036));
 sg13g2_a21oi_1 _32785_ (.A1(_22823_),
    .A2(net5141),
    .Y(_02452_),
    .B1(_02450_));
 sg13g2_a22oi_1 _32786_ (.Y(_00482_),
    .B1(_02451_),
    .B2(_02452_),
    .A2(net6420),
    .A1(_18089_));
 sg13g2_nand2_1 _32787_ (.Y(_02453_),
    .A(net3303),
    .B(net6420));
 sg13g2_a21oi_1 _32788_ (.A1(_22816_),
    .A2(net5948),
    .Y(_02454_),
    .B1(net7036));
 sg13g2_o21ai_1 _32789_ (.B1(_02454_),
    .Y(_02455_),
    .A1(_22840_),
    .A2(net5242));
 sg13g2_a21oi_1 _32790_ (.A1(_22823_),
    .A2(net5207),
    .Y(_02456_),
    .B1(_02455_));
 sg13g2_o21ai_1 _32791_ (.B1(net6491),
    .Y(_02457_),
    .A1(net1335),
    .A2(net7114));
 sg13g2_o21ai_1 _32792_ (.B1(_02453_),
    .Y(_00483_),
    .A1(_02456_),
    .A2(_02457_));
 sg13g2_nand2b_1 _32793_ (.Y(_02458_),
    .B(net6491),
    .A_N(net1450));
 sg13g2_a22oi_1 _32794_ (.Y(_02459_),
    .B1(_02458_),
    .B2(net6846),
    .A2(net5141),
    .A1(_22811_));
 sg13g2_a22oi_1 _32795_ (.Y(_02460_),
    .B1(net5081),
    .B2(_22816_),
    .A2(net5113),
    .A1(_22823_));
 sg13g2_a22oi_1 _32796_ (.Y(_00484_),
    .B1(_02459_),
    .B2(_02460_),
    .A2(net6420),
    .A1(_18088_));
 sg13g2_a221oi_1 _32797_ (.B2(net5081),
    .C1(net6421),
    .B1(_22811_),
    .A1(net1557),
    .Y(_02461_),
    .A2(net7037));
 sg13g2_a22oi_1 _32798_ (.Y(_02462_),
    .B1(net5113),
    .B2(_22816_),
    .A2(net5140),
    .A1(_22803_));
 sg13g2_a22oi_1 _32799_ (.Y(_00485_),
    .B1(_02461_),
    .B2(_02462_),
    .A2(net6422),
    .A1(_18087_));
 sg13g2_nand2_1 _32800_ (.Y(_02463_),
    .A(net2422),
    .B(net6424));
 sg13g2_a22oi_1 _32801_ (.Y(_02464_),
    .B1(net5907),
    .B2(_22803_),
    .A2(net5989),
    .A1(_22811_));
 sg13g2_nand2_1 _32802_ (.Y(_02465_),
    .A(net7117),
    .B(_02464_));
 sg13g2_a21oi_1 _32803_ (.A1(_22797_),
    .A2(net5955),
    .Y(_02466_),
    .B1(_02465_));
 sg13g2_o21ai_1 _32804_ (.B1(net6493),
    .Y(_02467_),
    .A1(net1343),
    .A2(net7117));
 sg13g2_o21ai_1 _32805_ (.B1(_02463_),
    .Y(_00486_),
    .A1(_02466_),
    .A2(_02467_));
 sg13g2_nor2_1 _32806_ (.A(_22790_),
    .B(net5127),
    .Y(_02468_));
 sg13g2_a221oi_1 _32807_ (.B2(net5084),
    .C1(_02468_),
    .B1(_22797_),
    .A1(net1318),
    .Y(_02469_),
    .A2(net7045));
 sg13g2_a22oi_1 _32808_ (.Y(_02470_),
    .B1(_22803_),
    .B2(net5103),
    .A2(net6432),
    .A1(net3632));
 sg13g2_o21ai_1 _32809_ (.B1(_02470_),
    .Y(_00487_),
    .A1(net6432),
    .A2(_02469_));
 sg13g2_nor2_1 _32810_ (.A(_22790_),
    .B(net5071),
    .Y(_02471_));
 sg13g2_a221oi_1 _32811_ (.B2(net5142),
    .C1(_02471_),
    .B1(_22779_),
    .A1(net1379),
    .Y(_02472_),
    .A2(net7047));
 sg13g2_a22oi_1 _32812_ (.Y(_02473_),
    .B1(_22797_),
    .B2(net5103),
    .A2(net6432),
    .A1(net3704));
 sg13g2_o21ai_1 _32813_ (.B1(_02473_),
    .Y(_00488_),
    .A1(net6432),
    .A2(_02472_));
 sg13g2_nor2_1 _32814_ (.A(net3532),
    .B(net6497),
    .Y(_02474_));
 sg13g2_nand2b_1 _32815_ (.Y(_02475_),
    .B(net5992),
    .A_N(_22790_));
 sg13g2_nand2b_1 _32816_ (.Y(_02476_),
    .B(net5958),
    .A_N(_22784_));
 sg13g2_a21oi_1 _32817_ (.A1(_02475_),
    .A2(_02476_),
    .Y(_02477_),
    .B1(net7045));
 sg13g2_a221oi_1 _32818_ (.B2(net5082),
    .C1(_02477_),
    .B1(_22779_),
    .A1(net1299),
    .Y(_02478_),
    .A2(net7047));
 sg13g2_a21oi_1 _32819_ (.A1(net6497),
    .A2(_02478_),
    .Y(_00489_),
    .B1(_02474_));
 sg13g2_nor2_1 _32820_ (.A(_22784_),
    .B(net5074),
    .Y(_02479_));
 sg13g2_a221oi_1 _32821_ (.B2(net5142),
    .C1(_02479_),
    .B1(_22766_),
    .A1(net1744),
    .Y(_02480_),
    .A2(net7048));
 sg13g2_a22oi_1 _32822_ (.Y(_02481_),
    .B1(_22779_),
    .B2(net5103),
    .A2(net6434),
    .A1(net3713));
 sg13g2_o21ai_1 _32823_ (.B1(_02481_),
    .Y(_00490_),
    .A1(net6434),
    .A2(_02480_));
 sg13g2_o21ai_1 _32824_ (.B1(net6857),
    .Y(_02482_),
    .A1(net1500),
    .A2(net6434));
 sg13g2_o21ai_1 _32825_ (.B1(_02482_),
    .Y(_02483_),
    .A1(_22784_),
    .A2(_02370_));
 sg13g2_a221oi_1 _32826_ (.B2(_22766_),
    .C1(_02483_),
    .B1(net5082),
    .A1(_22988_),
    .Y(_02484_),
    .A2(net5142));
 sg13g2_a21oi_1 _32827_ (.A1(_18086_),
    .A2(net6432),
    .Y(_00491_),
    .B1(_02484_));
 sg13g2_nand2b_1 _32828_ (.Y(_02485_),
    .B(net6495),
    .A_N(net1268));
 sg13g2_a22oi_1 _32829_ (.Y(_02486_),
    .B1(_02485_),
    .B2(net6857),
    .A2(net5082),
    .A1(_22988_));
 sg13g2_a22oi_1 _32830_ (.Y(_02487_),
    .B1(net5114),
    .B2(_22766_),
    .A2(net5143),
    .A1(_22997_));
 sg13g2_a22oi_1 _32831_ (.Y(_00492_),
    .B1(_02486_),
    .B2(_02487_),
    .A2(net6434),
    .A1(_18085_));
 sg13g2_nand2_1 _32832_ (.Y(_02488_),
    .A(net2832),
    .B(net6434));
 sg13g2_a21o_1 _32833_ (.A2(net5958),
    .A1(_22757_),
    .B1(net7049),
    .X(_02489_));
 sg13g2_a221oi_1 _32834_ (.B2(_22997_),
    .C1(_02489_),
    .B1(net5213),
    .A1(_22988_),
    .Y(_02490_),
    .A2(net5161));
 sg13g2_o21ai_1 _32835_ (.B1(net6495),
    .Y(_02491_),
    .A1(net1420),
    .A2(net7123));
 sg13g2_o21ai_1 _32836_ (.B1(_02488_),
    .Y(_00493_),
    .A1(_02490_),
    .A2(_02491_));
 sg13g2_and2_1 _32837_ (.A(net1345),
    .B(net7048),
    .X(_02492_));
 sg13g2_a221oi_1 _32838_ (.B2(_22757_),
    .C1(_02492_),
    .B1(net5082),
    .A1(_22751_),
    .Y(_02493_),
    .A2(net5143));
 sg13g2_a22oi_1 _32839_ (.Y(_02494_),
    .B1(_22997_),
    .B2(net5103),
    .A2(net6435),
    .A1(net3205));
 sg13g2_o21ai_1 _32840_ (.B1(_02494_),
    .Y(_00494_),
    .A1(net6435),
    .A2(_02493_));
 sg13g2_nand2b_1 _32841_ (.Y(_02495_),
    .B(net6495),
    .A_N(net1256));
 sg13g2_a22oi_1 _32842_ (.Y(_02496_),
    .B1(_02495_),
    .B2(net6857),
    .A2(net5144),
    .A1(_22730_));
 sg13g2_a22oi_1 _32843_ (.Y(_02497_),
    .B1(net5083),
    .B2(_22751_),
    .A2(net5115),
    .A1(_22757_));
 sg13g2_a22oi_1 _32844_ (.Y(_00495_),
    .B1(_02496_),
    .B2(_02497_),
    .A2(net6435),
    .A1(_18084_));
 sg13g2_nand2b_1 _32845_ (.Y(_02498_),
    .B(net6495),
    .A_N(net1264));
 sg13g2_a22oi_1 _32846_ (.Y(_02499_),
    .B1(_02498_),
    .B2(net6857),
    .A2(net5144),
    .A1(_22666_));
 sg13g2_a22oi_1 _32847_ (.Y(_02500_),
    .B1(net5085),
    .B2(_22730_),
    .A2(net5115),
    .A1(_22751_));
 sg13g2_a22oi_1 _32848_ (.Y(_00496_),
    .B1(_02499_),
    .B2(_02500_),
    .A2(net6434),
    .A1(_18083_));
 sg13g2_nand2_1 _32849_ (.Y(_02501_),
    .A(net1446),
    .B(net6435));
 sg13g2_a21o_1 _32850_ (.A2(net5958),
    .A1(_22742_),
    .B1(net7049),
    .X(_02502_));
 sg13g2_a221oi_1 _32851_ (.B2(_22666_),
    .C1(_02502_),
    .B1(net5213),
    .A1(_22730_),
    .Y(_02503_),
    .A2(net5161));
 sg13g2_o21ai_1 _32852_ (.B1(net6495),
    .Y(_02504_),
    .A1(\u_inv.input_reg[37] ),
    .A2(net7124));
 sg13g2_o21ai_1 _32853_ (.B1(_02501_),
    .Y(_00497_),
    .A1(_02503_),
    .A2(_02504_));
 sg13g2_a22oi_1 _32854_ (.Y(_02505_),
    .B1(net5085),
    .B2(_22742_),
    .A2(net5115),
    .A1(_22666_));
 sg13g2_a221oi_1 _32855_ (.B2(net5144),
    .C1(net6446),
    .B1(_22718_),
    .A1(net1351),
    .Y(_02506_),
    .A2(net7053));
 sg13g2_a22oi_1 _32856_ (.Y(_00498_),
    .B1(_02505_),
    .B2(_02506_),
    .A2(net6446),
    .A1(_18082_));
 sg13g2_a21oi_1 _32857_ (.A1(net1304),
    .A2(net7048),
    .Y(_02507_),
    .B1(net6434));
 sg13g2_a22oi_1 _32858_ (.Y(_02508_),
    .B1(net5908),
    .B2(_22718_),
    .A2(net5993),
    .A1(_22742_));
 sg13g2_nor2_1 _32859_ (.A(net7053),
    .B(_02508_),
    .Y(_02509_));
 sg13g2_a21oi_1 _32860_ (.A1(_22647_),
    .A2(net5144),
    .Y(_02510_),
    .B1(_02509_));
 sg13g2_a22oi_1 _32861_ (.Y(_00499_),
    .B1(_02507_),
    .B2(_02510_),
    .A2(net6434),
    .A1(_18081_));
 sg13g2_a21oi_1 _32862_ (.A1(net1590),
    .A2(net7053),
    .Y(_02511_),
    .B1(net6446));
 sg13g2_nand3_1 _32863_ (.B(net5993),
    .C(net5238),
    .A(_22718_),
    .Y(_02512_));
 sg13g2_nand2_1 _32864_ (.Y(_02513_),
    .A(_02511_),
    .B(_02512_));
 sg13g2_a221oi_1 _32865_ (.B2(_22647_),
    .C1(_02513_),
    .B1(net5085),
    .A1(_22634_),
    .Y(_02514_),
    .A2(net5144));
 sg13g2_a21oi_1 _32866_ (.A1(_18080_),
    .A2(net6446),
    .Y(_00500_),
    .B1(_02514_));
 sg13g2_nand2_1 _32867_ (.Y(_02515_),
    .A(net2439),
    .B(net6446));
 sg13g2_o21ai_1 _32868_ (.B1(net7129),
    .Y(_02516_),
    .A1(_22735_),
    .A2(net5930));
 sg13g2_a221oi_1 _32869_ (.B2(_22634_),
    .C1(_02516_),
    .B1(net5215),
    .A1(_22647_),
    .Y(_02517_),
    .A2(net5164));
 sg13g2_o21ai_1 _32870_ (.B1(net6500),
    .Y(_02518_),
    .A1(net2151),
    .A2(net7124));
 sg13g2_o21ai_1 _32871_ (.B1(_02515_),
    .Y(_00501_),
    .A1(_02517_),
    .A2(_02518_));
 sg13g2_a221oi_1 _32872_ (.B2(net5144),
    .C1(net6446),
    .B1(_22710_),
    .A1(net1755),
    .Y(_02519_),
    .A2(net7054));
 sg13g2_o21ai_1 _32873_ (.B1(_02519_),
    .Y(_02520_),
    .A1(_22735_),
    .A2(net5072));
 sg13g2_o21ai_1 _32874_ (.B1(_02520_),
    .Y(_02521_),
    .A1(net3738),
    .A2(net6500));
 sg13g2_o21ai_1 _32875_ (.B1(_02521_),
    .Y(_00502_),
    .A1(_22635_),
    .A2(net5065));
 sg13g2_nand2_1 _32876_ (.Y(_02522_),
    .A(net3267),
    .B(net6446));
 sg13g2_o21ai_1 _32877_ (.B1(net7129),
    .Y(_02523_),
    .A1(_22687_),
    .A2(net5930));
 sg13g2_a221oi_1 _32878_ (.B2(_22710_),
    .C1(_02523_),
    .B1(net5215),
    .A1(_22736_),
    .Y(_02524_),
    .A2(net5164));
 sg13g2_o21ai_1 _32879_ (.B1(net6500),
    .Y(_02525_),
    .A1(net1599),
    .A2(net7129));
 sg13g2_o21ai_1 _32880_ (.B1(_02522_),
    .Y(_00503_),
    .A1(_02524_),
    .A2(_02525_));
 sg13g2_nand2_1 _32881_ (.Y(_02526_),
    .A(net1971),
    .B(net6446));
 sg13g2_o21ai_1 _32882_ (.B1(net7129),
    .Y(_02527_),
    .A1(_22709_),
    .A2(net6006));
 sg13g2_a221oi_1 _32883_ (.B2(_22688_),
    .C1(_02527_),
    .B1(net5908),
    .A1(_23005_),
    .Y(_02528_),
    .A2(net5960));
 sg13g2_o21ai_1 _32884_ (.B1(net6500),
    .Y(_02529_),
    .A1(net1411),
    .A2(net7129));
 sg13g2_o21ai_1 _32885_ (.B1(_02526_),
    .Y(_00504_),
    .A1(_02528_),
    .A2(_02529_));
 sg13g2_nand2_1 _32886_ (.Y(_02530_),
    .A(net1284),
    .B(net6450));
 sg13g2_o21ai_1 _32887_ (.B1(net7129),
    .Y(_02531_),
    .A1(_22723_),
    .A2(net5930));
 sg13g2_a221oi_1 _32888_ (.B2(_23005_),
    .C1(_02531_),
    .B1(net5215),
    .A1(_22688_),
    .Y(_02532_),
    .A2(net5164));
 sg13g2_o21ai_1 _32889_ (.B1(net6500),
    .Y(_02533_),
    .A1(\u_inv.input_reg[45] ),
    .A2(net7129));
 sg13g2_o21ai_1 _32890_ (.B1(_02530_),
    .Y(_00505_),
    .A1(_02532_),
    .A2(_02533_));
 sg13g2_nor2_1 _32891_ (.A(_22723_),
    .B(net5072),
    .Y(_02534_));
 sg13g2_a221oi_1 _32892_ (.B2(net5146),
    .C1(_02534_),
    .B1(_22654_),
    .A1(net1349),
    .Y(_02535_),
    .A2(net7054));
 sg13g2_a22oi_1 _32893_ (.Y(_02536_),
    .B1(_23005_),
    .B2(net5108),
    .A2(net6450),
    .A1(net3663));
 sg13g2_o21ai_1 _32894_ (.B1(_02536_),
    .Y(_00506_),
    .A1(net6450),
    .A2(_02535_));
 sg13g2_a221oi_1 _32895_ (.B2(_22654_),
    .C1(net7058),
    .B1(net5216),
    .A1(_22642_),
    .Y(_02537_),
    .A2(net5961));
 sg13g2_o21ai_1 _32896_ (.B1(_02537_),
    .Y(_02538_),
    .A1(_22723_),
    .A2(net5243));
 sg13g2_o21ai_1 _32897_ (.B1(net6500),
    .Y(_02539_),
    .A1(net1523),
    .A2(net7130));
 sg13g2_nand2b_1 _32898_ (.Y(_02540_),
    .B(_02538_),
    .A_N(_02539_));
 sg13g2_o21ai_1 _32899_ (.B1(_02540_),
    .Y(_00507_),
    .A1(_18078_),
    .A2(net6500));
 sg13g2_nand2b_1 _32900_ (.Y(_02541_),
    .B(net6501),
    .A_N(net1262));
 sg13g2_a22oi_1 _32901_ (.Y(_02542_),
    .B1(_02541_),
    .B2(net6859),
    .A2(net5145),
    .A1(_22614_));
 sg13g2_a22oi_1 _32902_ (.Y(_02543_),
    .B1(net5086),
    .B2(_22642_),
    .A2(net5116),
    .A1(_22654_));
 sg13g2_a22oi_1 _32903_ (.Y(_00508_),
    .B1(_02542_),
    .B2(_02543_),
    .A2(net6451),
    .A1(_18077_));
 sg13g2_nand2_1 _32904_ (.Y(_02544_),
    .A(net1669),
    .B(net6451));
 sg13g2_o21ai_1 _32905_ (.B1(net7131),
    .Y(_02545_),
    .A1(_22701_),
    .A2(net5930));
 sg13g2_a221oi_1 _32906_ (.B2(_22614_),
    .C1(_02545_),
    .B1(net5216),
    .A1(_22642_),
    .Y(_02546_),
    .A2(net5165));
 sg13g2_o21ai_1 _32907_ (.B1(net6501),
    .Y(_02547_),
    .A1(net1477),
    .A2(net7129));
 sg13g2_o21ai_1 _32908_ (.B1(_02544_),
    .Y(_00509_),
    .A1(_02546_),
    .A2(_02547_));
 sg13g2_a221oi_1 _32909_ (.B2(net5145),
    .C1(net6451),
    .B1(_22695_),
    .A1(net1492),
    .Y(_02548_),
    .A2(net7058));
 sg13g2_nor2_1 _32910_ (.A(_22701_),
    .B(net5072),
    .Y(_02549_));
 sg13g2_a21oi_1 _32911_ (.A1(_22614_),
    .A2(net5115),
    .Y(_02550_),
    .B1(_02549_));
 sg13g2_a22oi_1 _32912_ (.Y(_00510_),
    .B1(_02548_),
    .B2(_02550_),
    .A2(net6451),
    .A1(_18076_));
 sg13g2_nand2_1 _32913_ (.Y(_02551_),
    .A(net2653),
    .B(net6451));
 sg13g2_o21ai_1 _32914_ (.B1(net7131),
    .Y(_02552_),
    .A1(_22701_),
    .A2(net6006));
 sg13g2_a221oi_1 _32915_ (.B2(_22695_),
    .C1(_02552_),
    .B1(net5908),
    .A1(_23011_),
    .Y(_02553_),
    .A2(net5961));
 sg13g2_o21ai_1 _32916_ (.B1(net6501),
    .Y(_02554_),
    .A1(net1490),
    .A2(net7131));
 sg13g2_o21ai_1 _32917_ (.B1(_02551_),
    .Y(_00511_),
    .A1(_02553_),
    .A2(_02554_));
 sg13g2_nand2_1 _32918_ (.Y(_02555_),
    .A(net2534),
    .B(net6451));
 sg13g2_o21ai_1 _32919_ (.B1(net7132),
    .Y(_02556_),
    .A1(_22582_),
    .A2(net5930));
 sg13g2_a221oi_1 _32920_ (.B2(_23011_),
    .C1(_02556_),
    .B1(net5216),
    .A1(_22695_),
    .Y(_02557_),
    .A2(net5164));
 sg13g2_o21ai_1 _32921_ (.B1(net6501),
    .Y(_02558_),
    .A1(net1541),
    .A2(net7131));
 sg13g2_o21ai_1 _32922_ (.B1(_02555_),
    .Y(_00512_),
    .A1(_02557_),
    .A2(_02558_));
 sg13g2_nand2_1 _32923_ (.Y(_02559_),
    .A(net3378),
    .B(net6452));
 sg13g2_o21ai_1 _32924_ (.B1(net7131),
    .Y(_02560_),
    .A1(_22620_),
    .A2(net5930));
 sg13g2_a221oi_1 _32925_ (.B2(_22583_),
    .C1(_02560_),
    .B1(net5216),
    .A1(_23011_),
    .Y(_02561_),
    .A2(net5164));
 sg13g2_o21ai_1 _32926_ (.B1(net6501),
    .Y(_02562_),
    .A1(net1890),
    .A2(net7131));
 sg13g2_o21ai_1 _32927_ (.B1(_02559_),
    .Y(_00513_),
    .A1(_02561_),
    .A2(_02562_));
 sg13g2_a22oi_1 _32928_ (.Y(_02563_),
    .B1(_22674_),
    .B2(net5149),
    .A2(net7059),
    .A1(net1467));
 sg13g2_o21ai_1 _32929_ (.B1(_02563_),
    .Y(_02564_),
    .A1(_22620_),
    .A2(net5073));
 sg13g2_a22oi_1 _32930_ (.Y(_02565_),
    .B1(_02564_),
    .B2(net6502),
    .A2(net5108),
    .A1(_22583_));
 sg13g2_o21ai_1 _32931_ (.B1(_02565_),
    .Y(_00514_),
    .A1(_18075_),
    .A2(net6502));
 sg13g2_nand2_1 _32932_ (.Y(_02566_),
    .A(net2300),
    .B(net6452));
 sg13g2_o21ai_1 _32933_ (.B1(net7132),
    .Y(_02567_),
    .A1(_22620_),
    .A2(net6006));
 sg13g2_a221oi_1 _32934_ (.B2(_22674_),
    .C1(_02567_),
    .B1(net5908),
    .A1(_22590_),
    .Y(_02568_),
    .A2(net5961));
 sg13g2_o21ai_1 _32935_ (.B1(net6502),
    .Y(_02569_),
    .A1(net1966),
    .A2(net7132));
 sg13g2_o21ai_1 _32936_ (.B1(_02566_),
    .Y(_00515_),
    .A1(_02568_),
    .A2(_02569_));
 sg13g2_nand2_1 _32937_ (.Y(_02570_),
    .A(net2879),
    .B(net6452));
 sg13g2_a22oi_1 _32938_ (.Y(_02571_),
    .B1(net5960),
    .B2(_23025_),
    .A2(net5166),
    .A1(_22674_));
 sg13g2_nand2_1 _32939_ (.Y(_02572_),
    .A(net7132),
    .B(_02571_));
 sg13g2_a21oi_1 _32940_ (.A1(_22590_),
    .A2(net5216),
    .Y(_02573_),
    .B1(_02572_));
 sg13g2_o21ai_1 _32941_ (.B1(net6501),
    .Y(_02574_),
    .A1(net1373),
    .A2(net7132));
 sg13g2_o21ai_1 _32942_ (.B1(_02570_),
    .Y(_00516_),
    .A1(_02573_),
    .A2(_02574_));
 sg13g2_a221oi_1 _32943_ (.B2(net5149),
    .C1(net6452),
    .B1(_22596_),
    .A1(net1597),
    .Y(_02575_),
    .A2(net7058));
 sg13g2_a22oi_1 _32944_ (.Y(_02576_),
    .B1(net5090),
    .B2(_23025_),
    .A2(net5117),
    .A1(_22590_));
 sg13g2_a22oi_1 _32945_ (.Y(_00517_),
    .B1(_02575_),
    .B2(_02576_),
    .A2(net6457),
    .A1(_18073_));
 sg13g2_nor2_1 _32946_ (.A(_23017_),
    .B(net5128),
    .Y(_02577_));
 sg13g2_a221oi_1 _32947_ (.B2(net5090),
    .C1(_02577_),
    .B1(_22596_),
    .A1(net1572),
    .Y(_02578_),
    .A2(net7059));
 sg13g2_a22oi_1 _32948_ (.Y(_02579_),
    .B1(_23025_),
    .B2(net5106),
    .A2(net6452),
    .A1(net3696));
 sg13g2_o21ai_1 _32949_ (.B1(net3697),
    .Y(_00518_),
    .A1(net6452),
    .A2(_02578_));
 sg13g2_a22oi_1 _32950_ (.Y(_02580_),
    .B1(_22558_),
    .B2(net5149),
    .A2(net7066),
    .A1(net1465));
 sg13g2_o21ai_1 _32951_ (.B1(_02580_),
    .Y(_02581_),
    .A1(_23017_),
    .A2(net5072));
 sg13g2_a22oi_1 _32952_ (.Y(_02582_),
    .B1(_02581_),
    .B2(net6507),
    .A2(net5106),
    .A1(_22596_));
 sg13g2_o21ai_1 _32953_ (.B1(_02582_),
    .Y(_00519_),
    .A1(_18072_),
    .A2(net6501));
 sg13g2_nand2_1 _32954_ (.Y(_02583_),
    .A(net1779),
    .B(net6457));
 sg13g2_o21ai_1 _32955_ (.B1(net7141),
    .Y(_02584_),
    .A1(_23017_),
    .A2(net6007));
 sg13g2_a221oi_1 _32956_ (.B2(_22558_),
    .C1(_02584_),
    .B1(net5915),
    .A1(_22543_),
    .Y(_02585_),
    .A2(net5963));
 sg13g2_o21ai_1 _32957_ (.B1(net6501),
    .Y(_02586_),
    .A1(net1670),
    .A2(net7131));
 sg13g2_o21ai_1 _32958_ (.B1(_02583_),
    .Y(_00520_),
    .A1(_02585_),
    .A2(_02586_));
 sg13g2_nor2_1 _32959_ (.A(_22602_),
    .B(net5128),
    .Y(_02587_));
 sg13g2_a221oi_1 _32960_ (.B2(net5117),
    .C1(net6457),
    .B1(_22558_),
    .A1(net1594),
    .Y(_02588_),
    .A2(net7066));
 sg13g2_a21oi_1 _32961_ (.A1(_22543_),
    .A2(net5088),
    .Y(_02589_),
    .B1(_02587_));
 sg13g2_a22oi_1 _32962_ (.Y(_00521_),
    .B1(_02588_),
    .B2(_02589_),
    .A2(net6457),
    .A1(_18071_));
 sg13g2_nor2_1 _32963_ (.A(_22602_),
    .B(net5072),
    .Y(_02590_));
 sg13g2_a221oi_1 _32964_ (.B2(net5149),
    .C1(_02590_),
    .B1(_22565_),
    .A1(net1825),
    .Y(_02591_),
    .A2(net7065));
 sg13g2_a22oi_1 _32965_ (.Y(_02592_),
    .B1(_22543_),
    .B2(net5106),
    .A2(net6458),
    .A1(net3666));
 sg13g2_o21ai_1 _32966_ (.B1(_02592_),
    .Y(_00522_),
    .A1(net6457),
    .A2(_02591_));
 sg13g2_o21ai_1 _32967_ (.B1(net6863),
    .Y(_02593_),
    .A1(net1417),
    .A2(net6457));
 sg13g2_nor2_1 _32968_ (.A(_22602_),
    .B(_02370_),
    .Y(_02594_));
 sg13g2_a221oi_1 _32969_ (.B2(_22565_),
    .C1(_02594_),
    .B1(net5088),
    .A1(_23060_),
    .Y(_02595_),
    .A2(net5147));
 sg13g2_a22oi_1 _32970_ (.Y(_00523_),
    .B1(_02593_),
    .B2(_02595_),
    .A2(net6457),
    .A1(_18070_));
 sg13g2_nor2_1 _32971_ (.A(_23059_),
    .B(net5072),
    .Y(_02596_));
 sg13g2_a221oi_1 _32972_ (.B2(net5147),
    .C1(_02596_),
    .B1(_23086_),
    .A1(net1616),
    .Y(_02597_),
    .A2(net7066));
 sg13g2_a22oi_1 _32973_ (.Y(_02598_),
    .B1(_22565_),
    .B2(net5106),
    .A2(net6458),
    .A1(net3657));
 sg13g2_o21ai_1 _32974_ (.B1(_02598_),
    .Y(_00524_),
    .A1(net6458),
    .A2(_02597_));
 sg13g2_nand2_1 _32975_ (.Y(_02599_),
    .A(net2494),
    .B(net6458));
 sg13g2_o21ai_1 _32976_ (.B1(net7141),
    .Y(_02600_),
    .A1(_22570_),
    .A2(net5933));
 sg13g2_a221oi_1 _32977_ (.B2(_23086_),
    .C1(_02600_),
    .B1(net5219),
    .A1(_23060_),
    .Y(_02601_),
    .A2(net5166));
 sg13g2_o21ai_1 _32978_ (.B1(net6507),
    .Y(_02602_),
    .A1(net1737),
    .A2(net7141));
 sg13g2_o21ai_1 _32979_ (.B1(_02599_),
    .Y(_00525_),
    .A1(_02601_),
    .A2(_02602_));
 sg13g2_nor2_1 _32980_ (.A(_22570_),
    .B(net5072),
    .Y(_02603_));
 sg13g2_a221oi_1 _32981_ (.B2(net5147),
    .C1(net6457),
    .B1(_22552_),
    .A1(net1601),
    .Y(_02604_),
    .A2(net7066));
 sg13g2_a21oi_1 _32982_ (.A1(_23086_),
    .A2(net5117),
    .Y(_02605_),
    .B1(_02603_));
 sg13g2_a22oi_1 _32983_ (.Y(_00526_),
    .B1(_02604_),
    .B2(_02605_),
    .A2(net6458),
    .A1(_18069_));
 sg13g2_a22oi_1 _32984_ (.Y(_02606_),
    .B1(net5915),
    .B2(_22552_),
    .A2(net5962),
    .A1(_22526_));
 sg13g2_o21ai_1 _32985_ (.B1(_02606_),
    .Y(_02607_),
    .A1(_22570_),
    .A2(net6006));
 sg13g2_a221oi_1 _32986_ (.B2(_02607_),
    .C1(net6458),
    .B1(net5238),
    .A1(net1757),
    .Y(_02608_),
    .A2(net7066));
 sg13g2_a21oi_1 _32987_ (.A1(_18068_),
    .A2(net6458),
    .Y(_00527_),
    .B1(_02608_));
 sg13g2_a221oi_1 _32988_ (.B2(net5087),
    .C1(net6461),
    .B1(_22526_),
    .A1(net1951),
    .Y(_02609_),
    .A2(net7068));
 sg13g2_o21ai_1 _32989_ (.B1(_02609_),
    .Y(_02610_),
    .A1(_22520_),
    .A2(net5126));
 sg13g2_o21ai_1 _32990_ (.B1(_02610_),
    .Y(_02611_),
    .A1(net3717),
    .A2(net6505));
 sg13g2_o21ai_1 _32991_ (.B1(_02611_),
    .Y(_00528_),
    .A1(_22551_),
    .A2(net5065));
 sg13g2_a22oi_1 _32992_ (.Y(_02612_),
    .B1(net5087),
    .B2(_22521_),
    .A2(net5147),
    .A1(_23041_));
 sg13g2_a221oi_1 _32993_ (.B2(net5117),
    .C1(net6461),
    .B1(_22526_),
    .A1(net1780),
    .Y(_02613_),
    .A2(net7068));
 sg13g2_a22oi_1 _32994_ (.Y(_00529_),
    .B1(_02612_),
    .B2(_02613_),
    .A2(net6461),
    .A1(_18067_));
 sg13g2_o21ai_1 _32995_ (.B1(net6863),
    .Y(_02614_),
    .A1(net1829),
    .A2(net6461));
 sg13g2_nor2_1 _32996_ (.A(_23040_),
    .B(net5073),
    .Y(_02615_));
 sg13g2_a221oi_1 _32997_ (.B2(_22521_),
    .C1(_02615_),
    .B1(net5117),
    .A1(_23050_),
    .Y(_02616_),
    .A2(net5148));
 sg13g2_a22oi_1 _32998_ (.Y(_00530_),
    .B1(_02614_),
    .B2(_02616_),
    .A2(net6461),
    .A1(_18066_));
 sg13g2_nand2_1 _32999_ (.Y(_02617_),
    .A(net3077),
    .B(net6461));
 sg13g2_o21ai_1 _33000_ (.B1(net7140),
    .Y(_02618_),
    .A1(_23035_),
    .A2(net5933));
 sg13g2_a221oi_1 _33001_ (.B2(_23050_),
    .C1(_02618_),
    .B1(net5219),
    .A1(_23041_),
    .Y(_02619_),
    .A2(net5166));
 sg13g2_o21ai_1 _33002_ (.B1(net6507),
    .Y(_02620_),
    .A1(net1584),
    .A2(net7141));
 sg13g2_o21ai_1 _33003_ (.B1(_02617_),
    .Y(_00531_),
    .A1(_02619_),
    .A2(_02620_));
 sg13g2_nor2_1 _33004_ (.A(_23035_),
    .B(net5073),
    .Y(_02621_));
 sg13g2_a221oi_1 _33005_ (.B2(net5147),
    .C1(_02621_),
    .B1(_23068_),
    .A1(net2085),
    .Y(_02622_),
    .A2(net7068));
 sg13g2_a22oi_1 _33006_ (.Y(_02623_),
    .B1(_23050_),
    .B2(net5106),
    .A2(net6466),
    .A1(net3647));
 sg13g2_o21ai_1 _33007_ (.B1(_02623_),
    .Y(_00532_),
    .A1(net6462),
    .A2(_02622_));
 sg13g2_a221oi_1 _33008_ (.B2(_23068_),
    .C1(net7068),
    .B1(net5219),
    .A1(_23114_),
    .Y(_02624_),
    .A2(net5962));
 sg13g2_o21ai_1 _33009_ (.B1(_02624_),
    .Y(_02625_),
    .A1(_23035_),
    .A2(net5243));
 sg13g2_o21ai_1 _33010_ (.B1(net6505),
    .Y(_02626_),
    .A1(net1471),
    .A2(net7140));
 sg13g2_nand2b_1 _33011_ (.Y(_02627_),
    .B(_02625_),
    .A_N(_02626_));
 sg13g2_o21ai_1 _33012_ (.B1(_02627_),
    .Y(_00533_),
    .A1(_18065_),
    .A2(net6505));
 sg13g2_nand2_1 _33013_ (.Y(_02628_),
    .A(net3188),
    .B(net6462));
 sg13g2_a22oi_1 _33014_ (.Y(_02629_),
    .B1(net5915),
    .B2(_23114_),
    .A2(net6001),
    .A1(_23068_));
 sg13g2_nand2_1 _33015_ (.Y(_02630_),
    .A(net7140),
    .B(_02629_));
 sg13g2_a21oi_1 _33016_ (.A1(_23156_),
    .A2(net5962),
    .Y(_02631_),
    .B1(_02630_));
 sg13g2_o21ai_1 _33017_ (.B1(net6505),
    .Y(_02632_),
    .A1(net2153),
    .A2(net7140));
 sg13g2_o21ai_1 _33018_ (.B1(_02628_),
    .Y(_00534_),
    .A1(_02631_),
    .A2(_02632_));
 sg13g2_nand2_1 _33019_ (.Y(_02633_),
    .A(net3317),
    .B(net6462));
 sg13g2_a22oi_1 _33020_ (.Y(_02634_),
    .B1(net5915),
    .B2(_23156_),
    .A2(net6001),
    .A1(_23114_));
 sg13g2_nand2_1 _33021_ (.Y(_02635_),
    .A(net7140),
    .B(_02634_));
 sg13g2_a21oi_1 _33022_ (.A1(_23175_),
    .A2(net5962),
    .Y(_02636_),
    .B1(_02635_));
 sg13g2_o21ai_1 _33023_ (.B1(net6505),
    .Y(_02637_),
    .A1(net1675),
    .A2(net7140));
 sg13g2_o21ai_1 _33024_ (.B1(_02633_),
    .Y(_00535_),
    .A1(_02636_),
    .A2(_02637_));
 sg13g2_nor2_1 _33025_ (.A(net7069),
    .B(_23169_),
    .Y(_02638_));
 sg13g2_nor2_1 _33026_ (.A(_23169_),
    .B(net5126),
    .Y(_02639_));
 sg13g2_a221oi_1 _33027_ (.B2(net5087),
    .C1(_02639_),
    .B1(_23175_),
    .A1(net2188),
    .Y(_02640_),
    .A2(net7069));
 sg13g2_a22oi_1 _33028_ (.Y(_02641_),
    .B1(_23156_),
    .B2(net5106),
    .A2(net6462),
    .A1(net3714));
 sg13g2_o21ai_1 _33029_ (.B1(_02641_),
    .Y(_00536_),
    .A1(net6466),
    .A2(_02640_));
 sg13g2_a221oi_1 _33030_ (.B2(net5147),
    .C1(net6460),
    .B1(_23091_),
    .A1(net1827),
    .Y(_02642_),
    .A2(net7068));
 sg13g2_a22oi_1 _33031_ (.Y(_02643_),
    .B1(_02638_),
    .B2(net5219),
    .A2(net5117),
    .A1(_23175_));
 sg13g2_a22oi_1 _33032_ (.Y(_00537_),
    .B1(_02642_),
    .B2(_02643_),
    .A2(net6461),
    .A1(_18064_));
 sg13g2_a221oi_1 _33033_ (.B2(_02638_),
    .C1(net6460),
    .B1(net5166),
    .A1(net2003),
    .Y(_02644_),
    .A2(net7069));
 sg13g2_inv_1 _33034_ (.Y(_02645_),
    .A(_02644_));
 sg13g2_a221oi_1 _33035_ (.B2(_23091_),
    .C1(_02645_),
    .B1(net5087),
    .A1(_23078_),
    .Y(_02646_),
    .A2(net5147));
 sg13g2_a21oi_1 _33036_ (.A1(_18063_),
    .A2(net6466),
    .Y(_00538_),
    .B1(_02646_));
 sg13g2_nand2_1 _33037_ (.Y(_02647_),
    .A(_23078_),
    .B(net5087));
 sg13g2_a22oi_1 _33038_ (.Y(_02648_),
    .B1(net5962),
    .B2(_23097_),
    .A2(net6001),
    .A1(_23091_));
 sg13g2_inv_1 _33039_ (.Y(_02649_),
    .A(_02648_));
 sg13g2_a221oi_1 _33040_ (.B2(_02649_),
    .C1(net6460),
    .B1(net5238),
    .A1(net1553),
    .Y(_02650_),
    .A2(net7066));
 sg13g2_a22oi_1 _33041_ (.Y(_00539_),
    .B1(_02647_),
    .B2(_02650_),
    .A2(net6460),
    .A1(_18062_));
 sg13g2_and2_1 _33042_ (.A(net1791),
    .B(net7069),
    .X(_02651_));
 sg13g2_a221oi_1 _33043_ (.B2(_23097_),
    .C1(_02651_),
    .B1(net5087),
    .A1(_23107_),
    .Y(_02652_),
    .A2(net5147));
 sg13g2_a22oi_1 _33044_ (.Y(_02653_),
    .B1(_23078_),
    .B2(net5106),
    .A2(net6462),
    .A1(net3627));
 sg13g2_o21ai_1 _33045_ (.B1(_02653_),
    .Y(_00540_),
    .A1(net6462),
    .A2(_02652_));
 sg13g2_nand2_1 _33046_ (.Y(_02654_),
    .A(net3185),
    .B(net6460));
 sg13g2_a21o_1 _33047_ (.A2(net5962),
    .A1(_23119_),
    .B1(net7069),
    .X(_02655_));
 sg13g2_a221oi_1 _33048_ (.B2(_23107_),
    .C1(_02655_),
    .B1(net5219),
    .A1(_23097_),
    .Y(_02656_),
    .A2(net5166));
 sg13g2_o21ai_1 _33049_ (.B1(net6505),
    .Y(_02657_),
    .A1(net1815),
    .A2(net7140));
 sg13g2_o21ai_1 _33050_ (.B1(_02654_),
    .Y(_00541_),
    .A1(_02656_),
    .A2(_02657_));
 sg13g2_a22oi_1 _33051_ (.Y(_02658_),
    .B1(net5087),
    .B2(_23119_),
    .A2(net5148),
    .A1(_23148_));
 sg13g2_a221oi_1 _33052_ (.B2(net5117),
    .C1(net6460),
    .B1(_23107_),
    .A1(net1771),
    .Y(_02659_),
    .A2(net7072));
 sg13g2_a22oi_1 _33053_ (.Y(_00542_),
    .B1(_02658_),
    .B2(_02659_),
    .A2(net6460),
    .A1(_18059_));
 sg13g2_and2_1 _33054_ (.A(net1423),
    .B(net7067),
    .X(_02660_));
 sg13g2_a221oi_1 _33055_ (.B2(_23148_),
    .C1(_02660_),
    .B1(net5087),
    .A1(_23188_),
    .Y(_02661_),
    .A2(net5148));
 sg13g2_a22oi_1 _33056_ (.Y(_02662_),
    .B1(_23119_),
    .B2(net5106),
    .A2(net6460),
    .A1(net3654));
 sg13g2_o21ai_1 _33057_ (.B1(_02662_),
    .Y(_00543_),
    .A1(net6463),
    .A2(_02661_));
 sg13g2_o21ai_1 _33058_ (.B1(net6863),
    .Y(_02663_),
    .A1(net1358),
    .A2(net6459));
 sg13g2_o21ai_1 _33059_ (.B1(_02663_),
    .Y(_02664_),
    .A1(_22461_),
    .A2(net5126));
 sg13g2_a221oi_1 _33060_ (.B2(_23188_),
    .C1(_02664_),
    .B1(net5088),
    .A1(_23148_),
    .Y(_02665_),
    .A2(net5117));
 sg13g2_a21oi_1 _33061_ (.A1(_18058_),
    .A2(net6462),
    .Y(_00544_),
    .B1(_02665_));
 sg13g2_nor2_1 _33062_ (.A(net3359),
    .B(net6506),
    .Y(_02666_));
 sg13g2_a22oi_1 _33063_ (.Y(_02667_),
    .B1(net5963),
    .B2(_23141_),
    .A2(net6001),
    .A1(_23188_));
 sg13g2_nor2_1 _33064_ (.A(net7072),
    .B(_02667_),
    .Y(_02668_));
 sg13g2_a221oi_1 _33065_ (.B2(net5088),
    .C1(_02668_),
    .B1(_22462_),
    .A1(net1934),
    .Y(_02669_),
    .A2(net7072));
 sg13g2_a21oi_1 _33066_ (.A1(net6506),
    .A2(_02669_),
    .Y(_00545_),
    .B1(_02666_));
 sg13g2_a221oi_1 _33067_ (.B2(net5088),
    .C1(net6464),
    .B1(_23141_),
    .A1(net1614),
    .Y(_02670_),
    .A2(net7072));
 sg13g2_a22oi_1 _33068_ (.Y(_02671_),
    .B1(net5118),
    .B2(_22462_),
    .A2(net5148),
    .A1(_22503_));
 sg13g2_a22oi_1 _33069_ (.Y(_00546_),
    .B1(_02670_),
    .B2(_02671_),
    .A2(net6463),
    .A1(_18057_));
 sg13g2_nand2_1 _33070_ (.Y(_02672_),
    .A(net1576),
    .B(net6464));
 sg13g2_o21ai_1 _33071_ (.B1(net7138),
    .Y(_02673_),
    .A1(_23181_),
    .A2(net5933));
 sg13g2_a221oi_1 _33072_ (.B2(_22503_),
    .C1(_02673_),
    .B1(net5219),
    .A1(_23141_),
    .Y(_02674_),
    .A2(net5166));
 sg13g2_o21ai_1 _33073_ (.B1(net6506),
    .Y(_02675_),
    .A1(net1371),
    .A2(net7138));
 sg13g2_o21ai_1 _33074_ (.B1(_02672_),
    .Y(_00547_),
    .A1(_02674_),
    .A2(_02675_));
 sg13g2_a21oi_1 _33075_ (.A1(_22503_),
    .A2(net6001),
    .Y(_02676_),
    .B1(net7072));
 sg13g2_o21ai_1 _33076_ (.B1(_02676_),
    .Y(_02677_),
    .A1(_23181_),
    .A2(net5881));
 sg13g2_a21oi_1 _33077_ (.A1(_22471_),
    .A2(net5962),
    .Y(_02678_),
    .B1(_02677_));
 sg13g2_o21ai_1 _33078_ (.B1(net6505),
    .Y(_02679_),
    .A1(net1460),
    .A2(net7138));
 sg13g2_nand2_1 _33079_ (.Y(_02680_),
    .A(net2529),
    .B(net6464));
 sg13g2_o21ai_1 _33080_ (.B1(_02680_),
    .Y(_00548_),
    .A1(_02678_),
    .A2(_02679_));
 sg13g2_nor2_1 _33081_ (.A(_22484_),
    .B(net5126),
    .Y(_02681_));
 sg13g2_a221oi_1 _33082_ (.B2(net5089),
    .C1(net6463),
    .B1(_22471_),
    .A1(net1435),
    .Y(_02682_),
    .A2(net7072));
 sg13g2_a21oi_1 _33083_ (.A1(_23182_),
    .A2(net5118),
    .Y(_02683_),
    .B1(_02681_));
 sg13g2_a22oi_1 _33084_ (.Y(_00549_),
    .B1(_02682_),
    .B2(_02683_),
    .A2(net6463),
    .A1(_18055_));
 sg13g2_a21oi_1 _33085_ (.A1(net1719),
    .A2(net7072),
    .Y(_02684_),
    .B1(net6465));
 sg13g2_nand2_1 _33086_ (.Y(_02685_),
    .A(_22471_),
    .B(net6001));
 sg13g2_o21ai_1 _33087_ (.B1(_02685_),
    .Y(_02686_),
    .A1(_22484_),
    .A2(net5881));
 sg13g2_a22oi_1 _33088_ (.Y(_02687_),
    .B1(_02686_),
    .B2(net7139),
    .A2(net5150),
    .A1(_22443_));
 sg13g2_a22oi_1 _33089_ (.Y(_00550_),
    .B1(_02684_),
    .B2(_02687_),
    .A2(net6465),
    .A1(_18054_));
 sg13g2_o21ai_1 _33090_ (.B1(net7139),
    .Y(_02688_),
    .A1(_22484_),
    .A2(net6007));
 sg13g2_a221oi_1 _33091_ (.B2(_22443_),
    .C1(_02688_),
    .B1(net5915),
    .A1(_23205_),
    .Y(_02689_),
    .A2(net5962));
 sg13g2_o21ai_1 _33092_ (.B1(net6505),
    .Y(_02690_),
    .A1(net1526),
    .A2(net7138));
 sg13g2_nand2_1 _33093_ (.Y(_02691_),
    .A(net3238),
    .B(net6465));
 sg13g2_o21ai_1 _33094_ (.B1(_02691_),
    .Y(_00551_),
    .A1(_02689_),
    .A2(_02690_));
 sg13g2_nor2_1 _33095_ (.A(_22427_),
    .B(net5126),
    .Y(_02692_));
 sg13g2_a221oi_1 _33096_ (.B2(net5089),
    .C1(_02692_),
    .B1(_23205_),
    .A1(net1533),
    .Y(_02693_),
    .A2(net7067));
 sg13g2_a22oi_1 _33097_ (.Y(_02694_),
    .B1(_22443_),
    .B2(net5107),
    .A2(net6463),
    .A1(net3678));
 sg13g2_o21ai_1 _33098_ (.B1(_02694_),
    .Y(_00552_),
    .A1(net6463),
    .A2(_02693_));
 sg13g2_nor2_1 _33099_ (.A(_22427_),
    .B(net5073),
    .Y(_02695_));
 sg13g2_a21oi_1 _33100_ (.A1(net2087),
    .A2(net7075),
    .Y(_02696_),
    .B1(net6463));
 sg13g2_a22oi_1 _33101_ (.Y(_02697_),
    .B1(net5963),
    .B2(_23193_),
    .A2(net6001),
    .A1(_23205_));
 sg13g2_nor2_1 _33102_ (.A(net7067),
    .B(_02697_),
    .Y(_02698_));
 sg13g2_nor2_1 _33103_ (.A(_02695_),
    .B(_02698_),
    .Y(_02699_));
 sg13g2_a22oi_1 _33104_ (.Y(_00553_),
    .B1(_02696_),
    .B2(_02699_),
    .A2(net6464),
    .A1(_18052_));
 sg13g2_a221oi_1 _33105_ (.B2(net5089),
    .C1(net6463),
    .B1(_23193_),
    .A1(net1608),
    .Y(_02700_),
    .A2(net7075));
 sg13g2_o21ai_1 _33106_ (.B1(_02700_),
    .Y(_02701_),
    .A1(_22492_),
    .A2(net5126));
 sg13g2_o21ai_1 _33107_ (.B1(_02701_),
    .Y(_02702_),
    .A1(net3724),
    .A2(net6506));
 sg13g2_o21ai_1 _33108_ (.B1(_02702_),
    .Y(_00554_),
    .A1(_22427_),
    .A2(net5065));
 sg13g2_nand2_1 _33109_ (.Y(_02703_),
    .A(net2545),
    .B(net6464));
 sg13g2_o21ai_1 _33110_ (.B1(net7141),
    .Y(_02704_),
    .A1(_22449_),
    .A2(net5933));
 sg13g2_a221oi_1 _33111_ (.B2(_22493_),
    .C1(_02704_),
    .B1(net5219),
    .A1(_23193_),
    .Y(_02705_),
    .A2(net5166));
 sg13g2_o21ai_1 _33112_ (.B1(net6506),
    .Y(_02706_),
    .A1(net1797),
    .A2(net7141));
 sg13g2_o21ai_1 _33113_ (.B1(_02703_),
    .Y(_00555_),
    .A1(_02705_),
    .A2(_02706_));
 sg13g2_nand2_1 _33114_ (.Y(_02707_),
    .A(net2528),
    .B(net6453));
 sg13g2_nor2_1 _33115_ (.A(_22449_),
    .B(net5120),
    .Y(_02708_));
 sg13g2_a221oi_1 _33116_ (.B2(_22436_),
    .C1(net7061),
    .B1(net5960),
    .A1(_22493_),
    .Y(_02709_),
    .A2(net5165));
 sg13g2_nor2b_1 _33117_ (.A(_02708_),
    .B_N(_02709_),
    .Y(_02710_));
 sg13g2_o21ai_1 _33118_ (.B1(net6502),
    .Y(_02711_),
    .A1(net1546),
    .A2(net7133));
 sg13g2_o21ai_1 _33119_ (.B1(_02707_),
    .Y(_00556_),
    .A1(_02710_),
    .A2(_02711_));
 sg13g2_nand2b_1 _33120_ (.Y(_02712_),
    .B(net5960),
    .A_N(_23199_));
 sg13g2_o21ai_1 _33121_ (.B1(net7133),
    .Y(_02713_),
    .A1(_22449_),
    .A2(net6006));
 sg13g2_a21oi_1 _33122_ (.A1(_22436_),
    .A2(net5908),
    .Y(_02714_),
    .B1(_02713_));
 sg13g2_o21ai_1 _33123_ (.B1(net6502),
    .Y(_02715_),
    .A1(net1365),
    .A2(net7133));
 sg13g2_a21oi_1 _33124_ (.A1(_02712_),
    .A2(_02714_),
    .Y(_02716_),
    .B1(_02715_));
 sg13g2_a21o_1 _33125_ (.A2(net6459),
    .A1(net2964),
    .B1(_02716_),
    .X(_00557_));
 sg13g2_nand2_1 _33126_ (.Y(_02717_),
    .A(net2735),
    .B(net6451));
 sg13g2_a21oi_1 _33127_ (.A1(_22436_),
    .A2(net5993),
    .Y(_02718_),
    .B1(net7060));
 sg13g2_o21ai_1 _33128_ (.B1(_02718_),
    .Y(_02719_),
    .A1(_23199_),
    .A2(net5881));
 sg13g2_a21oi_1 _33129_ (.A1(_22409_),
    .A2(net5960),
    .Y(_02720_),
    .B1(_02719_));
 sg13g2_o21ai_1 _33130_ (.B1(net6502),
    .Y(_02721_),
    .A1(net1658),
    .A2(net7131));
 sg13g2_o21ai_1 _33131_ (.B1(_02717_),
    .Y(_00558_),
    .A1(_02720_),
    .A2(_02721_));
 sg13g2_a221oi_1 _33132_ (.B2(_22409_),
    .C1(net7060),
    .B1(net5215),
    .A1(_22402_),
    .Y(_02722_),
    .A2(net5960));
 sg13g2_o21ai_1 _33133_ (.B1(_02722_),
    .Y(_02723_),
    .A1(_23199_),
    .A2(net5243));
 sg13g2_o21ai_1 _33134_ (.B1(net6502),
    .Y(_02724_),
    .A1(net1322),
    .A2(net7133));
 sg13g2_nor2b_1 _33135_ (.A(_02724_),
    .B_N(_02723_),
    .Y(_02725_));
 sg13g2_a21o_1 _33136_ (.A2(net6451),
    .A1(net3496),
    .B1(_02725_),
    .X(_00559_));
 sg13g2_nor2_1 _33137_ (.A(net3036),
    .B(net6503),
    .Y(_02726_));
 sg13g2_a22oi_1 _33138_ (.Y(_02727_),
    .B1(net5908),
    .B2(_22402_),
    .A2(net5993),
    .A1(_22409_));
 sg13g2_nor2_1 _33139_ (.A(net7060),
    .B(_02727_),
    .Y(_02728_));
 sg13g2_a221oi_1 _33140_ (.B2(net5145),
    .C1(_02728_),
    .B1(_22322_),
    .A1(net1945),
    .Y(_02729_),
    .A2(net7060));
 sg13g2_a21oi_1 _33141_ (.A1(net6503),
    .A2(_02729_),
    .Y(_00560_),
    .B1(_02726_));
 sg13g2_nand2_1 _33142_ (.Y(_02730_),
    .A(net2821),
    .B(net6453));
 sg13g2_o21ai_1 _33143_ (.B1(net7130),
    .Y(_02731_),
    .A1(_22477_),
    .A2(net5930));
 sg13g2_a221oi_1 _33144_ (.B2(_22322_),
    .C1(_02731_),
    .B1(net5215),
    .A1(_22402_),
    .Y(_02732_),
    .A2(net5164));
 sg13g2_o21ai_1 _33145_ (.B1(net6503),
    .Y(_02733_),
    .A1(net1800),
    .A2(net7130));
 sg13g2_o21ai_1 _33146_ (.B1(_02730_),
    .Y(_00561_),
    .A1(_02732_),
    .A2(_02733_));
 sg13g2_o21ai_1 _33147_ (.B1(net6859),
    .Y(_02734_),
    .A1(net1863),
    .A2(net6453));
 sg13g2_o21ai_1 _33148_ (.B1(_02734_),
    .Y(_02735_),
    .A1(_22360_),
    .A2(net5126));
 sg13g2_a221oi_1 _33149_ (.B2(_22478_),
    .C1(_02735_),
    .B1(net5086),
    .A1(_22322_),
    .Y(_02736_),
    .A2(net5116));
 sg13g2_a21oi_1 _33150_ (.A1(_18051_),
    .A2(net6453),
    .Y(_00562_),
    .B1(_02736_));
 sg13g2_nor2_1 _33151_ (.A(net3023),
    .B(net6500),
    .Y(_02737_));
 sg13g2_nor2_1 _33152_ (.A(_22360_),
    .B(net5881),
    .Y(_02738_));
 sg13g2_a21oi_1 _33153_ (.A1(_22373_),
    .A2(net5960),
    .Y(_02739_),
    .B1(_02738_));
 sg13g2_o21ai_1 _33154_ (.B1(_02739_),
    .Y(_02740_),
    .A1(_22477_),
    .A2(net6006));
 sg13g2_a22oi_1 _33155_ (.Y(_02741_),
    .B1(net5238),
    .B2(_02740_),
    .A2(net7056),
    .A1(net1409));
 sg13g2_a21oi_1 _33156_ (.A1(net6503),
    .A2(_02741_),
    .Y(_00563_),
    .B1(_02737_));
 sg13g2_a21oi_1 _33157_ (.A1(net1682),
    .A2(net7064),
    .Y(_02742_),
    .B1(net6448));
 sg13g2_nand2_1 _33158_ (.Y(_02743_),
    .A(_22373_),
    .B(net5908));
 sg13g2_o21ai_1 _33159_ (.B1(_02743_),
    .Y(_02744_),
    .A1(_22360_),
    .A2(net6006));
 sg13g2_a22oi_1 _33160_ (.Y(_02745_),
    .B1(_02744_),
    .B2(net7130),
    .A2(net5145),
    .A1(_22216_));
 sg13g2_a22oi_1 _33161_ (.Y(_00564_),
    .B1(_02742_),
    .B2(_02745_),
    .A2(net6448),
    .A1(_18050_));
 sg13g2_nand2_1 _33162_ (.Y(_02746_),
    .A(net1419),
    .B(net6453));
 sg13g2_o21ai_1 _33163_ (.B1(net7130),
    .Y(_02747_),
    .A1(_22366_),
    .A2(net5930));
 sg13g2_a221oi_1 _33164_ (.B2(_22216_),
    .C1(_02747_),
    .B1(net5215),
    .A1(_22373_),
    .Y(_02748_),
    .A2(net5164));
 sg13g2_o21ai_1 _33165_ (.B1(net6503),
    .Y(_02749_),
    .A1(net1363),
    .A2(net7130));
 sg13g2_o21ai_1 _33166_ (.B1(_02746_),
    .Y(_00565_),
    .A1(_02748_),
    .A2(_02749_));
 sg13g2_a22oi_1 _33167_ (.Y(_02750_),
    .B1(net5116),
    .B2(_22216_),
    .A2(net5145),
    .A1(_22349_));
 sg13g2_nor2_1 _33168_ (.A(net7056),
    .B(_22366_),
    .Y(_02751_));
 sg13g2_a221oi_1 _33169_ (.B2(_02751_),
    .C1(net6448),
    .B1(net5215),
    .A1(net2370),
    .Y(_02752_),
    .A2(net7056));
 sg13g2_a22oi_1 _33170_ (.Y(_00566_),
    .B1(_02750_),
    .B2(_02752_),
    .A2(net6448),
    .A1(_18048_));
 sg13g2_nand2b_1 _33171_ (.Y(_02753_),
    .B(net6504),
    .A_N(net1276));
 sg13g2_a22oi_1 _33172_ (.Y(_02754_),
    .B1(_02753_),
    .B2(net6859),
    .A2(_02751_),
    .A1(net5164));
 sg13g2_a22oi_1 _33173_ (.Y(_02755_),
    .B1(net5086),
    .B2(_22349_),
    .A2(net5145),
    .A1(_22394_));
 sg13g2_a22oi_1 _33174_ (.Y(_00567_),
    .B1(_02754_),
    .B2(_02755_),
    .A2(net6448),
    .A1(_18047_));
 sg13g2_and2_1 _33175_ (.A(net1689),
    .B(net7064),
    .X(_02756_));
 sg13g2_a221oi_1 _33176_ (.B2(_22394_),
    .C1(_02756_),
    .B1(net5086),
    .A1(_22297_),
    .Y(_02757_),
    .A2(net5146));
 sg13g2_a22oi_1 _33177_ (.Y(_02758_),
    .B1(_22349_),
    .B2(net5108),
    .A2(net6449),
    .A1(net3687));
 sg13g2_o21ai_1 _33178_ (.B1(_02758_),
    .Y(_00568_),
    .A1(net6449),
    .A2(_02757_));
 sg13g2_a221oi_1 _33179_ (.B2(net5115),
    .C1(net6447),
    .B1(_22394_),
    .A1(net1762),
    .Y(_02759_),
    .A2(net7064));
 sg13g2_a22oi_1 _33180_ (.Y(_02760_),
    .B1(net5085),
    .B2(_22297_),
    .A2(net5146),
    .A1(_22354_));
 sg13g2_a22oi_1 _33181_ (.Y(_00569_),
    .B1(_02759_),
    .B2(_02760_),
    .A2(net6448),
    .A1(_18046_));
 sg13g2_nor2_1 _33182_ (.A(_22336_),
    .B(net5126),
    .Y(_02761_));
 sg13g2_a221oi_1 _33183_ (.B2(net5085),
    .C1(net6448),
    .B1(_22354_),
    .A1(net1592),
    .Y(_02762_),
    .A2(net7064));
 sg13g2_a21oi_1 _33184_ (.A1(_22297_),
    .A2(net5116),
    .Y(_02763_),
    .B1(_02761_));
 sg13g2_a22oi_1 _33185_ (.Y(_00570_),
    .B1(_02762_),
    .B2(_02763_),
    .A2(net6448),
    .A1(_18045_));
 sg13g2_nand2_1 _33186_ (.Y(_02764_),
    .A(_22263_),
    .B(net5146));
 sg13g2_nand2_1 _33187_ (.Y(_02765_),
    .A(_22354_),
    .B(net5993));
 sg13g2_o21ai_1 _33188_ (.B1(_02765_),
    .Y(_02766_),
    .A1(_22336_),
    .A2(net5881));
 sg13g2_a221oi_1 _33189_ (.B2(_02766_),
    .C1(net6447),
    .B1(net5238),
    .A1(net1733),
    .Y(_02767_),
    .A2(net7055));
 sg13g2_a22oi_1 _33190_ (.Y(_00571_),
    .B1(_02764_),
    .B2(_02767_),
    .A2(net6447),
    .A1(_18044_));
 sg13g2_nand2_1 _33191_ (.Y(_02768_),
    .A(net2563),
    .B(net6449));
 sg13g2_a21oi_1 _33192_ (.A1(_23267_),
    .A2(net5960),
    .Y(_02769_),
    .B1(net7057));
 sg13g2_o21ai_1 _33193_ (.B1(_02769_),
    .Y(_02770_),
    .A1(_22336_),
    .A2(net5243));
 sg13g2_a21oi_1 _33194_ (.A1(_22263_),
    .A2(net5215),
    .Y(_02771_),
    .B1(_02770_));
 sg13g2_o21ai_1 _33195_ (.B1(net6504),
    .Y(_02772_),
    .A1(net1397),
    .A2(net7137));
 sg13g2_o21ai_1 _33196_ (.B1(_02768_),
    .Y(_00572_),
    .A1(_02771_),
    .A2(_02772_));
 sg13g2_nand2_1 _33197_ (.Y(_02773_),
    .A(_22328_),
    .B(net5146));
 sg13g2_a22oi_1 _33198_ (.Y(_02774_),
    .B1(net5908),
    .B2(_23267_),
    .A2(net5993),
    .A1(_22263_));
 sg13g2_inv_1 _33199_ (.Y(_02775_),
    .A(_02774_));
 sg13g2_a221oi_1 _33200_ (.B2(_02775_),
    .C1(net6447),
    .B1(_02345_),
    .A1(net1535),
    .Y(_02776_),
    .A2(net7055));
 sg13g2_a22oi_1 _33201_ (.Y(_00573_),
    .B1(_02773_),
    .B2(_02776_),
    .A2(net6447),
    .A1(_18043_));
 sg13g2_a221oi_1 _33202_ (.B2(net5146),
    .C1(net6447),
    .B1(_22236_),
    .A1(net1748),
    .Y(_02777_),
    .A2(net7055));
 sg13g2_a22oi_1 _33203_ (.Y(_02778_),
    .B1(net5085),
    .B2(_22328_),
    .A2(net5115),
    .A1(_23267_));
 sg13g2_a22oi_1 _33204_ (.Y(_00574_),
    .B1(_02777_),
    .B2(_02778_),
    .A2(net6447),
    .A1(_18042_));
 sg13g2_nor2_1 _33205_ (.A(_22235_),
    .B(net5072),
    .Y(_02779_));
 sg13g2_a221oi_1 _33206_ (.B2(net5146),
    .C1(_02779_),
    .B1(_23259_),
    .A1(net2015),
    .Y(_02780_),
    .A2(net7055));
 sg13g2_a22oi_1 _33207_ (.Y(_02781_),
    .B1(_22328_),
    .B2(net5108),
    .A2(net6449),
    .A1(net3728));
 sg13g2_o21ai_1 _33208_ (.B1(_02781_),
    .Y(_00575_),
    .A1(net6447),
    .A2(_02780_));
 sg13g2_nand2_1 _33209_ (.Y(_02782_),
    .A(net2143),
    .B(net6437));
 sg13g2_a22oi_1 _33210_ (.Y(_02783_),
    .B1(net5213),
    .B2(_23259_),
    .A2(net5958),
    .A1(_23328_));
 sg13g2_nand2_1 _33211_ (.Y(_02784_),
    .A(net7124),
    .B(_02783_));
 sg13g2_a21oi_1 _33212_ (.A1(_22236_),
    .A2(net5161),
    .Y(_02785_),
    .B1(_02784_));
 sg13g2_o21ai_1 _33213_ (.B1(net6495),
    .Y(_02786_),
    .A1(\u_inv.input_reg[116] ),
    .A2(net7124));
 sg13g2_o21ai_1 _33214_ (.B1(_02782_),
    .Y(_00576_),
    .A1(_02785_),
    .A2(_02786_));
 sg13g2_a22oi_1 _33215_ (.Y(_02787_),
    .B1(net5958),
    .B2(_22378_),
    .A2(net5161),
    .A1(_23259_));
 sg13g2_a21oi_1 _33216_ (.A1(_23328_),
    .A2(net5213),
    .Y(_02788_),
    .B1(net7050));
 sg13g2_o21ai_1 _33217_ (.B1(net6498),
    .Y(_02789_),
    .A1(net1429),
    .A2(net7126));
 sg13g2_a21o_1 _33218_ (.A2(_02788_),
    .A1(_02787_),
    .B1(_02789_),
    .X(_02790_));
 sg13g2_o21ai_1 _33219_ (.B1(_02790_),
    .Y(_00577_),
    .A1(_18041_),
    .A2(net6495));
 sg13g2_and2_1 _33220_ (.A(net1728),
    .B(net7055),
    .X(_02791_));
 sg13g2_a221oi_1 _33221_ (.B2(_22378_),
    .C1(_02791_),
    .B1(net5085),
    .A1(_22272_),
    .Y(_02792_),
    .A2(net5145));
 sg13g2_a22oi_1 _33222_ (.Y(_02793_),
    .B1(_23328_),
    .B2(net5103),
    .A2(net6436),
    .A1(net3745));
 sg13g2_o21ai_1 _33223_ (.B1(_02793_),
    .Y(_00578_),
    .A1(net6437),
    .A2(_02792_));
 sg13g2_nor2_1 _33224_ (.A(net2938),
    .B(net6495),
    .Y(_02794_));
 sg13g2_a22oi_1 _33225_ (.Y(_02795_),
    .B1(net5907),
    .B2(_22272_),
    .A2(net5992),
    .A1(_22378_));
 sg13g2_nor2_1 _33226_ (.A(net7050),
    .B(_02795_),
    .Y(_02796_));
 sg13g2_a221oi_1 _33227_ (.B2(net5144),
    .C1(_02796_),
    .B1(_23212_),
    .A1(net2569),
    .Y(_02797_),
    .A2(net7050));
 sg13g2_a21oi_1 _33228_ (.A1(net6496),
    .A2(_02797_),
    .Y(_00579_),
    .B1(_02794_));
 sg13g2_nand2b_1 _33229_ (.Y(_02798_),
    .B(net6498),
    .A_N(net1316));
 sg13g2_a22oi_1 _33230_ (.Y(_02799_),
    .B1(_02798_),
    .B2(net6857),
    .A2(net5144),
    .A1(_23320_));
 sg13g2_a22oi_1 _33231_ (.Y(_02800_),
    .B1(net5085),
    .B2(_23212_),
    .A2(net5115),
    .A1(_22272_));
 sg13g2_a22oi_1 _33232_ (.Y(_00580_),
    .B1(_02799_),
    .B2(_02800_),
    .A2(net6437),
    .A1(_18040_));
 sg13g2_nand2_1 _33233_ (.Y(_02801_),
    .A(net2844),
    .B(net6437));
 sg13g2_o21ai_1 _33234_ (.B1(net7124),
    .Y(_02802_),
    .A1(_22253_),
    .A2(net5928));
 sg13g2_a221oi_1 _33235_ (.B2(_23320_),
    .C1(_02802_),
    .B1(net5213),
    .A1(_23212_),
    .Y(_02803_),
    .A2(net5161));
 sg13g2_o21ai_1 _33236_ (.B1(net6499),
    .Y(_02804_),
    .A1(net2346),
    .A2(net7127));
 sg13g2_o21ai_1 _33237_ (.B1(_02801_),
    .Y(_00581_),
    .A1(_02803_),
    .A2(_02804_));
 sg13g2_a221oi_1 _33238_ (.B2(net5115),
    .C1(net6437),
    .B1(_23320_),
    .A1(net1656),
    .Y(_02805_),
    .A2(net7050));
 sg13g2_a22oi_1 _33239_ (.Y(_02806_),
    .B1(net5083),
    .B2(_22254_),
    .A2(net5142),
    .A1(_23220_));
 sg13g2_a22oi_1 _33240_ (.Y(_00582_),
    .B1(_02805_),
    .B2(_02806_),
    .A2(net6437),
    .A1(_18038_));
 sg13g2_nand2b_2 _33241_ (.Y(_02807_),
    .B(net6498),
    .A_N(net1258));
 sg13g2_a22oi_1 _33242_ (.Y(_02808_),
    .B1(_02807_),
    .B2(net6857),
    .A2(net5083),
    .A1(_23220_));
 sg13g2_a22oi_1 _33243_ (.Y(_02809_),
    .B1(net5114),
    .B2(_22254_),
    .A2(net5142),
    .A1(_23370_));
 sg13g2_a22oi_1 _33244_ (.Y(_00583_),
    .B1(_02808_),
    .B2(_02809_),
    .A2(net6436),
    .A1(_18037_));
 sg13g2_a221oi_1 _33245_ (.B2(net5082),
    .C1(net6436),
    .B1(_23370_),
    .A1(net3170),
    .Y(_02810_),
    .A2(net7051));
 sg13g2_nor2_1 _33246_ (.A(net7051),
    .B(_23474_),
    .Y(_02811_));
 sg13g2_a22oi_1 _33247_ (.Y(_02812_),
    .B1(_02811_),
    .B2(net5233),
    .A2(net5114),
    .A1(_23220_));
 sg13g2_a22oi_1 _33248_ (.Y(_00584_),
    .B1(_02810_),
    .B2(_02812_),
    .A2(net6436),
    .A1(_18036_));
 sg13g2_a221oi_1 _33249_ (.B2(net5114),
    .C1(net6436),
    .B1(_23370_),
    .A1(net3165),
    .Y(_02813_),
    .A2(net7051));
 sg13g2_a22oi_1 _33250_ (.Y(_02814_),
    .B1(net5213),
    .B2(_02811_),
    .A2(net5142),
    .A1(_22341_));
 sg13g2_a22oi_1 _33251_ (.Y(_00585_),
    .B1(_02813_),
    .B2(_02814_),
    .A2(net6436),
    .A1(_18035_));
 sg13g2_nand2b_1 _33252_ (.Y(_02815_),
    .B(net6496),
    .A_N(net2998));
 sg13g2_a22oi_1 _33253_ (.Y(_02816_),
    .B1(_02815_),
    .B2(net6857),
    .A2(net5082),
    .A1(_22341_));
 sg13g2_a22oi_1 _33254_ (.Y(_02817_),
    .B1(_02811_),
    .B2(net5161),
    .A2(net5142),
    .A1(_22282_));
 sg13g2_a22oi_1 _33255_ (.Y(_00586_),
    .B1(_02816_),
    .B2(_02817_),
    .A2(net6436),
    .A1(_18034_));
 sg13g2_nand2_1 _33256_ (.Y(_02818_),
    .A(net3167),
    .B(net6436));
 sg13g2_o21ai_1 _33257_ (.B1(net7122),
    .Y(_02819_),
    .A1(_23250_),
    .A2(net5928));
 sg13g2_a221oi_1 _33258_ (.B2(_22282_),
    .C1(_02819_),
    .B1(net5213),
    .A1(_22341_),
    .Y(_02820_),
    .A2(net5161));
 sg13g2_o21ai_1 _33259_ (.B1(net6496),
    .Y(_02821_),
    .A1(net1906),
    .A2(net7122));
 sg13g2_o21ai_1 _33260_ (.B1(_02818_),
    .Y(_00587_),
    .A1(_02820_),
    .A2(_02821_));
 sg13g2_nor2_1 _33261_ (.A(_23397_),
    .B(net5127),
    .Y(_02822_));
 sg13g2_a221oi_1 _33262_ (.B2(net5082),
    .C1(_02822_),
    .B1(_23251_),
    .A1(net2317),
    .Y(_02823_),
    .A2(net7046));
 sg13g2_a22oi_1 _33263_ (.Y(_02824_),
    .B1(_22282_),
    .B2(net5103),
    .A2(net6433),
    .A1(net3712));
 sg13g2_o21ai_1 _33264_ (.B1(_02824_),
    .Y(_00588_),
    .A1(net6433),
    .A2(_02823_));
 sg13g2_nand2_1 _33265_ (.Y(_02825_),
    .A(net2758),
    .B(net6433));
 sg13g2_nor2_1 _33266_ (.A(_23397_),
    .B(net5120),
    .Y(_02826_));
 sg13g2_a21oi_1 _33267_ (.A1(_22388_),
    .A2(net5958),
    .Y(_02827_),
    .B1(net7046));
 sg13g2_o21ai_1 _33268_ (.B1(_02827_),
    .Y(_02828_),
    .A1(_23250_),
    .A2(net5242));
 sg13g2_nor2_1 _33269_ (.A(_02826_),
    .B(_02828_),
    .Y(_02829_));
 sg13g2_o21ai_1 _33270_ (.B1(net6496),
    .Y(_02830_),
    .A1(net1640),
    .A2(net7122));
 sg13g2_o21ai_1 _33271_ (.B1(_02825_),
    .Y(_00589_),
    .A1(_02829_),
    .A2(_02830_));
 sg13g2_nand2_1 _33272_ (.Y(_02831_),
    .A(_22388_),
    .B(net5082));
 sg13g2_nand2_1 _33273_ (.Y(_02832_),
    .A(_23234_),
    .B(net5958));
 sg13g2_o21ai_1 _33274_ (.B1(_02832_),
    .Y(_02833_),
    .A1(_23397_),
    .A2(net6008));
 sg13g2_a221oi_1 _33275_ (.B2(_02833_),
    .C1(net6433),
    .B1(net5238),
    .A1(net2399),
    .Y(_02834_),
    .A2(net7046));
 sg13g2_a22oi_1 _33276_ (.Y(_00590_),
    .B1(_02831_),
    .B2(_02834_),
    .A2(net6433),
    .A1(_18033_));
 sg13g2_nand2_1 _33277_ (.Y(_02835_),
    .A(net2407),
    .B(net6432));
 sg13g2_a21o_1 _33278_ (.A2(net5958),
    .A1(_23403_),
    .B1(net7046),
    .X(_02836_));
 sg13g2_a221oi_1 _33279_ (.B2(_23234_),
    .C1(_02836_),
    .B1(net5213),
    .A1(_22388_),
    .Y(_02837_),
    .A2(net5161));
 sg13g2_o21ai_1 _33280_ (.B1(net6497),
    .Y(_02838_),
    .A1(net1381),
    .A2(net7122));
 sg13g2_o21ai_1 _33281_ (.B1(_02835_),
    .Y(_00591_),
    .A1(_02837_),
    .A2(_02838_));
 sg13g2_and2_1 _33282_ (.A(net1271),
    .B(net7046),
    .X(_02839_));
 sg13g2_a221oi_1 _33283_ (.B2(_23403_),
    .C1(_02839_),
    .B1(net5084),
    .A1(_23303_),
    .Y(_02840_),
    .A2(net5142));
 sg13g2_a22oi_1 _33284_ (.Y(_02841_),
    .B1(_23234_),
    .B2(net5103),
    .A2(net6432),
    .A1(net3637));
 sg13g2_o21ai_1 _33285_ (.B1(_02841_),
    .Y(_00592_),
    .A1(net6432),
    .A2(_02840_));
 sg13g2_nand2_1 _33286_ (.Y(_02842_),
    .A(net3459),
    .B(net6424));
 sg13g2_a22oi_1 _33287_ (.Y(_02843_),
    .B1(net5209),
    .B2(_23303_),
    .A2(net5955),
    .A1(_22222_));
 sg13g2_nand2_1 _33288_ (.Y(_02844_),
    .A(net7117),
    .B(_02843_));
 sg13g2_a21oi_1 _33289_ (.A1(_23403_),
    .A2(net5163),
    .Y(_02845_),
    .B1(_02844_));
 sg13g2_o21ai_1 _33290_ (.B1(net6494),
    .Y(_02846_),
    .A1(net1531),
    .A2(net7117));
 sg13g2_o21ai_1 _33291_ (.B1(_02842_),
    .Y(_00593_),
    .A1(_02845_),
    .A2(_02846_));
 sg13g2_nor2_1 _33292_ (.A(_23242_),
    .B(net5127),
    .Y(_02847_));
 sg13g2_a221oi_1 _33293_ (.B2(net5084),
    .C1(_02847_),
    .B1(_22222_),
    .A1(net1685),
    .Y(_02848_),
    .A2(net7043));
 sg13g2_a22oi_1 _33294_ (.Y(_02849_),
    .B1(_23303_),
    .B2(net5101),
    .A2(net6424),
    .A1(net3685));
 sg13g2_o21ai_1 _33295_ (.B1(_02849_),
    .Y(_00594_),
    .A1(net6424),
    .A2(_02848_));
 sg13g2_a21oi_1 _33296_ (.A1(net2552),
    .A2(net7043),
    .Y(_02850_),
    .B1(net6424));
 sg13g2_a22oi_1 _33297_ (.Y(_02851_),
    .B1(net5902),
    .B2(_23243_),
    .A2(net5989),
    .A1(_22222_));
 sg13g2_nor2_1 _33298_ (.A(net7043),
    .B(_02851_),
    .Y(_02852_));
 sg13g2_a21oi_1 _33299_ (.A1(_23409_),
    .A2(net5140),
    .Y(_02853_),
    .B1(_02852_));
 sg13g2_a22oi_1 _33300_ (.Y(_00595_),
    .B1(_02850_),
    .B2(_02853_),
    .A2(net6424),
    .A1(_18032_));
 sg13g2_nand2_1 _33301_ (.Y(_02854_),
    .A(_23312_),
    .B(net5141));
 sg13g2_a221oi_1 _33302_ (.B2(net5084),
    .C1(net6426),
    .B1(_23409_),
    .A1(net2600),
    .Y(_02855_),
    .A2(net7042));
 sg13g2_nand2_1 _33303_ (.Y(_02856_),
    .A(_02854_),
    .B(_02855_));
 sg13g2_o21ai_1 _33304_ (.B1(_02856_),
    .Y(_02857_),
    .A1(net3720),
    .A2(net6494));
 sg13g2_o21ai_1 _33305_ (.B1(_02857_),
    .Y(_00596_),
    .A1(_23242_),
    .A2(net5065));
 sg13g2_a221oi_1 _33306_ (.B2(net5113),
    .C1(net6426),
    .B1(_23409_),
    .A1(net2969),
    .Y(_02858_),
    .A2(net7042));
 sg13g2_nor2_1 _33307_ (.A(_22303_),
    .B(net5127),
    .Y(_02859_));
 sg13g2_a21oi_1 _33308_ (.A1(_23312_),
    .A2(net5081),
    .Y(_02860_),
    .B1(_02859_));
 sg13g2_a22oi_1 _33309_ (.Y(_00597_),
    .B1(_02858_),
    .B2(_02860_),
    .A2(net6426),
    .A1(_18031_));
 sg13g2_nor2_1 _33310_ (.A(_22303_),
    .B(net5071),
    .Y(_02861_));
 sg13g2_a221oi_1 _33311_ (.B2(net5143),
    .C1(_02861_),
    .B1(_23353_),
    .A1(net2229),
    .Y(_02862_),
    .A2(net7042));
 sg13g2_a22oi_1 _33312_ (.Y(_02863_),
    .B1(_23312_),
    .B2(net5101),
    .A2(net6426),
    .A1(net3630));
 sg13g2_o21ai_1 _33313_ (.B1(_02863_),
    .Y(_00598_),
    .A1(net6426),
    .A2(_02862_));
 sg13g2_a221oi_1 _33314_ (.B2(net5084),
    .C1(net6427),
    .B1(_23353_),
    .A1(net2473),
    .Y(_02864_),
    .A2(net7042));
 sg13g2_o21ai_1 _33315_ (.B1(_02864_),
    .Y(_02865_),
    .A1(_23273_),
    .A2(net5127));
 sg13g2_o21ai_1 _33316_ (.B1(_02865_),
    .Y(_02866_),
    .A1(net3737),
    .A2(net6494));
 sg13g2_o21ai_1 _33317_ (.B1(_02866_),
    .Y(_00599_),
    .A1(_22303_),
    .A2(net5065));
 sg13g2_nand2_1 _33318_ (.Y(_02867_),
    .A(net2595),
    .B(net6423));
 sg13g2_nor2_1 _33319_ (.A(_23273_),
    .B(net5121),
    .Y(_02868_));
 sg13g2_nor2_1 _33320_ (.A(_23352_),
    .B(net5242),
    .Y(_02869_));
 sg13g2_o21ai_1 _33321_ (.B1(net7115),
    .Y(_02870_),
    .A1(_22194_),
    .A2(net5926));
 sg13g2_nor3_1 _33322_ (.A(_02868_),
    .B(_02869_),
    .C(_02870_),
    .Y(_02871_));
 sg13g2_o21ai_1 _33323_ (.B1(net6492),
    .Y(_02872_),
    .A1(net1911),
    .A2(net7115));
 sg13g2_o21ai_1 _33324_ (.B1(_02867_),
    .Y(_00600_),
    .A1(_02871_),
    .A2(_02872_));
 sg13g2_nand2_1 _33325_ (.Y(_02873_),
    .A(_23226_),
    .B(net5140));
 sg13g2_nand2b_1 _33326_ (.Y(_02874_),
    .B(net5989),
    .A_N(_23273_));
 sg13g2_o21ai_1 _33327_ (.B1(_02874_),
    .Y(_02875_),
    .A1(_22194_),
    .A2(net5882));
 sg13g2_a221oi_1 _33328_ (.B2(_02875_),
    .C1(net6423),
    .B1(net5238),
    .A1(net2262),
    .Y(_02876_),
    .A2(net7038));
 sg13g2_a22oi_1 _33329_ (.Y(_00601_),
    .B1(_02873_),
    .B2(_02876_),
    .A2(net6423),
    .A1(_18029_));
 sg13g2_a21oi_1 _33330_ (.A1(net1960),
    .A2(net7038),
    .Y(_02877_),
    .B1(net6422));
 sg13g2_a22oi_1 _33331_ (.Y(_02878_),
    .B1(net5902),
    .B2(_23226_),
    .A2(net5952),
    .A1(_23342_));
 sg13g2_o21ai_1 _33332_ (.B1(_02878_),
    .Y(_02879_),
    .A1(_22194_),
    .A2(net6008));
 sg13g2_nand3_1 _33333_ (.B(net5268),
    .C(_02879_),
    .A(net7115),
    .Y(_02880_));
 sg13g2_a22oi_1 _33334_ (.Y(_00602_),
    .B1(_02877_),
    .B2(_02880_),
    .A2(net6423),
    .A1(_18028_));
 sg13g2_nand2_1 _33335_ (.Y(_02881_),
    .A(net3151),
    .B(net6421));
 sg13g2_o21ai_1 _33336_ (.B1(net7114),
    .Y(_02882_),
    .A1(_23488_),
    .A2(net5926));
 sg13g2_a221oi_1 _33337_ (.B2(_23342_),
    .C1(_02882_),
    .B1(net5209),
    .A1(_23226_),
    .Y(_02883_),
    .A2(net5163));
 sg13g2_o21ai_1 _33338_ (.B1(net6492),
    .Y(_02884_),
    .A1(net1337),
    .A2(net7115));
 sg13g2_o21ai_1 _33339_ (.B1(_02881_),
    .Y(_00603_),
    .A1(_02883_),
    .A2(_02884_));
 sg13g2_o21ai_1 _33340_ (.B1(net6850),
    .Y(_02885_),
    .A1(net2362),
    .A2(net6425));
 sg13g2_nand2_1 _33341_ (.Y(_02886_),
    .A(_23342_),
    .B(net5113));
 sg13g2_o21ai_1 _33342_ (.B1(_02885_),
    .Y(_02887_),
    .A1(_23488_),
    .A2(net5071));
 sg13g2_a21oi_1 _33343_ (.A1(_23503_),
    .A2(net5140),
    .Y(_02888_),
    .B1(_02887_));
 sg13g2_a22oi_1 _33344_ (.Y(_00604_),
    .B1(_02886_),
    .B2(_02888_),
    .A2(net6427),
    .A1(_18027_));
 sg13g2_nand2_1 _33345_ (.Y(_02889_),
    .A(net1473),
    .B(net6427));
 sg13g2_a21oi_1 _33346_ (.A1(_23279_),
    .A2(net5955),
    .Y(_02890_),
    .B1(net7040));
 sg13g2_o21ai_1 _33347_ (.B1(_02890_),
    .Y(_02891_),
    .A1(_23488_),
    .A2(net5242));
 sg13g2_a21oi_1 _33348_ (.A1(_23503_),
    .A2(net5211),
    .Y(_02892_),
    .B1(_02891_));
 sg13g2_o21ai_1 _33349_ (.B1(net6493),
    .Y(_02893_),
    .A1(\u_inv.input_reg[145] ),
    .A2(net7117));
 sg13g2_o21ai_1 _33350_ (.B1(_02889_),
    .Y(_00605_),
    .A1(_02892_),
    .A2(_02893_));
 sg13g2_nor2_1 _33351_ (.A(_22201_),
    .B(net5127),
    .Y(_02894_));
 sg13g2_a221oi_1 _33352_ (.B2(net5081),
    .C1(_02894_),
    .B1(_23279_),
    .A1(net2791),
    .Y(_02895_),
    .A2(net7040));
 sg13g2_a22oi_1 _33353_ (.Y(_02896_),
    .B1(_23503_),
    .B2(net5101),
    .A2(net6424),
    .A1(net3648));
 sg13g2_o21ai_1 _33354_ (.B1(_02896_),
    .Y(_00606_),
    .A1(net6424),
    .A2(_02895_));
 sg13g2_a22oi_1 _33355_ (.Y(_02897_),
    .B1(_22177_),
    .B2(net5140),
    .A2(net7039),
    .A1(net2495));
 sg13g2_o21ai_1 _33356_ (.B1(_02897_),
    .Y(_02898_),
    .A1(_22201_),
    .A2(net5071));
 sg13g2_a22oi_1 _33357_ (.Y(_02899_),
    .B1(_02898_),
    .B2(net6493),
    .A2(net5101),
    .A1(_23279_));
 sg13g2_o21ai_1 _33358_ (.B1(_02899_),
    .Y(_00607_),
    .A1(_18026_),
    .A2(net6493));
 sg13g2_nor2_1 _33359_ (.A(net7040),
    .B(_23512_),
    .Y(_02900_));
 sg13g2_a221oi_1 _33360_ (.B2(_02900_),
    .C1(net6425),
    .B1(net5228),
    .A1(net1885),
    .Y(_02901_),
    .A2(net7039));
 sg13g2_o21ai_1 _33361_ (.B1(_02901_),
    .Y(_02902_),
    .A1(_22176_),
    .A2(net5071));
 sg13g2_o21ai_1 _33362_ (.B1(_02902_),
    .Y(_02903_),
    .A1(net3734),
    .A2(net6493));
 sg13g2_o21ai_1 _33363_ (.B1(_02903_),
    .Y(_00608_),
    .A1(_22201_),
    .A2(net5065));
 sg13g2_a221oi_1 _33364_ (.B2(net5140),
    .C1(net6425),
    .B1(_23381_),
    .A1(net2892),
    .Y(_02904_),
    .A2(net7039));
 sg13g2_a22oi_1 _33365_ (.Y(_02905_),
    .B1(_02900_),
    .B2(net5211),
    .A2(net5113),
    .A1(_22177_));
 sg13g2_a22oi_1 _33366_ (.Y(_00609_),
    .B1(_02904_),
    .B2(_02905_),
    .A2(net6425),
    .A1(_18025_));
 sg13g2_nand2_1 _33367_ (.Y(_02906_),
    .A(_23381_),
    .B(net5081));
 sg13g2_a21oi_1 _33368_ (.A1(net1804),
    .A2(net7039),
    .Y(_02907_),
    .B1(net6425));
 sg13g2_a22oi_1 _33369_ (.Y(_02908_),
    .B1(_02900_),
    .B2(net5163),
    .A2(net5140),
    .A1(_23466_));
 sg13g2_nand3_1 _33370_ (.B(_02907_),
    .C(_02908_),
    .A(_02906_),
    .Y(_02909_));
 sg13g2_o21ai_1 _33371_ (.B1(_02909_),
    .Y(_02910_),
    .A1(net3563),
    .A2(net6493));
 sg13g2_inv_1 _33372_ (.Y(_00610_),
    .A(_02910_));
 sg13g2_nand2_1 _33373_ (.Y(_02911_),
    .A(net3230),
    .B(net6421));
 sg13g2_o21ai_1 _33374_ (.B1(net7114),
    .Y(_02912_),
    .A1(_23428_),
    .A2(net5926));
 sg13g2_a221oi_1 _33375_ (.B2(_23466_),
    .C1(_02912_),
    .B1(net5209),
    .A1(_23381_),
    .Y(_02913_),
    .A2(net5163));
 sg13g2_o21ai_1 _33376_ (.B1(net6491),
    .Y(_02914_),
    .A1(net2238),
    .A2(net7114));
 sg13g2_o21ai_1 _33377_ (.B1(_02911_),
    .Y(_00611_),
    .A1(_02913_),
    .A2(_02914_));
 sg13g2_o21ai_1 _33378_ (.B1(net6850),
    .Y(_02915_),
    .A1(net1498),
    .A2(net6425));
 sg13g2_nor2_1 _33379_ (.A(_23428_),
    .B(net5071),
    .Y(_02916_));
 sg13g2_a221oi_1 _33380_ (.B2(_23466_),
    .C1(_02916_),
    .B1(net5113),
    .A1(_01912_),
    .Y(_02917_),
    .A2(net5140));
 sg13g2_a22oi_1 _33381_ (.Y(_00612_),
    .B1(_02915_),
    .B2(_02917_),
    .A2(net6425),
    .A1(_18023_));
 sg13g2_nand2_1 _33382_ (.Y(_02918_),
    .A(net3358),
    .B(net6421));
 sg13g2_o21ai_1 _33383_ (.B1(net7114),
    .Y(_02919_),
    .A1(_23480_),
    .A2(net5926));
 sg13g2_a221oi_1 _33384_ (.B2(_01912_),
    .C1(_02919_),
    .B1(net5209),
    .A1(_23429_),
    .Y(_02920_),
    .A2(net5163));
 sg13g2_o21ai_1 _33385_ (.B1(net6491),
    .Y(_02921_),
    .A1(net1555),
    .A2(net7114));
 sg13g2_o21ai_1 _33386_ (.B1(_02918_),
    .Y(_00613_),
    .A1(_02920_),
    .A2(_02921_));
 sg13g2_nor2_1 _33387_ (.A(_23480_),
    .B(net5071),
    .Y(_02922_));
 sg13g2_a221oi_1 _33388_ (.B2(net5141),
    .C1(_02922_),
    .B1(_23449_),
    .A1(net2041),
    .Y(_02923_),
    .A2(net7037));
 sg13g2_a22oi_1 _33389_ (.Y(_02924_),
    .B1(_01912_),
    .B2(net5101),
    .A2(net6422),
    .A1(net3688));
 sg13g2_o21ai_1 _33390_ (.B1(_02924_),
    .Y(_00614_),
    .A1(net6422),
    .A2(_02923_));
 sg13g2_o21ai_1 _33391_ (.B1(net6846),
    .Y(_02925_),
    .A1(net2089),
    .A2(net6420));
 sg13g2_o21ai_1 _33392_ (.B1(_02925_),
    .Y(_02926_),
    .A1(_23480_),
    .A2(_02370_));
 sg13g2_a221oi_1 _33393_ (.B2(_23449_),
    .C1(_02926_),
    .B1(net5081),
    .A1(_23633_),
    .Y(_02927_),
    .A2(net5141));
 sg13g2_a21oi_1 _33394_ (.A1(_18021_),
    .A2(net6421),
    .Y(_00615_),
    .B1(_02927_));
 sg13g2_nand2b_1 _33395_ (.Y(_02928_),
    .B(net6491),
    .A_N(net1413));
 sg13g2_a22oi_1 _33396_ (.Y(_02929_),
    .B1(_02928_),
    .B2(net6850),
    .A2(net5081),
    .A1(_23633_));
 sg13g2_a22oi_1 _33397_ (.Y(_02930_),
    .B1(net5113),
    .B2(_23449_),
    .A2(net5141),
    .A1(_23564_));
 sg13g2_a22oi_1 _33398_ (.Y(_00616_),
    .B1(_02929_),
    .B2(_02930_),
    .A2(net6420),
    .A1(_18020_));
 sg13g2_nand2_1 _33399_ (.Y(_02931_),
    .A(net3391),
    .B(net6421));
 sg13g2_a21o_1 _33400_ (.A2(net5209),
    .A1(_23564_),
    .B1(net7037),
    .X(_02932_));
 sg13g2_a221oi_1 _33401_ (.B2(_23334_),
    .C1(_02932_),
    .B1(net5952),
    .A1(_23633_),
    .Y(_02933_),
    .A2(net5163));
 sg13g2_o21ai_1 _33402_ (.B1(net6491),
    .Y(_02934_),
    .A1(net2021),
    .A2(net7105));
 sg13g2_o21ai_1 _33403_ (.B1(_02931_),
    .Y(_00617_),
    .A1(_02933_),
    .A2(_02934_));
 sg13g2_nor2_1 _33404_ (.A(_23362_),
    .B(net5127),
    .Y(_02935_));
 sg13g2_a221oi_1 _33405_ (.B2(net5081),
    .C1(_02935_),
    .B1(_23334_),
    .A1(net1502),
    .Y(_02936_),
    .A2(net7036));
 sg13g2_a22oi_1 _33406_ (.Y(_02937_),
    .B1(_23564_),
    .B2(net5098),
    .A2(net6420),
    .A1(net3727));
 sg13g2_o21ai_1 _33407_ (.B1(_02937_),
    .Y(_00618_),
    .A1(net6421),
    .A2(_02936_));
 sg13g2_nand2b_1 _33408_ (.Y(_02938_),
    .B(net5209),
    .A_N(_23362_));
 sg13g2_a221oi_1 _33409_ (.B2(_23389_),
    .C1(net7036),
    .B1(net5952),
    .A1(_23334_),
    .Y(_02939_),
    .A2(net5163));
 sg13g2_o21ai_1 _33410_ (.B1(net6491),
    .Y(_02940_),
    .A1(net2048),
    .A2(net7105));
 sg13g2_a21oi_1 _33411_ (.A1(_02938_),
    .A2(_02939_),
    .Y(_02941_),
    .B1(_02940_));
 sg13g2_a21o_1 _33412_ (.A2(net6420),
    .A1(net3537),
    .B1(_02941_),
    .X(_00619_));
 sg13g2_nor2_1 _33413_ (.A(net3448),
    .B(net6488),
    .Y(_02942_));
 sg13g2_a22oi_1 _33414_ (.Y(_02943_),
    .B1(net5898),
    .B2(_23389_),
    .A2(net5948),
    .A1(_23457_));
 sg13g2_o21ai_1 _33415_ (.B1(_02943_),
    .Y(_02944_),
    .A1(_23362_),
    .A2(net6005));
 sg13g2_a22oi_1 _33416_ (.Y(_02945_),
    .B1(net5238),
    .B2(_02944_),
    .A2(net7033),
    .A1(net2477));
 sg13g2_a21oi_1 _33417_ (.A1(net6488),
    .A2(_02945_),
    .Y(_00620_),
    .B1(_02942_));
 sg13g2_nor2_1 _33418_ (.A(_23286_),
    .B(net5125),
    .Y(_02946_));
 sg13g2_a21oi_1 _33419_ (.A1(_23457_),
    .A2(net5080),
    .Y(_02947_),
    .B1(_02946_));
 sg13g2_a221oi_1 _33420_ (.B2(net5112),
    .C1(net6410),
    .B1(_23389_),
    .A1(net1561),
    .Y(_02948_),
    .A2(net7031));
 sg13g2_a22oi_1 _33421_ (.Y(_00621_),
    .B1(_02947_),
    .B2(_02948_),
    .A2(net6410),
    .A1(_18019_));
 sg13g2_nor2_1 _33422_ (.A(_23286_),
    .B(net5070),
    .Y(_02949_));
 sg13g2_a221oi_1 _33423_ (.B2(net5139),
    .C1(net6410),
    .B1(_23418_),
    .A1(net1454),
    .Y(_02950_),
    .A2(net7031));
 sg13g2_a21oi_1 _33424_ (.A1(_23457_),
    .A2(net5112),
    .Y(_02951_),
    .B1(_02949_));
 sg13g2_a22oi_1 _33425_ (.Y(_00622_),
    .B1(_02950_),
    .B2(_02951_),
    .A2(net6410),
    .A1(_18018_));
 sg13g2_a22oi_1 _33426_ (.Y(_02952_),
    .B1(net5892),
    .B2(_23418_),
    .A2(net5946),
    .A1(_23645_));
 sg13g2_o21ai_1 _33427_ (.B1(_02952_),
    .Y(_02953_),
    .A1(_23286_),
    .A2(net6004));
 sg13g2_a221oi_1 _33428_ (.B2(_02953_),
    .C1(net6410),
    .B1(net5237),
    .A1(\u_inv.input_reg[163] ),
    .Y(_02954_),
    .A2(net7031));
 sg13g2_a21oi_1 _33429_ (.A1(_18017_),
    .A2(net6410),
    .Y(_00623_),
    .B1(_02954_));
 sg13g2_nor2_1 _33430_ (.A(net3457),
    .B(net6487),
    .Y(_02955_));
 sg13g2_a22oi_1 _33431_ (.Y(_02956_),
    .B1(net5896),
    .B2(_23645_),
    .A2(net5977),
    .A1(_23418_));
 sg13g2_nor2_1 _33432_ (.A(net7029),
    .B(_02956_),
    .Y(_02957_));
 sg13g2_a221oi_1 _33433_ (.B2(net5138),
    .C1(_02957_),
    .B1(_22114_),
    .A1(net1980),
    .Y(_02958_),
    .A2(net7030));
 sg13g2_a21oi_1 _33434_ (.A1(net6487),
    .A2(_02958_),
    .Y(_00624_),
    .B1(_02955_));
 sg13g2_nand2_1 _33435_ (.Y(_02959_),
    .A(net1511),
    .B(net6402));
 sg13g2_o21ai_1 _33436_ (.B1(net7096),
    .Y(_02960_),
    .A1(_23620_),
    .A2(net5923));
 sg13g2_a221oi_1 _33437_ (.B2(_22114_),
    .C1(_02960_),
    .B1(net5203),
    .A1(_23645_),
    .Y(_02961_),
    .A2(net5158));
 sg13g2_o21ai_1 _33438_ (.B1(net6488),
    .Y(_02962_),
    .A1(\u_inv.input_reg[165] ),
    .A2(net7096));
 sg13g2_o21ai_1 _33439_ (.B1(_02959_),
    .Y(_00625_),
    .A1(_02961_),
    .A2(_02962_));
 sg13g2_nand2b_1 _33440_ (.Y(_02963_),
    .B(net6487),
    .A_N(net1356));
 sg13g2_a22oi_1 _33441_ (.Y(_02964_),
    .B1(_02963_),
    .B2(net6844),
    .A2(net5138),
    .A1(_23609_));
 sg13g2_nor2_1 _33442_ (.A(_23620_),
    .B(net5070),
    .Y(_02965_));
 sg13g2_a21oi_1 _33443_ (.A1(_22114_),
    .A2(net5112),
    .Y(_02966_),
    .B1(_02965_));
 sg13g2_a22oi_1 _33444_ (.Y(_00626_),
    .B1(_02964_),
    .B2(_02966_),
    .A2(net6402),
    .A1(_18015_));
 sg13g2_a21oi_1 _33445_ (.A1(net1516),
    .A2(net7030),
    .Y(_02967_),
    .B1(net6402));
 sg13g2_nand2_1 _33446_ (.Y(_02968_),
    .A(_23609_),
    .B(net5892));
 sg13g2_o21ai_1 _33447_ (.B1(_02968_),
    .Y(_02969_),
    .A1(_23620_),
    .A2(net6004));
 sg13g2_a22oi_1 _33448_ (.Y(_02970_),
    .B1(_02969_),
    .B2(net7096),
    .A2(net5138),
    .A1(_23574_));
 sg13g2_a22oi_1 _33449_ (.Y(_00627_),
    .B1(_02967_),
    .B2(_02970_),
    .A2(net6402),
    .A1(_18014_));
 sg13g2_nand2b_1 _33450_ (.Y(_02971_),
    .B(net5943),
    .A_N(_02177_));
 sg13g2_a221oi_1 _33451_ (.B2(_23574_),
    .C1(net7029),
    .B1(net5892),
    .A1(_23609_),
    .Y(_02972_),
    .A2(net5977));
 sg13g2_o21ai_1 _33452_ (.B1(net6486),
    .Y(_02973_),
    .A1(net2353),
    .A2(net7095));
 sg13g2_a21oi_1 _33453_ (.A1(_02971_),
    .A2(_02972_),
    .Y(_02974_),
    .B1(_02973_));
 sg13g2_a21o_1 _33454_ (.A2(net6402),
    .A1(net3587),
    .B1(_02974_),
    .X(_00628_));
 sg13g2_a22oi_1 _33455_ (.Y(_02975_),
    .B1(net5943),
    .B2(_01937_),
    .A2(net5977),
    .A1(_23574_));
 sg13g2_nor2_1 _33456_ (.A(net7025),
    .B(_02975_),
    .Y(_02976_));
 sg13g2_a21oi_1 _33457_ (.A1(net2639),
    .A2(net7025),
    .Y(_02977_),
    .B1(_02976_));
 sg13g2_o21ai_1 _33458_ (.B1(_02977_),
    .Y(_02978_),
    .A1(_02177_),
    .A2(net5070));
 sg13g2_mux2_1 _33459_ (.A0(net3631),
    .A1(_02978_),
    .S(net6486),
    .X(_00629_));
 sg13g2_nand2_1 _33460_ (.Y(_02979_),
    .A(_23519_),
    .B(net5137));
 sg13g2_a221oi_1 _33461_ (.B2(net5080),
    .C1(net6400),
    .B1(_01937_),
    .A1(net1930),
    .Y(_02980_),
    .A2(net7025));
 sg13g2_nand2_1 _33462_ (.Y(_02981_),
    .A(_02979_),
    .B(_02980_));
 sg13g2_o21ai_1 _33463_ (.B1(_02981_),
    .Y(_02982_),
    .A1(net3708),
    .A2(net6485));
 sg13g2_o21ai_1 _33464_ (.B1(_02982_),
    .Y(_00630_),
    .A1(_02177_),
    .A2(net5066));
 sg13g2_nand2_1 _33465_ (.Y(_02983_),
    .A(net2927),
    .B(net6400));
 sg13g2_o21ai_1 _33466_ (.B1(net7095),
    .Y(_02984_),
    .A1(_22059_),
    .A2(net5923));
 sg13g2_a221oi_1 _33467_ (.B2(_23519_),
    .C1(_02984_),
    .B1(net5203),
    .A1(_01937_),
    .Y(_02985_),
    .A2(net5158));
 sg13g2_o21ai_1 _33468_ (.B1(net6487),
    .Y(_02986_),
    .A1(net1519),
    .A2(net7098));
 sg13g2_o21ai_1 _33469_ (.B1(_02983_),
    .Y(_00631_),
    .A1(_02985_),
    .A2(_02986_));
 sg13g2_and2_1 _33470_ (.A(net1329),
    .B(net7028),
    .X(_02987_));
 sg13g2_a221oi_1 _33471_ (.B2(_22060_),
    .C1(_02987_),
    .B1(net5080),
    .A1(_02044_),
    .Y(_02988_),
    .A2(net5137));
 sg13g2_a22oi_1 _33472_ (.Y(_02989_),
    .B1(_23519_),
    .B2(net5097),
    .A2(net6399),
    .A1(net3710));
 sg13g2_o21ai_1 _33473_ (.B1(_02989_),
    .Y(_00632_),
    .A1(net6399),
    .A2(_02988_));
 sg13g2_a22oi_1 _33474_ (.Y(_02990_),
    .B1(net5891),
    .B2(_02044_),
    .A2(net5943),
    .A1(_23292_));
 sg13g2_o21ai_1 _33475_ (.B1(_02990_),
    .Y(_02991_),
    .A1(_22059_),
    .A2(net6005));
 sg13g2_a221oi_1 _33476_ (.B2(_02991_),
    .C1(net6401),
    .B1(net5237),
    .A1(net1287),
    .Y(_02992_),
    .A2(net7028));
 sg13g2_a21oi_1 _33477_ (.A1(_18012_),
    .A2(net6400),
    .Y(_00633_),
    .B1(_02992_));
 sg13g2_a22oi_1 _33478_ (.Y(_02993_),
    .B1(_23292_),
    .B2(net5080),
    .A2(net7028),
    .A1(net1630));
 sg13g2_o21ai_1 _33479_ (.B1(_02993_),
    .Y(_02994_),
    .A1(_23436_),
    .A2(net5125));
 sg13g2_a22oi_1 _33480_ (.Y(_02995_),
    .B1(_02994_),
    .B2(net6485),
    .A2(net5097),
    .A1(_02044_));
 sg13g2_o21ai_1 _33481_ (.B1(_02995_),
    .Y(_00634_),
    .A1(_18011_),
    .A2(net6485));
 sg13g2_a21oi_1 _33482_ (.A1(net1978),
    .A2(net7028),
    .Y(_02996_),
    .B1(net6401));
 sg13g2_a22oi_1 _33483_ (.Y(_02997_),
    .B1(net5891),
    .B2(_23437_),
    .A2(net5971),
    .A1(_23292_));
 sg13g2_nor2_1 _33484_ (.A(net7024),
    .B(_02997_),
    .Y(_02998_));
 sg13g2_a21oi_1 _33485_ (.A1(_23639_),
    .A2(net5137),
    .Y(_02999_),
    .B1(_02998_));
 sg13g2_a22oi_1 _33486_ (.Y(_00635_),
    .B1(_02996_),
    .B2(_02999_),
    .A2(net6399),
    .A1(_18010_));
 sg13g2_nand2b_1 _33487_ (.Y(_03000_),
    .B(net6485),
    .A_N(net1551));
 sg13g2_a22oi_1 _33488_ (.Y(_03001_),
    .B1(_03000_),
    .B2(net6837),
    .A2(net5079),
    .A1(_23639_));
 sg13g2_a22oi_1 _33489_ (.Y(_03002_),
    .B1(net5111),
    .B2(_23437_),
    .A2(net5137),
    .A1(_22081_));
 sg13g2_a22oi_1 _33490_ (.Y(_00636_),
    .B1(_03001_),
    .B2(_03002_),
    .A2(net6399),
    .A1(_18009_));
 sg13g2_a21oi_1 _33491_ (.A1(net1570),
    .A2(net7024),
    .Y(_03003_),
    .B1(net6399));
 sg13g2_nand2_1 _33492_ (.Y(_03004_),
    .A(_23639_),
    .B(net5971));
 sg13g2_o21ai_1 _33493_ (.B1(_03004_),
    .Y(_03005_),
    .A1(_23627_),
    .A2(net5920));
 sg13g2_a22oi_1 _33494_ (.Y(_03006_),
    .B1(_03005_),
    .B2(net7089),
    .A2(net5079),
    .A1(_22081_));
 sg13g2_a22oi_1 _33495_ (.Y(_00637_),
    .B1(_03003_),
    .B2(_03006_),
    .A2(net6399),
    .A1(_18008_));
 sg13g2_nor2_1 _33496_ (.A(_23627_),
    .B(net5069),
    .Y(_03007_));
 sg13g2_a221oi_1 _33497_ (.B2(net5134),
    .C1(_03007_),
    .B1(_01944_),
    .A1(net1404),
    .Y(_03008_),
    .A2(net7024));
 sg13g2_a22oi_1 _33498_ (.Y(_03009_),
    .B1(_22081_),
    .B2(net5095),
    .A2(net6400),
    .A1(net3695));
 sg13g2_o21ai_1 _33499_ (.B1(_03009_),
    .Y(_00638_),
    .A1(net6399),
    .A2(_03008_));
 sg13g2_nand2_1 _33500_ (.Y(_03010_),
    .A(net2830),
    .B(net6392));
 sg13g2_a21oi_1 _33501_ (.A1(_22009_),
    .A2(net5941),
    .Y(_03011_),
    .B1(net7020));
 sg13g2_o21ai_1 _33502_ (.B1(_03011_),
    .Y(_03012_),
    .A1(_23627_),
    .A2(net5241));
 sg13g2_a21oi_1 _33503_ (.A1(_01944_),
    .A2(net5202),
    .Y(_03013_),
    .B1(_03012_));
 sg13g2_o21ai_1 _33504_ (.B1(net6481),
    .Y(_03014_),
    .A1(net1581),
    .A2(net7089));
 sg13g2_o21ai_1 _33505_ (.B1(_03010_),
    .Y(_00639_),
    .A1(_03013_),
    .A2(_03014_));
 sg13g2_a21oi_1 _33506_ (.A1(net1544),
    .A2(net7022),
    .Y(_03015_),
    .B1(net6392));
 sg13g2_a22oi_1 _33507_ (.Y(_03016_),
    .B1(net5891),
    .B2(_22009_),
    .A2(net5971),
    .A1(_01944_));
 sg13g2_nor2_1 _33508_ (.A(net7020),
    .B(_03016_),
    .Y(_03017_));
 sg13g2_a21oi_1 _33509_ (.A1(_02081_),
    .A2(net5135),
    .Y(_03018_),
    .B1(_03017_));
 sg13g2_a22oi_1 _33510_ (.Y(_00640_),
    .B1(_03015_),
    .B2(_03018_),
    .A2(net6392),
    .A1(_18006_));
 sg13g2_nand2_1 _33511_ (.Y(_03019_),
    .A(net2372),
    .B(net6392));
 sg13g2_o21ai_1 _33512_ (.B1(net7089),
    .Y(_03020_),
    .A1(_23614_),
    .A2(net5920));
 sg13g2_a221oi_1 _33513_ (.B2(_02081_),
    .C1(_03020_),
    .B1(net5202),
    .A1(_22009_),
    .Y(_03021_),
    .A2(net5160));
 sg13g2_o21ai_1 _33514_ (.B1(net6481),
    .Y(_03022_),
    .A1(net1393),
    .A2(net7090));
 sg13g2_o21ai_1 _33515_ (.B1(_03019_),
    .Y(_00641_),
    .A1(_03021_),
    .A2(_03022_));
 sg13g2_a221oi_1 _33516_ (.B2(net5134),
    .C1(net6391),
    .B1(_23587_),
    .A1(net1835),
    .Y(_03023_),
    .A2(net7020));
 sg13g2_o21ai_1 _33517_ (.B1(_03023_),
    .Y(_03024_),
    .A1(_23614_),
    .A2(net5069));
 sg13g2_o21ai_1 _33518_ (.B1(_03024_),
    .Y(_03025_),
    .A1(net3731),
    .A2(net6482));
 sg13g2_o21ai_1 _33519_ (.B1(_03025_),
    .Y(_00642_),
    .A1(_02080_),
    .A2(net5066));
 sg13g2_o21ai_1 _33520_ (.B1(net6840),
    .Y(_03026_),
    .A1(net2289),
    .A2(net6392));
 sg13g2_nor2_1 _33521_ (.A(_23614_),
    .B(_02370_),
    .Y(_03027_));
 sg13g2_a221oi_1 _33522_ (.B2(_23587_),
    .C1(_03027_),
    .B1(net5079),
    .A1(_23554_),
    .Y(_03028_),
    .A2(net5135));
 sg13g2_a22oi_1 _33523_ (.Y(_00643_),
    .B1(_03026_),
    .B2(_03028_),
    .A2(net6392),
    .A1(_18005_));
 sg13g2_nor2_1 _33524_ (.A(_02186_),
    .B(net5124),
    .Y(_03029_));
 sg13g2_o21ai_1 _33525_ (.B1(net6837),
    .Y(_03030_),
    .A1(net1812),
    .A2(net6391));
 sg13g2_a221oi_1 _33526_ (.B2(_23554_),
    .C1(_03029_),
    .B1(net5079),
    .A1(_23587_),
    .Y(_03031_),
    .A2(net5111));
 sg13g2_a22oi_1 _33527_ (.Y(_00644_),
    .B1(_03030_),
    .B2(_03031_),
    .A2(net6391),
    .A1(_18004_));
 sg13g2_a221oi_1 _33528_ (.B2(net5111),
    .C1(net6391),
    .B1(_23554_),
    .A1(net1817),
    .Y(_03032_),
    .A2(net7021));
 sg13g2_nor2_1 _33529_ (.A(_02186_),
    .B(net5069),
    .Y(_03033_));
 sg13g2_a21oi_1 _33530_ (.A1(_23580_),
    .A2(net5134),
    .Y(_03034_),
    .B1(_03033_));
 sg13g2_a22oi_1 _33531_ (.Y(_00645_),
    .B1(_03032_),
    .B2(_03034_),
    .A2(net6391),
    .A1(_18003_));
 sg13g2_nand2_1 _33532_ (.Y(_03035_),
    .A(_21988_),
    .B(net5134));
 sg13g2_nand2_1 _33533_ (.Y(_03036_),
    .A(_23580_),
    .B(net5886));
 sg13g2_o21ai_1 _33534_ (.B1(_03036_),
    .Y(_03037_),
    .A1(_02186_),
    .A2(net6005));
 sg13g2_a221oi_1 _33535_ (.B2(_03037_),
    .C1(net6391),
    .B1(net5236),
    .A1(net2059),
    .Y(_03038_),
    .A2(net7021));
 sg13g2_a22oi_1 _33536_ (.Y(_00646_),
    .B1(_03035_),
    .B2(_03038_),
    .A2(net6391),
    .A1(_18002_));
 sg13g2_a22oi_1 _33537_ (.Y(_03039_),
    .B1(net5079),
    .B2(_21988_),
    .A2(net5111),
    .A1(_23580_));
 sg13g2_a221oi_1 _33538_ (.B2(net5134),
    .C1(net6390),
    .B1(_02127_),
    .A1(net2312),
    .Y(_03040_),
    .A2(net7017));
 sg13g2_a22oi_1 _33539_ (.Y(_00647_),
    .B1(_03039_),
    .B2(_03040_),
    .A2(net6388),
    .A1(_18001_));
 sg13g2_nand2_1 _33540_ (.Y(_03041_),
    .A(_02127_),
    .B(net5079));
 sg13g2_a22oi_1 _33541_ (.Y(_03042_),
    .B1(net5941),
    .B2(_02237_),
    .A2(net5970),
    .A1(_21988_));
 sg13g2_inv_1 _33542_ (.Y(_03043_),
    .A(_03042_));
 sg13g2_a221oi_1 _33543_ (.B2(_03043_),
    .C1(net6389),
    .B1(net5236),
    .A1(net1872),
    .Y(_03044_),
    .A2(net7022));
 sg13g2_a22oi_1 _33544_ (.Y(_00648_),
    .B1(_03041_),
    .B2(_03044_),
    .A2(net6388),
    .A1(_18000_));
 sg13g2_a22oi_1 _33545_ (.Y(_03045_),
    .B1(net5886),
    .B2(_02237_),
    .A2(net5970),
    .A1(_02127_));
 sg13g2_inv_1 _33546_ (.Y(_03046_),
    .A(_03045_));
 sg13g2_a221oi_1 _33547_ (.B2(_03046_),
    .C1(net6388),
    .B1(net5236),
    .A1(net2382),
    .Y(_03047_),
    .A2(net7017));
 sg13g2_o21ai_1 _33548_ (.B1(_03047_),
    .Y(_03048_),
    .A1(_23495_),
    .A2(net5124));
 sg13g2_o21ai_1 _33549_ (.B1(_03048_),
    .Y(_03049_),
    .A1(net3638),
    .A2(net6481));
 sg13g2_inv_1 _33550_ (.Y(_00649_),
    .A(_03049_));
 sg13g2_nor2_1 _33551_ (.A(_23495_),
    .B(net5069),
    .Y(_03050_));
 sg13g2_a221oi_1 _33552_ (.B2(net5134),
    .C1(_03050_),
    .B1(_01919_),
    .A1(net1999),
    .Y(_03051_),
    .A2(net7018));
 sg13g2_a22oi_1 _33553_ (.Y(_03052_),
    .B1(_02237_),
    .B2(net5095),
    .A2(net6389),
    .A1(net3700));
 sg13g2_o21ai_1 _33554_ (.B1(_03052_),
    .Y(_00650_),
    .A1(net6389),
    .A2(_03051_));
 sg13g2_nand2_1 _33555_ (.Y(_03053_),
    .A(net3355),
    .B(net6389));
 sg13g2_a21oi_1 _33556_ (.A1(_23544_),
    .A2(net5937),
    .Y(_03054_),
    .B1(net7019));
 sg13g2_o21ai_1 _33557_ (.B1(_03054_),
    .Y(_03055_),
    .A1(_23495_),
    .A2(net5240));
 sg13g2_a21oi_1 _33558_ (.A1(_01919_),
    .A2(net5197),
    .Y(_03056_),
    .B1(_03055_));
 sg13g2_o21ai_1 _33559_ (.B1(net6481),
    .Y(_03057_),
    .A1(net1462),
    .A2(net7088));
 sg13g2_o21ai_1 _33560_ (.B1(_03053_),
    .Y(_00651_),
    .A1(_03056_),
    .A2(_03057_));
 sg13g2_nand2b_1 _33561_ (.Y(_03058_),
    .B(net6481),
    .A_N(net1282));
 sg13g2_a22oi_1 _33562_ (.Y(_03059_),
    .B1(_03058_),
    .B2(net6836),
    .A2(net5078),
    .A1(_23544_));
 sg13g2_a22oi_1 _33563_ (.Y(_03060_),
    .B1(net5110),
    .B2(_01919_),
    .A2(net5130),
    .A1(_02115_));
 sg13g2_a22oi_1 _33564_ (.Y(_00652_),
    .B1(_03059_),
    .B2(_03060_),
    .A2(net6389),
    .A1(_17997_));
 sg13g2_a221oi_1 _33565_ (.B2(net5130),
    .C1(net6380),
    .B1(_01931_),
    .A1(net1806),
    .Y(_03061_),
    .A2(net7019));
 sg13g2_a22oi_1 _33566_ (.Y(_03062_),
    .B1(net5078),
    .B2(_02115_),
    .A2(net5110),
    .A1(_23544_));
 sg13g2_a22oi_1 _33567_ (.Y(_00653_),
    .B1(_03061_),
    .B2(_03062_),
    .A2(net6380),
    .A1(_17996_));
 sg13g2_nor2_1 _33568_ (.A(_22128_),
    .B(net5124),
    .Y(_03063_));
 sg13g2_a221oi_1 _33569_ (.B2(net5078),
    .C1(_03063_),
    .B1(_01931_),
    .A1(net1713),
    .Y(_03064_),
    .A2(net7005));
 sg13g2_a22oi_1 _33570_ (.Y(_03065_),
    .B1(_02115_),
    .B2(net5093),
    .A2(net6380),
    .A1(net3707));
 sg13g2_o21ai_1 _33571_ (.B1(_03065_),
    .Y(_00654_),
    .A1(net6380),
    .A2(_03064_));
 sg13g2_a22oi_1 _33572_ (.Y(_03066_),
    .B1(_02139_),
    .B2(net5130),
    .A2(net7004),
    .A1(net1783));
 sg13g2_o21ai_1 _33573_ (.B1(_03066_),
    .Y(_03067_),
    .A1(_22128_),
    .A2(net5069));
 sg13g2_a22oi_1 _33574_ (.Y(_03068_),
    .B1(_03067_),
    .B2(net6477),
    .A2(net5093),
    .A1(_01931_));
 sg13g2_o21ai_1 _33575_ (.B1(_03068_),
    .Y(_00655_),
    .A1(_17995_),
    .A2(net6477));
 sg13g2_o21ai_1 _33576_ (.B1(net6836),
    .Y(_03069_),
    .A1(net1704),
    .A2(net6380));
 sg13g2_o21ai_1 _33577_ (.B1(_03069_),
    .Y(_03070_),
    .A1(_22128_),
    .A2(_02370_));
 sg13g2_a221oi_1 _33578_ (.B2(_02139_),
    .C1(_03070_),
    .B1(net5078),
    .A1(_02216_),
    .Y(_03071_),
    .A2(net5130));
 sg13g2_a21oi_1 _33579_ (.A1(_17994_),
    .A2(net6380),
    .Y(_00656_),
    .B1(_03071_));
 sg13g2_a221oi_1 _33580_ (.B2(net5110),
    .C1(net6380),
    .B1(_02139_),
    .A1(net1833),
    .Y(_03072_),
    .A2(net7004));
 sg13g2_a22oi_1 _33581_ (.Y(_03073_),
    .B1(net5078),
    .B2(_02216_),
    .A2(net5130),
    .A1(_23601_));
 sg13g2_a22oi_1 _33582_ (.Y(_00657_),
    .B1(_03072_),
    .B2(_03073_),
    .A2(net6381),
    .A1(_17993_));
 sg13g2_a22oi_1 _33583_ (.Y(_03074_),
    .B1(net5884),
    .B2(_23601_),
    .A2(net5935),
    .A1(_22036_));
 sg13g2_a221oi_1 _33584_ (.B2(net5110),
    .C1(net6380),
    .B1(_02216_),
    .A1(net1456),
    .Y(_03075_),
    .A2(net7004));
 sg13g2_o21ai_1 _33585_ (.B1(_03075_),
    .Y(_03076_),
    .A1(net7005),
    .A2(_03074_));
 sg13g2_o21ai_1 _33586_ (.B1(_03076_),
    .Y(_03077_),
    .A1(net3531),
    .A2(net6477));
 sg13g2_inv_1 _33587_ (.Y(_00658_),
    .A(_03077_));
 sg13g2_nand2_1 _33588_ (.Y(_03078_),
    .A(net2380),
    .B(net6379));
 sg13g2_o21ai_1 _33589_ (.B1(net7080),
    .Y(_03079_),
    .A1(_02169_),
    .A2(net5918));
 sg13g2_a221oi_1 _33590_ (.B2(_22036_),
    .C1(_03079_),
    .B1(net5195),
    .A1(_23601_),
    .Y(_03080_),
    .A2(net5154));
 sg13g2_o21ai_1 _33591_ (.B1(net6477),
    .Y(_03081_),
    .A1(net1425),
    .A2(net7081));
 sg13g2_o21ai_1 _33592_ (.B1(_03078_),
    .Y(_00659_),
    .A1(_03080_),
    .A2(_03081_));
 sg13g2_nor2_1 _33593_ (.A(_02169_),
    .B(net5067),
    .Y(_03082_));
 sg13g2_a221oi_1 _33594_ (.B2(net5129),
    .C1(_03082_),
    .B1(_02262_),
    .A1(net1340),
    .Y(_03083_),
    .A2(net7003));
 sg13g2_a22oi_1 _33595_ (.Y(_03084_),
    .B1(_22036_),
    .B2(net5092),
    .A2(net6379),
    .A1(net3699));
 sg13g2_o21ai_1 _33596_ (.B1(_03084_),
    .Y(_00660_),
    .A1(net6381),
    .A2(_03083_));
 sg13g2_nor2_1 _33597_ (.A(_23534_),
    .B(net5918),
    .Y(_03085_));
 sg13g2_a21oi_1 _33598_ (.A1(_02262_),
    .A2(net5884),
    .Y(_03086_),
    .B1(_03085_));
 sg13g2_o21ai_1 _33599_ (.B1(_03086_),
    .Y(_03087_),
    .A1(_02169_),
    .A2(net6003));
 sg13g2_a221oi_1 _33600_ (.B2(_03087_),
    .C1(net6379),
    .B1(net5235),
    .A1(net2759),
    .Y(_03088_),
    .A2(net7003));
 sg13g2_a21oi_1 _33601_ (.A1(_17991_),
    .A2(net6381),
    .Y(_00661_),
    .B1(_03088_));
 sg13g2_o21ai_1 _33602_ (.B1(net6836),
    .Y(_03089_),
    .A1(net1660),
    .A2(net6379));
 sg13g2_o21ai_1 _33603_ (.B1(_03089_),
    .Y(_03090_),
    .A1(_23534_),
    .A2(net5067));
 sg13g2_a221oi_1 _33604_ (.B2(_02262_),
    .C1(_03090_),
    .B1(net5110),
    .A1(_23527_),
    .Y(_03091_),
    .A2(net5129));
 sg13g2_a21oi_1 _33605_ (.A1(_17990_),
    .A2(net6379),
    .Y(_00662_),
    .B1(_03091_));
 sg13g2_nand2_1 _33606_ (.Y(_03092_),
    .A(net3419),
    .B(net6379));
 sg13g2_o21ai_1 _33607_ (.B1(net7080),
    .Y(_03093_),
    .A1(_23534_),
    .A2(net5239));
 sg13g2_a221oi_1 _33608_ (.B2(_23527_),
    .C1(_03093_),
    .B1(net5195),
    .A1(_21960_),
    .Y(_03094_),
    .A2(net5935));
 sg13g2_o21ai_1 _33609_ (.B1(net6481),
    .Y(_03095_),
    .A1(net2785),
    .A2(net7081));
 sg13g2_o21ai_1 _33610_ (.B1(_03092_),
    .Y(_00663_),
    .A1(_03094_),
    .A2(_03095_));
 sg13g2_nor2_1 _33611_ (.A(_21932_),
    .B(net5123),
    .Y(_03096_));
 sg13g2_a221oi_1 _33612_ (.B2(net5077),
    .C1(_03096_),
    .B1(_21960_),
    .A1(net2484),
    .Y(_03097_),
    .A2(net6996));
 sg13g2_a22oi_1 _33613_ (.Y(_03098_),
    .B1(_23527_),
    .B2(net5092),
    .A2(net6372),
    .A1(net3736));
 sg13g2_o21ai_1 _33614_ (.B1(_03098_),
    .Y(_00664_),
    .A1(net6372),
    .A2(_03097_));
 sg13g2_nand2_1 _33615_ (.Y(_03099_),
    .A(net1926),
    .B(net6372));
 sg13g2_a22oi_1 _33616_ (.Y(_03100_),
    .B1(net5195),
    .B2(_21933_),
    .A2(net5935),
    .A1(_01925_));
 sg13g2_nand2_1 _33617_ (.Y(_03101_),
    .A(net7078),
    .B(_03100_));
 sg13g2_a21oi_1 _33618_ (.A1(_21960_),
    .A2(net5154),
    .Y(_03102_),
    .B1(_03101_));
 sg13g2_o21ai_1 _33619_ (.B1(net6477),
    .Y(_03103_),
    .A1(\u_inv.input_reg[205] ),
    .A2(net7080));
 sg13g2_o21ai_1 _33620_ (.B1(_03099_),
    .Y(_00665_),
    .A1(_03102_),
    .A2(_03103_));
 sg13g2_and2_1 _33621_ (.A(net1928),
    .B(net6996),
    .X(_03104_));
 sg13g2_a221oi_1 _33622_ (.B2(_01925_),
    .C1(_03104_),
    .B1(net5077),
    .A1(_22019_),
    .Y(_03105_),
    .A2(net5129));
 sg13g2_a22oi_1 _33623_ (.Y(_03106_),
    .B1(_21933_),
    .B2(net5092),
    .A2(net6372),
    .A1(net3711));
 sg13g2_o21ai_1 _33624_ (.B1(_03106_),
    .Y(_00666_),
    .A1(net6372),
    .A2(_03105_));
 sg13g2_nand2_1 _33625_ (.Y(_03107_),
    .A(net2843),
    .B(net6372));
 sg13g2_o21ai_1 _33626_ (.B1(net7078),
    .Y(_03108_),
    .A1(_02198_),
    .A2(net5918));
 sg13g2_a221oi_1 _33627_ (.B2(_22019_),
    .C1(_03108_),
    .B1(net5195),
    .A1(_01925_),
    .Y(_03109_),
    .A2(net5154));
 sg13g2_o21ai_1 _33628_ (.B1(net6477),
    .Y(_03110_),
    .A1(net2718),
    .A2(net7078));
 sg13g2_o21ai_1 _33629_ (.B1(_03107_),
    .Y(_00667_),
    .A1(_03109_),
    .A2(_03110_));
 sg13g2_nand2b_1 _33630_ (.Y(_03111_),
    .B(net6475),
    .A_N(net1481));
 sg13g2_a22oi_1 _33631_ (.Y(_03112_),
    .B1(_03111_),
    .B2(net6836),
    .A2(net5077),
    .A1(_02199_));
 sg13g2_a22oi_1 _33632_ (.Y(_03113_),
    .B1(net5110),
    .B2(_22019_),
    .A2(net5129),
    .A1(_01981_));
 sg13g2_a22oi_1 _33633_ (.Y(_00668_),
    .B1(_03112_),
    .B2(_03113_),
    .A2(net6372),
    .A1(_17986_));
 sg13g2_nand2_1 _33634_ (.Y(_03114_),
    .A(net2756),
    .B(net6372));
 sg13g2_o21ai_1 _33635_ (.B1(net7078),
    .Y(_03115_),
    .A1(_22141_),
    .A2(net5918));
 sg13g2_a221oi_1 _33636_ (.B2(_01981_),
    .C1(_03115_),
    .B1(net5195),
    .A1(_02199_),
    .Y(_03116_),
    .A2(net5154));
 sg13g2_o21ai_1 _33637_ (.B1(net6477),
    .Y(_03117_),
    .A1(net2301),
    .A2(net7078));
 sg13g2_o21ai_1 _33638_ (.B1(_03114_),
    .Y(_00669_),
    .A1(_03116_),
    .A2(_03117_));
 sg13g2_nor2_1 _33639_ (.A(_22150_),
    .B(net5123),
    .Y(_03118_));
 sg13g2_nand2_1 _33640_ (.Y(_03119_),
    .A(net1528),
    .B(net7003));
 sg13g2_o21ai_1 _33641_ (.B1(_03119_),
    .Y(_03120_),
    .A1(_22141_),
    .A2(net5067));
 sg13g2_o21ai_1 _33642_ (.B1(net6475),
    .Y(_03121_),
    .A1(_03118_),
    .A2(_03120_));
 sg13g2_a22oi_1 _33643_ (.Y(_03122_),
    .B1(_01981_),
    .B2(net5092),
    .A2(net6373),
    .A1(net3721));
 sg13g2_nand2_1 _33644_ (.Y(_00670_),
    .A(_03121_),
    .B(_03122_));
 sg13g2_nor2_1 _33645_ (.A(_22150_),
    .B(net5122),
    .Y(_03123_));
 sg13g2_a21oi_1 _33646_ (.A1(_02192_),
    .A2(net5935),
    .Y(_03124_),
    .B1(net6996));
 sg13g2_o21ai_1 _33647_ (.B1(_03124_),
    .Y(_03125_),
    .A1(_22141_),
    .A2(net5239));
 sg13g2_a21oi_1 _33648_ (.A1(_18614_),
    .A2(net7003),
    .Y(_03126_),
    .B1(net6379));
 sg13g2_o21ai_1 _33649_ (.B1(_03126_),
    .Y(_03127_),
    .A1(_03123_),
    .A2(_03125_));
 sg13g2_o21ai_1 _33650_ (.B1(_03127_),
    .Y(_00671_),
    .A1(_17985_),
    .A2(net6475));
 sg13g2_a22oi_1 _33651_ (.Y(_03128_),
    .B1(net5884),
    .B2(_02192_),
    .A2(net5935),
    .A1(_01998_));
 sg13g2_o21ai_1 _33652_ (.B1(_03128_),
    .Y(_03129_),
    .A1(_22150_),
    .A2(net6003));
 sg13g2_a221oi_1 _33653_ (.B2(_03129_),
    .C1(net6373),
    .B1(net5235),
    .A1(net1699),
    .Y(_03130_),
    .A2(net7003));
 sg13g2_a21oi_1 _33654_ (.A1(_17984_),
    .A2(net6374),
    .Y(_00672_),
    .B1(_03130_));
 sg13g2_nand2_1 _33655_ (.Y(_03131_),
    .A(net3326),
    .B(net6373));
 sg13g2_o21ai_1 _33656_ (.B1(net7078),
    .Y(_03132_),
    .A1(_21997_),
    .A2(net5918));
 sg13g2_a221oi_1 _33657_ (.B2(_01998_),
    .C1(_03132_),
    .B1(net5195),
    .A1(_02192_),
    .Y(_03133_),
    .A2(net5154));
 sg13g2_o21ai_1 _33658_ (.B1(net6477),
    .Y(_03134_),
    .A1(net2457),
    .A2(net7078));
 sg13g2_o21ai_1 _33659_ (.B1(_03131_),
    .Y(_00673_),
    .A1(_03133_),
    .A2(_03134_));
 sg13g2_nor2_1 _33660_ (.A(_02146_),
    .B(net5123),
    .Y(_03135_));
 sg13g2_a221oi_1 _33661_ (.B2(net5077),
    .C1(_03135_),
    .B1(_21998_),
    .A1(net2272),
    .Y(_03136_),
    .A2(net6996));
 sg13g2_a22oi_1 _33662_ (.Y(_03137_),
    .B1(_01998_),
    .B2(net5092),
    .A2(net6374),
    .A1(net3725));
 sg13g2_o21ai_1 _33663_ (.B1(_03137_),
    .Y(_00674_),
    .A1(net6374),
    .A2(_03136_));
 sg13g2_a22oi_1 _33664_ (.Y(_03138_),
    .B1(_01987_),
    .B2(net5129),
    .A2(net7006),
    .A1(net1628));
 sg13g2_o21ai_1 _33665_ (.B1(_03138_),
    .Y(_03139_),
    .A1(_02146_),
    .A2(net5067));
 sg13g2_a22oi_1 _33666_ (.Y(_03140_),
    .B1(_03139_),
    .B2(net6475),
    .A2(net5092),
    .A1(_21998_));
 sg13g2_o21ai_1 _33667_ (.B1(_03140_),
    .Y(_00675_),
    .A1(_17982_),
    .A2(net6475));
 sg13g2_nand2_1 _33668_ (.Y(_03141_),
    .A(net2052),
    .B(net6379));
 sg13g2_o21ai_1 _33669_ (.B1(net7078),
    .Y(_03142_),
    .A1(_02146_),
    .A2(net6003));
 sg13g2_a221oi_1 _33670_ (.B2(_01987_),
    .C1(_03142_),
    .B1(net5884),
    .A1(_21831_),
    .Y(_03143_),
    .A2(net5935));
 sg13g2_o21ai_1 _33671_ (.B1(net6478),
    .Y(_03144_),
    .A1(net1625),
    .A2(net7080));
 sg13g2_o21ai_1 _33672_ (.B1(_03141_),
    .Y(_00676_),
    .A1(_03143_),
    .A2(_03144_));
 sg13g2_a22oi_1 _33673_ (.Y(_03145_),
    .B1(net5936),
    .B2(_02162_),
    .A2(net5976),
    .A1(_01987_));
 sg13g2_o21ai_1 _33674_ (.B1(_03145_),
    .Y(_03146_),
    .A1(_21830_),
    .A2(net5122));
 sg13g2_nand2_1 _33675_ (.Y(_03147_),
    .A(net7079),
    .B(_03146_));
 sg13g2_a21oi_1 _33676_ (.A1(net1310),
    .A2(net7006),
    .Y(_03148_),
    .B1(net6382));
 sg13g2_a22oi_1 _33677_ (.Y(_00677_),
    .B1(_03147_),
    .B2(_03148_),
    .A2(net6373),
    .A1(_17980_));
 sg13g2_nand2_1 _33678_ (.Y(_03149_),
    .A(net2937),
    .B(net6375));
 sg13g2_a22oi_1 _33679_ (.Y(_03150_),
    .B1(net5196),
    .B2(_02162_),
    .A2(net5936),
    .A1(_02155_));
 sg13g2_nand2_1 _33680_ (.Y(_03151_),
    .A(net7079),
    .B(_03150_));
 sg13g2_a21oi_1 _33681_ (.A1(_21831_),
    .A2(net5154),
    .Y(_03152_),
    .B1(_03151_));
 sg13g2_o21ai_1 _33682_ (.B1(net6475),
    .Y(_03153_),
    .A1(net1469),
    .A2(net7080));
 sg13g2_o21ai_1 _33683_ (.B1(_03149_),
    .Y(_00678_),
    .A1(_03152_),
    .A2(_03153_));
 sg13g2_nand2_1 _33684_ (.Y(_03154_),
    .A(net1726),
    .B(net6377));
 sg13g2_a21o_1 _33685_ (.A2(net5935),
    .A1(_02222_),
    .B1(net7000),
    .X(_03155_));
 sg13g2_a221oi_1 _33686_ (.B2(_02155_),
    .C1(_03155_),
    .B1(net5195),
    .A1(_02162_),
    .Y(_03156_),
    .A2(net5155));
 sg13g2_o21ai_1 _33687_ (.B1(net6475),
    .Y(_03157_),
    .A1(\u_inv.input_reg[219] ),
    .A2(net7079));
 sg13g2_o21ai_1 _33688_ (.B1(_03154_),
    .Y(_00679_),
    .A1(_03156_),
    .A2(_03157_));
 sg13g2_nand2_1 _33689_ (.Y(_03158_),
    .A(_01972_),
    .B(net5223));
 sg13g2_o21ai_1 _33690_ (.B1(_03158_),
    .Y(_03159_),
    .A1(_02155_),
    .A2(net5239));
 sg13g2_o21ai_1 _33691_ (.B1(net7079),
    .Y(_03160_),
    .A1(_02222_),
    .A2(net5122));
 sg13g2_or2_1 _33692_ (.X(_03161_),
    .B(_03160_),
    .A(_03159_));
 sg13g2_a21oi_1 _33693_ (.A1(net1312),
    .A2(net7006),
    .Y(_03162_),
    .B1(net6382));
 sg13g2_a22oi_1 _33694_ (.Y(_00680_),
    .B1(_03161_),
    .B2(_03162_),
    .A2(net6375),
    .A1(_17978_));
 sg13g2_nor2_1 _33695_ (.A(_01972_),
    .B(net5067),
    .Y(_03163_));
 sg13g2_a221oi_1 _33696_ (.B2(net5129),
    .C1(_03163_),
    .B1(_23594_),
    .A1(net1868),
    .Y(_03164_),
    .A2(net7000));
 sg13g2_a22oi_1 _33697_ (.Y(_03165_),
    .B1(_02222_),
    .B2(net5092),
    .A2(net6375),
    .A1(net3702));
 sg13g2_o21ai_1 _33698_ (.B1(_03165_),
    .Y(_00681_),
    .A1(net6375),
    .A2(_03164_));
 sg13g2_nand2_1 _33699_ (.Y(_03166_),
    .A(_23594_),
    .B(net5195));
 sg13g2_o21ai_1 _33700_ (.B1(_03166_),
    .Y(_03167_),
    .A1(_01972_),
    .A2(net5239));
 sg13g2_a22oi_1 _33701_ (.Y(_03168_),
    .B1(_01904_),
    .B2(net5129),
    .A2(net7006),
    .A1(net1795));
 sg13g2_a22oi_1 _33702_ (.Y(_03169_),
    .B1(net6866),
    .B2(_03167_),
    .A2(net6375),
    .A1(net3609));
 sg13g2_o21ai_1 _33703_ (.B1(_03169_),
    .Y(_00682_),
    .A1(net6375),
    .A2(_03168_));
 sg13g2_a21oi_1 _33704_ (.A1(net2673),
    .A2(net7001),
    .Y(_03170_),
    .B1(net6375));
 sg13g2_a22oi_1 _33705_ (.Y(_03171_),
    .B1(net5884),
    .B2(_01904_),
    .A2(net5976),
    .A1(_23594_));
 sg13g2_nor2_1 _33706_ (.A(net7000),
    .B(_03171_),
    .Y(_03172_));
 sg13g2_a21oi_1 _33707_ (.A1(_22092_),
    .A2(net5129),
    .Y(_03173_),
    .B1(_03172_));
 sg13g2_a22oi_1 _33708_ (.Y(_00683_),
    .B1(_03170_),
    .B2(_03173_),
    .A2(net6378),
    .A1(_17977_));
 sg13g2_nand2_1 _33709_ (.Y(_03174_),
    .A(net2498),
    .B(net6377));
 sg13g2_a21oi_1 _33710_ (.A1(_02026_),
    .A2(net5936),
    .Y(_03175_),
    .B1(net7000));
 sg13g2_o21ai_1 _33711_ (.B1(_03175_),
    .Y(_03176_),
    .A1(_01903_),
    .A2(net5239));
 sg13g2_a21oi_1 _33712_ (.A1(_22092_),
    .A2(net5196),
    .Y(_03177_),
    .B1(_03176_));
 sg13g2_o21ai_1 _33713_ (.B1(net6476),
    .Y(_03178_),
    .A1(net1399),
    .A2(net7079));
 sg13g2_o21ai_1 _33714_ (.B1(_03174_),
    .Y(_00684_),
    .A1(_03177_),
    .A2(_03178_));
 sg13g2_a22oi_1 _33715_ (.Y(_03179_),
    .B1(net5885),
    .B2(_02026_),
    .A2(net5976),
    .A1(_22092_));
 sg13g2_inv_1 _33716_ (.Y(_03180_),
    .A(_03179_));
 sg13g2_a221oi_1 _33717_ (.B2(_03180_),
    .C1(net6375),
    .B1(net5235),
    .A1(net1838),
    .Y(_03181_),
    .A2(net7000));
 sg13g2_o21ai_1 _33718_ (.B1(_03181_),
    .Y(_03182_),
    .A1(_21971_),
    .A2(net5123));
 sg13g2_o21ai_1 _33719_ (.B1(_03182_),
    .Y(_03183_),
    .A1(net3752),
    .A2(net6476));
 sg13g2_inv_1 _33720_ (.Y(_00685_),
    .A(_03183_));
 sg13g2_nand2b_1 _33721_ (.Y(_03184_),
    .B(net5196),
    .A_N(_21971_));
 sg13g2_a221oi_1 _33722_ (.B2(_22101_),
    .C1(net7001),
    .B1(net5936),
    .A1(_02026_),
    .Y(_03185_),
    .A2(net5154));
 sg13g2_o21ai_1 _33723_ (.B1(net6476),
    .Y(_03186_),
    .A1(net1395),
    .A2(net7079));
 sg13g2_a21oi_1 _33724_ (.A1(_03184_),
    .A2(_03185_),
    .Y(_03187_),
    .B1(_03186_));
 sg13g2_a21o_1 _33725_ (.A2(net6376),
    .A1(net3369),
    .B1(_03187_),
    .X(_00686_));
 sg13g2_nand2_1 _33726_ (.Y(_03188_),
    .A(net2947),
    .B(net6377));
 sg13g2_a21oi_1 _33727_ (.A1(_02036_),
    .A2(net5936),
    .Y(_03189_),
    .B1(net7001));
 sg13g2_o21ai_1 _33728_ (.B1(_03189_),
    .Y(_03190_),
    .A1(_21971_),
    .A2(net5239));
 sg13g2_a21oi_1 _33729_ (.A1(_22101_),
    .A2(net5196),
    .Y(_03191_),
    .B1(_03190_));
 sg13g2_o21ai_1 _33730_ (.B1(net6475),
    .Y(_03192_),
    .A1(net1652),
    .A2(net7079));
 sg13g2_o21ai_1 _33731_ (.B1(_03188_),
    .Y(_00687_),
    .A1(_03191_),
    .A2(_03192_));
 sg13g2_and2_1 _33732_ (.A(net1559),
    .B(net7001),
    .X(_03193_));
 sg13g2_a221oi_1 _33733_ (.B2(_02036_),
    .C1(_03193_),
    .B1(net5075),
    .A1(_02254_),
    .Y(_03194_),
    .A2(net5131));
 sg13g2_a22oi_1 _33734_ (.Y(_03195_),
    .B1(_22101_),
    .B2(net5092),
    .A2(net6376),
    .A1(net3732));
 sg13g2_o21ai_1 _33735_ (.B1(_03195_),
    .Y(_00688_),
    .A1(net6376),
    .A2(_03194_));
 sg13g2_a221oi_1 _33736_ (.B2(net5075),
    .C1(net6376),
    .B1(_02254_),
    .A1(net1610),
    .Y(_03196_),
    .A2(net7001));
 sg13g2_nor2_1 _33737_ (.A(_22068_),
    .B(net5123),
    .Y(_03197_));
 sg13g2_a21oi_1 _33738_ (.A1(_02036_),
    .A2(net5110),
    .Y(_03198_),
    .B1(_03197_));
 sg13g2_a22oi_1 _33739_ (.Y(_00689_),
    .B1(_03196_),
    .B2(_03198_),
    .A2(net6376),
    .A1(_17974_));
 sg13g2_nor2_1 _33740_ (.A(_22068_),
    .B(net5068),
    .Y(_03199_));
 sg13g2_a221oi_1 _33741_ (.B2(net5131),
    .C1(_03199_),
    .B1(_02088_),
    .A1(net1401),
    .Y(_03200_),
    .A2(net7009));
 sg13g2_a22oi_1 _33742_ (.Y(_03201_),
    .B1(_02254_),
    .B2(net5093),
    .A2(net6378),
    .A1(net3705));
 sg13g2_o21ai_1 _33743_ (.B1(_03201_),
    .Y(_00690_),
    .A1(net6378),
    .A2(_03200_));
 sg13g2_nand2_1 _33744_ (.Y(_03202_),
    .A(net3130),
    .B(net6376));
 sg13g2_a21oi_1 _33745_ (.A1(_02018_),
    .A2(net5935),
    .Y(_03203_),
    .B1(net7009));
 sg13g2_o21ai_1 _33746_ (.B1(_03203_),
    .Y(_03204_),
    .A1(_22068_),
    .A2(net5239));
 sg13g2_a21oi_1 _33747_ (.A1(_02088_),
    .A2(net5196),
    .Y(_03205_),
    .B1(_03204_));
 sg13g2_o21ai_1 _33748_ (.B1(net6476),
    .Y(_03206_),
    .A1(net2093),
    .A2(net7079));
 sg13g2_o21ai_1 _33749_ (.B1(_03202_),
    .Y(_00691_),
    .A1(_03205_),
    .A2(_03206_));
 sg13g2_nand2_1 _33750_ (.Y(_03207_),
    .A(net3195),
    .B(net6376));
 sg13g2_o21ai_1 _33751_ (.B1(net7082),
    .Y(_03208_),
    .A1(_21862_),
    .A2(net5918));
 sg13g2_a221oi_1 _33752_ (.B2(_02018_),
    .C1(_03208_),
    .B1(net5196),
    .A1(_02088_),
    .Y(_03209_),
    .A2(net5154));
 sg13g2_o21ai_1 _33753_ (.B1(net6479),
    .Y(_03210_),
    .A1(net1385),
    .A2(net7082));
 sg13g2_o21ai_1 _33754_ (.B1(_03207_),
    .Y(_00692_),
    .A1(_03209_),
    .A2(_03210_));
 sg13g2_nand2_1 _33755_ (.Y(_03211_),
    .A(net2818),
    .B(net6376));
 sg13g2_a22oi_1 _33756_ (.Y(_03212_),
    .B1(net5198),
    .B2(_21863_),
    .A2(net5938),
    .A1(_21940_));
 sg13g2_nand2_1 _33757_ (.Y(_03213_),
    .A(net7082),
    .B(_03212_));
 sg13g2_a21oi_1 _33758_ (.A1(_02018_),
    .A2(net5155),
    .Y(_03214_),
    .B1(_03213_));
 sg13g2_o21ai_1 _33759_ (.B1(net6480),
    .Y(_03215_),
    .A1(net1377),
    .A2(net7082));
 sg13g2_o21ai_1 _33760_ (.B1(_03211_),
    .Y(_00693_),
    .A1(_03214_),
    .A2(_03215_));
 sg13g2_nor2_1 _33761_ (.A(_02062_),
    .B(net5123),
    .Y(_03216_));
 sg13g2_a221oi_1 _33762_ (.B2(net5075),
    .C1(_03216_),
    .B1(_21940_),
    .A1(net1514),
    .Y(_03217_),
    .A2(net7009));
 sg13g2_a22oi_1 _33763_ (.Y(_03218_),
    .B1(_21863_),
    .B2(net5094),
    .A2(net6384),
    .A1(net3746));
 sg13g2_o21ai_1 _33764_ (.B1(_03218_),
    .Y(_00694_),
    .A1(net6384),
    .A2(_03217_));
 sg13g2_nand2_1 _33765_ (.Y(_03219_),
    .A(net2874),
    .B(net6383));
 sg13g2_o21ai_1 _33766_ (.B1(net7082),
    .Y(_03220_),
    .A1(_01950_),
    .A2(net5919));
 sg13g2_a221oi_1 _33767_ (.B2(_02063_),
    .C1(_03220_),
    .B1(net5198),
    .A1(_21940_),
    .Y(_03221_),
    .A2(net5156));
 sg13g2_o21ai_1 _33768_ (.B1(net6480),
    .Y(_03222_),
    .A1(net1942),
    .A2(net7082));
 sg13g2_o21ai_1 _33769_ (.B1(_03219_),
    .Y(_00695_),
    .A1(_03221_),
    .A2(_03222_));
 sg13g2_o21ai_1 _33770_ (.B1(net6836),
    .Y(_03223_),
    .A1(net1438),
    .A2(net6383));
 sg13g2_a221oi_1 _33771_ (.B2(_01950_),
    .C1(net7009),
    .B1(net5198),
    .A1(_02062_),
    .Y(_03224_),
    .A2(net5156));
 sg13g2_o21ai_1 _33772_ (.B1(_03224_),
    .Y(_03225_),
    .A1(_21881_),
    .A2(net5151));
 sg13g2_a22oi_1 _33773_ (.Y(_00696_),
    .B1(_03223_),
    .B2(_03225_),
    .A2(net6383),
    .A1(_17972_));
 sg13g2_a221oi_1 _33774_ (.B2(net5132),
    .C1(net6383),
    .B1(_22027_),
    .A1(net1289),
    .Y(_03226_),
    .A2(net7009));
 sg13g2_o21ai_1 _33775_ (.B1(_03226_),
    .Y(_03227_),
    .A1(_21880_),
    .A2(net5068));
 sg13g2_o21ai_1 _33776_ (.B1(_03227_),
    .Y(_03228_),
    .A1(net3733),
    .A2(net6479));
 sg13g2_o21ai_1 _33777_ (.B1(_03228_),
    .Y(_00697_),
    .A1(_01950_),
    .A2(net5066));
 sg13g2_a221oi_1 _33778_ (.B2(net5075),
    .C1(net6383),
    .B1(_22027_),
    .A1(net1604),
    .Y(_03229_),
    .A2(net7009));
 sg13g2_o21ai_1 _33779_ (.B1(_03229_),
    .Y(_03230_),
    .A1(_22158_),
    .A2(net5123));
 sg13g2_o21ai_1 _33780_ (.B1(_03230_),
    .Y(_03231_),
    .A1(net3716),
    .A2(net6479));
 sg13g2_o21ai_1 _33781_ (.B1(_03231_),
    .Y(_00698_),
    .A1(_21880_),
    .A2(net5066));
 sg13g2_nor2_1 _33782_ (.A(_22158_),
    .B(net5068),
    .Y(_03232_));
 sg13g2_a221oi_1 _33783_ (.B2(net5132),
    .C1(_03232_),
    .B1(_21953_),
    .A1(net1333),
    .Y(_03233_),
    .A2(net7010));
 sg13g2_a22oi_1 _33784_ (.Y(_03234_),
    .B1(_22027_),
    .B2(net5094),
    .A2(net6383),
    .A1(net3730));
 sg13g2_o21ai_1 _33785_ (.B1(_03234_),
    .Y(_00699_),
    .A1(net6384),
    .A2(_03233_));
 sg13g2_a221oi_1 _33786_ (.B2(net5132),
    .C1(net6383),
    .B1(_01958_),
    .A1(net1327),
    .Y(_03235_),
    .A2(net7009));
 sg13g2_o21ai_1 _33787_ (.B1(_03235_),
    .Y(_03236_),
    .A1(_21952_),
    .A2(net5068));
 sg13g2_o21ai_1 _33788_ (.B1(_03236_),
    .Y(_03237_),
    .A1(net3735),
    .A2(net6479));
 sg13g2_o21ai_1 _33789_ (.B1(_03237_),
    .Y(_00700_),
    .A1(_22158_),
    .A2(net5066));
 sg13g2_nand2_1 _33790_ (.Y(_03238_),
    .A(net3501),
    .B(net6384));
 sg13g2_a22oi_1 _33791_ (.Y(_03239_),
    .B1(net5198),
    .B2(_01958_),
    .A2(net5938),
    .A1(_02105_));
 sg13g2_nand2_1 _33792_ (.Y(_03240_),
    .A(net7083),
    .B(_03239_));
 sg13g2_a21oi_1 _33793_ (.A1(_21953_),
    .A2(net5156),
    .Y(_03241_),
    .B1(_03240_));
 sg13g2_o21ai_1 _33794_ (.B1(net6479),
    .Y(_03242_),
    .A1(net1320),
    .A2(net7082));
 sg13g2_o21ai_1 _33795_ (.B1(_03238_),
    .Y(_00701_),
    .A1(_03241_),
    .A2(_03242_));
 sg13g2_a22oi_1 _33796_ (.Y(_03243_),
    .B1(_02105_),
    .B2(net5075),
    .A2(net7009),
    .A1(net1475));
 sg13g2_o21ai_1 _33797_ (.B1(_03243_),
    .Y(_03244_),
    .A1(_02207_),
    .A2(net5123));
 sg13g2_a22oi_1 _33798_ (.Y(_03245_),
    .B1(_03244_),
    .B2(net6479),
    .A2(net5094),
    .A1(_01958_));
 sg13g2_o21ai_1 _33799_ (.B1(_03245_),
    .Y(_00702_),
    .A1(_17969_),
    .A2(net6479));
 sg13g2_nand2_1 _33800_ (.Y(_03246_),
    .A(net1691),
    .B(net6384));
 sg13g2_o21ai_1 _33801_ (.B1(net7083),
    .Y(_03247_),
    .A1(_02005_),
    .A2(net5919));
 sg13g2_a221oi_1 _33802_ (.B2(_02208_),
    .C1(_03247_),
    .B1(net5198),
    .A1(_02105_),
    .Y(_03248_),
    .A2(net5156));
 sg13g2_o21ai_1 _33803_ (.B1(net6479),
    .Y(_03249_),
    .A1(net1427),
    .A2(net7082));
 sg13g2_o21ai_1 _33804_ (.B1(_03246_),
    .Y(_00703_),
    .A1(_03248_),
    .A2(_03249_));
 sg13g2_o21ai_1 _33805_ (.B1(net6836),
    .Y(_03250_),
    .A1(net1706),
    .A2(net6384));
 sg13g2_a221oi_1 _33806_ (.B2(_02005_),
    .C1(net7014),
    .B1(net5198),
    .A1(_21812_),
    .Y(_03251_),
    .A2(net5223));
 sg13g2_o21ai_1 _33807_ (.B1(_03251_),
    .Y(_03252_),
    .A1(_02208_),
    .A2(net5240));
 sg13g2_a22oi_1 _33808_ (.Y(_00704_),
    .B1(_03250_),
    .B2(_03252_),
    .A2(net6384),
    .A1(_17967_));
 sg13g2_a221oi_1 _33809_ (.B2(_21813_),
    .C1(net7013),
    .B1(net5885),
    .A1(_02071_),
    .Y(_03253_),
    .A2(net5938));
 sg13g2_o21ai_1 _33810_ (.B1(_03253_),
    .Y(_03254_),
    .A1(_02005_),
    .A2(net5240));
 sg13g2_o21ai_1 _33811_ (.B1(net6480),
    .Y(_03255_),
    .A1(net1564),
    .A2(net7084));
 sg13g2_nor2b_1 _33812_ (.A(_03255_),
    .B_N(_03254_),
    .Y(_03256_));
 sg13g2_a21o_1 _33813_ (.A2(net6386),
    .A1(net3401),
    .B1(_03256_),
    .X(_00705_));
 sg13g2_a22oi_1 _33814_ (.Y(_03257_),
    .B1(net5198),
    .B2(_02071_),
    .A2(net5976),
    .A1(_21813_));
 sg13g2_nor2_1 _33815_ (.A(net6836),
    .B(_03257_),
    .Y(_03258_));
 sg13g2_a22oi_1 _33816_ (.Y(_03259_),
    .B1(_02097_),
    .B2(net5132),
    .A2(net7014),
    .A1(net1367));
 sg13g2_a21oi_1 _33817_ (.A1(net3469),
    .A2(net6386),
    .Y(_03260_),
    .B1(_03258_));
 sg13g2_o21ai_1 _33818_ (.B1(_03260_),
    .Y(_00706_),
    .A1(net6386),
    .A2(_03259_));
 sg13g2_a22oi_1 _33819_ (.Y(_03261_),
    .B1(net5885),
    .B2(_02097_),
    .A2(net5976),
    .A1(_02071_));
 sg13g2_o21ai_1 _33820_ (.B1(_03261_),
    .Y(_03262_),
    .A1(_02244_),
    .A2(net5919));
 sg13g2_a221oi_1 _33821_ (.B2(_03262_),
    .C1(net6385),
    .B1(net5235),
    .A1(net1308),
    .Y(_03263_),
    .A2(net7014));
 sg13g2_a21oi_1 _33822_ (.A1(_17966_),
    .A2(net6386),
    .Y(_00707_),
    .B1(_03263_));
 sg13g2_o21ai_1 _33823_ (.B1(net6841),
    .Y(_03264_),
    .A1(net1715),
    .A2(net6385));
 sg13g2_a221oi_1 _33824_ (.B2(_02244_),
    .C1(net7013),
    .B1(net5198),
    .A1(_21843_),
    .Y(_03265_),
    .A2(net5223));
 sg13g2_o21ai_1 _33825_ (.B1(_03265_),
    .Y(_03266_),
    .A1(_02097_),
    .A2(net5240));
 sg13g2_a22oi_1 _33826_ (.Y(_00708_),
    .B1(_03264_),
    .B2(_03266_),
    .A2(net6385),
    .A1(_17965_));
 sg13g2_a22oi_1 _33827_ (.Y(_03267_),
    .B1(net5223),
    .B2(_02229_),
    .A2(net5156),
    .A1(_02244_));
 sg13g2_a21oi_1 _33828_ (.A1(_21843_),
    .A2(net5199),
    .Y(_03268_),
    .B1(net7013));
 sg13g2_a221oi_1 _33829_ (.B2(_03268_),
    .C1(net6387),
    .B1(_03267_),
    .A1(net1989),
    .Y(_03269_),
    .A2(net7013));
 sg13g2_a21oi_1 _33830_ (.A1(_17964_),
    .A2(net6386),
    .Y(_00709_),
    .B1(_03269_));
 sg13g2_nor2_1 _33831_ (.A(net3259),
    .B(net6480),
    .Y(_03270_));
 sg13g2_o21ai_1 _33832_ (.B1(net7084),
    .Y(_03271_),
    .A1(_02054_),
    .A2(net5151));
 sg13g2_a221oi_1 _33833_ (.B2(_02229_),
    .C1(_03271_),
    .B1(net5199),
    .A1(_21843_),
    .Y(_03272_),
    .A2(net5156));
 sg13g2_a21oi_1 _33834_ (.A1(net2323),
    .A2(net7013),
    .Y(_03273_),
    .B1(_03272_));
 sg13g2_a21oi_1 _33835_ (.A1(net6480),
    .A2(_03273_),
    .Y(_00710_),
    .B1(_03270_));
 sg13g2_o21ai_1 _33836_ (.B1(net6841),
    .Y(_03274_),
    .A1(net1963),
    .A2(net6385));
 sg13g2_a221oi_1 _33837_ (.B2(_02011_),
    .C1(net7013),
    .B1(net5223),
    .A1(_02229_),
    .Y(_03275_),
    .A2(net5156));
 sg13g2_o21ai_1 _33838_ (.B1(_03275_),
    .Y(_03276_),
    .A1(_02054_),
    .A2(net5122));
 sg13g2_a22oi_1 _33839_ (.Y(_00711_),
    .B1(_03274_),
    .B2(_03276_),
    .A2(net6386),
    .A1(_17963_));
 sg13g2_nor2_1 _33840_ (.A(net3418),
    .B(net6480),
    .Y(_03277_));
 sg13g2_nor2_1 _33841_ (.A(_02054_),
    .B(net5240),
    .Y(_03278_));
 sg13g2_a21oi_1 _33842_ (.A1(_21797_),
    .A2(net5223),
    .Y(_03279_),
    .B1(_03278_));
 sg13g2_a21oi_1 _33843_ (.A1(_02011_),
    .A2(net5199),
    .Y(_03280_),
    .B1(net7014));
 sg13g2_a22oi_1 _33844_ (.Y(_03281_),
    .B1(_03279_),
    .B2(_03280_),
    .A2(net7014),
    .A1(net2505));
 sg13g2_a21oi_1 _33845_ (.A1(net6484),
    .A2(_03281_),
    .Y(_00712_),
    .B1(_03277_));
 sg13g2_nand2_1 _33846_ (.Y(_03282_),
    .A(net3407),
    .B(net6385));
 sg13g2_nor2_1 _33847_ (.A(_02011_),
    .B(net5240),
    .Y(_03283_));
 sg13g2_nor2_1 _33848_ (.A(_21911_),
    .B(net5919),
    .Y(_03284_));
 sg13g2_o21ai_1 _33849_ (.B1(net7084),
    .Y(_03285_),
    .A1(_21797_),
    .A2(net5880));
 sg13g2_nor3_1 _33850_ (.A(_03283_),
    .B(_03284_),
    .C(_03285_),
    .Y(_03286_));
 sg13g2_o21ai_1 _33851_ (.B1(net6480),
    .Y(_03287_),
    .A1(net1314),
    .A2(net7084));
 sg13g2_o21ai_1 _33852_ (.B1(_03282_),
    .Y(_00713_),
    .A1(_03286_),
    .A2(_03287_));
 sg13g2_nor2_1 _33853_ (.A(_21911_),
    .B(net5880),
    .Y(_03288_));
 sg13g2_a21oi_1 _33854_ (.A1(_21907_),
    .A2(net5938),
    .Y(_03289_),
    .B1(_03288_));
 sg13g2_o21ai_1 _33855_ (.B1(_03289_),
    .Y(_03290_),
    .A1(_21797_),
    .A2(net6003));
 sg13g2_a221oi_1 _33856_ (.B2(_03290_),
    .C1(net6385),
    .B1(net5236),
    .A1(net1775),
    .Y(_03291_),
    .A2(net7013));
 sg13g2_a21oi_1 _33857_ (.A1(_17962_),
    .A2(net6386),
    .Y(_00714_),
    .B1(_03291_));
 sg13g2_a21oi_1 _33858_ (.A1(net1802),
    .A2(net7016),
    .Y(_03292_),
    .B1(net6385));
 sg13g2_o21ai_1 _33859_ (.B1(_03292_),
    .Y(_03293_),
    .A1(_21911_),
    .A2(_02370_));
 sg13g2_a21oi_1 _33860_ (.A1(_21907_),
    .A2(_02346_),
    .Y(_03294_),
    .B1(_03293_));
 sg13g2_a21oi_1 _33861_ (.A1(_17961_),
    .A2(net6383),
    .Y(_00715_),
    .B1(_03294_));
 sg13g2_a22oi_1 _33862_ (.Y(_03295_),
    .B1(_21907_),
    .B2(net6866),
    .A2(net6385),
    .A1(net2730));
 sg13g2_inv_1 _33863_ (.Y(_00716_),
    .A(_03295_));
 sg13g2_nor2_2 _33864_ (.A(_24689_[0]),
    .B(net5075),
    .Y(_03296_));
 sg13g2_o21ai_1 _33865_ (.B1(net3578),
    .Y(_03297_),
    .A1(_24689_[0]),
    .A2(net5075));
 sg13g2_mux2_1 _33866_ (.A0(net5075),
    .A1(_03296_),
    .S(net3578),
    .X(_00717_));
 sg13g2_nand3_1 _33867_ (.B(net1387),
    .C(net5076),
    .A(net3578),
    .Y(_03298_));
 sg13g2_nand2_1 _33868_ (.Y(_03299_),
    .A(net6606),
    .B(_03298_));
 sg13g2_a21oi_1 _33869_ (.A1(_18346_),
    .A2(_03297_),
    .Y(_00718_),
    .B1(_03299_));
 sg13g2_nand3_1 _33870_ (.B(net6606),
    .C(_03298_),
    .A(net1157),
    .Y(_03300_));
 sg13g2_o21ai_1 _33871_ (.B1(_03300_),
    .Y(_00719_),
    .A1(net1157),
    .A2(_03298_));
 sg13g2_nand2_1 _33872_ (.Y(_03301_),
    .A(net1164),
    .B(_03296_));
 sg13g2_nand3_1 _33873_ (.B(net1387),
    .C(net1157),
    .A(net3578),
    .Y(_03302_));
 sg13g2_nor2_1 _33874_ (.A(_18347_),
    .B(_03302_),
    .Y(_03303_));
 sg13g2_xnor2_1 _33875_ (.Y(_03304_),
    .A(_18347_),
    .B(_03302_));
 sg13g2_o21ai_1 _33876_ (.B1(_03301_),
    .Y(_00720_),
    .A1(net5067),
    .A2(_03304_));
 sg13g2_nand2_1 _33877_ (.Y(_03305_),
    .A(net1235),
    .B(_03296_));
 sg13g2_and2_1 _33878_ (.A(net1235),
    .B(_03303_),
    .X(_03306_));
 sg13g2_o21ai_1 _33879_ (.B1(net5076),
    .Y(_03307_),
    .A1(net1235),
    .A2(_03303_));
 sg13g2_o21ai_1 _33880_ (.B1(_03305_),
    .Y(_00721_),
    .A1(_03306_),
    .A2(_03307_));
 sg13g2_nand2_1 _33881_ (.Y(_03308_),
    .A(net1251),
    .B(_03296_));
 sg13g2_xnor2_1 _33882_ (.Y(_03309_),
    .A(net1251),
    .B(_03306_));
 sg13g2_o21ai_1 _33883_ (.B1(_03308_),
    .Y(_00722_),
    .A1(net5067),
    .A2(_03309_));
 sg13g2_nand2_1 _33884_ (.Y(_03310_),
    .A(net1255),
    .B(_03296_));
 sg13g2_nand3_1 _33885_ (.B(net1255),
    .C(_03306_),
    .A(net1251),
    .Y(_03311_));
 sg13g2_a21o_1 _33886_ (.A2(_03306_),
    .A1(net1251),
    .B1(net1255),
    .X(_03312_));
 sg13g2_nand3_1 _33887_ (.B(_03311_),
    .C(_03312_),
    .A(net5076),
    .Y(_03313_));
 sg13g2_nand2_1 _33888_ (.Y(_00723_),
    .A(_03310_),
    .B(_03313_));
 sg13g2_nand2_1 _33889_ (.Y(_03314_),
    .A(net1169),
    .B(_03296_));
 sg13g2_nor2_1 _33890_ (.A(_18349_),
    .B(_03311_),
    .Y(_03315_));
 sg13g2_xnor2_1 _33891_ (.Y(_03316_),
    .A(_18349_),
    .B(_03311_));
 sg13g2_o21ai_1 _33892_ (.B1(_03314_),
    .Y(_00724_),
    .A1(net5068),
    .A2(_03316_));
 sg13g2_nand2_1 _33893_ (.Y(_03317_),
    .A(net1286),
    .B(_03296_));
 sg13g2_xnor2_1 _33894_ (.Y(_03318_),
    .A(net1286),
    .B(_03315_));
 sg13g2_o21ai_1 _33895_ (.B1(_03317_),
    .Y(_00725_),
    .A1(net5067),
    .A2(_03318_));
 sg13g2_and3_1 _33896_ (.X(_03319_),
    .A(net1286),
    .B(net5076),
    .C(_03315_));
 sg13g2_o21ai_1 _33897_ (.B1(net6606),
    .Y(_03320_),
    .A1(net1149),
    .A2(_03319_));
 sg13g2_a21oi_1 _33898_ (.A1(net1149),
    .A2(_03319_),
    .Y(_00726_),
    .B1(_03320_));
 sg13g2_nor2_1 _33899_ (.A(net1187),
    .B(net7083),
    .Y(_03321_));
 sg13g2_a21oi_1 _33900_ (.A1(net1187),
    .A2(_19809_),
    .Y(_00727_),
    .B1(_03321_));
 sg13g2_a21o_1 _33901_ (.A2(_19809_),
    .A1(net1187),
    .B1(net3693),
    .X(_03322_));
 sg13g2_nand3_1 _33902_ (.B(net3693),
    .C(_19809_),
    .A(net1187),
    .Y(_03323_));
 sg13g2_and3_1 _33903_ (.X(_00728_),
    .A(net6606),
    .B(_03322_),
    .C(_03323_));
 sg13g2_nand4_1 _33904_ (.B(\perf_total[1] ),
    .C(net1266),
    .A(net1187),
    .Y(_03324_),
    .D(net7084));
 sg13g2_nand2_1 _33905_ (.Y(_03325_),
    .A(net6606),
    .B(_03324_));
 sg13g2_a21oi_1 _33906_ (.A1(_18351_),
    .A2(_03323_),
    .Y(_00729_),
    .B1(_03325_));
 sg13g2_nor2b_1 _33907_ (.A(net1161),
    .B_N(_03324_),
    .Y(_03326_));
 sg13g2_a21oi_1 _33908_ (.A1(net1161),
    .A2(_03325_),
    .Y(_00730_),
    .B1(_03326_));
 sg13g2_and4_1 _33909_ (.A(net1187),
    .B(\perf_total[1] ),
    .C(\perf_total[2] ),
    .D(net1161),
    .X(_03327_));
 sg13g2_a21oi_1 _33910_ (.A1(_19809_),
    .A2(_03327_),
    .Y(_03328_),
    .B1(net1193));
 sg13g2_and3_2 _33911_ (.X(_03329_),
    .A(net1193),
    .B(net7084),
    .C(_03327_));
 sg13g2_nor3_1 _33912_ (.A(_24689_[0]),
    .B(net1194),
    .C(_03329_),
    .Y(_00731_));
 sg13g2_a21oi_1 _33913_ (.A1(net1155),
    .A2(net6607),
    .Y(_03330_),
    .B1(_03329_));
 sg13g2_a21oi_1 _33914_ (.A1(net1155),
    .A2(_03329_),
    .Y(_00732_),
    .B1(_03330_));
 sg13g2_and3_2 _33915_ (.X(_03331_),
    .A(net1155),
    .B(net1183),
    .C(_03329_));
 sg13g2_a21oi_1 _33916_ (.A1(net1155),
    .A2(_03329_),
    .Y(_03332_),
    .B1(net1183));
 sg13g2_nor3_1 _33917_ (.A(_24689_[0]),
    .B(_03331_),
    .C(net1184),
    .Y(_00733_));
 sg13g2_a21oi_1 _33918_ (.A1(net1279),
    .A2(net6607),
    .Y(_03333_),
    .B1(_03331_));
 sg13g2_nand2_1 _33919_ (.Y(_03334_),
    .A(net1279),
    .B(_03331_));
 sg13g2_nor2b_1 _33920_ (.A(_03333_),
    .B_N(_03334_),
    .Y(_00734_));
 sg13g2_o21ai_1 _33921_ (.B1(net6607),
    .Y(_03335_),
    .A1(_18354_),
    .A2(_03334_));
 sg13g2_a21oi_1 _33922_ (.A1(_18354_),
    .A2(_03334_),
    .Y(_00735_),
    .B1(_03335_));
 sg13g2_nand4_1 _33923_ (.B(\perf_total[8] ),
    .C(_18355_),
    .A(net1279),
    .Y(_03336_),
    .D(_03331_));
 sg13g2_o21ai_1 _33924_ (.B1(net1280),
    .Y(_00736_),
    .A1(_18355_),
    .A2(_03335_));
 sg13g2_and2_1 _33925_ (.A(\u_inv.d_next[2] ),
    .B(\u_inv.d_reg[2] ),
    .X(_03337_));
 sg13g2_xor2_1 _33926_ (.B(\u_inv.d_reg[2] ),
    .A(\u_inv.d_next[2] ),
    .X(_03338_));
 sg13g2_nand2_1 _33927_ (.Y(_03339_),
    .A(\u_inv.d_next[1] ),
    .B(net7293));
 sg13g2_xnor2_1 _33928_ (.Y(_03340_),
    .A(\u_inv.d_next[1] ),
    .B(net7293));
 sg13g2_nand2b_1 _33929_ (.Y(_03341_),
    .B(net7294),
    .A_N(\u_inv.d_next[0] ));
 sg13g2_nor2b_1 _33930_ (.A(net7293),
    .B_N(\u_inv.d_next[1] ),
    .Y(_03342_));
 sg13g2_a21oi_1 _33931_ (.A1(_03340_),
    .A2(_03341_),
    .Y(_03343_),
    .B1(_03342_));
 sg13g2_xnor2_1 _33932_ (.Y(_03344_),
    .A(_03338_),
    .B(_03343_));
 sg13g2_nor2_1 _33933_ (.A(net6218),
    .B(_03344_),
    .Y(_03345_));
 sg13g2_nor2_1 _33934_ (.A(net7330),
    .B(\u_inv.d_next[2] ),
    .Y(_03346_));
 sg13g2_nand2_1 _33935_ (.Y(_03347_),
    .A(\u_inv.d_next[0] ),
    .B(net7294));
 sg13g2_o21ai_1 _33936_ (.B1(_03339_),
    .Y(_03348_),
    .A1(_03340_),
    .A2(_03347_));
 sg13g2_xnor2_1 _33937_ (.Y(_03349_),
    .A(_03338_),
    .B(_03348_));
 sg13g2_a21oi_1 _33938_ (.A1(net7330),
    .A2(_03349_),
    .Y(_03350_),
    .B1(_03346_));
 sg13g2_a21oi_2 _33939_ (.B1(_03345_),
    .Y(_03351_),
    .A2(_03350_),
    .A1(net6218));
 sg13g2_nand2_1 _33940_ (.Y(_03352_),
    .A(net7330),
    .B(net7294));
 sg13g2_xnor2_1 _33941_ (.Y(_03353_),
    .A(\u_inv.d_next[0] ),
    .B(_03352_));
 sg13g2_xor2_1 _33942_ (.B(_03352_),
    .A(\u_inv.d_next[0] ),
    .X(_03354_));
 sg13g2_xnor2_1 _33943_ (.Y(_03355_),
    .A(\u_inv.d_next[256] ),
    .B(\u_inv.d_reg[256] ));
 sg13g2_inv_1 _33944_ (.Y(_03356_),
    .A(_03355_));
 sg13g2_xor2_1 _33945_ (.B(\u_inv.d_reg[207] ),
    .A(\u_inv.d_next[207] ),
    .X(_03357_));
 sg13g2_nor2_1 _33946_ (.A(\u_inv.d_next[206] ),
    .B(\u_inv.d_reg[206] ),
    .Y(_03358_));
 sg13g2_nand2_1 _33947_ (.Y(_03359_),
    .A(\u_inv.d_next[206] ),
    .B(\u_inv.d_reg[206] ));
 sg13g2_xor2_1 _33948_ (.B(\u_inv.d_reg[206] ),
    .A(\u_inv.d_next[206] ),
    .X(_03360_));
 sg13g2_nand2_1 _33949_ (.Y(_03361_),
    .A(_03357_),
    .B(_03360_));
 sg13g2_nor2_1 _33950_ (.A(\u_inv.d_next[205] ),
    .B(\u_inv.d_reg[205] ),
    .Y(_03362_));
 sg13g2_nand2_1 _33951_ (.Y(_03363_),
    .A(\u_inv.d_next[205] ),
    .B(\u_inv.d_reg[205] ));
 sg13g2_nand2_1 _33952_ (.Y(_03364_),
    .A(\u_inv.d_next[204] ),
    .B(\u_inv.d_reg[204] ));
 sg13g2_inv_1 _33953_ (.Y(_03365_),
    .A(_03364_));
 sg13g2_o21ai_1 _33954_ (.B1(_03363_),
    .Y(_03366_),
    .A1(_03362_),
    .A2(_03364_));
 sg13g2_nand2b_2 _33955_ (.Y(_03367_),
    .B(_03363_),
    .A_N(_03362_));
 sg13g2_xnor2_1 _33956_ (.Y(_03368_),
    .A(\u_inv.d_next[204] ),
    .B(\u_inv.d_reg[204] ));
 sg13g2_inv_1 _33957_ (.Y(_03369_),
    .A(_03368_));
 sg13g2_nor2_1 _33958_ (.A(_03367_),
    .B(_03368_),
    .Y(_03370_));
 sg13g2_nand2_1 _33959_ (.Y(_03371_),
    .A(\u_inv.d_next[202] ),
    .B(\u_inv.d_reg[202] ));
 sg13g2_a21oi_1 _33960_ (.A1(_18116_),
    .A2(_18411_),
    .Y(_03372_),
    .B1(_03371_));
 sg13g2_a21oi_1 _33961_ (.A1(\u_inv.d_next[203] ),
    .A2(\u_inv.d_reg[203] ),
    .Y(_03373_),
    .B1(_03372_));
 sg13g2_xnor2_1 _33962_ (.Y(_03374_),
    .A(\u_inv.d_next[203] ),
    .B(\u_inv.d_reg[203] ));
 sg13g2_xnor2_1 _33963_ (.Y(_03375_),
    .A(\u_inv.d_next[202] ),
    .B(\u_inv.d_reg[202] ));
 sg13g2_or2_1 _33964_ (.X(_03376_),
    .B(_03375_),
    .A(_03374_));
 sg13g2_or2_1 _33965_ (.X(_03377_),
    .B(\u_inv.d_reg[201] ),
    .A(\u_inv.d_next[201] ));
 sg13g2_nand2_1 _33966_ (.Y(_03378_),
    .A(\u_inv.d_next[201] ),
    .B(\u_inv.d_reg[201] ));
 sg13g2_nand2_1 _33967_ (.Y(_03379_),
    .A(\u_inv.d_next[200] ),
    .B(\u_inv.d_reg[200] ));
 sg13g2_inv_1 _33968_ (.Y(_03380_),
    .A(_03379_));
 sg13g2_nand2_1 _33969_ (.Y(_03381_),
    .A(_03378_),
    .B(_03379_));
 sg13g2_nand2_1 _33970_ (.Y(_03382_),
    .A(_03377_),
    .B(_03381_));
 sg13g2_and2_1 _33971_ (.A(_03377_),
    .B(_03378_),
    .X(_03383_));
 sg13g2_nand2_1 _33972_ (.Y(_03384_),
    .A(_03377_),
    .B(_03378_));
 sg13g2_xor2_1 _33973_ (.B(\u_inv.d_reg[200] ),
    .A(\u_inv.d_next[200] ),
    .X(_03385_));
 sg13g2_and2_1 _33974_ (.A(_03383_),
    .B(_03385_),
    .X(_03386_));
 sg13g2_nor2_1 _33975_ (.A(\u_inv.d_next[199] ),
    .B(\u_inv.d_reg[199] ),
    .Y(_03387_));
 sg13g2_nand2_1 _33976_ (.Y(_03388_),
    .A(\u_inv.d_next[199] ),
    .B(\u_inv.d_reg[199] ));
 sg13g2_nor2b_2 _33977_ (.A(_03387_),
    .B_N(_03388_),
    .Y(_03389_));
 sg13g2_nand2b_1 _33978_ (.Y(_03390_),
    .B(_03388_),
    .A_N(_03387_));
 sg13g2_nand2_1 _33979_ (.Y(_03391_),
    .A(\u_inv.d_next[198] ),
    .B(\u_inv.d_reg[198] ));
 sg13g2_xor2_1 _33980_ (.B(\u_inv.d_reg[198] ),
    .A(\u_inv.d_next[198] ),
    .X(_03392_));
 sg13g2_nand2_1 _33981_ (.Y(_03393_),
    .A(_03389_),
    .B(_03392_));
 sg13g2_a22oi_1 _33982_ (.Y(_03394_),
    .B1(\u_inv.d_reg[196] ),
    .B2(\u_inv.d_next[196] ),
    .A2(\u_inv.d_reg[197] ),
    .A1(\u_inv.d_next[197] ));
 sg13g2_inv_1 _33983_ (.Y(_03395_),
    .A(_03394_));
 sg13g2_o21ai_1 _33984_ (.B1(_03395_),
    .Y(_03396_),
    .A1(\u_inv.d_next[197] ),
    .A2(\u_inv.d_reg[197] ));
 sg13g2_nor2_1 _33985_ (.A(_03393_),
    .B(_03396_),
    .Y(_03397_));
 sg13g2_o21ai_1 _33986_ (.B1(_03388_),
    .Y(_03398_),
    .A1(_03387_),
    .A2(_03391_));
 sg13g2_nor2_1 _33987_ (.A(_03397_),
    .B(_03398_),
    .Y(_03399_));
 sg13g2_o21ai_1 _33988_ (.B1(_03373_),
    .Y(_03400_),
    .A1(_03376_),
    .A2(_03382_));
 sg13g2_a21oi_1 _33989_ (.A1(_03370_),
    .A2(_03400_),
    .Y(_03401_),
    .B1(_03366_));
 sg13g2_nor2_1 _33990_ (.A(_03361_),
    .B(_03401_),
    .Y(_03402_));
 sg13g2_nor2_1 _33991_ (.A(_03361_),
    .B(_03376_),
    .Y(_03403_));
 sg13g2_nand3_1 _33992_ (.B(_03386_),
    .C(_03403_),
    .A(_03370_),
    .Y(_03404_));
 sg13g2_o21ai_1 _33993_ (.B1(_03359_),
    .Y(_03405_),
    .A1(_18115_),
    .A2(_18407_));
 sg13g2_o21ai_1 _33994_ (.B1(_03405_),
    .Y(_03406_),
    .A1(\u_inv.d_next[207] ),
    .A2(\u_inv.d_reg[207] ));
 sg13g2_nand2_1 _33995_ (.Y(_03407_),
    .A(\u_inv.d_next[195] ),
    .B(\u_inv.d_reg[195] ));
 sg13g2_nor2_1 _33996_ (.A(\u_inv.d_next[195] ),
    .B(\u_inv.d_reg[195] ),
    .Y(_03408_));
 sg13g2_xnor2_1 _33997_ (.Y(_03409_),
    .A(\u_inv.d_next[195] ),
    .B(\u_inv.d_reg[195] ));
 sg13g2_nand2_1 _33998_ (.Y(_03410_),
    .A(\u_inv.d_next[194] ),
    .B(\u_inv.d_reg[194] ));
 sg13g2_xnor2_1 _33999_ (.Y(_03411_),
    .A(\u_inv.d_next[194] ),
    .B(\u_inv.d_reg[194] ));
 sg13g2_nor2_1 _34000_ (.A(_03409_),
    .B(_03411_),
    .Y(_03412_));
 sg13g2_nand2b_1 _34001_ (.Y(_03413_),
    .B(\u_inv.d_reg[193] ),
    .A_N(\u_inv.d_next[193] ));
 sg13g2_nor2b_1 _34002_ (.A(\u_inv.d_reg[193] ),
    .B_N(\u_inv.d_next[193] ),
    .Y(_03414_));
 sg13g2_xnor2_1 _34003_ (.Y(_03415_),
    .A(\u_inv.d_next[193] ),
    .B(\u_inv.d_reg[193] ));
 sg13g2_xor2_1 _34004_ (.B(\u_inv.d_reg[193] ),
    .A(\u_inv.d_next[193] ),
    .X(_03416_));
 sg13g2_nand2_1 _34005_ (.Y(_03417_),
    .A(\u_inv.d_next[192] ),
    .B(\u_inv.d_reg[192] ));
 sg13g2_nand2_1 _34006_ (.Y(_03418_),
    .A(\u_inv.d_next[193] ),
    .B(\u_inv.d_reg[193] ));
 sg13g2_o21ai_1 _34007_ (.B1(_03418_),
    .Y(_03419_),
    .A1(_03415_),
    .A2(_03417_));
 sg13g2_o21ai_1 _34008_ (.B1(_03407_),
    .Y(_03420_),
    .A1(_03408_),
    .A2(_03410_));
 sg13g2_a21o_2 _34009_ (.A2(_03419_),
    .A1(_03412_),
    .B1(_03420_),
    .X(_03421_));
 sg13g2_xor2_1 _34010_ (.B(\u_inv.d_reg[197] ),
    .A(\u_inv.d_next[197] ),
    .X(_03422_));
 sg13g2_xnor2_1 _34011_ (.Y(_03423_),
    .A(\u_inv.d_next[197] ),
    .B(\u_inv.d_reg[197] ));
 sg13g2_xor2_1 _34012_ (.B(\u_inv.d_reg[196] ),
    .A(\u_inv.d_next[196] ),
    .X(_03424_));
 sg13g2_xnor2_1 _34013_ (.Y(_03425_),
    .A(\u_inv.d_next[196] ),
    .B(\u_inv.d_reg[196] ));
 sg13g2_nand2_1 _34014_ (.Y(_03426_),
    .A(_03422_),
    .B(_03424_));
 sg13g2_or2_1 _34015_ (.X(_03427_),
    .B(_03426_),
    .A(_03393_));
 sg13g2_or2_1 _34016_ (.X(_03428_),
    .B(_03427_),
    .A(_03404_));
 sg13g2_nor2b_1 _34017_ (.A(_03428_),
    .B_N(_03421_),
    .Y(_03429_));
 sg13g2_o21ai_1 _34018_ (.B1(_03406_),
    .Y(_03430_),
    .A1(_03399_),
    .A2(_03404_));
 sg13g2_nor3_2 _34019_ (.A(_03402_),
    .B(_03429_),
    .C(_03430_),
    .Y(_03431_));
 sg13g2_xnor2_1 _34020_ (.Y(_03432_),
    .A(\u_inv.d_next[221] ),
    .B(\u_inv.d_reg[221] ));
 sg13g2_nand2_1 _34021_ (.Y(_03433_),
    .A(\u_inv.d_next[220] ),
    .B(\u_inv.d_reg[220] ));
 sg13g2_xnor2_1 _34022_ (.Y(_03434_),
    .A(\u_inv.d_next[220] ),
    .B(\u_inv.d_reg[220] ));
 sg13g2_inv_1 _34023_ (.Y(_03435_),
    .A(_03434_));
 sg13g2_nor2_1 _34024_ (.A(_03432_),
    .B(_03434_),
    .Y(_03436_));
 sg13g2_xnor2_1 _34025_ (.Y(_03437_),
    .A(\u_inv.d_next[223] ),
    .B(\u_inv.d_reg[223] ));
 sg13g2_nand2_1 _34026_ (.Y(_03438_),
    .A(\u_inv.d_next[222] ),
    .B(\u_inv.d_reg[222] ));
 sg13g2_xnor2_1 _34027_ (.Y(_03439_),
    .A(\u_inv.d_next[222] ),
    .B(\u_inv.d_reg[222] ));
 sg13g2_inv_1 _34028_ (.Y(_03440_),
    .A(_03439_));
 sg13g2_nor4_1 _34029_ (.A(_03432_),
    .B(_03434_),
    .C(_03437_),
    .D(_03439_),
    .Y(_03441_));
 sg13g2_nor2_2 _34030_ (.A(\u_inv.d_next[219] ),
    .B(\u_inv.d_reg[219] ),
    .Y(_03442_));
 sg13g2_nand2_1 _34031_ (.Y(_03443_),
    .A(\u_inv.d_next[219] ),
    .B(\u_inv.d_reg[219] ));
 sg13g2_nor2b_2 _34032_ (.A(_03442_),
    .B_N(_03443_),
    .Y(_03444_));
 sg13g2_nand2b_1 _34033_ (.Y(_03445_),
    .B(_03443_),
    .A_N(_03442_));
 sg13g2_nand2_1 _34034_ (.Y(_03446_),
    .A(\u_inv.d_next[218] ),
    .B(_18396_));
 sg13g2_xor2_1 _34035_ (.B(\u_inv.d_reg[218] ),
    .A(\u_inv.d_next[218] ),
    .X(_03447_));
 sg13g2_nand2_1 _34036_ (.Y(_03448_),
    .A(_03444_),
    .B(_03447_));
 sg13g2_xor2_1 _34037_ (.B(\u_inv.d_reg[217] ),
    .A(\u_inv.d_next[217] ),
    .X(_03449_));
 sg13g2_xnor2_1 _34038_ (.Y(_03450_),
    .A(\u_inv.d_next[217] ),
    .B(\u_inv.d_reg[217] ));
 sg13g2_nand2_1 _34039_ (.Y(_03451_),
    .A(\u_inv.d_next[216] ),
    .B(\u_inv.d_reg[216] ));
 sg13g2_xor2_1 _34040_ (.B(\u_inv.d_reg[216] ),
    .A(\u_inv.d_next[216] ),
    .X(_03452_));
 sg13g2_nand2_1 _34041_ (.Y(_03453_),
    .A(_03449_),
    .B(_03452_));
 sg13g2_inv_1 _34042_ (.Y(_03454_),
    .A(_03453_));
 sg13g2_and4_1 _34043_ (.A(_03441_),
    .B(_03444_),
    .C(_03447_),
    .D(_03454_),
    .X(_03455_));
 sg13g2_xor2_1 _34044_ (.B(\u_inv.d_reg[215] ),
    .A(\u_inv.d_next[215] ),
    .X(_03456_));
 sg13g2_xnor2_1 _34045_ (.Y(_03457_),
    .A(\u_inv.d_next[215] ),
    .B(\u_inv.d_reg[215] ));
 sg13g2_nand2_1 _34046_ (.Y(_03458_),
    .A(\u_inv.d_next[214] ),
    .B(\u_inv.d_reg[214] ));
 sg13g2_xor2_1 _34047_ (.B(\u_inv.d_reg[214] ),
    .A(\u_inv.d_next[214] ),
    .X(_03459_));
 sg13g2_xnor2_1 _34048_ (.Y(_03460_),
    .A(\u_inv.d_next[214] ),
    .B(\u_inv.d_reg[214] ));
 sg13g2_nor2_1 _34049_ (.A(_03457_),
    .B(_03460_),
    .Y(_03461_));
 sg13g2_xor2_1 _34050_ (.B(\u_inv.d_reg[213] ),
    .A(\u_inv.d_next[213] ),
    .X(_03462_));
 sg13g2_xnor2_1 _34051_ (.Y(_03463_),
    .A(\u_inv.d_next[213] ),
    .B(\u_inv.d_reg[213] ));
 sg13g2_and2_1 _34052_ (.A(\u_inv.d_next[212] ),
    .B(\u_inv.d_reg[212] ),
    .X(_03464_));
 sg13g2_xor2_1 _34053_ (.B(\u_inv.d_reg[212] ),
    .A(\u_inv.d_next[212] ),
    .X(_03465_));
 sg13g2_and2_1 _34054_ (.A(_03462_),
    .B(_03465_),
    .X(_03466_));
 sg13g2_inv_1 _34055_ (.Y(_03467_),
    .A(_03466_));
 sg13g2_nand2_1 _34056_ (.Y(_03468_),
    .A(_03461_),
    .B(_03466_));
 sg13g2_xor2_1 _34057_ (.B(\u_inv.d_reg[211] ),
    .A(\u_inv.d_next[211] ),
    .X(_03469_));
 sg13g2_xor2_1 _34058_ (.B(\u_inv.d_reg[210] ),
    .A(\u_inv.d_next[210] ),
    .X(_03470_));
 sg13g2_and2_1 _34059_ (.A(_03469_),
    .B(_03470_),
    .X(_03471_));
 sg13g2_nand3_1 _34060_ (.B(_03466_),
    .C(_03471_),
    .A(_03461_),
    .Y(_03472_));
 sg13g2_xor2_1 _34061_ (.B(\u_inv.d_reg[209] ),
    .A(\u_inv.d_next[209] ),
    .X(_03473_));
 sg13g2_xnor2_1 _34062_ (.Y(_03474_),
    .A(\u_inv.d_next[209] ),
    .B(\u_inv.d_reg[209] ));
 sg13g2_xor2_1 _34063_ (.B(\u_inv.d_reg[208] ),
    .A(\u_inv.d_next[208] ),
    .X(_03475_));
 sg13g2_xnor2_1 _34064_ (.Y(_03476_),
    .A(\u_inv.d_next[208] ),
    .B(\u_inv.d_reg[208] ));
 sg13g2_nand2_1 _34065_ (.Y(_03477_),
    .A(_03473_),
    .B(_03475_));
 sg13g2_nor2_1 _34066_ (.A(_03472_),
    .B(_03477_),
    .Y(_03478_));
 sg13g2_inv_1 _34067_ (.Y(_03479_),
    .A(_03478_));
 sg13g2_nand2_1 _34068_ (.Y(_03480_),
    .A(_03455_),
    .B(_03478_));
 sg13g2_a21oi_1 _34069_ (.A1(_18110_),
    .A2(_18397_),
    .Y(_03481_),
    .B1(_03451_));
 sg13g2_a21oi_1 _34070_ (.A1(\u_inv.d_next[217] ),
    .A2(\u_inv.d_reg[217] ),
    .Y(_03482_),
    .B1(_03481_));
 sg13g2_nor2_1 _34071_ (.A(_03448_),
    .B(_03482_),
    .Y(_03483_));
 sg13g2_and2_1 _34072_ (.A(\u_inv.d_next[218] ),
    .B(\u_inv.d_reg[218] ),
    .X(_03484_));
 sg13g2_nand2_1 _34073_ (.Y(_03485_),
    .A(\u_inv.d_next[218] ),
    .B(\u_inv.d_reg[218] ));
 sg13g2_a21oi_2 _34074_ (.B1(_03442_),
    .Y(_03486_),
    .A2(_03485_),
    .A1(_03443_));
 sg13g2_o21ai_1 _34075_ (.B1(_03441_),
    .Y(_03487_),
    .A1(_03483_),
    .A2(_03486_));
 sg13g2_a21oi_1 _34076_ (.A1(_18108_),
    .A2(_18391_),
    .Y(_03488_),
    .B1(_03438_));
 sg13g2_a21oi_1 _34077_ (.A1(\u_inv.d_next[223] ),
    .A2(\u_inv.d_reg[223] ),
    .Y(_03489_),
    .B1(_03488_));
 sg13g2_o21ai_1 _34078_ (.B1(_03433_),
    .Y(_03490_),
    .A1(_18109_),
    .A2(_18393_));
 sg13g2_o21ai_1 _34079_ (.B1(_03490_),
    .Y(_03491_),
    .A1(\u_inv.d_next[221] ),
    .A2(\u_inv.d_reg[221] ));
 sg13g2_or3_1 _34080_ (.A(_03437_),
    .B(_03439_),
    .C(_03491_),
    .X(_03492_));
 sg13g2_nand3_1 _34081_ (.B(_03489_),
    .C(_03492_),
    .A(_03487_),
    .Y(_03493_));
 sg13g2_a22oi_1 _34082_ (.Y(_03494_),
    .B1(\u_inv.d_reg[208] ),
    .B2(\u_inv.d_next[208] ),
    .A2(\u_inv.d_reg[209] ),
    .A1(\u_inv.d_next[209] ));
 sg13g2_a21oi_2 _34083_ (.B1(_03494_),
    .Y(_03495_),
    .A2(_18405_),
    .A1(_18114_));
 sg13g2_a22oi_1 _34084_ (.Y(_03496_),
    .B1(\u_inv.d_reg[210] ),
    .B2(\u_inv.d_next[210] ),
    .A2(\u_inv.d_reg[211] ),
    .A1(\u_inv.d_next[211] ));
 sg13g2_inv_1 _34085_ (.Y(_03497_),
    .A(_03496_));
 sg13g2_o21ai_1 _34086_ (.B1(_03497_),
    .Y(_03498_),
    .A1(\u_inv.d_next[211] ),
    .A2(\u_inv.d_reg[211] ));
 sg13g2_a21oi_1 _34087_ (.A1(_18111_),
    .A2(_18399_),
    .Y(_03499_),
    .B1(_03458_));
 sg13g2_a21oi_1 _34088_ (.A1(\u_inv.d_next[215] ),
    .A2(\u_inv.d_reg[215] ),
    .Y(_03500_),
    .B1(_03499_));
 sg13g2_o21ai_1 _34089_ (.B1(_03464_),
    .Y(_03501_),
    .A1(\u_inv.d_next[213] ),
    .A2(\u_inv.d_reg[213] ));
 sg13g2_o21ai_1 _34090_ (.B1(_03501_),
    .Y(_03502_),
    .A1(_18112_),
    .A2(_18401_));
 sg13g2_nand2_1 _34091_ (.Y(_03503_),
    .A(_03471_),
    .B(_03495_));
 sg13g2_a21oi_1 _34092_ (.A1(_03498_),
    .A2(_03503_),
    .Y(_03504_),
    .B1(_03468_));
 sg13g2_a21oi_1 _34093_ (.A1(_03461_),
    .A2(_03502_),
    .Y(_03505_),
    .B1(_03504_));
 sg13g2_nand2_2 _34094_ (.Y(_03506_),
    .A(_03500_),
    .B(_03505_));
 sg13g2_a21oi_1 _34095_ (.A1(_03455_),
    .A2(_03506_),
    .Y(_03507_),
    .B1(_03493_));
 sg13g2_o21ai_1 _34096_ (.B1(_03507_),
    .Y(_03508_),
    .A1(_03431_),
    .A2(_03480_));
 sg13g2_nor2_1 _34097_ (.A(\u_inv.d_next[239] ),
    .B(\u_inv.d_reg[239] ),
    .Y(_03509_));
 sg13g2_nand2_1 _34098_ (.Y(_03510_),
    .A(\u_inv.d_next[239] ),
    .B(\u_inv.d_reg[239] ));
 sg13g2_nor2b_1 _34099_ (.A(_03509_),
    .B_N(_03510_),
    .Y(_03511_));
 sg13g2_nand2b_2 _34100_ (.Y(_03512_),
    .B(_03510_),
    .A_N(_03509_));
 sg13g2_nand2_1 _34101_ (.Y(_03513_),
    .A(\u_inv.d_next[238] ),
    .B(\u_inv.d_reg[238] ));
 sg13g2_xor2_1 _34102_ (.B(\u_inv.d_reg[238] ),
    .A(\u_inv.d_next[238] ),
    .X(_03514_));
 sg13g2_and2_1 _34103_ (.A(_03511_),
    .B(_03514_),
    .X(_03515_));
 sg13g2_nor2_1 _34104_ (.A(\u_inv.d_next[237] ),
    .B(\u_inv.d_reg[237] ),
    .Y(_03516_));
 sg13g2_nand2_1 _34105_ (.Y(_03517_),
    .A(\u_inv.d_next[237] ),
    .B(\u_inv.d_reg[237] ));
 sg13g2_nand2b_2 _34106_ (.Y(_03518_),
    .B(_03517_),
    .A_N(_03516_));
 sg13g2_nand2_1 _34107_ (.Y(_03519_),
    .A(\u_inv.d_next[236] ),
    .B(\u_inv.d_reg[236] ));
 sg13g2_xnor2_1 _34108_ (.Y(_03520_),
    .A(\u_inv.d_next[236] ),
    .B(\u_inv.d_reg[236] ));
 sg13g2_nor2_1 _34109_ (.A(_03518_),
    .B(_03520_),
    .Y(_03521_));
 sg13g2_and2_1 _34110_ (.A(_03515_),
    .B(_03521_),
    .X(_03522_));
 sg13g2_nor2_1 _34111_ (.A(\u_inv.d_next[233] ),
    .B(\u_inv.d_reg[233] ),
    .Y(_03523_));
 sg13g2_nand2_1 _34112_ (.Y(_03524_),
    .A(\u_inv.d_next[233] ),
    .B(\u_inv.d_reg[233] ));
 sg13g2_nor2b_2 _34113_ (.A(_03523_),
    .B_N(_03524_),
    .Y(_03525_));
 sg13g2_nand2b_1 _34114_ (.Y(_03526_),
    .B(_03524_),
    .A_N(_03523_));
 sg13g2_nand2_1 _34115_ (.Y(_03527_),
    .A(\u_inv.d_next[232] ),
    .B(\u_inv.d_reg[232] ));
 sg13g2_xor2_1 _34116_ (.B(\u_inv.d_reg[232] ),
    .A(\u_inv.d_next[232] ),
    .X(_03528_));
 sg13g2_xnor2_1 _34117_ (.Y(_03529_),
    .A(\u_inv.d_next[232] ),
    .B(\u_inv.d_reg[232] ));
 sg13g2_nor2_1 _34118_ (.A(_03526_),
    .B(_03529_),
    .Y(_03530_));
 sg13g2_nand2_1 _34119_ (.Y(_03531_),
    .A(\u_inv.d_next[235] ),
    .B(\u_inv.d_reg[235] ));
 sg13g2_nor2_1 _34120_ (.A(\u_inv.d_next[235] ),
    .B(\u_inv.d_reg[235] ),
    .Y(_03532_));
 sg13g2_xor2_1 _34121_ (.B(\u_inv.d_reg[235] ),
    .A(\u_inv.d_next[235] ),
    .X(_03533_));
 sg13g2_xnor2_1 _34122_ (.Y(_03534_),
    .A(\u_inv.d_next[235] ),
    .B(\u_inv.d_reg[235] ));
 sg13g2_nand2_1 _34123_ (.Y(_03535_),
    .A(\u_inv.d_next[234] ),
    .B(\u_inv.d_reg[234] ));
 sg13g2_xnor2_1 _34124_ (.Y(_03536_),
    .A(\u_inv.d_next[234] ),
    .B(\u_inv.d_reg[234] ));
 sg13g2_nor2_1 _34125_ (.A(_03534_),
    .B(_03536_),
    .Y(_03537_));
 sg13g2_nand3_1 _34126_ (.B(_03530_),
    .C(_03537_),
    .A(_03522_),
    .Y(_03538_));
 sg13g2_xor2_1 _34127_ (.B(\u_inv.d_reg[227] ),
    .A(\u_inv.d_next[227] ),
    .X(_03539_));
 sg13g2_and2_1 _34128_ (.A(\u_inv.d_next[226] ),
    .B(\u_inv.d_reg[226] ),
    .X(_03540_));
 sg13g2_xor2_1 _34129_ (.B(\u_inv.d_reg[226] ),
    .A(\u_inv.d_next[226] ),
    .X(_03541_));
 sg13g2_and2_1 _34130_ (.A(_03539_),
    .B(_03541_),
    .X(_03542_));
 sg13g2_nor2_1 _34131_ (.A(\u_inv.d_next[229] ),
    .B(\u_inv.d_reg[229] ),
    .Y(_03543_));
 sg13g2_nand2_1 _34132_ (.Y(_03544_),
    .A(\u_inv.d_next[229] ),
    .B(\u_inv.d_reg[229] ));
 sg13g2_nor2b_1 _34133_ (.A(_03543_),
    .B_N(_03544_),
    .Y(_03545_));
 sg13g2_nand2b_2 _34134_ (.Y(_03546_),
    .B(_03544_),
    .A_N(_03543_));
 sg13g2_nand2_1 _34135_ (.Y(_03547_),
    .A(\u_inv.d_next[228] ),
    .B(\u_inv.d_reg[228] ));
 sg13g2_xor2_1 _34136_ (.B(\u_inv.d_reg[228] ),
    .A(\u_inv.d_next[228] ),
    .X(_03548_));
 sg13g2_xnor2_1 _34137_ (.Y(_03549_),
    .A(\u_inv.d_next[228] ),
    .B(\u_inv.d_reg[228] ));
 sg13g2_nor2_1 _34138_ (.A(_03546_),
    .B(_03549_),
    .Y(_03550_));
 sg13g2_nand2_1 _34139_ (.Y(_03551_),
    .A(\u_inv.d_next[230] ),
    .B(\u_inv.d_reg[230] ));
 sg13g2_xnor2_1 _34140_ (.Y(_03552_),
    .A(\u_inv.d_next[230] ),
    .B(\u_inv.d_reg[230] ));
 sg13g2_nand2_1 _34141_ (.Y(_03553_),
    .A(\u_inv.d_next[231] ),
    .B(\u_inv.d_reg[231] ));
 sg13g2_nor2_1 _34142_ (.A(\u_inv.d_next[231] ),
    .B(\u_inv.d_reg[231] ),
    .Y(_03554_));
 sg13g2_xnor2_1 _34143_ (.Y(_03555_),
    .A(\u_inv.d_next[231] ),
    .B(\u_inv.d_reg[231] ));
 sg13g2_nor2_1 _34144_ (.A(_03552_),
    .B(_03555_),
    .Y(_03556_));
 sg13g2_and2_1 _34145_ (.A(_03550_),
    .B(_03556_),
    .X(_03557_));
 sg13g2_xnor2_1 _34146_ (.Y(_03558_),
    .A(\u_inv.d_next[224] ),
    .B(\u_inv.d_reg[224] ));
 sg13g2_nor2_1 _34147_ (.A(\u_inv.d_next[225] ),
    .B(\u_inv.d_reg[225] ),
    .Y(_03559_));
 sg13g2_xnor2_1 _34148_ (.Y(_03560_),
    .A(\u_inv.d_next[225] ),
    .B(\u_inv.d_reg[225] ));
 sg13g2_nor2_1 _34149_ (.A(_03558_),
    .B(_03560_),
    .Y(_03561_));
 sg13g2_or2_1 _34150_ (.X(_03562_),
    .B(_03560_),
    .A(_03558_));
 sg13g2_nand3_1 _34151_ (.B(_03557_),
    .C(_03561_),
    .A(_03542_),
    .Y(_03563_));
 sg13g2_nor2_2 _34152_ (.A(_03538_),
    .B(_03563_),
    .Y(_03564_));
 sg13g2_inv_1 _34153_ (.Y(_03565_),
    .A(_03564_));
 sg13g2_xor2_1 _34154_ (.B(\u_inv.d_reg[255] ),
    .A(\u_inv.d_next[255] ),
    .X(_03566_));
 sg13g2_xnor2_1 _34155_ (.Y(_03567_),
    .A(\u_inv.d_next[255] ),
    .B(\u_inv.d_reg[255] ));
 sg13g2_nand2_1 _34156_ (.Y(_03568_),
    .A(\u_inv.d_next[254] ),
    .B(\u_inv.d_reg[254] ));
 sg13g2_nor2_1 _34157_ (.A(\u_inv.d_next[254] ),
    .B(\u_inv.d_reg[254] ),
    .Y(_03569_));
 sg13g2_xor2_1 _34158_ (.B(\u_inv.d_reg[254] ),
    .A(\u_inv.d_next[254] ),
    .X(_03570_));
 sg13g2_and2_1 _34159_ (.A(_03566_),
    .B(_03570_),
    .X(_03571_));
 sg13g2_nand2_1 _34160_ (.Y(_03572_),
    .A(\u_inv.d_next[253] ),
    .B(\u_inv.d_reg[253] ));
 sg13g2_nor2_1 _34161_ (.A(\u_inv.d_next[253] ),
    .B(\u_inv.d_reg[253] ),
    .Y(_03573_));
 sg13g2_xor2_1 _34162_ (.B(\u_inv.d_reg[253] ),
    .A(\u_inv.d_next[253] ),
    .X(_03574_));
 sg13g2_xnor2_1 _34163_ (.Y(_03575_),
    .A(\u_inv.d_next[253] ),
    .B(\u_inv.d_reg[253] ));
 sg13g2_nand2_1 _34164_ (.Y(_03576_),
    .A(\u_inv.d_next[252] ),
    .B(\u_inv.d_reg[252] ));
 sg13g2_xor2_1 _34165_ (.B(\u_inv.d_reg[252] ),
    .A(\u_inv.d_next[252] ),
    .X(_03577_));
 sg13g2_xnor2_1 _34166_ (.Y(_03578_),
    .A(\u_inv.d_next[252] ),
    .B(\u_inv.d_reg[252] ));
 sg13g2_nor2_1 _34167_ (.A(_03575_),
    .B(_03578_),
    .Y(_03579_));
 sg13g2_and2_1 _34168_ (.A(_03571_),
    .B(_03579_),
    .X(_03580_));
 sg13g2_nand2_1 _34169_ (.Y(_03581_),
    .A(\u_inv.d_next[249] ),
    .B(\u_inv.d_reg[249] ));
 sg13g2_nor2_1 _34170_ (.A(\u_inv.d_next[249] ),
    .B(\u_inv.d_reg[249] ),
    .Y(_03582_));
 sg13g2_xor2_1 _34171_ (.B(\u_inv.d_reg[249] ),
    .A(\u_inv.d_next[249] ),
    .X(_03583_));
 sg13g2_nand2_1 _34172_ (.Y(_03584_),
    .A(\u_inv.d_next[248] ),
    .B(\u_inv.d_reg[248] ));
 sg13g2_xor2_1 _34173_ (.B(\u_inv.d_reg[248] ),
    .A(\u_inv.d_next[248] ),
    .X(_03585_));
 sg13g2_xnor2_1 _34174_ (.Y(_03586_),
    .A(\u_inv.d_next[248] ),
    .B(\u_inv.d_reg[248] ));
 sg13g2_and2_1 _34175_ (.A(_03583_),
    .B(_03585_),
    .X(_03587_));
 sg13g2_inv_1 _34176_ (.Y(_03588_),
    .A(_03587_));
 sg13g2_xnor2_1 _34177_ (.Y(_03589_),
    .A(\u_inv.d_next[251] ),
    .B(\u_inv.d_reg[251] ));
 sg13g2_nand2_1 _34178_ (.Y(_03590_),
    .A(\u_inv.d_next[250] ),
    .B(\u_inv.d_reg[250] ));
 sg13g2_xnor2_1 _34179_ (.Y(_03591_),
    .A(\u_inv.d_next[250] ),
    .B(\u_inv.d_reg[250] ));
 sg13g2_nor2_2 _34180_ (.A(_03589_),
    .B(_03591_),
    .Y(_03592_));
 sg13g2_xor2_1 _34181_ (.B(\u_inv.d_reg[245] ),
    .A(net7295),
    .X(_03593_));
 sg13g2_xnor2_1 _34182_ (.Y(_03594_),
    .A(net7295),
    .B(\u_inv.d_reg[245] ));
 sg13g2_nand2_1 _34183_ (.Y(_03595_),
    .A(\u_inv.d_next[244] ),
    .B(\u_inv.d_reg[244] ));
 sg13g2_xor2_1 _34184_ (.B(\u_inv.d_reg[244] ),
    .A(\u_inv.d_next[244] ),
    .X(_03596_));
 sg13g2_and2_1 _34185_ (.A(_03593_),
    .B(_03596_),
    .X(_03597_));
 sg13g2_xor2_1 _34186_ (.B(net7287),
    .A(\u_inv.d_next[241] ),
    .X(_03598_));
 sg13g2_xnor2_1 _34187_ (.Y(_03599_),
    .A(\u_inv.d_next[241] ),
    .B(net7287));
 sg13g2_and2_1 _34188_ (.A(\u_inv.d_next[246] ),
    .B(\u_inv.d_reg[246] ),
    .X(_03600_));
 sg13g2_xor2_1 _34189_ (.B(\u_inv.d_reg[246] ),
    .A(\u_inv.d_next[246] ),
    .X(_03601_));
 sg13g2_inv_1 _34190_ (.Y(_03602_),
    .A(_03601_));
 sg13g2_xor2_1 _34191_ (.B(\u_inv.d_reg[247] ),
    .A(\u_inv.d_next[247] ),
    .X(_03603_));
 sg13g2_nand2_1 _34192_ (.Y(_03604_),
    .A(_03601_),
    .B(_03603_));
 sg13g2_or2_1 _34193_ (.X(_03605_),
    .B(\u_inv.d_reg[243] ),
    .A(\u_inv.d_next[243] ));
 sg13g2_nand2_1 _34194_ (.Y(_03606_),
    .A(\u_inv.d_next[243] ),
    .B(\u_inv.d_reg[243] ));
 sg13g2_and2_1 _34195_ (.A(_03605_),
    .B(_03606_),
    .X(_03607_));
 sg13g2_nand2_1 _34196_ (.Y(_03608_),
    .A(_03605_),
    .B(_03606_));
 sg13g2_xnor2_1 _34197_ (.Y(_03609_),
    .A(\u_inv.d_next[242] ),
    .B(\u_inv.d_reg[242] ));
 sg13g2_nor2_1 _34198_ (.A(_03608_),
    .B(_03609_),
    .Y(_03610_));
 sg13g2_or2_1 _34199_ (.X(_03611_),
    .B(_03609_),
    .A(_03608_));
 sg13g2_and4_1 _34200_ (.A(_03597_),
    .B(_03598_),
    .C(_03601_),
    .D(_03603_),
    .X(_03612_));
 sg13g2_nand2_1 _34201_ (.Y(_03613_),
    .A(_03610_),
    .B(_03612_));
 sg13g2_xor2_1 _34202_ (.B(net7288),
    .A(\u_inv.d_next[240] ),
    .X(_03614_));
 sg13g2_xnor2_1 _34203_ (.Y(_03615_),
    .A(\u_inv.d_next[240] ),
    .B(net7288));
 sg13g2_a21oi_1 _34204_ (.A1(\u_inv.d_next[247] ),
    .A2(\u_inv.d_reg[247] ),
    .Y(_03616_),
    .B1(_03600_));
 sg13g2_a21oi_1 _34205_ (.A1(_18103_),
    .A2(_18367_),
    .Y(_03617_),
    .B1(_03616_));
 sg13g2_a21oi_1 _34206_ (.A1(_18104_),
    .A2(_18369_),
    .Y(_03618_),
    .B1(_03595_));
 sg13g2_a21oi_1 _34207_ (.A1(net7295),
    .A2(\u_inv.d_reg[245] ),
    .Y(_03619_),
    .B1(_03618_));
 sg13g2_a22oi_1 _34208_ (.Y(_03620_),
    .B1(net7288),
    .B2(\u_inv.d_next[240] ),
    .A2(net7287),
    .A1(\u_inv.d_next[241] ));
 sg13g2_inv_1 _34209_ (.Y(_03621_),
    .A(_03620_));
 sg13g2_o21ai_1 _34210_ (.B1(_03621_),
    .Y(_03622_),
    .A1(\u_inv.d_next[241] ),
    .A2(net7287));
 sg13g2_nor2_1 _34211_ (.A(_03611_),
    .B(_03622_),
    .Y(_03623_));
 sg13g2_nand3_1 _34212_ (.B(\u_inv.d_reg[242] ),
    .C(_03605_),
    .A(\u_inv.d_next[242] ),
    .Y(_03624_));
 sg13g2_nand2_2 _34213_ (.Y(_03625_),
    .A(_03606_),
    .B(_03624_));
 sg13g2_o21ai_1 _34214_ (.B1(_03597_),
    .Y(_03626_),
    .A1(_03623_),
    .A2(_03625_));
 sg13g2_a21oi_1 _34215_ (.A1(_03619_),
    .A2(_03626_),
    .Y(_03627_),
    .B1(_03604_));
 sg13g2_or2_1 _34216_ (.X(_03628_),
    .B(_03627_),
    .A(_03617_));
 sg13g2_inv_1 _34217_ (.Y(_03629_),
    .A(_03628_));
 sg13g2_o21ai_1 _34218_ (.B1(_03581_),
    .Y(_03630_),
    .A1(_03582_),
    .A2(_03584_));
 sg13g2_a21oi_1 _34219_ (.A1(_18102_),
    .A2(_18363_),
    .Y(_03631_),
    .B1(_03590_));
 sg13g2_a221oi_1 _34220_ (.B2(_03630_),
    .C1(_03631_),
    .B1(_03592_),
    .A1(\u_inv.d_next[251] ),
    .Y(_03632_),
    .A2(\u_inv.d_reg[251] ));
 sg13g2_inv_1 _34221_ (.Y(_03633_),
    .A(_03632_));
 sg13g2_o21ai_1 _34222_ (.B1(_03572_),
    .Y(_03634_),
    .A1(_03573_),
    .A2(_03576_));
 sg13g2_a21oi_1 _34223_ (.A1(_18101_),
    .A2(_18359_),
    .Y(_03635_),
    .B1(_03568_));
 sg13g2_a22oi_1 _34224_ (.Y(_03636_),
    .B1(\u_inv.d_reg[224] ),
    .B2(\u_inv.d_next[224] ),
    .A2(\u_inv.d_reg[225] ),
    .A1(\u_inv.d_next[225] ));
 sg13g2_or2_1 _34225_ (.X(_03637_),
    .B(_03636_),
    .A(_03559_));
 sg13g2_o21ai_1 _34226_ (.B1(_03540_),
    .Y(_03638_),
    .A1(\u_inv.d_next[227] ),
    .A2(\u_inv.d_reg[227] ));
 sg13g2_o21ai_1 _34227_ (.B1(_03638_),
    .Y(_03639_),
    .A1(_18107_),
    .A2(_18387_));
 sg13g2_a21oi_1 _34228_ (.A1(_03551_),
    .A2(_03553_),
    .Y(_03640_),
    .B1(_03554_));
 sg13g2_o21ai_1 _34229_ (.B1(_03544_),
    .Y(_03641_),
    .A1(_03543_),
    .A2(_03547_));
 sg13g2_nand2b_1 _34230_ (.Y(_03642_),
    .B(_03542_),
    .A_N(_03637_));
 sg13g2_nand2b_1 _34231_ (.Y(_03643_),
    .B(_03642_),
    .A_N(_03639_));
 sg13g2_a221oi_1 _34232_ (.B2(_03557_),
    .C1(_03640_),
    .B1(_03643_),
    .A1(_03556_),
    .Y(_03644_),
    .A2(_03641_));
 sg13g2_o21ai_1 _34233_ (.B1(_03517_),
    .Y(_03645_),
    .A1(_03516_),
    .A2(_03519_));
 sg13g2_o21ai_1 _34234_ (.B1(_03510_),
    .Y(_03646_),
    .A1(_03509_),
    .A2(_03513_));
 sg13g2_o21ai_1 _34235_ (.B1(_03524_),
    .Y(_03647_),
    .A1(_03523_),
    .A2(_03527_));
 sg13g2_a21oi_1 _34236_ (.A1(_03531_),
    .A2(_03535_),
    .Y(_03648_),
    .B1(_03532_));
 sg13g2_a21o_1 _34237_ (.A2(_03647_),
    .A1(_03537_),
    .B1(_03648_),
    .X(_03649_));
 sg13g2_a221oi_1 _34238_ (.B2(_03522_),
    .C1(_03646_),
    .B1(_03649_),
    .A1(_03515_),
    .Y(_03650_),
    .A2(_03645_));
 sg13g2_o21ai_1 _34239_ (.B1(_03650_),
    .Y(_03651_),
    .A1(_03538_),
    .A2(_03644_));
 sg13g2_inv_1 _34240_ (.Y(_03652_),
    .A(_03651_));
 sg13g2_nand3_1 _34241_ (.B(_03587_),
    .C(_03592_),
    .A(_03580_),
    .Y(_03653_));
 sg13g2_nor3_1 _34242_ (.A(_03613_),
    .B(_03615_),
    .C(_03653_),
    .Y(_03654_));
 sg13g2_nand2_1 _34243_ (.Y(_03655_),
    .A(_03651_),
    .B(_03654_));
 sg13g2_nand2b_1 _34244_ (.Y(_03656_),
    .B(_03628_),
    .A_N(_03653_));
 sg13g2_a221oi_1 _34245_ (.B2(_03633_),
    .C1(_03635_),
    .B1(_03580_),
    .A1(\u_inv.d_next[255] ),
    .Y(_03657_),
    .A2(\u_inv.d_reg[255] ));
 sg13g2_nand3_1 _34246_ (.B(_03656_),
    .C(_03657_),
    .A(_03655_),
    .Y(_03658_));
 sg13g2_and2_1 _34247_ (.A(_03564_),
    .B(_03654_),
    .X(_03659_));
 sg13g2_a22oi_1 _34248_ (.Y(_03660_),
    .B1(_03659_),
    .B2(_03508_),
    .A2(_03634_),
    .A1(_03571_));
 sg13g2_nand2b_2 _34249_ (.Y(_03661_),
    .B(_03660_),
    .A_N(_03658_));
 sg13g2_nor2_1 _34250_ (.A(\u_inv.d_next[161] ),
    .B(_18453_),
    .Y(_03662_));
 sg13g2_nand2_1 _34251_ (.Y(_03663_),
    .A(\u_inv.d_next[161] ),
    .B(_18453_));
 sg13g2_nor2b_2 _34252_ (.A(_03662_),
    .B_N(_03663_),
    .Y(_03664_));
 sg13g2_nand2b_2 _34253_ (.Y(_03665_),
    .B(_03663_),
    .A_N(_03662_));
 sg13g2_nand2_1 _34254_ (.Y(_03666_),
    .A(\u_inv.d_next[160] ),
    .B(\u_inv.d_reg[160] ));
 sg13g2_xor2_1 _34255_ (.B(\u_inv.d_reg[160] ),
    .A(\u_inv.d_next[160] ),
    .X(_03667_));
 sg13g2_xnor2_1 _34256_ (.Y(_03668_),
    .A(\u_inv.d_next[160] ),
    .B(\u_inv.d_reg[160] ));
 sg13g2_xnor2_1 _34257_ (.Y(_03669_),
    .A(\u_inv.d_next[163] ),
    .B(\u_inv.d_reg[163] ));
 sg13g2_nand2_1 _34258_ (.Y(_03670_),
    .A(\u_inv.d_next[162] ),
    .B(\u_inv.d_reg[162] ));
 sg13g2_xnor2_1 _34259_ (.Y(_03671_),
    .A(\u_inv.d_next[162] ),
    .B(\u_inv.d_reg[162] ));
 sg13g2_nor2_1 _34260_ (.A(_03669_),
    .B(_03671_),
    .Y(_03672_));
 sg13g2_nand3_1 _34261_ (.B(_03667_),
    .C(_03672_),
    .A(_03665_),
    .Y(_03673_));
 sg13g2_xor2_1 _34262_ (.B(\u_inv.d_reg[175] ),
    .A(\u_inv.d_next[175] ),
    .X(_03674_));
 sg13g2_nor2_1 _34263_ (.A(\u_inv.d_next[174] ),
    .B(\u_inv.d_reg[174] ),
    .Y(_03675_));
 sg13g2_nand2_1 _34264_ (.Y(_03676_),
    .A(\u_inv.d_next[174] ),
    .B(\u_inv.d_reg[174] ));
 sg13g2_nor2b_2 _34265_ (.A(_03675_),
    .B_N(_03676_),
    .Y(_03677_));
 sg13g2_nand2_1 _34266_ (.Y(_03678_),
    .A(_03674_),
    .B(_03677_));
 sg13g2_inv_1 _34267_ (.Y(_03679_),
    .A(_03678_));
 sg13g2_nor2_1 _34268_ (.A(\u_inv.d_next[173] ),
    .B(\u_inv.d_reg[173] ),
    .Y(_03680_));
 sg13g2_nand2_1 _34269_ (.Y(_03681_),
    .A(\u_inv.d_next[173] ),
    .B(\u_inv.d_reg[173] ));
 sg13g2_nor2b_1 _34270_ (.A(_03680_),
    .B_N(_03681_),
    .Y(_03682_));
 sg13g2_nand2b_2 _34271_ (.Y(_03683_),
    .B(_03681_),
    .A_N(_03680_));
 sg13g2_nand2_1 _34272_ (.Y(_03684_),
    .A(\u_inv.d_next[172] ),
    .B(\u_inv.d_reg[172] ));
 sg13g2_xor2_1 _34273_ (.B(\u_inv.d_reg[172] ),
    .A(\u_inv.d_next[172] ),
    .X(_03685_));
 sg13g2_inv_1 _34274_ (.Y(_03686_),
    .A(_03685_));
 sg13g2_nor2_1 _34275_ (.A(_03683_),
    .B(_03686_),
    .Y(_03687_));
 sg13g2_nor2b_1 _34276_ (.A(_03678_),
    .B_N(_03687_),
    .Y(_03688_));
 sg13g2_xor2_1 _34277_ (.B(\u_inv.d_reg[169] ),
    .A(\u_inv.d_next[169] ),
    .X(_03689_));
 sg13g2_xnor2_1 _34278_ (.Y(_03690_),
    .A(\u_inv.d_next[169] ),
    .B(\u_inv.d_reg[169] ));
 sg13g2_xnor2_1 _34279_ (.Y(_03691_),
    .A(\u_inv.d_next[168] ),
    .B(\u_inv.d_reg[168] ));
 sg13g2_inv_2 _34280_ (.Y(_03692_),
    .A(_03691_));
 sg13g2_nor2_1 _34281_ (.A(_03690_),
    .B(_03691_),
    .Y(_03693_));
 sg13g2_nor2_1 _34282_ (.A(\u_inv.d_next[171] ),
    .B(\u_inv.d_reg[171] ),
    .Y(_03694_));
 sg13g2_nand2_1 _34283_ (.Y(_03695_),
    .A(\u_inv.d_next[171] ),
    .B(\u_inv.d_reg[171] ));
 sg13g2_nor2b_2 _34284_ (.A(_03694_),
    .B_N(_03695_),
    .Y(_03696_));
 sg13g2_nand2b_1 _34285_ (.Y(_03697_),
    .B(_03695_),
    .A_N(_03694_));
 sg13g2_nand2_1 _34286_ (.Y(_03698_),
    .A(\u_inv.d_next[170] ),
    .B(\u_inv.d_reg[170] ));
 sg13g2_xnor2_1 _34287_ (.Y(_03699_),
    .A(\u_inv.d_next[170] ),
    .B(\u_inv.d_reg[170] ));
 sg13g2_nor2_1 _34288_ (.A(_03697_),
    .B(_03699_),
    .Y(_03700_));
 sg13g2_nand2_1 _34289_ (.Y(_03701_),
    .A(_03693_),
    .B(_03700_));
 sg13g2_nand3_1 _34290_ (.B(_03693_),
    .C(_03700_),
    .A(_03688_),
    .Y(_03702_));
 sg13g2_inv_1 _34291_ (.Y(_03703_),
    .A(_03702_));
 sg13g2_nand2_1 _34292_ (.Y(_03704_),
    .A(\u_inv.d_next[164] ),
    .B(\u_inv.d_reg[164] ));
 sg13g2_xnor2_1 _34293_ (.Y(_03705_),
    .A(\u_inv.d_next[164] ),
    .B(\u_inv.d_reg[164] ));
 sg13g2_nand2_1 _34294_ (.Y(_03706_),
    .A(\u_inv.d_next[166] ),
    .B(\u_inv.d_reg[166] ));
 sg13g2_xor2_1 _34295_ (.B(\u_inv.d_reg[166] ),
    .A(\u_inv.d_next[166] ),
    .X(_03707_));
 sg13g2_xnor2_1 _34296_ (.Y(_03708_),
    .A(\u_inv.d_next[166] ),
    .B(\u_inv.d_reg[166] ));
 sg13g2_nor2_1 _34297_ (.A(\u_inv.d_next[167] ),
    .B(\u_inv.d_reg[167] ),
    .Y(_03709_));
 sg13g2_xor2_1 _34298_ (.B(\u_inv.d_reg[167] ),
    .A(\u_inv.d_next[167] ),
    .X(_03710_));
 sg13g2_xnor2_1 _34299_ (.Y(_03711_),
    .A(\u_inv.d_next[167] ),
    .B(\u_inv.d_reg[167] ));
 sg13g2_nor2_1 _34300_ (.A(_03708_),
    .B(_03711_),
    .Y(_03712_));
 sg13g2_xnor2_1 _34301_ (.Y(_03713_),
    .A(\u_inv.d_next[165] ),
    .B(\u_inv.d_reg[165] ));
 sg13g2_nor2_1 _34302_ (.A(_03705_),
    .B(_03713_),
    .Y(_03714_));
 sg13g2_nand2_2 _34303_ (.Y(_03715_),
    .A(_03712_),
    .B(_03714_));
 sg13g2_inv_1 _34304_ (.Y(_03716_),
    .A(_03715_));
 sg13g2_nor3_1 _34305_ (.A(_03673_),
    .B(_03702_),
    .C(_03715_),
    .Y(_03717_));
 sg13g2_and2_1 _34306_ (.A(\u_inv.d_next[182] ),
    .B(\u_inv.d_reg[182] ),
    .X(_03718_));
 sg13g2_xor2_1 _34307_ (.B(\u_inv.d_reg[182] ),
    .A(\u_inv.d_next[182] ),
    .X(_03719_));
 sg13g2_xor2_1 _34308_ (.B(\u_inv.d_reg[183] ),
    .A(\u_inv.d_next[183] ),
    .X(_03720_));
 sg13g2_and2_1 _34309_ (.A(_03719_),
    .B(_03720_),
    .X(_03721_));
 sg13g2_xor2_1 _34310_ (.B(\u_inv.d_reg[181] ),
    .A(\u_inv.d_next[181] ),
    .X(_03722_));
 sg13g2_and2_1 _34311_ (.A(\u_inv.d_next[180] ),
    .B(\u_inv.d_reg[180] ),
    .X(_03723_));
 sg13g2_xor2_1 _34312_ (.B(\u_inv.d_reg[180] ),
    .A(\u_inv.d_next[180] ),
    .X(_03724_));
 sg13g2_and2_1 _34313_ (.A(_03722_),
    .B(_03724_),
    .X(_03725_));
 sg13g2_nand2_1 _34314_ (.Y(_03726_),
    .A(\u_inv.d_next[178] ),
    .B(\u_inv.d_reg[178] ));
 sg13g2_xnor2_1 _34315_ (.Y(_03727_),
    .A(\u_inv.d_next[178] ),
    .B(\u_inv.d_reg[178] ));
 sg13g2_inv_2 _34316_ (.Y(_03728_),
    .A(_03727_));
 sg13g2_nor2_1 _34317_ (.A(\u_inv.d_next[179] ),
    .B(\u_inv.d_reg[179] ),
    .Y(_03729_));
 sg13g2_nand2_1 _34318_ (.Y(_03730_),
    .A(\u_inv.d_next[179] ),
    .B(\u_inv.d_reg[179] ));
 sg13g2_nor2b_1 _34319_ (.A(_03729_),
    .B_N(_03730_),
    .Y(_03731_));
 sg13g2_nand2b_2 _34320_ (.Y(_03732_),
    .B(_03730_),
    .A_N(_03729_));
 sg13g2_nor2_1 _34321_ (.A(_03727_),
    .B(_03732_),
    .Y(_03733_));
 sg13g2_inv_1 _34322_ (.Y(_03734_),
    .A(_03733_));
 sg13g2_xnor2_1 _34323_ (.Y(_03735_),
    .A(\u_inv.d_next[177] ),
    .B(\u_inv.d_reg[177] ));
 sg13g2_nand2_1 _34324_ (.Y(_03736_),
    .A(\u_inv.d_next[176] ),
    .B(\u_inv.d_reg[176] ));
 sg13g2_xnor2_1 _34325_ (.Y(_03737_),
    .A(\u_inv.d_next[176] ),
    .B(\u_inv.d_reg[176] ));
 sg13g2_nor2_1 _34326_ (.A(_03735_),
    .B(_03737_),
    .Y(_03738_));
 sg13g2_nand4_1 _34327_ (.B(_03725_),
    .C(_03733_),
    .A(_03721_),
    .Y(_03739_),
    .D(_03738_));
 sg13g2_nand2_1 _34328_ (.Y(_03740_),
    .A(\u_inv.d_next[191] ),
    .B(\u_inv.d_reg[191] ));
 sg13g2_nor2_1 _34329_ (.A(\u_inv.d_next[191] ),
    .B(\u_inv.d_reg[191] ),
    .Y(_03741_));
 sg13g2_xor2_1 _34330_ (.B(\u_inv.d_reg[191] ),
    .A(\u_inv.d_next[191] ),
    .X(_03742_));
 sg13g2_xnor2_1 _34331_ (.Y(_03743_),
    .A(\u_inv.d_next[191] ),
    .B(\u_inv.d_reg[191] ));
 sg13g2_nand2_1 _34332_ (.Y(_03744_),
    .A(\u_inv.d_next[190] ),
    .B(\u_inv.d_reg[190] ));
 sg13g2_xnor2_1 _34333_ (.Y(_03745_),
    .A(\u_inv.d_next[190] ),
    .B(\u_inv.d_reg[190] ));
 sg13g2_inv_1 _34334_ (.Y(_03746_),
    .A(_03745_));
 sg13g2_nor2_1 _34335_ (.A(_03743_),
    .B(_03745_),
    .Y(_03747_));
 sg13g2_nand2_1 _34336_ (.Y(_03748_),
    .A(\u_inv.d_next[189] ),
    .B(\u_inv.d_reg[189] ));
 sg13g2_nor2_1 _34337_ (.A(\u_inv.d_next[189] ),
    .B(\u_inv.d_reg[189] ),
    .Y(_03749_));
 sg13g2_xnor2_1 _34338_ (.Y(_03750_),
    .A(\u_inv.d_next[189] ),
    .B(\u_inv.d_reg[189] ));
 sg13g2_nand2_1 _34339_ (.Y(_03751_),
    .A(\u_inv.d_next[188] ),
    .B(\u_inv.d_reg[188] ));
 sg13g2_xnor2_1 _34340_ (.Y(_03752_),
    .A(\u_inv.d_next[188] ),
    .B(\u_inv.d_reg[188] ));
 sg13g2_nor2_1 _34341_ (.A(_03750_),
    .B(_03752_),
    .Y(_03753_));
 sg13g2_and2_1 _34342_ (.A(_03747_),
    .B(_03753_),
    .X(_03754_));
 sg13g2_nor2_1 _34343_ (.A(\u_inv.d_next[187] ),
    .B(\u_inv.d_reg[187] ),
    .Y(_03755_));
 sg13g2_nand2_1 _34344_ (.Y(_03756_),
    .A(\u_inv.d_next[187] ),
    .B(\u_inv.d_reg[187] ));
 sg13g2_nand2b_2 _34345_ (.Y(_03757_),
    .B(_03756_),
    .A_N(_03755_));
 sg13g2_inv_2 _34346_ (.Y(_03758_),
    .A(_03757_));
 sg13g2_nand2_1 _34347_ (.Y(_03759_),
    .A(\u_inv.d_next[186] ),
    .B(\u_inv.d_reg[186] ));
 sg13g2_xnor2_1 _34348_ (.Y(_03760_),
    .A(\u_inv.d_next[186] ),
    .B(\u_inv.d_reg[186] ));
 sg13g2_nor2_1 _34349_ (.A(_03757_),
    .B(_03760_),
    .Y(_03761_));
 sg13g2_xor2_1 _34350_ (.B(\u_inv.d_reg[185] ),
    .A(\u_inv.d_next[185] ),
    .X(_03762_));
 sg13g2_xnor2_1 _34351_ (.Y(_03763_),
    .A(\u_inv.d_next[185] ),
    .B(\u_inv.d_reg[185] ));
 sg13g2_and2_1 _34352_ (.A(\u_inv.d_next[184] ),
    .B(\u_inv.d_reg[184] ),
    .X(_03764_));
 sg13g2_xor2_1 _34353_ (.B(\u_inv.d_reg[184] ),
    .A(\u_inv.d_next[184] ),
    .X(_03765_));
 sg13g2_and2_1 _34354_ (.A(_03762_),
    .B(_03765_),
    .X(_03766_));
 sg13g2_a21oi_1 _34355_ (.A1(\u_inv.d_next[183] ),
    .A2(\u_inv.d_reg[183] ),
    .Y(_03767_),
    .B1(_03718_));
 sg13g2_a21oi_1 _34356_ (.A1(_18118_),
    .A2(_18431_),
    .Y(_03768_),
    .B1(_03767_));
 sg13g2_a21oi_1 _34357_ (.A1(\u_inv.d_next[181] ),
    .A2(\u_inv.d_reg[181] ),
    .Y(_03769_),
    .B1(_03723_));
 sg13g2_a21oi_1 _34358_ (.A1(_18119_),
    .A2(_18433_),
    .Y(_03770_),
    .B1(_03769_));
 sg13g2_a22oi_1 _34359_ (.Y(_03771_),
    .B1(\u_inv.d_reg[176] ),
    .B2(\u_inv.d_next[176] ),
    .A2(\u_inv.d_reg[177] ),
    .A1(\u_inv.d_next[177] ));
 sg13g2_a21oi_1 _34360_ (.A1(_18121_),
    .A2(_18437_),
    .Y(_03772_),
    .B1(_03771_));
 sg13g2_a21oi_1 _34361_ (.A1(_03726_),
    .A2(_03730_),
    .Y(_03773_),
    .B1(_03729_));
 sg13g2_inv_1 _34362_ (.Y(_03774_),
    .A(_03773_));
 sg13g2_a21oi_1 _34363_ (.A1(_03733_),
    .A2(_03772_),
    .Y(_03775_),
    .B1(_03773_));
 sg13g2_nor2b_1 _34364_ (.A(_03775_),
    .B_N(_03725_),
    .Y(_03776_));
 sg13g2_o21ai_1 _34365_ (.B1(_03721_),
    .Y(_03777_),
    .A1(_03770_),
    .A2(_03776_));
 sg13g2_nor2b_1 _34366_ (.A(_03768_),
    .B_N(_03777_),
    .Y(_03778_));
 sg13g2_a21oi_1 _34367_ (.A1(\u_inv.d_next[185] ),
    .A2(\u_inv.d_reg[185] ),
    .Y(_03779_),
    .B1(_03764_));
 sg13g2_a21oi_1 _34368_ (.A1(_18117_),
    .A2(_18429_),
    .Y(_03780_),
    .B1(_03779_));
 sg13g2_a21oi_1 _34369_ (.A1(_03756_),
    .A2(_03759_),
    .Y(_03781_),
    .B1(_03755_));
 sg13g2_a21o_1 _34370_ (.A2(_03780_),
    .A1(_03761_),
    .B1(_03781_),
    .X(_03782_));
 sg13g2_o21ai_1 _34371_ (.B1(_03748_),
    .Y(_03783_),
    .A1(_03749_),
    .A2(_03751_));
 sg13g2_o21ai_1 _34372_ (.B1(_03740_),
    .Y(_03784_),
    .A1(_03741_),
    .A2(_03744_));
 sg13g2_a221oi_1 _34373_ (.B2(_03747_),
    .C1(_03784_),
    .B1(_03783_),
    .A1(_03754_),
    .Y(_03785_),
    .A2(_03782_));
 sg13g2_nand2_1 _34374_ (.Y(_03786_),
    .A(\u_inv.d_next[161] ),
    .B(\u_inv.d_reg[161] ));
 sg13g2_o21ai_1 _34375_ (.B1(_03786_),
    .Y(_03787_),
    .A1(_03664_),
    .A2(_03666_));
 sg13g2_a21oi_1 _34376_ (.A1(_18125_),
    .A2(_18451_),
    .Y(_03788_),
    .B1(_03670_));
 sg13g2_a221oi_1 _34377_ (.B2(_03787_),
    .C1(_03788_),
    .B1(_03672_),
    .A1(\u_inv.d_next[163] ),
    .Y(_03789_),
    .A2(\u_inv.d_reg[163] ));
 sg13g2_o21ai_1 _34378_ (.B1(_03681_),
    .Y(_03790_),
    .A1(_03680_),
    .A2(_03684_));
 sg13g2_a21oi_1 _34379_ (.A1(_18122_),
    .A2(_18439_),
    .Y(_03791_),
    .B1(_03676_));
 sg13g2_a221oi_1 _34380_ (.B2(_03790_),
    .C1(_03791_),
    .B1(_03679_),
    .A1(\u_inv.d_next[175] ),
    .Y(_03792_),
    .A2(\u_inv.d_reg[175] ));
 sg13g2_a22oi_1 _34381_ (.Y(_03793_),
    .B1(\u_inv.d_reg[168] ),
    .B2(\u_inv.d_next[168] ),
    .A2(\u_inv.d_reg[169] ),
    .A1(\u_inv.d_next[169] ));
 sg13g2_inv_1 _34382_ (.Y(_03794_),
    .A(_03793_));
 sg13g2_o21ai_1 _34383_ (.B1(_03794_),
    .Y(_03795_),
    .A1(\u_inv.d_next[169] ),
    .A2(\u_inv.d_reg[169] ));
 sg13g2_nor3_1 _34384_ (.A(_03697_),
    .B(_03699_),
    .C(_03795_),
    .Y(_03796_));
 sg13g2_o21ai_1 _34385_ (.B1(_03695_),
    .Y(_03797_),
    .A1(_03694_),
    .A2(_03698_));
 sg13g2_nor2_1 _34386_ (.A(_03796_),
    .B(_03797_),
    .Y(_03798_));
 sg13g2_o21ai_1 _34387_ (.B1(_03688_),
    .Y(_03799_),
    .A1(_03796_),
    .A2(_03797_));
 sg13g2_o21ai_1 _34388_ (.B1(_03704_),
    .Y(_03800_),
    .A1(_18124_),
    .A2(_18449_));
 sg13g2_o21ai_1 _34389_ (.B1(_03800_),
    .Y(_03801_),
    .A1(\u_inv.d_next[165] ),
    .A2(\u_inv.d_reg[165] ));
 sg13g2_inv_1 _34390_ (.Y(_03802_),
    .A(_03801_));
 sg13g2_a22oi_1 _34391_ (.Y(_03803_),
    .B1(_03712_),
    .B2(_03802_),
    .A2(\u_inv.d_reg[167] ),
    .A1(\u_inv.d_next[167] ));
 sg13g2_o21ai_1 _34392_ (.B1(_03803_),
    .Y(_03804_),
    .A1(_03706_),
    .A2(_03709_));
 sg13g2_nor2_1 _34393_ (.A(_03715_),
    .B(_03789_),
    .Y(_03805_));
 sg13g2_o21ai_1 _34394_ (.B1(_03703_),
    .Y(_03806_),
    .A1(_03804_),
    .A2(_03805_));
 sg13g2_nand3_1 _34395_ (.B(_03799_),
    .C(_03806_),
    .A(_03792_),
    .Y(_03807_));
 sg13g2_nand2_1 _34396_ (.Y(_03808_),
    .A(\u_inv.d_next[127] ),
    .B(\u_inv.d_reg[127] ));
 sg13g2_nor2_1 _34397_ (.A(\u_inv.d_next[127] ),
    .B(\u_inv.d_reg[127] ),
    .Y(_03809_));
 sg13g2_xor2_1 _34398_ (.B(\u_inv.d_reg[127] ),
    .A(\u_inv.d_next[127] ),
    .X(_03810_));
 sg13g2_xnor2_1 _34399_ (.Y(_03811_),
    .A(\u_inv.d_next[127] ),
    .B(\u_inv.d_reg[127] ));
 sg13g2_nand2_1 _34400_ (.Y(_03812_),
    .A(\u_inv.d_next[126] ),
    .B(\u_inv.d_reg[126] ));
 sg13g2_xor2_1 _34401_ (.B(\u_inv.d_reg[126] ),
    .A(\u_inv.d_next[126] ),
    .X(_03813_));
 sg13g2_xor2_1 _34402_ (.B(\u_inv.d_reg[125] ),
    .A(\u_inv.d_next[125] ),
    .X(_03814_));
 sg13g2_xnor2_1 _34403_ (.Y(_03815_),
    .A(\u_inv.d_next[125] ),
    .B(\u_inv.d_reg[125] ));
 sg13g2_and2_1 _34404_ (.A(\u_inv.d_next[124] ),
    .B(\u_inv.d_reg[124] ),
    .X(_03816_));
 sg13g2_xor2_1 _34405_ (.B(\u_inv.d_reg[124] ),
    .A(\u_inv.d_next[124] ),
    .X(_03817_));
 sg13g2_and2_1 _34406_ (.A(_03814_),
    .B(_03817_),
    .X(_03818_));
 sg13g2_nand3_1 _34407_ (.B(_03813_),
    .C(_03818_),
    .A(_03810_),
    .Y(_03819_));
 sg13g2_xor2_1 _34408_ (.B(\u_inv.d_reg[123] ),
    .A(\u_inv.d_next[123] ),
    .X(_03820_));
 sg13g2_nand2_1 _34409_ (.Y(_03821_),
    .A(\u_inv.d_next[122] ),
    .B(\u_inv.d_reg[122] ));
 sg13g2_nor2_1 _34410_ (.A(\u_inv.d_next[122] ),
    .B(\u_inv.d_reg[122] ),
    .Y(_03822_));
 sg13g2_xor2_1 _34411_ (.B(\u_inv.d_reg[122] ),
    .A(\u_inv.d_next[122] ),
    .X(_03823_));
 sg13g2_nand2_1 _34412_ (.Y(_03824_),
    .A(_03820_),
    .B(_03823_));
 sg13g2_nand2b_1 _34413_ (.Y(_03825_),
    .B(\u_inv.d_reg[121] ),
    .A_N(\u_inv.d_next[121] ));
 sg13g2_nor2b_1 _34414_ (.A(\u_inv.d_reg[121] ),
    .B_N(\u_inv.d_next[121] ),
    .Y(_03826_));
 sg13g2_xnor2_1 _34415_ (.Y(_03827_),
    .A(\u_inv.d_next[121] ),
    .B(\u_inv.d_reg[121] ));
 sg13g2_nand2_1 _34416_ (.Y(_03828_),
    .A(\u_inv.d_next[120] ),
    .B(\u_inv.d_reg[120] ));
 sg13g2_nand2_1 _34417_ (.Y(_03829_),
    .A(\u_inv.d_next[121] ),
    .B(\u_inv.d_reg[121] ));
 sg13g2_o21ai_1 _34418_ (.B1(_03829_),
    .Y(_03830_),
    .A1(_03827_),
    .A2(_03828_));
 sg13g2_nand2b_1 _34419_ (.Y(_03831_),
    .B(_03830_),
    .A_N(_03824_));
 sg13g2_a21oi_1 _34420_ (.A1(_18138_),
    .A2(_18491_),
    .Y(_03832_),
    .B1(_03821_));
 sg13g2_a21oi_1 _34421_ (.A1(\u_inv.d_next[123] ),
    .A2(\u_inv.d_reg[123] ),
    .Y(_03833_),
    .B1(_03832_));
 sg13g2_a21oi_1 _34422_ (.A1(_03831_),
    .A2(_03833_),
    .Y(_03834_),
    .B1(_03819_));
 sg13g2_a21oi_1 _34423_ (.A1(\u_inv.d_next[125] ),
    .A2(\u_inv.d_reg[125] ),
    .Y(_03835_),
    .B1(_03816_));
 sg13g2_a21oi_1 _34424_ (.A1(_18137_),
    .A2(_18489_),
    .Y(_03836_),
    .B1(_03835_));
 sg13g2_and3_1 _34425_ (.X(_03837_),
    .A(_03810_),
    .B(_03813_),
    .C(_03836_));
 sg13g2_o21ai_1 _34426_ (.B1(_03808_),
    .Y(_03838_),
    .A1(_03809_),
    .A2(_03812_));
 sg13g2_nor3_1 _34427_ (.A(_03834_),
    .B(_03837_),
    .C(_03838_),
    .Y(_03839_));
 sg13g2_nor2_1 _34428_ (.A(\u_inv.d_next[119] ),
    .B(\u_inv.d_reg[119] ),
    .Y(_03840_));
 sg13g2_nand2_1 _34429_ (.Y(_03841_),
    .A(\u_inv.d_next[119] ),
    .B(\u_inv.d_reg[119] ));
 sg13g2_nor2b_2 _34430_ (.A(_03840_),
    .B_N(_03841_),
    .Y(_03842_));
 sg13g2_nand2b_2 _34431_ (.Y(_03843_),
    .B(_03841_),
    .A_N(_03840_));
 sg13g2_nand2_1 _34432_ (.Y(_03844_),
    .A(\u_inv.d_next[118] ),
    .B(\u_inv.d_reg[118] ));
 sg13g2_xor2_1 _34433_ (.B(\u_inv.d_reg[118] ),
    .A(\u_inv.d_next[118] ),
    .X(_03845_));
 sg13g2_inv_1 _34434_ (.Y(_03846_),
    .A(_03845_));
 sg13g2_nor2b_2 _34435_ (.A(\u_inv.d_next[117] ),
    .B_N(\u_inv.d_reg[117] ),
    .Y(_03847_));
 sg13g2_nand2b_1 _34436_ (.Y(_03848_),
    .B(\u_inv.d_next[117] ),
    .A_N(\u_inv.d_reg[117] ));
 sg13g2_nor2b_2 _34437_ (.A(_03847_),
    .B_N(_03848_),
    .Y(_03849_));
 sg13g2_nand2b_1 _34438_ (.Y(_03850_),
    .B(_03848_),
    .A_N(_03847_));
 sg13g2_nand2_1 _34439_ (.Y(_03851_),
    .A(\u_inv.d_next[116] ),
    .B(\u_inv.d_reg[116] ));
 sg13g2_xor2_1 _34440_ (.B(\u_inv.d_reg[116] ),
    .A(\u_inv.d_next[116] ),
    .X(_03852_));
 sg13g2_and2_1 _34441_ (.A(_03850_),
    .B(_03852_),
    .X(_03853_));
 sg13g2_nand3_1 _34442_ (.B(_03845_),
    .C(_03853_),
    .A(_03842_),
    .Y(_03854_));
 sg13g2_xnor2_1 _34443_ (.Y(_03855_),
    .A(\u_inv.d_next[115] ),
    .B(\u_inv.d_reg[115] ));
 sg13g2_nand2_1 _34444_ (.Y(_03856_),
    .A(\u_inv.d_next[112] ),
    .B(\u_inv.d_reg[112] ));
 sg13g2_nor2_1 _34445_ (.A(\u_inv.d_next[113] ),
    .B(_18501_),
    .Y(_03857_));
 sg13g2_nand2_1 _34446_ (.Y(_03858_),
    .A(\u_inv.d_next[113] ),
    .B(_18501_));
 sg13g2_xor2_1 _34447_ (.B(\u_inv.d_reg[113] ),
    .A(\u_inv.d_next[113] ),
    .X(_03859_));
 sg13g2_nand2b_1 _34448_ (.Y(_03860_),
    .B(_03859_),
    .A_N(_03856_));
 sg13g2_nand2_1 _34449_ (.Y(_03861_),
    .A(\u_inv.d_next[113] ),
    .B(\u_inv.d_reg[113] ));
 sg13g2_and2_1 _34450_ (.A(_03860_),
    .B(_03861_),
    .X(_03862_));
 sg13g2_nand3b_1 _34451_ (.B(\u_inv.d_reg[114] ),
    .C(\u_inv.d_next[114] ),
    .Y(_03863_),
    .A_N(_03855_));
 sg13g2_xnor2_1 _34452_ (.Y(_03864_),
    .A(\u_inv.d_next[114] ),
    .B(\u_inv.d_reg[114] ));
 sg13g2_or2_1 _34453_ (.X(_03865_),
    .B(_03864_),
    .A(_03855_));
 sg13g2_o21ai_1 _34454_ (.B1(_03863_),
    .Y(_03866_),
    .A1(_03862_),
    .A2(_03865_));
 sg13g2_a21oi_1 _34455_ (.A1(\u_inv.d_next[115] ),
    .A2(\u_inv.d_reg[115] ),
    .Y(_03867_),
    .B1(_03866_));
 sg13g2_o21ai_1 _34456_ (.B1(_03841_),
    .Y(_03868_),
    .A1(_03840_),
    .A2(_03844_));
 sg13g2_nand2_1 _34457_ (.Y(_03869_),
    .A(\u_inv.d_next[117] ),
    .B(\u_inv.d_reg[117] ));
 sg13g2_o21ai_1 _34458_ (.B1(_03869_),
    .Y(_03870_),
    .A1(_03849_),
    .A2(_03851_));
 sg13g2_nand3_1 _34459_ (.B(_03845_),
    .C(_03870_),
    .A(_03842_),
    .Y(_03871_));
 sg13g2_o21ai_1 _34460_ (.B1(_03871_),
    .Y(_03872_),
    .A1(_03854_),
    .A2(_03867_));
 sg13g2_nor2_1 _34461_ (.A(_03868_),
    .B(_03872_),
    .Y(_03873_));
 sg13g2_xnor2_1 _34462_ (.Y(_03874_),
    .A(\u_inv.d_next[120] ),
    .B(\u_inv.d_reg[120] ));
 sg13g2_inv_1 _34463_ (.Y(_03875_),
    .A(_03874_));
 sg13g2_nor2_1 _34464_ (.A(_03827_),
    .B(_03874_),
    .Y(_03876_));
 sg13g2_xor2_1 _34465_ (.B(\u_inv.d_reg[111] ),
    .A(\u_inv.d_next[111] ),
    .X(_03877_));
 sg13g2_xnor2_1 _34466_ (.Y(_03878_),
    .A(\u_inv.d_next[111] ),
    .B(\u_inv.d_reg[111] ));
 sg13g2_nand2_1 _34467_ (.Y(_03879_),
    .A(\u_inv.d_next[110] ),
    .B(\u_inv.d_reg[110] ));
 sg13g2_xor2_1 _34468_ (.B(\u_inv.d_reg[110] ),
    .A(\u_inv.d_next[110] ),
    .X(_03880_));
 sg13g2_nand2_1 _34469_ (.Y(_03881_),
    .A(_03877_),
    .B(_03880_));
 sg13g2_nand2_1 _34470_ (.Y(_03882_),
    .A(\u_inv.d_next[108] ),
    .B(\u_inv.d_reg[108] ));
 sg13g2_xor2_1 _34471_ (.B(\u_inv.d_reg[108] ),
    .A(\u_inv.d_next[108] ),
    .X(_03883_));
 sg13g2_xnor2_1 _34472_ (.Y(_03884_),
    .A(\u_inv.d_next[108] ),
    .B(\u_inv.d_reg[108] ));
 sg13g2_nor2_1 _34473_ (.A(\u_inv.d_next[109] ),
    .B(_18505_),
    .Y(_03885_));
 sg13g2_nand2_1 _34474_ (.Y(_03886_),
    .A(\u_inv.d_next[109] ),
    .B(_18505_));
 sg13g2_xnor2_1 _34475_ (.Y(_03887_),
    .A(\u_inv.d_next[109] ),
    .B(\u_inv.d_reg[109] ));
 sg13g2_nand2b_1 _34476_ (.Y(_03888_),
    .B(_03886_),
    .A_N(_03885_));
 sg13g2_nor3_1 _34477_ (.A(_03881_),
    .B(_03884_),
    .C(_03887_),
    .Y(_03889_));
 sg13g2_nor2_1 _34478_ (.A(\u_inv.d_next[107] ),
    .B(_18507_),
    .Y(_03890_));
 sg13g2_xnor2_1 _34479_ (.Y(_03891_),
    .A(\u_inv.d_next[107] ),
    .B(\u_inv.d_reg[107] ));
 sg13g2_inv_2 _34480_ (.Y(_03892_),
    .A(_03891_));
 sg13g2_xnor2_1 _34481_ (.Y(_03893_),
    .A(\u_inv.d_next[106] ),
    .B(\u_inv.d_reg[106] ));
 sg13g2_inv_1 _34482_ (.Y(_03894_),
    .A(_03893_));
 sg13g2_nor2_1 _34483_ (.A(_03891_),
    .B(_03893_),
    .Y(_03895_));
 sg13g2_xor2_1 _34484_ (.B(\u_inv.d_reg[105] ),
    .A(\u_inv.d_next[105] ),
    .X(_03896_));
 sg13g2_and2_1 _34485_ (.A(\u_inv.d_next[104] ),
    .B(\u_inv.d_reg[104] ),
    .X(_03897_));
 sg13g2_xor2_1 _34486_ (.B(\u_inv.d_reg[104] ),
    .A(\u_inv.d_next[104] ),
    .X(_03898_));
 sg13g2_xnor2_1 _34487_ (.Y(_03899_),
    .A(\u_inv.d_next[104] ),
    .B(\u_inv.d_reg[104] ));
 sg13g2_nand2_1 _34488_ (.Y(_03900_),
    .A(_03896_),
    .B(_03898_));
 sg13g2_and4_1 _34489_ (.A(_03889_),
    .B(_03895_),
    .C(_03896_),
    .D(_03898_),
    .X(_03901_));
 sg13g2_inv_1 _34490_ (.Y(_03902_),
    .A(_03901_));
 sg13g2_nand2_1 _34491_ (.Y(_03903_),
    .A(\u_inv.d_next[100] ),
    .B(\u_inv.d_reg[100] ));
 sg13g2_xnor2_1 _34492_ (.Y(_03904_),
    .A(\u_inv.d_next[100] ),
    .B(\u_inv.d_reg[100] ));
 sg13g2_nor2_1 _34493_ (.A(\u_inv.d_next[101] ),
    .B(\u_inv.d_reg[101] ),
    .Y(_03905_));
 sg13g2_nand2_1 _34494_ (.Y(_03906_),
    .A(\u_inv.d_next[101] ),
    .B(\u_inv.d_reg[101] ));
 sg13g2_xor2_1 _34495_ (.B(\u_inv.d_reg[101] ),
    .A(\u_inv.d_next[101] ),
    .X(_03907_));
 sg13g2_inv_1 _34496_ (.Y(_03908_),
    .A(_03907_));
 sg13g2_nand2b_1 _34497_ (.Y(_03909_),
    .B(_03907_),
    .A_N(_03904_));
 sg13g2_nor2_1 _34498_ (.A(\u_inv.d_next[102] ),
    .B(\u_inv.d_reg[102] ),
    .Y(_03910_));
 sg13g2_xnor2_1 _34499_ (.Y(_03911_),
    .A(\u_inv.d_next[102] ),
    .B(\u_inv.d_reg[102] ));
 sg13g2_nand2b_1 _34500_ (.Y(_03912_),
    .B(\u_inv.d_reg[103] ),
    .A_N(\u_inv.d_next[103] ));
 sg13g2_xnor2_1 _34501_ (.Y(_03913_),
    .A(\u_inv.d_next[103] ),
    .B(\u_inv.d_reg[103] ));
 sg13g2_nor3_1 _34502_ (.A(_03909_),
    .B(_03911_),
    .C(_03913_),
    .Y(_03914_));
 sg13g2_nand2b_1 _34503_ (.Y(_03915_),
    .B(\u_inv.d_reg[99] ),
    .A_N(\u_inv.d_next[99] ));
 sg13g2_nor2b_1 _34504_ (.A(\u_inv.d_reg[99] ),
    .B_N(\u_inv.d_next[99] ),
    .Y(_03916_));
 sg13g2_xnor2_1 _34505_ (.Y(_03917_),
    .A(\u_inv.d_next[99] ),
    .B(\u_inv.d_reg[99] ));
 sg13g2_xor2_1 _34506_ (.B(\u_inv.d_reg[99] ),
    .A(\u_inv.d_next[99] ),
    .X(_03918_));
 sg13g2_nand2_1 _34507_ (.Y(_03919_),
    .A(\u_inv.d_next[98] ),
    .B(\u_inv.d_reg[98] ));
 sg13g2_or2_1 _34508_ (.X(_03920_),
    .B(\u_inv.d_reg[98] ),
    .A(\u_inv.d_next[98] ));
 sg13g2_nand2b_1 _34509_ (.Y(_03921_),
    .B(\u_inv.d_reg[97] ),
    .A_N(\u_inv.d_next[97] ));
 sg13g2_nor2b_1 _34510_ (.A(\u_inv.d_reg[97] ),
    .B_N(\u_inv.d_next[97] ),
    .Y(_03922_));
 sg13g2_xnor2_1 _34511_ (.Y(_03923_),
    .A(\u_inv.d_next[97] ),
    .B(\u_inv.d_reg[97] ));
 sg13g2_xor2_1 _34512_ (.B(\u_inv.d_reg[97] ),
    .A(\u_inv.d_next[97] ),
    .X(_03924_));
 sg13g2_nand2_1 _34513_ (.Y(_03925_),
    .A(\u_inv.d_next[96] ),
    .B(\u_inv.d_reg[96] ));
 sg13g2_nand2_1 _34514_ (.Y(_03926_),
    .A(\u_inv.d_next[97] ),
    .B(\u_inv.d_reg[97] ));
 sg13g2_o21ai_1 _34515_ (.B1(_03926_),
    .Y(_03927_),
    .A1(_03923_),
    .A2(_03925_));
 sg13g2_nor2_1 _34516_ (.A(_03917_),
    .B(_03919_),
    .Y(_03928_));
 sg13g2_xnor2_1 _34517_ (.Y(_03929_),
    .A(\u_inv.d_next[98] ),
    .B(\u_inv.d_reg[98] ));
 sg13g2_nor2_2 _34518_ (.A(_03917_),
    .B(_03929_),
    .Y(_03930_));
 sg13g2_a221oi_1 _34519_ (.B2(_03930_),
    .C1(_03928_),
    .B1(_03927_),
    .A1(\u_inv.d_next[99] ),
    .Y(_03931_),
    .A2(\u_inv.d_reg[99] ));
 sg13g2_inv_1 _34520_ (.Y(_03932_),
    .A(_03931_));
 sg13g2_o21ai_1 _34521_ (.B1(_03906_),
    .Y(_03933_),
    .A1(_03903_),
    .A2(_03905_));
 sg13g2_a21oi_1 _34522_ (.A1(\u_inv.d_next[102] ),
    .A2(\u_inv.d_reg[102] ),
    .Y(_03934_),
    .B1(_03933_));
 sg13g2_nor3_1 _34523_ (.A(_03910_),
    .B(_03913_),
    .C(_03934_),
    .Y(_03935_));
 sg13g2_a221oi_1 _34524_ (.B2(_03932_),
    .C1(_03935_),
    .B1(_03914_),
    .A1(\u_inv.d_next[103] ),
    .Y(_03936_),
    .A2(\u_inv.d_reg[103] ));
 sg13g2_and2_1 _34525_ (.A(\u_inv.d_next[105] ),
    .B(\u_inv.d_reg[105] ),
    .X(_03937_));
 sg13g2_a21o_1 _34526_ (.A2(_03897_),
    .A1(_03896_),
    .B1(_03937_),
    .X(_03938_));
 sg13g2_a21oi_1 _34527_ (.A1(\u_inv.d_next[106] ),
    .A2(\u_inv.d_reg[106] ),
    .Y(_03939_),
    .B1(_03938_));
 sg13g2_o21ai_1 _34528_ (.B1(_03892_),
    .Y(_03940_),
    .A1(\u_inv.d_next[106] ),
    .A2(\u_inv.d_reg[106] ));
 sg13g2_nand2_1 _34529_ (.Y(_03941_),
    .A(\u_inv.d_next[107] ),
    .B(\u_inv.d_reg[107] ));
 sg13g2_o21ai_1 _34530_ (.B1(_03941_),
    .Y(_03942_),
    .A1(_03939_),
    .A2(_03940_));
 sg13g2_nor2_1 _34531_ (.A(_03882_),
    .B(_03887_),
    .Y(_03943_));
 sg13g2_a21oi_1 _34532_ (.A1(\u_inv.d_next[109] ),
    .A2(\u_inv.d_reg[109] ),
    .Y(_03944_),
    .B1(_03943_));
 sg13g2_inv_1 _34533_ (.Y(_03945_),
    .A(_03944_));
 sg13g2_a21oi_1 _34534_ (.A1(_18141_),
    .A2(_18503_),
    .Y(_03946_),
    .B1(_03879_));
 sg13g2_a21oi_1 _34535_ (.A1(\u_inv.d_next[111] ),
    .A2(\u_inv.d_reg[111] ),
    .Y(_03947_),
    .B1(_03946_));
 sg13g2_o21ai_1 _34536_ (.B1(_03947_),
    .Y(_03948_),
    .A1(_03881_),
    .A2(_03944_));
 sg13g2_a21oi_1 _34537_ (.A1(_03889_),
    .A2(_03942_),
    .Y(_03949_),
    .B1(_03948_));
 sg13g2_o21ai_1 _34538_ (.B1(_03949_),
    .Y(_03950_),
    .A1(_03902_),
    .A2(_03936_));
 sg13g2_xor2_1 _34539_ (.B(\u_inv.d_reg[112] ),
    .A(\u_inv.d_next[112] ),
    .X(_03951_));
 sg13g2_xnor2_1 _34540_ (.Y(_03952_),
    .A(\u_inv.d_next[112] ),
    .B(\u_inv.d_reg[112] ));
 sg13g2_nand2_1 _34541_ (.Y(_03953_),
    .A(_03859_),
    .B(_03951_));
 sg13g2_or2_1 _34542_ (.X(_03954_),
    .B(_03953_),
    .A(_03865_));
 sg13g2_or2_1 _34543_ (.X(_03955_),
    .B(_03954_),
    .A(_03854_));
 sg13g2_nand2_1 _34544_ (.Y(_03956_),
    .A(\u_inv.d_next[94] ),
    .B(\u_inv.d_reg[94] ));
 sg13g2_xnor2_1 _34545_ (.Y(_03957_),
    .A(\u_inv.d_next[94] ),
    .B(\u_inv.d_reg[94] ));
 sg13g2_inv_1 _34546_ (.Y(_03958_),
    .A(_03957_));
 sg13g2_xor2_1 _34547_ (.B(\u_inv.d_reg[95] ),
    .A(\u_inv.d_next[95] ),
    .X(_03959_));
 sg13g2_xnor2_1 _34548_ (.Y(_03960_),
    .A(\u_inv.d_next[95] ),
    .B(\u_inv.d_reg[95] ));
 sg13g2_nor2_1 _34549_ (.A(_03957_),
    .B(_03960_),
    .Y(_03961_));
 sg13g2_xor2_1 _34550_ (.B(\u_inv.d_reg[93] ),
    .A(\u_inv.d_next[93] ),
    .X(_03962_));
 sg13g2_xnor2_1 _34551_ (.Y(_03963_),
    .A(\u_inv.d_next[92] ),
    .B(\u_inv.d_reg[92] ));
 sg13g2_inv_1 _34552_ (.Y(_03964_),
    .A(_03963_));
 sg13g2_nand3_1 _34553_ (.B(_03962_),
    .C(_03964_),
    .A(_03961_),
    .Y(_03965_));
 sg13g2_nand2b_1 _34554_ (.Y(_03966_),
    .B(\u_inv.d_reg[91] ),
    .A_N(\u_inv.d_next[91] ));
 sg13g2_nand2b_1 _34555_ (.Y(_03967_),
    .B(\u_inv.d_next[91] ),
    .A_N(\u_inv.d_reg[91] ));
 sg13g2_and2_1 _34556_ (.A(_03966_),
    .B(_03967_),
    .X(_03968_));
 sg13g2_nand2_1 _34557_ (.Y(_03969_),
    .A(_03966_),
    .B(_03967_));
 sg13g2_nor2_1 _34558_ (.A(\u_inv.d_next[90] ),
    .B(\u_inv.d_reg[90] ),
    .Y(_03970_));
 sg13g2_and2_1 _34559_ (.A(\u_inv.d_next[90] ),
    .B(\u_inv.d_reg[90] ),
    .X(_03971_));
 sg13g2_nand2_1 _34560_ (.Y(_03972_),
    .A(\u_inv.d_next[90] ),
    .B(\u_inv.d_reg[90] ));
 sg13g2_nand2b_2 _34561_ (.Y(_03973_),
    .B(_03972_),
    .A_N(_03970_));
 sg13g2_nor2_1 _34562_ (.A(_03968_),
    .B(_03973_),
    .Y(_03974_));
 sg13g2_xnor2_1 _34563_ (.Y(_03975_),
    .A(\u_inv.d_next[89] ),
    .B(\u_inv.d_reg[89] ));
 sg13g2_xor2_1 _34564_ (.B(\u_inv.d_reg[89] ),
    .A(\u_inv.d_next[89] ),
    .X(_03976_));
 sg13g2_and2_1 _34565_ (.A(\u_inv.d_next[88] ),
    .B(\u_inv.d_reg[88] ),
    .X(_03977_));
 sg13g2_xor2_1 _34566_ (.B(\u_inv.d_reg[88] ),
    .A(\u_inv.d_next[88] ),
    .X(_03978_));
 sg13g2_and2_1 _34567_ (.A(_03976_),
    .B(_03978_),
    .X(_03979_));
 sg13g2_nand3b_1 _34568_ (.B(_03974_),
    .C(_03979_),
    .Y(_03980_),
    .A_N(_03965_));
 sg13g2_xnor2_1 _34569_ (.Y(_03981_),
    .A(\u_inv.d_next[83] ),
    .B(\u_inv.d_reg[83] ));
 sg13g2_xnor2_1 _34570_ (.Y(_03982_),
    .A(\u_inv.d_next[81] ),
    .B(net7290));
 sg13g2_xor2_1 _34571_ (.B(net7290),
    .A(\u_inv.d_next[81] ),
    .X(_03983_));
 sg13g2_nor2_1 _34572_ (.A(\u_inv.d_next[82] ),
    .B(\u_inv.d_reg[82] ),
    .Y(_03984_));
 sg13g2_nand2_1 _34573_ (.Y(_03985_),
    .A(\u_inv.d_next[82] ),
    .B(\u_inv.d_reg[82] ));
 sg13g2_nand2b_2 _34574_ (.Y(_03986_),
    .B(_03985_),
    .A_N(_03984_));
 sg13g2_nand2_1 _34575_ (.Y(_03987_),
    .A(\u_inv.d_next[80] ),
    .B(\u_inv.d_reg[80] ));
 sg13g2_xnor2_1 _34576_ (.Y(_03988_),
    .A(\u_inv.d_next[80] ),
    .B(\u_inv.d_reg[80] ));
 sg13g2_inv_2 _34577_ (.Y(_03989_),
    .A(_03988_));
 sg13g2_nor4_1 _34578_ (.A(_03981_),
    .B(_03982_),
    .C(_03986_),
    .D(_03988_),
    .Y(_03990_));
 sg13g2_xnor2_1 _34579_ (.Y(_03991_),
    .A(\u_inv.d_next[85] ),
    .B(\u_inv.d_reg[85] ));
 sg13g2_nand2_1 _34580_ (.Y(_03992_),
    .A(\u_inv.d_next[84] ),
    .B(\u_inv.d_reg[84] ));
 sg13g2_xnor2_1 _34581_ (.Y(_03993_),
    .A(\u_inv.d_next[84] ),
    .B(\u_inv.d_reg[84] ));
 sg13g2_nor2_1 _34582_ (.A(_03991_),
    .B(_03993_),
    .Y(_03994_));
 sg13g2_nand2_1 _34583_ (.Y(_03995_),
    .A(\u_inv.d_next[86] ),
    .B(\u_inv.d_reg[86] ));
 sg13g2_xor2_1 _34584_ (.B(\u_inv.d_reg[86] ),
    .A(\u_inv.d_next[86] ),
    .X(_03996_));
 sg13g2_xnor2_1 _34585_ (.Y(_03997_),
    .A(\u_inv.d_next[86] ),
    .B(\u_inv.d_reg[86] ));
 sg13g2_nand2_1 _34586_ (.Y(_03998_),
    .A(\u_inv.d_next[87] ),
    .B(_18527_));
 sg13g2_xnor2_1 _34587_ (.Y(_03999_),
    .A(\u_inv.d_next[87] ),
    .B(\u_inv.d_reg[87] ));
 sg13g2_xor2_1 _34588_ (.B(\u_inv.d_reg[87] ),
    .A(\u_inv.d_next[87] ),
    .X(_04000_));
 sg13g2_nor4_1 _34589_ (.A(_03991_),
    .B(_03993_),
    .C(_03997_),
    .D(_03999_),
    .Y(_04001_));
 sg13g2_nand3_1 _34590_ (.B(_03996_),
    .C(_04000_),
    .A(_03994_),
    .Y(_04002_));
 sg13g2_nand3b_1 _34591_ (.B(_03990_),
    .C(_04001_),
    .Y(_04003_),
    .A_N(_03980_));
 sg13g2_and2_1 _34592_ (.A(\u_inv.d_next[68] ),
    .B(\u_inv.d_reg[68] ),
    .X(_04004_));
 sg13g2_nand2_1 _34593_ (.Y(_04005_),
    .A(\u_inv.d_next[68] ),
    .B(\u_inv.d_reg[68] ));
 sg13g2_xor2_1 _34594_ (.B(\u_inv.d_reg[68] ),
    .A(\u_inv.d_next[68] ),
    .X(_04006_));
 sg13g2_and2_1 _34595_ (.A(\u_inv.d_next[69] ),
    .B(\u_inv.d_reg[69] ),
    .X(_04007_));
 sg13g2_or2_1 _34596_ (.X(_04008_),
    .B(\u_inv.d_reg[69] ),
    .A(\u_inv.d_next[69] ));
 sg13g2_xor2_1 _34597_ (.B(\u_inv.d_reg[69] ),
    .A(\u_inv.d_next[69] ),
    .X(_04009_));
 sg13g2_nand2b_1 _34598_ (.Y(_04010_),
    .B(_04008_),
    .A_N(_04007_));
 sg13g2_nand2_1 _34599_ (.Y(_04011_),
    .A(_04006_),
    .B(_04009_));
 sg13g2_nand2_1 _34600_ (.Y(_04012_),
    .A(net7297),
    .B(\u_inv.d_reg[70] ));
 sg13g2_xor2_1 _34601_ (.B(\u_inv.d_reg[70] ),
    .A(net7297),
    .X(_04013_));
 sg13g2_xnor2_1 _34602_ (.Y(_04014_),
    .A(net7297),
    .B(\u_inv.d_reg[70] ));
 sg13g2_nor2b_1 _34603_ (.A(\u_inv.d_next[71] ),
    .B_N(\u_inv.d_reg[71] ),
    .Y(_04015_));
 sg13g2_nand2b_1 _34604_ (.Y(_04016_),
    .B(\u_inv.d_next[71] ),
    .A_N(\u_inv.d_reg[71] ));
 sg13g2_nor2b_2 _34605_ (.A(_04015_),
    .B_N(_04016_),
    .Y(_04017_));
 sg13g2_xor2_1 _34606_ (.B(\u_inv.d_reg[71] ),
    .A(\u_inv.d_next[71] ),
    .X(_04018_));
 sg13g2_nor3_2 _34607_ (.A(_04011_),
    .B(_04014_),
    .C(_04017_),
    .Y(_04019_));
 sg13g2_nand2_1 _34608_ (.Y(_04020_),
    .A(\u_inv.d_next[67] ),
    .B(\u_inv.d_reg[67] ));
 sg13g2_nand2_1 _34609_ (.Y(_04021_),
    .A(\u_inv.d_next[66] ),
    .B(\u_inv.d_reg[66] ));
 sg13g2_nand2b_1 _34610_ (.Y(_04022_),
    .B(\u_inv.d_reg[65] ),
    .A_N(\u_inv.d_next[65] ));
 sg13g2_nor2b_1 _34611_ (.A(\u_inv.d_reg[65] ),
    .B_N(\u_inv.d_next[65] ),
    .Y(_04023_));
 sg13g2_xor2_1 _34612_ (.B(\u_inv.d_reg[65] ),
    .A(\u_inv.d_next[65] ),
    .X(_04024_));
 sg13g2_and2_1 _34613_ (.A(\u_inv.d_next[64] ),
    .B(\u_inv.d_reg[64] ),
    .X(_04025_));
 sg13g2_and2_1 _34614_ (.A(_04024_),
    .B(_04025_),
    .X(_04026_));
 sg13g2_and2_1 _34615_ (.A(\u_inv.d_next[65] ),
    .B(\u_inv.d_reg[65] ),
    .X(_04027_));
 sg13g2_a221oi_1 _34616_ (.B2(_04025_),
    .C1(_04027_),
    .B1(_04024_),
    .A1(\u_inv.d_next[66] ),
    .Y(_04028_),
    .A2(\u_inv.d_reg[66] ));
 sg13g2_xnor2_1 _34617_ (.Y(_04029_),
    .A(\u_inv.d_next[67] ),
    .B(\u_inv.d_reg[67] ));
 sg13g2_a21o_1 _34618_ (.A2(_18548_),
    .A1(_18159_),
    .B1(_04029_),
    .X(_04030_));
 sg13g2_xnor2_1 _34619_ (.Y(_04031_),
    .A(\u_inv.d_next[66] ),
    .B(\u_inv.d_reg[66] ));
 sg13g2_o21ai_1 _34620_ (.B1(_04020_),
    .Y(_04032_),
    .A1(_04028_),
    .A2(_04030_));
 sg13g2_nand2_1 _34621_ (.Y(_04033_),
    .A(\u_inv.d_next[71] ),
    .B(\u_inv.d_reg[71] ));
 sg13g2_a21oi_1 _34622_ (.A1(_04004_),
    .A2(_04008_),
    .Y(_04034_),
    .B1(_04007_));
 sg13g2_a221oi_1 _34623_ (.B2(_04008_),
    .C1(_04007_),
    .B1(_04004_),
    .A1(net7297),
    .Y(_04035_),
    .A2(\u_inv.d_reg[70] ));
 sg13g2_o21ai_1 _34624_ (.B1(_04018_),
    .Y(_04036_),
    .A1(net7297),
    .A2(\u_inv.d_reg[70] ));
 sg13g2_o21ai_1 _34625_ (.B1(_04033_),
    .Y(_04037_),
    .A1(_04035_),
    .A2(_04036_));
 sg13g2_a21o_1 _34626_ (.A2(_04032_),
    .A1(_04019_),
    .B1(_04037_),
    .X(_04038_));
 sg13g2_xnor2_1 _34627_ (.Y(_04039_),
    .A(\u_inv.d_next[77] ),
    .B(\u_inv.d_reg[77] ));
 sg13g2_nand2_1 _34628_ (.Y(_04040_),
    .A(\u_inv.d_next[76] ),
    .B(\u_inv.d_reg[76] ));
 sg13g2_xnor2_1 _34629_ (.Y(_04041_),
    .A(\u_inv.d_next[76] ),
    .B(\u_inv.d_reg[76] ));
 sg13g2_nand2_1 _34630_ (.Y(_04042_),
    .A(\u_inv.d_next[78] ),
    .B(\u_inv.d_reg[78] ));
 sg13g2_xor2_1 _34631_ (.B(\u_inv.d_reg[78] ),
    .A(\u_inv.d_next[78] ),
    .X(_04043_));
 sg13g2_xnor2_1 _34632_ (.Y(_04044_),
    .A(\u_inv.d_next[78] ),
    .B(\u_inv.d_reg[78] ));
 sg13g2_nor2b_1 _34633_ (.A(\u_inv.d_next[79] ),
    .B_N(\u_inv.d_reg[79] ),
    .Y(_04045_));
 sg13g2_nand2b_1 _34634_ (.Y(_04046_),
    .B(\u_inv.d_next[79] ),
    .A_N(\u_inv.d_reg[79] ));
 sg13g2_nor2b_2 _34635_ (.A(_04045_),
    .B_N(_04046_),
    .Y(_04047_));
 sg13g2_nor4_1 _34636_ (.A(_04039_),
    .B(_04041_),
    .C(_04044_),
    .D(_04047_),
    .Y(_04048_));
 sg13g2_xnor2_1 _34637_ (.Y(_04049_),
    .A(\u_inv.d_next[75] ),
    .B(\u_inv.d_reg[75] ));
 sg13g2_xor2_1 _34638_ (.B(\u_inv.d_reg[75] ),
    .A(\u_inv.d_next[75] ),
    .X(_04050_));
 sg13g2_and2_1 _34639_ (.A(\u_inv.d_next[74] ),
    .B(\u_inv.d_reg[74] ),
    .X(_04051_));
 sg13g2_xor2_1 _34640_ (.B(\u_inv.d_reg[74] ),
    .A(\u_inv.d_next[74] ),
    .X(_04052_));
 sg13g2_xnor2_1 _34641_ (.Y(_04053_),
    .A(\u_inv.d_next[74] ),
    .B(\u_inv.d_reg[74] ));
 sg13g2_nand2_1 _34642_ (.Y(_04054_),
    .A(\u_inv.d_next[73] ),
    .B(\u_inv.d_reg[73] ));
 sg13g2_nor2_1 _34643_ (.A(\u_inv.d_next[73] ),
    .B(\u_inv.d_reg[73] ),
    .Y(_04055_));
 sg13g2_xnor2_1 _34644_ (.Y(_04056_),
    .A(\u_inv.d_next[73] ),
    .B(\u_inv.d_reg[73] ));
 sg13g2_nand2_1 _34645_ (.Y(_04057_),
    .A(\u_inv.d_next[72] ),
    .B(\u_inv.d_reg[72] ));
 sg13g2_xor2_1 _34646_ (.B(\u_inv.d_reg[72] ),
    .A(\u_inv.d_next[72] ),
    .X(_04058_));
 sg13g2_xnor2_1 _34647_ (.Y(_04059_),
    .A(\u_inv.d_next[72] ),
    .B(\u_inv.d_reg[72] ));
 sg13g2_nor4_1 _34648_ (.A(_04049_),
    .B(_04053_),
    .C(_04056_),
    .D(_04059_),
    .Y(_04060_));
 sg13g2_and2_1 _34649_ (.A(_04048_),
    .B(_04060_),
    .X(_04061_));
 sg13g2_nand2_1 _34650_ (.Y(_04062_),
    .A(_04038_),
    .B(_04061_));
 sg13g2_nand2_1 _34651_ (.Y(_04063_),
    .A(\u_inv.d_next[75] ),
    .B(\u_inv.d_reg[75] ));
 sg13g2_o21ai_1 _34652_ (.B1(_04054_),
    .Y(_04064_),
    .A1(_04055_),
    .A2(_04057_));
 sg13g2_inv_1 _34653_ (.Y(_04065_),
    .A(_04064_));
 sg13g2_a21oi_1 _34654_ (.A1(_04052_),
    .A2(_04064_),
    .Y(_04066_),
    .B1(_04051_));
 sg13g2_o21ai_1 _34655_ (.B1(_04063_),
    .Y(_04067_),
    .A1(_04049_),
    .A2(_04066_));
 sg13g2_a22oi_1 _34656_ (.Y(_04068_),
    .B1(\u_inv.d_reg[76] ),
    .B2(\u_inv.d_next[76] ),
    .A2(\u_inv.d_reg[77] ),
    .A1(\u_inv.d_next[77] ));
 sg13g2_a21oi_1 _34657_ (.A1(_18154_),
    .A2(_18537_),
    .Y(_04069_),
    .B1(_04068_));
 sg13g2_nand2_1 _34658_ (.Y(_04070_),
    .A(_04043_),
    .B(_04069_));
 sg13g2_a21oi_1 _34659_ (.A1(_04042_),
    .A2(_04070_),
    .Y(_04071_),
    .B1(_04047_));
 sg13g2_a221oi_1 _34660_ (.B2(_04067_),
    .C1(_04071_),
    .B1(_04048_),
    .A1(\u_inv.d_next[79] ),
    .Y(_04072_),
    .A2(\u_inv.d_reg[79] ));
 sg13g2_nand2_1 _34661_ (.Y(_04073_),
    .A(_04062_),
    .B(_04072_));
 sg13g2_a21oi_1 _34662_ (.A1(_04062_),
    .A2(_04072_),
    .Y(_04074_),
    .B1(_04003_));
 sg13g2_and2_1 _34663_ (.A(\u_inv.d_next[91] ),
    .B(\u_inv.d_reg[91] ),
    .X(_04075_));
 sg13g2_nand2_1 _34664_ (.Y(_04076_),
    .A(_03976_),
    .B(_03977_));
 sg13g2_nand2_1 _34665_ (.Y(_04077_),
    .A(\u_inv.d_next[89] ),
    .B(\u_inv.d_reg[89] ));
 sg13g2_and2_1 _34666_ (.A(_04076_),
    .B(_04077_),
    .X(_04078_));
 sg13g2_a21oi_1 _34667_ (.A1(_03972_),
    .A2(_04078_),
    .Y(_04079_),
    .B1(_03970_));
 sg13g2_a21oi_2 _34668_ (.B1(_04075_),
    .Y(_04080_),
    .A2(_04079_),
    .A1(_03969_));
 sg13g2_and3_1 _34669_ (.X(_04081_),
    .A(\u_inv.d_next[92] ),
    .B(\u_inv.d_reg[92] ),
    .C(_03962_));
 sg13g2_a21o_1 _34670_ (.A2(\u_inv.d_reg[93] ),
    .A1(\u_inv.d_next[93] ),
    .B1(_04081_),
    .X(_04082_));
 sg13g2_a21oi_1 _34671_ (.A1(_18147_),
    .A2(_18519_),
    .Y(_04083_),
    .B1(_03956_));
 sg13g2_a221oi_1 _34672_ (.B2(_04082_),
    .C1(_04083_),
    .B1(_03961_),
    .A1(\u_inv.d_next[95] ),
    .Y(_04084_),
    .A2(\u_inv.d_reg[95] ));
 sg13g2_o21ai_1 _34673_ (.B1(_04084_),
    .Y(_04085_),
    .A1(_03965_),
    .A2(_04080_));
 sg13g2_nand2_1 _34674_ (.Y(_04086_),
    .A(\u_inv.d_next[83] ),
    .B(\u_inv.d_reg[83] ));
 sg13g2_nor2_1 _34675_ (.A(_03982_),
    .B(_03987_),
    .Y(_04087_));
 sg13g2_a21oi_1 _34676_ (.A1(\u_inv.d_next[81] ),
    .A2(net7290),
    .Y(_04088_),
    .B1(_04087_));
 sg13g2_a221oi_1 _34677_ (.B2(\u_inv.d_next[81] ),
    .C1(_04087_),
    .B1(net7290),
    .A1(\u_inv.d_next[82] ),
    .Y(_04089_),
    .A2(\u_inv.d_reg[82] ));
 sg13g2_or2_1 _34678_ (.X(_04090_),
    .B(_03984_),
    .A(_03981_));
 sg13g2_o21ai_1 _34679_ (.B1(_04086_),
    .Y(_04091_),
    .A1(_04089_),
    .A2(_04090_));
 sg13g2_o21ai_1 _34680_ (.B1(_03992_),
    .Y(_04092_),
    .A1(_18150_),
    .A2(_18529_));
 sg13g2_o21ai_1 _34681_ (.B1(_04092_),
    .Y(_04093_),
    .A1(\u_inv.d_next[85] ),
    .A2(\u_inv.d_reg[85] ));
 sg13g2_o21ai_1 _34682_ (.B1(_04000_),
    .Y(_04094_),
    .A1(\u_inv.d_next[86] ),
    .A2(\u_inv.d_reg[86] ));
 sg13g2_a21oi_1 _34683_ (.A1(_03995_),
    .A2(_04093_),
    .Y(_04095_),
    .B1(_04094_));
 sg13g2_a221oi_1 _34684_ (.B2(_04091_),
    .C1(_04095_),
    .B1(_04001_),
    .A1(\u_inv.d_next[87] ),
    .Y(_04096_),
    .A2(\u_inv.d_reg[87] ));
 sg13g2_nor2_1 _34685_ (.A(_03980_),
    .B(_04096_),
    .Y(_04097_));
 sg13g2_nor3_2 _34686_ (.A(_04074_),
    .B(_04085_),
    .C(_04097_),
    .Y(_04098_));
 sg13g2_nand2_1 _34687_ (.Y(_04099_),
    .A(\u_inv.d_next[63] ),
    .B(\u_inv.d_reg[63] ));
 sg13g2_nor2_1 _34688_ (.A(\u_inv.d_next[63] ),
    .B(\u_inv.d_reg[63] ),
    .Y(_04100_));
 sg13g2_xnor2_1 _34689_ (.Y(_04101_),
    .A(\u_inv.d_next[63] ),
    .B(\u_inv.d_reg[63] ));
 sg13g2_nand2_1 _34690_ (.Y(_04102_),
    .A(\u_inv.d_next[62] ),
    .B(\u_inv.d_reg[62] ));
 sg13g2_xnor2_1 _34691_ (.Y(_04103_),
    .A(\u_inv.d_next[62] ),
    .B(\u_inv.d_reg[62] ));
 sg13g2_or2_1 _34692_ (.X(_04104_),
    .B(_04103_),
    .A(_04101_));
 sg13g2_xnor2_1 _34693_ (.Y(_04105_),
    .A(\u_inv.d_next[61] ),
    .B(\u_inv.d_reg[61] ));
 sg13g2_nand2_1 _34694_ (.Y(_04106_),
    .A(\u_inv.d_next[60] ),
    .B(\u_inv.d_reg[60] ));
 sg13g2_xor2_1 _34695_ (.B(\u_inv.d_reg[60] ),
    .A(\u_inv.d_next[60] ),
    .X(_04107_));
 sg13g2_nand2b_1 _34696_ (.Y(_04108_),
    .B(_04107_),
    .A_N(_04105_));
 sg13g2_nor2_1 _34697_ (.A(_04104_),
    .B(_04108_),
    .Y(_04109_));
 sg13g2_nor2_1 _34698_ (.A(\u_inv.d_next[59] ),
    .B(_18555_),
    .Y(_04110_));
 sg13g2_xnor2_1 _34699_ (.Y(_04111_),
    .A(\u_inv.d_next[59] ),
    .B(\u_inv.d_reg[59] ));
 sg13g2_nand2_1 _34700_ (.Y(_04112_),
    .A(\u_inv.d_next[58] ),
    .B(\u_inv.d_reg[58] ));
 sg13g2_xnor2_1 _34701_ (.Y(_04113_),
    .A(\u_inv.d_next[58] ),
    .B(\u_inv.d_reg[58] ));
 sg13g2_inv_1 _34702_ (.Y(_04114_),
    .A(_04113_));
 sg13g2_nor2_1 _34703_ (.A(_04111_),
    .B(_04113_),
    .Y(_04115_));
 sg13g2_inv_1 _34704_ (.Y(_04116_),
    .A(_04115_));
 sg13g2_nor2b_1 _34705_ (.A(\u_inv.d_next[57] ),
    .B_N(\u_inv.d_reg[57] ),
    .Y(_04117_));
 sg13g2_nand2b_1 _34706_ (.Y(_04118_),
    .B(\u_inv.d_next[57] ),
    .A_N(\u_inv.d_reg[57] ));
 sg13g2_nor2b_1 _34707_ (.A(_04117_),
    .B_N(_04118_),
    .Y(_04119_));
 sg13g2_nand2b_2 _34708_ (.Y(_04120_),
    .B(_04118_),
    .A_N(_04117_));
 sg13g2_nand2_1 _34709_ (.Y(_04121_),
    .A(\u_inv.d_next[56] ),
    .B(\u_inv.d_reg[56] ));
 sg13g2_xor2_1 _34710_ (.B(\u_inv.d_reg[56] ),
    .A(\u_inv.d_next[56] ),
    .X(_04122_));
 sg13g2_xnor2_1 _34711_ (.Y(_04123_),
    .A(\u_inv.d_next[56] ),
    .B(\u_inv.d_reg[56] ));
 sg13g2_nor2_1 _34712_ (.A(_04119_),
    .B(_04123_),
    .Y(_04124_));
 sg13g2_nand3_1 _34713_ (.B(_04115_),
    .C(_04124_),
    .A(_04109_),
    .Y(_04125_));
 sg13g2_and2_1 _34714_ (.A(\u_inv.d_next[52] ),
    .B(\u_inv.d_reg[52] ),
    .X(_04126_));
 sg13g2_xor2_1 _34715_ (.B(\u_inv.d_reg[52] ),
    .A(\u_inv.d_next[52] ),
    .X(_04127_));
 sg13g2_xnor2_1 _34716_ (.Y(_04128_),
    .A(\u_inv.d_next[52] ),
    .B(\u_inv.d_reg[52] ));
 sg13g2_and2_1 _34717_ (.A(\u_inv.d_next[53] ),
    .B(\u_inv.d_reg[53] ),
    .X(_04129_));
 sg13g2_nand2_1 _34718_ (.Y(_04130_),
    .A(\u_inv.d_next[53] ),
    .B(\u_inv.d_reg[53] ));
 sg13g2_or2_1 _34719_ (.X(_04131_),
    .B(\u_inv.d_reg[53] ),
    .A(\u_inv.d_next[53] ));
 sg13g2_nand2_2 _34720_ (.Y(_04132_),
    .A(_04130_),
    .B(_04131_));
 sg13g2_nor2_1 _34721_ (.A(_18162_),
    .B(\u_inv.d_reg[55] ),
    .Y(_04133_));
 sg13g2_xnor2_1 _34722_ (.Y(_04134_),
    .A(\u_inv.d_next[55] ),
    .B(\u_inv.d_reg[55] ));
 sg13g2_or2_1 _34723_ (.X(_04135_),
    .B(\u_inv.d_reg[54] ),
    .A(\u_inv.d_next[54] ));
 sg13g2_nand2_2 _34724_ (.Y(_04136_),
    .A(\u_inv.d_next[54] ),
    .B(\u_inv.d_reg[54] ));
 sg13g2_nand2_2 _34725_ (.Y(_04137_),
    .A(_04135_),
    .B(_04136_));
 sg13g2_inv_1 _34726_ (.Y(_04138_),
    .A(_04137_));
 sg13g2_nor4_1 _34727_ (.A(_04128_),
    .B(_04132_),
    .C(_04134_),
    .D(_04137_),
    .Y(_04139_));
 sg13g2_nor2_1 _34728_ (.A(\u_inv.d_next[51] ),
    .B(_18563_),
    .Y(_04140_));
 sg13g2_xnor2_1 _34729_ (.Y(_04141_),
    .A(\u_inv.d_next[51] ),
    .B(\u_inv.d_reg[51] ));
 sg13g2_xor2_1 _34730_ (.B(\u_inv.d_reg[51] ),
    .A(\u_inv.d_next[51] ),
    .X(_04142_));
 sg13g2_and2_1 _34731_ (.A(net7298),
    .B(\u_inv.d_reg[50] ),
    .X(_04143_));
 sg13g2_xor2_1 _34732_ (.B(\u_inv.d_reg[50] ),
    .A(net7298),
    .X(_04144_));
 sg13g2_xnor2_1 _34733_ (.Y(_04145_),
    .A(net7298),
    .B(\u_inv.d_reg[50] ));
 sg13g2_xor2_1 _34734_ (.B(\u_inv.d_reg[49] ),
    .A(\u_inv.d_next[49] ),
    .X(_04146_));
 sg13g2_and2_1 _34735_ (.A(\u_inv.d_next[48] ),
    .B(\u_inv.d_reg[48] ),
    .X(_04147_));
 sg13g2_nand2_1 _34736_ (.Y(_04148_),
    .A(\u_inv.d_next[48] ),
    .B(\u_inv.d_reg[48] ));
 sg13g2_xor2_1 _34737_ (.B(\u_inv.d_reg[48] ),
    .A(\u_inv.d_next[48] ),
    .X(_04149_));
 sg13g2_and2_1 _34738_ (.A(_04146_),
    .B(_04149_),
    .X(_04150_));
 sg13g2_and3_1 _34739_ (.X(_04151_),
    .A(_04142_),
    .B(_04144_),
    .C(_04150_));
 sg13g2_nand2_1 _34740_ (.Y(_04152_),
    .A(_04139_),
    .B(_04151_));
 sg13g2_inv_1 _34741_ (.Y(_04153_),
    .A(_04152_));
 sg13g2_nor2_2 _34742_ (.A(_04125_),
    .B(_04152_),
    .Y(_04154_));
 sg13g2_nand2_1 _34743_ (.Y(_04155_),
    .A(\u_inv.d_next[57] ),
    .B(\u_inv.d_reg[57] ));
 sg13g2_o21ai_1 _34744_ (.B1(_04155_),
    .Y(_04156_),
    .A1(_04119_),
    .A2(_04121_));
 sg13g2_nor2_1 _34745_ (.A(_04111_),
    .B(_04112_),
    .Y(_04157_));
 sg13g2_a221oi_1 _34746_ (.B2(_04156_),
    .C1(_04157_),
    .B1(_04115_),
    .A1(\u_inv.d_next[59] ),
    .Y(_04158_),
    .A2(\u_inv.d_reg[59] ));
 sg13g2_nor2b_1 _34747_ (.A(_04158_),
    .B_N(_04109_),
    .Y(_04159_));
 sg13g2_or2_1 _34748_ (.X(_04160_),
    .B(_04106_),
    .A(_04105_));
 sg13g2_nand2_1 _34749_ (.Y(_04161_),
    .A(\u_inv.d_next[61] ),
    .B(\u_inv.d_reg[61] ));
 sg13g2_and2_1 _34750_ (.A(_04160_),
    .B(_04161_),
    .X(_04162_));
 sg13g2_nor2_1 _34751_ (.A(_04104_),
    .B(_04162_),
    .Y(_04163_));
 sg13g2_o21ai_1 _34752_ (.B1(_04099_),
    .Y(_04164_),
    .A1(_04100_),
    .A2(_04102_));
 sg13g2_nand2_1 _34753_ (.Y(_04165_),
    .A(\u_inv.d_next[51] ),
    .B(\u_inv.d_reg[51] ));
 sg13g2_and2_1 _34754_ (.A(_04146_),
    .B(_04147_),
    .X(_04166_));
 sg13g2_and2_1 _34755_ (.A(\u_inv.d_next[49] ),
    .B(\u_inv.d_reg[49] ),
    .X(_04167_));
 sg13g2_nor2_1 _34756_ (.A(_04166_),
    .B(_04167_),
    .Y(_04168_));
 sg13g2_a221oi_1 _34757_ (.B2(_04147_),
    .C1(_04167_),
    .B1(_04146_),
    .A1(net7298),
    .Y(_04169_),
    .A2(\u_inv.d_reg[50] ));
 sg13g2_o21ai_1 _34758_ (.B1(_04142_),
    .Y(_04170_),
    .A1(net7298),
    .A2(\u_inv.d_reg[50] ));
 sg13g2_o21ai_1 _34759_ (.B1(_04165_),
    .Y(_04171_),
    .A1(_04169_),
    .A2(_04170_));
 sg13g2_a21o_1 _34760_ (.A2(_04131_),
    .A1(_04126_),
    .B1(_04129_),
    .X(_04172_));
 sg13g2_a21oi_1 _34761_ (.A1(_04126_),
    .A2(_04131_),
    .Y(_04173_),
    .B1(_04129_));
 sg13g2_a21oi_1 _34762_ (.A1(_04136_),
    .A2(_04173_),
    .Y(_04174_),
    .B1(_04134_));
 sg13g2_nor2_1 _34763_ (.A(_18162_),
    .B(_18559_),
    .Y(_04175_));
 sg13g2_a221oi_1 _34764_ (.B2(_04135_),
    .C1(_04175_),
    .B1(_04174_),
    .A1(_04139_),
    .Y(_04176_),
    .A2(_04171_));
 sg13g2_inv_1 _34765_ (.Y(_04177_),
    .A(_04176_));
 sg13g2_nor2_1 _34766_ (.A(_04125_),
    .B(_04176_),
    .Y(_04178_));
 sg13g2_xor2_1 _34767_ (.B(\u_inv.d_reg[44] ),
    .A(\u_inv.d_next[44] ),
    .X(_04179_));
 sg13g2_nand2_1 _34768_ (.Y(_04180_),
    .A(\u_inv.d_next[45] ),
    .B(\u_inv.d_reg[45] ));
 sg13g2_nor2_1 _34769_ (.A(\u_inv.d_next[45] ),
    .B(\u_inv.d_reg[45] ),
    .Y(_04181_));
 sg13g2_nand2_1 _34770_ (.Y(_04182_),
    .A(_18166_),
    .B(_18569_));
 sg13g2_xor2_1 _34771_ (.B(\u_inv.d_reg[45] ),
    .A(\u_inv.d_next[45] ),
    .X(_04183_));
 sg13g2_nand2_1 _34772_ (.Y(_04184_),
    .A(_04179_),
    .B(_04183_));
 sg13g2_xnor2_1 _34773_ (.Y(_04185_),
    .A(\u_inv.d_next[47] ),
    .B(\u_inv.d_reg[47] ));
 sg13g2_or2_1 _34774_ (.X(_04186_),
    .B(\u_inv.d_reg[46] ),
    .A(\u_inv.d_next[46] ));
 sg13g2_and2_1 _34775_ (.A(\u_inv.d_next[46] ),
    .B(\u_inv.d_reg[46] ),
    .X(_04187_));
 sg13g2_nand2_1 _34776_ (.Y(_04188_),
    .A(\u_inv.d_next[46] ),
    .B(\u_inv.d_reg[46] ));
 sg13g2_nand2_2 _34777_ (.Y(_04189_),
    .A(_04186_),
    .B(_04188_));
 sg13g2_or3_1 _34778_ (.A(_04184_),
    .B(_04185_),
    .C(_04189_),
    .X(_04190_));
 sg13g2_xnor2_1 _34779_ (.Y(_04191_),
    .A(\u_inv.d_next[43] ),
    .B(\u_inv.d_reg[43] ));
 sg13g2_nand2_1 _34780_ (.Y(_04192_),
    .A(\u_inv.d_next[42] ),
    .B(\u_inv.d_reg[42] ));
 sg13g2_xor2_1 _34781_ (.B(\u_inv.d_reg[42] ),
    .A(\u_inv.d_next[42] ),
    .X(_04193_));
 sg13g2_inv_1 _34782_ (.Y(_04194_),
    .A(_04193_));
 sg13g2_nand2b_1 _34783_ (.Y(_04195_),
    .B(_04193_),
    .A_N(_04191_));
 sg13g2_nor2_1 _34784_ (.A(\u_inv.d_next[41] ),
    .B(\u_inv.d_reg[41] ),
    .Y(_04196_));
 sg13g2_xor2_1 _34785_ (.B(\u_inv.d_reg[41] ),
    .A(\u_inv.d_next[41] ),
    .X(_04197_));
 sg13g2_and2_1 _34786_ (.A(\u_inv.d_next[40] ),
    .B(\u_inv.d_reg[40] ),
    .X(_04198_));
 sg13g2_xor2_1 _34787_ (.B(\u_inv.d_reg[40] ),
    .A(\u_inv.d_next[40] ),
    .X(_04199_));
 sg13g2_nand2_1 _34788_ (.Y(_04200_),
    .A(_04197_),
    .B(_04199_));
 sg13g2_nor3_1 _34789_ (.A(_04190_),
    .B(_04195_),
    .C(_04200_),
    .Y(_04201_));
 sg13g2_inv_1 _34790_ (.Y(_04202_),
    .A(_04201_));
 sg13g2_xnor2_1 _34791_ (.Y(_04203_),
    .A(\u_inv.d_next[29] ),
    .B(\u_inv.d_reg[29] ));
 sg13g2_xnor2_1 _34792_ (.Y(_04204_),
    .A(\u_inv.d_next[28] ),
    .B(\u_inv.d_reg[28] ));
 sg13g2_nor2_1 _34793_ (.A(_04203_),
    .B(_04204_),
    .Y(_04205_));
 sg13g2_xnor2_1 _34794_ (.Y(_04206_),
    .A(\u_inv.d_next[31] ),
    .B(\u_inv.d_reg[31] ));
 sg13g2_nor2_1 _34795_ (.A(\u_inv.d_next[30] ),
    .B(\u_inv.d_reg[30] ),
    .Y(_04207_));
 sg13g2_xnor2_1 _34796_ (.Y(_04208_),
    .A(\u_inv.d_next[30] ),
    .B(\u_inv.d_reg[30] ));
 sg13g2_nor4_1 _34797_ (.A(_04203_),
    .B(_04204_),
    .C(_04206_),
    .D(_04208_),
    .Y(_04209_));
 sg13g2_nand2b_1 _34798_ (.Y(_04210_),
    .B(\u_inv.d_reg[27] ),
    .A_N(\u_inv.d_next[27] ));
 sg13g2_nand2b_1 _34799_ (.Y(_04211_),
    .B(\u_inv.d_next[27] ),
    .A_N(\u_inv.d_reg[27] ));
 sg13g2_and2_1 _34800_ (.A(_04210_),
    .B(_04211_),
    .X(_04212_));
 sg13g2_nand2_1 _34801_ (.Y(_04213_),
    .A(\u_inv.d_next[26] ),
    .B(\u_inv.d_reg[26] ));
 sg13g2_xnor2_1 _34802_ (.Y(_04214_),
    .A(\u_inv.d_next[26] ),
    .B(\u_inv.d_reg[26] ));
 sg13g2_nor2_1 _34803_ (.A(_04212_),
    .B(_04214_),
    .Y(_04215_));
 sg13g2_nor2_1 _34804_ (.A(\u_inv.d_next[25] ),
    .B(\u_inv.d_reg[25] ),
    .Y(_04216_));
 sg13g2_xnor2_1 _34805_ (.Y(_04217_),
    .A(\u_inv.d_next[25] ),
    .B(\u_inv.d_reg[25] ));
 sg13g2_xnor2_1 _34806_ (.Y(_04218_),
    .A(\u_inv.d_next[24] ),
    .B(\u_inv.d_reg[24] ));
 sg13g2_nor2_1 _34807_ (.A(_04217_),
    .B(_04218_),
    .Y(_04219_));
 sg13g2_nand2_1 _34808_ (.Y(_04220_),
    .A(_04215_),
    .B(_04219_));
 sg13g2_nand3_1 _34809_ (.B(_04215_),
    .C(_04219_),
    .A(_04209_),
    .Y(_04221_));
 sg13g2_a22oi_1 _34810_ (.Y(_04222_),
    .B1(\u_inv.d_reg[28] ),
    .B2(\u_inv.d_next[28] ),
    .A2(\u_inv.d_reg[29] ),
    .A1(\u_inv.d_next[29] ));
 sg13g2_a21oi_1 _34811_ (.A1(_18175_),
    .A2(_18585_),
    .Y(_04223_),
    .B1(_04222_));
 sg13g2_a21oi_1 _34812_ (.A1(\u_inv.d_next[30] ),
    .A2(\u_inv.d_reg[30] ),
    .Y(_04224_),
    .B1(_04223_));
 sg13g2_nor3_1 _34813_ (.A(_04206_),
    .B(_04207_),
    .C(_04224_),
    .Y(_04225_));
 sg13g2_a21oi_1 _34814_ (.A1(\u_inv.d_next[31] ),
    .A2(\u_inv.d_reg[31] ),
    .Y(_04226_),
    .B1(_04225_));
 sg13g2_nand2_1 _34815_ (.Y(_04227_),
    .A(\u_inv.d_next[27] ),
    .B(\u_inv.d_reg[27] ));
 sg13g2_a22oi_1 _34816_ (.Y(_04228_),
    .B1(\u_inv.d_reg[24] ),
    .B2(\u_inv.d_next[24] ),
    .A2(\u_inv.d_reg[25] ),
    .A1(\u_inv.d_next[25] ));
 sg13g2_or2_1 _34817_ (.X(_04229_),
    .B(_04228_),
    .A(_04216_));
 sg13g2_nor3_1 _34818_ (.A(_04214_),
    .B(_04216_),
    .C(_04228_),
    .Y(_04230_));
 sg13g2_a21oi_1 _34819_ (.A1(\u_inv.d_next[26] ),
    .A2(\u_inv.d_reg[26] ),
    .Y(_04231_),
    .B1(_04230_));
 sg13g2_o21ai_1 _34820_ (.B1(_04227_),
    .Y(_04232_),
    .A1(_04212_),
    .A2(_04231_));
 sg13g2_inv_1 _34821_ (.Y(_04233_),
    .A(_04232_));
 sg13g2_nand2_1 _34822_ (.Y(_04234_),
    .A(_04209_),
    .B(_04232_));
 sg13g2_nor2_1 _34823_ (.A(\u_inv.d_next[13] ),
    .B(\u_inv.d_reg[13] ),
    .Y(_04235_));
 sg13g2_nand2_1 _34824_ (.Y(_04236_),
    .A(\u_inv.d_next[13] ),
    .B(\u_inv.d_reg[13] ));
 sg13g2_xor2_1 _34825_ (.B(\u_inv.d_reg[13] ),
    .A(\u_inv.d_next[13] ),
    .X(_04237_));
 sg13g2_nand2_1 _34826_ (.Y(_04238_),
    .A(\u_inv.d_next[12] ),
    .B(\u_inv.d_reg[12] ));
 sg13g2_xor2_1 _34827_ (.B(\u_inv.d_reg[12] ),
    .A(\u_inv.d_next[12] ),
    .X(_04239_));
 sg13g2_xnor2_1 _34828_ (.Y(_04240_),
    .A(\u_inv.d_next[12] ),
    .B(\u_inv.d_reg[12] ));
 sg13g2_nand2_1 _34829_ (.Y(_04241_),
    .A(_04237_),
    .B(_04239_));
 sg13g2_nor2_1 _34830_ (.A(\u_inv.d_next[14] ),
    .B(\u_inv.d_reg[14] ),
    .Y(_04242_));
 sg13g2_nand2_2 _34831_ (.Y(_04243_),
    .A(\u_inv.d_next[14] ),
    .B(\u_inv.d_reg[14] ));
 sg13g2_nor2b_2 _34832_ (.A(_04242_),
    .B_N(_04243_),
    .Y(_04244_));
 sg13g2_nand2b_2 _34833_ (.Y(_04245_),
    .B(_04243_),
    .A_N(_04242_));
 sg13g2_nand2b_1 _34834_ (.Y(_04246_),
    .B(\u_inv.d_reg[15] ),
    .A_N(\u_inv.d_next[15] ));
 sg13g2_nand2b_1 _34835_ (.Y(_04247_),
    .B(\u_inv.d_next[15] ),
    .A_N(\u_inv.d_reg[15] ));
 sg13g2_and2_1 _34836_ (.A(_04246_),
    .B(_04247_),
    .X(_04248_));
 sg13g2_nor3_1 _34837_ (.A(_04241_),
    .B(_04245_),
    .C(_04248_),
    .Y(_04249_));
 sg13g2_nand2_1 _34838_ (.Y(_04250_),
    .A(\u_inv.d_next[11] ),
    .B(\u_inv.d_reg[11] ));
 sg13g2_nor2b_1 _34839_ (.A(\u_inv.d_reg[11] ),
    .B_N(\u_inv.d_next[11] ),
    .Y(_04251_));
 sg13g2_nand2b_1 _34840_ (.Y(_04252_),
    .B(\u_inv.d_reg[11] ),
    .A_N(\u_inv.d_next[11] ));
 sg13g2_nor2b_2 _34841_ (.A(_04251_),
    .B_N(_04252_),
    .Y(_04253_));
 sg13g2_and2_1 _34842_ (.A(\u_inv.d_next[10] ),
    .B(net7292),
    .X(_04254_));
 sg13g2_xnor2_1 _34843_ (.Y(_04255_),
    .A(\u_inv.d_next[9] ),
    .B(\u_inv.d_reg[9] ));
 sg13g2_nand2_1 _34844_ (.Y(_04256_),
    .A(\u_inv.d_next[8] ),
    .B(\u_inv.d_reg[8] ));
 sg13g2_nand2_1 _34845_ (.Y(_04257_),
    .A(\u_inv.d_next[9] ),
    .B(\u_inv.d_reg[9] ));
 sg13g2_o21ai_1 _34846_ (.B1(_04257_),
    .Y(_04258_),
    .A1(_04255_),
    .A2(_04256_));
 sg13g2_xor2_1 _34847_ (.B(net7292),
    .A(\u_inv.d_next[10] ),
    .X(_04259_));
 sg13g2_xnor2_1 _34848_ (.Y(_04260_),
    .A(\u_inv.d_next[10] ),
    .B(net7292));
 sg13g2_a21oi_1 _34849_ (.A1(_04258_),
    .A2(_04259_),
    .Y(_04261_),
    .B1(_04254_));
 sg13g2_o21ai_1 _34850_ (.B1(_04250_),
    .Y(_04262_),
    .A1(_04253_),
    .A2(_04261_));
 sg13g2_o21ai_1 _34851_ (.B1(_04236_),
    .Y(_04263_),
    .A1(_04235_),
    .A2(_04238_));
 sg13g2_nand2_1 _34852_ (.Y(_04264_),
    .A(_04244_),
    .B(_04263_));
 sg13g2_a21oi_1 _34853_ (.A1(_04243_),
    .A2(_04264_),
    .Y(_04265_),
    .B1(_04248_));
 sg13g2_a221oi_1 _34854_ (.B2(_04262_),
    .C1(_04265_),
    .B1(_04249_),
    .A1(\u_inv.d_next[15] ),
    .Y(_04266_),
    .A2(\u_inv.d_reg[15] ));
 sg13g2_nand2b_1 _34855_ (.Y(_04267_),
    .B(\u_inv.d_reg[5] ),
    .A_N(\u_inv.d_next[5] ));
 sg13g2_nor2b_1 _34856_ (.A(\u_inv.d_reg[5] ),
    .B_N(\u_inv.d_next[5] ),
    .Y(_04268_));
 sg13g2_xnor2_1 _34857_ (.Y(_04269_),
    .A(\u_inv.d_next[5] ),
    .B(\u_inv.d_reg[5] ));
 sg13g2_nor2_1 _34858_ (.A(\u_inv.d_next[3] ),
    .B(\u_inv.d_reg[3] ),
    .Y(_04270_));
 sg13g2_a21oi_1 _34859_ (.A1(_03338_),
    .A2(_03348_),
    .Y(_04271_),
    .B1(_03337_));
 sg13g2_a221oi_1 _34860_ (.B2(_03348_),
    .C1(_03337_),
    .B1(_03338_),
    .A1(\u_inv.d_next[3] ),
    .Y(_04272_),
    .A2(\u_inv.d_reg[3] ));
 sg13g2_nand2_1 _34861_ (.Y(_04273_),
    .A(\u_inv.d_next[4] ),
    .B(\u_inv.d_reg[4] ));
 sg13g2_xor2_1 _34862_ (.B(\u_inv.d_reg[4] ),
    .A(\u_inv.d_next[4] ),
    .X(_04274_));
 sg13g2_xnor2_1 _34863_ (.Y(_04275_),
    .A(\u_inv.d_next[4] ),
    .B(\u_inv.d_reg[4] ));
 sg13g2_or3_1 _34864_ (.A(_04270_),
    .B(_04272_),
    .C(_04275_),
    .X(_04276_));
 sg13g2_nor2_1 _34865_ (.A(_04269_),
    .B(_04276_),
    .Y(_04277_));
 sg13g2_nand2b_2 _34866_ (.Y(_04278_),
    .B(\u_inv.d_reg[7] ),
    .A_N(\u_inv.d_next[7] ));
 sg13g2_xnor2_1 _34867_ (.Y(_04279_),
    .A(\u_inv.d_next[7] ),
    .B(\u_inv.d_reg[7] ));
 sg13g2_and2_1 _34868_ (.A(\u_inv.d_next[6] ),
    .B(\u_inv.d_reg[6] ),
    .X(_04280_));
 sg13g2_xor2_1 _34869_ (.B(\u_inv.d_reg[6] ),
    .A(\u_inv.d_next[6] ),
    .X(_04281_));
 sg13g2_nand3b_1 _34870_ (.B(_04274_),
    .C(_04281_),
    .Y(_04282_),
    .A_N(_04269_));
 sg13g2_nor4_1 _34871_ (.A(_04270_),
    .B(_04272_),
    .C(_04279_),
    .D(_04282_),
    .Y(_04283_));
 sg13g2_nand2_1 _34872_ (.Y(_04284_),
    .A(\u_inv.d_next[7] ),
    .B(\u_inv.d_reg[7] ));
 sg13g2_nand2_1 _34873_ (.Y(_04285_),
    .A(\u_inv.d_next[5] ),
    .B(\u_inv.d_reg[5] ));
 sg13g2_o21ai_1 _34874_ (.B1(_04285_),
    .Y(_04286_),
    .A1(_04269_),
    .A2(_04273_));
 sg13g2_a21oi_1 _34875_ (.A1(_04281_),
    .A2(_04286_),
    .Y(_04287_),
    .B1(_04280_));
 sg13g2_o21ai_1 _34876_ (.B1(_04284_),
    .Y(_04288_),
    .A1(_04279_),
    .A2(_04287_));
 sg13g2_nor2_1 _34877_ (.A(_04283_),
    .B(_04288_),
    .Y(_04289_));
 sg13g2_xnor2_1 _34878_ (.Y(_04290_),
    .A(\u_inv.d_next[8] ),
    .B(\u_inv.d_reg[8] ));
 sg13g2_or2_1 _34879_ (.X(_04291_),
    .B(_04290_),
    .A(_04289_));
 sg13g2_nor2_2 _34880_ (.A(_04255_),
    .B(_04291_),
    .Y(_04292_));
 sg13g2_nor2_1 _34881_ (.A(_04253_),
    .B(_04260_),
    .Y(_04293_));
 sg13g2_nor4_1 _34882_ (.A(_04253_),
    .B(_04255_),
    .C(_04260_),
    .D(_04290_),
    .Y(_04294_));
 sg13g2_and2_1 _34883_ (.A(_04249_),
    .B(_04294_),
    .X(_04295_));
 sg13g2_o21ai_1 _34884_ (.B1(_04295_),
    .Y(_04296_),
    .A1(_04283_),
    .A2(_04288_));
 sg13g2_nand2_1 _34885_ (.Y(_04297_),
    .A(_04266_),
    .B(_04296_));
 sg13g2_nand2_1 _34886_ (.Y(_04298_),
    .A(\u_inv.d_next[20] ),
    .B(\u_inv.d_reg[20] ));
 sg13g2_xnor2_1 _34887_ (.Y(_04299_),
    .A(\u_inv.d_next[20] ),
    .B(\u_inv.d_reg[20] ));
 sg13g2_nor2_1 _34888_ (.A(\u_inv.d_next[21] ),
    .B(\u_inv.d_reg[21] ),
    .Y(_04300_));
 sg13g2_xor2_1 _34889_ (.B(\u_inv.d_reg[21] ),
    .A(\u_inv.d_next[21] ),
    .X(_04301_));
 sg13g2_nand2b_1 _34890_ (.Y(_04302_),
    .B(_04301_),
    .A_N(_04299_));
 sg13g2_nor2b_1 _34891_ (.A(\u_inv.d_next[23] ),
    .B_N(\u_inv.d_reg[23] ),
    .Y(_04303_));
 sg13g2_nand2b_1 _34892_ (.Y(_04304_),
    .B(\u_inv.d_next[23] ),
    .A_N(\u_inv.d_reg[23] ));
 sg13g2_nor2b_2 _34893_ (.A(_04303_),
    .B_N(_04304_),
    .Y(_04305_));
 sg13g2_xor2_1 _34894_ (.B(\u_inv.d_reg[23] ),
    .A(\u_inv.d_next[23] ),
    .X(_04306_));
 sg13g2_nand2_1 _34895_ (.Y(_04307_),
    .A(\u_inv.d_next[22] ),
    .B(net7291));
 sg13g2_xor2_1 _34896_ (.B(net7291),
    .A(\u_inv.d_next[22] ),
    .X(_04308_));
 sg13g2_xnor2_1 _34897_ (.Y(_04309_),
    .A(\u_inv.d_next[22] ),
    .B(net7291));
 sg13g2_nor3_1 _34898_ (.A(_04302_),
    .B(_04305_),
    .C(_04309_),
    .Y(_04310_));
 sg13g2_xnor2_1 _34899_ (.Y(_04311_),
    .A(\u_inv.d_next[19] ),
    .B(\u_inv.d_reg[19] ));
 sg13g2_nand2b_1 _34900_ (.Y(_04312_),
    .B(\u_inv.d_reg[17] ),
    .A_N(\u_inv.d_next[17] ));
 sg13g2_nor2b_1 _34901_ (.A(\u_inv.d_reg[17] ),
    .B_N(\u_inv.d_next[17] ),
    .Y(_04313_));
 sg13g2_xnor2_1 _34902_ (.Y(_04314_),
    .A(\u_inv.d_next[17] ),
    .B(\u_inv.d_reg[17] ));
 sg13g2_xor2_1 _34903_ (.B(\u_inv.d_reg[17] ),
    .A(\u_inv.d_next[17] ),
    .X(_04315_));
 sg13g2_nand2_1 _34904_ (.Y(_04316_),
    .A(net7299),
    .B(\u_inv.d_reg[18] ));
 sg13g2_nor2_1 _34905_ (.A(net7299),
    .B(\u_inv.d_reg[18] ),
    .Y(_04317_));
 sg13g2_xnor2_1 _34906_ (.Y(_04318_),
    .A(net7299),
    .B(\u_inv.d_reg[18] ));
 sg13g2_inv_1 _34907_ (.Y(_04319_),
    .A(_04318_));
 sg13g2_and2_1 _34908_ (.A(\u_inv.d_next[16] ),
    .B(\u_inv.d_reg[16] ),
    .X(_04320_));
 sg13g2_xor2_1 _34909_ (.B(\u_inv.d_reg[16] ),
    .A(\u_inv.d_next[16] ),
    .X(_04321_));
 sg13g2_or2_1 _34910_ (.X(_04322_),
    .B(_04317_),
    .A(_04311_));
 sg13g2_nor2_1 _34911_ (.A(_04311_),
    .B(_04318_),
    .Y(_04323_));
 sg13g2_nand4_1 _34912_ (.B(_04315_),
    .C(_04321_),
    .A(_04310_),
    .Y(_04324_),
    .D(_04323_));
 sg13g2_a21oi_1 _34913_ (.A1(_04266_),
    .A2(_04296_),
    .Y(_04325_),
    .B1(_04324_));
 sg13g2_nand2_1 _34914_ (.Y(_04326_),
    .A(\u_inv.d_next[19] ),
    .B(\u_inv.d_reg[19] ));
 sg13g2_and2_1 _34915_ (.A(\u_inv.d_next[17] ),
    .B(\u_inv.d_reg[17] ),
    .X(_04327_));
 sg13g2_a21o_1 _34916_ (.A2(_04320_),
    .A1(_04315_),
    .B1(_04327_),
    .X(_04328_));
 sg13g2_a221oi_1 _34917_ (.B2(_04320_),
    .C1(_04327_),
    .B1(_04315_),
    .A1(net7299),
    .Y(_04329_),
    .A2(\u_inv.d_reg[18] ));
 sg13g2_o21ai_1 _34918_ (.B1(_04326_),
    .Y(_04330_),
    .A1(_04322_),
    .A2(_04329_));
 sg13g2_a22oi_1 _34919_ (.Y(_04331_),
    .B1(\u_inv.d_reg[20] ),
    .B2(\u_inv.d_next[20] ),
    .A2(\u_inv.d_reg[21] ),
    .A1(\u_inv.d_next[21] ));
 sg13g2_or2_1 _34920_ (.X(_04332_),
    .B(_04331_),
    .A(_04300_));
 sg13g2_o21ai_1 _34921_ (.B1(_04306_),
    .Y(_04333_),
    .A1(\u_inv.d_next[22] ),
    .A2(net7291));
 sg13g2_a21oi_1 _34922_ (.A1(_04307_),
    .A2(_04332_),
    .Y(_04334_),
    .B1(_04333_));
 sg13g2_a221oi_1 _34923_ (.B2(_04330_),
    .C1(_04334_),
    .B1(_04310_),
    .A1(\u_inv.d_next[23] ),
    .Y(_04335_),
    .A2(\u_inv.d_reg[23] ));
 sg13g2_or2_1 _34924_ (.X(_04336_),
    .B(_04335_),
    .A(_04221_));
 sg13g2_nand3_1 _34925_ (.B(_04234_),
    .C(_04336_),
    .A(_04226_),
    .Y(_04337_));
 sg13g2_or2_1 _34926_ (.X(_04338_),
    .B(_04324_),
    .A(_04221_));
 sg13g2_a21oi_2 _34927_ (.B1(_04338_),
    .Y(_04339_),
    .A2(_04296_),
    .A1(_04266_));
 sg13g2_nor2_1 _34928_ (.A(_04337_),
    .B(_04339_),
    .Y(_04340_));
 sg13g2_nor2_1 _34929_ (.A(\u_inv.d_next[37] ),
    .B(\u_inv.d_reg[37] ),
    .Y(_04341_));
 sg13g2_xnor2_1 _34930_ (.Y(_04342_),
    .A(\u_inv.d_next[37] ),
    .B(\u_inv.d_reg[37] ));
 sg13g2_nand2_1 _34931_ (.Y(_04343_),
    .A(\u_inv.d_next[36] ),
    .B(\u_inv.d_reg[36] ));
 sg13g2_xor2_1 _34932_ (.B(\u_inv.d_reg[36] ),
    .A(\u_inv.d_next[36] ),
    .X(_04344_));
 sg13g2_inv_1 _34933_ (.Y(_04345_),
    .A(_04344_));
 sg13g2_nor2b_1 _34934_ (.A(_04342_),
    .B_N(_04344_),
    .Y(_04346_));
 sg13g2_nor2b_1 _34935_ (.A(\u_inv.d_next[39] ),
    .B_N(\u_inv.d_reg[39] ),
    .Y(_04347_));
 sg13g2_nand2b_1 _34936_ (.Y(_04348_),
    .B(\u_inv.d_next[39] ),
    .A_N(\u_inv.d_reg[39] ));
 sg13g2_xnor2_1 _34937_ (.Y(_04349_),
    .A(\u_inv.d_next[39] ),
    .B(\u_inv.d_reg[39] ));
 sg13g2_nand2b_2 _34938_ (.Y(_04350_),
    .B(_04348_),
    .A_N(_04347_));
 sg13g2_nand2_1 _34939_ (.Y(_04351_),
    .A(\u_inv.d_next[38] ),
    .B(\u_inv.d_reg[38] ));
 sg13g2_xor2_1 _34940_ (.B(\u_inv.d_reg[38] ),
    .A(\u_inv.d_next[38] ),
    .X(_04352_));
 sg13g2_xnor2_1 _34941_ (.Y(_04353_),
    .A(\u_inv.d_next[38] ),
    .B(\u_inv.d_reg[38] ));
 sg13g2_nand3_1 _34942_ (.B(_04350_),
    .C(_04352_),
    .A(_04346_),
    .Y(_04354_));
 sg13g2_nand2b_1 _34943_ (.Y(_04355_),
    .B(\u_inv.d_reg[35] ),
    .A_N(\u_inv.d_next[35] ));
 sg13g2_nor2b_1 _34944_ (.A(\u_inv.d_reg[35] ),
    .B_N(\u_inv.d_next[35] ),
    .Y(_04356_));
 sg13g2_xnor2_1 _34945_ (.Y(_04357_),
    .A(\u_inv.d_next[35] ),
    .B(\u_inv.d_reg[35] ));
 sg13g2_xnor2_1 _34946_ (.Y(_04358_),
    .A(\u_inv.d_next[34] ),
    .B(\u_inv.d_reg[34] ));
 sg13g2_nor2_1 _34947_ (.A(_04357_),
    .B(_04358_),
    .Y(_04359_));
 sg13g2_or2_1 _34948_ (.X(_04360_),
    .B(_04358_),
    .A(_04357_));
 sg13g2_xnor2_1 _34949_ (.Y(_04361_),
    .A(\u_inv.d_next[33] ),
    .B(\u_inv.d_reg[33] ));
 sg13g2_inv_1 _34950_ (.Y(_04362_),
    .A(net6995));
 sg13g2_nand2_2 _34951_ (.Y(_04363_),
    .A(\u_inv.d_next[32] ),
    .B(\u_inv.d_reg[32] ));
 sg13g2_or2_1 _34952_ (.X(_04364_),
    .B(\u_inv.d_reg[32] ),
    .A(\u_inv.d_next[32] ));
 sg13g2_nand2_2 _34953_ (.Y(_04365_),
    .A(_04363_),
    .B(_04364_));
 sg13g2_nor4_1 _34954_ (.A(_04354_),
    .B(_04360_),
    .C(_04361_),
    .D(_04365_),
    .Y(_04366_));
 sg13g2_o21ai_1 _34955_ (.B1(_04366_),
    .Y(_04367_),
    .A1(_04337_),
    .A2(_04339_));
 sg13g2_nor2_1 _34956_ (.A(net6995),
    .B(_04363_),
    .Y(_04368_));
 sg13g2_nand2_1 _34957_ (.Y(_04369_),
    .A(\u_inv.d_next[33] ),
    .B(\u_inv.d_reg[33] ));
 sg13g2_nor2b_1 _34958_ (.A(_04368_),
    .B_N(_04369_),
    .Y(_04370_));
 sg13g2_o21ai_1 _34959_ (.B1(_04369_),
    .Y(_04371_),
    .A1(net6995),
    .A2(_04363_));
 sg13g2_nor3_1 _34960_ (.A(_18172_),
    .B(_18580_),
    .C(_04357_),
    .Y(_04372_));
 sg13g2_a221oi_1 _34961_ (.B2(_04371_),
    .C1(_04372_),
    .B1(_04359_),
    .A1(\u_inv.d_next[35] ),
    .Y(_04373_),
    .A2(\u_inv.d_reg[35] ));
 sg13g2_nor2_1 _34962_ (.A(_04354_),
    .B(_04373_),
    .Y(_04374_));
 sg13g2_a22oi_1 _34963_ (.Y(_04375_),
    .B1(\u_inv.d_reg[36] ),
    .B2(\u_inv.d_next[36] ),
    .A2(\u_inv.d_reg[37] ),
    .A1(\u_inv.d_next[37] ));
 sg13g2_nor2_1 _34964_ (.A(_04341_),
    .B(_04375_),
    .Y(_04376_));
 sg13g2_o21ai_1 _34965_ (.B1(_04351_),
    .Y(_04377_),
    .A1(_04341_),
    .A2(_04375_));
 sg13g2_a21oi_1 _34966_ (.A1(_18170_),
    .A2(_18576_),
    .Y(_04378_),
    .B1(_04349_));
 sg13g2_a22oi_1 _34967_ (.Y(_04379_),
    .B1(_04377_),
    .B2(_04378_),
    .A2(\u_inv.d_reg[39] ),
    .A1(\u_inv.d_next[39] ));
 sg13g2_nor2b_1 _34968_ (.A(_04374_),
    .B_N(_04379_),
    .Y(_04380_));
 sg13g2_o21ai_1 _34969_ (.B1(_04379_),
    .Y(_04381_),
    .A1(_04354_),
    .A2(_04373_));
 sg13g2_a22oi_1 _34970_ (.Y(_04382_),
    .B1(\u_inv.d_reg[44] ),
    .B2(\u_inv.d_next[44] ),
    .A2(\u_inv.d_reg[45] ),
    .A1(\u_inv.d_next[45] ));
 sg13g2_or2_1 _34971_ (.X(_04383_),
    .B(_04382_),
    .A(_04181_));
 sg13g2_o21ai_1 _34972_ (.B1(_04188_),
    .Y(_04384_),
    .A1(_04181_),
    .A2(_04382_));
 sg13g2_nor2b_1 _34973_ (.A(_04185_),
    .B_N(_04186_),
    .Y(_04385_));
 sg13g2_a22oi_1 _34974_ (.Y(_04386_),
    .B1(_04384_),
    .B2(_04385_),
    .A2(\u_inv.d_reg[47] ),
    .A1(\u_inv.d_next[47] ));
 sg13g2_a22oi_1 _34975_ (.Y(_04387_),
    .B1(\u_inv.d_reg[40] ),
    .B2(\u_inv.d_next[40] ),
    .A2(\u_inv.d_reg[41] ),
    .A1(\u_inv.d_next[41] ));
 sg13g2_nor2_1 _34976_ (.A(_04196_),
    .B(_04387_),
    .Y(_04388_));
 sg13g2_o21ai_1 _34977_ (.B1(_04192_),
    .Y(_04389_),
    .A1(_04196_),
    .A2(_04387_));
 sg13g2_a21oi_1 _34978_ (.A1(_18169_),
    .A2(_18572_),
    .Y(_04390_),
    .B1(_04191_));
 sg13g2_a22oi_1 _34979_ (.Y(_04391_),
    .B1(_04389_),
    .B2(_04390_),
    .A2(\u_inv.d_reg[43] ),
    .A1(\u_inv.d_next[43] ));
 sg13g2_o21ai_1 _34980_ (.B1(_04386_),
    .Y(_04392_),
    .A1(_04190_),
    .A2(_04391_));
 sg13g2_a21o_2 _34981_ (.A2(_04381_),
    .A1(_04201_),
    .B1(_04392_),
    .X(_04393_));
 sg13g2_inv_1 _34982_ (.Y(_04394_),
    .A(_04393_));
 sg13g2_a21o_1 _34983_ (.A2(_04393_),
    .A1(_04154_),
    .B1(_04178_),
    .X(_04395_));
 sg13g2_nor4_2 _34984_ (.A(_04159_),
    .B(_04163_),
    .C(_04164_),
    .Y(_04396_),
    .D(_04395_));
 sg13g2_and3_1 _34985_ (.X(_04397_),
    .A(_04154_),
    .B(_04201_),
    .C(_04366_));
 sg13g2_o21ai_1 _34986_ (.B1(_04397_),
    .Y(_04398_),
    .A1(_04339_),
    .A2(_04337_));
 sg13g2_nand2_1 _34987_ (.Y(_04399_),
    .A(_04396_),
    .B(net1071));
 sg13g2_and2_1 _34988_ (.A(_04396_),
    .B(net1071),
    .X(_04400_));
 sg13g2_xor2_1 _34989_ (.B(\u_inv.d_reg[64] ),
    .A(\u_inv.d_next[64] ),
    .X(_04401_));
 sg13g2_nand2_1 _34990_ (.Y(_04402_),
    .A(_04024_),
    .B(_04401_));
 sg13g2_nor3_1 _34991_ (.A(_04029_),
    .B(_04031_),
    .C(_04402_),
    .Y(_04403_));
 sg13g2_inv_1 _34992_ (.Y(_04404_),
    .A(_04403_));
 sg13g2_and3_2 _34993_ (.X(_04405_),
    .A(_04019_),
    .B(_04061_),
    .C(_04403_));
 sg13g2_inv_1 _34994_ (.Y(_04406_),
    .A(_04405_));
 sg13g2_nand2b_2 _34995_ (.Y(_04407_),
    .B(_04405_),
    .A_N(_04003_));
 sg13g2_o21ai_1 _34996_ (.B1(_04098_),
    .Y(_04408_),
    .A1(_04400_),
    .A2(_04407_));
 sg13g2_xnor2_1 _34997_ (.Y(_04409_),
    .A(\u_inv.d_next[96] ),
    .B(\u_inv.d_reg[96] ));
 sg13g2_nor2_2 _34998_ (.A(_03923_),
    .B(_04409_),
    .Y(_04410_));
 sg13g2_nand4_1 _34999_ (.B(_03914_),
    .C(_03930_),
    .A(_03901_),
    .Y(_04411_),
    .D(_04410_));
 sg13g2_inv_1 _35000_ (.Y(_04412_),
    .A(_04411_));
 sg13g2_or4_1 _35001_ (.A(_03819_),
    .B(_03824_),
    .C(_03827_),
    .D(_03874_),
    .X(_04413_));
 sg13g2_nor3_1 _35002_ (.A(_03955_),
    .B(_04411_),
    .C(_04413_),
    .Y(_04414_));
 sg13g2_inv_1 _35003_ (.Y(_04415_),
    .A(_04414_));
 sg13g2_o21ai_1 _35004_ (.B1(_03839_),
    .Y(_04416_),
    .A1(_04098_),
    .A2(_04415_));
 sg13g2_nand2b_1 _35005_ (.Y(_04417_),
    .B(_04414_),
    .A_N(_04407_));
 sg13g2_a21oi_1 _35006_ (.A1(_04396_),
    .A2(net1070),
    .Y(_04418_),
    .B1(_04417_));
 sg13g2_nand2b_1 _35007_ (.Y(_04419_),
    .B(_03950_),
    .A_N(_03955_));
 sg13g2_a21oi_1 _35008_ (.A1(_03873_),
    .A2(_04419_),
    .Y(_04420_),
    .B1(_04413_));
 sg13g2_nor3_2 _35009_ (.A(_04416_),
    .B(_04420_),
    .C(_04418_),
    .Y(_04421_));
 sg13g2_or3_1 _35010_ (.A(_04416_),
    .B(_04418_),
    .C(_04420_),
    .X(_04422_));
 sg13g2_xor2_1 _35011_ (.B(\u_inv.d_reg[151] ),
    .A(\u_inv.d_next[151] ),
    .X(_04423_));
 sg13g2_xnor2_1 _35012_ (.Y(_04424_),
    .A(\u_inv.d_next[151] ),
    .B(\u_inv.d_reg[151] ));
 sg13g2_nand2_1 _35013_ (.Y(_04425_),
    .A(\u_inv.d_next[150] ),
    .B(\u_inv.d_reg[150] ));
 sg13g2_xor2_1 _35014_ (.B(\u_inv.d_reg[150] ),
    .A(\u_inv.d_next[150] ),
    .X(_04426_));
 sg13g2_xnor2_1 _35015_ (.Y(_04427_),
    .A(\u_inv.d_next[150] ),
    .B(\u_inv.d_reg[150] ));
 sg13g2_nand2_1 _35016_ (.Y(_04428_),
    .A(_04423_),
    .B(_04426_));
 sg13g2_xnor2_1 _35017_ (.Y(_04429_),
    .A(\u_inv.d_next[149] ),
    .B(\u_inv.d_reg[149] ));
 sg13g2_nand2_1 _35018_ (.Y(_04430_),
    .A(\u_inv.d_next[148] ),
    .B(\u_inv.d_reg[148] ));
 sg13g2_xnor2_1 _35019_ (.Y(_04431_),
    .A(\u_inv.d_next[148] ),
    .B(\u_inv.d_reg[148] ));
 sg13g2_inv_1 _35020_ (.Y(_04432_),
    .A(_04431_));
 sg13g2_nor2_1 _35021_ (.A(_04429_),
    .B(_04431_),
    .Y(_04433_));
 sg13g2_nor2b_1 _35022_ (.A(_04428_),
    .B_N(_04433_),
    .Y(_04434_));
 sg13g2_nor2_1 _35023_ (.A(\u_inv.d_next[147] ),
    .B(\u_inv.d_reg[147] ),
    .Y(_04435_));
 sg13g2_xor2_1 _35024_ (.B(\u_inv.d_reg[147] ),
    .A(\u_inv.d_next[147] ),
    .X(_04436_));
 sg13g2_xnor2_1 _35025_ (.Y(_04437_),
    .A(\u_inv.d_next[147] ),
    .B(\u_inv.d_reg[147] ));
 sg13g2_xnor2_1 _35026_ (.Y(_04438_),
    .A(\u_inv.d_next[146] ),
    .B(\u_inv.d_reg[146] ));
 sg13g2_nor2_1 _35027_ (.A(_04437_),
    .B(_04438_),
    .Y(_04439_));
 sg13g2_inv_1 _35028_ (.Y(_04440_),
    .A(_04439_));
 sg13g2_nor2b_1 _35029_ (.A(\u_inv.d_next[145] ),
    .B_N(\u_inv.d_reg[145] ),
    .Y(_04441_));
 sg13g2_nand2b_1 _35030_ (.Y(_04442_),
    .B(\u_inv.d_next[145] ),
    .A_N(\u_inv.d_reg[145] ));
 sg13g2_nor2b_1 _35031_ (.A(_04441_),
    .B_N(_04442_),
    .Y(_04443_));
 sg13g2_xor2_1 _35032_ (.B(\u_inv.d_reg[145] ),
    .A(\u_inv.d_next[145] ),
    .X(_04444_));
 sg13g2_nand2_1 _35033_ (.Y(_04445_),
    .A(\u_inv.d_next[144] ),
    .B(\u_inv.d_reg[144] ));
 sg13g2_xor2_1 _35034_ (.B(\u_inv.d_reg[144] ),
    .A(\u_inv.d_next[144] ),
    .X(_04446_));
 sg13g2_inv_1 _35035_ (.Y(_04447_),
    .A(_04446_));
 sg13g2_nand2_1 _35036_ (.Y(_04448_),
    .A(_04444_),
    .B(_04446_));
 sg13g2_nand4_1 _35037_ (.B(_04439_),
    .C(_04444_),
    .A(_04434_),
    .Y(_04449_),
    .D(_04446_));
 sg13g2_nand2_1 _35038_ (.Y(_04450_),
    .A(\u_inv.d_next[158] ),
    .B(\u_inv.d_reg[158] ));
 sg13g2_xnor2_1 _35039_ (.Y(_04451_),
    .A(\u_inv.d_next[158] ),
    .B(\u_inv.d_reg[158] ));
 sg13g2_xnor2_1 _35040_ (.Y(_04452_),
    .A(\u_inv.d_next[159] ),
    .B(\u_inv.d_reg[159] ));
 sg13g2_nor2_1 _35041_ (.A(_04451_),
    .B(_04452_),
    .Y(_04453_));
 sg13g2_nor2_1 _35042_ (.A(\u_inv.d_next[157] ),
    .B(\u_inv.d_reg[157] ),
    .Y(_04454_));
 sg13g2_xor2_1 _35043_ (.B(\u_inv.d_reg[157] ),
    .A(\u_inv.d_next[157] ),
    .X(_04455_));
 sg13g2_xnor2_1 _35044_ (.Y(_04456_),
    .A(\u_inv.d_next[157] ),
    .B(\u_inv.d_reg[157] ));
 sg13g2_nand2_1 _35045_ (.Y(_04457_),
    .A(\u_inv.d_next[156] ),
    .B(\u_inv.d_reg[156] ));
 sg13g2_xor2_1 _35046_ (.B(\u_inv.d_reg[156] ),
    .A(\u_inv.d_next[156] ),
    .X(_04458_));
 sg13g2_and2_1 _35047_ (.A(_04455_),
    .B(_04458_),
    .X(_04459_));
 sg13g2_nand2_1 _35048_ (.Y(_04460_),
    .A(_04453_),
    .B(_04459_));
 sg13g2_nor2_1 _35049_ (.A(\u_inv.d_next[155] ),
    .B(\u_inv.d_reg[155] ),
    .Y(_04461_));
 sg13g2_nand2_2 _35050_ (.Y(_04462_),
    .A(\u_inv.d_next[155] ),
    .B(\u_inv.d_reg[155] ));
 sg13g2_nor2b_1 _35051_ (.A(_04461_),
    .B_N(_04462_),
    .Y(_04463_));
 sg13g2_nand2b_2 _35052_ (.Y(_04464_),
    .B(_04462_),
    .A_N(_04461_));
 sg13g2_nand2_2 _35053_ (.Y(_04465_),
    .A(\u_inv.d_next[154] ),
    .B(\u_inv.d_reg[154] ));
 sg13g2_xor2_1 _35054_ (.B(\u_inv.d_reg[154] ),
    .A(\u_inv.d_next[154] ),
    .X(_04466_));
 sg13g2_nand2_1 _35055_ (.Y(_04467_),
    .A(_04463_),
    .B(_04466_));
 sg13g2_nand2_1 _35056_ (.Y(_04468_),
    .A(\u_inv.d_next[153] ),
    .B(\u_inv.d_reg[153] ));
 sg13g2_nor2_1 _35057_ (.A(\u_inv.d_next[153] ),
    .B(\u_inv.d_reg[153] ),
    .Y(_04469_));
 sg13g2_xnor2_1 _35058_ (.Y(_04470_),
    .A(\u_inv.d_next[153] ),
    .B(\u_inv.d_reg[153] ));
 sg13g2_nand2_1 _35059_ (.Y(_04471_),
    .A(\u_inv.d_next[152] ),
    .B(\u_inv.d_reg[152] ));
 sg13g2_xnor2_1 _35060_ (.Y(_04472_),
    .A(\u_inv.d_next[152] ),
    .B(\u_inv.d_reg[152] ));
 sg13g2_nor2_1 _35061_ (.A(_04470_),
    .B(_04472_),
    .Y(_04473_));
 sg13g2_nor4_1 _35062_ (.A(_04460_),
    .B(_04467_),
    .C(_04470_),
    .D(_04472_),
    .Y(_04474_));
 sg13g2_nand2b_2 _35063_ (.Y(_04475_),
    .B(_04474_),
    .A_N(_04449_));
 sg13g2_xor2_1 _35064_ (.B(\u_inv.d_reg[143] ),
    .A(\u_inv.d_next[143] ),
    .X(_04476_));
 sg13g2_nand2_1 _35065_ (.Y(_04477_),
    .A(\u_inv.d_next[142] ),
    .B(\u_inv.d_reg[142] ));
 sg13g2_nor2_1 _35066_ (.A(\u_inv.d_next[142] ),
    .B(\u_inv.d_reg[142] ),
    .Y(_04478_));
 sg13g2_xor2_1 _35067_ (.B(\u_inv.d_reg[142] ),
    .A(\u_inv.d_next[142] ),
    .X(_04479_));
 sg13g2_xor2_1 _35068_ (.B(\u_inv.d_reg[141] ),
    .A(\u_inv.d_next[141] ),
    .X(_04480_));
 sg13g2_and2_1 _35069_ (.A(\u_inv.d_next[140] ),
    .B(\u_inv.d_reg[140] ),
    .X(_04481_));
 sg13g2_xor2_1 _35070_ (.B(\u_inv.d_reg[140] ),
    .A(\u_inv.d_next[140] ),
    .X(_04482_));
 sg13g2_and2_1 _35071_ (.A(_04480_),
    .B(_04482_),
    .X(_04483_));
 sg13g2_and3_1 _35072_ (.X(_04484_),
    .A(_04476_),
    .B(_04479_),
    .C(_04483_));
 sg13g2_xor2_1 _35073_ (.B(\u_inv.d_reg[139] ),
    .A(\u_inv.d_next[139] ),
    .X(_04485_));
 sg13g2_xnor2_1 _35074_ (.Y(_04486_),
    .A(\u_inv.d_next[139] ),
    .B(\u_inv.d_reg[139] ));
 sg13g2_and2_1 _35075_ (.A(\u_inv.d_next[138] ),
    .B(\u_inv.d_reg[138] ),
    .X(_04487_));
 sg13g2_xor2_1 _35076_ (.B(\u_inv.d_reg[138] ),
    .A(\u_inv.d_next[138] ),
    .X(_04488_));
 sg13g2_and2_1 _35077_ (.A(_04485_),
    .B(_04488_),
    .X(_04489_));
 sg13g2_nand2_1 _35078_ (.Y(_04490_),
    .A(_04485_),
    .B(_04488_));
 sg13g2_xnor2_1 _35079_ (.Y(_04491_),
    .A(\u_inv.d_next[137] ),
    .B(\u_inv.d_reg[137] ));
 sg13g2_nand2_1 _35080_ (.Y(_04492_),
    .A(\u_inv.d_next[136] ),
    .B(\u_inv.d_reg[136] ));
 sg13g2_xnor2_1 _35081_ (.Y(_04493_),
    .A(\u_inv.d_next[136] ),
    .B(\u_inv.d_reg[136] ));
 sg13g2_nor2_1 _35082_ (.A(_04491_),
    .B(_04493_),
    .Y(_04494_));
 sg13g2_nand3_1 _35083_ (.B(_04489_),
    .C(_04494_),
    .A(_04484_),
    .Y(_04495_));
 sg13g2_nor2_1 _35084_ (.A(\u_inv.d_next[135] ),
    .B(\u_inv.d_reg[135] ),
    .Y(_04496_));
 sg13g2_xor2_1 _35085_ (.B(\u_inv.d_reg[135] ),
    .A(\u_inv.d_next[135] ),
    .X(_04497_));
 sg13g2_xnor2_1 _35086_ (.Y(_04498_),
    .A(\u_inv.d_next[135] ),
    .B(\u_inv.d_reg[135] ));
 sg13g2_nand2_1 _35087_ (.Y(_04499_),
    .A(\u_inv.d_next[134] ),
    .B(\u_inv.d_reg[134] ));
 sg13g2_xor2_1 _35088_ (.B(\u_inv.d_reg[134] ),
    .A(\u_inv.d_next[134] ),
    .X(_04500_));
 sg13g2_xnor2_1 _35089_ (.Y(_04501_),
    .A(\u_inv.d_next[134] ),
    .B(\u_inv.d_reg[134] ));
 sg13g2_xnor2_1 _35090_ (.Y(_04502_),
    .A(\u_inv.d_next[133] ),
    .B(\u_inv.d_reg[133] ));
 sg13g2_xor2_1 _35091_ (.B(\u_inv.d_reg[133] ),
    .A(\u_inv.d_next[133] ),
    .X(_04503_));
 sg13g2_and2_1 _35092_ (.A(\u_inv.d_next[132] ),
    .B(\u_inv.d_reg[132] ),
    .X(_04504_));
 sg13g2_xor2_1 _35093_ (.B(\u_inv.d_reg[132] ),
    .A(\u_inv.d_next[132] ),
    .X(_04505_));
 sg13g2_xnor2_1 _35094_ (.Y(_04506_),
    .A(\u_inv.d_next[132] ),
    .B(\u_inv.d_reg[132] ));
 sg13g2_nand2_1 _35095_ (.Y(_04507_),
    .A(_04503_),
    .B(_04505_));
 sg13g2_nor3_1 _35096_ (.A(_04498_),
    .B(_04501_),
    .C(_04507_),
    .Y(_04508_));
 sg13g2_nand2_1 _35097_ (.Y(_04509_),
    .A(net7296),
    .B(net7289));
 sg13g2_xor2_1 _35098_ (.B(net7289),
    .A(net7296),
    .X(_04510_));
 sg13g2_xnor2_1 _35099_ (.Y(_04511_),
    .A(net7296),
    .B(net7289));
 sg13g2_xnor2_1 _35100_ (.Y(_04512_),
    .A(\u_inv.d_next[131] ),
    .B(\u_inv.d_reg[131] ));
 sg13g2_xor2_1 _35101_ (.B(\u_inv.d_reg[131] ),
    .A(\u_inv.d_next[131] ),
    .X(_04513_));
 sg13g2_nor2b_1 _35102_ (.A(\u_inv.d_next[129] ),
    .B_N(\u_inv.d_reg[129] ),
    .Y(_04514_));
 sg13g2_nand2b_1 _35103_ (.Y(_04515_),
    .B(\u_inv.d_next[129] ),
    .A_N(\u_inv.d_reg[129] ));
 sg13g2_xnor2_1 _35104_ (.Y(_04516_),
    .A(\u_inv.d_next[129] ),
    .B(\u_inv.d_reg[129] ));
 sg13g2_nand2b_1 _35105_ (.Y(_04517_),
    .B(_04515_),
    .A_N(_04514_));
 sg13g2_o21ai_1 _35106_ (.B1(_04513_),
    .Y(_04518_),
    .A1(net7296),
    .A2(net7289));
 sg13g2_nor3_2 _35107_ (.A(_04511_),
    .B(_04512_),
    .C(_04516_),
    .Y(_04519_));
 sg13g2_nand2_1 _35108_ (.Y(_04520_),
    .A(\u_inv.d_next[128] ),
    .B(\u_inv.d_reg[128] ));
 sg13g2_xor2_1 _35109_ (.B(\u_inv.d_reg[128] ),
    .A(\u_inv.d_next[128] ),
    .X(_04521_));
 sg13g2_inv_1 _35110_ (.Y(_04522_),
    .A(net6994));
 sg13g2_and3_2 _35111_ (.X(_04523_),
    .A(_04508_),
    .B(_04519_),
    .C(net6994));
 sg13g2_nand3_1 _35112_ (.B(_04519_),
    .C(net6994),
    .A(_04508_),
    .Y(_04524_));
 sg13g2_nor3_2 _35113_ (.A(_04475_),
    .B(_04495_),
    .C(_04524_),
    .Y(_04525_));
 sg13g2_nand2_1 _35114_ (.Y(_04526_),
    .A(\u_inv.d_next[131] ),
    .B(\u_inv.d_reg[131] ));
 sg13g2_nor2_1 _35115_ (.A(_04516_),
    .B(_04520_),
    .Y(_04527_));
 sg13g2_a21oi_1 _35116_ (.A1(\u_inv.d_next[129] ),
    .A2(\u_inv.d_reg[129] ),
    .Y(_04528_),
    .B1(_04527_));
 sg13g2_a221oi_1 _35117_ (.B2(\u_inv.d_next[129] ),
    .C1(_04527_),
    .B1(\u_inv.d_reg[129] ),
    .A1(net7296),
    .Y(_04529_),
    .A2(net7289));
 sg13g2_o21ai_1 _35118_ (.B1(_04526_),
    .Y(_04530_),
    .A1(_04518_),
    .A2(_04529_));
 sg13g2_and2_1 _35119_ (.A(\u_inv.d_next[133] ),
    .B(\u_inv.d_reg[133] ),
    .X(_04531_));
 sg13g2_a21oi_1 _35120_ (.A1(_04503_),
    .A2(_04504_),
    .Y(_04532_),
    .B1(_04531_));
 sg13g2_nand3b_1 _35121_ (.B(_04500_),
    .C(_04497_),
    .Y(_04533_),
    .A_N(_04532_));
 sg13g2_o21ai_1 _35122_ (.B1(_04533_),
    .Y(_04534_),
    .A1(_04496_),
    .A2(_04499_));
 sg13g2_a221oi_1 _35123_ (.B2(_04530_),
    .C1(_04534_),
    .B1(_04508_),
    .A1(\u_inv.d_next[135] ),
    .Y(_04535_),
    .A2(\u_inv.d_reg[135] ));
 sg13g2_inv_1 _35124_ (.Y(_04536_),
    .A(_04535_));
 sg13g2_or2_1 _35125_ (.X(_04537_),
    .B(_04535_),
    .A(_04495_));
 sg13g2_a21oi_1 _35126_ (.A1(\u_inv.d_next[141] ),
    .A2(\u_inv.d_reg[141] ),
    .Y(_04538_),
    .B1(_04481_));
 sg13g2_a21oi_1 _35127_ (.A1(_18131_),
    .A2(_18473_),
    .Y(_04539_),
    .B1(_04538_));
 sg13g2_nand3_1 _35128_ (.B(_04479_),
    .C(_04539_),
    .A(_04476_),
    .Y(_04540_));
 sg13g2_a21oi_1 _35129_ (.A1(_18130_),
    .A2(_18471_),
    .Y(_04541_),
    .B1(_04477_));
 sg13g2_nor2_1 _35130_ (.A(_04491_),
    .B(_04492_),
    .Y(_04542_));
 sg13g2_a21oi_1 _35131_ (.A1(\u_inv.d_next[137] ),
    .A2(\u_inv.d_reg[137] ),
    .Y(_04543_),
    .B1(_04542_));
 sg13g2_a21oi_1 _35132_ (.A1(\u_inv.d_next[139] ),
    .A2(\u_inv.d_reg[139] ),
    .Y(_04544_),
    .B1(_04487_));
 sg13g2_inv_1 _35133_ (.Y(_04545_),
    .A(_04544_));
 sg13g2_o21ai_1 _35134_ (.B1(_04545_),
    .Y(_04546_),
    .A1(\u_inv.d_next[139] ),
    .A2(\u_inv.d_reg[139] ));
 sg13g2_inv_1 _35135_ (.Y(_04547_),
    .A(_04546_));
 sg13g2_o21ai_1 _35136_ (.B1(_04546_),
    .Y(_04548_),
    .A1(_04490_),
    .A2(_04543_));
 sg13g2_a221oi_1 _35137_ (.B2(_04548_),
    .C1(_04541_),
    .B1(_04484_),
    .A1(\u_inv.d_next[143] ),
    .Y(_04549_),
    .A2(\u_inv.d_reg[143] ));
 sg13g2_and3_2 _35138_ (.X(_04550_),
    .A(_04537_),
    .B(_04540_),
    .C(_04549_));
 sg13g2_o21ai_1 _35139_ (.B1(_04468_),
    .Y(_04551_),
    .A1(_04469_),
    .A2(_04471_));
 sg13g2_inv_1 _35140_ (.Y(_04552_),
    .A(_04551_));
 sg13g2_nor2_1 _35141_ (.A(_04467_),
    .B(_04552_),
    .Y(_04553_));
 sg13g2_a21oi_2 _35142_ (.B1(_04461_),
    .Y(_04554_),
    .A2(_04465_),
    .A1(_04462_));
 sg13g2_nor2_1 _35143_ (.A(_04553_),
    .B(_04554_),
    .Y(_04555_));
 sg13g2_a22oi_1 _35144_ (.Y(_04556_),
    .B1(\u_inv.d_reg[156] ),
    .B2(\u_inv.d_next[156] ),
    .A2(\u_inv.d_reg[157] ),
    .A1(\u_inv.d_next[157] ));
 sg13g2_nor2_1 _35145_ (.A(_04454_),
    .B(_04556_),
    .Y(_04557_));
 sg13g2_or2_1 _35146_ (.X(_04558_),
    .B(_04556_),
    .A(_04454_));
 sg13g2_a21oi_1 _35147_ (.A1(_18126_),
    .A2(_18455_),
    .Y(_04559_),
    .B1(_04450_));
 sg13g2_a221oi_1 _35148_ (.B2(_04557_),
    .C1(_04559_),
    .B1(_04453_),
    .A1(\u_inv.d_next[159] ),
    .Y(_04560_),
    .A2(\u_inv.d_reg[159] ));
 sg13g2_o21ai_1 _35149_ (.B1(_04560_),
    .Y(_04561_),
    .A1(_04460_),
    .A2(_04555_));
 sg13g2_nand2b_1 _35150_ (.Y(_04562_),
    .B(_04444_),
    .A_N(_04445_));
 sg13g2_nand2_1 _35151_ (.Y(_04563_),
    .A(\u_inv.d_next[145] ),
    .B(\u_inv.d_reg[145] ));
 sg13g2_and2_1 _35152_ (.A(_04562_),
    .B(_04563_),
    .X(_04564_));
 sg13g2_a22oi_1 _35153_ (.Y(_04565_),
    .B1(\u_inv.d_reg[146] ),
    .B2(\u_inv.d_next[146] ),
    .A2(\u_inv.d_reg[147] ),
    .A1(\u_inv.d_next[147] ));
 sg13g2_or2_1 _35154_ (.X(_04566_),
    .B(_04565_),
    .A(_04435_));
 sg13g2_nor2_1 _35155_ (.A(_04435_),
    .B(_04565_),
    .Y(_04567_));
 sg13g2_o21ai_1 _35156_ (.B1(_04566_),
    .Y(_04568_),
    .A1(_04440_),
    .A2(_04564_));
 sg13g2_a21oi_1 _35157_ (.A1(_18127_),
    .A2(_18463_),
    .Y(_04569_),
    .B1(_04425_));
 sg13g2_a22oi_1 _35158_ (.Y(_04570_),
    .B1(\u_inv.d_reg[148] ),
    .B2(\u_inv.d_next[148] ),
    .A2(\u_inv.d_reg[149] ),
    .A1(\u_inv.d_next[149] ));
 sg13g2_a21o_1 _35159_ (.A2(_18465_),
    .A1(_18129_),
    .B1(_04570_),
    .X(_04571_));
 sg13g2_a221oi_1 _35160_ (.B2(_04568_),
    .C1(_04569_),
    .B1(_04434_),
    .A1(\u_inv.d_next[151] ),
    .Y(_04572_),
    .A2(\u_inv.d_reg[151] ));
 sg13g2_o21ai_1 _35161_ (.B1(_04572_),
    .Y(_04573_),
    .A1(_04428_),
    .A2(_04571_));
 sg13g2_a21oi_1 _35162_ (.A1(_04474_),
    .A2(_04573_),
    .Y(_04574_),
    .B1(_04561_));
 sg13g2_o21ai_1 _35163_ (.B1(_04574_),
    .Y(_04575_),
    .A1(_04475_),
    .A2(_04550_));
 sg13g2_nand3_1 _35164_ (.B(_03761_),
    .C(_03766_),
    .A(_03754_),
    .Y(_04576_));
 sg13g2_o21ai_1 _35165_ (.B1(_03785_),
    .Y(_04577_),
    .A1(_03778_),
    .A2(_04576_));
 sg13g2_nor2_2 _35166_ (.A(_03739_),
    .B(_04576_),
    .Y(_04578_));
 sg13g2_inv_1 _35167_ (.Y(_04579_),
    .A(_04578_));
 sg13g2_nor4_1 _35168_ (.A(_03673_),
    .B(_03702_),
    .C(_03715_),
    .D(_04579_),
    .Y(_04580_));
 sg13g2_a221oi_1 _35169_ (.B2(_04575_),
    .C1(_04577_),
    .B1(_04580_),
    .A1(_03807_),
    .Y(_04581_),
    .A2(_04578_));
 sg13g2_nand2_1 _35170_ (.Y(_04582_),
    .A(_04525_),
    .B(_04580_));
 sg13g2_o21ai_1 _35171_ (.B1(_04581_),
    .Y(_04583_),
    .A1(_04582_),
    .A2(net1109));
 sg13g2_xor2_1 _35172_ (.B(\u_inv.d_reg[192] ),
    .A(\u_inv.d_next[192] ),
    .X(_04584_));
 sg13g2_and3_2 _35173_ (.X(_04585_),
    .A(_03412_),
    .B(_03416_),
    .C(_04584_));
 sg13g2_inv_1 _35174_ (.Y(_04586_),
    .A(_04585_));
 sg13g2_nor3_1 _35175_ (.A(_03428_),
    .B(_03480_),
    .C(_04586_),
    .Y(_04587_));
 sg13g2_and2_1 _35176_ (.A(_03659_),
    .B(_04587_),
    .X(_04588_));
 sg13g2_a21o_2 _35177_ (.A2(_04588_),
    .A1(net1080),
    .B1(_03661_),
    .X(_04589_));
 sg13g2_nand3_1 _35178_ (.B(_03356_),
    .C(_04589_),
    .A(net7327),
    .Y(_04590_));
 sg13g2_o21ai_1 _35179_ (.B1(net6216),
    .Y(_04591_),
    .A1(net7327),
    .A2(\u_inv.d_next[256] ));
 sg13g2_a21oi_1 _35180_ (.A1(_18100_),
    .A2(_18358_),
    .Y(_04592_),
    .B1(_04591_));
 sg13g2_and2_1 _35181_ (.A(_04590_),
    .B(_04592_),
    .X(_04593_));
 sg13g2_nor2_1 _35182_ (.A(_03574_),
    .B(_03577_),
    .Y(_04594_));
 sg13g2_nor4_1 _35183_ (.A(_03566_),
    .B(_03570_),
    .C(_03574_),
    .D(_03577_),
    .Y(_04595_));
 sg13g2_nand2_1 _35184_ (.Y(_04596_),
    .A(_03589_),
    .B(_03591_));
 sg13g2_nand2b_2 _35185_ (.Y(_04597_),
    .B(_03586_),
    .A_N(_03583_));
 sg13g2_nor2_1 _35186_ (.A(_04596_),
    .B(_04597_),
    .Y(_04598_));
 sg13g2_and2_1 _35187_ (.A(_04595_),
    .B(_04598_),
    .X(_04599_));
 sg13g2_nor2_1 _35188_ (.A(_03593_),
    .B(_03596_),
    .Y(_04600_));
 sg13g2_nor4_1 _35189_ (.A(_03593_),
    .B(_03596_),
    .C(_03601_),
    .D(_03603_),
    .Y(_04601_));
 sg13g2_nor2_1 _35190_ (.A(_03598_),
    .B(_03614_),
    .Y(_04602_));
 sg13g2_and3_1 _35191_ (.X(_04603_),
    .A(_03608_),
    .B(_03609_),
    .C(_04602_));
 sg13g2_and2_1 _35192_ (.A(_04601_),
    .B(_04603_),
    .X(_04604_));
 sg13g2_nand2_1 _35193_ (.Y(_04605_),
    .A(_04599_),
    .B(_04604_));
 sg13g2_nor2_1 _35194_ (.A(_03511_),
    .B(_03514_),
    .Y(_04606_));
 sg13g2_and2_1 _35195_ (.A(_03518_),
    .B(_03520_),
    .X(_04607_));
 sg13g2_nand2_1 _35196_ (.Y(_04608_),
    .A(_04606_),
    .B(_04607_));
 sg13g2_and2_1 _35197_ (.A(_03534_),
    .B(_03536_),
    .X(_04609_));
 sg13g2_nand2_1 _35198_ (.Y(_04610_),
    .A(_03526_),
    .B(_03529_));
 sg13g2_nand3_1 _35199_ (.B(_03529_),
    .C(_04609_),
    .A(_03526_),
    .Y(_04611_));
 sg13g2_nor2_1 _35200_ (.A(_04608_),
    .B(_04611_),
    .Y(_04612_));
 sg13g2_nand2_1 _35201_ (.Y(_04613_),
    .A(_03546_),
    .B(_03549_));
 sg13g2_nand4_1 _35202_ (.B(_03549_),
    .C(_03552_),
    .A(_03546_),
    .Y(_04614_),
    .D(_03555_));
 sg13g2_nor2_1 _35203_ (.A(_03539_),
    .B(_03541_),
    .Y(_04615_));
 sg13g2_and2_1 _35204_ (.A(_03558_),
    .B(_03560_),
    .X(_04616_));
 sg13g2_nand2_1 _35205_ (.Y(_04617_),
    .A(_04615_),
    .B(_04616_));
 sg13g2_nor2_2 _35206_ (.A(_04614_),
    .B(_04617_),
    .Y(_04618_));
 sg13g2_nand2_2 _35207_ (.Y(_04619_),
    .A(_04612_),
    .B(_04618_));
 sg13g2_or2_1 _35208_ (.X(_04620_),
    .B(_04619_),
    .A(_04605_));
 sg13g2_and2_1 _35209_ (.A(_03432_),
    .B(_03434_),
    .X(_04621_));
 sg13g2_nand3_1 _35210_ (.B(_03439_),
    .C(_04621_),
    .A(_03437_),
    .Y(_04622_));
 sg13g2_nor2_1 _35211_ (.A(_03444_),
    .B(_03447_),
    .Y(_04623_));
 sg13g2_nor2_1 _35212_ (.A(_03449_),
    .B(_03452_),
    .Y(_04624_));
 sg13g2_nand2_1 _35213_ (.Y(_04625_),
    .A(_04623_),
    .B(_04624_));
 sg13g2_nor2_1 _35214_ (.A(_04622_),
    .B(_04625_),
    .Y(_04626_));
 sg13g2_nor2_1 _35215_ (.A(_03462_),
    .B(_03465_),
    .Y(_04627_));
 sg13g2_inv_1 _35216_ (.Y(_04628_),
    .A(_04627_));
 sg13g2_nor2_1 _35217_ (.A(_03456_),
    .B(_03459_),
    .Y(_04629_));
 sg13g2_and2_1 _35218_ (.A(_04627_),
    .B(_04629_),
    .X(_04630_));
 sg13g2_inv_1 _35219_ (.Y(_04631_),
    .A(_04630_));
 sg13g2_nor2_1 _35220_ (.A(_03469_),
    .B(_03470_),
    .Y(_04632_));
 sg13g2_nor2_2 _35221_ (.A(_03473_),
    .B(_03475_),
    .Y(_04633_));
 sg13g2_and3_2 _35222_ (.X(_04634_),
    .A(_04630_),
    .B(_04632_),
    .C(_04633_));
 sg13g2_nand2_1 _35223_ (.Y(_04635_),
    .A(_04626_),
    .B(_04634_));
 sg13g2_nor2_1 _35224_ (.A(_03357_),
    .B(_03360_),
    .Y(_04636_));
 sg13g2_and2_1 _35225_ (.A(_03367_),
    .B(_03368_),
    .X(_04637_));
 sg13g2_and2_1 _35226_ (.A(_04636_),
    .B(_04637_),
    .X(_04638_));
 sg13g2_inv_1 _35227_ (.Y(_04639_),
    .A(_04638_));
 sg13g2_nand2_1 _35228_ (.Y(_04640_),
    .A(_03374_),
    .B(_03375_));
 sg13g2_or2_1 _35229_ (.X(_04641_),
    .B(_03385_),
    .A(_03383_));
 sg13g2_nor3_1 _35230_ (.A(_04639_),
    .B(_04640_),
    .C(_04641_),
    .Y(_04642_));
 sg13g2_nor2_1 _35231_ (.A(_03422_),
    .B(_03424_),
    .Y(_04643_));
 sg13g2_nor2_1 _35232_ (.A(_03389_),
    .B(_03392_),
    .Y(_04644_));
 sg13g2_and2_1 _35233_ (.A(_04643_),
    .B(_04644_),
    .X(_04645_));
 sg13g2_nand2_1 _35234_ (.Y(_04646_),
    .A(_04643_),
    .B(_04644_));
 sg13g2_nand2b_1 _35235_ (.Y(_04647_),
    .B(_03415_),
    .A_N(_04584_));
 sg13g2_nand2_1 _35236_ (.Y(_04648_),
    .A(_03409_),
    .B(_03411_));
 sg13g2_or2_1 _35237_ (.X(_04649_),
    .B(_04648_),
    .A(_04647_));
 sg13g2_nor2_1 _35238_ (.A(_04646_),
    .B(_04649_),
    .Y(_04650_));
 sg13g2_nand2_1 _35239_ (.Y(_04651_),
    .A(_04642_),
    .B(_04650_));
 sg13g2_or2_1 _35240_ (.X(_04652_),
    .B(_04651_),
    .A(_04635_));
 sg13g2_inv_1 _35241_ (.Y(_04653_),
    .A(_04652_));
 sg13g2_or2_1 _35242_ (.X(_04654_),
    .B(_04652_),
    .A(_04620_));
 sg13g2_nand2_1 _35243_ (.Y(_04655_),
    .A(\u_inv.d_next[198] ),
    .B(_18416_));
 sg13g2_nor2b_1 _35244_ (.A(\u_inv.d_reg[196] ),
    .B_N(\u_inv.d_next[196] ),
    .Y(_04656_));
 sg13g2_nor2b_1 _35245_ (.A(\u_inv.d_reg[197] ),
    .B_N(\u_inv.d_next[197] ),
    .Y(_04657_));
 sg13g2_a21o_1 _35246_ (.A2(_04656_),
    .A1(_03423_),
    .B1(_04657_),
    .X(_04658_));
 sg13g2_nor2_1 _35247_ (.A(_03389_),
    .B(_04655_),
    .Y(_04659_));
 sg13g2_a221oi_1 _35248_ (.B2(_04658_),
    .C1(_04659_),
    .B1(_04644_),
    .A1(\u_inv.d_next[199] ),
    .Y(_04660_),
    .A2(_18415_));
 sg13g2_inv_1 _35249_ (.Y(_04661_),
    .A(_04660_));
 sg13g2_nor2b_1 _35250_ (.A(\u_inv.d_reg[192] ),
    .B_N(\u_inv.d_next[192] ),
    .Y(_04662_));
 sg13g2_a21oi_1 _35251_ (.A1(_03413_),
    .A2(_04662_),
    .Y(_04663_),
    .B1(_03414_));
 sg13g2_nor2b_1 _35252_ (.A(\u_inv.d_reg[194] ),
    .B_N(\u_inv.d_next[194] ),
    .Y(_04664_));
 sg13g2_nand2_1 _35253_ (.Y(_04665_),
    .A(\u_inv.d_next[195] ),
    .B(_18419_));
 sg13g2_o21ai_1 _35254_ (.B1(_04665_),
    .Y(_04666_),
    .A1(_04648_),
    .A2(_04663_));
 sg13g2_a21oi_1 _35255_ (.A1(_03409_),
    .A2(_04664_),
    .Y(_04667_),
    .B1(_04666_));
 sg13g2_o21ai_1 _35256_ (.B1(_04660_),
    .Y(_04668_),
    .A1(_04646_),
    .A2(_04667_));
 sg13g2_nand2_1 _35257_ (.Y(_04669_),
    .A(_04642_),
    .B(_04668_));
 sg13g2_nand2_1 _35258_ (.Y(_04670_),
    .A(\u_inv.d_next[200] ),
    .B(_18414_));
 sg13g2_nor2_1 _35259_ (.A(_03383_),
    .B(_04670_),
    .Y(_04671_));
 sg13g2_a21oi_1 _35260_ (.A1(\u_inv.d_next[201] ),
    .A2(_18413_),
    .Y(_04672_),
    .B1(_04671_));
 sg13g2_nor2_1 _35261_ (.A(_18116_),
    .B(\u_inv.d_reg[203] ),
    .Y(_04673_));
 sg13g2_nor2b_1 _35262_ (.A(\u_inv.d_reg[202] ),
    .B_N(\u_inv.d_next[202] ),
    .Y(_04674_));
 sg13g2_a21oi_1 _35263_ (.A1(_03374_),
    .A2(_04674_),
    .Y(_04675_),
    .B1(_04673_));
 sg13g2_o21ai_1 _35264_ (.B1(_04675_),
    .Y(_04676_),
    .A1(_04640_),
    .A2(_04672_));
 sg13g2_nand2_1 _35265_ (.Y(_04677_),
    .A(\u_inv.d_next[204] ),
    .B(_18410_));
 sg13g2_nor2b_1 _35266_ (.A(_04677_),
    .B_N(_03367_),
    .Y(_04678_));
 sg13g2_a21oi_1 _35267_ (.A1(\u_inv.d_next[205] ),
    .A2(_18409_),
    .Y(_04679_),
    .B1(_04678_));
 sg13g2_nor2b_1 _35268_ (.A(_04679_),
    .B_N(_04636_),
    .Y(_04680_));
 sg13g2_nor2b_1 _35269_ (.A(\u_inv.d_reg[206] ),
    .B_N(\u_inv.d_next[206] ),
    .Y(_04681_));
 sg13g2_nand2b_1 _35270_ (.Y(_04682_),
    .B(_04681_),
    .A_N(_03357_));
 sg13g2_a221oi_1 _35271_ (.B2(_04676_),
    .C1(_04680_),
    .B1(_04638_),
    .A1(\u_inv.d_next[207] ),
    .Y(_04683_),
    .A2(_18407_));
 sg13g2_and3_1 _35272_ (.X(_04684_),
    .A(_04669_),
    .B(_04682_),
    .C(_04683_));
 sg13g2_nor2_1 _35273_ (.A(_04635_),
    .B(_04684_),
    .Y(_04685_));
 sg13g2_nor2b_1 _35274_ (.A(\u_inv.d_reg[208] ),
    .B_N(\u_inv.d_next[208] ),
    .Y(_04686_));
 sg13g2_nand2_1 _35275_ (.Y(_04687_),
    .A(_03474_),
    .B(_04686_));
 sg13g2_o21ai_1 _35276_ (.B1(_04687_),
    .Y(_04688_),
    .A1(_18114_),
    .A2(\u_inv.d_reg[209] ));
 sg13g2_nand2_1 _35277_ (.Y(_04689_),
    .A(\u_inv.d_next[210] ),
    .B(_18404_));
 sg13g2_nor2_1 _35278_ (.A(_03469_),
    .B(_04689_),
    .Y(_04690_));
 sg13g2_a221oi_1 _35279_ (.B2(_04688_),
    .C1(_04690_),
    .B1(_04632_),
    .A1(\u_inv.d_next[211] ),
    .Y(_04691_),
    .A2(_18403_));
 sg13g2_nor2b_1 _35280_ (.A(\u_inv.d_reg[212] ),
    .B_N(\u_inv.d_next[212] ),
    .Y(_04692_));
 sg13g2_nand2_1 _35281_ (.Y(_04693_),
    .A(_03463_),
    .B(_04692_));
 sg13g2_o21ai_1 _35282_ (.B1(_04693_),
    .Y(_04694_),
    .A1(_18112_),
    .A2(\u_inv.d_reg[213] ));
 sg13g2_nand2_1 _35283_ (.Y(_04695_),
    .A(\u_inv.d_next[214] ),
    .B(_18400_));
 sg13g2_nor2_1 _35284_ (.A(_03456_),
    .B(_04695_),
    .Y(_04696_));
 sg13g2_a221oi_1 _35285_ (.B2(_04694_),
    .C1(_04696_),
    .B1(_04629_),
    .A1(\u_inv.d_next[215] ),
    .Y(_04697_),
    .A2(_18399_));
 sg13g2_o21ai_1 _35286_ (.B1(_04697_),
    .Y(_04698_),
    .A1(_04631_),
    .A2(_04691_));
 sg13g2_nor2_1 _35287_ (.A(_18108_),
    .B(\u_inv.d_reg[223] ),
    .Y(_04699_));
 sg13g2_nand2_1 _35288_ (.Y(_04700_),
    .A(\u_inv.d_next[222] ),
    .B(_18392_));
 sg13g2_nor2b_1 _35289_ (.A(\u_inv.d_reg[220] ),
    .B_N(\u_inv.d_next[220] ),
    .Y(_04701_));
 sg13g2_nor2_1 _35290_ (.A(_18109_),
    .B(\u_inv.d_reg[221] ),
    .Y(_04702_));
 sg13g2_a21oi_1 _35291_ (.A1(_03432_),
    .A2(_04701_),
    .Y(_04703_),
    .B1(_04702_));
 sg13g2_o21ai_1 _35292_ (.B1(_04700_),
    .Y(_04704_),
    .A1(_03440_),
    .A2(_04703_));
 sg13g2_a221oi_1 _35293_ (.B2(_03437_),
    .C1(_04699_),
    .B1(_04704_),
    .A1(_04626_),
    .Y(_04705_),
    .A2(_04698_));
 sg13g2_nand2_1 _35294_ (.Y(_04706_),
    .A(\u_inv.d_next[216] ),
    .B(_18398_));
 sg13g2_nor2_1 _35295_ (.A(_03449_),
    .B(_04706_),
    .Y(_04707_));
 sg13g2_a21oi_1 _35296_ (.A1(\u_inv.d_next[217] ),
    .A2(_18397_),
    .Y(_04708_),
    .B1(_04707_));
 sg13g2_inv_1 _35297_ (.Y(_04709_),
    .A(_04708_));
 sg13g2_nor2_1 _35298_ (.A(_03444_),
    .B(_03446_),
    .Y(_04710_));
 sg13g2_a221oi_1 _35299_ (.B2(_04709_),
    .C1(_04710_),
    .B1(_04623_),
    .A1(\u_inv.d_next[219] ),
    .Y(_04711_),
    .A2(_18395_));
 sg13g2_o21ai_1 _35300_ (.B1(_04705_),
    .Y(_04712_),
    .A1(_04622_),
    .A2(_04711_));
 sg13g2_nor2_1 _35301_ (.A(_04685_),
    .B(_04712_),
    .Y(_04713_));
 sg13g2_inv_1 _35302_ (.Y(_04714_),
    .A(_04713_));
 sg13g2_or2_1 _35303_ (.X(_04715_),
    .B(_04713_),
    .A(_04620_));
 sg13g2_nand2_1 _35304_ (.Y(_04716_),
    .A(\u_inv.d_next[226] ),
    .B(_18388_));
 sg13g2_nor2b_1 _35305_ (.A(\u_inv.d_reg[224] ),
    .B_N(\u_inv.d_next[224] ),
    .Y(_04717_));
 sg13g2_nor2b_1 _35306_ (.A(\u_inv.d_reg[225] ),
    .B_N(\u_inv.d_next[225] ),
    .Y(_04718_));
 sg13g2_a21o_1 _35307_ (.A2(_04717_),
    .A1(_03560_),
    .B1(_04718_),
    .X(_04719_));
 sg13g2_nor2_1 _35308_ (.A(_03539_),
    .B(_04716_),
    .Y(_04720_));
 sg13g2_a221oi_1 _35309_ (.B2(_04719_),
    .C1(_04720_),
    .B1(_04615_),
    .A1(\u_inv.d_next[227] ),
    .Y(_04721_),
    .A2(_18387_));
 sg13g2_nor2b_1 _35310_ (.A(\u_inv.d_reg[231] ),
    .B_N(\u_inv.d_next[231] ),
    .Y(_04722_));
 sg13g2_nand2_1 _35311_ (.Y(_04723_),
    .A(\u_inv.d_next[230] ),
    .B(_18384_));
 sg13g2_nor2b_1 _35312_ (.A(\u_inv.d_reg[228] ),
    .B_N(\u_inv.d_next[228] ),
    .Y(_04724_));
 sg13g2_nor2b_1 _35313_ (.A(\u_inv.d_reg[229] ),
    .B_N(\u_inv.d_next[229] ),
    .Y(_04725_));
 sg13g2_a21o_1 _35314_ (.A2(_04724_),
    .A1(_03546_),
    .B1(_04725_),
    .X(_04726_));
 sg13g2_nand2_1 _35315_ (.Y(_04727_),
    .A(_03552_),
    .B(_04726_));
 sg13g2_nand2_1 _35316_ (.Y(_04728_),
    .A(_04723_),
    .B(_04727_));
 sg13g2_a21oi_1 _35317_ (.A1(_03555_),
    .A2(_04728_),
    .Y(_04729_),
    .B1(_04722_));
 sg13g2_o21ai_1 _35318_ (.B1(_04729_),
    .Y(_04730_),
    .A1(_04614_),
    .A2(_04721_));
 sg13g2_nor2b_1 _35319_ (.A(\u_inv.d_reg[236] ),
    .B_N(\u_inv.d_next[236] ),
    .Y(_04731_));
 sg13g2_nand2_1 _35320_ (.Y(_04732_),
    .A(_03518_),
    .B(_04731_));
 sg13g2_o21ai_1 _35321_ (.B1(_04732_),
    .Y(_04733_),
    .A1(_18106_),
    .A2(\u_inv.d_reg[237] ));
 sg13g2_nor2b_1 _35322_ (.A(\u_inv.d_reg[238] ),
    .B_N(\u_inv.d_next[238] ),
    .Y(_04734_));
 sg13g2_nand2_1 _35323_ (.Y(_04735_),
    .A(\u_inv.d_next[238] ),
    .B(_18376_));
 sg13g2_nor2b_1 _35324_ (.A(\u_inv.d_reg[235] ),
    .B_N(\u_inv.d_next[235] ),
    .Y(_04736_));
 sg13g2_nor2b_1 _35325_ (.A(\u_inv.d_reg[234] ),
    .B_N(\u_inv.d_next[234] ),
    .Y(_04737_));
 sg13g2_nand2_1 _35326_ (.Y(_04738_),
    .A(\u_inv.d_next[232] ),
    .B(_18382_));
 sg13g2_nand2_1 _35327_ (.Y(_04739_),
    .A(\u_inv.d_next[233] ),
    .B(_18381_));
 sg13g2_o21ai_1 _35328_ (.B1(_04739_),
    .Y(_04740_),
    .A1(_03525_),
    .A2(_04738_));
 sg13g2_inv_1 _35329_ (.Y(_04741_),
    .A(_04740_));
 sg13g2_a221oi_1 _35330_ (.B2(_04609_),
    .C1(_04736_),
    .B1(_04740_),
    .A1(_03534_),
    .Y(_04742_),
    .A2(_04737_));
 sg13g2_a22oi_1 _35331_ (.Y(_04743_),
    .B1(_04606_),
    .B2(_04733_),
    .A2(_18375_),
    .A1(\u_inv.d_next[239] ));
 sg13g2_o21ai_1 _35332_ (.B1(_04743_),
    .Y(_04744_),
    .A1(_04608_),
    .A2(_04742_));
 sg13g2_a221oi_1 _35333_ (.B2(_03512_),
    .C1(_04744_),
    .B1(_04734_),
    .A1(_04612_),
    .Y(_04745_),
    .A2(_04730_));
 sg13g2_or2_1 _35334_ (.X(_04746_),
    .B(_04745_),
    .A(_04605_));
 sg13g2_nand2_1 _35335_ (.Y(_04747_),
    .A(\u_inv.d_next[243] ),
    .B(_18371_));
 sg13g2_nor2_1 _35336_ (.A(_18105_),
    .B(\u_inv.d_reg[242] ),
    .Y(_04748_));
 sg13g2_nor2b_1 _35337_ (.A(net7288),
    .B_N(\u_inv.d_next[240] ),
    .Y(_04749_));
 sg13g2_nor2b_1 _35338_ (.A(\u_inv.d_reg[241] ),
    .B_N(\u_inv.d_next[241] ),
    .Y(_04750_));
 sg13g2_a21o_1 _35339_ (.A2(_04749_),
    .A1(_03599_),
    .B1(_04750_),
    .X(_04751_));
 sg13g2_a21oi_1 _35340_ (.A1(_03609_),
    .A2(_04751_),
    .Y(_04752_),
    .B1(_04748_));
 sg13g2_o21ai_1 _35341_ (.B1(_04747_),
    .Y(_04753_),
    .A1(_03607_),
    .A2(_04752_));
 sg13g2_nand2_1 _35342_ (.Y(_04754_),
    .A(_04601_),
    .B(_04753_));
 sg13g2_nand2_1 _35343_ (.Y(_04755_),
    .A(\u_inv.d_next[247] ),
    .B(_18367_));
 sg13g2_nand2_1 _35344_ (.Y(_04756_),
    .A(\u_inv.d_next[246] ),
    .B(_18368_));
 sg13g2_nand2_1 _35345_ (.Y(_04757_),
    .A(\u_inv.d_next[244] ),
    .B(_18370_));
 sg13g2_nor2_1 _35346_ (.A(_03593_),
    .B(_04757_),
    .Y(_04758_));
 sg13g2_a21oi_1 _35347_ (.A1(net7295),
    .A2(_18369_),
    .Y(_04759_),
    .B1(_04758_));
 sg13g2_o21ai_1 _35348_ (.B1(_04756_),
    .Y(_04760_),
    .A1(_03601_),
    .A2(_04759_));
 sg13g2_nand2b_1 _35349_ (.Y(_04761_),
    .B(_04760_),
    .A_N(_03603_));
 sg13g2_nand3_1 _35350_ (.B(_04755_),
    .C(_04761_),
    .A(_04754_),
    .Y(_04762_));
 sg13g2_nand2_1 _35351_ (.Y(_04763_),
    .A(\u_inv.d_next[248] ),
    .B(_18366_));
 sg13g2_nand2_1 _35352_ (.Y(_04764_),
    .A(\u_inv.d_next[249] ),
    .B(_18365_));
 sg13g2_o21ai_1 _35353_ (.B1(_04764_),
    .Y(_04765_),
    .A1(_03583_),
    .A2(_04763_));
 sg13g2_inv_1 _35354_ (.Y(_04766_),
    .A(_04765_));
 sg13g2_nor2_1 _35355_ (.A(_18102_),
    .B(\u_inv.d_reg[251] ),
    .Y(_04767_));
 sg13g2_nor2b_1 _35356_ (.A(\u_inv.d_reg[250] ),
    .B_N(\u_inv.d_next[250] ),
    .Y(_04768_));
 sg13g2_a21oi_1 _35357_ (.A1(_03589_),
    .A2(_04768_),
    .Y(_04769_),
    .B1(_04767_));
 sg13g2_o21ai_1 _35358_ (.B1(_04769_),
    .Y(_04770_),
    .A1(_04596_),
    .A2(_04766_));
 sg13g2_nand2_1 _35359_ (.Y(_04771_),
    .A(\u_inv.d_next[254] ),
    .B(_18360_));
 sg13g2_nand2_1 _35360_ (.Y(_04772_),
    .A(\u_inv.d_next[252] ),
    .B(_18362_));
 sg13g2_nor2_1 _35361_ (.A(_03574_),
    .B(_04772_),
    .Y(_04773_));
 sg13g2_a21oi_1 _35362_ (.A1(\u_inv.d_next[253] ),
    .A2(_18361_),
    .Y(_04774_),
    .B1(_04773_));
 sg13g2_o21ai_1 _35363_ (.B1(_04771_),
    .Y(_04775_),
    .A1(_03570_),
    .A2(_04774_));
 sg13g2_nor2b_1 _35364_ (.A(\u_inv.d_reg[255] ),
    .B_N(\u_inv.d_next[255] ),
    .Y(_04776_));
 sg13g2_a21o_1 _35365_ (.A2(_04775_),
    .A1(_03567_),
    .B1(_04776_),
    .X(_04777_));
 sg13g2_a221oi_1 _35366_ (.B2(_04595_),
    .C1(_04777_),
    .B1(_04770_),
    .A1(_04599_),
    .Y(_04778_),
    .A2(_04762_));
 sg13g2_nand2b_1 _35367_ (.Y(_04779_),
    .B(_04105_),
    .A_N(_04107_));
 sg13g2_nand2_1 _35368_ (.Y(_04780_),
    .A(_04101_),
    .B(_04103_));
 sg13g2_nor2_1 _35369_ (.A(_04779_),
    .B(_04780_),
    .Y(_04781_));
 sg13g2_and2_1 _35370_ (.A(_04111_),
    .B(_04113_),
    .X(_04782_));
 sg13g2_nand2_1 _35371_ (.Y(_04783_),
    .A(\u_inv.d_next[56] ),
    .B(_18558_));
 sg13g2_o21ai_1 _35372_ (.B1(_04118_),
    .Y(_04784_),
    .A1(_04117_),
    .A2(_04783_));
 sg13g2_nand2_1 _35373_ (.Y(_04785_),
    .A(\u_inv.d_next[58] ),
    .B(_18556_));
 sg13g2_a22oi_1 _35374_ (.Y(_04786_),
    .B1(_04782_),
    .B2(_04784_),
    .A2(_18555_),
    .A1(\u_inv.d_next[59] ));
 sg13g2_o21ai_1 _35375_ (.B1(_04786_),
    .Y(_04787_),
    .A1(_04110_),
    .A2(_04785_));
 sg13g2_nor2b_1 _35376_ (.A(\u_inv.d_reg[62] ),
    .B_N(\u_inv.d_next[62] ),
    .Y(_04788_));
 sg13g2_nand2_1 _35377_ (.Y(_04789_),
    .A(_04101_),
    .B(_04788_));
 sg13g2_nand2_1 _35378_ (.Y(_04790_),
    .A(\u_inv.d_next[60] ),
    .B(_18554_));
 sg13g2_o21ai_1 _35379_ (.B1(_04790_),
    .Y(_04791_),
    .A1(_18161_),
    .A2(\u_inv.d_reg[61] ));
 sg13g2_o21ai_1 _35380_ (.B1(_04791_),
    .Y(_04792_),
    .A1(\u_inv.d_next[61] ),
    .A2(_18553_));
 sg13g2_o21ai_1 _35381_ (.B1(_04789_),
    .Y(_04793_),
    .A1(_04780_),
    .A2(_04792_));
 sg13g2_a221oi_1 _35382_ (.B2(_04787_),
    .C1(_04793_),
    .B1(_04781_),
    .A1(\u_inv.d_next[63] ),
    .Y(_04794_),
    .A2(_18551_));
 sg13g2_nor2_1 _35383_ (.A(_04120_),
    .B(_04122_),
    .Y(_04795_));
 sg13g2_inv_1 _35384_ (.Y(_04796_),
    .A(_04795_));
 sg13g2_nand3_1 _35385_ (.B(_04782_),
    .C(_04795_),
    .A(_04781_),
    .Y(_04797_));
 sg13g2_nand2_1 _35386_ (.Y(_04798_),
    .A(\u_inv.d_next[48] ),
    .B(_18566_));
 sg13g2_o21ai_1 _35387_ (.B1(_04798_),
    .Y(_04799_),
    .A1(_18164_),
    .A2(\u_inv.d_reg[49] ));
 sg13g2_o21ai_1 _35388_ (.B1(_04799_),
    .Y(_04800_),
    .A1(\u_inv.d_next[49] ),
    .A2(_18565_));
 sg13g2_nand4_1 _35389_ (.B(_04132_),
    .C(_04134_),
    .A(_04128_),
    .Y(_04801_),
    .D(_04137_));
 sg13g2_nor2_1 _35390_ (.A(_04142_),
    .B(_04144_),
    .Y(_04802_));
 sg13g2_inv_1 _35391_ (.Y(_04803_),
    .A(_04802_));
 sg13g2_nor2b_1 _35392_ (.A(\u_inv.d_reg[50] ),
    .B_N(net7298),
    .Y(_04804_));
 sg13g2_a21oi_1 _35393_ (.A1(\u_inv.d_next[51] ),
    .A2(_18563_),
    .Y(_04805_),
    .B1(_04804_));
 sg13g2_or2_1 _35394_ (.X(_04806_),
    .B(_04805_),
    .A(_04140_));
 sg13g2_nand2_2 _35395_ (.Y(_04807_),
    .A(\u_inv.d_next[54] ),
    .B(_18560_));
 sg13g2_a21oi_1 _35396_ (.A1(_18162_),
    .A2(\u_inv.d_reg[55] ),
    .Y(_04808_),
    .B1(_04807_));
 sg13g2_nand2_1 _35397_ (.Y(_04809_),
    .A(\u_inv.d_next[52] ),
    .B(_18562_));
 sg13g2_nor2b_1 _35398_ (.A(_04809_),
    .B_N(_04132_),
    .Y(_04810_));
 sg13g2_a21o_1 _35399_ (.A2(_18561_),
    .A1(\u_inv.d_next[53] ),
    .B1(_04810_),
    .X(_04811_));
 sg13g2_and3_1 _35400_ (.X(_04812_),
    .A(_04134_),
    .B(_04137_),
    .C(_04811_));
 sg13g2_o21ai_1 _35401_ (.B1(_04806_),
    .Y(_04813_),
    .A1(_04800_),
    .A2(_04803_));
 sg13g2_nor2b_1 _35402_ (.A(_04801_),
    .B_N(_04813_),
    .Y(_04814_));
 sg13g2_nor4_2 _35403_ (.A(_04133_),
    .B(_04808_),
    .C(_04812_),
    .Y(_04815_),
    .D(_04814_));
 sg13g2_nor2_1 _35404_ (.A(_04146_),
    .B(_04149_),
    .Y(_04816_));
 sg13g2_nand3b_1 _35405_ (.B(_04802_),
    .C(_04816_),
    .Y(_04817_),
    .A_N(_04801_));
 sg13g2_inv_1 _35406_ (.Y(_04818_),
    .A(_04817_));
 sg13g2_or2_1 _35407_ (.X(_04819_),
    .B(_04199_),
    .A(_04197_));
 sg13g2_nand2_1 _35408_ (.Y(_04820_),
    .A(_04185_),
    .B(_04189_));
 sg13g2_nor3_1 _35409_ (.A(_04179_),
    .B(_04183_),
    .C(_04820_),
    .Y(_04821_));
 sg13g2_nor2b_1 _35410_ (.A(_04193_),
    .B_N(_04191_),
    .Y(_04822_));
 sg13g2_nand2_1 _35411_ (.Y(_04823_),
    .A(_04821_),
    .B(_04822_));
 sg13g2_nor2_1 _35412_ (.A(_04819_),
    .B(_04823_),
    .Y(_04824_));
 sg13g2_nand2_1 _35413_ (.Y(_04825_),
    .A(_04342_),
    .B(_04345_));
 sg13g2_inv_1 _35414_ (.Y(_04826_),
    .A(_04825_));
 sg13g2_nor3_1 _35415_ (.A(_04350_),
    .B(_04352_),
    .C(_04825_),
    .Y(_04827_));
 sg13g2_and2_1 _35416_ (.A(_04357_),
    .B(_04358_),
    .X(_04828_));
 sg13g2_nor2b_1 _35417_ (.A(\u_inv.d_reg[32] ),
    .B_N(\u_inv.d_next[32] ),
    .Y(_04829_));
 sg13g2_o21ai_1 _35418_ (.B1(_04829_),
    .Y(_04830_),
    .A1(\u_inv.d_next[33] ),
    .A2(_18581_));
 sg13g2_o21ai_1 _35419_ (.B1(_04830_),
    .Y(_04831_),
    .A1(_18173_),
    .A2(\u_inv.d_reg[33] ));
 sg13g2_nor2b_1 _35420_ (.A(\u_inv.d_reg[34] ),
    .B_N(\u_inv.d_next[34] ),
    .Y(_04832_));
 sg13g2_o21ai_1 _35421_ (.B1(_04355_),
    .Y(_04833_),
    .A1(_04356_),
    .A2(_04832_));
 sg13g2_inv_1 _35422_ (.Y(_04834_),
    .A(_04833_));
 sg13g2_a21oi_1 _35423_ (.A1(_04828_),
    .A2(_04831_),
    .Y(_04835_),
    .B1(_04834_));
 sg13g2_nand2b_1 _35424_ (.Y(_04836_),
    .B(_04827_),
    .A_N(_04835_));
 sg13g2_nand2_1 _35425_ (.Y(_04837_),
    .A(\u_inv.d_next[38] ),
    .B(_18576_));
 sg13g2_o21ai_1 _35426_ (.B1(_04348_),
    .Y(_04838_),
    .A1(_04347_),
    .A2(_04837_));
 sg13g2_nor2_1 _35427_ (.A(_18171_),
    .B(\u_inv.d_reg[36] ),
    .Y(_04839_));
 sg13g2_nor2b_1 _35428_ (.A(\u_inv.d_reg[37] ),
    .B_N(\u_inv.d_next[37] ),
    .Y(_04840_));
 sg13g2_a21o_1 _35429_ (.A2(_04839_),
    .A1(_04342_),
    .B1(_04840_),
    .X(_04841_));
 sg13g2_nand3_1 _35430_ (.B(_04353_),
    .C(_04841_),
    .A(_04349_),
    .Y(_04842_));
 sg13g2_nand3b_1 _35431_ (.B(_04842_),
    .C(_04836_),
    .Y(_04843_),
    .A_N(_04838_));
 sg13g2_inv_1 _35432_ (.Y(_04844_),
    .A(_04843_));
 sg13g2_nand2_1 _35433_ (.Y(_04845_),
    .A(\u_inv.d_next[40] ),
    .B(_18574_));
 sg13g2_nor2_1 _35434_ (.A(_04197_),
    .B(_04845_),
    .Y(_04846_));
 sg13g2_a21oi_1 _35435_ (.A1(\u_inv.d_next[41] ),
    .A2(_18573_),
    .Y(_04847_),
    .B1(_04846_));
 sg13g2_inv_1 _35436_ (.Y(_04848_),
    .A(_04847_));
 sg13g2_nand2_1 _35437_ (.Y(_04849_),
    .A(\u_inv.d_next[44] ),
    .B(_18570_));
 sg13g2_nand2_1 _35438_ (.Y(_04850_),
    .A(\u_inv.d_next[45] ),
    .B(_18569_));
 sg13g2_o21ai_1 _35439_ (.B1(_04850_),
    .Y(_04851_),
    .A1(_04183_),
    .A2(_04849_));
 sg13g2_inv_1 _35440_ (.Y(_04852_),
    .A(_04851_));
 sg13g2_nand2_1 _35441_ (.Y(_04853_),
    .A(\u_inv.d_next[46] ),
    .B(_18568_));
 sg13g2_a21oi_1 _35442_ (.A1(_18165_),
    .A2(\u_inv.d_reg[47] ),
    .Y(_04854_),
    .B1(_04853_));
 sg13g2_nor2_1 _35443_ (.A(_18169_),
    .B(\u_inv.d_reg[42] ),
    .Y(_04855_));
 sg13g2_a21oi_1 _35444_ (.A1(\u_inv.d_next[43] ),
    .A2(_18571_),
    .Y(_04856_),
    .B1(_04855_));
 sg13g2_a21oi_1 _35445_ (.A1(_18168_),
    .A2(\u_inv.d_reg[43] ),
    .Y(_04857_),
    .B1(_04856_));
 sg13g2_inv_1 _35446_ (.Y(_04858_),
    .A(_04857_));
 sg13g2_a221oi_1 _35447_ (.B2(_04857_),
    .C1(_04854_),
    .B1(_04821_),
    .A1(\u_inv.d_next[47] ),
    .Y(_04859_),
    .A2(_18567_));
 sg13g2_o21ai_1 _35448_ (.B1(_04859_),
    .Y(_04860_),
    .A1(_04820_),
    .A2(_04852_));
 sg13g2_a21oi_1 _35449_ (.A1(_04824_),
    .A2(_04843_),
    .Y(_04861_),
    .B1(_04860_));
 sg13g2_o21ai_1 _35450_ (.B1(_04861_),
    .Y(_04862_),
    .A1(_04823_),
    .A2(_04847_));
 sg13g2_and2_1 _35451_ (.A(_04206_),
    .B(_04208_),
    .X(_04863_));
 sg13g2_nand2_1 _35452_ (.Y(_04864_),
    .A(_04203_),
    .B(_04204_));
 sg13g2_and3_1 _35453_ (.X(_04865_),
    .A(_04203_),
    .B(_04204_),
    .C(_04863_));
 sg13g2_and2_1 _35454_ (.A(_04212_),
    .B(_04214_),
    .X(_04866_));
 sg13g2_and2_1 _35455_ (.A(_04217_),
    .B(_04218_),
    .X(_04867_));
 sg13g2_inv_1 _35456_ (.Y(_04868_),
    .A(_04867_));
 sg13g2_and3_1 _35457_ (.X(_04869_),
    .A(_04865_),
    .B(_04866_),
    .C(_04867_));
 sg13g2_nor2_1 _35458_ (.A(_18176_),
    .B(\u_inv.d_reg[28] ),
    .Y(_04870_));
 sg13g2_nand2_1 _35459_ (.Y(_04871_),
    .A(_04203_),
    .B(_04870_));
 sg13g2_o21ai_1 _35460_ (.B1(_04871_),
    .Y(_04872_),
    .A1(_18175_),
    .A2(\u_inv.d_reg[29] ));
 sg13g2_nand2_1 _35461_ (.Y(_04873_),
    .A(\u_inv.d_next[30] ),
    .B(_18584_));
 sg13g2_a21oi_1 _35462_ (.A1(_18174_),
    .A2(\u_inv.d_reg[31] ),
    .Y(_04874_),
    .B1(_04873_));
 sg13g2_a221oi_1 _35463_ (.B2(_04872_),
    .C1(_04874_),
    .B1(_04863_),
    .A1(\u_inv.d_next[31] ),
    .Y(_04875_),
    .A2(_18583_));
 sg13g2_nor2b_1 _35464_ (.A(\u_inv.d_reg[24] ),
    .B_N(\u_inv.d_next[24] ),
    .Y(_04876_));
 sg13g2_nor2b_1 _35465_ (.A(\u_inv.d_reg[25] ),
    .B_N(\u_inv.d_next[25] ),
    .Y(_04877_));
 sg13g2_a21o_1 _35466_ (.A2(_04876_),
    .A1(_04217_),
    .B1(_04877_),
    .X(_04878_));
 sg13g2_nand2_1 _35467_ (.Y(_04879_),
    .A(\u_inv.d_next[26] ),
    .B(_18588_));
 sg13g2_and2_1 _35468_ (.A(_04211_),
    .B(_04879_),
    .X(_04880_));
 sg13g2_nand2_1 _35469_ (.Y(_04881_),
    .A(_04211_),
    .B(_04879_));
 sg13g2_a22oi_1 _35470_ (.Y(_04882_),
    .B1(_04881_),
    .B2(_04210_),
    .A2(_04878_),
    .A1(_04866_));
 sg13g2_nand2b_1 _35471_ (.Y(_04883_),
    .B(_04865_),
    .A_N(_04882_));
 sg13g2_nor2_1 _35472_ (.A(_04237_),
    .B(_04239_),
    .Y(_04884_));
 sg13g2_nand3_1 _35473_ (.B(_04248_),
    .C(_04884_),
    .A(_04245_),
    .Y(_04885_));
 sg13g2_nand2_1 _35474_ (.Y(_04886_),
    .A(_04253_),
    .B(_04260_));
 sg13g2_nor2_1 _35475_ (.A(_04885_),
    .B(_04886_),
    .Y(_04887_));
 sg13g2_nand2_1 _35476_ (.Y(_04888_),
    .A(\u_inv.d_next[12] ),
    .B(_18602_));
 sg13g2_nor2_1 _35477_ (.A(_04237_),
    .B(_04888_),
    .Y(_04889_));
 sg13g2_nand2_1 _35478_ (.Y(_04890_),
    .A(\u_inv.d_next[13] ),
    .B(_18601_));
 sg13g2_o21ai_1 _35479_ (.B1(_04890_),
    .Y(_04891_),
    .A1(_04237_),
    .A2(_04888_));
 sg13g2_nand3_1 _35480_ (.B(_04248_),
    .C(_04891_),
    .A(_04245_),
    .Y(_04892_));
 sg13g2_nand3_1 _35481_ (.B(_18600_),
    .C(_04246_),
    .A(\u_inv.d_next[14] ),
    .Y(_04893_));
 sg13g2_nor2b_1 _35482_ (.A(net7292),
    .B_N(\u_inv.d_next[10] ),
    .Y(_04894_));
 sg13g2_o21ai_1 _35483_ (.B1(_04252_),
    .Y(_04895_),
    .A1(_04251_),
    .A2(_04894_));
 sg13g2_nor2_1 _35484_ (.A(_04885_),
    .B(_04895_),
    .Y(_04896_));
 sg13g2_nor2b_1 _35485_ (.A(\u_inv.d_reg[6] ),
    .B_N(\u_inv.d_next[6] ),
    .Y(_04897_));
 sg13g2_a21oi_1 _35486_ (.A1(\u_inv.d_next[7] ),
    .A2(_18607_),
    .Y(_04898_),
    .B1(_04897_));
 sg13g2_nor2b_1 _35487_ (.A(\u_inv.d_reg[4] ),
    .B_N(\u_inv.d_next[4] ),
    .Y(_04899_));
 sg13g2_nor2b_1 _35488_ (.A(\u_inv.d_reg[3] ),
    .B_N(\u_inv.d_next[3] ),
    .Y(_04900_));
 sg13g2_xnor2_1 _35489_ (.Y(_04901_),
    .A(\u_inv.d_next[3] ),
    .B(\u_inv.d_reg[3] ));
 sg13g2_nand2_1 _35490_ (.Y(_04902_),
    .A(\u_inv.d_next[2] ),
    .B(_18612_));
 sg13g2_o21ai_1 _35491_ (.B1(_04902_),
    .Y(_04903_),
    .A1(_03338_),
    .A2(_03343_));
 sg13g2_a21oi_1 _35492_ (.A1(_04901_),
    .A2(_04903_),
    .Y(_04904_),
    .B1(_04900_));
 sg13g2_nor2_1 _35493_ (.A(_04274_),
    .B(_04904_),
    .Y(_04905_));
 sg13g2_nor2_1 _35494_ (.A(_04899_),
    .B(_04905_),
    .Y(_04906_));
 sg13g2_a21oi_1 _35495_ (.A1(_04267_),
    .A2(_04899_),
    .Y(_04907_),
    .B1(_04268_));
 sg13g2_nand3b_1 _35496_ (.B(_04269_),
    .C(_04275_),
    .Y(_04908_),
    .A_N(_04904_));
 sg13g2_a21o_1 _35497_ (.A2(_04908_),
    .A1(_04907_),
    .B1(_04281_),
    .X(_04909_));
 sg13g2_nand2_1 _35498_ (.Y(_04910_),
    .A(_04281_),
    .B(_04898_));
 sg13g2_nand3_1 _35499_ (.B(_04907_),
    .C(_04908_),
    .A(_04898_),
    .Y(_04911_));
 sg13g2_and3_2 _35500_ (.X(_04912_),
    .A(_04278_),
    .B(_04910_),
    .C(_04911_));
 sg13g2_and2_1 _35501_ (.A(_04255_),
    .B(_04290_),
    .X(_04913_));
 sg13g2_nor2b_1 _35502_ (.A(\u_inv.d_reg[8] ),
    .B_N(\u_inv.d_next[8] ),
    .Y(_04914_));
 sg13g2_a21oi_1 _35503_ (.A1(\u_inv.d_next[9] ),
    .A2(_18605_),
    .Y(_04915_),
    .B1(_04914_));
 sg13g2_a21oi_1 _35504_ (.A1(_18180_),
    .A2(\u_inv.d_reg[9] ),
    .Y(_04916_),
    .B1(_04915_));
 sg13g2_and2_1 _35505_ (.A(_04887_),
    .B(_04913_),
    .X(_04917_));
 sg13g2_and4_1 _35506_ (.A(_04278_),
    .B(_04910_),
    .C(_04911_),
    .D(_04917_),
    .X(_04918_));
 sg13g2_nand4_1 _35507_ (.B(_04910_),
    .C(_04911_),
    .A(_04278_),
    .Y(_04919_),
    .D(_04917_));
 sg13g2_a21oi_1 _35508_ (.A1(_04887_),
    .A2(_04916_),
    .Y(_04920_),
    .B1(_04896_));
 sg13g2_nand4_1 _35509_ (.B(_04892_),
    .C(_04893_),
    .A(_04247_),
    .Y(_04921_),
    .D(_04920_));
 sg13g2_inv_1 _35510_ (.Y(_04922_),
    .A(_04921_));
 sg13g2_nor2_1 _35511_ (.A(_04918_),
    .B(_04921_),
    .Y(_04923_));
 sg13g2_nor2_1 _35512_ (.A(_04306_),
    .B(_04308_),
    .Y(_04924_));
 sg13g2_nor3_1 _35513_ (.A(_04301_),
    .B(_04306_),
    .C(_04308_),
    .Y(_04925_));
 sg13g2_and2_1 _35514_ (.A(_04299_),
    .B(_04925_),
    .X(_04926_));
 sg13g2_nand2_1 _35515_ (.Y(_04927_),
    .A(_04311_),
    .B(_04318_));
 sg13g2_nor2_1 _35516_ (.A(_04315_),
    .B(_04321_),
    .Y(_04928_));
 sg13g2_and4_1 _35517_ (.A(_04311_),
    .B(_04318_),
    .C(_04926_),
    .D(_04928_),
    .X(_04929_));
 sg13g2_o21ai_1 _35518_ (.B1(_04929_),
    .Y(_04930_),
    .A1(_04918_),
    .A2(_04921_));
 sg13g2_nor2b_1 _35519_ (.A(\u_inv.d_reg[16] ),
    .B_N(\u_inv.d_next[16] ),
    .Y(_04931_));
 sg13g2_a21oi_2 _35520_ (.B1(_04313_),
    .Y(_04932_),
    .A2(_04931_),
    .A1(_04312_));
 sg13g2_a22oi_1 _35521_ (.Y(_04933_),
    .B1(_18596_),
    .B2(net7299),
    .A2(_18595_),
    .A1(\u_inv.d_next[19] ));
 sg13g2_a21oi_1 _35522_ (.A1(_18178_),
    .A2(\u_inv.d_reg[19] ),
    .Y(_04934_),
    .B1(_04933_));
 sg13g2_nand2_1 _35523_ (.Y(_04935_),
    .A(\u_inv.d_next[22] ),
    .B(_18592_));
 sg13g2_o21ai_1 _35524_ (.B1(_04304_),
    .Y(_04936_),
    .A1(_04303_),
    .A2(_04935_));
 sg13g2_nand2_1 _35525_ (.Y(_04937_),
    .A(\u_inv.d_next[20] ),
    .B(_18594_));
 sg13g2_nor2_1 _35526_ (.A(_04301_),
    .B(_04937_),
    .Y(_04938_));
 sg13g2_nor2b_1 _35527_ (.A(\u_inv.d_reg[21] ),
    .B_N(\u_inv.d_next[21] ),
    .Y(_04939_));
 sg13g2_o21ai_1 _35528_ (.B1(_04924_),
    .Y(_04940_),
    .A1(_04938_),
    .A2(_04939_));
 sg13g2_nor2_1 _35529_ (.A(_04927_),
    .B(_04932_),
    .Y(_04941_));
 sg13g2_o21ai_1 _35530_ (.B1(_04926_),
    .Y(_04942_),
    .A1(_04934_),
    .A2(_04941_));
 sg13g2_nand3b_1 _35531_ (.B(_04940_),
    .C(_04942_),
    .Y(_04943_),
    .A_N(_04936_));
 sg13g2_inv_1 _35532_ (.Y(_04944_),
    .A(_04943_));
 sg13g2_nand2_1 _35533_ (.Y(_04945_),
    .A(_04869_),
    .B(_04943_));
 sg13g2_and3_2 _35534_ (.X(_04946_),
    .A(_04875_),
    .B(_04883_),
    .C(_04945_));
 sg13g2_inv_1 _35535_ (.Y(_04947_),
    .A(_04946_));
 sg13g2_nand2_1 _35536_ (.Y(_04948_),
    .A(_04869_),
    .B(_04929_));
 sg13g2_a21oi_2 _35537_ (.B1(_04948_),
    .Y(_04949_),
    .A2(_04922_),
    .A1(_04919_));
 sg13g2_a21o_2 _35538_ (.A2(_04922_),
    .A1(_04919_),
    .B1(_04948_),
    .X(_04950_));
 sg13g2_nand2_1 _35539_ (.Y(_04951_),
    .A(_04946_),
    .B(_04950_));
 sg13g2_and4_1 _35540_ (.A(net6995),
    .B(_04365_),
    .C(_04827_),
    .D(_04828_),
    .X(_04952_));
 sg13g2_and2_1 _35541_ (.A(_04824_),
    .B(_04952_),
    .X(_04953_));
 sg13g2_inv_1 _35542_ (.Y(_04954_),
    .A(_04953_));
 sg13g2_a21oi_1 _35543_ (.A1(_04946_),
    .A2(_04950_),
    .Y(_04955_),
    .B1(_04954_));
 sg13g2_nor2_1 _35544_ (.A(_04862_),
    .B(_04955_),
    .Y(_04956_));
 sg13g2_o21ai_1 _35545_ (.B1(_04818_),
    .Y(_04957_),
    .A1(_04862_),
    .A2(_04955_));
 sg13g2_nand2_1 _35546_ (.Y(_04958_),
    .A(_04815_),
    .B(_04957_));
 sg13g2_o21ai_1 _35547_ (.B1(_04794_),
    .Y(_04959_),
    .A1(_04797_),
    .A2(_04815_));
 sg13g2_nor2_1 _35548_ (.A(_04797_),
    .B(_04817_),
    .Y(_04960_));
 sg13g2_nand2_1 _35549_ (.Y(_04961_),
    .A(_04953_),
    .B(_04960_));
 sg13g2_a21oi_2 _35550_ (.B1(_04961_),
    .Y(_04962_),
    .A2(_04950_),
    .A1(_04946_));
 sg13g2_and2_1 _35551_ (.A(_04862_),
    .B(_04960_),
    .X(_04963_));
 sg13g2_nor3_2 _35552_ (.A(_04959_),
    .B(_04962_),
    .C(_04963_),
    .Y(_04964_));
 sg13g2_or3_1 _35553_ (.A(_04959_),
    .B(_04962_),
    .C(_04963_),
    .X(_04965_));
 sg13g2_nor2_1 _35554_ (.A(_03810_),
    .B(_03813_),
    .Y(_04966_));
 sg13g2_nor2_1 _35555_ (.A(_03814_),
    .B(_03817_),
    .Y(_04967_));
 sg13g2_or2_1 _35556_ (.X(_04968_),
    .B(_03817_),
    .A(_03814_));
 sg13g2_nand2_1 _35557_ (.Y(_04969_),
    .A(_04966_),
    .B(_04967_));
 sg13g2_nor2_1 _35558_ (.A(_03820_),
    .B(_03823_),
    .Y(_04970_));
 sg13g2_and2_1 _35559_ (.A(_03827_),
    .B(_03874_),
    .X(_04971_));
 sg13g2_and4_1 _35560_ (.A(_04966_),
    .B(_04967_),
    .C(_04970_),
    .D(_04971_),
    .X(_04972_));
 sg13g2_nor2_1 _35561_ (.A(_03850_),
    .B(_03852_),
    .Y(_04973_));
 sg13g2_inv_1 _35562_ (.Y(_04974_),
    .A(_04973_));
 sg13g2_nor2_1 _35563_ (.A(_03842_),
    .B(_03845_),
    .Y(_04975_));
 sg13g2_nand2_1 _35564_ (.Y(_04976_),
    .A(_04973_),
    .B(_04975_));
 sg13g2_and2_1 _35565_ (.A(_03855_),
    .B(_03864_),
    .X(_04977_));
 sg13g2_nand2_1 _35566_ (.Y(_04978_),
    .A(_03855_),
    .B(_03864_));
 sg13g2_nor4_1 _35567_ (.A(_03859_),
    .B(_03951_),
    .C(_04976_),
    .D(_04978_),
    .Y(_04979_));
 sg13g2_nand2_1 _35568_ (.Y(_04980_),
    .A(_04972_),
    .B(_04979_));
 sg13g2_inv_1 _35569_ (.Y(_04981_),
    .A(_04980_));
 sg13g2_nor2_1 _35570_ (.A(_03877_),
    .B(_03880_),
    .Y(_04982_));
 sg13g2_nor2_1 _35571_ (.A(_03883_),
    .B(_03888_),
    .Y(_04983_));
 sg13g2_and2_1 _35572_ (.A(_04982_),
    .B(_04983_),
    .X(_04984_));
 sg13g2_nor2_2 _35573_ (.A(_03892_),
    .B(_03894_),
    .Y(_04985_));
 sg13g2_nor2_1 _35574_ (.A(_03896_),
    .B(_03898_),
    .Y(_04986_));
 sg13g2_nand2b_1 _35575_ (.Y(_04987_),
    .B(_03899_),
    .A_N(_03896_));
 sg13g2_nand3_1 _35576_ (.B(_04985_),
    .C(_04986_),
    .A(_04984_),
    .Y(_04988_));
 sg13g2_and2_1 _35577_ (.A(_03911_),
    .B(_03913_),
    .X(_04989_));
 sg13g2_nand3_1 _35578_ (.B(_03908_),
    .C(_04989_),
    .A(_03904_),
    .Y(_04990_));
 sg13g2_nand2_1 _35579_ (.Y(_04991_),
    .A(_03917_),
    .B(_03929_));
 sg13g2_or2_1 _35580_ (.X(_04992_),
    .B(_04991_),
    .A(_04990_));
 sg13g2_and2_1 _35581_ (.A(_03923_),
    .B(_04409_),
    .X(_04993_));
 sg13g2_nand2b_1 _35582_ (.Y(_04994_),
    .B(_04993_),
    .A_N(_04992_));
 sg13g2_nor2_2 _35583_ (.A(_04988_),
    .B(_04994_),
    .Y(_04995_));
 sg13g2_nand2_1 _35584_ (.Y(_04996_),
    .A(_04981_),
    .B(_04995_));
 sg13g2_nand2_1 _35585_ (.Y(_04997_),
    .A(_03997_),
    .B(_03999_));
 sg13g2_nand2_1 _35586_ (.Y(_04998_),
    .A(_03991_),
    .B(_03993_));
 sg13g2_inv_1 _35587_ (.Y(_04999_),
    .A(_04998_));
 sg13g2_nor2_1 _35588_ (.A(_04997_),
    .B(_04998_),
    .Y(_05000_));
 sg13g2_nand2_1 _35589_ (.Y(_05001_),
    .A(_03981_),
    .B(_03986_));
 sg13g2_nand2_1 _35590_ (.Y(_05002_),
    .A(_03982_),
    .B(_03988_));
 sg13g2_nor4_1 _35591_ (.A(_04997_),
    .B(_04998_),
    .C(_05001_),
    .D(_05002_),
    .Y(_05003_));
 sg13g2_nor2_1 _35592_ (.A(_03958_),
    .B(_03959_),
    .Y(_05004_));
 sg13g2_nor2_1 _35593_ (.A(_03962_),
    .B(_03964_),
    .Y(_05005_));
 sg13g2_nand2_1 _35594_ (.Y(_05006_),
    .A(_05004_),
    .B(_05005_));
 sg13g2_nand2_1 _35595_ (.Y(_05007_),
    .A(_03968_),
    .B(_03973_));
 sg13g2_nand2b_1 _35596_ (.Y(_05008_),
    .B(_03975_),
    .A_N(_03978_));
 sg13g2_or2_1 _35597_ (.X(_05009_),
    .B(_05008_),
    .A(_05007_));
 sg13g2_nor2_1 _35598_ (.A(_05006_),
    .B(_05009_),
    .Y(_05010_));
 sg13g2_nand2_1 _35599_ (.Y(_05011_),
    .A(_05003_),
    .B(_05010_));
 sg13g2_inv_1 _35600_ (.Y(_05012_),
    .A(_05011_));
 sg13g2_nor2_1 _35601_ (.A(_04013_),
    .B(_04018_),
    .Y(_05013_));
 sg13g2_nor4_1 _35602_ (.A(_04006_),
    .B(_04009_),
    .C(_04013_),
    .D(_04018_),
    .Y(_05014_));
 sg13g2_and2_1 _35603_ (.A(_04029_),
    .B(_04031_),
    .X(_05015_));
 sg13g2_nand2_1 _35604_ (.Y(_05016_),
    .A(_05014_),
    .B(_05015_));
 sg13g2_nand2_1 _35605_ (.Y(_05017_),
    .A(_04044_),
    .B(_04047_));
 sg13g2_nand2_1 _35606_ (.Y(_05018_),
    .A(_04039_),
    .B(_04041_));
 sg13g2_inv_1 _35607_ (.Y(_05019_),
    .A(_05018_));
 sg13g2_nand2b_1 _35608_ (.Y(_05020_),
    .B(_05019_),
    .A_N(_05017_));
 sg13g2_inv_1 _35609_ (.Y(_05021_),
    .A(_05020_));
 sg13g2_nand2_1 _35610_ (.Y(_05022_),
    .A(_04056_),
    .B(_04059_));
 sg13g2_inv_1 _35611_ (.Y(_05023_),
    .A(_05022_));
 sg13g2_nand2_1 _35612_ (.Y(_05024_),
    .A(_04049_),
    .B(_04053_));
 sg13g2_nor3_1 _35613_ (.A(_05020_),
    .B(_05022_),
    .C(_05024_),
    .Y(_05025_));
 sg13g2_or2_1 _35614_ (.X(_05026_),
    .B(_04401_),
    .A(_04024_));
 sg13g2_nor2_1 _35615_ (.A(_05016_),
    .B(_05026_),
    .Y(_05027_));
 sg13g2_nand2_1 _35616_ (.Y(_05028_),
    .A(_05025_),
    .B(_05027_));
 sg13g2_inv_2 _35617_ (.Y(_05029_),
    .A(_05028_));
 sg13g2_nand2_2 _35618_ (.Y(_05030_),
    .A(_05012_),
    .B(_05029_));
 sg13g2_nor2_1 _35619_ (.A(_04996_),
    .B(_05030_),
    .Y(_05031_));
 sg13g2_nor2b_1 _35620_ (.A(\u_inv.d_reg[64] ),
    .B_N(\u_inv.d_next[64] ),
    .Y(_05032_));
 sg13g2_a21oi_1 _35621_ (.A1(_04022_),
    .A2(_05032_),
    .Y(_05033_),
    .B1(_04023_));
 sg13g2_nor2_1 _35622_ (.A(_18159_),
    .B(\u_inv.d_reg[66] ),
    .Y(_05034_));
 sg13g2_o21ai_1 _35623_ (.B1(_05034_),
    .Y(_05035_),
    .A1(\u_inv.d_next[67] ),
    .A2(_18547_));
 sg13g2_o21ai_1 _35624_ (.B1(_05035_),
    .Y(_05036_),
    .A1(_18158_),
    .A2(\u_inv.d_reg[67] ));
 sg13g2_nand2_1 _35625_ (.Y(_05037_),
    .A(net7297),
    .B(_18544_));
 sg13g2_o21ai_1 _35626_ (.B1(_04016_),
    .Y(_05038_),
    .A1(_04015_),
    .A2(_05037_));
 sg13g2_nand2_1 _35627_ (.Y(_05039_),
    .A(\u_inv.d_next[68] ),
    .B(_18546_));
 sg13g2_nand2_1 _35628_ (.Y(_05040_),
    .A(\u_inv.d_next[69] ),
    .B(_18545_));
 sg13g2_o21ai_1 _35629_ (.B1(_05040_),
    .Y(_05041_),
    .A1(_04009_),
    .A2(_05039_));
 sg13g2_a221oi_1 _35630_ (.B2(_05013_),
    .C1(_05038_),
    .B1(_05041_),
    .A1(_05014_),
    .Y(_05042_),
    .A2(_05036_));
 sg13g2_o21ai_1 _35631_ (.B1(_05042_),
    .Y(_05043_),
    .A1(_05016_),
    .A2(_05033_));
 sg13g2_nand2_1 _35632_ (.Y(_05044_),
    .A(\u_inv.d_next[76] ),
    .B(_18538_));
 sg13g2_nor2b_1 _35633_ (.A(_05044_),
    .B_N(_04039_),
    .Y(_05045_));
 sg13g2_a21oi_1 _35634_ (.A1(\u_inv.d_next[77] ),
    .A2(_18537_),
    .Y(_05046_),
    .B1(_05045_));
 sg13g2_nand2_1 _35635_ (.Y(_05047_),
    .A(\u_inv.d_next[78] ),
    .B(_18536_));
 sg13g2_o21ai_1 _35636_ (.B1(_04046_),
    .Y(_05048_),
    .A1(_04045_),
    .A2(_05047_));
 sg13g2_nor2_1 _35637_ (.A(_18157_),
    .B(\u_inv.d_reg[72] ),
    .Y(_05049_));
 sg13g2_nor2b_1 _35638_ (.A(\u_inv.d_reg[73] ),
    .B_N(\u_inv.d_next[73] ),
    .Y(_05050_));
 sg13g2_a21oi_2 _35639_ (.B1(_05050_),
    .Y(_05051_),
    .A2(_05049_),
    .A1(_04056_));
 sg13g2_nor2_1 _35640_ (.A(_05024_),
    .B(_05051_),
    .Y(_05052_));
 sg13g2_nor2b_1 _35641_ (.A(\u_inv.d_reg[74] ),
    .B_N(\u_inv.d_next[74] ),
    .Y(_05053_));
 sg13g2_o21ai_1 _35642_ (.B1(_05053_),
    .Y(_05054_),
    .A1(\u_inv.d_next[75] ),
    .A2(_18539_));
 sg13g2_o21ai_1 _35643_ (.B1(_05054_),
    .Y(_05055_),
    .A1(_18156_),
    .A2(\u_inv.d_reg[75] ));
 sg13g2_or2_1 _35644_ (.X(_05056_),
    .B(_05055_),
    .A(_05052_));
 sg13g2_a221oi_1 _35645_ (.B2(_05021_),
    .C1(_05048_),
    .B1(_05056_),
    .A1(_05025_),
    .Y(_05057_),
    .A2(_05043_));
 sg13g2_o21ai_1 _35646_ (.B1(_05057_),
    .Y(_05058_),
    .A1(_05017_),
    .A2(_05046_));
 sg13g2_nand2_1 _35647_ (.Y(_05059_),
    .A(\u_inv.d_next[88] ),
    .B(_18526_));
 sg13g2_o21ai_1 _35648_ (.B1(_05059_),
    .Y(_05060_),
    .A1(_18149_),
    .A2(\u_inv.d_reg[89] ));
 sg13g2_o21ai_1 _35649_ (.B1(_05060_),
    .Y(_05061_),
    .A1(\u_inv.d_next[89] ),
    .A2(_18525_));
 sg13g2_nor2b_1 _35650_ (.A(\u_inv.d_reg[90] ),
    .B_N(\u_inv.d_next[90] ),
    .Y(_05062_));
 sg13g2_o21ai_1 _35651_ (.B1(_03967_),
    .Y(_05063_),
    .A1(_05007_),
    .A2(_05061_));
 sg13g2_a21oi_1 _35652_ (.A1(_03966_),
    .A2(_05062_),
    .Y(_05064_),
    .B1(_05063_));
 sg13g2_nor2b_1 _35653_ (.A(\u_inv.d_reg[92] ),
    .B_N(\u_inv.d_next[92] ),
    .Y(_05065_));
 sg13g2_a21oi_1 _35654_ (.A1(\u_inv.d_next[93] ),
    .A2(_18521_),
    .Y(_05066_),
    .B1(_05065_));
 sg13g2_a21oi_1 _35655_ (.A1(_18148_),
    .A2(\u_inv.d_reg[93] ),
    .Y(_05067_),
    .B1(_05066_));
 sg13g2_nand2_1 _35656_ (.Y(_05068_),
    .A(\u_inv.d_next[94] ),
    .B(_18520_));
 sg13g2_nor2_1 _35657_ (.A(_03959_),
    .B(_05068_),
    .Y(_05069_));
 sg13g2_a221oi_1 _35658_ (.B2(_05067_),
    .C1(_05069_),
    .B1(_05004_),
    .A1(\u_inv.d_next[95] ),
    .Y(_05070_),
    .A2(_18519_));
 sg13g2_o21ai_1 _35659_ (.B1(_05070_),
    .Y(_05071_),
    .A1(_05006_),
    .A2(_05064_));
 sg13g2_nand2_1 _35660_ (.Y(_05072_),
    .A(\u_inv.d_next[80] ),
    .B(_18534_));
 sg13g2_o21ai_1 _35661_ (.B1(_05072_),
    .Y(_05073_),
    .A1(_18152_),
    .A2(net7290));
 sg13g2_o21ai_1 _35662_ (.B1(_05073_),
    .Y(_05074_),
    .A1(\u_inv.d_next[81] ),
    .A2(_18533_));
 sg13g2_nor2_1 _35663_ (.A(_05001_),
    .B(_05074_),
    .Y(_05075_));
 sg13g2_nor2b_1 _35664_ (.A(\u_inv.d_reg[82] ),
    .B_N(\u_inv.d_next[82] ),
    .Y(_05076_));
 sg13g2_o21ai_1 _35665_ (.B1(_05076_),
    .Y(_05077_),
    .A1(\u_inv.d_next[83] ),
    .A2(_18531_));
 sg13g2_o21ai_1 _35666_ (.B1(_05077_),
    .Y(_05078_),
    .A1(_18151_),
    .A2(\u_inv.d_reg[83] ));
 sg13g2_o21ai_1 _35667_ (.B1(_05000_),
    .Y(_05079_),
    .A1(_05075_),
    .A2(_05078_));
 sg13g2_nor2b_1 _35668_ (.A(\u_inv.d_reg[86] ),
    .B_N(\u_inv.d_next[86] ),
    .Y(_05080_));
 sg13g2_o21ai_1 _35669_ (.B1(_05080_),
    .Y(_05081_),
    .A1(\u_inv.d_next[87] ),
    .A2(_18527_));
 sg13g2_nor2b_1 _35670_ (.A(\u_inv.d_reg[84] ),
    .B_N(\u_inv.d_next[84] ),
    .Y(_05082_));
 sg13g2_nand2_1 _35671_ (.Y(_05083_),
    .A(\u_inv.d_next[84] ),
    .B(_18530_));
 sg13g2_nor2_1 _35672_ (.A(_18150_),
    .B(\u_inv.d_reg[85] ),
    .Y(_05084_));
 sg13g2_a21oi_1 _35673_ (.A1(_03991_),
    .A2(_05082_),
    .Y(_05085_),
    .B1(_05084_));
 sg13g2_or2_1 _35674_ (.X(_05086_),
    .B(_05085_),
    .A(_04997_));
 sg13g2_nand4_1 _35675_ (.B(_05079_),
    .C(_05081_),
    .A(_03998_),
    .Y(_05087_),
    .D(_05086_));
 sg13g2_a221oi_1 _35676_ (.B2(_05010_),
    .C1(_05071_),
    .B1(_05087_),
    .A1(_05012_),
    .Y(_05088_),
    .A2(_05058_));
 sg13g2_nand2_1 _35677_ (.Y(_05089_),
    .A(\u_inv.d_next[112] ),
    .B(_18502_));
 sg13g2_a21oi_2 _35678_ (.B1(_03857_),
    .Y(_05090_),
    .A2(_05089_),
    .A1(_03858_));
 sg13g2_nand2_1 _35679_ (.Y(_05091_),
    .A(_04977_),
    .B(_05090_));
 sg13g2_nor2b_1 _35680_ (.A(\u_inv.d_reg[114] ),
    .B_N(\u_inv.d_next[114] ),
    .Y(_05092_));
 sg13g2_a21oi_1 _35681_ (.A1(\u_inv.d_next[115] ),
    .A2(_18499_),
    .Y(_05093_),
    .B1(_05092_));
 sg13g2_a21o_2 _35682_ (.A2(\u_inv.d_reg[115] ),
    .A1(_18140_),
    .B1(_05093_),
    .X(_05094_));
 sg13g2_a21oi_1 _35683_ (.A1(_05091_),
    .A2(_05094_),
    .Y(_05095_),
    .B1(_04976_));
 sg13g2_nand2_1 _35684_ (.Y(_05096_),
    .A(\u_inv.d_next[118] ),
    .B(_18496_));
 sg13g2_nor2_1 _35685_ (.A(_03842_),
    .B(_05096_),
    .Y(_05097_));
 sg13g2_a21oi_1 _35686_ (.A1(\u_inv.d_next[119] ),
    .A2(_18495_),
    .Y(_05098_),
    .B1(_05097_));
 sg13g2_nor2b_1 _35687_ (.A(\u_inv.d_reg[116] ),
    .B_N(\u_inv.d_next[116] ),
    .Y(_05099_));
 sg13g2_nand2_1 _35688_ (.Y(_05100_),
    .A(\u_inv.d_next[116] ),
    .B(_18498_));
 sg13g2_o21ai_1 _35689_ (.B1(_03848_),
    .Y(_05101_),
    .A1(_03847_),
    .A2(_05100_));
 sg13g2_a21oi_1 _35690_ (.A1(_04975_),
    .A2(_05101_),
    .Y(_05102_),
    .B1(_05095_));
 sg13g2_nand2_1 _35691_ (.Y(_05103_),
    .A(_05098_),
    .B(_05102_));
 sg13g2_nor2b_1 _35692_ (.A(\u_inv.d_reg[120] ),
    .B_N(\u_inv.d_next[120] ),
    .Y(_05104_));
 sg13g2_a21o_1 _35693_ (.A2(_05104_),
    .A1(_03825_),
    .B1(_03826_),
    .X(_05105_));
 sg13g2_nand2_1 _35694_ (.Y(_05106_),
    .A(\u_inv.d_next[122] ),
    .B(_18492_));
 sg13g2_nor2_1 _35695_ (.A(_03820_),
    .B(_05106_),
    .Y(_05107_));
 sg13g2_a221oi_1 _35696_ (.B2(_05105_),
    .C1(_05107_),
    .B1(_04970_),
    .A1(\u_inv.d_next[123] ),
    .Y(_05108_),
    .A2(_18491_));
 sg13g2_nand2_1 _35697_ (.Y(_05109_),
    .A(\u_inv.d_next[124] ),
    .B(_18490_));
 sg13g2_nand2_1 _35698_ (.Y(_05110_),
    .A(\u_inv.d_next[125] ),
    .B(_18489_));
 sg13g2_o21ai_1 _35699_ (.B1(_05110_),
    .Y(_05111_),
    .A1(_03814_),
    .A2(_05109_));
 sg13g2_inv_1 _35700_ (.Y(_05112_),
    .A(_05111_));
 sg13g2_nand2_1 _35701_ (.Y(_05113_),
    .A(\u_inv.d_next[126] ),
    .B(_18488_));
 sg13g2_nor2_1 _35702_ (.A(_03810_),
    .B(_05113_),
    .Y(_05114_));
 sg13g2_a221oi_1 _35703_ (.B2(_05111_),
    .C1(_05114_),
    .B1(_04966_),
    .A1(\u_inv.d_next[127] ),
    .Y(_05115_),
    .A2(_18487_));
 sg13g2_o21ai_1 _35704_ (.B1(_05115_),
    .Y(_05116_),
    .A1(_04969_),
    .A2(_05108_));
 sg13g2_nor2b_1 _35705_ (.A(\u_inv.d_reg[96] ),
    .B_N(\u_inv.d_next[96] ),
    .Y(_05117_));
 sg13g2_a21oi_1 _35706_ (.A1(_03921_),
    .A2(_05117_),
    .Y(_05118_),
    .B1(_03922_));
 sg13g2_inv_1 _35707_ (.Y(_05119_),
    .A(_05118_));
 sg13g2_nor2_1 _35708_ (.A(_04992_),
    .B(_05118_),
    .Y(_05120_));
 sg13g2_nor2b_1 _35709_ (.A(\u_inv.d_reg[100] ),
    .B_N(\u_inv.d_next[100] ),
    .Y(_05121_));
 sg13g2_nand2_1 _35710_ (.Y(_05122_),
    .A(_03908_),
    .B(_05121_));
 sg13g2_nand2_1 _35711_ (.Y(_05123_),
    .A(\u_inv.d_next[101] ),
    .B(_18513_));
 sg13g2_nand2_1 _35712_ (.Y(_05124_),
    .A(_05122_),
    .B(_05123_));
 sg13g2_nor2b_1 _35713_ (.A(\u_inv.d_reg[102] ),
    .B_N(\u_inv.d_next[102] ),
    .Y(_05125_));
 sg13g2_and2_1 _35714_ (.A(_03912_),
    .B(_05125_),
    .X(_05126_));
 sg13g2_a221oi_1 _35715_ (.B2(_05124_),
    .C1(_05126_),
    .B1(_04989_),
    .A1(\u_inv.d_next[103] ),
    .Y(_05127_),
    .A2(_18511_));
 sg13g2_nor2b_2 _35716_ (.A(\u_inv.d_reg[98] ),
    .B_N(\u_inv.d_next[98] ),
    .Y(_05128_));
 sg13g2_o21ai_1 _35717_ (.B1(_03915_),
    .Y(_05129_),
    .A1(_03916_),
    .A2(_05128_));
 sg13g2_o21ai_1 _35718_ (.B1(_05127_),
    .Y(_05130_),
    .A1(_04990_),
    .A2(_05129_));
 sg13g2_nor2_2 _35719_ (.A(_05120_),
    .B(_05130_),
    .Y(_05131_));
 sg13g2_nor2_1 _35720_ (.A(_18146_),
    .B(\u_inv.d_reg[104] ),
    .Y(_05132_));
 sg13g2_a21oi_1 _35721_ (.A1(\u_inv.d_next[105] ),
    .A2(_18509_),
    .Y(_05133_),
    .B1(_05132_));
 sg13g2_a21oi_1 _35722_ (.A1(_18145_),
    .A2(\u_inv.d_reg[105] ),
    .Y(_05134_),
    .B1(_05133_));
 sg13g2_nand2_1 _35723_ (.Y(_05135_),
    .A(\u_inv.d_next[106] ),
    .B(_18508_));
 sg13g2_a22oi_1 _35724_ (.Y(_05136_),
    .B1(_04985_),
    .B2(_05134_),
    .A2(_18507_),
    .A1(\u_inv.d_next[107] ));
 sg13g2_o21ai_1 _35725_ (.B1(_05136_),
    .Y(_05137_),
    .A1(_03890_),
    .A2(_05135_));
 sg13g2_nand2_1 _35726_ (.Y(_05138_),
    .A(\u_inv.d_next[108] ),
    .B(_18506_));
 sg13g2_o21ai_1 _35727_ (.B1(_03886_),
    .Y(_05139_),
    .A1(_03885_),
    .A2(_05138_));
 sg13g2_nand2_1 _35728_ (.Y(_05140_),
    .A(\u_inv.d_next[111] ),
    .B(_18503_));
 sg13g2_nand2_1 _35729_ (.Y(_05141_),
    .A(\u_inv.d_next[110] ),
    .B(_18504_));
 sg13g2_o21ai_1 _35730_ (.B1(_05140_),
    .Y(_05142_),
    .A1(_03877_),
    .A2(_05141_));
 sg13g2_a221oi_1 _35731_ (.B2(_04982_),
    .C1(_05142_),
    .B1(_05139_),
    .A1(_04984_),
    .Y(_05143_),
    .A2(_05137_));
 sg13g2_o21ai_1 _35732_ (.B1(_05143_),
    .Y(_05144_),
    .A1(_04988_),
    .A2(_05131_));
 sg13g2_a221oi_1 _35733_ (.B2(_04981_),
    .C1(_05116_),
    .B1(_05144_),
    .A1(_04972_),
    .Y(_05145_),
    .A2(_05103_));
 sg13g2_o21ai_1 _35734_ (.B1(_05145_),
    .Y(_05146_),
    .A1(_04996_),
    .A2(_05088_));
 sg13g2_a21oi_2 _35735_ (.B1(_05146_),
    .Y(_05147_),
    .A2(_04965_),
    .A1(_05031_));
 sg13g2_a21o_2 _35736_ (.A2(_05031_),
    .A1(_04965_),
    .B1(_05146_),
    .X(_05148_));
 sg13g2_nor2_1 _35737_ (.A(_03674_),
    .B(_03677_),
    .Y(_05149_));
 sg13g2_nor2_1 _35738_ (.A(_03682_),
    .B(_03685_),
    .Y(_05150_));
 sg13g2_nand2_1 _35739_ (.Y(_05151_),
    .A(_05149_),
    .B(_05150_));
 sg13g2_nand2_1 _35740_ (.Y(_05152_),
    .A(_03697_),
    .B(_03699_));
 sg13g2_nor2_1 _35741_ (.A(_03689_),
    .B(_03692_),
    .Y(_05153_));
 sg13g2_nor4_1 _35742_ (.A(_03689_),
    .B(_03692_),
    .C(_05151_),
    .D(_05152_),
    .Y(_05154_));
 sg13g2_nand2_1 _35743_ (.Y(_05155_),
    .A(_03664_),
    .B(_03668_));
 sg13g2_nand4_1 _35744_ (.B(_03668_),
    .C(_03669_),
    .A(_03664_),
    .Y(_05156_),
    .D(_03671_));
 sg13g2_and2_1 _35745_ (.A(_03705_),
    .B(_03713_),
    .X(_05157_));
 sg13g2_nor2_1 _35746_ (.A(_03707_),
    .B(_03710_),
    .Y(_05158_));
 sg13g2_nand2_1 _35747_ (.Y(_05159_),
    .A(_05157_),
    .B(_05158_));
 sg13g2_nor2_1 _35748_ (.A(_05156_),
    .B(_05159_),
    .Y(_05160_));
 sg13g2_nand2_2 _35749_ (.Y(_05161_),
    .A(_05154_),
    .B(_05160_));
 sg13g2_nand2_1 _35750_ (.Y(_05162_),
    .A(_03743_),
    .B(_03745_));
 sg13g2_nand2_1 _35751_ (.Y(_05163_),
    .A(_03750_),
    .B(_03752_));
 sg13g2_inv_1 _35752_ (.Y(_05164_),
    .A(_05163_));
 sg13g2_nor2_1 _35753_ (.A(_05162_),
    .B(_05163_),
    .Y(_05165_));
 sg13g2_nand2_1 _35754_ (.Y(_05166_),
    .A(_03757_),
    .B(_03760_));
 sg13g2_or2_1 _35755_ (.X(_05167_),
    .B(_03765_),
    .A(_03762_));
 sg13g2_nor4_1 _35756_ (.A(_05162_),
    .B(_05163_),
    .C(_05166_),
    .D(_05167_),
    .Y(_05168_));
 sg13g2_nor2_1 _35757_ (.A(_03722_),
    .B(_03724_),
    .Y(_05169_));
 sg13g2_nor4_1 _35758_ (.A(_03719_),
    .B(_03720_),
    .C(_03722_),
    .D(_03724_),
    .Y(_05170_));
 sg13g2_and2_1 _35759_ (.A(_03735_),
    .B(_03737_),
    .X(_05171_));
 sg13g2_and3_2 _35760_ (.X(_05172_),
    .A(_03727_),
    .B(_03732_),
    .C(_05171_));
 sg13g2_and2_1 _35761_ (.A(_05170_),
    .B(_05172_),
    .X(_05173_));
 sg13g2_nand2_1 _35762_ (.Y(_05174_),
    .A(_05168_),
    .B(_05173_));
 sg13g2_nor2_1 _35763_ (.A(_05161_),
    .B(_05174_),
    .Y(_05175_));
 sg13g2_nor2_1 _35764_ (.A(_04455_),
    .B(_04458_),
    .Y(_05176_));
 sg13g2_inv_1 _35765_ (.Y(_05177_),
    .A(_05176_));
 sg13g2_and2_1 _35766_ (.A(_04451_),
    .B(_04452_),
    .X(_05178_));
 sg13g2_nand2_1 _35767_ (.Y(_05179_),
    .A(_05176_),
    .B(_05178_));
 sg13g2_or2_1 _35768_ (.X(_05180_),
    .B(_04466_),
    .A(_04463_));
 sg13g2_and2_1 _35769_ (.A(_04470_),
    .B(_04472_),
    .X(_05181_));
 sg13g2_nand3_1 _35770_ (.B(_05178_),
    .C(_05181_),
    .A(_05176_),
    .Y(_05182_));
 sg13g2_nor2_1 _35771_ (.A(_05180_),
    .B(_05182_),
    .Y(_05183_));
 sg13g2_and2_1 _35772_ (.A(_04429_),
    .B(_04431_),
    .X(_05184_));
 sg13g2_and3_1 _35773_ (.X(_05185_),
    .A(_04424_),
    .B(_04427_),
    .C(_05184_));
 sg13g2_nand2_1 _35774_ (.Y(_05186_),
    .A(_04437_),
    .B(_04438_));
 sg13g2_nand2_1 _35775_ (.Y(_05187_),
    .A(_04443_),
    .B(_04447_));
 sg13g2_nor2_1 _35776_ (.A(_05186_),
    .B(_05187_),
    .Y(_05188_));
 sg13g2_and2_1 _35777_ (.A(_05185_),
    .B(_05188_),
    .X(_05189_));
 sg13g2_inv_1 _35778_ (.Y(_05190_),
    .A(_05189_));
 sg13g2_nor2_1 _35779_ (.A(_04476_),
    .B(_04479_),
    .Y(_05191_));
 sg13g2_nor2_1 _35780_ (.A(_04480_),
    .B(_04482_),
    .Y(_05192_));
 sg13g2_and2_1 _35781_ (.A(_05191_),
    .B(_05192_),
    .X(_05193_));
 sg13g2_and2_1 _35782_ (.A(_04491_),
    .B(_04493_),
    .X(_05194_));
 sg13g2_nor2_1 _35783_ (.A(_04485_),
    .B(_04488_),
    .Y(_05195_));
 sg13g2_nand3_1 _35784_ (.B(_05194_),
    .C(_05195_),
    .A(_05193_),
    .Y(_05196_));
 sg13g2_nor2_1 _35785_ (.A(_04503_),
    .B(_04505_),
    .Y(_05197_));
 sg13g2_nor2_1 _35786_ (.A(_04497_),
    .B(_04500_),
    .Y(_05198_));
 sg13g2_nand2_1 _35787_ (.Y(_05199_),
    .A(_05197_),
    .B(_05198_));
 sg13g2_nor2_1 _35788_ (.A(_04510_),
    .B(_04513_),
    .Y(_05200_));
 sg13g2_nand2_1 _35789_ (.Y(_05201_),
    .A(_04511_),
    .B(_04512_));
 sg13g2_nor2_1 _35790_ (.A(_04517_),
    .B(net6994),
    .Y(_05202_));
 sg13g2_nand4_1 _35791_ (.B(_05198_),
    .C(_05200_),
    .A(_05197_),
    .Y(_05203_),
    .D(_05202_));
 sg13g2_nor2_2 _35792_ (.A(_05196_),
    .B(_05203_),
    .Y(_05204_));
 sg13g2_and3_2 _35793_ (.X(_05205_),
    .A(_05183_),
    .B(_05189_),
    .C(_05204_));
 sg13g2_and2_1 _35794_ (.A(_05175_),
    .B(_05205_),
    .X(_05206_));
 sg13g2_nand2_1 _35795_ (.Y(_05207_),
    .A(_05175_),
    .B(_05205_));
 sg13g2_nand2b_1 _35796_ (.Y(_05208_),
    .B(\u_inv.d_next[128] ),
    .A_N(\u_inv.d_reg[128] ));
 sg13g2_o21ai_1 _35797_ (.B1(_04515_),
    .Y(_05209_),
    .A1(_04514_),
    .A2(_05208_));
 sg13g2_nand2_1 _35798_ (.Y(_05210_),
    .A(_05200_),
    .B(_05209_));
 sg13g2_nand2b_1 _35799_ (.Y(_05211_),
    .B(net7296),
    .A_N(net7289));
 sg13g2_a21oi_1 _35800_ (.A1(_18135_),
    .A2(\u_inv.d_reg[131] ),
    .Y(_05212_),
    .B1(_05211_));
 sg13g2_a21oi_1 _35801_ (.A1(\u_inv.d_next[131] ),
    .A2(_18483_),
    .Y(_05213_),
    .B1(_05212_));
 sg13g2_a21oi_1 _35802_ (.A1(_05210_),
    .A2(_05213_),
    .Y(_05214_),
    .B1(_05199_));
 sg13g2_nor2b_1 _35803_ (.A(\u_inv.d_reg[132] ),
    .B_N(\u_inv.d_next[132] ),
    .Y(_05215_));
 sg13g2_a21oi_1 _35804_ (.A1(\u_inv.d_next[133] ),
    .A2(_18481_),
    .Y(_05216_),
    .B1(_05215_));
 sg13g2_a21oi_1 _35805_ (.A1(_18134_),
    .A2(\u_inv.d_reg[133] ),
    .Y(_05217_),
    .B1(_05216_));
 sg13g2_nand2_1 _35806_ (.Y(_05218_),
    .A(\u_inv.d_next[134] ),
    .B(_18480_));
 sg13g2_nor2_1 _35807_ (.A(_04497_),
    .B(_05218_),
    .Y(_05219_));
 sg13g2_a221oi_1 _35808_ (.B2(_05217_),
    .C1(_05219_),
    .B1(_05198_),
    .A1(\u_inv.d_next[135] ),
    .Y(_05220_),
    .A2(_18479_));
 sg13g2_nor2b_2 _35809_ (.A(_05214_),
    .B_N(_05220_),
    .Y(_05221_));
 sg13g2_nand2_1 _35810_ (.Y(_05222_),
    .A(\u_inv.d_next[140] ),
    .B(_18474_));
 sg13g2_nand2_1 _35811_ (.Y(_05223_),
    .A(\u_inv.d_next[141] ),
    .B(_18473_));
 sg13g2_o21ai_1 _35812_ (.B1(_05223_),
    .Y(_05224_),
    .A1(_04480_),
    .A2(_05222_));
 sg13g2_nand2_1 _35813_ (.Y(_05225_),
    .A(\u_inv.d_next[143] ),
    .B(_18471_));
 sg13g2_nand2_1 _35814_ (.Y(_05226_),
    .A(\u_inv.d_next[142] ),
    .B(_18472_));
 sg13g2_o21ai_1 _35815_ (.B1(_05225_),
    .Y(_05227_),
    .A1(_04476_),
    .A2(_05226_));
 sg13g2_nand2_1 _35816_ (.Y(_05228_),
    .A(\u_inv.d_next[138] ),
    .B(_18476_));
 sg13g2_nand2_1 _35817_ (.Y(_05229_),
    .A(\u_inv.d_next[139] ),
    .B(_18475_));
 sg13g2_o21ai_1 _35818_ (.B1(_05229_),
    .Y(_05230_),
    .A1(_04485_),
    .A2(_05228_));
 sg13g2_nor2b_1 _35819_ (.A(\u_inv.d_reg[136] ),
    .B_N(\u_inv.d_next[136] ),
    .Y(_05231_));
 sg13g2_a21oi_1 _35820_ (.A1(\u_inv.d_next[137] ),
    .A2(_18477_),
    .Y(_05232_),
    .B1(_05231_));
 sg13g2_a21oi_1 _35821_ (.A1(_18132_),
    .A2(\u_inv.d_reg[137] ),
    .Y(_05233_),
    .B1(_05232_));
 sg13g2_a21o_1 _35822_ (.A2(_05233_),
    .A1(_05195_),
    .B1(_05230_),
    .X(_05234_));
 sg13g2_a221oi_1 _35823_ (.B2(_05193_),
    .C1(_05227_),
    .B1(_05234_),
    .A1(_05191_),
    .Y(_05235_),
    .A2(_05224_));
 sg13g2_o21ai_1 _35824_ (.B1(_05235_),
    .Y(_05236_),
    .A1(_05196_),
    .A2(_05221_));
 sg13g2_nand3_1 _35825_ (.B(_05189_),
    .C(_05236_),
    .A(_05183_),
    .Y(_05237_));
 sg13g2_nor2b_1 _35826_ (.A(\u_inv.d_reg[152] ),
    .B_N(\u_inv.d_next[152] ),
    .Y(_05238_));
 sg13g2_nor2b_1 _35827_ (.A(\u_inv.d_reg[153] ),
    .B_N(\u_inv.d_next[153] ),
    .Y(_05239_));
 sg13g2_a21oi_1 _35828_ (.A1(_04470_),
    .A2(_05238_),
    .Y(_05240_),
    .B1(_05239_));
 sg13g2_inv_1 _35829_ (.Y(_05241_),
    .A(_05240_));
 sg13g2_nand2_1 _35830_ (.Y(_05242_),
    .A(\u_inv.d_next[154] ),
    .B(_18460_));
 sg13g2_nand2b_1 _35831_ (.Y(_05243_),
    .B(_04464_),
    .A_N(_05242_));
 sg13g2_o21ai_1 _35832_ (.B1(_05243_),
    .Y(_05244_),
    .A1(_05180_),
    .A2(_05240_));
 sg13g2_a21oi_1 _35833_ (.A1(\u_inv.d_next[155] ),
    .A2(_18459_),
    .Y(_05245_),
    .B1(_05244_));
 sg13g2_nor2_1 _35834_ (.A(_05179_),
    .B(_05245_),
    .Y(_05246_));
 sg13g2_nand2_1 _35835_ (.Y(_05247_),
    .A(\u_inv.d_next[158] ),
    .B(_18456_));
 sg13g2_nor2b_1 _35836_ (.A(\u_inv.d_reg[156] ),
    .B_N(\u_inv.d_next[156] ),
    .Y(_05248_));
 sg13g2_nor2b_1 _35837_ (.A(\u_inv.d_reg[157] ),
    .B_N(\u_inv.d_next[157] ),
    .Y(_05249_));
 sg13g2_a21o_1 _35838_ (.A2(_05248_),
    .A1(_04456_),
    .B1(_05249_),
    .X(_05250_));
 sg13g2_nand3_1 _35839_ (.B(_18456_),
    .C(_04452_),
    .A(\u_inv.d_next[158] ),
    .Y(_05251_));
 sg13g2_nand2b_1 _35840_ (.Y(_05252_),
    .B(\u_inv.d_next[144] ),
    .A_N(\u_inv.d_reg[144] ));
 sg13g2_o21ai_1 _35841_ (.B1(_04442_),
    .Y(_05253_),
    .A1(_04441_),
    .A2(_05252_));
 sg13g2_inv_1 _35842_ (.Y(_05254_),
    .A(_05253_));
 sg13g2_nand2_1 _35843_ (.Y(_05255_),
    .A(\u_inv.d_next[147] ),
    .B(_18467_));
 sg13g2_nor2b_1 _35844_ (.A(\u_inv.d_reg[146] ),
    .B_N(\u_inv.d_next[146] ),
    .Y(_05256_));
 sg13g2_a21oi_1 _35845_ (.A1(_04438_),
    .A2(_05253_),
    .Y(_05257_),
    .B1(_05256_));
 sg13g2_o21ai_1 _35846_ (.B1(_05255_),
    .Y(_05258_),
    .A1(_04436_),
    .A2(_05257_));
 sg13g2_nor2b_1 _35847_ (.A(\u_inv.d_reg[148] ),
    .B_N(\u_inv.d_next[148] ),
    .Y(_05259_));
 sg13g2_nor2_1 _35848_ (.A(_18129_),
    .B(\u_inv.d_reg[149] ),
    .Y(_05260_));
 sg13g2_a21oi_1 _35849_ (.A1(_04429_),
    .A2(_05259_),
    .Y(_05261_),
    .B1(_05260_));
 sg13g2_nor2_1 _35850_ (.A(_18128_),
    .B(\u_inv.d_reg[150] ),
    .Y(_05262_));
 sg13g2_nor2_1 _35851_ (.A(_04426_),
    .B(_05261_),
    .Y(_05263_));
 sg13g2_nor2_1 _35852_ (.A(_05262_),
    .B(_05263_),
    .Y(_05264_));
 sg13g2_a22oi_1 _35853_ (.Y(_05265_),
    .B1(_05185_),
    .B2(_05258_),
    .A2(_18463_),
    .A1(\u_inv.d_next[151] ));
 sg13g2_o21ai_1 _35854_ (.B1(_05265_),
    .Y(_05266_),
    .A1(_04423_),
    .A2(_05264_));
 sg13g2_inv_1 _35855_ (.Y(_05267_),
    .A(_05266_));
 sg13g2_nand2_1 _35856_ (.Y(_05268_),
    .A(_05183_),
    .B(_05266_));
 sg13g2_a221oi_1 _35857_ (.B2(_05250_),
    .C1(_05246_),
    .B1(_05178_),
    .A1(\u_inv.d_next[159] ),
    .Y(_05269_),
    .A2(_18455_));
 sg13g2_nand4_1 _35858_ (.B(_05251_),
    .C(_05268_),
    .A(_05237_),
    .Y(_05270_),
    .D(_05269_));
 sg13g2_nand2_1 _35859_ (.Y(_05271_),
    .A(_05175_),
    .B(_05270_));
 sg13g2_nand2_1 _35860_ (.Y(_05272_),
    .A(\u_inv.d_next[179] ),
    .B(_18435_));
 sg13g2_nand2_1 _35861_ (.Y(_05273_),
    .A(\u_inv.d_next[178] ),
    .B(_18436_));
 sg13g2_nor2b_1 _35862_ (.A(\u_inv.d_reg[176] ),
    .B_N(\u_inv.d_next[176] ),
    .Y(_05274_));
 sg13g2_nor2_1 _35863_ (.A(_18121_),
    .B(\u_inv.d_reg[177] ),
    .Y(_05275_));
 sg13g2_a21o_1 _35864_ (.A2(_05274_),
    .A1(_03735_),
    .B1(_05275_),
    .X(_05276_));
 sg13g2_nand2_1 _35865_ (.Y(_05277_),
    .A(_03727_),
    .B(_05276_));
 sg13g2_and2_1 _35866_ (.A(_05273_),
    .B(_05277_),
    .X(_05278_));
 sg13g2_o21ai_1 _35867_ (.B1(_05272_),
    .Y(_05279_),
    .A1(_03731_),
    .A2(_05278_));
 sg13g2_nand2_1 _35868_ (.Y(_05280_),
    .A(_05170_),
    .B(_05279_));
 sg13g2_nand2_1 _35869_ (.Y(_05281_),
    .A(\u_inv.d_next[183] ),
    .B(_18431_));
 sg13g2_nand2_1 _35870_ (.Y(_05282_),
    .A(\u_inv.d_next[182] ),
    .B(_18432_));
 sg13g2_nand2_1 _35871_ (.Y(_05283_),
    .A(\u_inv.d_next[180] ),
    .B(_18434_));
 sg13g2_nor2_1 _35872_ (.A(_03722_),
    .B(_05283_),
    .Y(_05284_));
 sg13g2_a21oi_1 _35873_ (.A1(\u_inv.d_next[181] ),
    .A2(_18433_),
    .Y(_05285_),
    .B1(_05284_));
 sg13g2_o21ai_1 _35874_ (.B1(_05282_),
    .Y(_05286_),
    .A1(_03719_),
    .A2(_05285_));
 sg13g2_nand2b_1 _35875_ (.Y(_05287_),
    .B(_05286_),
    .A_N(_03720_));
 sg13g2_nand3_1 _35876_ (.B(_05281_),
    .C(_05287_),
    .A(_05280_),
    .Y(_05288_));
 sg13g2_nand2_1 _35877_ (.Y(_05289_),
    .A(\u_inv.d_next[187] ),
    .B(_18427_));
 sg13g2_nor2b_1 _35878_ (.A(\u_inv.d_reg[186] ),
    .B_N(\u_inv.d_next[186] ),
    .Y(_05290_));
 sg13g2_nand2_1 _35879_ (.Y(_05291_),
    .A(\u_inv.d_next[184] ),
    .B(_18430_));
 sg13g2_nand2_1 _35880_ (.Y(_05292_),
    .A(\u_inv.d_next[185] ),
    .B(_18429_));
 sg13g2_o21ai_1 _35881_ (.B1(_05292_),
    .Y(_05293_),
    .A1(_03762_),
    .A2(_05291_));
 sg13g2_inv_1 _35882_ (.Y(_05294_),
    .A(_05293_));
 sg13g2_a21oi_1 _35883_ (.A1(_03760_),
    .A2(_05293_),
    .Y(_05295_),
    .B1(_05290_));
 sg13g2_o21ai_1 _35884_ (.B1(_05289_),
    .Y(_05296_),
    .A1(_03758_),
    .A2(_05295_));
 sg13g2_nand2_1 _35885_ (.Y(_05297_),
    .A(\u_inv.d_next[188] ),
    .B(_18426_));
 sg13g2_nor2b_1 _35886_ (.A(_05297_),
    .B_N(_03750_),
    .Y(_05298_));
 sg13g2_a21oi_1 _35887_ (.A1(\u_inv.d_next[189] ),
    .A2(_18425_),
    .Y(_05299_),
    .B1(_05298_));
 sg13g2_nor2b_1 _35888_ (.A(\u_inv.d_reg[190] ),
    .B_N(\u_inv.d_next[190] ),
    .Y(_05300_));
 sg13g2_nand2_1 _35889_ (.Y(_05301_),
    .A(_03743_),
    .B(_05300_));
 sg13g2_nand2_1 _35890_ (.Y(_05302_),
    .A(\u_inv.d_next[191] ),
    .B(_18423_));
 sg13g2_nand2_1 _35891_ (.Y(_05303_),
    .A(\u_inv.d_next[160] ),
    .B(_18454_));
 sg13g2_o21ai_1 _35892_ (.B1(_03663_),
    .Y(_05304_),
    .A1(_03662_),
    .A2(_05303_));
 sg13g2_inv_1 _35893_ (.Y(_05305_),
    .A(_05304_));
 sg13g2_nor2_1 _35894_ (.A(_18125_),
    .B(\u_inv.d_reg[163] ),
    .Y(_05306_));
 sg13g2_nor2b_1 _35895_ (.A(\u_inv.d_reg[162] ),
    .B_N(\u_inv.d_next[162] ),
    .Y(_05307_));
 sg13g2_a21o_1 _35896_ (.A2(_05304_),
    .A1(_03671_),
    .B1(_05307_),
    .X(_05308_));
 sg13g2_a21oi_1 _35897_ (.A1(_03669_),
    .A2(_05308_),
    .Y(_05309_),
    .B1(_05306_));
 sg13g2_nor2b_1 _35898_ (.A(\u_inv.d_reg[164] ),
    .B_N(\u_inv.d_next[164] ),
    .Y(_05310_));
 sg13g2_nor2_1 _35899_ (.A(_18124_),
    .B(\u_inv.d_reg[165] ),
    .Y(_05311_));
 sg13g2_a21o_1 _35900_ (.A2(_05310_),
    .A1(_03713_),
    .B1(_05311_),
    .X(_05312_));
 sg13g2_nand2_1 _35901_ (.Y(_05313_),
    .A(\u_inv.d_next[166] ),
    .B(_18448_));
 sg13g2_nor2_1 _35902_ (.A(_03710_),
    .B(_05313_),
    .Y(_05314_));
 sg13g2_a221oi_1 _35903_ (.B2(_05312_),
    .C1(_05314_),
    .B1(_05158_),
    .A1(\u_inv.d_next[167] ),
    .Y(_05315_),
    .A2(_18447_));
 sg13g2_o21ai_1 _35904_ (.B1(_05315_),
    .Y(_05316_),
    .A1(_05159_),
    .A2(_05309_));
 sg13g2_nand2_1 _35905_ (.Y(_05317_),
    .A(\u_inv.d_next[168] ),
    .B(_18446_));
 sg13g2_nor2_1 _35906_ (.A(_03689_),
    .B(_05317_),
    .Y(_05318_));
 sg13g2_a21o_1 _35907_ (.A2(_18445_),
    .A1(\u_inv.d_next[169] ),
    .B1(_05318_),
    .X(_05319_));
 sg13g2_nor2b_1 _35908_ (.A(\u_inv.d_reg[170] ),
    .B_N(\u_inv.d_next[170] ),
    .Y(_05320_));
 sg13g2_a21oi_1 _35909_ (.A1(_03699_),
    .A2(_05319_),
    .Y(_05321_),
    .B1(_05320_));
 sg13g2_nor2_1 _35910_ (.A(_03696_),
    .B(_05321_),
    .Y(_05322_));
 sg13g2_a21oi_1 _35911_ (.A1(\u_inv.d_next[171] ),
    .A2(_18443_),
    .Y(_05323_),
    .B1(_05322_));
 sg13g2_nor2b_1 _35912_ (.A(\u_inv.d_reg[172] ),
    .B_N(\u_inv.d_next[172] ),
    .Y(_05324_));
 sg13g2_nor2b_1 _35913_ (.A(\u_inv.d_reg[173] ),
    .B_N(\u_inv.d_next[173] ),
    .Y(_05325_));
 sg13g2_a21o_1 _35914_ (.A2(_05324_),
    .A1(_03683_),
    .B1(_05325_),
    .X(_05326_));
 sg13g2_nand2_1 _35915_ (.Y(_05327_),
    .A(\u_inv.d_next[174] ),
    .B(_18440_));
 sg13g2_nand2_1 _35916_ (.Y(_05328_),
    .A(\u_inv.d_next[175] ),
    .B(_18439_));
 sg13g2_o21ai_1 _35917_ (.B1(_05328_),
    .Y(_05329_),
    .A1(_03674_),
    .A2(_05327_));
 sg13g2_a221oi_1 _35918_ (.B2(_05149_),
    .C1(_05329_),
    .B1(_05326_),
    .A1(_05154_),
    .Y(_05330_),
    .A2(_05316_));
 sg13g2_o21ai_1 _35919_ (.B1(_05330_),
    .Y(_05331_),
    .A1(_05151_),
    .A2(_05323_));
 sg13g2_inv_1 _35920_ (.Y(_05332_),
    .A(_05331_));
 sg13g2_nand2b_1 _35921_ (.Y(_05333_),
    .B(_05331_),
    .A_N(_05174_));
 sg13g2_o21ai_1 _35922_ (.B1(_05301_),
    .Y(_05334_),
    .A1(_05162_),
    .A2(_05299_));
 sg13g2_a221oi_1 _35923_ (.B2(_05165_),
    .C1(_05334_),
    .B1(_05296_),
    .A1(_05168_),
    .Y(_05335_),
    .A2(_05288_));
 sg13g2_nand4_1 _35924_ (.B(_05302_),
    .C(_05333_),
    .A(_05271_),
    .Y(_05336_),
    .D(_05335_));
 sg13g2_nor3_1 _35925_ (.A(_04654_),
    .B(net1104),
    .C(_05207_),
    .Y(_05337_));
 sg13g2_nand2b_1 _35926_ (.Y(_05338_),
    .B(_05336_),
    .A_N(_04654_));
 sg13g2_nand4_1 _35927_ (.B(_04746_),
    .C(_04778_),
    .A(_04715_),
    .Y(_05339_),
    .D(_05338_));
 sg13g2_o21ai_1 _35928_ (.B1(_03355_),
    .Y(_05340_),
    .A1(_05337_),
    .A2(_05339_));
 sg13g2_a21oi_2 _35929_ (.B1(net6216),
    .Y(_05341_),
    .A2(\u_inv.d_reg[256] ),
    .A1(_18100_));
 sg13g2_a21oi_1 _35930_ (.A1(_05340_),
    .A2(_05341_),
    .Y(_05342_),
    .B1(_04593_));
 sg13g2_a21o_1 _35931_ (.A2(_05341_),
    .A1(_05340_),
    .B1(_04593_),
    .X(_05343_));
 sg13g2_nand2_2 _35932_ (.Y(_05344_),
    .A(net6801),
    .B(net5845));
 sg13g2_nand2_1 _35933_ (.Y(_05345_),
    .A(\u_inv.d_reg[0] ),
    .B(net6299));
 sg13g2_xnor2_1 _35934_ (.Y(_05346_),
    .A(_03340_),
    .B(_03347_));
 sg13g2_nand2_1 _35935_ (.Y(_05347_),
    .A(net7330),
    .B(_05346_));
 sg13g2_o21ai_1 _35936_ (.B1(_05347_),
    .Y(_05348_),
    .A1(net7330),
    .A2(\u_inv.d_next[1] ));
 sg13g2_xnor2_1 _35937_ (.Y(_05349_),
    .A(_05345_),
    .B(_05348_));
 sg13g2_nor2_1 _35938_ (.A(_05344_),
    .B(_05349_),
    .Y(_05350_));
 sg13g2_xor2_1 _35939_ (.B(_05349_),
    .A(_05344_),
    .X(_05351_));
 sg13g2_xnor2_1 _35940_ (.Y(_05352_),
    .A(_05344_),
    .B(_05349_));
 sg13g2_a21oi_2 _35941_ (.B1(_05336_),
    .Y(_05353_),
    .A2(_05206_),
    .A1(_05148_));
 sg13g2_a21o_2 _35942_ (.A2(_05206_),
    .A1(_05148_),
    .B1(_05336_),
    .X(_05354_));
 sg13g2_a21oi_2 _35943_ (.B1(_04714_),
    .Y(_05355_),
    .A2(_05354_),
    .A1(_04653_));
 sg13g2_o21ai_1 _35944_ (.B1(_04713_),
    .Y(_05356_),
    .A1(_04652_),
    .A2(_05353_));
 sg13g2_o21ai_1 _35945_ (.B1(_04745_),
    .Y(_05357_),
    .A1(_04619_),
    .A2(_05355_));
 sg13g2_a21oi_2 _35946_ (.B1(_04762_),
    .Y(_05358_),
    .A2(_05357_),
    .A1(_04604_));
 sg13g2_nor3_2 _35947_ (.A(_04596_),
    .B(_04597_),
    .C(_05358_),
    .Y(_05359_));
 sg13g2_nor2_1 _35948_ (.A(_04770_),
    .B(_05359_),
    .Y(_05360_));
 sg13g2_o21ai_1 _35949_ (.B1(_04594_),
    .Y(_05361_),
    .A1(_04770_),
    .A2(_05359_));
 sg13g2_a21o_1 _35950_ (.A2(_05361_),
    .A1(_04774_),
    .B1(_03570_),
    .X(_05362_));
 sg13g2_nand3_1 _35951_ (.B(_04774_),
    .C(_05361_),
    .A(_03570_),
    .Y(_05363_));
 sg13g2_and2_1 _35952_ (.A(_05362_),
    .B(_05363_),
    .X(_05364_));
 sg13g2_a21oi_2 _35953_ (.B1(_03508_),
    .Y(_05365_),
    .A2(_04587_),
    .A1(net1081));
 sg13g2_o21ai_1 _35954_ (.B1(_03652_),
    .Y(_05366_),
    .A1(_03565_),
    .A2(_05365_));
 sg13g2_and2_1 _35955_ (.A(_03614_),
    .B(_05366_),
    .X(_05367_));
 sg13g2_nand4_1 _35956_ (.B(_03612_),
    .C(_03614_),
    .A(_03610_),
    .Y(_05368_),
    .D(_05366_));
 sg13g2_and2_1 _35957_ (.A(_03629_),
    .B(_05368_),
    .X(_05369_));
 sg13g2_nand2b_1 _35958_ (.Y(_05370_),
    .B(_03585_),
    .A_N(_05369_));
 sg13g2_a21oi_1 _35959_ (.A1(_03629_),
    .A2(_05368_),
    .Y(_05371_),
    .B1(_03588_));
 sg13g2_a21oi_1 _35960_ (.A1(_03592_),
    .A2(_05371_),
    .Y(_05372_),
    .B1(_03633_));
 sg13g2_a21o_1 _35961_ (.A2(_05371_),
    .A1(_03592_),
    .B1(_03633_),
    .X(_05373_));
 sg13g2_a21oi_1 _35962_ (.A1(_03579_),
    .A2(_05373_),
    .Y(_05374_),
    .B1(_03634_));
 sg13g2_xor2_1 _35963_ (.B(_05374_),
    .A(_03570_),
    .X(_05375_));
 sg13g2_o21ai_1 _35964_ (.B1(net6206),
    .Y(_05376_),
    .A1(net7316),
    .A2(\u_inv.d_next[254] ));
 sg13g2_a21oi_1 _35965_ (.A1(net7316),
    .A2(_05375_),
    .Y(_05377_),
    .B1(_05376_));
 sg13g2_a21oi_1 _35966_ (.A1(net6285),
    .A2(_05364_),
    .Y(_05378_),
    .B1(_05377_));
 sg13g2_or2_1 _35967_ (.X(_05379_),
    .B(_05378_),
    .A(net5836));
 sg13g2_xnor2_1 _35968_ (.Y(_05380_),
    .A(net5836),
    .B(_05378_));
 sg13g2_o21ai_1 _35969_ (.B1(_03568_),
    .Y(_05381_),
    .A1(_03569_),
    .A2(_05374_));
 sg13g2_xnor2_1 _35970_ (.Y(_05382_),
    .A(_03567_),
    .B(_05381_));
 sg13g2_nand2_1 _35971_ (.Y(_05383_),
    .A(net7316),
    .B(_05382_));
 sg13g2_nand2_1 _35972_ (.Y(_05384_),
    .A(net7194),
    .B(\u_inv.d_next[255] ));
 sg13g2_and3_1 _35973_ (.X(_05385_),
    .A(net6206),
    .B(_05383_),
    .C(_05384_));
 sg13g2_nand3_1 _35974_ (.B(_05383_),
    .C(_05384_),
    .A(net6208),
    .Y(_05386_));
 sg13g2_and3_1 _35975_ (.X(_05387_),
    .A(_03567_),
    .B(_04771_),
    .C(_05362_));
 sg13g2_a21oi_1 _35976_ (.A1(_04771_),
    .A2(_05362_),
    .Y(_05388_),
    .B1(_03567_));
 sg13g2_nor3_1 _35977_ (.A(net6206),
    .B(_05387_),
    .C(_05388_),
    .Y(_05389_));
 sg13g2_or3_1 _35978_ (.A(net6206),
    .B(_05387_),
    .C(_05388_),
    .X(_05390_));
 sg13g2_nor3_1 _35979_ (.A(net5836),
    .B(_05385_),
    .C(_05389_),
    .Y(_05391_));
 sg13g2_nand3_1 _35980_ (.B(_05386_),
    .C(_05390_),
    .A(net5774),
    .Y(_05392_));
 sg13g2_a21oi_1 _35981_ (.A1(_05386_),
    .A2(_05390_),
    .Y(_05393_),
    .B1(net5774));
 sg13g2_nor2_1 _35982_ (.A(_05391_),
    .B(_05393_),
    .Y(_05394_));
 sg13g2_o21ai_1 _35983_ (.B1(_03576_),
    .Y(_05395_),
    .A1(_03578_),
    .A2(_05372_));
 sg13g2_nand2b_1 _35984_ (.Y(_05396_),
    .B(_03575_),
    .A_N(_05395_));
 sg13g2_a21oi_1 _35985_ (.A1(_03574_),
    .A2(_05395_),
    .Y(_05397_),
    .B1(net7185));
 sg13g2_a221oi_1 _35986_ (.B2(_05397_),
    .C1(net6285),
    .B1(_05396_),
    .A1(net7185),
    .Y(_05398_),
    .A2(\u_inv.d_next[253] ));
 sg13g2_o21ai_1 _35987_ (.B1(_03578_),
    .Y(_05399_),
    .A1(_04770_),
    .A2(_05359_));
 sg13g2_and3_1 _35988_ (.X(_05400_),
    .A(_03575_),
    .B(_04772_),
    .C(_05399_));
 sg13g2_a21oi_1 _35989_ (.A1(_04772_),
    .A2(_05399_),
    .Y(_05401_),
    .B1(_03575_));
 sg13g2_nor3_1 _35990_ (.A(net6206),
    .B(_05400_),
    .C(_05401_),
    .Y(_05402_));
 sg13g2_or3_1 _35991_ (.A(net5836),
    .B(_05398_),
    .C(_05402_),
    .X(_05403_));
 sg13g2_o21ai_1 _35992_ (.B1(net5836),
    .Y(_05404_),
    .A1(_05398_),
    .A2(_05402_));
 sg13g2_xnor2_1 _35993_ (.Y(_05405_),
    .A(_03578_),
    .B(_05360_));
 sg13g2_xnor2_1 _35994_ (.Y(_05406_),
    .A(_03578_),
    .B(_05372_));
 sg13g2_o21ai_1 _35995_ (.B1(net6206),
    .Y(_05407_),
    .A1(net7316),
    .A2(\u_inv.d_next[252] ));
 sg13g2_a21oi_1 _35996_ (.A1(net7316),
    .A2(_05406_),
    .Y(_05408_),
    .B1(_05407_));
 sg13g2_a21oi_2 _35997_ (.B1(_05408_),
    .Y(_05409_),
    .A2(_05405_),
    .A1(net6285));
 sg13g2_nor2_1 _35998_ (.A(net5836),
    .B(_05409_),
    .Y(_05410_));
 sg13g2_inv_1 _35999_ (.Y(_05411_),
    .A(_05410_));
 sg13g2_xnor2_1 _36000_ (.Y(_05412_),
    .A(net5774),
    .B(_05409_));
 sg13g2_and3_1 _36001_ (.X(_05413_),
    .A(_05403_),
    .B(_05404_),
    .C(_05412_));
 sg13g2_nand3_1 _36002_ (.B(_05404_),
    .C(_05412_),
    .A(_05403_),
    .Y(_05414_));
 sg13g2_nor4_2 _36003_ (.A(_05380_),
    .B(_05391_),
    .C(_05393_),
    .Y(_05415_),
    .D(_05414_));
 sg13g2_o21ai_1 _36004_ (.B1(_04766_),
    .Y(_05416_),
    .A1(_04597_),
    .A2(_05358_));
 sg13g2_xnor2_1 _36005_ (.Y(_05417_),
    .A(_03591_),
    .B(_05416_));
 sg13g2_or2_1 _36006_ (.X(_05418_),
    .B(_05371_),
    .A(_03630_));
 sg13g2_nand2b_1 _36007_ (.Y(_05419_),
    .B(_03591_),
    .A_N(_05418_));
 sg13g2_nand2b_1 _36008_ (.Y(_05420_),
    .B(_05418_),
    .A_N(_03591_));
 sg13g2_nand3_1 _36009_ (.B(_05419_),
    .C(_05420_),
    .A(net7316),
    .Y(_05421_));
 sg13g2_a21oi_1 _36010_ (.A1(net7185),
    .A2(\u_inv.d_next[250] ),
    .Y(_05422_),
    .B1(net6285));
 sg13g2_a22oi_1 _36011_ (.Y(_05423_),
    .B1(_05421_),
    .B2(_05422_),
    .A2(_05417_),
    .A1(net6285));
 sg13g2_nand2_1 _36012_ (.Y(_05424_),
    .A(net5774),
    .B(_05423_));
 sg13g2_or2_1 _36013_ (.X(_05425_),
    .B(_05423_),
    .A(net5774));
 sg13g2_and2_1 _36014_ (.A(_05424_),
    .B(_05425_),
    .X(_05426_));
 sg13g2_a21o_1 _36015_ (.A2(_05420_),
    .A1(_03590_),
    .B1(_03589_),
    .X(_05427_));
 sg13g2_nand3_1 _36016_ (.B(_03590_),
    .C(_05420_),
    .A(_03589_),
    .Y(_05428_));
 sg13g2_nand3_1 _36017_ (.B(_05427_),
    .C(_05428_),
    .A(net7316),
    .Y(_05429_));
 sg13g2_a21oi_1 _36018_ (.A1(net7185),
    .A2(\u_inv.d_next[251] ),
    .Y(_05430_),
    .B1(net6285));
 sg13g2_a21oi_1 _36019_ (.A1(_03591_),
    .A2(_05416_),
    .Y(_05431_),
    .B1(_04768_));
 sg13g2_or2_1 _36020_ (.X(_05432_),
    .B(_05431_),
    .A(_03589_));
 sg13g2_a21oi_1 _36021_ (.A1(_03589_),
    .A2(_05431_),
    .Y(_05433_),
    .B1(net6206));
 sg13g2_a22oi_1 _36022_ (.Y(_05434_),
    .B1(_05432_),
    .B2(_05433_),
    .A2(_05430_),
    .A1(_05429_));
 sg13g2_xnor2_1 _36023_ (.Y(_05435_),
    .A(net5774),
    .B(_05434_));
 sg13g2_nand3b_1 _36024_ (.B(_05425_),
    .C(_05424_),
    .Y(_05436_),
    .A_N(_05435_));
 sg13g2_o21ai_1 _36025_ (.B1(_03584_),
    .Y(_05437_),
    .A1(_03586_),
    .A2(_05369_));
 sg13g2_o21ai_1 _36026_ (.B1(net7319),
    .Y(_05438_),
    .A1(_03583_),
    .A2(_05437_));
 sg13g2_a21o_1 _36027_ (.A2(_05437_),
    .A1(_03583_),
    .B1(_05438_),
    .X(_05439_));
 sg13g2_a21oi_1 _36028_ (.A1(net7185),
    .A2(\u_inv.d_next[249] ),
    .Y(_05440_),
    .B1(net6285));
 sg13g2_o21ai_1 _36029_ (.B1(_04763_),
    .Y(_05441_),
    .A1(_03585_),
    .A2(_05358_));
 sg13g2_or2_1 _36030_ (.X(_05442_),
    .B(_05441_),
    .A(_03583_));
 sg13g2_a21oi_1 _36031_ (.A1(_03583_),
    .A2(_05441_),
    .Y(_05443_),
    .B1(net6206));
 sg13g2_a22oi_1 _36032_ (.Y(_05444_),
    .B1(_05442_),
    .B2(_05443_),
    .A2(_05440_),
    .A1(_05439_));
 sg13g2_nand2_1 _36033_ (.Y(_05445_),
    .A(net5774),
    .B(_05444_));
 sg13g2_xnor2_1 _36034_ (.Y(_05446_),
    .A(net5774),
    .B(_05444_));
 sg13g2_xnor2_1 _36035_ (.Y(_05447_),
    .A(_03585_),
    .B(_05358_));
 sg13g2_a21oi_1 _36036_ (.A1(_03586_),
    .A2(_05369_),
    .Y(_05448_),
    .B1(net7187));
 sg13g2_a221oi_1 _36037_ (.B2(_05448_),
    .C1(net6288),
    .B1(_05370_),
    .A1(net7187),
    .Y(_05449_),
    .A2(\u_inv.d_next[248] ));
 sg13g2_a21oi_2 _36038_ (.B1(_05449_),
    .Y(_05450_),
    .A2(_05447_),
    .A1(net6288));
 sg13g2_nand2_1 _36039_ (.Y(_05451_),
    .A(net5776),
    .B(_05450_));
 sg13g2_xnor2_1 _36040_ (.Y(_05452_),
    .A(net5836),
    .B(_05450_));
 sg13g2_inv_1 _36041_ (.Y(_05453_),
    .A(_05452_));
 sg13g2_nand2b_1 _36042_ (.Y(_05454_),
    .B(_05452_),
    .A_N(_05446_));
 sg13g2_nor2_2 _36043_ (.A(_05436_),
    .B(_05454_),
    .Y(_05455_));
 sg13g2_inv_1 _36044_ (.Y(_05456_),
    .A(_05455_));
 sg13g2_a21oi_1 _36045_ (.A1(_04603_),
    .A2(_05357_),
    .Y(_05457_),
    .B1(_04753_));
 sg13g2_a21o_1 _36046_ (.A2(_05357_),
    .A1(_04603_),
    .B1(_04753_),
    .X(_05458_));
 sg13g2_a221oi_1 _36047_ (.B2(_05458_),
    .C1(_04758_),
    .B1(_04600_),
    .A1(net7295),
    .Y(_05459_),
    .A2(_18369_));
 sg13g2_a21oi_1 _36048_ (.A1(_03601_),
    .A2(_05459_),
    .Y(_05460_),
    .B1(net6209));
 sg13g2_o21ai_1 _36049_ (.B1(_05460_),
    .Y(_05461_),
    .A1(_03601_),
    .A2(_05459_));
 sg13g2_a21o_1 _36050_ (.A2(\u_inv.d_reg[240] ),
    .A1(\u_inv.d_next[240] ),
    .B1(_05367_),
    .X(_05462_));
 sg13g2_nand3_1 _36051_ (.B(_03614_),
    .C(_05366_),
    .A(_03598_),
    .Y(_05463_));
 sg13g2_a21oi_1 _36052_ (.A1(_03622_),
    .A2(_05463_),
    .Y(_05464_),
    .B1(_03611_));
 sg13g2_o21ai_1 _36053_ (.B1(_03597_),
    .Y(_05465_),
    .A1(_03625_),
    .A2(_05464_));
 sg13g2_and3_1 _36054_ (.X(_05466_),
    .A(_03602_),
    .B(_03619_),
    .C(_05465_));
 sg13g2_a21oi_1 _36055_ (.A1(_03619_),
    .A2(_05465_),
    .Y(_05467_),
    .B1(_03602_));
 sg13g2_nor2_1 _36056_ (.A(_05466_),
    .B(_05467_),
    .Y(_05468_));
 sg13g2_nor2_1 _36057_ (.A(net7187),
    .B(_05468_),
    .Y(_05469_));
 sg13g2_o21ai_1 _36058_ (.B1(net6209),
    .Y(_05470_),
    .A1(net7322),
    .A2(\u_inv.d_next[246] ));
 sg13g2_o21ai_1 _36059_ (.B1(_05461_),
    .Y(_05471_),
    .A1(_05469_),
    .A2(_05470_));
 sg13g2_nand2_1 _36060_ (.Y(_05472_),
    .A(net5775),
    .B(_05471_));
 sg13g2_inv_1 _36061_ (.Y(_05473_),
    .A(_05472_));
 sg13g2_xnor2_1 _36062_ (.Y(_05474_),
    .A(net5836),
    .B(_05471_));
 sg13g2_xnor2_1 _36063_ (.Y(_05475_),
    .A(net5775),
    .B(_05471_));
 sg13g2_or3_1 _36064_ (.A(_03600_),
    .B(_03603_),
    .C(_05467_),
    .X(_05476_));
 sg13g2_o21ai_1 _36065_ (.B1(_03603_),
    .Y(_05477_),
    .A1(_03600_),
    .A2(_05467_));
 sg13g2_nand3_1 _36066_ (.B(_05476_),
    .C(_05477_),
    .A(net7322),
    .Y(_05478_));
 sg13g2_a21oi_1 _36067_ (.A1(net7187),
    .A2(\u_inv.d_next[247] ),
    .Y(_05479_),
    .B1(net6288));
 sg13g2_o21ai_1 _36068_ (.B1(_04756_),
    .Y(_05480_),
    .A1(_03601_),
    .A2(_05459_));
 sg13g2_or2_1 _36069_ (.X(_05481_),
    .B(_05480_),
    .A(_03603_));
 sg13g2_a21oi_1 _36070_ (.A1(_03603_),
    .A2(_05480_),
    .Y(_05482_),
    .B1(net6209));
 sg13g2_a22oi_1 _36071_ (.Y(_05483_),
    .B1(_05481_),
    .B2(_05482_),
    .A2(_05479_),
    .A1(_05478_));
 sg13g2_xnor2_1 _36072_ (.Y(_05484_),
    .A(net5775),
    .B(_05483_));
 sg13g2_xnor2_1 _36073_ (.Y(_05485_),
    .A(_03596_),
    .B(_05457_));
 sg13g2_o21ai_1 _36074_ (.B1(_03596_),
    .Y(_05486_),
    .A1(_03625_),
    .A2(_05464_));
 sg13g2_nor3_1 _36075_ (.A(_03596_),
    .B(_03625_),
    .C(_05464_),
    .Y(_05487_));
 sg13g2_nand3b_1 _36076_ (.B(net7322),
    .C(_05486_),
    .Y(_05488_),
    .A_N(_05487_));
 sg13g2_a21oi_1 _36077_ (.A1(net7187),
    .A2(\u_inv.d_next[244] ),
    .Y(_05489_),
    .B1(net6288));
 sg13g2_a22oi_1 _36078_ (.Y(_05490_),
    .B1(_05488_),
    .B2(_05489_),
    .A2(_05485_),
    .A1(net6288));
 sg13g2_nand2_1 _36079_ (.Y(_05491_),
    .A(net5775),
    .B(_05490_));
 sg13g2_xnor2_1 _36080_ (.Y(_05492_),
    .A(net5775),
    .B(_05490_));
 sg13g2_a21oi_1 _36081_ (.A1(_03595_),
    .A2(_05486_),
    .Y(_05493_),
    .B1(_03594_));
 sg13g2_nand3_1 _36082_ (.B(_03595_),
    .C(_05486_),
    .A(_03594_),
    .Y(_05494_));
 sg13g2_nand3b_1 _36083_ (.B(_05494_),
    .C(net7322),
    .Y(_05495_),
    .A_N(_05493_));
 sg13g2_a21oi_1 _36084_ (.A1(net7187),
    .A2(net7295),
    .Y(_05496_),
    .B1(net6289));
 sg13g2_o21ai_1 _36085_ (.B1(_04757_),
    .Y(_05497_),
    .A1(_03596_),
    .A2(_05457_));
 sg13g2_nand2b_1 _36086_ (.Y(_05498_),
    .B(_03594_),
    .A_N(_05497_));
 sg13g2_a21oi_1 _36087_ (.A1(_03593_),
    .A2(_05497_),
    .Y(_05499_),
    .B1(net6209));
 sg13g2_a22oi_1 _36088_ (.Y(_05500_),
    .B1(_05498_),
    .B2(_05499_),
    .A2(_05496_),
    .A1(_05495_));
 sg13g2_xnor2_1 _36089_ (.Y(_05501_),
    .A(net5775),
    .B(_05500_));
 sg13g2_or2_1 _36090_ (.X(_05502_),
    .B(_05501_),
    .A(_05492_));
 sg13g2_nor3_1 _36091_ (.A(_05475_),
    .B(_05484_),
    .C(_05502_),
    .Y(_05503_));
 sg13g2_a21o_1 _36092_ (.A2(_05357_),
    .A1(_04602_),
    .B1(_04751_),
    .X(_05504_));
 sg13g2_xor2_1 _36093_ (.B(_05504_),
    .A(_03609_),
    .X(_05505_));
 sg13g2_a21oi_1 _36094_ (.A1(_03622_),
    .A2(_05463_),
    .Y(_05506_),
    .B1(_03609_));
 sg13g2_nand3_1 _36095_ (.B(_03622_),
    .C(_05463_),
    .A(_03609_),
    .Y(_05507_));
 sg13g2_nor2b_1 _36096_ (.A(_05506_),
    .B_N(_05507_),
    .Y(_05508_));
 sg13g2_a21oi_1 _36097_ (.A1(net7322),
    .A2(_05508_),
    .Y(_05509_),
    .B1(net6289));
 sg13g2_o21ai_1 _36098_ (.B1(_05509_),
    .Y(_05510_),
    .A1(net7322),
    .A2(_18105_));
 sg13g2_o21ai_1 _36099_ (.B1(_05510_),
    .Y(_05511_),
    .A1(net6209),
    .A2(_05505_));
 sg13g2_nand2b_1 _36100_ (.Y(_05512_),
    .B(net5782),
    .A_N(_05511_));
 sg13g2_xnor2_1 _36101_ (.Y(_05513_),
    .A(net5782),
    .B(_05511_));
 sg13g2_xnor2_1 _36102_ (.Y(_05514_),
    .A(net5837),
    .B(_05511_));
 sg13g2_a21oi_1 _36103_ (.A1(\u_inv.d_next[242] ),
    .A2(\u_inv.d_reg[242] ),
    .Y(_05515_),
    .B1(_05506_));
 sg13g2_xnor2_1 _36104_ (.Y(_05516_),
    .A(_03607_),
    .B(_05515_));
 sg13g2_a21o_1 _36105_ (.A2(\u_inv.d_next[243] ),
    .A1(net7188),
    .B1(net6289),
    .X(_05517_));
 sg13g2_a21oi_1 _36106_ (.A1(net7322),
    .A2(_05516_),
    .Y(_05518_),
    .B1(_05517_));
 sg13g2_a21oi_1 _36107_ (.A1(_03609_),
    .A2(_05504_),
    .Y(_05519_),
    .B1(_04748_));
 sg13g2_nand2b_1 _36108_ (.Y(_05520_),
    .B(_03607_),
    .A_N(_05519_));
 sg13g2_a21oi_1 _36109_ (.A1(_03608_),
    .A2(_05519_),
    .Y(_05521_),
    .B1(net6209));
 sg13g2_a21o_2 _36110_ (.A2(_05521_),
    .A1(_05520_),
    .B1(_05518_),
    .X(_05522_));
 sg13g2_xnor2_1 _36111_ (.Y(_05523_),
    .A(net5837),
    .B(_05522_));
 sg13g2_nor2_2 _36112_ (.A(_05514_),
    .B(_05523_),
    .Y(_05524_));
 sg13g2_a21oi_1 _36113_ (.A1(_03615_),
    .A2(_05357_),
    .Y(_05525_),
    .B1(_04749_));
 sg13g2_o21ai_1 _36114_ (.B1(net6289),
    .Y(_05526_),
    .A1(_03599_),
    .A2(_05525_));
 sg13g2_a21oi_1 _36115_ (.A1(_03599_),
    .A2(_05525_),
    .Y(_05527_),
    .B1(_05526_));
 sg13g2_a21oi_1 _36116_ (.A1(_03598_),
    .A2(_05462_),
    .Y(_05528_),
    .B1(net7188));
 sg13g2_o21ai_1 _36117_ (.B1(_05528_),
    .Y(_05529_),
    .A1(_03598_),
    .A2(_05462_));
 sg13g2_a21oi_1 _36118_ (.A1(net7187),
    .A2(\u_inv.d_next[241] ),
    .Y(_05530_),
    .B1(net6288));
 sg13g2_a21oi_1 _36119_ (.A1(_05529_),
    .A2(_05530_),
    .Y(_05531_),
    .B1(_05527_));
 sg13g2_nand2_1 _36120_ (.Y(_05532_),
    .A(net5777),
    .B(_05531_));
 sg13g2_xnor2_1 _36121_ (.Y(_05533_),
    .A(net5777),
    .B(_05531_));
 sg13g2_nor2_1 _36122_ (.A(net7187),
    .B(_05367_),
    .Y(_05534_));
 sg13g2_o21ai_1 _36123_ (.B1(_05534_),
    .Y(_05535_),
    .A1(_03614_),
    .A2(_05366_));
 sg13g2_xnor2_1 _36124_ (.Y(_05536_),
    .A(_03615_),
    .B(_05357_));
 sg13g2_a21oi_1 _36125_ (.A1(net7188),
    .A2(\u_inv.d_next[240] ),
    .Y(_05537_),
    .B1(net6288));
 sg13g2_a22oi_1 _36126_ (.Y(_05538_),
    .B1(_05537_),
    .B2(_05535_),
    .A2(_05536_),
    .A1(net6288));
 sg13g2_nand2_1 _36127_ (.Y(_05539_),
    .A(net5777),
    .B(_05538_));
 sg13g2_xnor2_1 _36128_ (.Y(_05540_),
    .A(net5837),
    .B(_05538_));
 sg13g2_nor2b_1 _36129_ (.A(_05533_),
    .B_N(_05540_),
    .Y(_05541_));
 sg13g2_inv_1 _36130_ (.Y(_05542_),
    .A(_05541_));
 sg13g2_and3_1 _36131_ (.X(_05543_),
    .A(_05503_),
    .B(_05524_),
    .C(_05541_));
 sg13g2_a21oi_2 _36132_ (.B1(_04730_),
    .Y(_05544_),
    .A2(_05356_),
    .A1(_04618_));
 sg13g2_o21ai_1 _36133_ (.B1(_04742_),
    .Y(_05545_),
    .A1(_04611_),
    .A2(_05544_));
 sg13g2_a21oi_1 _36134_ (.A1(_04607_),
    .A2(_05545_),
    .Y(_05546_),
    .B1(_04733_));
 sg13g2_xnor2_1 _36135_ (.Y(_05547_),
    .A(_03514_),
    .B(_05546_));
 sg13g2_nor2_1 _36136_ (.A(_03558_),
    .B(_05365_),
    .Y(_05548_));
 sg13g2_o21ai_1 _36137_ (.B1(_03644_),
    .Y(_05549_),
    .A1(_03563_),
    .A2(_05365_));
 sg13g2_a21oi_1 _36138_ (.A1(_03530_),
    .A2(_05549_),
    .Y(_05550_),
    .B1(_03647_));
 sg13g2_a21o_1 _36139_ (.A2(_05549_),
    .A1(_03530_),
    .B1(_03647_),
    .X(_05551_));
 sg13g2_a21o_2 _36140_ (.A2(_05551_),
    .A1(_03537_),
    .B1(_03648_),
    .X(_05552_));
 sg13g2_a21oi_1 _36141_ (.A1(_03521_),
    .A2(_05552_),
    .Y(_05553_),
    .B1(_03645_));
 sg13g2_nand2b_1 _36142_ (.Y(_05554_),
    .B(_03514_),
    .A_N(_05553_));
 sg13g2_xnor2_1 _36143_ (.Y(_05555_),
    .A(_03514_),
    .B(_05553_));
 sg13g2_nand2_1 _36144_ (.Y(_05556_),
    .A(net7191),
    .B(\u_inv.d_next[238] ));
 sg13g2_a21oi_1 _36145_ (.A1(net7321),
    .A2(_05555_),
    .Y(_05557_),
    .B1(net6293));
 sg13g2_a22oi_1 _36146_ (.Y(_05558_),
    .B1(_05556_),
    .B2(_05557_),
    .A2(_05547_),
    .A1(net6293));
 sg13g2_nand2_1 _36147_ (.Y(_05559_),
    .A(net5777),
    .B(_05558_));
 sg13g2_xnor2_1 _36148_ (.Y(_05560_),
    .A(net5777),
    .B(_05558_));
 sg13g2_nand3_1 _36149_ (.B(_03513_),
    .C(_05554_),
    .A(_03512_),
    .Y(_05561_));
 sg13g2_a21o_1 _36150_ (.A2(_05554_),
    .A1(_03513_),
    .B1(_03512_),
    .X(_05562_));
 sg13g2_nand3_1 _36151_ (.B(_05561_),
    .C(_05562_),
    .A(net7321),
    .Y(_05563_));
 sg13g2_a21oi_1 _36152_ (.A1(net7191),
    .A2(\u_inv.d_next[239] ),
    .Y(_05564_),
    .B1(net6292));
 sg13g2_o21ai_1 _36153_ (.B1(_04735_),
    .Y(_05565_),
    .A1(_03514_),
    .A2(_05546_));
 sg13g2_nand2b_1 _36154_ (.Y(_05566_),
    .B(_03512_),
    .A_N(_05565_));
 sg13g2_a21oi_1 _36155_ (.A1(_03511_),
    .A2(_05565_),
    .Y(_05567_),
    .B1(net6210));
 sg13g2_a22oi_1 _36156_ (.Y(_05568_),
    .B1(_05566_),
    .B2(_05567_),
    .A2(_05564_),
    .A1(_05563_));
 sg13g2_xnor2_1 _36157_ (.Y(_05569_),
    .A(net5777),
    .B(_05568_));
 sg13g2_nor2_1 _36158_ (.A(_05560_),
    .B(_05569_),
    .Y(_05570_));
 sg13g2_xnor2_1 _36159_ (.Y(_05571_),
    .A(_03520_),
    .B(_05545_));
 sg13g2_nand2b_1 _36160_ (.Y(_05572_),
    .B(_05552_),
    .A_N(_03520_));
 sg13g2_xnor2_1 _36161_ (.Y(_05573_),
    .A(_03520_),
    .B(_05552_));
 sg13g2_nand2_1 _36162_ (.Y(_05574_),
    .A(net7191),
    .B(\u_inv.d_next[236] ));
 sg13g2_a21oi_1 _36163_ (.A1(net7321),
    .A2(_05573_),
    .Y(_05575_),
    .B1(net6292));
 sg13g2_a22oi_1 _36164_ (.Y(_05576_),
    .B1(_05574_),
    .B2(_05575_),
    .A2(_05571_),
    .A1(net6292));
 sg13g2_nand2_1 _36165_ (.Y(_05577_),
    .A(net5777),
    .B(_05576_));
 sg13g2_inv_1 _36166_ (.Y(_05578_),
    .A(_05577_));
 sg13g2_xnor2_1 _36167_ (.Y(_05579_),
    .A(net5778),
    .B(_05576_));
 sg13g2_inv_1 _36168_ (.Y(_05580_),
    .A(_05579_));
 sg13g2_a21o_1 _36169_ (.A2(_05572_),
    .A1(_03519_),
    .B1(_03518_),
    .X(_05581_));
 sg13g2_nand3_1 _36170_ (.B(_03519_),
    .C(_05572_),
    .A(_03518_),
    .Y(_05582_));
 sg13g2_nand3_1 _36171_ (.B(_05581_),
    .C(_05582_),
    .A(net7321),
    .Y(_05583_));
 sg13g2_a21oi_1 _36172_ (.A1(net7190),
    .A2(\u_inv.d_next[237] ),
    .Y(_05584_),
    .B1(net6292));
 sg13g2_a21oi_1 _36173_ (.A1(_03520_),
    .A2(_05545_),
    .Y(_05585_),
    .B1(_04731_));
 sg13g2_or2_1 _36174_ (.X(_05586_),
    .B(_05585_),
    .A(_03518_));
 sg13g2_a21oi_1 _36175_ (.A1(_03518_),
    .A2(_05585_),
    .Y(_05587_),
    .B1(net6210));
 sg13g2_a22oi_1 _36176_ (.Y(_05588_),
    .B1(_05586_),
    .B2(_05587_),
    .A2(_05584_),
    .A1(_05583_));
 sg13g2_xnor2_1 _36177_ (.Y(_05589_),
    .A(net5778),
    .B(_05588_));
 sg13g2_or2_1 _36178_ (.X(_05590_),
    .B(_05589_),
    .A(_05579_));
 sg13g2_inv_1 _36179_ (.Y(_05591_),
    .A(_05590_));
 sg13g2_nor3_1 _36180_ (.A(_05560_),
    .B(_05569_),
    .C(_05590_),
    .Y(_05592_));
 sg13g2_nand2_1 _36181_ (.Y(_05593_),
    .A(_03528_),
    .B(_05549_));
 sg13g2_xnor2_1 _36182_ (.Y(_05594_),
    .A(_03528_),
    .B(_05549_));
 sg13g2_o21ai_1 _36183_ (.B1(net6210),
    .Y(_05595_),
    .A1(net7320),
    .A2(\u_inv.d_next[232] ));
 sg13g2_a21oi_1 _36184_ (.A1(net7321),
    .A2(_05594_),
    .Y(_05596_),
    .B1(_05595_));
 sg13g2_xnor2_1 _36185_ (.Y(_05597_),
    .A(_03529_),
    .B(_05544_));
 sg13g2_a21oi_2 _36186_ (.B1(_05596_),
    .Y(_05598_),
    .A2(_05597_),
    .A1(net6290));
 sg13g2_or2_1 _36187_ (.X(_05599_),
    .B(_05598_),
    .A(net5837));
 sg13g2_xnor2_1 _36188_ (.Y(_05600_),
    .A(net5781),
    .B(_05598_));
 sg13g2_o21ai_1 _36189_ (.B1(_04738_),
    .Y(_05601_),
    .A1(_03528_),
    .A2(_05544_));
 sg13g2_o21ai_1 _36190_ (.B1(net6291),
    .Y(_05602_),
    .A1(_03525_),
    .A2(_05601_));
 sg13g2_a21oi_1 _36191_ (.A1(_03525_),
    .A2(_05601_),
    .Y(_05603_),
    .B1(_05602_));
 sg13g2_nand2_1 _36192_ (.Y(_05604_),
    .A(_03527_),
    .B(_05593_));
 sg13g2_a21oi_1 _36193_ (.A1(_03525_),
    .A2(_05604_),
    .Y(_05605_),
    .B1(net7190));
 sg13g2_o21ai_1 _36194_ (.B1(_05605_),
    .Y(_05606_),
    .A1(_03525_),
    .A2(_05604_));
 sg13g2_a21oi_1 _36195_ (.A1(net7190),
    .A2(\u_inv.d_next[233] ),
    .Y(_05607_),
    .B1(net6290));
 sg13g2_a21oi_1 _36196_ (.A1(_05606_),
    .A2(_05607_),
    .Y(_05608_),
    .B1(_05603_));
 sg13g2_nand2_1 _36197_ (.Y(_05609_),
    .A(net5778),
    .B(_05608_));
 sg13g2_xnor2_1 _36198_ (.Y(_05610_),
    .A(net5837),
    .B(_05608_));
 sg13g2_and2_1 _36199_ (.A(_05600_),
    .B(_05610_),
    .X(_05611_));
 sg13g2_a21oi_1 _36200_ (.A1(_03536_),
    .A2(_05550_),
    .Y(_05612_),
    .B1(net7190));
 sg13g2_o21ai_1 _36201_ (.B1(_05612_),
    .Y(_05613_),
    .A1(_03536_),
    .A2(_05550_));
 sg13g2_o21ai_1 _36202_ (.B1(_04741_),
    .Y(_05614_),
    .A1(_04610_),
    .A2(_05544_));
 sg13g2_xnor2_1 _36203_ (.Y(_05615_),
    .A(_03536_),
    .B(_05614_));
 sg13g2_a21oi_1 _36204_ (.A1(net7190),
    .A2(\u_inv.d_next[234] ),
    .Y(_05616_),
    .B1(net6292));
 sg13g2_a22oi_1 _36205_ (.Y(_05617_),
    .B1(_05616_),
    .B2(_05613_),
    .A2(_05615_),
    .A1(net6292));
 sg13g2_nand2_1 _36206_ (.Y(_05618_),
    .A(net5778),
    .B(_05617_));
 sg13g2_xnor2_1 _36207_ (.Y(_05619_),
    .A(net5778),
    .B(_05617_));
 sg13g2_a21oi_1 _36208_ (.A1(_03536_),
    .A2(_05614_),
    .Y(_05620_),
    .B1(_04737_));
 sg13g2_nand2b_1 _36209_ (.Y(_05621_),
    .B(_03533_),
    .A_N(_05620_));
 sg13g2_a21oi_1 _36210_ (.A1(_03534_),
    .A2(_05620_),
    .Y(_05622_),
    .B1(net6210));
 sg13g2_o21ai_1 _36211_ (.B1(_03535_),
    .Y(_05623_),
    .A1(_03536_),
    .A2(_05550_));
 sg13g2_a21oi_1 _36212_ (.A1(_03533_),
    .A2(_05623_),
    .Y(_05624_),
    .B1(net7190));
 sg13g2_o21ai_1 _36213_ (.B1(_05624_),
    .Y(_05625_),
    .A1(_03533_),
    .A2(_05623_));
 sg13g2_a21oi_1 _36214_ (.A1(net7190),
    .A2(\u_inv.d_next[235] ),
    .Y(_05626_),
    .B1(net6292));
 sg13g2_a22oi_1 _36215_ (.Y(_05627_),
    .B1(_05625_),
    .B2(_05626_),
    .A2(_05622_),
    .A1(_05621_));
 sg13g2_xnor2_1 _36216_ (.Y(_05628_),
    .A(net5778),
    .B(_05627_));
 sg13g2_or2_1 _36217_ (.X(_05629_),
    .B(_05628_),
    .A(_05619_));
 sg13g2_inv_1 _36218_ (.Y(_05630_),
    .A(_05629_));
 sg13g2_a21oi_1 _36219_ (.A1(\u_inv.d_next[224] ),
    .A2(\u_inv.d_reg[224] ),
    .Y(_05631_),
    .B1(_05548_));
 sg13g2_o21ai_1 _36220_ (.B1(_03637_),
    .Y(_05632_),
    .A1(_03562_),
    .A2(_05365_));
 sg13g2_a21o_1 _36221_ (.A2(_05632_),
    .A1(_03542_),
    .B1(_03639_),
    .X(_05633_));
 sg13g2_a21oi_1 _36222_ (.A1(_03550_),
    .A2(_05633_),
    .Y(_05634_),
    .B1(_03641_));
 sg13g2_or2_1 _36223_ (.X(_05635_),
    .B(_05634_),
    .A(_03552_));
 sg13g2_nand3_1 _36224_ (.B(_03555_),
    .C(_05635_),
    .A(_03551_),
    .Y(_05636_));
 sg13g2_a21o_1 _36225_ (.A2(_05635_),
    .A1(_03551_),
    .B1(_03555_),
    .X(_05637_));
 sg13g2_nand3_1 _36226_ (.B(_05636_),
    .C(_05637_),
    .A(net7320),
    .Y(_05638_));
 sg13g2_nand2_1 _36227_ (.Y(_05639_),
    .A(net7189),
    .B(\u_inv.d_next[231] ));
 sg13g2_nand3_1 _36228_ (.B(_05638_),
    .C(_05639_),
    .A(net6209),
    .Y(_05640_));
 sg13g2_nand3_1 _36229_ (.B(_04616_),
    .C(_05356_),
    .A(_04615_),
    .Y(_05641_));
 sg13g2_a21oi_1 _36230_ (.A1(_04721_),
    .A2(_05641_),
    .Y(_05642_),
    .B1(_04613_));
 sg13g2_nor2_1 _36231_ (.A(_04726_),
    .B(_05642_),
    .Y(_05643_));
 sg13g2_o21ai_1 _36232_ (.B1(_03552_),
    .Y(_05644_),
    .A1(_04726_),
    .A2(_05642_));
 sg13g2_a21o_1 _36233_ (.A2(_05644_),
    .A1(_04723_),
    .B1(_03555_),
    .X(_05645_));
 sg13g2_nand3_1 _36234_ (.B(_04723_),
    .C(_05644_),
    .A(_03555_),
    .Y(_05646_));
 sg13g2_nand3_1 _36235_ (.B(_05645_),
    .C(_05646_),
    .A(net6290),
    .Y(_05647_));
 sg13g2_and3_2 _36236_ (.X(_05648_),
    .A(net5779),
    .B(_05640_),
    .C(_05647_));
 sg13g2_a21oi_1 _36237_ (.A1(_05640_),
    .A2(_05647_),
    .Y(_05649_),
    .B1(net5779));
 sg13g2_or2_1 _36238_ (.X(_05650_),
    .B(_05649_),
    .A(_05648_));
 sg13g2_xor2_1 _36239_ (.B(_05643_),
    .A(_03552_),
    .X(_05651_));
 sg13g2_nand2_1 _36240_ (.Y(_05652_),
    .A(_03552_),
    .B(_05634_));
 sg13g2_nand3_1 _36241_ (.B(_05635_),
    .C(_05652_),
    .A(net7320),
    .Y(_05653_));
 sg13g2_a21oi_1 _36242_ (.A1(net7189),
    .A2(\u_inv.d_next[230] ),
    .Y(_05654_),
    .B1(net6290));
 sg13g2_a22oi_1 _36243_ (.Y(_05655_),
    .B1(_05653_),
    .B2(_05654_),
    .A2(_05651_),
    .A1(net6290));
 sg13g2_and2_1 _36244_ (.A(net5779),
    .B(_05655_),
    .X(_05656_));
 sg13g2_xnor2_1 _36245_ (.Y(_05657_),
    .A(net5779),
    .B(_05655_));
 sg13g2_nor3_1 _36246_ (.A(_05648_),
    .B(_05649_),
    .C(_05657_),
    .Y(_05658_));
 sg13g2_a21oi_1 _36247_ (.A1(_04721_),
    .A2(_05641_),
    .Y(_05659_),
    .B1(_03548_));
 sg13g2_nand3_1 _36248_ (.B(_04721_),
    .C(_05641_),
    .A(_03548_),
    .Y(_05660_));
 sg13g2_nand2b_1 _36249_ (.Y(_05661_),
    .B(_05660_),
    .A_N(_05659_));
 sg13g2_nand2_1 _36250_ (.Y(_05662_),
    .A(_03548_),
    .B(_05633_));
 sg13g2_o21ai_1 _36251_ (.B1(net7320),
    .Y(_05663_),
    .A1(_03548_),
    .A2(_05633_));
 sg13g2_nand2b_1 _36252_ (.Y(_05664_),
    .B(_05662_),
    .A_N(_05663_));
 sg13g2_a21oi_1 _36253_ (.A1(net7189),
    .A2(\u_inv.d_next[228] ),
    .Y(_05665_),
    .B1(net6290));
 sg13g2_a22oi_1 _36254_ (.Y(_05666_),
    .B1(_05664_),
    .B2(_05665_),
    .A2(_05661_),
    .A1(net6290));
 sg13g2_nand2_1 _36255_ (.Y(_05667_),
    .A(net5780),
    .B(_05666_));
 sg13g2_xnor2_1 _36256_ (.Y(_05668_),
    .A(net5837),
    .B(_05666_));
 sg13g2_inv_1 _36257_ (.Y(_05669_),
    .A(_05668_));
 sg13g2_a21oi_1 _36258_ (.A1(_03547_),
    .A2(_05662_),
    .Y(_05670_),
    .B1(_03546_));
 sg13g2_nand3_1 _36259_ (.B(_03547_),
    .C(_05662_),
    .A(_03546_),
    .Y(_05671_));
 sg13g2_nand2_1 _36260_ (.Y(_05672_),
    .A(net7320),
    .B(_05671_));
 sg13g2_a21oi_1 _36261_ (.A1(net7191),
    .A2(\u_inv.d_next[229] ),
    .Y(_05673_),
    .B1(net6291));
 sg13g2_o21ai_1 _36262_ (.B1(_05673_),
    .Y(_05674_),
    .A1(_05670_),
    .A2(_05672_));
 sg13g2_o21ai_1 _36263_ (.B1(_03545_),
    .Y(_05675_),
    .A1(_04724_),
    .A2(_05659_));
 sg13g2_or3_1 _36264_ (.A(_03545_),
    .B(_04724_),
    .C(_05659_),
    .X(_05676_));
 sg13g2_nand3_1 _36265_ (.B(_05675_),
    .C(_05676_),
    .A(net6290),
    .Y(_05677_));
 sg13g2_a21o_1 _36266_ (.A2(_05677_),
    .A1(_05674_),
    .B1(net5780),
    .X(_05678_));
 sg13g2_nand3_1 _36267_ (.B(_05674_),
    .C(_05677_),
    .A(net5780),
    .Y(_05679_));
 sg13g2_and2_1 _36268_ (.A(_05678_),
    .B(_05679_),
    .X(_05680_));
 sg13g2_nand3_1 _36269_ (.B(_05678_),
    .C(_05679_),
    .A(_05668_),
    .Y(_05681_));
 sg13g2_nor4_1 _36270_ (.A(_05648_),
    .B(_05649_),
    .C(_05657_),
    .D(_05681_),
    .Y(_05682_));
 sg13g2_a21oi_1 _36271_ (.A1(_04616_),
    .A2(_05356_),
    .Y(_05683_),
    .B1(_04719_));
 sg13g2_xnor2_1 _36272_ (.Y(_05684_),
    .A(_03541_),
    .B(_05683_));
 sg13g2_o21ai_1 _36273_ (.B1(net7320),
    .Y(_05685_),
    .A1(_03541_),
    .A2(_05632_));
 sg13g2_a21o_1 _36274_ (.A2(_05632_),
    .A1(_03541_),
    .B1(_05685_),
    .X(_05686_));
 sg13g2_a21oi_1 _36275_ (.A1(net7189),
    .A2(\u_inv.d_next[226] ),
    .Y(_05687_),
    .B1(net6291));
 sg13g2_a22oi_1 _36276_ (.Y(_05688_),
    .B1(_05686_),
    .B2(_05687_),
    .A2(_05684_),
    .A1(net6291));
 sg13g2_nand2_1 _36277_ (.Y(_05689_),
    .A(net5779),
    .B(_05688_));
 sg13g2_xnor2_1 _36278_ (.Y(_05690_),
    .A(net5838),
    .B(_05688_));
 sg13g2_inv_1 _36279_ (.Y(_05691_),
    .A(_05690_));
 sg13g2_a21oi_1 _36280_ (.A1(_03541_),
    .A2(_05632_),
    .Y(_05692_),
    .B1(_03540_));
 sg13g2_xnor2_1 _36281_ (.Y(_05693_),
    .A(_03539_),
    .B(_05692_));
 sg13g2_nand2_1 _36282_ (.Y(_05694_),
    .A(net7320),
    .B(_05693_));
 sg13g2_a21oi_1 _36283_ (.A1(net7189),
    .A2(\u_inv.d_next[227] ),
    .Y(_05695_),
    .B1(net6281));
 sg13g2_o21ai_1 _36284_ (.B1(_04716_),
    .Y(_05696_),
    .A1(_03541_),
    .A2(_05683_));
 sg13g2_or2_1 _36285_ (.X(_05697_),
    .B(_05696_),
    .A(_03539_));
 sg13g2_a21oi_1 _36286_ (.A1(_03539_),
    .A2(_05696_),
    .Y(_05698_),
    .B1(net6209));
 sg13g2_a22oi_1 _36287_ (.Y(_05699_),
    .B1(_05697_),
    .B2(_05698_),
    .A2(_05695_),
    .A1(_05694_));
 sg13g2_xnor2_1 _36288_ (.Y(_05700_),
    .A(net5838),
    .B(_05699_));
 sg13g2_and2_1 _36289_ (.A(_05690_),
    .B(_05700_),
    .X(_05701_));
 sg13g2_a21oi_1 _36290_ (.A1(_03560_),
    .A2(_05631_),
    .Y(_05702_),
    .B1(net7189));
 sg13g2_o21ai_1 _36291_ (.B1(_05702_),
    .Y(_05703_),
    .A1(_03560_),
    .A2(_05631_));
 sg13g2_a21oi_1 _36292_ (.A1(net7189),
    .A2(\u_inv.d_next[225] ),
    .Y(_05704_),
    .B1(net6281));
 sg13g2_a21oi_1 _36293_ (.A1(_03558_),
    .A2(_05356_),
    .Y(_05705_),
    .B1(_04717_));
 sg13g2_or2_1 _36294_ (.X(_05706_),
    .B(_05705_),
    .A(_03560_));
 sg13g2_a21oi_1 _36295_ (.A1(_03560_),
    .A2(_05705_),
    .Y(_05707_),
    .B1(net6210));
 sg13g2_a22oi_1 _36296_ (.Y(_05708_),
    .B1(_05706_),
    .B2(_05707_),
    .A2(_05704_),
    .A1(_05703_));
 sg13g2_nand2_1 _36297_ (.Y(_05709_),
    .A(net5779),
    .B(_05708_));
 sg13g2_xnor2_1 _36298_ (.Y(_05710_),
    .A(net5779),
    .B(_05708_));
 sg13g2_nand2_1 _36299_ (.Y(_05711_),
    .A(_03558_),
    .B(_05365_));
 sg13g2_nand3b_1 _36300_ (.B(_05711_),
    .C(net7320),
    .Y(_05712_),
    .A_N(_05548_));
 sg13g2_xnor2_1 _36301_ (.Y(_05713_),
    .A(_03558_),
    .B(_05356_));
 sg13g2_a21oi_1 _36302_ (.A1(net7189),
    .A2(\u_inv.d_next[224] ),
    .Y(_05714_),
    .B1(net6281));
 sg13g2_a22oi_1 _36303_ (.Y(_05715_),
    .B1(_05714_),
    .B2(_05712_),
    .A2(_05713_),
    .A1(net6291));
 sg13g2_nand2_1 _36304_ (.Y(_05716_),
    .A(net5779),
    .B(_05715_));
 sg13g2_xnor2_1 _36305_ (.Y(_05717_),
    .A(net5837),
    .B(_05715_));
 sg13g2_nor2b_1 _36306_ (.A(_05710_),
    .B_N(_05717_),
    .Y(_05718_));
 sg13g2_inv_1 _36307_ (.Y(_05719_),
    .A(_05718_));
 sg13g2_and3_2 _36308_ (.X(_05720_),
    .A(_05682_),
    .B(_05701_),
    .C(_05718_));
 sg13g2_and4_1 _36309_ (.A(_05592_),
    .B(_05611_),
    .C(_05630_),
    .D(_05720_),
    .X(_05721_));
 sg13g2_nand4_1 _36310_ (.B(_05455_),
    .C(_05543_),
    .A(_05415_),
    .Y(_05722_),
    .D(_05721_));
 sg13g2_o21ai_1 _36311_ (.B1(_04684_),
    .Y(_05723_),
    .A1(_04651_),
    .A2(_05353_));
 sg13g2_a21oi_2 _36312_ (.B1(_04698_),
    .Y(_05724_),
    .A2(_05723_),
    .A1(_04634_));
 sg13g2_a21o_1 _36313_ (.A2(_05723_),
    .A1(_04634_),
    .B1(_04698_),
    .X(_05725_));
 sg13g2_o21ai_1 _36314_ (.B1(_04711_),
    .Y(_05726_),
    .A1(_04625_),
    .A2(_05724_));
 sg13g2_a221oi_1 _36315_ (.B2(_04621_),
    .C1(_04702_),
    .B1(_05726_),
    .A1(_03432_),
    .Y(_05727_),
    .A2(_04701_));
 sg13g2_xnor2_1 _36316_ (.Y(_05728_),
    .A(_03440_),
    .B(_05727_));
 sg13g2_nand2_1 _36317_ (.Y(_05729_),
    .A(net1080),
    .B(_04584_));
 sg13g2_nand3b_1 _36318_ (.B(net1081),
    .C(_04585_),
    .Y(_05730_),
    .A_N(_03428_));
 sg13g2_a21oi_1 _36319_ (.A1(_03431_),
    .A2(_05730_),
    .Y(_05731_),
    .B1(_03479_));
 sg13g2_o21ai_1 _36320_ (.B1(_03454_),
    .Y(_05732_),
    .A1(_03506_),
    .A2(_05731_));
 sg13g2_nand2_1 _36321_ (.Y(_05733_),
    .A(_03482_),
    .B(_05732_));
 sg13g2_a21oi_1 _36322_ (.A1(_03482_),
    .A2(_05732_),
    .Y(_05734_),
    .B1(_03448_));
 sg13g2_o21ai_1 _36323_ (.B1(_03436_),
    .Y(_05735_),
    .A1(_03486_),
    .A2(_05734_));
 sg13g2_nand3_1 _36324_ (.B(_03491_),
    .C(_05735_),
    .A(_03439_),
    .Y(_05736_));
 sg13g2_a21o_1 _36325_ (.A2(_05735_),
    .A1(_03491_),
    .B1(_03439_),
    .X(_05737_));
 sg13g2_nand3_1 _36326_ (.B(_05736_),
    .C(_05737_),
    .A(net7323),
    .Y(_05738_));
 sg13g2_a21oi_1 _36327_ (.A1(net7192),
    .A2(\u_inv.d_next[222] ),
    .Y(_05739_),
    .B1(net6294));
 sg13g2_a22oi_1 _36328_ (.Y(_05740_),
    .B1(_05738_),
    .B2(_05739_),
    .A2(_05728_),
    .A1(net6294));
 sg13g2_nand2_1 _36329_ (.Y(_05741_),
    .A(net5783),
    .B(_05740_));
 sg13g2_xnor2_1 _36330_ (.Y(_05742_),
    .A(net5783),
    .B(_05740_));
 sg13g2_a21o_1 _36331_ (.A2(_05737_),
    .A1(_03438_),
    .B1(_03437_),
    .X(_05743_));
 sg13g2_nand3_1 _36332_ (.B(_03438_),
    .C(_05737_),
    .A(_03437_),
    .Y(_05744_));
 sg13g2_nand3_1 _36333_ (.B(_05743_),
    .C(_05744_),
    .A(net7323),
    .Y(_05745_));
 sg13g2_a21oi_1 _36334_ (.A1(net7192),
    .A2(\u_inv.d_next[223] ),
    .Y(_05746_),
    .B1(net6295));
 sg13g2_o21ai_1 _36335_ (.B1(_04700_),
    .Y(_05747_),
    .A1(_03440_),
    .A2(_05727_));
 sg13g2_xnor2_1 _36336_ (.Y(_05748_),
    .A(_03437_),
    .B(_05747_));
 sg13g2_a22oi_1 _36337_ (.Y(_05749_),
    .B1(_05748_),
    .B2(net6294),
    .A2(_05746_),
    .A1(_05745_));
 sg13g2_xnor2_1 _36338_ (.Y(_05750_),
    .A(net5838),
    .B(_05749_));
 sg13g2_xnor2_1 _36339_ (.Y(_05751_),
    .A(net5783),
    .B(_05749_));
 sg13g2_nor2_1 _36340_ (.A(_05742_),
    .B(_05751_),
    .Y(_05752_));
 sg13g2_o21ai_1 _36341_ (.B1(_03435_),
    .Y(_05753_),
    .A1(_03486_),
    .A2(_05734_));
 sg13g2_a21o_1 _36342_ (.A2(_05753_),
    .A1(_03433_),
    .B1(_03432_),
    .X(_05754_));
 sg13g2_nand3_1 _36343_ (.B(_03433_),
    .C(_05753_),
    .A(_03432_),
    .Y(_05755_));
 sg13g2_nand3_1 _36344_ (.B(_05754_),
    .C(_05755_),
    .A(net7323),
    .Y(_05756_));
 sg13g2_a21oi_1 _36345_ (.A1(net7192),
    .A2(\u_inv.d_next[221] ),
    .Y(_05757_),
    .B1(net6294));
 sg13g2_a21oi_1 _36346_ (.A1(_03434_),
    .A2(_05726_),
    .Y(_05758_),
    .B1(_04701_));
 sg13g2_xor2_1 _36347_ (.B(_05758_),
    .A(_03432_),
    .X(_05759_));
 sg13g2_a22oi_1 _36348_ (.Y(_05760_),
    .B1(_05759_),
    .B2(net6294),
    .A2(_05757_),
    .A1(_05756_));
 sg13g2_nand2_1 _36349_ (.Y(_05761_),
    .A(net5785),
    .B(_05760_));
 sg13g2_xnor2_1 _36350_ (.Y(_05762_),
    .A(net5785),
    .B(_05760_));
 sg13g2_xnor2_1 _36351_ (.Y(_05763_),
    .A(_03434_),
    .B(_05726_));
 sg13g2_or3_1 _36352_ (.A(_03435_),
    .B(_03486_),
    .C(_05734_),
    .X(_05764_));
 sg13g2_nand3_1 _36353_ (.B(_05753_),
    .C(_05764_),
    .A(net7323),
    .Y(_05765_));
 sg13g2_a21oi_1 _36354_ (.A1(net7192),
    .A2(\u_inv.d_next[220] ),
    .Y(_05766_),
    .B1(net6294));
 sg13g2_a22oi_1 _36355_ (.Y(_05767_),
    .B1(_05765_),
    .B2(_05766_),
    .A2(_05763_),
    .A1(net6294));
 sg13g2_nand2_1 _36356_ (.Y(_05768_),
    .A(net5783),
    .B(_05767_));
 sg13g2_xnor2_1 _36357_ (.Y(_05769_),
    .A(net5783),
    .B(_05767_));
 sg13g2_nor2_1 _36358_ (.A(_05762_),
    .B(_05769_),
    .Y(_05770_));
 sg13g2_nor4_1 _36359_ (.A(_05742_),
    .B(_05751_),
    .C(_05762_),
    .D(_05769_),
    .Y(_05771_));
 sg13g2_nand3b_1 _36360_ (.B(_05750_),
    .C(_05770_),
    .Y(_05772_),
    .A_N(_05742_));
 sg13g2_a21oi_1 _36361_ (.A1(_03447_),
    .A2(_05733_),
    .Y(_05773_),
    .B1(_03484_));
 sg13g2_a21oi_1 _36362_ (.A1(_03445_),
    .A2(_05773_),
    .Y(_05774_),
    .B1(net7192));
 sg13g2_o21ai_1 _36363_ (.B1(_05774_),
    .Y(_05775_),
    .A1(_03445_),
    .A2(_05773_));
 sg13g2_a21oi_1 _36364_ (.A1(net7193),
    .A2(\u_inv.d_next[219] ),
    .Y(_05776_),
    .B1(net6294));
 sg13g2_a21oi_1 _36365_ (.A1(_04624_),
    .A2(_05725_),
    .Y(_05777_),
    .B1(_04709_));
 sg13g2_o21ai_1 _36366_ (.B1(_03446_),
    .Y(_05778_),
    .A1(_03447_),
    .A2(_05777_));
 sg13g2_nand2b_1 _36367_ (.Y(_05779_),
    .B(_03445_),
    .A_N(_05778_));
 sg13g2_a21oi_1 _36368_ (.A1(_03444_),
    .A2(_05778_),
    .Y(_05780_),
    .B1(net6211));
 sg13g2_a22oi_1 _36369_ (.Y(_05781_),
    .B1(_05779_),
    .B2(_05780_),
    .A2(_05776_),
    .A1(_05775_));
 sg13g2_nand2_1 _36370_ (.Y(_05782_),
    .A(net5783),
    .B(_05781_));
 sg13g2_xnor2_1 _36371_ (.Y(_05783_),
    .A(net5838),
    .B(_05781_));
 sg13g2_o21ai_1 _36372_ (.B1(net6295),
    .Y(_05784_),
    .A1(_03447_),
    .A2(_05777_));
 sg13g2_a21oi_1 _36373_ (.A1(_03447_),
    .A2(_05777_),
    .Y(_05785_),
    .B1(_05784_));
 sg13g2_xnor2_1 _36374_ (.Y(_05786_),
    .A(_03447_),
    .B(_05733_));
 sg13g2_o21ai_1 _36375_ (.B1(net6211),
    .Y(_05787_),
    .A1(net7323),
    .A2(\u_inv.d_next[218] ));
 sg13g2_a21oi_1 _36376_ (.A1(net7323),
    .A2(_05786_),
    .Y(_05788_),
    .B1(_05787_));
 sg13g2_nor2_1 _36377_ (.A(_05785_),
    .B(_05788_),
    .Y(_05789_));
 sg13g2_o21ai_1 _36378_ (.B1(net5784),
    .Y(_05790_),
    .A1(_05785_),
    .A2(_05788_));
 sg13g2_xnor2_1 _36379_ (.Y(_05791_),
    .A(net5783),
    .B(_05789_));
 sg13g2_and2_1 _36380_ (.A(_05783_),
    .B(_05791_),
    .X(_05792_));
 sg13g2_nand2_1 _36381_ (.Y(_05793_),
    .A(_05783_),
    .B(_05791_));
 sg13g2_xnor2_1 _36382_ (.Y(_05794_),
    .A(_03452_),
    .B(_05724_));
 sg13g2_nor3_1 _36383_ (.A(_03452_),
    .B(_03506_),
    .C(_05731_),
    .Y(_05795_));
 sg13g2_o21ai_1 _36384_ (.B1(_03452_),
    .Y(_05796_),
    .A1(_03506_),
    .A2(_05731_));
 sg13g2_nand3b_1 _36385_ (.B(_05796_),
    .C(net7323),
    .Y(_05797_),
    .A_N(_05795_));
 sg13g2_a21oi_1 _36386_ (.A1(net7192),
    .A2(\u_inv.d_next[216] ),
    .Y(_05798_),
    .B1(net6295));
 sg13g2_a22oi_1 _36387_ (.Y(_05799_),
    .B1(_05797_),
    .B2(_05798_),
    .A2(_05794_),
    .A1(net6295));
 sg13g2_nand2_1 _36388_ (.Y(_05800_),
    .A(net5784),
    .B(_05799_));
 sg13g2_xnor2_1 _36389_ (.Y(_05801_),
    .A(net5838),
    .B(_05799_));
 sg13g2_nand2_1 _36390_ (.Y(_05802_),
    .A(_03451_),
    .B(_05796_));
 sg13g2_a21oi_1 _36391_ (.A1(_03449_),
    .A2(_05802_),
    .Y(_05803_),
    .B1(net7192));
 sg13g2_o21ai_1 _36392_ (.B1(_05803_),
    .Y(_05804_),
    .A1(_03449_),
    .A2(_05802_));
 sg13g2_a21oi_1 _36393_ (.A1(net7192),
    .A2(\u_inv.d_next[217] ),
    .Y(_05805_),
    .B1(net6295));
 sg13g2_o21ai_1 _36394_ (.B1(_04706_),
    .Y(_05806_),
    .A1(_03452_),
    .A2(_05724_));
 sg13g2_nand2b_1 _36395_ (.Y(_05807_),
    .B(_03450_),
    .A_N(_05806_));
 sg13g2_a21oi_1 _36396_ (.A1(_03449_),
    .A2(_05806_),
    .Y(_05808_),
    .B1(net6211));
 sg13g2_a22oi_1 _36397_ (.Y(_05809_),
    .B1(_05807_),
    .B2(_05808_),
    .A2(_05805_),
    .A1(_05804_));
 sg13g2_nand2_1 _36398_ (.Y(_05810_),
    .A(net5784),
    .B(_05809_));
 sg13g2_xnor2_1 _36399_ (.Y(_05811_),
    .A(net5785),
    .B(_05809_));
 sg13g2_inv_1 _36400_ (.Y(_05812_),
    .A(_05811_));
 sg13g2_nand2_1 _36401_ (.Y(_05813_),
    .A(_05801_),
    .B(_05812_));
 sg13g2_nand2_1 _36402_ (.Y(_05814_),
    .A(_04633_),
    .B(_05723_));
 sg13g2_nand2_1 _36403_ (.Y(_05815_),
    .A(_04687_),
    .B(_05814_));
 sg13g2_a21oi_1 _36404_ (.A1(_04633_),
    .A2(_05723_),
    .Y(_05816_),
    .B1(_04688_));
 sg13g2_nand3_1 _36405_ (.B(_04633_),
    .C(_05723_),
    .A(_04632_),
    .Y(_05817_));
 sg13g2_a21oi_1 _36406_ (.A1(_04691_),
    .A2(_05817_),
    .Y(_05818_),
    .B1(_04628_));
 sg13g2_o21ai_1 _36407_ (.B1(_03460_),
    .Y(_05819_),
    .A1(_04694_),
    .A2(_05818_));
 sg13g2_nor3_1 _36408_ (.A(_03460_),
    .B(_04694_),
    .C(_05818_),
    .Y(_05820_));
 sg13g2_nor2_1 _36409_ (.A(net6219),
    .B(_05820_),
    .Y(_05821_));
 sg13g2_a21oi_1 _36410_ (.A1(_03431_),
    .A2(_05730_),
    .Y(_05822_),
    .B1(_03476_));
 sg13g2_a21oi_1 _36411_ (.A1(_03431_),
    .A2(_05730_),
    .Y(_05823_),
    .B1(_03477_));
 sg13g2_nor2_1 _36412_ (.A(_03495_),
    .B(_05823_),
    .Y(_05824_));
 sg13g2_o21ai_1 _36413_ (.B1(_03471_),
    .Y(_05825_),
    .A1(_03495_),
    .A2(_05823_));
 sg13g2_nand2_1 _36414_ (.Y(_05826_),
    .A(_03498_),
    .B(_05825_));
 sg13g2_a21oi_1 _36415_ (.A1(_03498_),
    .A2(_05825_),
    .Y(_05827_),
    .B1(_03467_));
 sg13g2_nor3_1 _36416_ (.A(_03459_),
    .B(_03502_),
    .C(_05827_),
    .Y(_05828_));
 sg13g2_o21ai_1 _36417_ (.B1(_03459_),
    .Y(_05829_),
    .A1(_03502_),
    .A2(_05827_));
 sg13g2_nand2_1 _36418_ (.Y(_05830_),
    .A(net7334),
    .B(_05829_));
 sg13g2_nand2_1 _36419_ (.Y(_05831_),
    .A(net7198),
    .B(\u_inv.d_next[214] ));
 sg13g2_o21ai_1 _36420_ (.B1(_05831_),
    .Y(_05832_),
    .A1(_05828_),
    .A2(_05830_));
 sg13g2_a22oi_1 _36421_ (.Y(_05833_),
    .B1(_05832_),
    .B2(net6219),
    .A2(_05821_),
    .A1(_05819_));
 sg13g2_or2_1 _36422_ (.X(_05834_),
    .B(_05833_),
    .A(net5838));
 sg13g2_xnor2_1 _36423_ (.Y(_05835_),
    .A(net5838),
    .B(_05833_));
 sg13g2_inv_1 _36424_ (.Y(_05836_),
    .A(_05835_));
 sg13g2_a21o_1 _36425_ (.A2(_05829_),
    .A1(_03458_),
    .B1(_03457_),
    .X(_05837_));
 sg13g2_nand3_1 _36426_ (.B(_03458_),
    .C(_05829_),
    .A(_03457_),
    .Y(_05838_));
 sg13g2_nand3_1 _36427_ (.B(_05837_),
    .C(_05838_),
    .A(net7334),
    .Y(_05839_));
 sg13g2_nand2_1 _36428_ (.Y(_05840_),
    .A(net7198),
    .B(\u_inv.d_next[215] ));
 sg13g2_nand3_1 _36429_ (.B(_05839_),
    .C(_05840_),
    .A(net6219),
    .Y(_05841_));
 sg13g2_nand3_1 _36430_ (.B(_04695_),
    .C(_05819_),
    .A(_03457_),
    .Y(_05842_));
 sg13g2_a21o_1 _36431_ (.A2(_05819_),
    .A1(_04695_),
    .B1(_03457_),
    .X(_05843_));
 sg13g2_nand3_1 _36432_ (.B(_05842_),
    .C(_05843_),
    .A(net6303),
    .Y(_05844_));
 sg13g2_nand2_1 _36433_ (.Y(_05845_),
    .A(_05841_),
    .B(_05844_));
 sg13g2_a21oi_1 _36434_ (.A1(_05841_),
    .A2(_05844_),
    .Y(_05846_),
    .B1(net5784));
 sg13g2_and3_1 _36435_ (.X(_05847_),
    .A(net5784),
    .B(_05841_),
    .C(_05844_));
 sg13g2_nor2_1 _36436_ (.A(_05846_),
    .B(_05847_),
    .Y(_05848_));
 sg13g2_nor3_1 _36437_ (.A(_05835_),
    .B(_05846_),
    .C(_05847_),
    .Y(_05849_));
 sg13g2_a21oi_1 _36438_ (.A1(_03465_),
    .A2(_05826_),
    .Y(_05850_),
    .B1(_03464_));
 sg13g2_xnor2_1 _36439_ (.Y(_05851_),
    .A(_03463_),
    .B(_05850_));
 sg13g2_a21oi_1 _36440_ (.A1(net7198),
    .A2(\u_inv.d_next[213] ),
    .Y(_05852_),
    .B1(net6303));
 sg13g2_o21ai_1 _36441_ (.B1(_05852_),
    .Y(_05853_),
    .A1(net7198),
    .A2(_05851_));
 sg13g2_a21oi_1 _36442_ (.A1(_04691_),
    .A2(_05817_),
    .Y(_05854_),
    .B1(_03465_));
 sg13g2_o21ai_1 _36443_ (.B1(_03462_),
    .Y(_05855_),
    .A1(_04692_),
    .A2(_05854_));
 sg13g2_or3_1 _36444_ (.A(_03462_),
    .B(_04692_),
    .C(_05854_),
    .X(_05856_));
 sg13g2_nand3_1 _36445_ (.B(_05855_),
    .C(_05856_),
    .A(net6303),
    .Y(_05857_));
 sg13g2_nand2_1 _36446_ (.Y(_05858_),
    .A(_05853_),
    .B(_05857_));
 sg13g2_nand3_1 _36447_ (.B(_05853_),
    .C(_05857_),
    .A(net5787),
    .Y(_05859_));
 sg13g2_a21o_1 _36448_ (.A2(_05857_),
    .A1(_05853_),
    .B1(net5787),
    .X(_05860_));
 sg13g2_nand2_1 _36449_ (.Y(_05861_),
    .A(net5787),
    .B(_05858_));
 sg13g2_nand3_1 _36450_ (.B(_05853_),
    .C(_05857_),
    .A(net5840),
    .Y(_05862_));
 sg13g2_nand2_1 _36451_ (.Y(_05863_),
    .A(_05859_),
    .B(_05860_));
 sg13g2_nand3_1 _36452_ (.B(_04691_),
    .C(_05817_),
    .A(_03465_),
    .Y(_05864_));
 sg13g2_nor2_1 _36453_ (.A(net6219),
    .B(_05854_),
    .Y(_05865_));
 sg13g2_xnor2_1 _36454_ (.Y(_05866_),
    .A(_03465_),
    .B(_05826_));
 sg13g2_o21ai_1 _36455_ (.B1(net6219),
    .Y(_05867_),
    .A1(net7334),
    .A2(\u_inv.d_next[212] ));
 sg13g2_a21oi_1 _36456_ (.A1(net7334),
    .A2(_05866_),
    .Y(_05868_),
    .B1(_05867_));
 sg13g2_a21o_2 _36457_ (.A2(_05865_),
    .A1(_05864_),
    .B1(_05868_),
    .X(_05869_));
 sg13g2_nand2_1 _36458_ (.Y(_05870_),
    .A(net5787),
    .B(_05869_));
 sg13g2_xnor2_1 _36459_ (.Y(_05871_),
    .A(net5840),
    .B(_05869_));
 sg13g2_xnor2_1 _36460_ (.Y(_05872_),
    .A(net5787),
    .B(_05869_));
 sg13g2_nand3_1 _36461_ (.B(_05860_),
    .C(_05871_),
    .A(_05859_),
    .Y(_05873_));
 sg13g2_nor4_1 _36462_ (.A(_05835_),
    .B(_05846_),
    .C(_05847_),
    .D(_05873_),
    .Y(_05874_));
 sg13g2_xor2_1 _36463_ (.B(_05816_),
    .A(_03470_),
    .X(_05875_));
 sg13g2_o21ai_1 _36464_ (.B1(_03470_),
    .Y(_05876_),
    .A1(_03495_),
    .A2(_05823_));
 sg13g2_xor2_1 _36465_ (.B(_05824_),
    .A(_03470_),
    .X(_05877_));
 sg13g2_a21oi_1 _36466_ (.A1(net7198),
    .A2(\u_inv.d_next[210] ),
    .Y(_05878_),
    .B1(net6303));
 sg13g2_o21ai_1 _36467_ (.B1(_05878_),
    .Y(_05879_),
    .A1(net7199),
    .A2(_05877_));
 sg13g2_o21ai_1 _36468_ (.B1(_05879_),
    .Y(_05880_),
    .A1(net6219),
    .A2(_05875_));
 sg13g2_nor2_1 _36469_ (.A(net5840),
    .B(_05880_),
    .Y(_05881_));
 sg13g2_nand2b_1 _36470_ (.Y(_05882_),
    .B(net5787),
    .A_N(_05880_));
 sg13g2_nand2_1 _36471_ (.Y(_05883_),
    .A(net5840),
    .B(_05880_));
 sg13g2_xnor2_1 _36472_ (.Y(_05884_),
    .A(net5840),
    .B(_05880_));
 sg13g2_o21ai_1 _36473_ (.B1(_05876_),
    .Y(_05885_),
    .A1(_18113_),
    .A2(_18404_));
 sg13g2_a21oi_1 _36474_ (.A1(_03469_),
    .A2(_05885_),
    .Y(_05886_),
    .B1(net7198));
 sg13g2_o21ai_1 _36475_ (.B1(_05886_),
    .Y(_05887_),
    .A1(_03469_),
    .A2(_05885_));
 sg13g2_a21oi_1 _36476_ (.A1(net7198),
    .A2(\u_inv.d_next[211] ),
    .Y(_05888_),
    .B1(net6303));
 sg13g2_o21ai_1 _36477_ (.B1(_04689_),
    .Y(_05889_),
    .A1(_03470_),
    .A2(_05816_));
 sg13g2_or2_1 _36478_ (.X(_05890_),
    .B(_05889_),
    .A(_03469_));
 sg13g2_a21oi_1 _36479_ (.A1(_03469_),
    .A2(_05889_),
    .Y(_05891_),
    .B1(net6220));
 sg13g2_a22oi_1 _36480_ (.Y(_05892_),
    .B1(_05890_),
    .B2(_05891_),
    .A2(_05888_),
    .A1(_05887_));
 sg13g2_nand2_1 _36481_ (.Y(_05893_),
    .A(net5787),
    .B(_05892_));
 sg13g2_xnor2_1 _36482_ (.Y(_05894_),
    .A(net5787),
    .B(_05892_));
 sg13g2_a21oi_1 _36483_ (.A1(\u_inv.d_next[208] ),
    .A2(\u_inv.d_reg[208] ),
    .Y(_05895_),
    .B1(_05822_));
 sg13g2_xnor2_1 _36484_ (.Y(_05896_),
    .A(_03473_),
    .B(_05895_));
 sg13g2_o21ai_1 _36485_ (.B1(net6219),
    .Y(_05897_),
    .A1(net7334),
    .A2(_18114_));
 sg13g2_a21oi_1 _36486_ (.A1(net7334),
    .A2(_05896_),
    .Y(_05898_),
    .B1(_05897_));
 sg13g2_nor2_1 _36487_ (.A(_03474_),
    .B(_04686_),
    .Y(_05899_));
 sg13g2_a21oi_1 _36488_ (.A1(_03476_),
    .A2(_05723_),
    .Y(_05900_),
    .B1(net6219));
 sg13g2_a221oi_1 _36489_ (.B2(_05900_),
    .C1(_05898_),
    .B1(_05899_),
    .A1(net6303),
    .Y(_05901_),
    .A2(_05815_));
 sg13g2_xnor2_1 _36490_ (.Y(_05902_),
    .A(net5788),
    .B(_05901_));
 sg13g2_xnor2_1 _36491_ (.Y(_05903_),
    .A(_03476_),
    .B(_05723_));
 sg13g2_nand3_1 _36492_ (.B(_03476_),
    .C(_05730_),
    .A(_03431_),
    .Y(_05904_));
 sg13g2_nand3b_1 _36493_ (.B(_05904_),
    .C(net7334),
    .Y(_05905_),
    .A_N(_05822_));
 sg13g2_a21oi_1 _36494_ (.A1(net7198),
    .A2(\u_inv.d_next[208] ),
    .Y(_05906_),
    .B1(net6303));
 sg13g2_a22oi_1 _36495_ (.Y(_05907_),
    .B1(_05905_),
    .B2(_05906_),
    .A2(_05903_),
    .A1(net6303));
 sg13g2_nand2_1 _36496_ (.Y(_05908_),
    .A(net5788),
    .B(_05907_));
 sg13g2_xnor2_1 _36497_ (.Y(_05909_),
    .A(net5844),
    .B(_05907_));
 sg13g2_nor2b_1 _36498_ (.A(_05902_),
    .B_N(_05909_),
    .Y(_05910_));
 sg13g2_inv_1 _36499_ (.Y(_05911_),
    .A(_05910_));
 sg13g2_nor3_1 _36500_ (.A(_05884_),
    .B(_05894_),
    .C(_05911_),
    .Y(_05912_));
 sg13g2_nand2_1 _36501_ (.Y(_05913_),
    .A(_05874_),
    .B(_05912_));
 sg13g2_inv_1 _36502_ (.Y(_05914_),
    .A(_05913_));
 sg13g2_or4_1 _36503_ (.A(_05772_),
    .B(_05793_),
    .C(_05813_),
    .D(_05913_),
    .X(_05915_));
 sg13g2_o21ai_1 _36504_ (.B1(_04667_),
    .Y(_05916_),
    .A1(_04649_),
    .A2(_05353_));
 sg13g2_a21oi_2 _36505_ (.B1(_04661_),
    .Y(_05917_),
    .A2(_05916_),
    .A1(_04645_));
 sg13g2_nor3_1 _36506_ (.A(_04640_),
    .B(_04641_),
    .C(_05917_),
    .Y(_05918_));
 sg13g2_o21ai_1 _36507_ (.B1(_04637_),
    .Y(_05919_),
    .A1(_04676_),
    .A2(_05918_));
 sg13g2_a21oi_1 _36508_ (.A1(_04679_),
    .A2(_05919_),
    .Y(_05920_),
    .B1(_03360_));
 sg13g2_nand3_1 _36509_ (.B(_04679_),
    .C(_05919_),
    .A(_03360_),
    .Y(_05921_));
 sg13g2_nor2b_1 _36510_ (.A(_05920_),
    .B_N(_05921_),
    .Y(_05922_));
 sg13g2_a21oi_2 _36511_ (.B1(_03421_),
    .Y(_05923_),
    .A2(_04585_),
    .A1(net1080));
 sg13g2_o21ai_1 _36512_ (.B1(_03396_),
    .Y(_05924_),
    .A1(_03426_),
    .A2(_05923_));
 sg13g2_o21ai_1 _36513_ (.B1(_03399_),
    .Y(_05925_),
    .A1(_03427_),
    .A2(_05923_));
 sg13g2_a22oi_1 _36514_ (.Y(_05926_),
    .B1(_03386_),
    .B2(_05925_),
    .A2(_03381_),
    .A1(_03377_));
 sg13g2_o21ai_1 _36515_ (.B1(_03373_),
    .Y(_05927_),
    .A1(_03376_),
    .A2(_05926_));
 sg13g2_a21oi_1 _36516_ (.A1(_03370_),
    .A2(_05927_),
    .Y(_05928_),
    .B1(_03366_));
 sg13g2_xor2_1 _36517_ (.B(_05928_),
    .A(_03360_),
    .X(_05929_));
 sg13g2_o21ai_1 _36518_ (.B1(net6220),
    .Y(_05930_),
    .A1(net7333),
    .A2(\u_inv.d_next[206] ));
 sg13g2_a21oi_1 _36519_ (.A1(net7333),
    .A2(_05929_),
    .Y(_05931_),
    .B1(_05930_));
 sg13g2_a21oi_1 _36520_ (.A1(net6302),
    .A2(_05922_),
    .Y(_05932_),
    .B1(_05931_));
 sg13g2_or2_1 _36521_ (.X(_05933_),
    .B(_05932_),
    .A(net5840));
 sg13g2_xnor2_1 _36522_ (.Y(_05934_),
    .A(net5840),
    .B(_05932_));
 sg13g2_o21ai_1 _36523_ (.B1(_03359_),
    .Y(_05935_),
    .A1(_03358_),
    .A2(_05928_));
 sg13g2_a21oi_1 _36524_ (.A1(_03357_),
    .A2(_05935_),
    .Y(_05936_),
    .B1(net7199));
 sg13g2_o21ai_1 _36525_ (.B1(_05936_),
    .Y(_05937_),
    .A1(_03357_),
    .A2(_05935_));
 sg13g2_nand2_1 _36526_ (.Y(_05938_),
    .A(net7199),
    .B(\u_inv.d_next[207] ));
 sg13g2_nand3_1 _36527_ (.B(_05937_),
    .C(_05938_),
    .A(net6220),
    .Y(_05939_));
 sg13g2_or3_1 _36528_ (.A(_03357_),
    .B(_04681_),
    .C(_05920_),
    .X(_05940_));
 sg13g2_o21ai_1 _36529_ (.B1(_03357_),
    .Y(_05941_),
    .A1(_04681_),
    .A2(_05920_));
 sg13g2_nand3_1 _36530_ (.B(_05940_),
    .C(_05941_),
    .A(net6302),
    .Y(_05942_));
 sg13g2_and3_1 _36531_ (.X(_05943_),
    .A(net5788),
    .B(_05939_),
    .C(_05942_));
 sg13g2_nand3_1 _36532_ (.B(_05939_),
    .C(_05942_),
    .A(net5789),
    .Y(_05944_));
 sg13g2_a21oi_1 _36533_ (.A1(_05939_),
    .A2(_05942_),
    .Y(_05945_),
    .B1(net5788));
 sg13g2_nor2_1 _36534_ (.A(_05943_),
    .B(_05945_),
    .Y(_05946_));
 sg13g2_nor3_1 _36535_ (.A(_05934_),
    .B(_05943_),
    .C(_05945_),
    .Y(_05947_));
 sg13g2_a21oi_1 _36536_ (.A1(_03369_),
    .A2(_05927_),
    .Y(_05948_),
    .B1(_03365_));
 sg13g2_o21ai_1 _36537_ (.B1(net7333),
    .Y(_05949_),
    .A1(_03367_),
    .A2(_05948_));
 sg13g2_a21o_1 _36538_ (.A2(_05948_),
    .A1(_03367_),
    .B1(_05949_),
    .X(_05950_));
 sg13g2_nand2_1 _36539_ (.Y(_05951_),
    .A(net7199),
    .B(\u_inv.d_next[205] ));
 sg13g2_nand3_1 _36540_ (.B(_05950_),
    .C(_05951_),
    .A(net6222),
    .Y(_05952_));
 sg13g2_o21ai_1 _36541_ (.B1(_03368_),
    .Y(_05953_),
    .A1(_04676_),
    .A2(_05918_));
 sg13g2_a21o_1 _36542_ (.A2(_05953_),
    .A1(_04677_),
    .B1(_03367_),
    .X(_05954_));
 sg13g2_nand3_1 _36543_ (.B(_04677_),
    .C(_05953_),
    .A(_03367_),
    .Y(_05955_));
 sg13g2_nand3_1 _36544_ (.B(_05954_),
    .C(_05955_),
    .A(net6301),
    .Y(_05956_));
 sg13g2_a21o_1 _36545_ (.A2(_05956_),
    .A1(_05952_),
    .B1(net5789),
    .X(_05957_));
 sg13g2_nand3_1 _36546_ (.B(_05952_),
    .C(_05956_),
    .A(net5789),
    .Y(_05958_));
 sg13g2_nand2_1 _36547_ (.Y(_05959_),
    .A(_05957_),
    .B(_05958_));
 sg13g2_or3_1 _36548_ (.A(_03368_),
    .B(_04676_),
    .C(_05918_),
    .X(_05960_));
 sg13g2_and2_1 _36549_ (.A(net6302),
    .B(_05953_),
    .X(_05961_));
 sg13g2_xnor2_1 _36550_ (.Y(_05962_),
    .A(_03369_),
    .B(_05927_));
 sg13g2_o21ai_1 _36551_ (.B1(net6220),
    .Y(_05963_),
    .A1(net7338),
    .A2(\u_inv.d_next[204] ));
 sg13g2_a21oi_1 _36552_ (.A1(net7338),
    .A2(_05962_),
    .Y(_05964_),
    .B1(_05963_));
 sg13g2_a21oi_2 _36553_ (.B1(_05964_),
    .Y(_05965_),
    .A2(_05961_),
    .A1(_05960_));
 sg13g2_nor2_1 _36554_ (.A(net5841),
    .B(_05965_),
    .Y(_05966_));
 sg13g2_xnor2_1 _36555_ (.Y(_05967_),
    .A(net5789),
    .B(_05965_));
 sg13g2_nor2b_1 _36556_ (.A(_05959_),
    .B_N(_05967_),
    .Y(_05968_));
 sg13g2_nand3_1 _36557_ (.B(_05958_),
    .C(_05967_),
    .A(_05957_),
    .Y(_05969_));
 sg13g2_nor4_1 _36558_ (.A(_05934_),
    .B(_05943_),
    .C(_05945_),
    .D(_05969_),
    .Y(_05970_));
 sg13g2_o21ai_1 _36559_ (.B1(_04672_),
    .Y(_05971_),
    .A1(_04641_),
    .A2(_05917_));
 sg13g2_xnor2_1 _36560_ (.Y(_05972_),
    .A(_03375_),
    .B(_05971_));
 sg13g2_xor2_1 _36561_ (.B(_05926_),
    .A(_03375_),
    .X(_05973_));
 sg13g2_nand2_1 _36562_ (.Y(_05974_),
    .A(net7199),
    .B(\u_inv.d_next[202] ));
 sg13g2_a21oi_1 _36563_ (.A1(net7333),
    .A2(_05973_),
    .Y(_05975_),
    .B1(net6301));
 sg13g2_a22oi_1 _36564_ (.Y(_05976_),
    .B1(_05974_),
    .B2(_05975_),
    .A2(_05972_),
    .A1(net6301));
 sg13g2_and2_1 _36565_ (.A(net5790),
    .B(_05976_),
    .X(_05977_));
 sg13g2_xnor2_1 _36566_ (.Y(_05978_),
    .A(net5841),
    .B(_05976_));
 sg13g2_a21oi_1 _36567_ (.A1(_03375_),
    .A2(_05971_),
    .Y(_05979_),
    .B1(_04674_));
 sg13g2_or2_1 _36568_ (.X(_05980_),
    .B(_05979_),
    .A(_03374_));
 sg13g2_a21oi_1 _36569_ (.A1(_03374_),
    .A2(_05979_),
    .Y(_05981_),
    .B1(net6220));
 sg13g2_o21ai_1 _36570_ (.B1(_03371_),
    .Y(_05982_),
    .A1(_03375_),
    .A2(_05926_));
 sg13g2_xnor2_1 _36571_ (.Y(_05983_),
    .A(_03374_),
    .B(_05982_));
 sg13g2_nand2_1 _36572_ (.Y(_05984_),
    .A(net7199),
    .B(\u_inv.d_next[203] ));
 sg13g2_a21oi_1 _36573_ (.A1(net7333),
    .A2(_05983_),
    .Y(_05985_),
    .B1(net6301));
 sg13g2_a22oi_1 _36574_ (.Y(_05986_),
    .B1(_05984_),
    .B2(_05985_),
    .A2(_05981_),
    .A1(_05980_));
 sg13g2_xnor2_1 _36575_ (.Y(_05987_),
    .A(net5841),
    .B(_05986_));
 sg13g2_nand2_1 _36576_ (.Y(_05988_),
    .A(_05978_),
    .B(_05987_));
 sg13g2_xnor2_1 _36577_ (.Y(_05989_),
    .A(_03385_),
    .B(_05925_));
 sg13g2_o21ai_1 _36578_ (.B1(net6220),
    .Y(_05990_),
    .A1(net7333),
    .A2(\u_inv.d_next[200] ));
 sg13g2_a21oi_1 _36579_ (.A1(net7333),
    .A2(_05989_),
    .Y(_05991_),
    .B1(_05990_));
 sg13g2_xor2_1 _36580_ (.B(_05917_),
    .A(_03385_),
    .X(_05992_));
 sg13g2_a21oi_2 _36581_ (.B1(_05991_),
    .Y(_05993_),
    .A2(_05992_),
    .A1(net6302));
 sg13g2_or2_1 _36582_ (.X(_05994_),
    .B(_05993_),
    .A(net5840));
 sg13g2_xnor2_1 _36583_ (.Y(_05995_),
    .A(net5789),
    .B(_05993_));
 sg13g2_a21oi_1 _36584_ (.A1(_03385_),
    .A2(_05925_),
    .Y(_05996_),
    .B1(_03380_));
 sg13g2_o21ai_1 _36585_ (.B1(net7333),
    .Y(_05997_),
    .A1(_03384_),
    .A2(_05996_));
 sg13g2_a21o_1 _36586_ (.A2(_05996_),
    .A1(_03384_),
    .B1(_05997_),
    .X(_05998_));
 sg13g2_a21oi_1 _36587_ (.A1(net7199),
    .A2(\u_inv.d_next[201] ),
    .Y(_05999_),
    .B1(net6301));
 sg13g2_o21ai_1 _36588_ (.B1(_04670_),
    .Y(_06000_),
    .A1(_03385_),
    .A2(_05917_));
 sg13g2_nand2b_1 _36589_ (.Y(_06001_),
    .B(_03384_),
    .A_N(_06000_));
 sg13g2_a21oi_1 _36590_ (.A1(_03383_),
    .A2(_06000_),
    .Y(_06002_),
    .B1(net6220));
 sg13g2_a22oi_1 _36591_ (.Y(_06003_),
    .B1(_06001_),
    .B2(_06002_),
    .A2(_05999_),
    .A1(_05998_));
 sg13g2_nand2_1 _36592_ (.Y(_06004_),
    .A(net5790),
    .B(_06003_));
 sg13g2_xnor2_1 _36593_ (.Y(_06005_),
    .A(net5789),
    .B(_06003_));
 sg13g2_inv_1 _36594_ (.Y(_06006_),
    .A(_06005_));
 sg13g2_nand2_1 _36595_ (.Y(_06007_),
    .A(_05995_),
    .B(_06006_));
 sg13g2_inv_1 _36596_ (.Y(_06008_),
    .A(_06007_));
 sg13g2_nor2_1 _36597_ (.A(_05988_),
    .B(_06007_),
    .Y(_06009_));
 sg13g2_and2_1 _36598_ (.A(_05970_),
    .B(_06009_),
    .X(_06010_));
 sg13g2_nand2_1 _36599_ (.Y(_06011_),
    .A(_03392_),
    .B(_05924_));
 sg13g2_o21ai_1 _36600_ (.B1(net7335),
    .Y(_06012_),
    .A1(_03392_),
    .A2(_05924_));
 sg13g2_nand2b_1 _36601_ (.Y(_06013_),
    .B(_06011_),
    .A_N(_06012_));
 sg13g2_a21oi_1 _36602_ (.A1(_04643_),
    .A2(_05916_),
    .Y(_06014_),
    .B1(_04658_));
 sg13g2_xnor2_1 _36603_ (.Y(_06015_),
    .A(_03392_),
    .B(_06014_));
 sg13g2_a21oi_1 _36604_ (.A1(net7200),
    .A2(\u_inv.d_next[198] ),
    .Y(_06016_),
    .B1(net6301));
 sg13g2_a22oi_1 _36605_ (.Y(_06017_),
    .B1(_06016_),
    .B2(_06013_),
    .A2(_06015_),
    .A1(net6301));
 sg13g2_and2_1 _36606_ (.A(net5789),
    .B(_06017_),
    .X(_06018_));
 sg13g2_xnor2_1 _36607_ (.Y(_06019_),
    .A(net5791),
    .B(_06017_));
 sg13g2_inv_1 _36608_ (.Y(_06020_),
    .A(_06019_));
 sg13g2_nand3_1 _36609_ (.B(_03391_),
    .C(_06011_),
    .A(_03390_),
    .Y(_06021_));
 sg13g2_a21oi_1 _36610_ (.A1(_03391_),
    .A2(_06011_),
    .Y(_06022_),
    .B1(_03390_));
 sg13g2_nand2_1 _36611_ (.Y(_06023_),
    .A(net7335),
    .B(_06021_));
 sg13g2_a21oi_1 _36612_ (.A1(net7200),
    .A2(\u_inv.d_next[199] ),
    .Y(_06024_),
    .B1(net6301));
 sg13g2_o21ai_1 _36613_ (.B1(_06024_),
    .Y(_06025_),
    .A1(_06022_),
    .A2(_06023_));
 sg13g2_o21ai_1 _36614_ (.B1(_04655_),
    .Y(_06026_),
    .A1(_03392_),
    .A2(_06014_));
 sg13g2_xnor2_1 _36615_ (.Y(_06027_),
    .A(_03389_),
    .B(_06026_));
 sg13g2_o21ai_1 _36616_ (.B1(_06025_),
    .Y(_06028_),
    .A1(net6221),
    .A2(_06027_));
 sg13g2_nand2b_1 _36617_ (.Y(_06029_),
    .B(net5789),
    .A_N(_06028_));
 sg13g2_xnor2_1 _36618_ (.Y(_06030_),
    .A(net5791),
    .B(_06028_));
 sg13g2_nand2_1 _36619_ (.Y(_06031_),
    .A(_06020_),
    .B(_06030_));
 sg13g2_a21oi_1 _36620_ (.A1(_03425_),
    .A2(_05916_),
    .Y(_06032_),
    .B1(_04656_));
 sg13g2_o21ai_1 _36621_ (.B1(net6304),
    .Y(_06033_),
    .A1(_03423_),
    .A2(_06032_));
 sg13g2_a21oi_1 _36622_ (.A1(_03423_),
    .A2(_06032_),
    .Y(_06034_),
    .B1(_06033_));
 sg13g2_nor2_1 _36623_ (.A(_03425_),
    .B(_05923_),
    .Y(_06035_));
 sg13g2_a21o_1 _36624_ (.A2(\u_inv.d_reg[196] ),
    .A1(\u_inv.d_next[196] ),
    .B1(_06035_),
    .X(_06036_));
 sg13g2_o21ai_1 _36625_ (.B1(net7335),
    .Y(_06037_),
    .A1(_03422_),
    .A2(_06036_));
 sg13g2_a21o_1 _36626_ (.A2(_06036_),
    .A1(_03422_),
    .B1(_06037_),
    .X(_06038_));
 sg13g2_a21oi_1 _36627_ (.A1(net7200),
    .A2(\u_inv.d_next[197] ),
    .Y(_06039_),
    .B1(net6304));
 sg13g2_a21oi_2 _36628_ (.B1(_06034_),
    .Y(_06040_),
    .A2(_06039_),
    .A1(_06038_));
 sg13g2_inv_1 _36629_ (.Y(_06041_),
    .A(_06040_));
 sg13g2_xnor2_1 _36630_ (.Y(_06042_),
    .A(net5843),
    .B(_06040_));
 sg13g2_nand2_1 _36631_ (.Y(_06043_),
    .A(_03425_),
    .B(_05923_));
 sg13g2_nor2_1 _36632_ (.A(net7200),
    .B(_06035_),
    .Y(_06044_));
 sg13g2_xnor2_1 _36633_ (.Y(_06045_),
    .A(_03425_),
    .B(_05916_));
 sg13g2_a221oi_1 _36634_ (.B2(_06044_),
    .C1(net6304),
    .B1(_06043_),
    .A1(net7200),
    .Y(_06046_),
    .A2(\u_inv.d_next[196] ));
 sg13g2_a21oi_2 _36635_ (.B1(_06046_),
    .Y(_06047_),
    .A2(_06045_),
    .A1(net6304));
 sg13g2_nand2_1 _36636_ (.Y(_06048_),
    .A(net5791),
    .B(_06047_));
 sg13g2_xnor2_1 _36637_ (.Y(_06049_),
    .A(net5842),
    .B(_06047_));
 sg13g2_nand4_1 _36638_ (.B(_06030_),
    .C(_06042_),
    .A(_06020_),
    .Y(_06050_),
    .D(_06049_));
 sg13g2_o21ai_1 _36639_ (.B1(_04663_),
    .Y(_06051_),
    .A1(_04647_),
    .A2(_05353_));
 sg13g2_xor2_1 _36640_ (.B(_06051_),
    .A(_03411_),
    .X(_06052_));
 sg13g2_a21o_1 _36641_ (.A2(_05729_),
    .A1(_03417_),
    .B1(_03415_),
    .X(_06053_));
 sg13g2_a21o_1 _36642_ (.A2(_06053_),
    .A1(_03418_),
    .B1(_03411_),
    .X(_06054_));
 sg13g2_nand3_1 _36643_ (.B(_03418_),
    .C(_06053_),
    .A(_03411_),
    .Y(_06055_));
 sg13g2_nand3_1 _36644_ (.B(_06054_),
    .C(_06055_),
    .A(net7335),
    .Y(_06056_));
 sg13g2_a21oi_1 _36645_ (.A1(net7200),
    .A2(\u_inv.d_next[194] ),
    .Y(_06057_),
    .B1(net6304));
 sg13g2_nand2_1 _36646_ (.Y(_06058_),
    .A(_06056_),
    .B(_06057_));
 sg13g2_o21ai_1 _36647_ (.B1(_06058_),
    .Y(_06059_),
    .A1(net6221),
    .A2(_06052_));
 sg13g2_nor2_1 _36648_ (.A(net5842),
    .B(_06059_),
    .Y(_06060_));
 sg13g2_xnor2_1 _36649_ (.Y(_06061_),
    .A(net5791),
    .B(_06059_));
 sg13g2_inv_1 _36650_ (.Y(_06062_),
    .A(_06061_));
 sg13g2_a21o_1 _36651_ (.A2(_06054_),
    .A1(_03410_),
    .B1(_03409_),
    .X(_06063_));
 sg13g2_nand3_1 _36652_ (.B(_03410_),
    .C(_06054_),
    .A(_03409_),
    .Y(_06064_));
 sg13g2_nand3_1 _36653_ (.B(_06063_),
    .C(_06064_),
    .A(net7335),
    .Y(_06065_));
 sg13g2_a21oi_1 _36654_ (.A1(net7200),
    .A2(\u_inv.d_next[195] ),
    .Y(_06066_),
    .B1(net6304));
 sg13g2_a21oi_1 _36655_ (.A1(_03411_),
    .A2(_06051_),
    .Y(_06067_),
    .B1(_04664_));
 sg13g2_or2_1 _36656_ (.X(_06068_),
    .B(_06067_),
    .A(_03409_));
 sg13g2_a21oi_1 _36657_ (.A1(_03409_),
    .A2(_06067_),
    .Y(_06069_),
    .B1(net6221));
 sg13g2_a22oi_1 _36658_ (.Y(_06070_),
    .B1(_06068_),
    .B2(_06069_),
    .A2(_06066_),
    .A1(_06065_));
 sg13g2_xnor2_1 _36659_ (.Y(_06071_),
    .A(net5842),
    .B(_06070_));
 sg13g2_nand2_1 _36660_ (.Y(_06072_),
    .A(_06061_),
    .B(_06071_));
 sg13g2_xnor2_1 _36661_ (.Y(_06073_),
    .A(net1080),
    .B(_04584_));
 sg13g2_o21ai_1 _36662_ (.B1(net6221),
    .Y(_06074_),
    .A1(net7335),
    .A2(\u_inv.d_next[192] ));
 sg13g2_a21oi_1 _36663_ (.A1(net7335),
    .A2(_06073_),
    .Y(_06075_),
    .B1(_06074_));
 sg13g2_nor2_1 _36664_ (.A(_04584_),
    .B(_05353_),
    .Y(_06076_));
 sg13g2_xnor2_1 _36665_ (.Y(_06077_),
    .A(_04584_),
    .B(_05354_));
 sg13g2_a21oi_2 _36666_ (.B1(_06075_),
    .Y(_06078_),
    .A2(_06077_),
    .A1(net6304));
 sg13g2_nor2_1 _36667_ (.A(net5843),
    .B(_06078_),
    .Y(_06079_));
 sg13g2_or2_1 _36668_ (.X(_06080_),
    .B(_06076_),
    .A(_04662_));
 sg13g2_a21oi_1 _36669_ (.A1(_03416_),
    .A2(_06080_),
    .Y(_06081_),
    .B1(net6221));
 sg13g2_o21ai_1 _36670_ (.B1(_06081_),
    .Y(_06082_),
    .A1(_03416_),
    .A2(_06080_));
 sg13g2_nand3_1 _36671_ (.B(_03417_),
    .C(_05729_),
    .A(_03415_),
    .Y(_06083_));
 sg13g2_nand3_1 _36672_ (.B(_06053_),
    .C(_06083_),
    .A(net7335),
    .Y(_06084_));
 sg13g2_a21oi_1 _36673_ (.A1(net7200),
    .A2(\u_inv.d_next[193] ),
    .Y(_06085_),
    .B1(net6304));
 sg13g2_nand2_1 _36674_ (.Y(_06086_),
    .A(_06084_),
    .B(_06085_));
 sg13g2_nand2_2 _36675_ (.Y(_06087_),
    .A(_06082_),
    .B(_06086_));
 sg13g2_a21o_1 _36676_ (.A2(_06087_),
    .A1(_06078_),
    .B1(net5842),
    .X(_06088_));
 sg13g2_a21oi_1 _36677_ (.A1(net5791),
    .A2(_06070_),
    .Y(_06089_),
    .B1(_06060_));
 sg13g2_o21ai_1 _36678_ (.B1(_06089_),
    .Y(_06090_),
    .A1(_06072_),
    .A2(_06088_));
 sg13g2_nor2b_1 _36679_ (.A(_06050_),
    .B_N(_06090_),
    .Y(_06091_));
 sg13g2_o21ai_1 _36680_ (.B1(net5791),
    .Y(_06092_),
    .A1(_06040_),
    .A2(_06047_));
 sg13g2_o21ai_1 _36681_ (.B1(_06029_),
    .Y(_06093_),
    .A1(_06031_),
    .A2(_06092_));
 sg13g2_or3_1 _36682_ (.A(_06018_),
    .B(_06091_),
    .C(_06093_),
    .X(_06094_));
 sg13g2_nand3_1 _36683_ (.B(_06009_),
    .C(_06094_),
    .A(_05970_),
    .Y(_06095_));
 sg13g2_and2_1 _36684_ (.A(_05994_),
    .B(_06004_),
    .X(_06096_));
 sg13g2_a21oi_1 _36685_ (.A1(net5790),
    .A2(_05986_),
    .Y(_06097_),
    .B1(_05977_));
 sg13g2_o21ai_1 _36686_ (.B1(_06097_),
    .Y(_06098_),
    .A1(_05988_),
    .A2(_06096_));
 sg13g2_inv_1 _36687_ (.Y(_06099_),
    .A(_06098_));
 sg13g2_nand2_1 _36688_ (.Y(_06100_),
    .A(_05933_),
    .B(_05944_));
 sg13g2_o21ai_1 _36689_ (.B1(_05958_),
    .Y(_06101_),
    .A1(net5841),
    .A2(_05965_));
 sg13g2_a221oi_1 _36690_ (.B2(_05947_),
    .C1(_06100_),
    .B1(_06101_),
    .A1(_05970_),
    .Y(_06102_),
    .A2(_06098_));
 sg13g2_nand2_2 _36691_ (.Y(_06103_),
    .A(_06095_),
    .B(_06102_));
 sg13g2_a21o_2 _36692_ (.A2(_06102_),
    .A1(_06095_),
    .B1(_05915_),
    .X(_06104_));
 sg13g2_nand2_1 _36693_ (.Y(_06105_),
    .A(_05800_),
    .B(_05810_));
 sg13g2_nand3_1 _36694_ (.B(_05791_),
    .C(_06105_),
    .A(_05783_),
    .Y(_06106_));
 sg13g2_nand3_1 _36695_ (.B(_05790_),
    .C(_06106_),
    .A(_05782_),
    .Y(_06107_));
 sg13g2_o21ai_1 _36696_ (.B1(net5783),
    .Y(_06108_),
    .A1(_05740_),
    .A2(_05749_));
 sg13g2_nand2_1 _36697_ (.Y(_06109_),
    .A(_05761_),
    .B(_05768_));
 sg13g2_a22oi_1 _36698_ (.Y(_06110_),
    .B1(_06109_),
    .B2(_05752_),
    .A2(_06107_),
    .A1(_05771_));
 sg13g2_o21ai_1 _36699_ (.B1(net5788),
    .Y(_06111_),
    .A1(_05901_),
    .A2(_05907_));
 sg13g2_or3_1 _36700_ (.A(_05884_),
    .B(_05894_),
    .C(_06111_),
    .X(_06112_));
 sg13g2_and3_1 _36701_ (.X(_06113_),
    .A(_05882_),
    .B(_05893_),
    .C(_06112_));
 sg13g2_nand3_1 _36702_ (.B(_05893_),
    .C(_06112_),
    .A(_05882_),
    .Y(_06114_));
 sg13g2_nand2_1 _36703_ (.Y(_06115_),
    .A(_05859_),
    .B(_05870_));
 sg13g2_o21ai_1 _36704_ (.B1(_05834_),
    .Y(_06116_),
    .A1(net5839),
    .A2(_05845_));
 sg13g2_a221oi_1 _36705_ (.B2(_05849_),
    .C1(_06116_),
    .B1(_06115_),
    .A1(_05874_),
    .Y(_06117_),
    .A2(_06114_));
 sg13g2_or4_1 _36706_ (.A(_05772_),
    .B(_05793_),
    .C(_05813_),
    .D(_06117_),
    .X(_06118_));
 sg13g2_and3_1 _36707_ (.X(_06119_),
    .A(_06108_),
    .B(_06110_),
    .C(_06118_));
 sg13g2_and2_1 _36708_ (.A(_06104_),
    .B(_06119_),
    .X(_06120_));
 sg13g2_a21oi_1 _36709_ (.A1(_06104_),
    .A2(_06119_),
    .Y(_06121_),
    .B1(_05722_));
 sg13g2_nand2_1 _36710_ (.Y(_06122_),
    .A(_05532_),
    .B(_05539_));
 sg13g2_a21oi_1 _36711_ (.A1(_05511_),
    .A2(_05522_),
    .Y(_06123_),
    .B1(net5837));
 sg13g2_a21o_2 _36712_ (.A2(_06122_),
    .A1(_05524_),
    .B1(_06123_),
    .X(_06124_));
 sg13g2_o21ai_1 _36713_ (.B1(net5775),
    .Y(_06125_),
    .A1(_05471_),
    .A2(_05483_));
 sg13g2_o21ai_1 _36714_ (.B1(net5775),
    .Y(_06126_),
    .A1(_05490_),
    .A2(_05500_));
 sg13g2_nor3_1 _36715_ (.A(_05475_),
    .B(_05484_),
    .C(_06126_),
    .Y(_06127_));
 sg13g2_a21oi_1 _36716_ (.A1(_05503_),
    .A2(_06124_),
    .Y(_06128_),
    .B1(_06127_));
 sg13g2_nand2_1 _36717_ (.Y(_06129_),
    .A(_06125_),
    .B(_06128_));
 sg13g2_inv_1 _36718_ (.Y(_06130_),
    .A(_06129_));
 sg13g2_and3_1 _36719_ (.X(_06131_),
    .A(_05415_),
    .B(_05455_),
    .C(_06129_));
 sg13g2_nand2_1 _36720_ (.Y(_06132_),
    .A(_05445_),
    .B(_05451_));
 sg13g2_inv_1 _36721_ (.Y(_06133_),
    .A(_06132_));
 sg13g2_o21ai_1 _36722_ (.B1(net5776),
    .Y(_06134_),
    .A1(_05423_),
    .A2(_05434_));
 sg13g2_o21ai_1 _36723_ (.B1(_06134_),
    .Y(_06135_),
    .A1(_05436_),
    .A2(_06133_));
 sg13g2_nand2_1 _36724_ (.Y(_06136_),
    .A(_05415_),
    .B(_06135_));
 sg13g2_and2_1 _36725_ (.A(_05403_),
    .B(_05411_),
    .X(_06137_));
 sg13g2_or4_1 _36726_ (.A(_05380_),
    .B(_05391_),
    .C(_05393_),
    .D(_06137_),
    .X(_06138_));
 sg13g2_nand4_1 _36727_ (.B(_05392_),
    .C(_06136_),
    .A(_05379_),
    .Y(_06139_),
    .D(_06138_));
 sg13g2_and2_1 _36728_ (.A(_05599_),
    .B(_05609_),
    .X(_06140_));
 sg13g2_o21ai_1 _36729_ (.B1(net5778),
    .Y(_06141_),
    .A1(_05617_),
    .A2(_05627_));
 sg13g2_o21ai_1 _36730_ (.B1(_06141_),
    .Y(_06142_),
    .A1(_05629_),
    .A2(_06140_));
 sg13g2_inv_1 _36731_ (.Y(_06143_),
    .A(_06142_));
 sg13g2_nand2_1 _36732_ (.Y(_06144_),
    .A(_05592_),
    .B(_06142_));
 sg13g2_o21ai_1 _36733_ (.B1(net5777),
    .Y(_06145_),
    .A1(_05558_),
    .A2(_05568_));
 sg13g2_a21o_1 _36734_ (.A2(_05588_),
    .A1(net5778),
    .B1(_05578_),
    .X(_06146_));
 sg13g2_nand2_1 _36735_ (.Y(_06147_),
    .A(_05570_),
    .B(_06146_));
 sg13g2_nand2_1 _36736_ (.Y(_06148_),
    .A(_05709_),
    .B(_05716_));
 sg13g2_nand3_1 _36737_ (.B(_05700_),
    .C(_06148_),
    .A(_05690_),
    .Y(_06149_));
 sg13g2_o21ai_1 _36738_ (.B1(net5780),
    .Y(_06150_),
    .A1(_05688_),
    .A2(_05699_));
 sg13g2_nand2_1 _36739_ (.Y(_06151_),
    .A(_06149_),
    .B(_06150_));
 sg13g2_or2_1 _36740_ (.X(_06152_),
    .B(_05656_),
    .A(_05648_));
 sg13g2_nand2_1 _36741_ (.Y(_06153_),
    .A(_05667_),
    .B(_05679_));
 sg13g2_inv_1 _36742_ (.Y(_06154_),
    .A(_06153_));
 sg13g2_a22oi_1 _36743_ (.Y(_06155_),
    .B1(_06153_),
    .B2(_05658_),
    .A2(_06151_),
    .A1(_05682_));
 sg13g2_a221oi_1 _36744_ (.B2(_05658_),
    .C1(_06152_),
    .B1(_06153_),
    .A1(_05682_),
    .Y(_06156_),
    .A2(_06151_));
 sg13g2_nand2b_2 _36745_ (.Y(_06157_),
    .B(_06155_),
    .A_N(_06152_));
 sg13g2_nor4_1 _36746_ (.A(_05560_),
    .B(_05569_),
    .C(_05590_),
    .D(_05629_),
    .Y(_06158_));
 sg13g2_nand3b_1 _36747_ (.B(_06158_),
    .C(_05611_),
    .Y(_06159_),
    .A_N(_06156_));
 sg13g2_and4_1 _36748_ (.A(_06144_),
    .B(_06145_),
    .C(_06147_),
    .D(_06159_),
    .X(_06160_));
 sg13g2_nand4_1 _36749_ (.B(_06145_),
    .C(_06147_),
    .A(_06144_),
    .Y(_06161_),
    .D(_06159_));
 sg13g2_and4_1 _36750_ (.A(_05415_),
    .B(_05455_),
    .C(_05543_),
    .D(_06161_),
    .X(_06162_));
 sg13g2_and3_1 _36751_ (.X(_06163_),
    .A(_05503_),
    .B(_05524_),
    .C(_05541_));
 sg13g2_nand3_1 _36752_ (.B(_05720_),
    .C(_06158_),
    .A(_05611_),
    .Y(_06164_));
 sg13g2_nor4_2 _36753_ (.A(_06121_),
    .B(_06131_),
    .C(_06139_),
    .Y(_06165_),
    .D(_06162_));
 sg13g2_a21oi_2 _36754_ (.B1(_05270_),
    .Y(_06166_),
    .A2(_05205_),
    .A1(_05148_));
 sg13g2_o21ai_1 _36755_ (.B1(_05309_),
    .Y(_06167_),
    .A1(_05156_),
    .A2(_06166_));
 sg13g2_a21oi_1 _36756_ (.A1(_05157_),
    .A2(_06167_),
    .Y(_06168_),
    .B1(_05312_));
 sg13g2_xnor2_1 _36757_ (.Y(_06169_),
    .A(_03707_),
    .B(_06168_));
 sg13g2_a21oi_2 _36758_ (.B1(_04575_),
    .Y(_06170_),
    .A2(_04525_),
    .A1(_04422_));
 sg13g2_a21o_2 _36759_ (.A2(_04525_),
    .A1(_04422_),
    .B1(_04575_),
    .X(_06171_));
 sg13g2_nor2_1 _36760_ (.A(_03668_),
    .B(_06170_),
    .Y(_06172_));
 sg13g2_a21oi_1 _36761_ (.A1(_03665_),
    .A2(_06172_),
    .Y(_06173_),
    .B1(_03787_));
 sg13g2_nor2_1 _36762_ (.A(_03673_),
    .B(_06170_),
    .Y(_06174_));
 sg13g2_nor2b_1 _36763_ (.A(_06174_),
    .B_N(_03789_),
    .Y(_06175_));
 sg13g2_o21ai_1 _36764_ (.B1(_03789_),
    .Y(_06176_),
    .A1(_03673_),
    .A2(_06170_));
 sg13g2_nand2b_1 _36765_ (.Y(_06177_),
    .B(_06176_),
    .A_N(_03705_));
 sg13g2_nand2_1 _36766_ (.Y(_06178_),
    .A(_03714_),
    .B(_06176_));
 sg13g2_nand3_1 _36767_ (.B(_03801_),
    .C(_06178_),
    .A(_03708_),
    .Y(_06179_));
 sg13g2_a21o_1 _36768_ (.A2(_06178_),
    .A1(_03801_),
    .B1(_03708_),
    .X(_06180_));
 sg13g2_nand3_1 _36769_ (.B(_06179_),
    .C(_06180_),
    .A(net7348),
    .Y(_06181_));
 sg13g2_a21oi_1 _36770_ (.A1(net7208),
    .A2(\u_inv.d_next[166] ),
    .Y(_06182_),
    .B1(net6316));
 sg13g2_a22oi_1 _36771_ (.Y(_06183_),
    .B1(_06181_),
    .B2(_06182_),
    .A2(_06169_),
    .A1(net6316));
 sg13g2_nand2_1 _36772_ (.Y(_06184_),
    .A(net5800),
    .B(_06183_));
 sg13g2_xnor2_1 _36773_ (.Y(_06185_),
    .A(net5800),
    .B(_06183_));
 sg13g2_nand3_1 _36774_ (.B(_03711_),
    .C(_06180_),
    .A(_03706_),
    .Y(_06186_));
 sg13g2_a21o_1 _36775_ (.A2(_06180_),
    .A1(_03706_),
    .B1(_03711_),
    .X(_06187_));
 sg13g2_nand3_1 _36776_ (.B(_06186_),
    .C(_06187_),
    .A(net7348),
    .Y(_06188_));
 sg13g2_a21oi_1 _36777_ (.A1(net7208),
    .A2(\u_inv.d_next[167] ),
    .Y(_06189_),
    .B1(net6316));
 sg13g2_o21ai_1 _36778_ (.B1(_05313_),
    .Y(_06190_),
    .A1(_03707_),
    .A2(_06168_));
 sg13g2_nand2b_1 _36779_ (.Y(_06191_),
    .B(_03711_),
    .A_N(_06190_));
 sg13g2_a21oi_1 _36780_ (.A1(_03710_),
    .A2(_06190_),
    .Y(_06192_),
    .B1(net6228));
 sg13g2_a22oi_1 _36781_ (.Y(_06193_),
    .B1(_06191_),
    .B2(_06192_),
    .A2(_06189_),
    .A1(_06188_));
 sg13g2_nand2_1 _36782_ (.Y(_06194_),
    .A(net5801),
    .B(_06193_));
 sg13g2_xnor2_1 _36783_ (.Y(_06195_),
    .A(net5801),
    .B(_06193_));
 sg13g2_nor2_1 _36784_ (.A(_06185_),
    .B(_06195_),
    .Y(_06196_));
 sg13g2_a21oi_1 _36785_ (.A1(_03705_),
    .A2(_06167_),
    .Y(_06197_),
    .B1(_05310_));
 sg13g2_o21ai_1 _36786_ (.B1(net6316),
    .Y(_06198_),
    .A1(_03713_),
    .A2(_06197_));
 sg13g2_a21oi_1 _36787_ (.A1(_03713_),
    .A2(_06197_),
    .Y(_06199_),
    .B1(_06198_));
 sg13g2_nand2_1 _36788_ (.Y(_06200_),
    .A(_03704_),
    .B(_06177_));
 sg13g2_xnor2_1 _36789_ (.Y(_06201_),
    .A(_03713_),
    .B(_06200_));
 sg13g2_o21ai_1 _36790_ (.B1(net6228),
    .Y(_06202_),
    .A1(net7348),
    .A2(_18124_));
 sg13g2_a21oi_1 _36791_ (.A1(net7348),
    .A2(_06201_),
    .Y(_06203_),
    .B1(_06202_));
 sg13g2_nor2_1 _36792_ (.A(_06199_),
    .B(_06203_),
    .Y(_06204_));
 sg13g2_nand2_1 _36793_ (.Y(_06205_),
    .A(net5799),
    .B(_06204_));
 sg13g2_xnor2_1 _36794_ (.Y(_06206_),
    .A(net5849),
    .B(_06204_));
 sg13g2_a21oi_1 _36795_ (.A1(_03705_),
    .A2(_06175_),
    .Y(_06207_),
    .B1(net7207));
 sg13g2_xnor2_1 _36796_ (.Y(_06208_),
    .A(_03705_),
    .B(_06167_));
 sg13g2_a221oi_1 _36797_ (.B2(_06207_),
    .C1(net6315),
    .B1(_06177_),
    .A1(net7207),
    .Y(_06209_),
    .A2(\u_inv.d_next[164] ));
 sg13g2_a21oi_2 _36798_ (.B1(_06209_),
    .Y(_06210_),
    .A2(_06208_),
    .A1(net6315));
 sg13g2_nand2_1 _36799_ (.Y(_06211_),
    .A(net5800),
    .B(_06210_));
 sg13g2_xnor2_1 _36800_ (.Y(_06212_),
    .A(net5801),
    .B(_06210_));
 sg13g2_nor3_1 _36801_ (.A(_06185_),
    .B(_06195_),
    .C(_06212_),
    .Y(_06213_));
 sg13g2_nand2_1 _36802_ (.Y(_06214_),
    .A(_06206_),
    .B(_06213_));
 sg13g2_xnor2_1 _36803_ (.Y(_06215_),
    .A(_03668_),
    .B(_06170_));
 sg13g2_o21ai_1 _36804_ (.B1(net6228),
    .Y(_06216_),
    .A1(net7348),
    .A2(\u_inv.d_next[160] ));
 sg13g2_a21oi_1 _36805_ (.A1(net7348),
    .A2(_06215_),
    .Y(_06217_),
    .B1(_06216_));
 sg13g2_xnor2_1 _36806_ (.Y(_06218_),
    .A(_03668_),
    .B(_06166_));
 sg13g2_a21oi_1 _36807_ (.A1(net6315),
    .A2(_06218_),
    .Y(_06219_),
    .B1(_06217_));
 sg13g2_nor2_1 _36808_ (.A(net5850),
    .B(_06219_),
    .Y(_06220_));
 sg13g2_xnor2_1 _36809_ (.Y(_06221_),
    .A(net5849),
    .B(_06219_));
 sg13g2_o21ai_1 _36810_ (.B1(_05305_),
    .Y(_06222_),
    .A1(_05155_),
    .A2(_06166_));
 sg13g2_xor2_1 _36811_ (.B(_06222_),
    .A(_03671_),
    .X(_06223_));
 sg13g2_or2_1 _36812_ (.X(_06224_),
    .B(_06173_),
    .A(_03671_));
 sg13g2_a21oi_1 _36813_ (.A1(_03671_),
    .A2(_06173_),
    .Y(_06225_),
    .B1(net7208));
 sg13g2_nand2_1 _36814_ (.Y(_06226_),
    .A(_06224_),
    .B(_06225_));
 sg13g2_a21oi_1 _36815_ (.A1(net7207),
    .A2(\u_inv.d_next[162] ),
    .Y(_06227_),
    .B1(net6315));
 sg13g2_nand2_1 _36816_ (.Y(_06228_),
    .A(_06226_),
    .B(_06227_));
 sg13g2_o21ai_1 _36817_ (.B1(_06228_),
    .Y(_06229_),
    .A1(net6228),
    .A2(_06223_));
 sg13g2_nand2b_1 _36818_ (.Y(_06230_),
    .B(net5801),
    .A_N(_06229_));
 sg13g2_xnor2_1 _36819_ (.Y(_06231_),
    .A(net5801),
    .B(_06229_));
 sg13g2_inv_1 _36820_ (.Y(_06232_),
    .A(_06231_));
 sg13g2_a21oi_1 _36821_ (.A1(_03671_),
    .A2(_06222_),
    .Y(_06233_),
    .B1(_05307_));
 sg13g2_or2_1 _36822_ (.X(_06234_),
    .B(_06233_),
    .A(_03669_));
 sg13g2_a21oi_1 _36823_ (.A1(_03669_),
    .A2(_06233_),
    .Y(_06235_),
    .B1(net6228));
 sg13g2_a21o_1 _36824_ (.A2(_06224_),
    .A1(_03670_),
    .B1(_03669_),
    .X(_06236_));
 sg13g2_nand3_1 _36825_ (.B(_03670_),
    .C(_06224_),
    .A(_03669_),
    .Y(_06237_));
 sg13g2_nand3_1 _36826_ (.B(_06236_),
    .C(_06237_),
    .A(net7348),
    .Y(_06238_));
 sg13g2_a21oi_1 _36827_ (.A1(net7207),
    .A2(\u_inv.d_next[163] ),
    .Y(_06239_),
    .B1(net6315));
 sg13g2_a22oi_1 _36828_ (.Y(_06240_),
    .B1(_06238_),
    .B2(_06239_),
    .A2(_06235_),
    .A1(_06234_));
 sg13g2_nand2_1 _36829_ (.Y(_06241_),
    .A(net5801),
    .B(_06240_));
 sg13g2_xnor2_1 _36830_ (.Y(_06242_),
    .A(net5850),
    .B(_06240_));
 sg13g2_nand2_1 _36831_ (.Y(_06243_),
    .A(_06231_),
    .B(_06242_));
 sg13g2_o21ai_1 _36832_ (.B1(_05303_),
    .Y(_06244_),
    .A1(_03667_),
    .A2(_06166_));
 sg13g2_o21ai_1 _36833_ (.B1(net6315),
    .Y(_06245_),
    .A1(_03665_),
    .A2(_06244_));
 sg13g2_a21oi_1 _36834_ (.A1(_03665_),
    .A2(_06244_),
    .Y(_06246_),
    .B1(_06245_));
 sg13g2_nand2_1 _36835_ (.Y(_06247_),
    .A(_03664_),
    .B(_03666_));
 sg13g2_o21ai_1 _36836_ (.B1(net7349),
    .Y(_06248_),
    .A1(_03664_),
    .A2(_03666_));
 sg13g2_a21oi_1 _36837_ (.A1(_03665_),
    .A2(_06172_),
    .Y(_06249_),
    .B1(_06248_));
 sg13g2_o21ai_1 _36838_ (.B1(_06249_),
    .Y(_06250_),
    .A1(_06172_),
    .A2(_06247_));
 sg13g2_a21oi_1 _36839_ (.A1(net7207),
    .A2(\u_inv.d_next[161] ),
    .Y(_06251_),
    .B1(net6315));
 sg13g2_a21oi_1 _36840_ (.A1(_06250_),
    .A2(_06251_),
    .Y(_06252_),
    .B1(_06246_));
 sg13g2_xnor2_1 _36841_ (.Y(_06253_),
    .A(net5799),
    .B(_06252_));
 sg13g2_nor2_1 _36842_ (.A(_06243_),
    .B(_06253_),
    .Y(_06254_));
 sg13g2_or2_1 _36843_ (.X(_06255_),
    .B(_06253_),
    .A(_06221_));
 sg13g2_inv_1 _36844_ (.Y(_06256_),
    .A(_06255_));
 sg13g2_nor3_1 _36845_ (.A(_06214_),
    .B(_06243_),
    .C(_06255_),
    .Y(_06257_));
 sg13g2_inv_1 _36846_ (.Y(_06258_),
    .A(_06257_));
 sg13g2_nor3_1 _36847_ (.A(_05156_),
    .B(_05159_),
    .C(_06166_),
    .Y(_06259_));
 sg13g2_nor2_1 _36848_ (.A(_05316_),
    .B(_06259_),
    .Y(_06260_));
 sg13g2_o21ai_1 _36849_ (.B1(_05153_),
    .Y(_06261_),
    .A1(_05316_),
    .A2(_06259_));
 sg13g2_o21ai_1 _36850_ (.B1(_05323_),
    .Y(_06262_),
    .A1(_05152_),
    .A2(_06261_));
 sg13g2_a21oi_1 _36851_ (.A1(_05150_),
    .A2(_06262_),
    .Y(_06263_),
    .B1(_05326_));
 sg13g2_xnor2_1 _36852_ (.Y(_06264_),
    .A(_03677_),
    .B(_06263_));
 sg13g2_a21oi_2 _36853_ (.B1(_03804_),
    .Y(_06265_),
    .A2(_06176_),
    .A1(_03716_));
 sg13g2_nand2b_1 _36854_ (.Y(_06266_),
    .B(_03693_),
    .A_N(_06265_));
 sg13g2_o21ai_1 _36855_ (.B1(_03798_),
    .Y(_06267_),
    .A1(_03701_),
    .A2(_06265_));
 sg13g2_a21oi_1 _36856_ (.A1(_03687_),
    .A2(_06267_),
    .Y(_06268_),
    .B1(_03790_));
 sg13g2_xnor2_1 _36857_ (.Y(_06269_),
    .A(_03677_),
    .B(_06268_));
 sg13g2_nand2_1 _36858_ (.Y(_06270_),
    .A(net7205),
    .B(\u_inv.d_next[174] ));
 sg13g2_a21oi_1 _36859_ (.A1(net7347),
    .A2(_06269_),
    .Y(_06271_),
    .B1(net6313));
 sg13g2_a22oi_1 _36860_ (.Y(_06272_),
    .B1(_06270_),
    .B2(_06271_),
    .A2(_06264_),
    .A1(net6313));
 sg13g2_nand2_1 _36861_ (.Y(_06273_),
    .A(net5799),
    .B(_06272_));
 sg13g2_xnor2_1 _36862_ (.Y(_06274_),
    .A(net5799),
    .B(_06272_));
 sg13g2_inv_1 _36863_ (.Y(_06275_),
    .A(_06274_));
 sg13g2_o21ai_1 _36864_ (.B1(_03676_),
    .Y(_06276_),
    .A1(_03675_),
    .A2(_06268_));
 sg13g2_a21oi_1 _36865_ (.A1(_03674_),
    .A2(_06276_),
    .Y(_06277_),
    .B1(net7205));
 sg13g2_o21ai_1 _36866_ (.B1(_06277_),
    .Y(_06278_),
    .A1(_03674_),
    .A2(_06276_));
 sg13g2_a21oi_1 _36867_ (.A1(net7205),
    .A2(\u_inv.d_next[175] ),
    .Y(_06279_),
    .B1(net6314));
 sg13g2_nand2_1 _36868_ (.Y(_06280_),
    .A(_06278_),
    .B(_06279_));
 sg13g2_o21ai_1 _36869_ (.B1(_05327_),
    .Y(_06281_),
    .A1(_03677_),
    .A2(_06263_));
 sg13g2_xnor2_1 _36870_ (.Y(_06282_),
    .A(_03674_),
    .B(_06281_));
 sg13g2_o21ai_1 _36871_ (.B1(_06280_),
    .Y(_06283_),
    .A1(net6229),
    .A2(_06282_));
 sg13g2_xnor2_1 _36872_ (.Y(_06284_),
    .A(net5851),
    .B(_06283_));
 sg13g2_nor2_1 _36873_ (.A(_06274_),
    .B(_06284_),
    .Y(_06285_));
 sg13g2_nand2_1 _36874_ (.Y(_06286_),
    .A(_03685_),
    .B(_06267_));
 sg13g2_xnor2_1 _36875_ (.Y(_06287_),
    .A(_03685_),
    .B(_06267_));
 sg13g2_o21ai_1 _36876_ (.B1(net6229),
    .Y(_06288_),
    .A1(net7347),
    .A2(\u_inv.d_next[172] ));
 sg13g2_a21o_1 _36877_ (.A2(_06287_),
    .A1(net7346),
    .B1(_06288_),
    .X(_06289_));
 sg13g2_xnor2_1 _36878_ (.Y(_06290_),
    .A(_03686_),
    .B(_06262_));
 sg13g2_o21ai_1 _36879_ (.B1(_06289_),
    .Y(_06291_),
    .A1(net6229),
    .A2(_06290_));
 sg13g2_nand2_1 _36880_ (.Y(_06292_),
    .A(net5799),
    .B(_06291_));
 sg13g2_xnor2_1 _36881_ (.Y(_06293_),
    .A(net5799),
    .B(_06291_));
 sg13g2_and2_1 _36882_ (.A(_03684_),
    .B(_06286_),
    .X(_06294_));
 sg13g2_a21oi_1 _36883_ (.A1(_03683_),
    .A2(_06294_),
    .Y(_06295_),
    .B1(net7205));
 sg13g2_o21ai_1 _36884_ (.B1(_06295_),
    .Y(_06296_),
    .A1(_03683_),
    .A2(_06294_));
 sg13g2_a21oi_1 _36885_ (.A1(net7205),
    .A2(\u_inv.d_next[173] ),
    .Y(_06297_),
    .B1(net6313));
 sg13g2_a21oi_1 _36886_ (.A1(_03686_),
    .A2(_06262_),
    .Y(_06298_),
    .B1(_05324_));
 sg13g2_nand2b_1 _36887_ (.Y(_06299_),
    .B(_03682_),
    .A_N(_06298_));
 sg13g2_a21oi_1 _36888_ (.A1(_03683_),
    .A2(_06298_),
    .Y(_06300_),
    .B1(net6229));
 sg13g2_a22oi_1 _36889_ (.Y(_06301_),
    .B1(_06299_),
    .B2(_06300_),
    .A2(_06297_),
    .A1(_06296_));
 sg13g2_nand2_1 _36890_ (.Y(_06302_),
    .A(net5799),
    .B(_06301_));
 sg13g2_or2_1 _36891_ (.X(_06303_),
    .B(_06301_),
    .A(net5849));
 sg13g2_nand2_1 _36892_ (.Y(_06304_),
    .A(net5849),
    .B(_06301_));
 sg13g2_xnor2_1 _36893_ (.Y(_06305_),
    .A(net5849),
    .B(_06301_));
 sg13g2_nand2b_1 _36894_ (.Y(_06306_),
    .B(_06305_),
    .A_N(_06293_));
 sg13g2_nor3_1 _36895_ (.A(_06274_),
    .B(_06284_),
    .C(_06306_),
    .Y(_06307_));
 sg13g2_a21o_1 _36896_ (.A2(_06266_),
    .A1(_03795_),
    .B1(_03699_),
    .X(_06308_));
 sg13g2_nand2_1 _36897_ (.Y(_06309_),
    .A(_03698_),
    .B(_06308_));
 sg13g2_o21ai_1 _36898_ (.B1(net7347),
    .Y(_06310_),
    .A1(_03696_),
    .A2(_06309_));
 sg13g2_a21o_1 _36899_ (.A2(_06309_),
    .A1(_03696_),
    .B1(_06310_),
    .X(_06311_));
 sg13g2_a21oi_1 _36900_ (.A1(net7205),
    .A2(\u_inv.d_next[171] ),
    .Y(_06312_),
    .B1(net6313));
 sg13g2_nor2b_1 _36901_ (.A(_05318_),
    .B_N(_06261_),
    .Y(_06313_));
 sg13g2_nand2b_1 _36902_ (.Y(_06314_),
    .B(_06261_),
    .A_N(_05319_));
 sg13g2_a21oi_1 _36903_ (.A1(_03699_),
    .A2(_06314_),
    .Y(_06315_),
    .B1(_05320_));
 sg13g2_xnor2_1 _36904_ (.Y(_06316_),
    .A(_03696_),
    .B(_06315_));
 sg13g2_a22oi_1 _36905_ (.Y(_06317_),
    .B1(_06316_),
    .B2(net6314),
    .A2(_06312_),
    .A1(_06311_));
 sg13g2_xnor2_1 _36906_ (.Y(_06318_),
    .A(net5800),
    .B(_06317_));
 sg13g2_nand3_1 _36907_ (.B(_03795_),
    .C(_06266_),
    .A(_03699_),
    .Y(_06319_));
 sg13g2_nand3_1 _36908_ (.B(_06308_),
    .C(_06319_),
    .A(net7347),
    .Y(_06320_));
 sg13g2_nand2_1 _36909_ (.Y(_06321_),
    .A(net7205),
    .B(\u_inv.d_next[170] ));
 sg13g2_a21oi_1 _36910_ (.A1(_06320_),
    .A2(_06321_),
    .Y(_06322_),
    .B1(net6313));
 sg13g2_xor2_1 _36911_ (.B(_06314_),
    .A(_03699_),
    .X(_06323_));
 sg13g2_a21oi_2 _36912_ (.B1(_06322_),
    .Y(_06324_),
    .A2(_06323_),
    .A1(net6314));
 sg13g2_nor2_1 _36913_ (.A(net5849),
    .B(_06324_),
    .Y(_06325_));
 sg13g2_xnor2_1 _36914_ (.Y(_06326_),
    .A(net5849),
    .B(_06324_));
 sg13g2_nor2_1 _36915_ (.A(_06318_),
    .B(_06326_),
    .Y(_06327_));
 sg13g2_nand2b_1 _36916_ (.Y(_06328_),
    .B(_03692_),
    .A_N(_06265_));
 sg13g2_o21ai_1 _36917_ (.B1(_06328_),
    .Y(_06329_),
    .A1(_18123_),
    .A2(_18446_));
 sg13g2_o21ai_1 _36918_ (.B1(net7348),
    .Y(_06330_),
    .A1(_03689_),
    .A2(_06329_));
 sg13g2_a21oi_1 _36919_ (.A1(_03689_),
    .A2(_06329_),
    .Y(_06331_),
    .B1(_06330_));
 sg13g2_a21oi_1 _36920_ (.A1(net7205),
    .A2(\u_inv.d_next[169] ),
    .Y(_06332_),
    .B1(_06331_));
 sg13g2_o21ai_1 _36921_ (.B1(_05317_),
    .Y(_06333_),
    .A1(_03692_),
    .A2(_06260_));
 sg13g2_o21ai_1 _36922_ (.B1(_06313_),
    .Y(_06334_),
    .A1(_03690_),
    .A2(_06333_));
 sg13g2_mux2_1 _36923_ (.A0(_06332_),
    .A1(_06334_),
    .S(net6314),
    .X(_06335_));
 sg13g2_nor2_1 _36924_ (.A(net5849),
    .B(_06335_),
    .Y(_06336_));
 sg13g2_xnor2_1 _36925_ (.Y(_06337_),
    .A(net5800),
    .B(_06335_));
 sg13g2_inv_1 _36926_ (.Y(_06338_),
    .A(_06337_));
 sg13g2_xnor2_1 _36927_ (.Y(_06339_),
    .A(_03692_),
    .B(_06260_));
 sg13g2_a21oi_1 _36928_ (.A1(_03691_),
    .A2(_06265_),
    .Y(_06340_),
    .B1(net7208));
 sg13g2_nand2_1 _36929_ (.Y(_06341_),
    .A(_06328_),
    .B(_06340_));
 sg13g2_a21oi_1 _36930_ (.A1(net7207),
    .A2(\u_inv.d_next[168] ),
    .Y(_06342_),
    .B1(net6314));
 sg13g2_a22oi_1 _36931_ (.Y(_06343_),
    .B1(_06341_),
    .B2(_06342_),
    .A2(_06339_),
    .A1(net6313));
 sg13g2_and2_1 _36932_ (.A(net5800),
    .B(_06343_),
    .X(_06344_));
 sg13g2_xnor2_1 _36933_ (.Y(_06345_),
    .A(net5800),
    .B(_06343_));
 sg13g2_nor2_1 _36934_ (.A(_06338_),
    .B(_06345_),
    .Y(_06346_));
 sg13g2_and2_1 _36935_ (.A(_06327_),
    .B(_06346_),
    .X(_06347_));
 sg13g2_nand4_1 _36936_ (.B(_06307_),
    .C(_06327_),
    .A(_06257_),
    .Y(_06348_),
    .D(_06346_));
 sg13g2_o21ai_1 _36937_ (.B1(_05332_),
    .Y(_06349_),
    .A1(_05161_),
    .A2(_06166_));
 sg13g2_a21oi_2 _36938_ (.B1(_05288_),
    .Y(_06350_),
    .A2(_06349_),
    .A1(_05173_));
 sg13g2_nor3_1 _36939_ (.A(_05166_),
    .B(_05167_),
    .C(_06350_),
    .Y(_06351_));
 sg13g2_nor2_1 _36940_ (.A(_05296_),
    .B(_06351_),
    .Y(_06352_));
 sg13g2_o21ai_1 _36941_ (.B1(_05164_),
    .Y(_06353_),
    .A1(_05296_),
    .A2(_06351_));
 sg13g2_a21oi_1 _36942_ (.A1(_05299_),
    .A2(_06353_),
    .Y(_06354_),
    .B1(_03746_));
 sg13g2_nand3_1 _36943_ (.B(_05299_),
    .C(_06353_),
    .A(_03746_),
    .Y(_06355_));
 sg13g2_nand2b_1 _36944_ (.Y(_06356_),
    .B(_06355_),
    .A_N(_06354_));
 sg13g2_a21oi_2 _36945_ (.B1(_03807_),
    .Y(_06357_),
    .A2(_06171_),
    .A1(_03717_));
 sg13g2_a21o_2 _36946_ (.A2(_06171_),
    .A1(_03717_),
    .B1(_03807_),
    .X(_06358_));
 sg13g2_o21ai_1 _36947_ (.B1(_03778_),
    .Y(_06359_),
    .A1(_03739_),
    .A2(_06357_));
 sg13g2_a21o_2 _36948_ (.A2(_06359_),
    .A1(_03766_),
    .B1(_03780_),
    .X(_06360_));
 sg13g2_a21oi_1 _36949_ (.A1(_03761_),
    .A2(_06360_),
    .Y(_06361_),
    .B1(_03781_));
 sg13g2_a21o_1 _36950_ (.A2(_06360_),
    .A1(_03761_),
    .B1(_03781_),
    .X(_06362_));
 sg13g2_a21oi_1 _36951_ (.A1(_03753_),
    .A2(_06362_),
    .Y(_06363_),
    .B1(_03783_));
 sg13g2_a21oi_1 _36952_ (.A1(_03745_),
    .A2(_06363_),
    .Y(_06364_),
    .B1(net7201));
 sg13g2_o21ai_1 _36953_ (.B1(_06364_),
    .Y(_06365_),
    .A1(_03745_),
    .A2(_06363_));
 sg13g2_a21oi_1 _36954_ (.A1(net7201),
    .A2(\u_inv.d_next[190] ),
    .Y(_06366_),
    .B1(net6305));
 sg13g2_a22oi_1 _36955_ (.Y(_06367_),
    .B1(_06365_),
    .B2(_06366_),
    .A2(_06356_),
    .A1(net6305));
 sg13g2_and2_1 _36956_ (.A(net5792),
    .B(_06367_),
    .X(_06368_));
 sg13g2_xnor2_1 _36957_ (.Y(_06369_),
    .A(net5792),
    .B(_06367_));
 sg13g2_o21ai_1 _36958_ (.B1(_03742_),
    .Y(_06370_),
    .A1(_05300_),
    .A2(_06354_));
 sg13g2_nor3_1 _36959_ (.A(_03742_),
    .B(_05300_),
    .C(_06354_),
    .Y(_06371_));
 sg13g2_nand3b_1 _36960_ (.B(net6306),
    .C(_06370_),
    .Y(_06372_),
    .A_N(_06371_));
 sg13g2_o21ai_1 _36961_ (.B1(_03744_),
    .Y(_06373_),
    .A1(_03745_),
    .A2(_06363_));
 sg13g2_a21oi_1 _36962_ (.A1(_03742_),
    .A2(_06373_),
    .Y(_06374_),
    .B1(net7201));
 sg13g2_o21ai_1 _36963_ (.B1(_06374_),
    .Y(_06375_),
    .A1(_03742_),
    .A2(_06373_));
 sg13g2_nand2_1 _36964_ (.Y(_06376_),
    .A(net7201),
    .B(\u_inv.d_next[191] ));
 sg13g2_nand3_1 _36965_ (.B(_06375_),
    .C(_06376_),
    .A(net6222),
    .Y(_06377_));
 sg13g2_and3_2 _36966_ (.X(_06378_),
    .A(net5791),
    .B(_06372_),
    .C(_06377_));
 sg13g2_a21oi_1 _36967_ (.A1(_06372_),
    .A2(_06377_),
    .Y(_06379_),
    .B1(net5792));
 sg13g2_nor2_1 _36968_ (.A(_06378_),
    .B(_06379_),
    .Y(_06380_));
 sg13g2_o21ai_1 _36969_ (.B1(_03752_),
    .Y(_06381_),
    .A1(_05296_),
    .A2(_06351_));
 sg13g2_a21o_1 _36970_ (.A2(_06381_),
    .A1(_05297_),
    .B1(_03750_),
    .X(_06382_));
 sg13g2_nand3_1 _36971_ (.B(_05297_),
    .C(_06381_),
    .A(_03750_),
    .Y(_06383_));
 sg13g2_nand3_1 _36972_ (.B(_06382_),
    .C(_06383_),
    .A(net6306),
    .Y(_06384_));
 sg13g2_o21ai_1 _36973_ (.B1(_03751_),
    .Y(_06385_),
    .A1(_03752_),
    .A2(_06361_));
 sg13g2_xor2_1 _36974_ (.B(_06385_),
    .A(_03750_),
    .X(_06386_));
 sg13g2_a21oi_1 _36975_ (.A1(net7202),
    .A2(\u_inv.d_next[189] ),
    .Y(_06387_),
    .B1(net6306));
 sg13g2_o21ai_1 _36976_ (.B1(_06387_),
    .Y(_06388_),
    .A1(net7202),
    .A2(_06386_));
 sg13g2_and2_1 _36977_ (.A(_06384_),
    .B(_06388_),
    .X(_06389_));
 sg13g2_nand3_1 _36978_ (.B(_06384_),
    .C(_06388_),
    .A(net5792),
    .Y(_06390_));
 sg13g2_a21o_1 _36979_ (.A2(_06388_),
    .A1(_06384_),
    .B1(net5792),
    .X(_06391_));
 sg13g2_nand2_1 _36980_ (.Y(_06392_),
    .A(_06390_),
    .B(_06391_));
 sg13g2_xnor2_1 _36981_ (.Y(_06393_),
    .A(_03752_),
    .B(_06361_));
 sg13g2_o21ai_1 _36982_ (.B1(net6222),
    .Y(_06394_),
    .A1(net7337),
    .A2(\u_inv.d_next[188] ));
 sg13g2_a21oi_1 _36983_ (.A1(net7337),
    .A2(_06393_),
    .Y(_06395_),
    .B1(_06394_));
 sg13g2_xnor2_1 _36984_ (.Y(_06396_),
    .A(_03752_),
    .B(_06352_));
 sg13g2_a21oi_2 _36985_ (.B1(_06395_),
    .Y(_06397_),
    .A2(_06396_),
    .A1(net6305));
 sg13g2_nor2_1 _36986_ (.A(net5844),
    .B(_06397_),
    .Y(_06398_));
 sg13g2_xnor2_1 _36987_ (.Y(_06399_),
    .A(net5792),
    .B(_06397_));
 sg13g2_nand3_1 _36988_ (.B(_06391_),
    .C(_06399_),
    .A(_06390_),
    .Y(_06400_));
 sg13g2_nor4_2 _36989_ (.A(_06369_),
    .B(_06378_),
    .C(_06379_),
    .Y(_06401_),
    .D(_06400_));
 sg13g2_nand2b_1 _36990_ (.Y(_06402_),
    .B(_06360_),
    .A_N(_03760_));
 sg13g2_nand2_1 _36991_ (.Y(_06403_),
    .A(_03759_),
    .B(_06402_));
 sg13g2_o21ai_1 _36992_ (.B1(net7336),
    .Y(_06404_),
    .A1(_03758_),
    .A2(_06403_));
 sg13g2_a21o_1 _36993_ (.A2(_06403_),
    .A1(_03758_),
    .B1(_06404_),
    .X(_06405_));
 sg13g2_a21oi_1 _36994_ (.A1(net7201),
    .A2(\u_inv.d_next[187] ),
    .Y(_06406_),
    .B1(net6305));
 sg13g2_o21ai_1 _36995_ (.B1(_05294_),
    .Y(_06407_),
    .A1(_05167_),
    .A2(_06350_));
 sg13g2_a21oi_1 _36996_ (.A1(_03760_),
    .A2(_06407_),
    .Y(_06408_),
    .B1(_05290_));
 sg13g2_xnor2_1 _36997_ (.Y(_06409_),
    .A(_03758_),
    .B(_06408_));
 sg13g2_a22oi_1 _36998_ (.Y(_06410_),
    .B1(_06409_),
    .B2(net6305),
    .A2(_06406_),
    .A1(_06405_));
 sg13g2_nand2_1 _36999_ (.Y(_06411_),
    .A(net5798),
    .B(_06410_));
 sg13g2_xnor2_1 _37000_ (.Y(_06412_),
    .A(net5798),
    .B(_06410_));
 sg13g2_xor2_1 _37001_ (.B(_06360_),
    .A(_03760_),
    .X(_06413_));
 sg13g2_o21ai_1 _37002_ (.B1(net6222),
    .Y(_06414_),
    .A1(net7337),
    .A2(\u_inv.d_next[186] ));
 sg13g2_a21oi_1 _37003_ (.A1(net7336),
    .A2(_06413_),
    .Y(_06415_),
    .B1(_06414_));
 sg13g2_xor2_1 _37004_ (.B(_06407_),
    .A(_03760_),
    .X(_06416_));
 sg13g2_a21oi_1 _37005_ (.A1(net6305),
    .A2(_06416_),
    .Y(_06417_),
    .B1(_06415_));
 sg13g2_or2_1 _37006_ (.X(_06418_),
    .B(_06417_),
    .A(net5844));
 sg13g2_xnor2_1 _37007_ (.Y(_06419_),
    .A(net5796),
    .B(_06417_));
 sg13g2_nor2b_1 _37008_ (.A(_06412_),
    .B_N(_06419_),
    .Y(_06420_));
 sg13g2_a21oi_1 _37009_ (.A1(_03765_),
    .A2(_06359_),
    .Y(_06421_),
    .B1(_03764_));
 sg13g2_a21oi_1 _37010_ (.A1(_03763_),
    .A2(_06421_),
    .Y(_06422_),
    .B1(net7201));
 sg13g2_o21ai_1 _37011_ (.B1(_06422_),
    .Y(_06423_),
    .A1(_03763_),
    .A2(_06421_));
 sg13g2_a21oi_1 _37012_ (.A1(net7201),
    .A2(\u_inv.d_next[185] ),
    .Y(_06424_),
    .B1(net6305));
 sg13g2_o21ai_1 _37013_ (.B1(_05291_),
    .Y(_06425_),
    .A1(_03765_),
    .A2(_06350_));
 sg13g2_nand2b_1 _37014_ (.Y(_06426_),
    .B(_03763_),
    .A_N(_06425_));
 sg13g2_a21oi_1 _37015_ (.A1(_03762_),
    .A2(_06425_),
    .Y(_06427_),
    .B1(net6221));
 sg13g2_a22oi_1 _37016_ (.Y(_06428_),
    .B1(_06426_),
    .B2(_06427_),
    .A2(_06424_),
    .A1(_06423_));
 sg13g2_nand2_1 _37017_ (.Y(_06429_),
    .A(net5797),
    .B(_06428_));
 sg13g2_xnor2_1 _37018_ (.Y(_06430_),
    .A(net5843),
    .B(_06428_));
 sg13g2_xnor2_1 _37019_ (.Y(_06431_),
    .A(_03765_),
    .B(_06359_));
 sg13g2_o21ai_1 _37020_ (.B1(net6221),
    .Y(_06432_),
    .A1(net7336),
    .A2(\u_inv.d_next[184] ));
 sg13g2_a21o_1 _37021_ (.A2(_06431_),
    .A1(net7336),
    .B1(_06432_),
    .X(_06433_));
 sg13g2_xnor2_1 _37022_ (.Y(_06434_),
    .A(_03765_),
    .B(_06350_));
 sg13g2_o21ai_1 _37023_ (.B1(_06433_),
    .Y(_06435_),
    .A1(net6221),
    .A2(_06434_));
 sg13g2_nand2_1 _37024_ (.Y(_06436_),
    .A(net5796),
    .B(_06435_));
 sg13g2_nor2_1 _37025_ (.A(net5797),
    .B(_06435_),
    .Y(_06437_));
 sg13g2_xnor2_1 _37026_ (.Y(_06438_),
    .A(net5843),
    .B(_06435_));
 sg13g2_nand2_1 _37027_ (.Y(_06439_),
    .A(_06430_),
    .B(_06438_));
 sg13g2_and3_2 _37028_ (.X(_06440_),
    .A(_06420_),
    .B(_06430_),
    .C(_06438_));
 sg13g2_inv_1 _37029_ (.Y(_06441_),
    .A(_06440_));
 sg13g2_nand2_2 _37030_ (.Y(_06442_),
    .A(_06401_),
    .B(_06440_));
 sg13g2_a21oi_1 _37031_ (.A1(_05172_),
    .A2(_06349_),
    .Y(_06443_),
    .B1(_05279_));
 sg13g2_a21o_1 _37032_ (.A2(_06349_),
    .A1(_05172_),
    .B1(_05279_),
    .X(_06444_));
 sg13g2_a221oi_1 _37033_ (.B2(_06444_),
    .C1(_05284_),
    .B1(_05169_),
    .A1(\u_inv.d_next[181] ),
    .Y(_06445_),
    .A2(_18433_));
 sg13g2_o21ai_1 _37034_ (.B1(_05282_),
    .Y(_06446_),
    .A1(_03719_),
    .A2(_06445_));
 sg13g2_or2_1 _37035_ (.X(_06447_),
    .B(_06446_),
    .A(_03720_));
 sg13g2_a21oi_1 _37036_ (.A1(_03720_),
    .A2(_06446_),
    .Y(_06448_),
    .B1(net6229));
 sg13g2_a21oi_2 _37037_ (.B1(_03772_),
    .Y(_06449_),
    .A2(_06358_),
    .A1(_03738_));
 sg13g2_o21ai_1 _37038_ (.B1(_03774_),
    .Y(_06450_),
    .A1(_03734_),
    .A2(_06449_));
 sg13g2_a21oi_1 _37039_ (.A1(_03725_),
    .A2(_06450_),
    .Y(_06451_),
    .B1(_03770_));
 sg13g2_nor2b_1 _37040_ (.A(_06451_),
    .B_N(_03719_),
    .Y(_06452_));
 sg13g2_or3_1 _37041_ (.A(_03718_),
    .B(_03720_),
    .C(_06452_),
    .X(_06453_));
 sg13g2_o21ai_1 _37042_ (.B1(_03720_),
    .Y(_06454_),
    .A1(_03718_),
    .A2(_06452_));
 sg13g2_nand3_1 _37043_ (.B(_06453_),
    .C(_06454_),
    .A(net7346),
    .Y(_06455_));
 sg13g2_a21oi_1 _37044_ (.A1(net7206),
    .A2(\u_inv.d_next[183] ),
    .Y(_06456_),
    .B1(net6311));
 sg13g2_a22oi_1 _37045_ (.Y(_06457_),
    .B1(_06455_),
    .B2(_06456_),
    .A2(_06448_),
    .A1(_06447_));
 sg13g2_nand2_1 _37046_ (.Y(_06458_),
    .A(net5796),
    .B(_06457_));
 sg13g2_xnor2_1 _37047_ (.Y(_06459_),
    .A(net5796),
    .B(_06457_));
 sg13g2_nand2b_1 _37048_ (.Y(_06460_),
    .B(_06451_),
    .A_N(_03719_));
 sg13g2_nand3b_1 _37049_ (.B(_06460_),
    .C(net7346),
    .Y(_06461_),
    .A_N(_06452_));
 sg13g2_xnor2_1 _37050_ (.Y(_06462_),
    .A(_03719_),
    .B(_06445_));
 sg13g2_a21oi_1 _37051_ (.A1(net7206),
    .A2(\u_inv.d_next[182] ),
    .Y(_06463_),
    .B1(net6311));
 sg13g2_a22oi_1 _37052_ (.Y(_06464_),
    .B1(_06463_),
    .B2(_06461_),
    .A2(_06462_),
    .A1(net6311));
 sg13g2_nand2_1 _37053_ (.Y(_06465_),
    .A(net5796),
    .B(_06464_));
 sg13g2_xnor2_1 _37054_ (.Y(_06466_),
    .A(net5796),
    .B(_06464_));
 sg13g2_nor2_1 _37055_ (.A(_06459_),
    .B(_06466_),
    .Y(_06467_));
 sg13g2_xnor2_1 _37056_ (.Y(_06468_),
    .A(_03724_),
    .B(_06443_));
 sg13g2_or2_1 _37057_ (.X(_06469_),
    .B(_06450_),
    .A(_03724_));
 sg13g2_a21oi_1 _37058_ (.A1(_03724_),
    .A2(_06450_),
    .Y(_06470_),
    .B1(net7206));
 sg13g2_nand2_1 _37059_ (.Y(_06471_),
    .A(net7206),
    .B(\u_inv.d_next[180] ));
 sg13g2_a21oi_1 _37060_ (.A1(_06469_),
    .A2(_06470_),
    .Y(_06472_),
    .B1(net6311));
 sg13g2_a22oi_1 _37061_ (.Y(_06473_),
    .B1(_06471_),
    .B2(_06472_),
    .A2(_06468_),
    .A1(net6311));
 sg13g2_nand2_1 _37062_ (.Y(_06474_),
    .A(net5798),
    .B(_06473_));
 sg13g2_xnor2_1 _37063_ (.Y(_06475_),
    .A(net5796),
    .B(_06473_));
 sg13g2_o21ai_1 _37064_ (.B1(_05283_),
    .Y(_06476_),
    .A1(_03724_),
    .A2(_06443_));
 sg13g2_o21ai_1 _37065_ (.B1(net6311),
    .Y(_06477_),
    .A1(_03722_),
    .A2(_06476_));
 sg13g2_a21oi_1 _37066_ (.A1(_03722_),
    .A2(_06476_),
    .Y(_06478_),
    .B1(_06477_));
 sg13g2_a21oi_1 _37067_ (.A1(_03724_),
    .A2(_06450_),
    .Y(_06479_),
    .B1(_03723_));
 sg13g2_xnor2_1 _37068_ (.Y(_06480_),
    .A(_03722_),
    .B(_06479_));
 sg13g2_o21ai_1 _37069_ (.B1(net6229),
    .Y(_06481_),
    .A1(net7346),
    .A2(_18119_));
 sg13g2_a21oi_1 _37070_ (.A1(net7346),
    .A2(_06480_),
    .Y(_06482_),
    .B1(_06481_));
 sg13g2_nor2_1 _37071_ (.A(_06478_),
    .B(_06482_),
    .Y(_06483_));
 sg13g2_nand2_1 _37072_ (.Y(_06484_),
    .A(net5798),
    .B(_06483_));
 sg13g2_xnor2_1 _37073_ (.Y(_06485_),
    .A(net5796),
    .B(_06483_));
 sg13g2_nor2_1 _37074_ (.A(_06475_),
    .B(_06485_),
    .Y(_06486_));
 sg13g2_nor4_1 _37075_ (.A(_06459_),
    .B(_06466_),
    .C(_06475_),
    .D(_06485_),
    .Y(_06487_));
 sg13g2_a21oi_1 _37076_ (.A1(_05171_),
    .A2(_06349_),
    .Y(_06488_),
    .B1(_05276_));
 sg13g2_xnor2_1 _37077_ (.Y(_06489_),
    .A(_03728_),
    .B(_06488_));
 sg13g2_xnor2_1 _37078_ (.Y(_06490_),
    .A(_03728_),
    .B(_06449_));
 sg13g2_nand2_1 _37079_ (.Y(_06491_),
    .A(net7206),
    .B(\u_inv.d_next[178] ));
 sg13g2_a21oi_1 _37080_ (.A1(net7346),
    .A2(_06490_),
    .Y(_06492_),
    .B1(net6311));
 sg13g2_a22oi_1 _37081_ (.Y(_06493_),
    .B1(_06491_),
    .B2(_06492_),
    .A2(_06489_),
    .A1(net6312));
 sg13g2_nand2_1 _37082_ (.Y(_06494_),
    .A(net5797),
    .B(_06493_));
 sg13g2_xnor2_1 _37083_ (.Y(_06495_),
    .A(net5797),
    .B(_06493_));
 sg13g2_o21ai_1 _37084_ (.B1(_05273_),
    .Y(_06496_),
    .A1(_03728_),
    .A2(_06488_));
 sg13g2_nand2b_1 _37085_ (.Y(_06497_),
    .B(_03732_),
    .A_N(_06496_));
 sg13g2_a21oi_1 _37086_ (.A1(_03731_),
    .A2(_06496_),
    .Y(_06498_),
    .B1(net6229));
 sg13g2_o21ai_1 _37087_ (.B1(_03726_),
    .Y(_06499_),
    .A1(_03727_),
    .A2(_06449_));
 sg13g2_xnor2_1 _37088_ (.Y(_06500_),
    .A(_03732_),
    .B(_06499_));
 sg13g2_nand2_1 _37089_ (.Y(_06501_),
    .A(net7206),
    .B(\u_inv.d_next[179] ));
 sg13g2_a21oi_1 _37090_ (.A1(net7346),
    .A2(_06500_),
    .Y(_06502_),
    .B1(net6312));
 sg13g2_a22oi_1 _37091_ (.Y(_06503_),
    .B1(_06501_),
    .B2(_06502_),
    .A2(_06498_),
    .A1(_06497_));
 sg13g2_xnor2_1 _37092_ (.Y(_06504_),
    .A(net5851),
    .B(_06503_));
 sg13g2_nor2b_1 _37093_ (.A(_06495_),
    .B_N(_06504_),
    .Y(_06505_));
 sg13g2_nand2b_1 _37094_ (.Y(_06506_),
    .B(_06504_),
    .A_N(_06495_));
 sg13g2_xnor2_1 _37095_ (.Y(_06507_),
    .A(_03737_),
    .B(_06349_));
 sg13g2_nand2b_1 _37096_ (.Y(_06508_),
    .B(_06358_),
    .A_N(_03737_));
 sg13g2_a21oi_1 _37097_ (.A1(_03737_),
    .A2(_06357_),
    .Y(_06509_),
    .B1(net7206));
 sg13g2_a221oi_1 _37098_ (.B2(_06509_),
    .C1(net6312),
    .B1(_06508_),
    .A1(net7209),
    .Y(_06510_),
    .A2(\u_inv.d_next[176] ));
 sg13g2_a21oi_2 _37099_ (.B1(_06510_),
    .Y(_06511_),
    .A2(_06507_),
    .A1(net6311));
 sg13g2_nand2_1 _37100_ (.Y(_06512_),
    .A(net5797),
    .B(_06511_));
 sg13g2_xnor2_1 _37101_ (.Y(_06513_),
    .A(net5797),
    .B(_06511_));
 sg13g2_a21oi_1 _37102_ (.A1(_03737_),
    .A2(_06349_),
    .Y(_06514_),
    .B1(_05274_));
 sg13g2_a21oi_1 _37103_ (.A1(_03735_),
    .A2(_06514_),
    .Y(_06515_),
    .B1(net6229));
 sg13g2_o21ai_1 _37104_ (.B1(_06515_),
    .Y(_06516_),
    .A1(_03735_),
    .A2(_06514_));
 sg13g2_nand3_1 _37105_ (.B(_03736_),
    .C(_06508_),
    .A(_03735_),
    .Y(_06517_));
 sg13g2_a21o_1 _37106_ (.A2(_06508_),
    .A1(_03736_),
    .B1(_03735_),
    .X(_06518_));
 sg13g2_nand3_1 _37107_ (.B(_06517_),
    .C(_06518_),
    .A(net7347),
    .Y(_06519_));
 sg13g2_o21ai_1 _37108_ (.B1(_06519_),
    .Y(_06520_),
    .A1(net7346),
    .A2(_18121_));
 sg13g2_o21ai_1 _37109_ (.B1(_06516_),
    .Y(_06521_),
    .A1(net6312),
    .A2(_06520_));
 sg13g2_nor2_1 _37110_ (.A(net5851),
    .B(_06521_),
    .Y(_06522_));
 sg13g2_xnor2_1 _37111_ (.Y(_06523_),
    .A(net5851),
    .B(_06521_));
 sg13g2_nor2_1 _37112_ (.A(_06513_),
    .B(_06523_),
    .Y(_06524_));
 sg13g2_nand2_1 _37113_ (.Y(_06525_),
    .A(_04422_),
    .B(net6994));
 sg13g2_nand3_1 _37114_ (.B(_04517_),
    .C(_04521_),
    .A(_04422_),
    .Y(_06526_));
 sg13g2_nand3_1 _37115_ (.B(_04519_),
    .C(net6994),
    .A(_04422_),
    .Y(_06527_));
 sg13g2_nand3b_1 _37116_ (.B(_04523_),
    .C(_04422_),
    .Y(_06528_),
    .A_N(_04495_));
 sg13g2_a21oi_1 _37117_ (.A1(_04550_),
    .A2(_06528_),
    .Y(_06529_),
    .B1(_04447_));
 sg13g2_a21o_2 _37118_ (.A2(_06528_),
    .A1(_04550_),
    .B1(_04448_),
    .X(_06530_));
 sg13g2_a21oi_1 _37119_ (.A1(_04564_),
    .A2(_06530_),
    .Y(_06531_),
    .B1(_04440_));
 sg13g2_o21ai_1 _37120_ (.B1(_04433_),
    .Y(_06532_),
    .A1(_04567_),
    .A2(_06531_));
 sg13g2_a21o_1 _37121_ (.A2(_06532_),
    .A1(_04571_),
    .B1(_04427_),
    .X(_06533_));
 sg13g2_a21oi_1 _37122_ (.A1(_04425_),
    .A2(_06533_),
    .Y(_06534_),
    .B1(_04424_));
 sg13g2_nand3_1 _37123_ (.B(_04425_),
    .C(_06533_),
    .A(_04424_),
    .Y(_06535_));
 sg13g2_nor2_1 _37124_ (.A(net7215),
    .B(_06534_),
    .Y(_06536_));
 sg13g2_a221oi_1 _37125_ (.B2(_06536_),
    .C1(net6325),
    .B1(_06535_),
    .A1(net7215),
    .Y(_06537_),
    .A2(\u_inv.d_next[151] ));
 sg13g2_a21oi_2 _37126_ (.B1(_05236_),
    .Y(_06538_),
    .A2(_05204_),
    .A1(_05148_));
 sg13g2_nor3_1 _37127_ (.A(_05186_),
    .B(_05187_),
    .C(_06538_),
    .Y(_06539_));
 sg13g2_o21ai_1 _37128_ (.B1(_05184_),
    .Y(_06540_),
    .A1(_05258_),
    .A2(_06539_));
 sg13g2_a21oi_1 _37129_ (.A1(_05261_),
    .A2(_06540_),
    .Y(_06541_),
    .B1(_04426_));
 sg13g2_nor3_1 _37130_ (.A(_04423_),
    .B(_05262_),
    .C(_06541_),
    .Y(_06542_));
 sg13g2_o21ai_1 _37131_ (.B1(_04423_),
    .Y(_06543_),
    .A1(_05262_),
    .A2(_06541_));
 sg13g2_nor2_1 _37132_ (.A(net6239),
    .B(_06542_),
    .Y(_06544_));
 sg13g2_a21o_1 _37133_ (.A2(_06544_),
    .A1(_06543_),
    .B1(_06537_),
    .X(_06545_));
 sg13g2_inv_1 _37134_ (.Y(_06546_),
    .A(_06545_));
 sg13g2_xnor2_1 _37135_ (.Y(_06547_),
    .A(net5805),
    .B(_06545_));
 sg13g2_nand3_1 _37136_ (.B(_05261_),
    .C(_06540_),
    .A(_04426_),
    .Y(_06548_));
 sg13g2_nor2_1 _37137_ (.A(net6239),
    .B(_06541_),
    .Y(_06549_));
 sg13g2_nand3_1 _37138_ (.B(_04571_),
    .C(_06532_),
    .A(_04427_),
    .Y(_06550_));
 sg13g2_nand3_1 _37139_ (.B(_06533_),
    .C(_06550_),
    .A(net7363),
    .Y(_06551_));
 sg13g2_o21ai_1 _37140_ (.B1(_06551_),
    .Y(_06552_),
    .A1(net7363),
    .A2(_18128_));
 sg13g2_a22oi_1 _37141_ (.Y(_06553_),
    .B1(_06552_),
    .B2(net6239),
    .A2(_06549_),
    .A1(_06548_));
 sg13g2_nor2_1 _37142_ (.A(net5856),
    .B(_06553_),
    .Y(_06554_));
 sg13g2_xnor2_1 _37143_ (.Y(_06555_),
    .A(net5805),
    .B(_06553_));
 sg13g2_nor3_1 _37144_ (.A(_04431_),
    .B(_05258_),
    .C(_06539_),
    .Y(_06556_));
 sg13g2_o21ai_1 _37145_ (.B1(_04431_),
    .Y(_06557_),
    .A1(_05258_),
    .A2(_06539_));
 sg13g2_nand2b_1 _37146_ (.Y(_06558_),
    .B(_06557_),
    .A_N(_06556_));
 sg13g2_o21ai_1 _37147_ (.B1(_04432_),
    .Y(_06559_),
    .A1(_04567_),
    .A2(_06531_));
 sg13g2_nor3_1 _37148_ (.A(_04432_),
    .B(_04567_),
    .C(_06531_),
    .Y(_06560_));
 sg13g2_nor2_1 _37149_ (.A(net7214),
    .B(_06560_),
    .Y(_06561_));
 sg13g2_a221oi_1 _37150_ (.B2(_06561_),
    .C1(net6326),
    .B1(_06559_),
    .A1(net7214),
    .Y(_06562_),
    .A2(\u_inv.d_next[148] ));
 sg13g2_a21oi_2 _37151_ (.B1(_06562_),
    .Y(_06563_),
    .A2(_06558_),
    .A1(net6326));
 sg13g2_nand2_1 _37152_ (.Y(_06564_),
    .A(net5805),
    .B(_06563_));
 sg13g2_xnor2_1 _37153_ (.Y(_06565_),
    .A(net5805),
    .B(_06563_));
 sg13g2_inv_1 _37154_ (.Y(_06566_),
    .A(_06565_));
 sg13g2_a21o_1 _37155_ (.A2(_06559_),
    .A1(_04430_),
    .B1(_04429_),
    .X(_06567_));
 sg13g2_nand3_1 _37156_ (.B(_04430_),
    .C(_06559_),
    .A(_04429_),
    .Y(_06568_));
 sg13g2_nand3_1 _37157_ (.B(_06567_),
    .C(_06568_),
    .A(net7363),
    .Y(_06569_));
 sg13g2_a21oi_1 _37158_ (.A1(net7218),
    .A2(\u_inv.d_next[149] ),
    .Y(_06570_),
    .B1(net6327));
 sg13g2_nand2b_1 _37159_ (.Y(_06571_),
    .B(_06557_),
    .A_N(_05259_));
 sg13g2_xnor2_1 _37160_ (.Y(_06572_),
    .A(_04429_),
    .B(_06571_));
 sg13g2_a22oi_1 _37161_ (.Y(_06573_),
    .B1(_06572_),
    .B2(net6327),
    .A2(_06570_),
    .A1(_06569_));
 sg13g2_xnor2_1 _37162_ (.Y(_06574_),
    .A(net5805),
    .B(_06573_));
 sg13g2_nor2_1 _37163_ (.A(_06565_),
    .B(_06574_),
    .Y(_06575_));
 sg13g2_a21oi_1 _37164_ (.A1(_04564_),
    .A2(_06530_),
    .Y(_06576_),
    .B1(_04438_));
 sg13g2_a21oi_1 _37165_ (.A1(\u_inv.d_next[146] ),
    .A2(\u_inv.d_reg[146] ),
    .Y(_06577_),
    .B1(_06576_));
 sg13g2_a21oi_1 _37166_ (.A1(_04437_),
    .A2(_06577_),
    .Y(_06578_),
    .B1(net7214));
 sg13g2_o21ai_1 _37167_ (.B1(_06578_),
    .Y(_06579_),
    .A1(_04437_),
    .A2(_06577_));
 sg13g2_a21oi_1 _37168_ (.A1(net7214),
    .A2(\u_inv.d_next[147] ),
    .Y(_06580_),
    .B1(net6326));
 sg13g2_o21ai_1 _37169_ (.B1(_05254_),
    .Y(_06581_),
    .A1(_05187_),
    .A2(_06538_));
 sg13g2_a21oi_1 _37170_ (.A1(_04438_),
    .A2(_06581_),
    .Y(_06582_),
    .B1(_05256_));
 sg13g2_nand2b_1 _37171_ (.Y(_06583_),
    .B(_04436_),
    .A_N(_06582_));
 sg13g2_a21oi_1 _37172_ (.A1(_04437_),
    .A2(_06582_),
    .Y(_06584_),
    .B1(net6239));
 sg13g2_a22oi_1 _37173_ (.Y(_06585_),
    .B1(_06583_),
    .B2(_06584_),
    .A2(_06580_),
    .A1(_06579_));
 sg13g2_nand2_1 _37174_ (.Y(_06586_),
    .A(net5806),
    .B(_06585_));
 sg13g2_xnor2_1 _37175_ (.Y(_06587_),
    .A(net5856),
    .B(_06585_));
 sg13g2_xnor2_1 _37176_ (.Y(_06588_),
    .A(_04438_),
    .B(_06581_));
 sg13g2_nand3_1 _37177_ (.B(_04564_),
    .C(_06530_),
    .A(_04438_),
    .Y(_06589_));
 sg13g2_nand3b_1 _37178_ (.B(_06589_),
    .C(net7363),
    .Y(_06590_),
    .A_N(_06576_));
 sg13g2_a21oi_1 _37179_ (.A1(net7214),
    .A2(\u_inv.d_next[146] ),
    .Y(_06591_),
    .B1(net6326));
 sg13g2_a22oi_1 _37180_ (.Y(_06592_),
    .B1(_06590_),
    .B2(_06591_),
    .A2(_06588_),
    .A1(net6326));
 sg13g2_nand2_1 _37181_ (.Y(_06593_),
    .A(net5806),
    .B(_06592_));
 sg13g2_xnor2_1 _37182_ (.Y(_06594_),
    .A(net5856),
    .B(_06592_));
 sg13g2_nand3b_1 _37183_ (.B(_04443_),
    .C(_04445_),
    .Y(_06595_),
    .A_N(_06529_));
 sg13g2_nand4_1 _37184_ (.B(_04562_),
    .C(_06530_),
    .A(net7363),
    .Y(_06596_),
    .D(_06595_));
 sg13g2_a21oi_1 _37185_ (.A1(net7214),
    .A2(\u_inv.d_next[145] ),
    .Y(_06597_),
    .B1(net6326));
 sg13g2_o21ai_1 _37186_ (.B1(_05252_),
    .Y(_06598_),
    .A1(_04446_),
    .A2(_06538_));
 sg13g2_or2_1 _37187_ (.X(_06599_),
    .B(_06598_),
    .A(_04444_));
 sg13g2_a21oi_1 _37188_ (.A1(_04444_),
    .A2(_06598_),
    .Y(_06600_),
    .B1(net6239));
 sg13g2_a22oi_1 _37189_ (.Y(_06601_),
    .B1(_06599_),
    .B2(_06600_),
    .A2(_06597_),
    .A1(_06596_));
 sg13g2_nand2_1 _37190_ (.Y(_06602_),
    .A(net5805),
    .B(_06601_));
 sg13g2_xnor2_1 _37191_ (.Y(_06603_),
    .A(net5856),
    .B(_06601_));
 sg13g2_o21ai_1 _37192_ (.B1(net6326),
    .Y(_06604_),
    .A1(_04446_),
    .A2(_06538_));
 sg13g2_a21o_1 _37193_ (.A2(_06538_),
    .A1(_04446_),
    .B1(_06604_),
    .X(_06605_));
 sg13g2_nand3_1 _37194_ (.B(_04550_),
    .C(_06528_),
    .A(_04447_),
    .Y(_06606_));
 sg13g2_nor2_1 _37195_ (.A(net7214),
    .B(_06529_),
    .Y(_06607_));
 sg13g2_a22oi_1 _37196_ (.Y(_06608_),
    .B1(_06606_),
    .B2(_06607_),
    .A2(\u_inv.d_next[144] ),
    .A1(net7214));
 sg13g2_o21ai_1 _37197_ (.B1(_06605_),
    .Y(_06609_),
    .A1(net6326),
    .A2(_06608_));
 sg13g2_nand2_1 _37198_ (.Y(_06610_),
    .A(net5806),
    .B(_06609_));
 sg13g2_xnor2_1 _37199_ (.Y(_06611_),
    .A(net5856),
    .B(_06609_));
 sg13g2_nand4_1 _37200_ (.B(_06594_),
    .C(_06603_),
    .A(_06587_),
    .Y(_06612_),
    .D(_06611_));
 sg13g2_inv_1 _37201_ (.Y(_06613_),
    .A(_06612_));
 sg13g2_nand4_1 _37202_ (.B(_06555_),
    .C(_06575_),
    .A(_06547_),
    .Y(_06614_),
    .D(_06613_));
 sg13g2_a21oi_1 _37203_ (.A1(_04550_),
    .A2(_06528_),
    .Y(_06615_),
    .B1(_04449_));
 sg13g2_or2_1 _37204_ (.X(_06616_),
    .B(_06615_),
    .A(_04573_));
 sg13g2_o21ai_1 _37205_ (.B1(_04473_),
    .Y(_06617_),
    .A1(_04573_),
    .A2(_06615_));
 sg13g2_and2_1 _37206_ (.A(_04552_),
    .B(_06617_),
    .X(_06618_));
 sg13g2_a21oi_1 _37207_ (.A1(_04552_),
    .A2(_06617_),
    .Y(_06619_),
    .B1(_04467_));
 sg13g2_o21ai_1 _37208_ (.B1(_04459_),
    .Y(_06620_),
    .A1(_04554_),
    .A2(_06619_));
 sg13g2_nand3_1 _37209_ (.B(_04558_),
    .C(_06620_),
    .A(_04451_),
    .Y(_06621_));
 sg13g2_a21o_1 _37210_ (.A2(_06620_),
    .A1(_04558_),
    .B1(_04451_),
    .X(_06622_));
 sg13g2_a21oi_1 _37211_ (.A1(_06621_),
    .A2(_06622_),
    .Y(_06623_),
    .B1(net7207));
 sg13g2_o21ai_1 _37212_ (.B1(net6228),
    .Y(_06624_),
    .A1(net7349),
    .A2(\u_inv.d_next[158] ));
 sg13g2_nor2_1 _37213_ (.A(_06623_),
    .B(_06624_),
    .Y(_06625_));
 sg13g2_o21ai_1 _37214_ (.B1(_05267_),
    .Y(_06626_),
    .A1(_05190_),
    .A2(_06538_));
 sg13g2_nand3b_1 _37215_ (.B(_05181_),
    .C(_06626_),
    .Y(_06627_),
    .A_N(_05180_));
 sg13g2_a21oi_1 _37216_ (.A1(_05245_),
    .A2(_06627_),
    .Y(_06628_),
    .B1(_05177_));
 sg13g2_nor3_1 _37217_ (.A(_04451_),
    .B(_05250_),
    .C(_06628_),
    .Y(_06629_));
 sg13g2_o21ai_1 _37218_ (.B1(_04451_),
    .Y(_06630_),
    .A1(_05250_),
    .A2(_06628_));
 sg13g2_nor2b_1 _37219_ (.A(_06629_),
    .B_N(_06630_),
    .Y(_06631_));
 sg13g2_a21oi_2 _37220_ (.B1(_06625_),
    .Y(_06632_),
    .A2(_06631_),
    .A1(net6315));
 sg13g2_or2_1 _37221_ (.X(_06633_),
    .B(_06632_),
    .A(net5855));
 sg13g2_xnor2_1 _37222_ (.Y(_06634_),
    .A(net5804),
    .B(_06632_));
 sg13g2_xnor2_1 _37223_ (.Y(_06635_),
    .A(net5855),
    .B(_06632_));
 sg13g2_a21o_1 _37224_ (.A2(_06630_),
    .A1(_05247_),
    .B1(_04452_),
    .X(_06636_));
 sg13g2_nand3_1 _37225_ (.B(_05247_),
    .C(_06630_),
    .A(_04452_),
    .Y(_06637_));
 sg13g2_nand3_1 _37226_ (.B(_06636_),
    .C(_06637_),
    .A(net6316),
    .Y(_06638_));
 sg13g2_nand3_1 _37227_ (.B(_04452_),
    .C(_06622_),
    .A(_04450_),
    .Y(_06639_));
 sg13g2_a21o_1 _37228_ (.A2(_06622_),
    .A1(_04450_),
    .B1(_04452_),
    .X(_06640_));
 sg13g2_nand3_1 _37229_ (.B(_06639_),
    .C(_06640_),
    .A(net7349),
    .Y(_06641_));
 sg13g2_nand2_1 _37230_ (.Y(_06642_),
    .A(net7207),
    .B(\u_inv.d_next[159] ));
 sg13g2_nand3_1 _37231_ (.B(_06641_),
    .C(_06642_),
    .A(net6228),
    .Y(_06643_));
 sg13g2_nand2_1 _37232_ (.Y(_06644_),
    .A(_06638_),
    .B(_06643_));
 sg13g2_nand3_1 _37233_ (.B(_06638_),
    .C(_06643_),
    .A(net5804),
    .Y(_06645_));
 sg13g2_a21oi_1 _37234_ (.A1(_06638_),
    .A2(_06643_),
    .Y(_06646_),
    .B1(net5804));
 sg13g2_xnor2_1 _37235_ (.Y(_06647_),
    .A(net5855),
    .B(_06644_));
 sg13g2_nor2_1 _37236_ (.A(_06635_),
    .B(_06647_),
    .Y(_06648_));
 sg13g2_nand3b_1 _37237_ (.B(_06634_),
    .C(_06645_),
    .Y(_06649_),
    .A_N(_06646_));
 sg13g2_a21oi_1 _37238_ (.A1(_05245_),
    .A2(_06627_),
    .Y(_06650_),
    .B1(_04458_));
 sg13g2_o21ai_1 _37239_ (.B1(_04455_),
    .Y(_06651_),
    .A1(_05248_),
    .A2(_06650_));
 sg13g2_nor3_1 _37240_ (.A(_04455_),
    .B(_05248_),
    .C(_06650_),
    .Y(_06652_));
 sg13g2_nand2_1 _37241_ (.Y(_06653_),
    .A(net6316),
    .B(_06651_));
 sg13g2_o21ai_1 _37242_ (.B1(_04458_),
    .Y(_06654_),
    .A1(_04554_),
    .A2(_06619_));
 sg13g2_a21o_1 _37243_ (.A2(_06654_),
    .A1(_04457_),
    .B1(_04456_),
    .X(_06655_));
 sg13g2_nand3_1 _37244_ (.B(_04457_),
    .C(_06654_),
    .A(_04456_),
    .Y(_06656_));
 sg13g2_nand3_1 _37245_ (.B(_06655_),
    .C(_06656_),
    .A(net7349),
    .Y(_06657_));
 sg13g2_nand2_1 _37246_ (.Y(_06658_),
    .A(net7208),
    .B(\u_inv.d_next[157] ));
 sg13g2_nand3_1 _37247_ (.B(_06657_),
    .C(_06658_),
    .A(net6228),
    .Y(_06659_));
 sg13g2_o21ai_1 _37248_ (.B1(_06659_),
    .Y(_06660_),
    .A1(_06652_),
    .A2(_06653_));
 sg13g2_xnor2_1 _37249_ (.Y(_06661_),
    .A(net5855),
    .B(_06660_));
 sg13g2_nand3_1 _37250_ (.B(_05245_),
    .C(_06627_),
    .A(_04458_),
    .Y(_06662_));
 sg13g2_nor2b_1 _37251_ (.A(_06650_),
    .B_N(_06662_),
    .Y(_06663_));
 sg13g2_nor3_1 _37252_ (.A(_04458_),
    .B(_04554_),
    .C(_06619_),
    .Y(_06664_));
 sg13g2_nand2_1 _37253_ (.Y(_06665_),
    .A(net7349),
    .B(_06654_));
 sg13g2_a21oi_1 _37254_ (.A1(net7208),
    .A2(\u_inv.d_next[156] ),
    .Y(_06666_),
    .B1(net6316));
 sg13g2_o21ai_1 _37255_ (.B1(_06666_),
    .Y(_06667_),
    .A1(_06664_),
    .A2(_06665_));
 sg13g2_o21ai_1 _37256_ (.B1(_06667_),
    .Y(_06668_),
    .A1(net6230),
    .A2(_06663_));
 sg13g2_nor2_1 _37257_ (.A(net5855),
    .B(_06668_),
    .Y(_06669_));
 sg13g2_xnor2_1 _37258_ (.Y(_06670_),
    .A(net5855),
    .B(_06668_));
 sg13g2_inv_1 _37259_ (.Y(_06671_),
    .A(_06670_));
 sg13g2_nor2_1 _37260_ (.A(_06661_),
    .B(_06670_),
    .Y(_06672_));
 sg13g2_nand2b_1 _37261_ (.Y(_06673_),
    .B(_06671_),
    .A_N(_06661_));
 sg13g2_nor2_1 _37262_ (.A(_06649_),
    .B(_06673_),
    .Y(_06674_));
 sg13g2_a21oi_1 _37263_ (.A1(_05181_),
    .A2(_06626_),
    .Y(_06675_),
    .B1(_05241_));
 sg13g2_o21ai_1 _37264_ (.B1(_05242_),
    .Y(_06676_),
    .A1(_04466_),
    .A2(_06675_));
 sg13g2_nand2b_1 _37265_ (.Y(_06677_),
    .B(_04464_),
    .A_N(_06676_));
 sg13g2_a21oi_1 _37266_ (.A1(_04463_),
    .A2(_06676_),
    .Y(_06678_),
    .B1(net6239));
 sg13g2_nand2b_1 _37267_ (.Y(_06679_),
    .B(_04466_),
    .A_N(_06618_));
 sg13g2_a21oi_1 _37268_ (.A1(_04465_),
    .A2(_06679_),
    .Y(_06680_),
    .B1(_04464_));
 sg13g2_nand3_1 _37269_ (.B(_04465_),
    .C(_06679_),
    .A(_04464_),
    .Y(_06681_));
 sg13g2_nand3b_1 _37270_ (.B(_06681_),
    .C(net7363),
    .Y(_06682_),
    .A_N(_06680_));
 sg13g2_a21oi_1 _37271_ (.A1(net7215),
    .A2(\u_inv.d_next[155] ),
    .Y(_06683_),
    .B1(net6325));
 sg13g2_a22oi_1 _37272_ (.Y(_06684_),
    .B1(_06682_),
    .B2(_06683_),
    .A2(_06678_),
    .A1(_06677_));
 sg13g2_xnor2_1 _37273_ (.Y(_06685_),
    .A(net5804),
    .B(_06684_));
 sg13g2_nand2b_1 _37274_ (.Y(_06686_),
    .B(_06618_),
    .A_N(_04466_));
 sg13g2_nand3_1 _37275_ (.B(_06679_),
    .C(_06686_),
    .A(net7363),
    .Y(_06687_));
 sg13g2_xnor2_1 _37276_ (.Y(_06688_),
    .A(_04466_),
    .B(_06675_));
 sg13g2_a21oi_1 _37277_ (.A1(net7215),
    .A2(\u_inv.d_next[154] ),
    .Y(_06689_),
    .B1(net6325));
 sg13g2_a22oi_1 _37278_ (.Y(_06690_),
    .B1(_06689_),
    .B2(_06687_),
    .A2(_06688_),
    .A1(net6325));
 sg13g2_nand2_1 _37279_ (.Y(_06691_),
    .A(net5804),
    .B(_06690_));
 sg13g2_xnor2_1 _37280_ (.Y(_06692_),
    .A(net5804),
    .B(_06690_));
 sg13g2_or2_1 _37281_ (.X(_06693_),
    .B(_06692_),
    .A(_06685_));
 sg13g2_nand2b_1 _37282_ (.Y(_06694_),
    .B(_04472_),
    .A_N(_06616_));
 sg13g2_nand2b_1 _37283_ (.Y(_06695_),
    .B(_06616_),
    .A_N(_04472_));
 sg13g2_nand3_1 _37284_ (.B(_06694_),
    .C(_06695_),
    .A(net7363),
    .Y(_06696_));
 sg13g2_xnor2_1 _37285_ (.Y(_06697_),
    .A(_04472_),
    .B(_06626_));
 sg13g2_a21oi_1 _37286_ (.A1(net7215),
    .A2(\u_inv.d_next[152] ),
    .Y(_06698_),
    .B1(net6325));
 sg13g2_a22oi_1 _37287_ (.Y(_06699_),
    .B1(_06698_),
    .B2(_06696_),
    .A2(_06697_),
    .A1(net6325));
 sg13g2_nand2_1 _37288_ (.Y(_06700_),
    .A(net5807),
    .B(_06699_));
 sg13g2_xnor2_1 _37289_ (.Y(_06701_),
    .A(net5855),
    .B(_06699_));
 sg13g2_inv_1 _37290_ (.Y(_06702_),
    .A(_06701_));
 sg13g2_a21oi_1 _37291_ (.A1(_04471_),
    .A2(_06695_),
    .Y(_06703_),
    .B1(_04470_));
 sg13g2_nand3_1 _37292_ (.B(_04471_),
    .C(_06695_),
    .A(_04470_),
    .Y(_06704_));
 sg13g2_nor2_1 _37293_ (.A(net7215),
    .B(_06703_),
    .Y(_06705_));
 sg13g2_a221oi_1 _37294_ (.B2(_06705_),
    .C1(net6325),
    .B1(_06704_),
    .A1(net7215),
    .Y(_06706_),
    .A2(\u_inv.d_next[153] ));
 sg13g2_a21oi_1 _37295_ (.A1(_04472_),
    .A2(_06626_),
    .Y(_06707_),
    .B1(_05238_));
 sg13g2_xor2_1 _37296_ (.B(_06707_),
    .A(_04470_),
    .X(_06708_));
 sg13g2_a21o_2 _37297_ (.A2(_06708_),
    .A1(net6325),
    .B1(_06706_),
    .X(_06709_));
 sg13g2_nor2_1 _37298_ (.A(net5856),
    .B(_06709_),
    .Y(_06710_));
 sg13g2_xnor2_1 _37299_ (.Y(_06711_),
    .A(net5807),
    .B(_06709_));
 sg13g2_and2_1 _37300_ (.A(_06701_),
    .B(_06711_),
    .X(_06712_));
 sg13g2_nand2b_1 _37301_ (.Y(_06713_),
    .B(_06712_),
    .A_N(_06693_));
 sg13g2_nor3_1 _37302_ (.A(_06649_),
    .B(_06673_),
    .C(_06713_),
    .Y(_06714_));
 sg13g2_nor4_1 _37303_ (.A(_06614_),
    .B(_06649_),
    .C(_06673_),
    .D(_06713_),
    .Y(_06715_));
 sg13g2_nand2b_2 _37304_ (.Y(_06716_),
    .B(_06527_),
    .A_N(_04530_));
 sg13g2_nand2b_1 _37305_ (.Y(_06717_),
    .B(_06716_),
    .A_N(_04507_));
 sg13g2_nand2_1 _37306_ (.Y(_06718_),
    .A(_04532_),
    .B(_06717_));
 sg13g2_nand2_1 _37307_ (.Y(_06719_),
    .A(_04500_),
    .B(_06718_));
 sg13g2_xnor2_1 _37308_ (.Y(_06720_),
    .A(_04500_),
    .B(_06718_));
 sg13g2_o21ai_1 _37309_ (.B1(net6247),
    .Y(_06721_),
    .A1(net7374),
    .A2(\u_inv.d_next[134] ));
 sg13g2_a21oi_1 _37310_ (.A1(net7374),
    .A2(_06720_),
    .Y(_06722_),
    .B1(_06721_));
 sg13g2_a21oi_1 _37311_ (.A1(_05148_),
    .A2(_05202_),
    .Y(_06723_),
    .B1(_05209_));
 sg13g2_o21ai_1 _37312_ (.B1(_05213_),
    .Y(_06724_),
    .A1(_05201_),
    .A2(_06723_));
 sg13g2_a21oi_1 _37313_ (.A1(_05197_),
    .A2(_06724_),
    .Y(_06725_),
    .B1(_05217_));
 sg13g2_xnor2_1 _37314_ (.Y(_06726_),
    .A(_04501_),
    .B(_06725_));
 sg13g2_a21oi_1 _37315_ (.A1(net6342),
    .A2(_06726_),
    .Y(_06727_),
    .B1(_06722_));
 sg13g2_nor2_1 _37316_ (.A(net5862),
    .B(_06727_),
    .Y(_06728_));
 sg13g2_nand2_1 _37317_ (.Y(_06729_),
    .A(net5862),
    .B(_06727_));
 sg13g2_nand2b_1 _37318_ (.Y(_06730_),
    .B(_06729_),
    .A_N(_06728_));
 sg13g2_o21ai_1 _37319_ (.B1(_05218_),
    .Y(_06731_),
    .A1(_04500_),
    .A2(_06725_));
 sg13g2_nand2b_1 _37320_ (.Y(_06732_),
    .B(_04498_),
    .A_N(_06731_));
 sg13g2_a21oi_1 _37321_ (.A1(_04497_),
    .A2(_06731_),
    .Y(_06733_),
    .B1(net6247));
 sg13g2_a21o_1 _37322_ (.A2(_06719_),
    .A1(_04499_),
    .B1(_04498_),
    .X(_06734_));
 sg13g2_nand3_1 _37323_ (.B(_04499_),
    .C(_06719_),
    .A(_04498_),
    .Y(_06735_));
 sg13g2_nand3_1 _37324_ (.B(_06734_),
    .C(_06735_),
    .A(net7374),
    .Y(_06736_));
 sg13g2_a21oi_1 _37325_ (.A1(net7222),
    .A2(\u_inv.d_next[135] ),
    .Y(_06737_),
    .B1(net6337));
 sg13g2_a22oi_1 _37326_ (.Y(_06738_),
    .B1(_06736_),
    .B2(_06737_),
    .A2(_06733_),
    .A1(_06732_));
 sg13g2_xnor2_1 _37327_ (.Y(_06739_),
    .A(net5814),
    .B(_06738_));
 sg13g2_nor2_1 _37328_ (.A(_06730_),
    .B(_06739_),
    .Y(_06740_));
 sg13g2_xnor2_1 _37329_ (.Y(_06741_),
    .A(_04505_),
    .B(_06716_));
 sg13g2_o21ai_1 _37330_ (.B1(net6248),
    .Y(_06742_),
    .A1(net7374),
    .A2(\u_inv.d_next[132] ));
 sg13g2_a21oi_1 _37331_ (.A1(net7374),
    .A2(_06741_),
    .Y(_06743_),
    .B1(_06742_));
 sg13g2_xnor2_1 _37332_ (.Y(_06744_),
    .A(_04505_),
    .B(_06724_));
 sg13g2_a21oi_2 _37333_ (.B1(_06743_),
    .Y(_06745_),
    .A2(_06744_),
    .A1(net6337));
 sg13g2_a21oi_1 _37334_ (.A1(_04505_),
    .A2(_06716_),
    .Y(_06746_),
    .B1(_04503_));
 sg13g2_nand2b_1 _37335_ (.Y(_06747_),
    .B(_06746_),
    .A_N(_04504_));
 sg13g2_a21oi_1 _37336_ (.A1(_04503_),
    .A2(_04504_),
    .Y(_06748_),
    .B1(net7222));
 sg13g2_nand3_1 _37337_ (.B(_06747_),
    .C(_06748_),
    .A(_06717_),
    .Y(_06749_));
 sg13g2_a21oi_1 _37338_ (.A1(net7222),
    .A2(\u_inv.d_next[133] ),
    .Y(_06750_),
    .B1(net6342));
 sg13g2_a21oi_1 _37339_ (.A1(_04506_),
    .A2(_06724_),
    .Y(_06751_),
    .B1(_05215_));
 sg13g2_or2_1 _37340_ (.X(_06752_),
    .B(_06751_),
    .A(_04502_));
 sg13g2_a21oi_1 _37341_ (.A1(_04502_),
    .A2(_06751_),
    .Y(_06753_),
    .B1(net6248));
 sg13g2_a22oi_1 _37342_ (.Y(_06754_),
    .B1(_06752_),
    .B2(_06753_),
    .A2(_06750_),
    .A1(_06749_));
 sg13g2_inv_1 _37343_ (.Y(_06755_),
    .A(_06754_));
 sg13g2_a21o_1 _37344_ (.A2(_06755_),
    .A1(_06745_),
    .B1(net5862),
    .X(_06756_));
 sg13g2_xnor2_1 _37345_ (.Y(_06757_),
    .A(net5862),
    .B(_06745_));
 sg13g2_xnor2_1 _37346_ (.Y(_06758_),
    .A(net5814),
    .B(_06754_));
 sg13g2_or2_1 _37347_ (.X(_06759_),
    .B(_06758_),
    .A(_06757_));
 sg13g2_a21o_1 _37348_ (.A2(_06526_),
    .A1(_04528_),
    .B1(_04511_),
    .X(_06760_));
 sg13g2_a21oi_1 _37349_ (.A1(_04509_),
    .A2(_06760_),
    .Y(_06761_),
    .B1(_04512_));
 sg13g2_nand3_1 _37350_ (.B(_04512_),
    .C(_06760_),
    .A(_04509_),
    .Y(_06762_));
 sg13g2_nor2_1 _37351_ (.A(net7221),
    .B(_06761_),
    .Y(_06763_));
 sg13g2_a221oi_1 _37352_ (.B2(_06763_),
    .C1(net6337),
    .B1(_06762_),
    .A1(net7222),
    .Y(_06764_),
    .A2(\u_inv.d_next[131] ));
 sg13g2_o21ai_1 _37353_ (.B1(_05211_),
    .Y(_06765_),
    .A1(_04510_),
    .A2(_06723_));
 sg13g2_xnor2_1 _37354_ (.Y(_06766_),
    .A(_04512_),
    .B(_06765_));
 sg13g2_a21o_2 _37355_ (.A2(_06766_),
    .A1(net6337),
    .B1(_06764_),
    .X(_06767_));
 sg13g2_nor2_1 _37356_ (.A(net5862),
    .B(_06767_),
    .Y(_06768_));
 sg13g2_xnor2_1 _37357_ (.Y(_06769_),
    .A(net5864),
    .B(_06767_));
 sg13g2_xnor2_1 _37358_ (.Y(_06770_),
    .A(_04510_),
    .B(_06723_));
 sg13g2_nand3_1 _37359_ (.B(_04528_),
    .C(_06526_),
    .A(_04511_),
    .Y(_06771_));
 sg13g2_nand3_1 _37360_ (.B(_06760_),
    .C(_06771_),
    .A(net7376),
    .Y(_06772_));
 sg13g2_a21oi_1 _37361_ (.A1(net7222),
    .A2(net7296),
    .Y(_06773_),
    .B1(net6337));
 sg13g2_a22oi_1 _37362_ (.Y(_06774_),
    .B1(_06772_),
    .B2(_06773_),
    .A2(_06770_),
    .A1(net6337));
 sg13g2_and2_1 _37363_ (.A(net5814),
    .B(_06774_),
    .X(_06775_));
 sg13g2_xnor2_1 _37364_ (.Y(_06776_),
    .A(net5862),
    .B(_06774_));
 sg13g2_inv_1 _37365_ (.Y(_06777_),
    .A(_06776_));
 sg13g2_nand3_1 _37366_ (.B(_04520_),
    .C(_06525_),
    .A(_04516_),
    .Y(_06778_));
 sg13g2_nor2_1 _37367_ (.A(net7225),
    .B(_04527_),
    .Y(_06779_));
 sg13g2_nand3_1 _37368_ (.B(_06778_),
    .C(_06779_),
    .A(_06526_),
    .Y(_06780_));
 sg13g2_a21oi_1 _37369_ (.A1(net7225),
    .A2(\u_inv.d_next[129] ),
    .Y(_06781_),
    .B1(net6341));
 sg13g2_o21ai_1 _37370_ (.B1(_05208_),
    .Y(_06782_),
    .A1(net6994),
    .A2(net1104));
 sg13g2_xnor2_1 _37371_ (.Y(_06783_),
    .A(_04516_),
    .B(_06782_));
 sg13g2_a22oi_1 _37372_ (.Y(_06784_),
    .B1(_06783_),
    .B2(net6341),
    .A2(_06781_),
    .A1(_06780_));
 sg13g2_inv_1 _37373_ (.Y(_06785_),
    .A(_06784_));
 sg13g2_a21oi_1 _37374_ (.A1(net1109),
    .A2(_04522_),
    .Y(_06786_),
    .B1(net7225));
 sg13g2_xnor2_1 _37375_ (.Y(_06787_),
    .A(net6994),
    .B(net1104));
 sg13g2_a221oi_1 _37376_ (.B2(_06786_),
    .C1(net6341),
    .B1(_06525_),
    .A1(net7225),
    .Y(_06788_),
    .A2(\u_inv.d_next[128] ));
 sg13g2_a21oi_2 _37377_ (.B1(_06788_),
    .Y(_06789_),
    .A2(_06787_),
    .A1(net6341));
 sg13g2_nand2_1 _37378_ (.Y(_06790_),
    .A(net5819),
    .B(_06789_));
 sg13g2_o21ai_1 _37379_ (.B1(net5819),
    .Y(_06791_),
    .A1(_06784_),
    .A2(_06789_));
 sg13g2_nor3_1 _37380_ (.A(_06769_),
    .B(_06777_),
    .C(_06791_),
    .Y(_06792_));
 sg13g2_nor3_1 _37381_ (.A(_06768_),
    .B(_06775_),
    .C(_06792_),
    .Y(_06793_));
 sg13g2_o21ai_1 _37382_ (.B1(_06756_),
    .Y(_06794_),
    .A1(_06759_),
    .A2(_06793_));
 sg13g2_a221oi_1 _37383_ (.B2(_06794_),
    .C1(_06728_),
    .B1(_06740_),
    .A1(net5814),
    .Y(_06795_),
    .A2(_06738_));
 sg13g2_o21ai_1 _37384_ (.B1(_05221_),
    .Y(_06796_),
    .A1(net1104),
    .A2(_05203_));
 sg13g2_a21oi_1 _37385_ (.A1(_05194_),
    .A2(_06796_),
    .Y(_06797_),
    .B1(_05233_));
 sg13g2_a21o_2 _37386_ (.A2(_06796_),
    .A1(_05194_),
    .B1(_05233_),
    .X(_06798_));
 sg13g2_a21oi_1 _37387_ (.A1(_05195_),
    .A2(_06798_),
    .Y(_06799_),
    .B1(_05230_));
 sg13g2_a21o_1 _37388_ (.A2(_06798_),
    .A1(_05195_),
    .B1(_05230_),
    .X(_06800_));
 sg13g2_a21oi_1 _37389_ (.A1(_05192_),
    .A2(_06800_),
    .Y(_06801_),
    .B1(_05224_));
 sg13g2_xnor2_1 _37390_ (.Y(_06802_),
    .A(_04479_),
    .B(_06801_));
 sg13g2_a21oi_1 _37391_ (.A1(_04422_),
    .A2(_04523_),
    .Y(_06803_),
    .B1(_04536_));
 sg13g2_or2_1 _37392_ (.X(_06804_),
    .B(_06803_),
    .A(_04493_));
 sg13g2_o21ai_1 _37393_ (.B1(_04543_),
    .Y(_06805_),
    .A1(_04491_),
    .A2(_06804_));
 sg13g2_a21o_2 _37394_ (.A2(_06805_),
    .A1(_04489_),
    .B1(_04547_),
    .X(_06806_));
 sg13g2_a21oi_1 _37395_ (.A1(_04483_),
    .A2(_06806_),
    .Y(_06807_),
    .B1(_04539_));
 sg13g2_xnor2_1 _37396_ (.Y(_06808_),
    .A(_04479_),
    .B(_06807_));
 sg13g2_nand2_1 _37397_ (.Y(_06809_),
    .A(net7364),
    .B(_06808_));
 sg13g2_a21oi_1 _37398_ (.A1(net7216),
    .A2(\u_inv.d_next[142] ),
    .Y(_06810_),
    .B1(net6328));
 sg13g2_a22oi_1 _37399_ (.Y(_06811_),
    .B1(_06809_),
    .B2(_06810_),
    .A2(_06802_),
    .A1(net6328));
 sg13g2_nand2_1 _37400_ (.Y(_06812_),
    .A(net5813),
    .B(_06811_));
 sg13g2_xnor2_1 _37401_ (.Y(_06813_),
    .A(net5863),
    .B(_06811_));
 sg13g2_o21ai_1 _37402_ (.B1(_04477_),
    .Y(_06814_),
    .A1(_04478_),
    .A2(_06807_));
 sg13g2_a21oi_1 _37403_ (.A1(_04476_),
    .A2(_06814_),
    .Y(_06815_),
    .B1(net7217));
 sg13g2_o21ai_1 _37404_ (.B1(_06815_),
    .Y(_06816_),
    .A1(_04476_),
    .A2(_06814_));
 sg13g2_a21oi_1 _37405_ (.A1(net7217),
    .A2(\u_inv.d_next[143] ),
    .Y(_06817_),
    .B1(net6329));
 sg13g2_o21ai_1 _37406_ (.B1(_05226_),
    .Y(_06818_),
    .A1(_04479_),
    .A2(_06801_));
 sg13g2_or2_1 _37407_ (.X(_06819_),
    .B(_06818_),
    .A(_04476_));
 sg13g2_a21oi_1 _37408_ (.A1(_04476_),
    .A2(_06818_),
    .Y(_06820_),
    .B1(net6239));
 sg13g2_a22oi_1 _37409_ (.Y(_06821_),
    .B1(_06819_),
    .B2(_06820_),
    .A2(_06817_),
    .A1(_06816_));
 sg13g2_nand2_1 _37410_ (.Y(_06822_),
    .A(net5814),
    .B(_06821_));
 sg13g2_xnor2_1 _37411_ (.Y(_06823_),
    .A(net5863),
    .B(_06821_));
 sg13g2_a21oi_1 _37412_ (.A1(_04482_),
    .A2(_06806_),
    .Y(_06824_),
    .B1(_04481_));
 sg13g2_xnor2_1 _37413_ (.Y(_06825_),
    .A(_04480_),
    .B(_06824_));
 sg13g2_nand2_1 _37414_ (.Y(_06826_),
    .A(net7216),
    .B(\u_inv.d_next[141] ));
 sg13g2_a21oi_1 _37415_ (.A1(net7364),
    .A2(_06825_),
    .Y(_06827_),
    .B1(net6328));
 sg13g2_o21ai_1 _37416_ (.B1(_05222_),
    .Y(_06828_),
    .A1(_04482_),
    .A2(_06799_));
 sg13g2_or2_1 _37417_ (.X(_06829_),
    .B(_06828_),
    .A(_04480_));
 sg13g2_a21oi_1 _37418_ (.A1(_04480_),
    .A2(_06828_),
    .Y(_06830_),
    .B1(net6239));
 sg13g2_a22oi_1 _37419_ (.Y(_06831_),
    .B1(_06829_),
    .B2(_06830_),
    .A2(_06827_),
    .A1(_06826_));
 sg13g2_nand2_1 _37420_ (.Y(_06832_),
    .A(net5813),
    .B(_06831_));
 sg13g2_xnor2_1 _37421_ (.Y(_06833_),
    .A(net5863),
    .B(_06831_));
 sg13g2_xnor2_1 _37422_ (.Y(_06834_),
    .A(_04482_),
    .B(_06799_));
 sg13g2_a21oi_1 _37423_ (.A1(_04482_),
    .A2(_06806_),
    .Y(_06835_),
    .B1(net7216));
 sg13g2_o21ai_1 _37424_ (.B1(_06835_),
    .Y(_06836_),
    .A1(_04482_),
    .A2(_06806_));
 sg13g2_a21oi_1 _37425_ (.A1(net7216),
    .A2(\u_inv.d_next[140] ),
    .Y(_06837_),
    .B1(net6328));
 sg13g2_a22oi_1 _37426_ (.Y(_06838_),
    .B1(_06836_),
    .B2(_06837_),
    .A2(_06834_),
    .A1(net6328));
 sg13g2_nand2_1 _37427_ (.Y(_06839_),
    .A(net5813),
    .B(_06838_));
 sg13g2_xnor2_1 _37428_ (.Y(_06840_),
    .A(net5863),
    .B(_06838_));
 sg13g2_inv_1 _37429_ (.Y(_06841_),
    .A(_06840_));
 sg13g2_and2_1 _37430_ (.A(_06833_),
    .B(_06840_),
    .X(_06842_));
 sg13g2_inv_1 _37431_ (.Y(_06843_),
    .A(_06842_));
 sg13g2_nand3_1 _37432_ (.B(_06823_),
    .C(_06842_),
    .A(_06813_),
    .Y(_06844_));
 sg13g2_a21oi_1 _37433_ (.A1(_04488_),
    .A2(_06805_),
    .Y(_06845_),
    .B1(_04487_));
 sg13g2_nand2b_1 _37434_ (.Y(_06846_),
    .B(_04485_),
    .A_N(_06845_));
 sg13g2_a21oi_1 _37435_ (.A1(_04486_),
    .A2(_06845_),
    .Y(_06847_),
    .B1(net7216));
 sg13g2_nand2_1 _37436_ (.Y(_06848_),
    .A(net7216),
    .B(\u_inv.d_next[139] ));
 sg13g2_a21oi_1 _37437_ (.A1(_06846_),
    .A2(_06847_),
    .Y(_06849_),
    .B1(net6328));
 sg13g2_o21ai_1 _37438_ (.B1(_05228_),
    .Y(_06850_),
    .A1(_04488_),
    .A2(_06797_));
 sg13g2_nand2b_1 _37439_ (.Y(_06851_),
    .B(_04486_),
    .A_N(_06850_));
 sg13g2_a21oi_1 _37440_ (.A1(_04485_),
    .A2(_06850_),
    .Y(_06852_),
    .B1(net6240));
 sg13g2_a22oi_1 _37441_ (.Y(_06853_),
    .B1(_06851_),
    .B2(_06852_),
    .A2(_06849_),
    .A1(_06848_));
 sg13g2_nand2_1 _37442_ (.Y(_06854_),
    .A(net5813),
    .B(_06853_));
 sg13g2_xnor2_1 _37443_ (.Y(_06855_),
    .A(net5863),
    .B(_06853_));
 sg13g2_xnor2_1 _37444_ (.Y(_06856_),
    .A(_04488_),
    .B(_06798_));
 sg13g2_xnor2_1 _37445_ (.Y(_06857_),
    .A(_04488_),
    .B(_06805_));
 sg13g2_o21ai_1 _37446_ (.B1(net6240),
    .Y(_06858_),
    .A1(net7364),
    .A2(\u_inv.d_next[138] ));
 sg13g2_a21oi_1 _37447_ (.A1(net7364),
    .A2(_06857_),
    .Y(_06859_),
    .B1(_06858_));
 sg13g2_a21oi_1 _37448_ (.A1(net6328),
    .A2(_06856_),
    .Y(_06860_),
    .B1(_06859_));
 sg13g2_or2_1 _37449_ (.X(_06861_),
    .B(_06860_),
    .A(net5863));
 sg13g2_xnor2_1 _37450_ (.Y(_06862_),
    .A(net5813),
    .B(_06860_));
 sg13g2_inv_1 _37451_ (.Y(_06863_),
    .A(_06862_));
 sg13g2_nand2_1 _37452_ (.Y(_06864_),
    .A(_06855_),
    .B(_06862_));
 sg13g2_xnor2_1 _37453_ (.Y(_06865_),
    .A(_04493_),
    .B(_06796_));
 sg13g2_a21oi_1 _37454_ (.A1(_04493_),
    .A2(_06803_),
    .Y(_06866_),
    .B1(net7216));
 sg13g2_a221oi_1 _37455_ (.B2(_06866_),
    .C1(net6328),
    .B1(_06804_),
    .A1(net7216),
    .Y(_06867_),
    .A2(\u_inv.d_next[136] ));
 sg13g2_a21oi_2 _37456_ (.B1(_06867_),
    .Y(_06868_),
    .A2(_06865_),
    .A1(net6329));
 sg13g2_nand2_1 _37457_ (.Y(_06869_),
    .A(net5813),
    .B(_06868_));
 sg13g2_xnor2_1 _37458_ (.Y(_06870_),
    .A(net5863),
    .B(_06868_));
 sg13g2_and2_1 _37459_ (.A(_04491_),
    .B(_04492_),
    .X(_06871_));
 sg13g2_nor2_1 _37460_ (.A(net7217),
    .B(_04542_),
    .Y(_06872_));
 sg13g2_o21ai_1 _37461_ (.B1(_06872_),
    .Y(_06873_),
    .A1(_04491_),
    .A2(_06804_));
 sg13g2_a21o_1 _37462_ (.A2(_06871_),
    .A1(_06804_),
    .B1(_06873_),
    .X(_06874_));
 sg13g2_a21oi_1 _37463_ (.A1(_04493_),
    .A2(_06796_),
    .Y(_06875_),
    .B1(_05231_));
 sg13g2_o21ai_1 _37464_ (.B1(net6329),
    .Y(_06876_),
    .A1(_04491_),
    .A2(_06875_));
 sg13g2_a21oi_1 _37465_ (.A1(_04491_),
    .A2(_06875_),
    .Y(_06877_),
    .B1(_06876_));
 sg13g2_a21oi_1 _37466_ (.A1(net7217),
    .A2(\u_inv.d_next[137] ),
    .Y(_06878_),
    .B1(net6329));
 sg13g2_a21o_2 _37467_ (.A2(_06878_),
    .A1(_06874_),
    .B1(_06877_),
    .X(_06879_));
 sg13g2_xnor2_1 _37468_ (.Y(_06880_),
    .A(net5813),
    .B(_06879_));
 sg13g2_and2_1 _37469_ (.A(_06870_),
    .B(_06880_),
    .X(_06881_));
 sg13g2_inv_1 _37470_ (.Y(_06882_),
    .A(_06881_));
 sg13g2_nor4_2 _37471_ (.A(_06795_),
    .B(_06844_),
    .C(_06864_),
    .Y(_06883_),
    .D(_06882_));
 sg13g2_o21ai_1 _37472_ (.B1(_06869_),
    .Y(_06884_),
    .A1(net5863),
    .A2(_06879_));
 sg13g2_nand3_1 _37473_ (.B(_06862_),
    .C(_06884_),
    .A(_06855_),
    .Y(_06885_));
 sg13g2_nand3_1 _37474_ (.B(_06861_),
    .C(_06885_),
    .A(_06854_),
    .Y(_06886_));
 sg13g2_inv_1 _37475_ (.Y(_06887_),
    .A(_06886_));
 sg13g2_nand4_1 _37476_ (.B(_06823_),
    .C(_06842_),
    .A(_06813_),
    .Y(_06888_),
    .D(_06886_));
 sg13g2_nand2_1 _37477_ (.Y(_06889_),
    .A(_06832_),
    .B(_06839_));
 sg13g2_nand3_1 _37478_ (.B(_06823_),
    .C(_06889_),
    .A(_06813_),
    .Y(_06890_));
 sg13g2_nand4_1 _37479_ (.B(_06822_),
    .C(_06888_),
    .A(_06812_),
    .Y(_06891_),
    .D(_06890_));
 sg13g2_nand4_1 _37480_ (.B(_06823_),
    .C(_06842_),
    .A(_06813_),
    .Y(_06892_),
    .D(_06881_));
 sg13g2_nor2_1 _37481_ (.A(_06883_),
    .B(_06891_),
    .Y(_06893_));
 sg13g2_o21ai_1 _37482_ (.B1(_06715_),
    .Y(_06894_),
    .A1(_06883_),
    .A2(_06891_));
 sg13g2_a21oi_1 _37483_ (.A1(net5804),
    .A2(_06699_),
    .Y(_06895_),
    .B1(_06710_));
 sg13g2_o21ai_1 _37484_ (.B1(net5804),
    .Y(_06896_),
    .A1(_06684_),
    .A2(_06690_));
 sg13g2_o21ai_1 _37485_ (.B1(_06896_),
    .Y(_06897_),
    .A1(_06693_),
    .A2(_06895_));
 sg13g2_inv_1 _37486_ (.Y(_06898_),
    .A(_06897_));
 sg13g2_a21oi_1 _37487_ (.A1(_06660_),
    .A2(_06668_),
    .Y(_06899_),
    .B1(net5855));
 sg13g2_nand2_1 _37488_ (.Y(_06900_),
    .A(_06633_),
    .B(_06645_));
 sg13g2_a221oi_1 _37489_ (.B2(_06648_),
    .C1(_06900_),
    .B1(_06899_),
    .A1(_06674_),
    .Y(_06901_),
    .A2(_06897_));
 sg13g2_nand2_1 _37490_ (.Y(_06902_),
    .A(_06602_),
    .B(_06610_));
 sg13g2_nand3_1 _37491_ (.B(_06594_),
    .C(_06902_),
    .A(_06587_),
    .Y(_06903_));
 sg13g2_nand3_1 _37492_ (.B(_06593_),
    .C(_06903_),
    .A(_06586_),
    .Y(_06904_));
 sg13g2_nand4_1 _37493_ (.B(_06555_),
    .C(_06575_),
    .A(_06547_),
    .Y(_06905_),
    .D(_06904_));
 sg13g2_a21oi_1 _37494_ (.A1(net5805),
    .A2(_06546_),
    .Y(_06906_),
    .B1(_06554_));
 sg13g2_o21ai_1 _37495_ (.B1(net5805),
    .Y(_06907_),
    .A1(_06563_),
    .A2(_06573_));
 sg13g2_nand3b_1 _37496_ (.B(_06555_),
    .C(_06547_),
    .Y(_06908_),
    .A_N(_06907_));
 sg13g2_nand3_1 _37497_ (.B(_06906_),
    .C(_06908_),
    .A(_06905_),
    .Y(_06909_));
 sg13g2_nand2_1 _37498_ (.Y(_06910_),
    .A(_06714_),
    .B(_06909_));
 sg13g2_and3_2 _37499_ (.X(_06911_),
    .A(_06894_),
    .B(_06901_),
    .C(_06910_));
 sg13g2_nand3_1 _37500_ (.B(_06901_),
    .C(_06910_),
    .A(_06894_),
    .Y(_06912_));
 sg13g2_a21oi_1 _37501_ (.A1(net5798),
    .A2(_06511_),
    .Y(_06913_),
    .B1(_06522_));
 sg13g2_o21ai_1 _37502_ (.B1(net5797),
    .Y(_06914_),
    .A1(_06493_),
    .A2(_06503_));
 sg13g2_o21ai_1 _37503_ (.B1(_06914_),
    .Y(_06915_),
    .A1(_06506_),
    .A2(_06913_));
 sg13g2_inv_1 _37504_ (.Y(_06916_),
    .A(_06915_));
 sg13g2_nand2_1 _37505_ (.Y(_06917_),
    .A(_06458_),
    .B(_06465_));
 sg13g2_nand2_1 _37506_ (.Y(_06918_),
    .A(_06474_),
    .B(_06484_));
 sg13g2_a221oi_1 _37507_ (.B2(_06467_),
    .C1(_06917_),
    .B1(_06918_),
    .A1(_06487_),
    .Y(_06919_),
    .A2(_06915_));
 sg13g2_nand3b_1 _37508_ (.B(_06440_),
    .C(_06401_),
    .Y(_06920_),
    .A_N(_06919_));
 sg13g2_nand2_1 _37509_ (.Y(_06921_),
    .A(_06429_),
    .B(_06436_));
 sg13g2_nand2_1 _37510_ (.Y(_06922_),
    .A(_06411_),
    .B(_06418_));
 sg13g2_a21o_1 _37511_ (.A2(_06921_),
    .A1(_06420_),
    .B1(_06922_),
    .X(_06923_));
 sg13g2_nand2_1 _37512_ (.Y(_06924_),
    .A(_06401_),
    .B(_06923_));
 sg13g2_nor2_1 _37513_ (.A(_06368_),
    .B(_06378_),
    .Y(_06925_));
 sg13g2_a21oi_1 _37514_ (.A1(net5792),
    .A2(_06389_),
    .Y(_06926_),
    .B1(_06398_));
 sg13g2_or4_1 _37515_ (.A(_06369_),
    .B(_06378_),
    .C(_06379_),
    .D(_06926_),
    .X(_06927_));
 sg13g2_nand4_1 _37516_ (.B(_06924_),
    .C(_06925_),
    .A(_06920_),
    .Y(_06928_),
    .D(_06927_));
 sg13g2_a21o_1 _37517_ (.A2(_06252_),
    .A1(net5799),
    .B1(_06220_),
    .X(_06929_));
 sg13g2_nand3_1 _37518_ (.B(_06242_),
    .C(_06929_),
    .A(_06231_),
    .Y(_06930_));
 sg13g2_nand3_1 _37519_ (.B(_06241_),
    .C(_06930_),
    .A(_06230_),
    .Y(_06931_));
 sg13g2_inv_1 _37520_ (.Y(_06932_),
    .A(_06931_));
 sg13g2_nand2_1 _37521_ (.Y(_06933_),
    .A(_06184_),
    .B(_06194_));
 sg13g2_nand2_1 _37522_ (.Y(_06934_),
    .A(_06205_),
    .B(_06211_));
 sg13g2_a21oi_1 _37523_ (.A1(_06196_),
    .A2(_06934_),
    .Y(_06935_),
    .B1(_06933_));
 sg13g2_o21ai_1 _37524_ (.B1(_06935_),
    .Y(_06936_),
    .A1(_06214_),
    .A2(_06932_));
 sg13g2_nand4_1 _37525_ (.B(_06327_),
    .C(_06346_),
    .A(_06307_),
    .Y(_06937_),
    .D(_06936_));
 sg13g2_nand2_1 _37526_ (.Y(_06938_),
    .A(_06292_),
    .B(_06302_));
 sg13g2_o21ai_1 _37527_ (.B1(_06273_),
    .Y(_06939_),
    .A1(net5850),
    .A2(_06283_));
 sg13g2_a21oi_1 _37528_ (.A1(_06285_),
    .A2(_06938_),
    .Y(_06940_),
    .B1(_06939_));
 sg13g2_nor2_1 _37529_ (.A(_06336_),
    .B(_06344_),
    .Y(_06941_));
 sg13g2_or2_1 _37530_ (.X(_06942_),
    .B(_06344_),
    .A(_06336_));
 sg13g2_a221oi_1 _37531_ (.B2(_06942_),
    .C1(_06325_),
    .B1(_06327_),
    .A1(net5800),
    .Y(_06943_),
    .A2(_06317_));
 sg13g2_nand2b_1 _37532_ (.Y(_06944_),
    .B(_06307_),
    .A_N(_06943_));
 sg13g2_nand3_1 _37533_ (.B(_06940_),
    .C(_06944_),
    .A(_06937_),
    .Y(_06945_));
 sg13g2_and3_1 _37534_ (.X(_06946_),
    .A(_06487_),
    .B(_06505_),
    .C(_06524_));
 sg13g2_inv_1 _37535_ (.Y(_06947_),
    .A(_06946_));
 sg13g2_nor2_1 _37536_ (.A(_06442_),
    .B(_06947_),
    .Y(_06948_));
 sg13g2_nor3_1 _37537_ (.A(_06348_),
    .B(_06442_),
    .C(_06947_),
    .Y(_06949_));
 sg13g2_a221oi_1 _37538_ (.B2(_06912_),
    .C1(_06928_),
    .B1(_06949_),
    .A1(_06945_),
    .Y(_06950_),
    .A2(_06948_));
 sg13g2_a21oi_2 _37539_ (.B1(_04404_),
    .Y(_06951_),
    .A2(net1071),
    .A1(_04396_));
 sg13g2_a21oi_1 _37540_ (.A1(_04019_),
    .A2(_06951_),
    .Y(_06952_),
    .B1(_04038_));
 sg13g2_a21o_2 _37541_ (.A2(_06951_),
    .A1(_04019_),
    .B1(_04038_),
    .X(_06953_));
 sg13g2_a21oi_1 _37542_ (.A1(_04396_),
    .A2(net1071),
    .Y(_06954_),
    .B1(_04406_));
 sg13g2_nor2_1 _37543_ (.A(_04073_),
    .B(_06954_),
    .Y(_06955_));
 sg13g2_nor2b_1 _37544_ (.A(_06955_),
    .B_N(_03990_),
    .Y(_06956_));
 sg13g2_o21ai_1 _37545_ (.B1(_03990_),
    .Y(_06957_),
    .A1(_04073_),
    .A2(_06954_));
 sg13g2_o21ai_1 _37546_ (.B1(_04096_),
    .Y(_06958_),
    .A1(_04002_),
    .A2(_06957_));
 sg13g2_nand2_1 _37547_ (.Y(_06959_),
    .A(_03979_),
    .B(_06958_));
 sg13g2_nand3_1 _37548_ (.B(_03979_),
    .C(_06958_),
    .A(_03974_),
    .Y(_06960_));
 sg13g2_a21oi_2 _37549_ (.B1(_03963_),
    .Y(_06961_),
    .A2(_06960_),
    .A1(_04080_));
 sg13g2_a21oi_1 _37550_ (.A1(_03962_),
    .A2(_06961_),
    .Y(_06962_),
    .B1(_04082_));
 sg13g2_o21ai_1 _37551_ (.B1(_03956_),
    .Y(_06963_),
    .A1(_03957_),
    .A2(_06962_));
 sg13g2_a21oi_1 _37552_ (.A1(_03959_),
    .A2(_06963_),
    .Y(_06964_),
    .B1(net7232));
 sg13g2_o21ai_1 _37553_ (.B1(_06964_),
    .Y(_06965_),
    .A1(_03959_),
    .A2(_06963_));
 sg13g2_a21oi_1 _37554_ (.A1(net7232),
    .A2(\u_inv.d_next[95] ),
    .Y(_06966_),
    .B1(net6353));
 sg13g2_a21oi_1 _37555_ (.A1(_04965_),
    .A2(_05029_),
    .Y(_06967_),
    .B1(_05058_));
 sg13g2_a21o_2 _37556_ (.A2(_05029_),
    .A1(_04965_),
    .B1(_05058_),
    .X(_06968_));
 sg13g2_a21oi_2 _37557_ (.B1(_05087_),
    .Y(_06969_),
    .A2(_06968_),
    .A1(_05003_));
 sg13g2_o21ai_1 _37558_ (.B1(_05064_),
    .Y(_06970_),
    .A1(_05009_),
    .A2(_06969_));
 sg13g2_a21oi_1 _37559_ (.A1(_05005_),
    .A2(_06970_),
    .Y(_06971_),
    .B1(_05067_));
 sg13g2_o21ai_1 _37560_ (.B1(_05068_),
    .Y(_06972_),
    .A1(_03958_),
    .A2(_06971_));
 sg13g2_nand2b_1 _37561_ (.Y(_06973_),
    .B(_03960_),
    .A_N(_06972_));
 sg13g2_a21oi_1 _37562_ (.A1(_03959_),
    .A2(_06972_),
    .Y(_06974_),
    .B1(net6257));
 sg13g2_a22oi_1 _37563_ (.Y(_06975_),
    .B1(_06973_),
    .B2(_06974_),
    .A2(_06966_),
    .A1(_06965_));
 sg13g2_xnor2_1 _37564_ (.Y(_06976_),
    .A(net5824),
    .B(_06975_));
 sg13g2_xnor2_1 _37565_ (.Y(_06977_),
    .A(_03958_),
    .B(_06971_));
 sg13g2_o21ai_1 _37566_ (.B1(net7392),
    .Y(_06978_),
    .A1(_03957_),
    .A2(_06962_));
 sg13g2_a21o_1 _37567_ (.A2(_06962_),
    .A1(_03957_),
    .B1(_06978_),
    .X(_06979_));
 sg13g2_a21oi_1 _37568_ (.A1(net7232),
    .A2(\u_inv.d_next[94] ),
    .Y(_06980_),
    .B1(net6353));
 sg13g2_a22oi_1 _37569_ (.Y(_06981_),
    .B1(_06979_),
    .B2(_06980_),
    .A2(_06977_),
    .A1(net6353));
 sg13g2_nand2_1 _37570_ (.Y(_06982_),
    .A(net5824),
    .B(_06981_));
 sg13g2_xnor2_1 _37571_ (.Y(_06983_),
    .A(net5824),
    .B(_06981_));
 sg13g2_nor2_1 _37572_ (.A(_06976_),
    .B(_06983_),
    .Y(_06984_));
 sg13g2_a21o_1 _37573_ (.A2(_06970_),
    .A1(_03963_),
    .B1(_05065_),
    .X(_06985_));
 sg13g2_o21ai_1 _37574_ (.B1(net6353),
    .Y(_06986_),
    .A1(_03962_),
    .A2(_06985_));
 sg13g2_a21oi_1 _37575_ (.A1(_03962_),
    .A2(_06985_),
    .Y(_06987_),
    .B1(_06986_));
 sg13g2_a21oi_1 _37576_ (.A1(\u_inv.d_next[92] ),
    .A2(\u_inv.d_reg[92] ),
    .Y(_06988_),
    .B1(_03962_));
 sg13g2_nand2b_1 _37577_ (.Y(_06989_),
    .B(_06988_),
    .A_N(_06961_));
 sg13g2_nand2b_1 _37578_ (.Y(_06990_),
    .B(net7392),
    .A_N(_04081_));
 sg13g2_a21oi_1 _37579_ (.A1(_03962_),
    .A2(_06961_),
    .Y(_06991_),
    .B1(_06990_));
 sg13g2_a22oi_1 _37580_ (.Y(_06992_),
    .B1(_06989_),
    .B2(_06991_),
    .A2(\u_inv.d_next[93] ),
    .A1(net7232));
 sg13g2_a21oi_2 _37581_ (.B1(_06987_),
    .Y(_06993_),
    .A2(_06992_),
    .A1(net6257));
 sg13g2_nand2_1 _37582_ (.Y(_06994_),
    .A(net5824),
    .B(_06993_));
 sg13g2_xnor2_1 _37583_ (.Y(_06995_),
    .A(net5824),
    .B(_06993_));
 sg13g2_xnor2_1 _37584_ (.Y(_06996_),
    .A(_03963_),
    .B(_06970_));
 sg13g2_nand3_1 _37585_ (.B(_04080_),
    .C(_06960_),
    .A(_03963_),
    .Y(_06997_));
 sg13g2_nor2_1 _37586_ (.A(net7231),
    .B(_06961_),
    .Y(_06998_));
 sg13g2_a221oi_1 _37587_ (.B2(_06998_),
    .C1(net6352),
    .B1(_06997_),
    .A1(net7231),
    .Y(_06999_),
    .A2(\u_inv.d_next[92] ));
 sg13g2_a21oi_2 _37588_ (.B1(_06999_),
    .Y(_07000_),
    .A2(_06996_),
    .A1(net6352));
 sg13g2_nand2_1 _37589_ (.Y(_07001_),
    .A(net5824),
    .B(_07000_));
 sg13g2_xnor2_1 _37590_ (.Y(_07002_),
    .A(net5870),
    .B(_07000_));
 sg13g2_nor2b_1 _37591_ (.A(_06995_),
    .B_N(_07002_),
    .Y(_07003_));
 sg13g2_o21ai_1 _37592_ (.B1(_05061_),
    .Y(_07004_),
    .A1(_05008_),
    .A2(_06969_));
 sg13g2_xnor2_1 _37593_ (.Y(_07005_),
    .A(_03973_),
    .B(_07004_));
 sg13g2_nand3_1 _37594_ (.B(_04078_),
    .C(_06959_),
    .A(_03973_),
    .Y(_07006_));
 sg13g2_a21oi_1 _37595_ (.A1(_04078_),
    .A2(_06959_),
    .Y(_07007_),
    .B1(_03973_));
 sg13g2_nand3b_1 _37596_ (.B(net7393),
    .C(_07006_),
    .Y(_07008_),
    .A_N(_07007_));
 sg13g2_a21oi_1 _37597_ (.A1(net7231),
    .A2(\u_inv.d_next[90] ),
    .Y(_07009_),
    .B1(net6352));
 sg13g2_a22oi_1 _37598_ (.Y(_07010_),
    .B1(_07008_),
    .B2(_07009_),
    .A2(_07005_),
    .A1(net6352));
 sg13g2_nand2_1 _37599_ (.Y(_07011_),
    .A(net5823),
    .B(_07010_));
 sg13g2_xnor2_1 _37600_ (.Y(_07012_),
    .A(net5870),
    .B(_07010_));
 sg13g2_inv_1 _37601_ (.Y(_07013_),
    .A(_07012_));
 sg13g2_o21ai_1 _37602_ (.B1(_03969_),
    .Y(_07014_),
    .A1(_03971_),
    .A2(_07007_));
 sg13g2_nor3_1 _37603_ (.A(_03969_),
    .B(_03971_),
    .C(_07007_),
    .Y(_07015_));
 sg13g2_nand2_1 _37604_ (.Y(_07016_),
    .A(net7393),
    .B(_07014_));
 sg13g2_a21oi_1 _37605_ (.A1(net7231),
    .A2(\u_inv.d_next[91] ),
    .Y(_07017_),
    .B1(net6352));
 sg13g2_o21ai_1 _37606_ (.B1(_07017_),
    .Y(_07018_),
    .A1(_07015_),
    .A2(_07016_));
 sg13g2_a21oi_1 _37607_ (.A1(_03973_),
    .A2(_07004_),
    .Y(_07019_),
    .B1(_05062_));
 sg13g2_and2_1 _37608_ (.A(_03968_),
    .B(_07019_),
    .X(_07020_));
 sg13g2_o21ai_1 _37609_ (.B1(net6352),
    .Y(_07021_),
    .A1(_03968_),
    .A2(_07019_));
 sg13g2_o21ai_1 _37610_ (.B1(_07018_),
    .Y(_07022_),
    .A1(_07020_),
    .A2(_07021_));
 sg13g2_nand2b_1 _37611_ (.Y(_07023_),
    .B(net5823),
    .A_N(_07022_));
 sg13g2_xnor2_1 _37612_ (.Y(_07024_),
    .A(net5823),
    .B(_07022_));
 sg13g2_o21ai_1 _37613_ (.B1(_05059_),
    .Y(_07025_),
    .A1(_03978_),
    .A2(_06969_));
 sg13g2_or2_1 _37614_ (.X(_07026_),
    .B(_07025_),
    .A(_03976_));
 sg13g2_a21oi_1 _37615_ (.A1(_03976_),
    .A2(_07025_),
    .Y(_07027_),
    .B1(net6257));
 sg13g2_a21oi_1 _37616_ (.A1(_03978_),
    .A2(_06958_),
    .Y(_07028_),
    .B1(_03977_));
 sg13g2_nand2_1 _37617_ (.Y(_07029_),
    .A(_03975_),
    .B(_07028_));
 sg13g2_nand4_1 _37618_ (.B(_04076_),
    .C(_06959_),
    .A(net7393),
    .Y(_07030_),
    .D(_07029_));
 sg13g2_a21oi_1 _37619_ (.A1(net7231),
    .A2(\u_inv.d_next[89] ),
    .Y(_07031_),
    .B1(net6351));
 sg13g2_a22oi_1 _37620_ (.Y(_07032_),
    .B1(_07030_),
    .B2(_07031_),
    .A2(_07027_),
    .A1(_07026_));
 sg13g2_nand2_1 _37621_ (.Y(_07033_),
    .A(net5823),
    .B(_07032_));
 sg13g2_nor2_1 _37622_ (.A(net5823),
    .B(_07032_),
    .Y(_07034_));
 sg13g2_xnor2_1 _37623_ (.Y(_07035_),
    .A(net5823),
    .B(_07032_));
 sg13g2_inv_1 _37624_ (.Y(_07036_),
    .A(_07035_));
 sg13g2_xnor2_1 _37625_ (.Y(_07037_),
    .A(_03978_),
    .B(_06969_));
 sg13g2_xnor2_1 _37626_ (.Y(_07038_),
    .A(_03978_),
    .B(_06958_));
 sg13g2_o21ai_1 _37627_ (.B1(net6257),
    .Y(_07039_),
    .A1(net7393),
    .A2(\u_inv.d_next[88] ));
 sg13g2_a21o_1 _37628_ (.A2(_07038_),
    .A1(net7393),
    .B1(_07039_),
    .X(_07040_));
 sg13g2_o21ai_1 _37629_ (.B1(_07040_),
    .Y(_07041_),
    .A1(net6257),
    .A2(_07037_));
 sg13g2_nand2_1 _37630_ (.Y(_07042_),
    .A(net5823),
    .B(_07041_));
 sg13g2_xnor2_1 _37631_ (.Y(_07043_),
    .A(net5870),
    .B(_07041_));
 sg13g2_nand4_1 _37632_ (.B(_07024_),
    .C(_07036_),
    .A(_07012_),
    .Y(_07044_),
    .D(_07043_));
 sg13g2_inv_1 _37633_ (.Y(_07045_),
    .A(_07044_));
 sg13g2_and3_2 _37634_ (.X(_07046_),
    .A(_06984_),
    .B(_07003_),
    .C(_07045_));
 sg13g2_nand3_1 _37635_ (.B(_03988_),
    .C(_06968_),
    .A(_03982_),
    .Y(_07047_));
 sg13g2_nand2_1 _37636_ (.Y(_07048_),
    .A(_05074_),
    .B(_07047_));
 sg13g2_a21oi_1 _37637_ (.A1(_05074_),
    .A2(_07047_),
    .Y(_07049_),
    .B1(_05001_));
 sg13g2_nor2_1 _37638_ (.A(_05078_),
    .B(_07049_),
    .Y(_07050_));
 sg13g2_o21ai_1 _37639_ (.B1(_04999_),
    .Y(_07051_),
    .A1(_05078_),
    .A2(_07049_));
 sg13g2_nand2_1 _37640_ (.Y(_07052_),
    .A(_05085_),
    .B(_07051_));
 sg13g2_a21oi_1 _37641_ (.A1(_05085_),
    .A2(_07051_),
    .Y(_07053_),
    .B1(_03996_));
 sg13g2_xnor2_1 _37642_ (.Y(_07054_),
    .A(_03997_),
    .B(_07052_));
 sg13g2_nor2_1 _37643_ (.A(_04091_),
    .B(_06956_),
    .Y(_07055_));
 sg13g2_o21ai_1 _37644_ (.B1(_03994_),
    .Y(_07056_),
    .A1(_04091_),
    .A2(_06956_));
 sg13g2_nand2_1 _37645_ (.Y(_07057_),
    .A(_04093_),
    .B(_07056_));
 sg13g2_nand2_1 _37646_ (.Y(_07058_),
    .A(_03996_),
    .B(_07057_));
 sg13g2_o21ai_1 _37647_ (.B1(net7393),
    .Y(_07059_),
    .A1(_03996_),
    .A2(_07057_));
 sg13g2_nand2b_1 _37648_ (.Y(_07060_),
    .B(_07058_),
    .A_N(_07059_));
 sg13g2_a21oi_1 _37649_ (.A1(net7231),
    .A2(\u_inv.d_next[86] ),
    .Y(_07061_),
    .B1(net6350));
 sg13g2_a22oi_1 _37650_ (.Y(_07062_),
    .B1(_07060_),
    .B2(_07061_),
    .A2(_07054_),
    .A1(net6350));
 sg13g2_nand2_1 _37651_ (.Y(_07063_),
    .A(net5821),
    .B(_07062_));
 sg13g2_xnor2_1 _37652_ (.Y(_07064_),
    .A(net5867),
    .B(_07062_));
 sg13g2_xnor2_1 _37653_ (.Y(_07065_),
    .A(net5821),
    .B(_07062_));
 sg13g2_nand2_1 _37654_ (.Y(_07066_),
    .A(_03995_),
    .B(_07058_));
 sg13g2_o21ai_1 _37655_ (.B1(net7393),
    .Y(_07067_),
    .A1(_04000_),
    .A2(_07066_));
 sg13g2_a21o_1 _37656_ (.A2(_07066_),
    .A1(_04000_),
    .B1(_07067_),
    .X(_07068_));
 sg13g2_nand2_1 _37657_ (.Y(_07069_),
    .A(net7231),
    .B(\u_inv.d_next[87] ));
 sg13g2_nand3_1 _37658_ (.B(_07068_),
    .C(_07069_),
    .A(net6257),
    .Y(_07070_));
 sg13g2_o21ai_1 _37659_ (.B1(_04000_),
    .Y(_07071_),
    .A1(_05080_),
    .A2(_07053_));
 sg13g2_or3_1 _37660_ (.A(_04000_),
    .B(_05080_),
    .C(_07053_),
    .X(_07072_));
 sg13g2_nand3_1 _37661_ (.B(_07071_),
    .C(_07072_),
    .A(net6350),
    .Y(_07073_));
 sg13g2_nand2_1 _37662_ (.Y(_07074_),
    .A(_07070_),
    .B(_07073_));
 sg13g2_and3_1 _37663_ (.X(_07075_),
    .A(net5821),
    .B(_07070_),
    .C(_07073_));
 sg13g2_a21oi_1 _37664_ (.A1(_07070_),
    .A2(_07073_),
    .Y(_07076_),
    .B1(net5821));
 sg13g2_or2_1 _37665_ (.X(_07077_),
    .B(_07076_),
    .A(_07075_));
 sg13g2_nor3_1 _37666_ (.A(_07065_),
    .B(_07075_),
    .C(_07076_),
    .Y(_07078_));
 sg13g2_o21ai_1 _37667_ (.B1(_03993_),
    .Y(_07079_),
    .A1(_05078_),
    .A2(_07049_));
 sg13g2_a21o_1 _37668_ (.A2(_07079_),
    .A1(_05083_),
    .B1(_03991_),
    .X(_07080_));
 sg13g2_nand3_1 _37669_ (.B(_05083_),
    .C(_07079_),
    .A(_03991_),
    .Y(_07081_));
 sg13g2_nand3_1 _37670_ (.B(_07080_),
    .C(_07081_),
    .A(net6350),
    .Y(_07082_));
 sg13g2_or2_1 _37671_ (.X(_07083_),
    .B(_07055_),
    .A(_03993_));
 sg13g2_a21oi_1 _37672_ (.A1(_03992_),
    .A2(_07083_),
    .Y(_07084_),
    .B1(_03991_));
 sg13g2_nand3_1 _37673_ (.B(_03992_),
    .C(_07083_),
    .A(_03991_),
    .Y(_07085_));
 sg13g2_nand2_1 _37674_ (.Y(_07086_),
    .A(net7393),
    .B(_07085_));
 sg13g2_a21oi_1 _37675_ (.A1(net7234),
    .A2(\u_inv.d_next[85] ),
    .Y(_07087_),
    .B1(net6350));
 sg13g2_o21ai_1 _37676_ (.B1(_07087_),
    .Y(_07088_),
    .A1(_07084_),
    .A2(_07086_));
 sg13g2_nand2_1 _37677_ (.Y(_07089_),
    .A(_07082_),
    .B(_07088_));
 sg13g2_nand2_1 _37678_ (.Y(_07090_),
    .A(net5822),
    .B(_07089_));
 sg13g2_nand3_1 _37679_ (.B(_07082_),
    .C(_07088_),
    .A(net5867),
    .Y(_07091_));
 sg13g2_xnor2_1 _37680_ (.Y(_07092_),
    .A(net5867),
    .B(_07089_));
 sg13g2_xor2_1 _37681_ (.B(_07050_),
    .A(_03993_),
    .X(_07093_));
 sg13g2_a21oi_1 _37682_ (.A1(_03993_),
    .A2(_07055_),
    .Y(_07094_),
    .B1(net7231));
 sg13g2_a221oi_1 _37683_ (.B2(_07094_),
    .C1(net6350),
    .B1(_07083_),
    .A1(net7234),
    .Y(_07095_),
    .A2(\u_inv.d_next[84] ));
 sg13g2_a21oi_2 _37684_ (.B1(_07095_),
    .Y(_07096_),
    .A2(_07093_),
    .A1(net6350));
 sg13g2_nand2_1 _37685_ (.Y(_07097_),
    .A(net5821),
    .B(_07096_));
 sg13g2_xnor2_1 _37686_ (.Y(_07098_),
    .A(net5821),
    .B(_07096_));
 sg13g2_nor2_1 _37687_ (.A(_07092_),
    .B(_07098_),
    .Y(_07099_));
 sg13g2_nand2_1 _37688_ (.Y(_07100_),
    .A(_07078_),
    .B(_07099_));
 sg13g2_o21ai_1 _37689_ (.B1(_03989_),
    .Y(_07101_),
    .A1(_04073_),
    .A2(_06954_));
 sg13g2_nand2b_1 _37690_ (.Y(_07102_),
    .B(_03983_),
    .A_N(_07101_));
 sg13g2_a21o_1 _37691_ (.A2(_07102_),
    .A1(_04088_),
    .B1(_03986_),
    .X(_07103_));
 sg13g2_a21oi_1 _37692_ (.A1(_03985_),
    .A2(_07103_),
    .Y(_07104_),
    .B1(_03981_));
 sg13g2_nand3_1 _37693_ (.B(_03985_),
    .C(_07103_),
    .A(_03981_),
    .Y(_07105_));
 sg13g2_nor2_1 _37694_ (.A(net7238),
    .B(_07104_),
    .Y(_07106_));
 sg13g2_a221oi_1 _37695_ (.B2(_07106_),
    .C1(net6350),
    .B1(_07105_),
    .A1(net7238),
    .Y(_07107_),
    .A2(\u_inv.d_next[83] ));
 sg13g2_a21oi_1 _37696_ (.A1(_03986_),
    .A2(_07048_),
    .Y(_07108_),
    .B1(_05076_));
 sg13g2_xor2_1 _37697_ (.B(_07108_),
    .A(_03981_),
    .X(_07109_));
 sg13g2_a21o_2 _37698_ (.A2(_07109_),
    .A1(net6351),
    .B1(_07107_),
    .X(_07110_));
 sg13g2_xnor2_1 _37699_ (.Y(_07111_),
    .A(net5867),
    .B(_07110_));
 sg13g2_nand3_1 _37700_ (.B(_04088_),
    .C(_07102_),
    .A(_03986_),
    .Y(_07112_));
 sg13g2_a21oi_1 _37701_ (.A1(_07103_),
    .A2(_07112_),
    .Y(_07113_),
    .B1(net7234));
 sg13g2_o21ai_1 _37702_ (.B1(net6267),
    .Y(_07114_),
    .A1(net7405),
    .A2(\u_inv.d_next[82] ));
 sg13g2_nor2_1 _37703_ (.A(_07113_),
    .B(_07114_),
    .Y(_07115_));
 sg13g2_xor2_1 _37704_ (.B(_07048_),
    .A(_03986_),
    .X(_07116_));
 sg13g2_a21oi_2 _37705_ (.B1(_07115_),
    .Y(_07117_),
    .A2(_07116_),
    .A1(net6351));
 sg13g2_or2_1 _37706_ (.X(_07118_),
    .B(_07117_),
    .A(net5867));
 sg13g2_xnor2_1 _37707_ (.Y(_07119_),
    .A(net5867),
    .B(_07117_));
 sg13g2_nor2_1 _37708_ (.A(_07111_),
    .B(_07119_),
    .Y(_07120_));
 sg13g2_nand2_1 _37709_ (.Y(_07121_),
    .A(_03988_),
    .B(_06955_));
 sg13g2_nand3_1 _37710_ (.B(_07101_),
    .C(_07121_),
    .A(net7405),
    .Y(_07122_));
 sg13g2_xnor2_1 _37711_ (.Y(_07123_),
    .A(_03989_),
    .B(_06967_));
 sg13g2_a21oi_1 _37712_ (.A1(net7238),
    .A2(\u_inv.d_next[80] ),
    .Y(_07124_),
    .B1(net6362));
 sg13g2_a22oi_1 _37713_ (.Y(_07125_),
    .B1(_07124_),
    .B2(_07122_),
    .A2(_07123_),
    .A1(net6362));
 sg13g2_and2_1 _37714_ (.A(net5822),
    .B(_07125_),
    .X(_07126_));
 sg13g2_xnor2_1 _37715_ (.Y(_07127_),
    .A(net5867),
    .B(_07125_));
 sg13g2_inv_1 _37716_ (.Y(_07128_),
    .A(_07127_));
 sg13g2_nand3_1 _37717_ (.B(_03987_),
    .C(_07101_),
    .A(_03982_),
    .Y(_07129_));
 sg13g2_o21ai_1 _37718_ (.B1(net7405),
    .Y(_07130_),
    .A1(_03982_),
    .A2(_03987_));
 sg13g2_nor2b_1 _37719_ (.A(_07130_),
    .B_N(_07102_),
    .Y(_07131_));
 sg13g2_a22oi_1 _37720_ (.Y(_07132_),
    .B1(_07129_),
    .B2(_07131_),
    .A2(\u_inv.d_next[81] ),
    .A1(net7238));
 sg13g2_o21ai_1 _37721_ (.B1(_05072_),
    .Y(_07133_),
    .A1(_03989_),
    .A2(_06967_));
 sg13g2_o21ai_1 _37722_ (.B1(net6362),
    .Y(_07134_),
    .A1(_03983_),
    .A2(_07133_));
 sg13g2_a21oi_1 _37723_ (.A1(_03983_),
    .A2(_07133_),
    .Y(_07135_),
    .B1(_07134_));
 sg13g2_a21oi_2 _37724_ (.B1(_07135_),
    .Y(_07136_),
    .A2(_07132_),
    .A1(net6267));
 sg13g2_xnor2_1 _37725_ (.Y(_07137_),
    .A(net5871),
    .B(_07136_));
 sg13g2_and3_1 _37726_ (.X(_07138_),
    .A(_07120_),
    .B(_07127_),
    .C(_07137_));
 sg13g2_and3_2 _37727_ (.X(_07139_),
    .A(_07078_),
    .B(_07099_),
    .C(_07138_));
 sg13g2_inv_1 _37728_ (.Y(_07140_),
    .A(_07139_));
 sg13g2_and2_1 _37729_ (.A(_07046_),
    .B(_07139_),
    .X(_07141_));
 sg13g2_nand2b_1 _37730_ (.Y(_07142_),
    .B(_04965_),
    .A_N(_04401_));
 sg13g2_nor3_2 _37731_ (.A(_04964_),
    .B(_05016_),
    .C(_05026_),
    .Y(_07143_));
 sg13g2_nor2_1 _37732_ (.A(_05043_),
    .B(_07143_),
    .Y(_07144_));
 sg13g2_o21ai_1 _37733_ (.B1(_05023_),
    .Y(_07145_),
    .A1(_05043_),
    .A2(_07143_));
 sg13g2_a21oi_1 _37734_ (.A1(_05051_),
    .A2(_07145_),
    .Y(_07146_),
    .B1(_05024_));
 sg13g2_nor2_1 _37735_ (.A(_05055_),
    .B(_07146_),
    .Y(_07147_));
 sg13g2_o21ai_1 _37736_ (.B1(_05019_),
    .Y(_07148_),
    .A1(_05055_),
    .A2(_07146_));
 sg13g2_nand3_1 _37737_ (.B(_05046_),
    .C(_07148_),
    .A(_04043_),
    .Y(_07149_));
 sg13g2_a21o_1 _37738_ (.A2(_07148_),
    .A1(_05046_),
    .B1(_04043_),
    .X(_07150_));
 sg13g2_a21oi_1 _37739_ (.A1(_07149_),
    .A2(_07150_),
    .Y(_07151_),
    .B1(net6268));
 sg13g2_nand2_1 _37740_ (.Y(_07152_),
    .A(_04058_),
    .B(_06953_));
 sg13g2_or2_1 _37741_ (.X(_07153_),
    .B(_07152_),
    .A(_04056_));
 sg13g2_a21oi_1 _37742_ (.A1(_04060_),
    .A2(_06953_),
    .Y(_07154_),
    .B1(_04067_));
 sg13g2_nor3_1 _37743_ (.A(_04039_),
    .B(_04041_),
    .C(_07154_),
    .Y(_07155_));
 sg13g2_o21ai_1 _37744_ (.B1(_04043_),
    .Y(_07156_),
    .A1(_04069_),
    .A2(_07155_));
 sg13g2_nor3_1 _37745_ (.A(_04043_),
    .B(_04069_),
    .C(_07155_),
    .Y(_07157_));
 sg13g2_nor2_1 _37746_ (.A(net7240),
    .B(_07157_),
    .Y(_07158_));
 sg13g2_nand2_1 _37747_ (.Y(_07159_),
    .A(net7240),
    .B(\u_inv.d_next[78] ));
 sg13g2_a21oi_1 _37748_ (.A1(_07156_),
    .A2(_07158_),
    .Y(_07160_),
    .B1(net6364));
 sg13g2_a21oi_2 _37749_ (.B1(_07151_),
    .Y(_07161_),
    .A2(_07160_),
    .A1(_07159_));
 sg13g2_nand2_1 _37750_ (.Y(_07162_),
    .A(net5827),
    .B(_07161_));
 sg13g2_xnor2_1 _37751_ (.Y(_07163_),
    .A(net5827),
    .B(_07161_));
 sg13g2_a21oi_1 _37752_ (.A1(_05047_),
    .A2(_07150_),
    .Y(_07164_),
    .B1(_04047_));
 sg13g2_nand3_1 _37753_ (.B(_05047_),
    .C(_07150_),
    .A(_04047_),
    .Y(_07165_));
 sg13g2_nand3b_1 _37754_ (.B(_07165_),
    .C(net6364),
    .Y(_07166_),
    .A_N(_07164_));
 sg13g2_a21o_1 _37755_ (.A2(_07156_),
    .A1(_04042_),
    .B1(_04047_),
    .X(_07167_));
 sg13g2_nand3_1 _37756_ (.B(_04047_),
    .C(_07156_),
    .A(_04042_),
    .Y(_07168_));
 sg13g2_nand3_1 _37757_ (.B(_07167_),
    .C(_07168_),
    .A(net7407),
    .Y(_07169_));
 sg13g2_nand2_1 _37758_ (.Y(_07170_),
    .A(net7243),
    .B(\u_inv.d_next[79] ));
 sg13g2_nand3_1 _37759_ (.B(_07169_),
    .C(_07170_),
    .A(net6268),
    .Y(_07171_));
 sg13g2_and3_1 _37760_ (.X(_07172_),
    .A(net5827),
    .B(_07166_),
    .C(_07171_));
 sg13g2_a21oi_1 _37761_ (.A1(_07166_),
    .A2(_07171_),
    .Y(_07173_),
    .B1(net5827));
 sg13g2_or2_1 _37762_ (.X(_07174_),
    .B(_07173_),
    .A(_07172_));
 sg13g2_nor3_1 _37763_ (.A(_07163_),
    .B(_07172_),
    .C(_07173_),
    .Y(_07175_));
 sg13g2_or2_1 _37764_ (.X(_07176_),
    .B(_07154_),
    .A(_04041_));
 sg13g2_xnor2_1 _37765_ (.Y(_07177_),
    .A(_04041_),
    .B(_07154_));
 sg13g2_o21ai_1 _37766_ (.B1(net6265),
    .Y(_07178_),
    .A1(net7403),
    .A2(\u_inv.d_next[76] ));
 sg13g2_a21oi_1 _37767_ (.A1(net7407),
    .A2(_07177_),
    .Y(_07179_),
    .B1(_07178_));
 sg13g2_o21ai_1 _37768_ (.B1(_04041_),
    .Y(_07180_),
    .A1(_05055_),
    .A2(_07146_));
 sg13g2_xnor2_1 _37769_ (.Y(_07181_),
    .A(_04041_),
    .B(_07147_));
 sg13g2_a21oi_2 _37770_ (.B1(_07179_),
    .Y(_07182_),
    .A2(_07181_),
    .A1(net6364));
 sg13g2_nor2_1 _37771_ (.A(net5872),
    .B(_07182_),
    .Y(_07183_));
 sg13g2_xnor2_1 _37772_ (.Y(_07184_),
    .A(net5827),
    .B(_07182_));
 sg13g2_a21o_1 _37773_ (.A2(_07180_),
    .A1(_05044_),
    .B1(_04039_),
    .X(_07185_));
 sg13g2_nand3_1 _37774_ (.B(_05044_),
    .C(_07180_),
    .A(_04039_),
    .Y(_07186_));
 sg13g2_nand3_1 _37775_ (.B(_07185_),
    .C(_07186_),
    .A(net6364),
    .Y(_07187_));
 sg13g2_nand3_1 _37776_ (.B(_04040_),
    .C(_07176_),
    .A(_04039_),
    .Y(_07188_));
 sg13g2_a21o_1 _37777_ (.A2(_07176_),
    .A1(_04040_),
    .B1(_04039_),
    .X(_07189_));
 sg13g2_nand3_1 _37778_ (.B(_07188_),
    .C(_07189_),
    .A(net7403),
    .Y(_07190_));
 sg13g2_nand2_1 _37779_ (.Y(_07191_),
    .A(net7236),
    .B(\u_inv.d_next[77] ));
 sg13g2_nand3_1 _37780_ (.B(_07190_),
    .C(_07191_),
    .A(net6268),
    .Y(_07192_));
 sg13g2_nand2_1 _37781_ (.Y(_07193_),
    .A(_07187_),
    .B(_07192_));
 sg13g2_nand3_1 _37782_ (.B(_07187_),
    .C(_07192_),
    .A(net5827),
    .Y(_07194_));
 sg13g2_a21oi_1 _37783_ (.A1(_07187_),
    .A2(_07192_),
    .Y(_07195_),
    .B1(net5827));
 sg13g2_xnor2_1 _37784_ (.Y(_07196_),
    .A(net5827),
    .B(_07193_));
 sg13g2_and2_1 _37785_ (.A(_07184_),
    .B(_07196_),
    .X(_07197_));
 sg13g2_nand3b_1 _37786_ (.B(_07184_),
    .C(_07194_),
    .Y(_07198_),
    .A_N(_07195_));
 sg13g2_nor4_1 _37787_ (.A(_07163_),
    .B(_07172_),
    .C(_07173_),
    .D(_07198_),
    .Y(_07199_));
 sg13g2_nor2_1 _37788_ (.A(_04058_),
    .B(_07144_),
    .Y(_07200_));
 sg13g2_nor2_1 _37789_ (.A(_05049_),
    .B(_07200_),
    .Y(_07201_));
 sg13g2_o21ai_1 _37790_ (.B1(net6364),
    .Y(_07202_),
    .A1(_04056_),
    .A2(_07201_));
 sg13g2_a21oi_1 _37791_ (.A1(_04056_),
    .A2(_07201_),
    .Y(_07203_),
    .B1(_07202_));
 sg13g2_a21o_1 _37792_ (.A2(_07152_),
    .A1(_04057_),
    .B1(_04056_),
    .X(_07204_));
 sg13g2_nand3_1 _37793_ (.B(_04057_),
    .C(_07152_),
    .A(_04056_),
    .Y(_07205_));
 sg13g2_nand3_1 _37794_ (.B(_07204_),
    .C(_07205_),
    .A(net7408),
    .Y(_07206_));
 sg13g2_a21oi_1 _37795_ (.A1(net7240),
    .A2(\u_inv.d_next[73] ),
    .Y(_07207_),
    .B1(net6365));
 sg13g2_a21oi_2 _37796_ (.B1(_07203_),
    .Y(_07208_),
    .A2(_07207_),
    .A1(_07206_));
 sg13g2_xnor2_1 _37797_ (.Y(_07209_),
    .A(net5828),
    .B(_07208_));
 sg13g2_xnor2_1 _37798_ (.Y(_07210_),
    .A(_04059_),
    .B(_06952_));
 sg13g2_o21ai_1 _37799_ (.B1(net6268),
    .Y(_07211_),
    .A1(net7407),
    .A2(\u_inv.d_next[72] ));
 sg13g2_a21oi_1 _37800_ (.A1(net7408),
    .A2(_07210_),
    .Y(_07212_),
    .B1(_07211_));
 sg13g2_xnor2_1 _37801_ (.Y(_07213_),
    .A(_04059_),
    .B(_07144_));
 sg13g2_a21oi_1 _37802_ (.A1(net6365),
    .A2(_07213_),
    .Y(_07214_),
    .B1(_07212_));
 sg13g2_nor2_1 _37803_ (.A(net5873),
    .B(_07214_),
    .Y(_07215_));
 sg13g2_inv_1 _37804_ (.Y(_07216_),
    .A(_07215_));
 sg13g2_xnor2_1 _37805_ (.Y(_07217_),
    .A(net5873),
    .B(_07214_));
 sg13g2_nor2_1 _37806_ (.A(_07209_),
    .B(_07217_),
    .Y(_07218_));
 sg13g2_a21oi_1 _37807_ (.A1(_05051_),
    .A2(_07145_),
    .Y(_07219_),
    .B1(_04052_));
 sg13g2_o21ai_1 _37808_ (.B1(_04050_),
    .Y(_07220_),
    .A1(_05053_),
    .A2(_07219_));
 sg13g2_nor3_1 _37809_ (.A(_04050_),
    .B(_05053_),
    .C(_07219_),
    .Y(_07221_));
 sg13g2_nand3b_1 _37810_ (.B(net6364),
    .C(_07220_),
    .Y(_07222_),
    .A_N(_07221_));
 sg13g2_a21oi_1 _37811_ (.A1(_04065_),
    .A2(_07153_),
    .Y(_07223_),
    .B1(_04053_));
 sg13g2_nor2_1 _37812_ (.A(_04051_),
    .B(_07223_),
    .Y(_07224_));
 sg13g2_o21ai_1 _37813_ (.B1(net7408),
    .Y(_07225_),
    .A1(_04049_),
    .A2(_07224_));
 sg13g2_a21oi_1 _37814_ (.A1(_04049_),
    .A2(_07224_),
    .Y(_07226_),
    .B1(_07225_));
 sg13g2_o21ai_1 _37815_ (.B1(net6268),
    .Y(_07227_),
    .A1(net7408),
    .A2(_18156_));
 sg13g2_o21ai_1 _37816_ (.B1(_07222_),
    .Y(_07228_),
    .A1(_07226_),
    .A2(_07227_));
 sg13g2_xnor2_1 _37817_ (.Y(_07229_),
    .A(net5873),
    .B(_07228_));
 sg13g2_nand3_1 _37818_ (.B(_04065_),
    .C(_07153_),
    .A(_04053_),
    .Y(_07230_));
 sg13g2_nor2_1 _37819_ (.A(net7240),
    .B(_07223_),
    .Y(_07231_));
 sg13g2_nand3_1 _37820_ (.B(_05051_),
    .C(_07145_),
    .A(_04052_),
    .Y(_07232_));
 sg13g2_nand2b_1 _37821_ (.Y(_07233_),
    .B(_07232_),
    .A_N(_07219_));
 sg13g2_a221oi_1 _37822_ (.B2(_07231_),
    .C1(net6364),
    .B1(_07230_),
    .A1(net7240),
    .Y(_07234_),
    .A2(\u_inv.d_next[74] ));
 sg13g2_a21o_2 _37823_ (.A2(_07233_),
    .A1(net6364),
    .B1(_07234_),
    .X(_07235_));
 sg13g2_nor2_1 _37824_ (.A(net5873),
    .B(_07235_),
    .Y(_07236_));
 sg13g2_xnor2_1 _37825_ (.Y(_07237_),
    .A(net5873),
    .B(_07235_));
 sg13g2_nor2_1 _37826_ (.A(_07229_),
    .B(_07237_),
    .Y(_07238_));
 sg13g2_or2_1 _37827_ (.X(_07239_),
    .B(_07237_),
    .A(_07229_));
 sg13g2_nand3_1 _37828_ (.B(_07218_),
    .C(_07238_),
    .A(_07199_),
    .Y(_07240_));
 sg13g2_o21ai_1 _37829_ (.B1(_05033_),
    .Y(_07241_),
    .A1(_04964_),
    .A2(_05026_));
 sg13g2_a21oi_2 _37830_ (.B1(_05036_),
    .Y(_07242_),
    .A2(_07241_),
    .A1(_05015_));
 sg13g2_nor3_1 _37831_ (.A(_04006_),
    .B(_04009_),
    .C(_07242_),
    .Y(_07243_));
 sg13g2_o21ai_1 _37832_ (.B1(_04014_),
    .Y(_07244_),
    .A1(_05041_),
    .A2(_07243_));
 sg13g2_a21o_1 _37833_ (.A2(_07244_),
    .A1(_05037_),
    .B1(_04017_),
    .X(_07245_));
 sg13g2_nand3_1 _37834_ (.B(_05037_),
    .C(_07244_),
    .A(_04017_),
    .Y(_07246_));
 sg13g2_nand3_1 _37835_ (.B(_07245_),
    .C(_07246_),
    .A(net6365),
    .Y(_07247_));
 sg13g2_nor2_1 _37836_ (.A(_04032_),
    .B(_06951_),
    .Y(_07248_));
 sg13g2_or2_1 _37837_ (.X(_07249_),
    .B(_07248_),
    .A(_04011_));
 sg13g2_a21o_1 _37838_ (.A2(_07249_),
    .A1(_04034_),
    .B1(_04014_),
    .X(_07250_));
 sg13g2_nand3_1 _37839_ (.B(_04017_),
    .C(_07250_),
    .A(_04012_),
    .Y(_07251_));
 sg13g2_a21oi_1 _37840_ (.A1(_04012_),
    .A2(_07250_),
    .Y(_07252_),
    .B1(_04017_));
 sg13g2_nand2_1 _37841_ (.Y(_07253_),
    .A(net7407),
    .B(_07251_));
 sg13g2_a21oi_1 _37842_ (.A1(net7240),
    .A2(\u_inv.d_next[71] ),
    .Y(_07254_),
    .B1(net6365));
 sg13g2_o21ai_1 _37843_ (.B1(_07254_),
    .Y(_07255_),
    .A1(_07252_),
    .A2(_07253_));
 sg13g2_and3_2 _37844_ (.X(_07256_),
    .A(net5829),
    .B(_07247_),
    .C(_07255_));
 sg13g2_a21oi_1 _37845_ (.A1(_07247_),
    .A2(_07255_),
    .Y(_07257_),
    .B1(net5829));
 sg13g2_nor2_1 _37846_ (.A(_07256_),
    .B(_07257_),
    .Y(_07258_));
 sg13g2_or3_1 _37847_ (.A(_04014_),
    .B(_05041_),
    .C(_07243_),
    .X(_07259_));
 sg13g2_and2_1 _37848_ (.A(_07244_),
    .B(_07259_),
    .X(_07260_));
 sg13g2_nand3_1 _37849_ (.B(_04034_),
    .C(_07249_),
    .A(_04014_),
    .Y(_07261_));
 sg13g2_nand3_1 _37850_ (.B(_07250_),
    .C(_07261_),
    .A(net7407),
    .Y(_07262_));
 sg13g2_nand2_1 _37851_ (.Y(_07263_),
    .A(net7240),
    .B(net7297));
 sg13g2_a21oi_1 _37852_ (.A1(_07262_),
    .A2(_07263_),
    .Y(_07264_),
    .B1(net6365));
 sg13g2_a21oi_2 _37853_ (.B1(_07264_),
    .Y(_07265_),
    .A2(_07260_),
    .A1(net6365));
 sg13g2_nor2_1 _37854_ (.A(net5872),
    .B(_07265_),
    .Y(_07266_));
 sg13g2_xnor2_1 _37855_ (.Y(_07267_),
    .A(net5872),
    .B(_07265_));
 sg13g2_inv_1 _37856_ (.Y(_07268_),
    .A(_07267_));
 sg13g2_nor3_1 _37857_ (.A(_07256_),
    .B(_07257_),
    .C(_07267_),
    .Y(_07269_));
 sg13g2_o21ai_1 _37858_ (.B1(_05039_),
    .Y(_07270_),
    .A1(_04006_),
    .A2(_07242_));
 sg13g2_nand2b_1 _37859_ (.Y(_07271_),
    .B(_04010_),
    .A_N(_07270_));
 sg13g2_a21oi_1 _37860_ (.A1(_04009_),
    .A2(_07270_),
    .Y(_07272_),
    .B1(net6268));
 sg13g2_o21ai_1 _37861_ (.B1(_04006_),
    .Y(_07273_),
    .A1(_04032_),
    .A2(_06951_));
 sg13g2_a21o_1 _37862_ (.A2(_07273_),
    .A1(_04005_),
    .B1(_04010_),
    .X(_07274_));
 sg13g2_nand3_1 _37863_ (.B(_04010_),
    .C(_07273_),
    .A(_04005_),
    .Y(_07275_));
 sg13g2_nand3_1 _37864_ (.B(_07274_),
    .C(_07275_),
    .A(net7407),
    .Y(_07276_));
 sg13g2_a21oi_1 _37865_ (.A1(net7240),
    .A2(\u_inv.d_next[69] ),
    .Y(_07277_),
    .B1(net6365));
 sg13g2_a22oi_1 _37866_ (.Y(_07278_),
    .B1(_07276_),
    .B2(_07277_),
    .A2(_07272_),
    .A1(_07271_));
 sg13g2_inv_1 _37867_ (.Y(_07279_),
    .A(_07278_));
 sg13g2_xor2_1 _37868_ (.B(_07248_),
    .A(_04006_),
    .X(_07280_));
 sg13g2_o21ai_1 _37869_ (.B1(net6268),
    .Y(_07281_),
    .A1(net7407),
    .A2(\u_inv.d_next[68] ));
 sg13g2_a21oi_1 _37870_ (.A1(net7407),
    .A2(_07280_),
    .Y(_07282_),
    .B1(_07281_));
 sg13g2_xor2_1 _37871_ (.B(_07242_),
    .A(_04006_),
    .X(_07283_));
 sg13g2_a21oi_2 _37872_ (.B1(_07282_),
    .Y(_07284_),
    .A2(_07283_),
    .A1(net6365));
 sg13g2_a21o_1 _37873_ (.A2(_07284_),
    .A1(_07279_),
    .B1(net5872),
    .X(_07285_));
 sg13g2_nor4_1 _37874_ (.A(_07256_),
    .B(_07257_),
    .C(_07267_),
    .D(_07285_),
    .Y(_07286_));
 sg13g2_or3_1 _37875_ (.A(_07256_),
    .B(_07266_),
    .C(_07286_),
    .X(_07287_));
 sg13g2_xnor2_1 _37876_ (.Y(_07288_),
    .A(net5872),
    .B(_07278_));
 sg13g2_xnor2_1 _37877_ (.Y(_07289_),
    .A(net5829),
    .B(_07284_));
 sg13g2_and3_2 _37878_ (.X(_07290_),
    .A(_07269_),
    .B(_07288_),
    .C(_07289_));
 sg13g2_nand3_1 _37879_ (.B(_07288_),
    .C(_07289_),
    .A(_07269_),
    .Y(_07291_));
 sg13g2_xor2_1 _37880_ (.B(_07241_),
    .A(_04031_),
    .X(_07292_));
 sg13g2_nor2_1 _37881_ (.A(_04400_),
    .B(_04402_),
    .Y(_07293_));
 sg13g2_or3_1 _37882_ (.A(_04026_),
    .B(_04027_),
    .C(_07293_),
    .X(_07294_));
 sg13g2_nand2b_1 _37883_ (.Y(_07295_),
    .B(_07294_),
    .A_N(_04031_));
 sg13g2_xor2_1 _37884_ (.B(_07294_),
    .A(_04031_),
    .X(_07296_));
 sg13g2_a21oi_1 _37885_ (.A1(net7238),
    .A2(\u_inv.d_next[66] ),
    .Y(_07297_),
    .B1(net6362));
 sg13g2_o21ai_1 _37886_ (.B1(_07297_),
    .Y(_07298_),
    .A1(net7238),
    .A2(_07296_));
 sg13g2_o21ai_1 _37887_ (.B1(_07298_),
    .Y(_07299_),
    .A1(net6267),
    .A2(_07292_));
 sg13g2_nor2_1 _37888_ (.A(net5874),
    .B(_07299_),
    .Y(_07300_));
 sg13g2_xnor2_1 _37889_ (.Y(_07301_),
    .A(net5831),
    .B(_07299_));
 sg13g2_a21oi_1 _37890_ (.A1(_04031_),
    .A2(_07241_),
    .Y(_07302_),
    .B1(_05034_));
 sg13g2_o21ai_1 _37891_ (.B1(net6362),
    .Y(_07303_),
    .A1(_04029_),
    .A2(_07302_));
 sg13g2_a21oi_1 _37892_ (.A1(_04029_),
    .A2(_07302_),
    .Y(_07304_),
    .B1(_07303_));
 sg13g2_a21oi_1 _37893_ (.A1(_04021_),
    .A2(_07295_),
    .Y(_07305_),
    .B1(_04029_));
 sg13g2_nand3_1 _37894_ (.B(_04029_),
    .C(_07295_),
    .A(_04021_),
    .Y(_07306_));
 sg13g2_nor2_1 _37895_ (.A(net7238),
    .B(_07305_),
    .Y(_07307_));
 sg13g2_a221oi_1 _37896_ (.B2(_07307_),
    .C1(net6362),
    .B1(_07306_),
    .A1(net7238),
    .Y(_07308_),
    .A2(\u_inv.d_next[67] ));
 sg13g2_or2_1 _37897_ (.X(_07309_),
    .B(_07308_),
    .A(_07304_));
 sg13g2_xnor2_1 _37898_ (.Y(_07310_),
    .A(net5831),
    .B(_07309_));
 sg13g2_nand2_1 _37899_ (.Y(_07311_),
    .A(_07301_),
    .B(_07310_));
 sg13g2_nand2b_1 _37900_ (.Y(_07312_),
    .B(_07142_),
    .A_N(_05032_));
 sg13g2_or2_1 _37901_ (.X(_07313_),
    .B(_07312_),
    .A(_04024_));
 sg13g2_a21oi_1 _37902_ (.A1(_04024_),
    .A2(_07312_),
    .Y(_07314_),
    .B1(net6267));
 sg13g2_a21oi_1 _37903_ (.A1(_04399_),
    .A2(_04401_),
    .Y(_07315_),
    .B1(_04025_));
 sg13g2_nor2b_1 _37904_ (.A(_04024_),
    .B_N(_07315_),
    .Y(_07316_));
 sg13g2_nor4_1 _37905_ (.A(net7239),
    .B(_04026_),
    .C(_07293_),
    .D(_07316_),
    .Y(_07317_));
 sg13g2_a21oi_1 _37906_ (.A1(net7239),
    .A2(\u_inv.d_next[65] ),
    .Y(_07318_),
    .B1(_07317_));
 sg13g2_a22oi_1 _37907_ (.Y(_07319_),
    .B1(_07318_),
    .B2(net6267),
    .A2(_07314_),
    .A1(_07313_));
 sg13g2_xnor2_1 _37908_ (.Y(_07320_),
    .A(_04399_),
    .B(_04401_));
 sg13g2_nor2_1 _37909_ (.A(net7405),
    .B(\u_inv.d_next[64] ),
    .Y(_07321_));
 sg13g2_a21oi_1 _37910_ (.A1(net7405),
    .A2(_07320_),
    .Y(_07322_),
    .B1(_07321_));
 sg13g2_a21oi_1 _37911_ (.A1(_04401_),
    .A2(_04964_),
    .Y(_07323_),
    .B1(net6267));
 sg13g2_a22oi_1 _37912_ (.Y(_07324_),
    .B1(_07323_),
    .B2(_07142_),
    .A2(_07322_),
    .A1(net6267));
 sg13g2_nor2_1 _37913_ (.A(net5874),
    .B(_07324_),
    .Y(_07325_));
 sg13g2_inv_1 _37914_ (.Y(_07326_),
    .A(_07325_));
 sg13g2_a21oi_1 _37915_ (.A1(net5833),
    .A2(_07319_),
    .Y(_07327_),
    .B1(_07325_));
 sg13g2_nor2_1 _37916_ (.A(_07311_),
    .B(_07327_),
    .Y(_07328_));
 sg13g2_a21o_1 _37917_ (.A2(_07309_),
    .A1(_07299_),
    .B1(net5874),
    .X(_07329_));
 sg13g2_nor2b_1 _37918_ (.A(_07328_),
    .B_N(_07329_),
    .Y(_07330_));
 sg13g2_o21ai_1 _37919_ (.B1(_07329_),
    .Y(_07331_),
    .A1(_07311_),
    .A2(_07327_));
 sg13g2_a21oi_1 _37920_ (.A1(_07290_),
    .A2(_07331_),
    .Y(_07332_),
    .B1(_07287_));
 sg13g2_nor2_1 _37921_ (.A(_07240_),
    .B(_07332_),
    .Y(_07333_));
 sg13g2_nand2b_1 _37922_ (.Y(_07334_),
    .B(_07194_),
    .A_N(_07183_));
 sg13g2_a21o_1 _37923_ (.A2(_07161_),
    .A1(net5828),
    .B1(_07172_),
    .X(_07335_));
 sg13g2_a21oi_2 _37924_ (.B1(_07215_),
    .Y(_07336_),
    .A2(_07208_),
    .A1(net5828));
 sg13g2_nor2_1 _37925_ (.A(_07239_),
    .B(_07336_),
    .Y(_07337_));
 sg13g2_a21o_1 _37926_ (.A2(_07235_),
    .A1(_07228_),
    .B1(net5873),
    .X(_07338_));
 sg13g2_nor2b_1 _37927_ (.A(_07337_),
    .B_N(_07338_),
    .Y(_07339_));
 sg13g2_o21ai_1 _37928_ (.B1(_07338_),
    .Y(_07340_),
    .A1(_07239_),
    .A2(_07336_));
 sg13g2_a221oi_1 _37929_ (.B2(_07199_),
    .C1(_07335_),
    .B1(_07340_),
    .A1(_07175_),
    .Y(_07341_),
    .A2(_07334_));
 sg13g2_nor2b_2 _37930_ (.A(_07333_),
    .B_N(_07341_),
    .Y(_07342_));
 sg13g2_o21ai_1 _37931_ (.B1(_07341_),
    .Y(_07343_),
    .A1(_07240_),
    .A2(_07332_));
 sg13g2_nand2_1 _37932_ (.Y(_07344_),
    .A(_07033_),
    .B(_07042_));
 sg13g2_inv_1 _37933_ (.Y(_07345_),
    .A(_07344_));
 sg13g2_nand3_1 _37934_ (.B(_07024_),
    .C(_07344_),
    .A(_07012_),
    .Y(_07346_));
 sg13g2_nand3_1 _37935_ (.B(_07023_),
    .C(_07346_),
    .A(_07011_),
    .Y(_07347_));
 sg13g2_nand3_1 _37936_ (.B(_07003_),
    .C(_07347_),
    .A(_06984_),
    .Y(_07348_));
 sg13g2_nand2_1 _37937_ (.Y(_07349_),
    .A(_06994_),
    .B(_07001_));
 sg13g2_a22oi_1 _37938_ (.Y(_07350_),
    .B1(_06984_),
    .B2(_07349_),
    .A2(_06975_),
    .A1(net5823));
 sg13g2_nand3_1 _37939_ (.B(_07348_),
    .C(_07350_),
    .A(_06982_),
    .Y(_07351_));
 sg13g2_a21o_1 _37940_ (.A2(_07136_),
    .A1(net5822),
    .B1(_07126_),
    .X(_07352_));
 sg13g2_o21ai_1 _37941_ (.B1(_07118_),
    .Y(_07353_),
    .A1(net5871),
    .A2(_07110_));
 sg13g2_a21oi_2 _37942_ (.B1(_07353_),
    .Y(_07354_),
    .A2(_07352_),
    .A1(_07120_));
 sg13g2_o21ai_1 _37943_ (.B1(_07097_),
    .Y(_07355_),
    .A1(net5867),
    .A2(_07089_));
 sg13g2_a221oi_1 _37944_ (.B2(_07355_),
    .C1(_07075_),
    .B1(_07078_),
    .A1(net5821),
    .Y(_07356_),
    .A2(_07062_));
 sg13g2_o21ai_1 _37945_ (.B1(_07356_),
    .Y(_07357_),
    .A1(_07100_),
    .A2(_07354_));
 sg13g2_a221oi_1 _37946_ (.B2(_07046_),
    .C1(_07351_),
    .B1(_07357_),
    .A1(_07141_),
    .Y(_07358_),
    .A2(_07343_));
 sg13g2_a21oi_2 _37947_ (.B1(_04796_),
    .Y(_07359_),
    .A2(_04957_),
    .A1(_04815_));
 sg13g2_nor2_1 _37948_ (.A(_04784_),
    .B(_07359_),
    .Y(_07360_));
 sg13g2_a21oi_2 _37949_ (.B1(_04787_),
    .Y(_07361_),
    .A2(_07359_),
    .A1(_04782_));
 sg13g2_o21ai_1 _37950_ (.B1(_04792_),
    .Y(_07362_),
    .A1(_04779_),
    .A2(_07361_));
 sg13g2_xnor2_1 _37951_ (.Y(_07363_),
    .A(_04103_),
    .B(_07362_));
 sg13g2_o21ai_1 _37952_ (.B1(_04394_),
    .Y(_07364_),
    .A1(_04202_),
    .A2(_04367_));
 sg13g2_nand2_1 _37953_ (.Y(_07365_),
    .A(_04150_),
    .B(_07364_));
 sg13g2_a21oi_1 _37954_ (.A1(_04151_),
    .A2(_07364_),
    .Y(_07366_),
    .B1(_04171_));
 sg13g2_a21oi_2 _37955_ (.B1(_04177_),
    .Y(_07367_),
    .A2(_07364_),
    .A1(_04153_));
 sg13g2_nor2b_1 _37956_ (.A(_07367_),
    .B_N(_04124_),
    .Y(_07368_));
 sg13g2_nand2b_1 _37957_ (.Y(_07369_),
    .B(_04124_),
    .A_N(_07367_));
 sg13g2_o21ai_1 _37958_ (.B1(_04158_),
    .Y(_07370_),
    .A1(_04116_),
    .A2(_07369_));
 sg13g2_nand2_1 _37959_ (.Y(_07371_),
    .A(_04107_),
    .B(_07370_));
 sg13g2_nand2b_1 _37960_ (.Y(_07372_),
    .B(_07370_),
    .A_N(_04108_));
 sg13g2_nand3_1 _37961_ (.B(_04162_),
    .C(_07372_),
    .A(_04103_),
    .Y(_07373_));
 sg13g2_a21o_1 _37962_ (.A2(_07372_),
    .A1(_04162_),
    .B1(_04103_),
    .X(_07374_));
 sg13g2_nand3_1 _37963_ (.B(_07373_),
    .C(_07374_),
    .A(net7391),
    .Y(_07375_));
 sg13g2_a21oi_1 _37964_ (.A1(net7223),
    .A2(\u_inv.d_next[62] ),
    .Y(_07376_),
    .B1(net6338));
 sg13g2_a22oi_1 _37965_ (.Y(_07377_),
    .B1(_07375_),
    .B2(_07376_),
    .A2(_07363_),
    .A1(net6338));
 sg13g2_nand2_1 _37966_ (.Y(_07378_),
    .A(net5815),
    .B(_07377_));
 sg13g2_xnor2_1 _37967_ (.Y(_07379_),
    .A(net5816),
    .B(_07377_));
 sg13g2_a21o_1 _37968_ (.A2(_07374_),
    .A1(_04102_),
    .B1(_04101_),
    .X(_07380_));
 sg13g2_nand3_1 _37969_ (.B(_04102_),
    .C(_07374_),
    .A(_04101_),
    .Y(_07381_));
 sg13g2_nand3_1 _37970_ (.B(_07380_),
    .C(_07381_),
    .A(net7375),
    .Y(_07382_));
 sg13g2_a21oi_1 _37971_ (.A1(net7223),
    .A2(\u_inv.d_next[63] ),
    .Y(_07383_),
    .B1(net6339));
 sg13g2_a21oi_1 _37972_ (.A1(_04103_),
    .A2(_07362_),
    .Y(_07384_),
    .B1(_04788_));
 sg13g2_or2_1 _37973_ (.X(_07385_),
    .B(_07384_),
    .A(_04101_));
 sg13g2_a21oi_1 _37974_ (.A1(_04101_),
    .A2(_07384_),
    .Y(_07386_),
    .B1(net6248));
 sg13g2_a22oi_1 _37975_ (.Y(_07387_),
    .B1(_07385_),
    .B2(_07386_),
    .A2(_07383_),
    .A1(_07382_));
 sg13g2_nand2_1 _37976_ (.Y(_07388_),
    .A(net5816),
    .B(_07387_));
 sg13g2_xnor2_1 _37977_ (.Y(_07389_),
    .A(net5816),
    .B(_07387_));
 sg13g2_nand3_1 _37978_ (.B(_04106_),
    .C(_07371_),
    .A(_04105_),
    .Y(_07390_));
 sg13g2_nand4_1 _37979_ (.B(_04160_),
    .C(_07372_),
    .A(net7391),
    .Y(_07391_),
    .D(_07390_));
 sg13g2_a21oi_1 _37980_ (.A1(net7230),
    .A2(\u_inv.d_next[61] ),
    .Y(_07392_),
    .B1(net6339));
 sg13g2_o21ai_1 _37981_ (.B1(_04790_),
    .Y(_07393_),
    .A1(_04107_),
    .A2(_07361_));
 sg13g2_xnor2_1 _37982_ (.Y(_07394_),
    .A(_04105_),
    .B(_07393_));
 sg13g2_a22oi_1 _37983_ (.Y(_07395_),
    .B1(_07394_),
    .B2(net6339),
    .A2(_07392_),
    .A1(_07391_));
 sg13g2_xnor2_1 _37984_ (.Y(_07396_),
    .A(net5865),
    .B(_07395_));
 sg13g2_o21ai_1 _37985_ (.B1(net6349),
    .Y(_07397_),
    .A1(_04107_),
    .A2(_07361_));
 sg13g2_a21o_1 _37986_ (.A2(_07361_),
    .A1(_04107_),
    .B1(_07397_),
    .X(_07398_));
 sg13g2_nor2_1 _37987_ (.A(_04107_),
    .B(_07370_),
    .Y(_07399_));
 sg13g2_nor2_1 _37988_ (.A(net7230),
    .B(_07399_),
    .Y(_07400_));
 sg13g2_a22oi_1 _37989_ (.Y(_07401_),
    .B1(_07371_),
    .B2(_07400_),
    .A2(\u_inv.d_next[60] ),
    .A1(net7230));
 sg13g2_o21ai_1 _37990_ (.B1(_07398_),
    .Y(_07402_),
    .A1(net6339),
    .A2(_07401_));
 sg13g2_nand2_1 _37991_ (.Y(_07403_),
    .A(net5817),
    .B(_07402_));
 sg13g2_inv_1 _37992_ (.Y(_07404_),
    .A(_07403_));
 sg13g2_xnor2_1 _37993_ (.Y(_07405_),
    .A(net5866),
    .B(_07402_));
 sg13g2_nand2_1 _37994_ (.Y(_07406_),
    .A(_07396_),
    .B(_07405_));
 sg13g2_or3_1 _37995_ (.A(_07379_),
    .B(_07389_),
    .C(_07406_),
    .X(_07407_));
 sg13g2_o21ai_1 _37996_ (.B1(_04114_),
    .Y(_07408_),
    .A1(_04156_),
    .A2(_07368_));
 sg13g2_a21oi_1 _37997_ (.A1(_04112_),
    .A2(_07408_),
    .Y(_07409_),
    .B1(_04111_));
 sg13g2_nand3_1 _37998_ (.B(_04112_),
    .C(_07408_),
    .A(_04111_),
    .Y(_07410_));
 sg13g2_nor2_1 _37999_ (.A(net7223),
    .B(_07409_),
    .Y(_07411_));
 sg13g2_a221oi_1 _38000_ (.B2(_07411_),
    .C1(net6338),
    .B1(_07410_),
    .A1(net7224),
    .Y(_07412_),
    .A2(\u_inv.d_next[59] ));
 sg13g2_o21ai_1 _38001_ (.B1(_04113_),
    .Y(_07413_),
    .A1(_04784_),
    .A2(_07359_));
 sg13g2_a21oi_1 _38002_ (.A1(_04785_),
    .A2(_07413_),
    .Y(_07414_),
    .B1(_04111_));
 sg13g2_nand3_1 _38003_ (.B(_04785_),
    .C(_07413_),
    .A(_04111_),
    .Y(_07415_));
 sg13g2_nor2_1 _38004_ (.A(net6248),
    .B(_07414_),
    .Y(_07416_));
 sg13g2_a21o_2 _38005_ (.A2(_07416_),
    .A1(_07415_),
    .B1(_07412_),
    .X(_07417_));
 sg13g2_xnor2_1 _38006_ (.Y(_07418_),
    .A(net5865),
    .B(_07417_));
 sg13g2_xnor2_1 _38007_ (.Y(_07419_),
    .A(_04113_),
    .B(_07360_));
 sg13g2_nand3b_1 _38008_ (.B(_07369_),
    .C(_04113_),
    .Y(_07420_),
    .A_N(_04156_));
 sg13g2_nand3_1 _38009_ (.B(_07408_),
    .C(_07420_),
    .A(net7375),
    .Y(_07421_));
 sg13g2_nand2_1 _38010_ (.Y(_07422_),
    .A(net7224),
    .B(\u_inv.d_next[58] ));
 sg13g2_a21oi_1 _38011_ (.A1(_07421_),
    .A2(_07422_),
    .Y(_07423_),
    .B1(net6338));
 sg13g2_a21oi_2 _38012_ (.B1(_07423_),
    .Y(_07424_),
    .A2(_07419_),
    .A1(net6338));
 sg13g2_nor2_1 _38013_ (.A(net5865),
    .B(_07424_),
    .Y(_07425_));
 sg13g2_xnor2_1 _38014_ (.Y(_07426_),
    .A(net5865),
    .B(_07424_));
 sg13g2_or2_1 _38015_ (.X(_07427_),
    .B(_07426_),
    .A(_07418_));
 sg13g2_nand2_1 _38016_ (.Y(_07428_),
    .A(_04123_),
    .B(_04958_));
 sg13g2_xnor2_1 _38017_ (.Y(_07429_),
    .A(_04123_),
    .B(_04958_));
 sg13g2_xnor2_1 _38018_ (.Y(_07430_),
    .A(_04122_),
    .B(_07367_));
 sg13g2_nand2_1 _38019_ (.Y(_07431_),
    .A(net7375),
    .B(_07430_));
 sg13g2_a21oi_1 _38020_ (.A1(net7224),
    .A2(\u_inv.d_next[56] ),
    .Y(_07432_),
    .B1(net6338));
 sg13g2_a22oi_1 _38021_ (.Y(_07433_),
    .B1(_07431_),
    .B2(_07432_),
    .A2(_07429_),
    .A1(net6340));
 sg13g2_xnor2_1 _38022_ (.Y(_07434_),
    .A(net5865),
    .B(_07433_));
 sg13g2_and2_1 _38023_ (.A(_04783_),
    .B(_07428_),
    .X(_07435_));
 sg13g2_xnor2_1 _38024_ (.Y(_07436_),
    .A(_04120_),
    .B(_07435_));
 sg13g2_o21ai_1 _38025_ (.B1(_04121_),
    .Y(_07437_),
    .A1(_04123_),
    .A2(_07367_));
 sg13g2_a21oi_1 _38026_ (.A1(_04120_),
    .A2(_07437_),
    .Y(_07438_),
    .B1(net7224));
 sg13g2_o21ai_1 _38027_ (.B1(_07438_),
    .Y(_07439_),
    .A1(_04120_),
    .A2(_07437_));
 sg13g2_a21oi_1 _38028_ (.A1(net7224),
    .A2(\u_inv.d_next[57] ),
    .Y(_07440_),
    .B1(net6338));
 sg13g2_a22oi_1 _38029_ (.Y(_07441_),
    .B1(_07439_),
    .B2(_07440_),
    .A2(_07436_),
    .A1(net6338));
 sg13g2_xnor2_1 _38030_ (.Y(_07442_),
    .A(net5815),
    .B(_07441_));
 sg13g2_inv_1 _38031_ (.Y(_07443_),
    .A(_07442_));
 sg13g2_nand2_1 _38032_ (.Y(_07444_),
    .A(_07434_),
    .B(_07443_));
 sg13g2_inv_1 _38033_ (.Y(_07445_),
    .A(_07444_));
 sg13g2_nor3_1 _38034_ (.A(_07407_),
    .B(_07427_),
    .C(_07444_),
    .Y(_07446_));
 sg13g2_nor3_1 _38035_ (.A(_04128_),
    .B(_04132_),
    .C(_07366_),
    .Y(_07447_));
 sg13g2_or3_1 _38036_ (.A(_04138_),
    .B(_04172_),
    .C(_07447_),
    .X(_07448_));
 sg13g2_o21ai_1 _38037_ (.B1(_04138_),
    .Y(_07449_),
    .A1(_04172_),
    .A2(_07447_));
 sg13g2_nand3_1 _38038_ (.B(_07448_),
    .C(_07449_),
    .A(net7375),
    .Y(_07450_));
 sg13g2_o21ai_1 _38039_ (.B1(_07450_),
    .Y(_07451_),
    .A1(net7375),
    .A2(_18163_));
 sg13g2_o21ai_1 _38040_ (.B1(_04816_),
    .Y(_07452_),
    .A1(_04862_),
    .A2(_04955_));
 sg13g2_nand2_1 _38041_ (.Y(_07453_),
    .A(_04800_),
    .B(_07452_));
 sg13g2_a21o_1 _38042_ (.A2(_07452_),
    .A1(_04800_),
    .B1(_04803_),
    .X(_07454_));
 sg13g2_and2_1 _38043_ (.A(_04806_),
    .B(_07454_),
    .X(_07455_));
 sg13g2_nand2b_1 _38044_ (.Y(_07456_),
    .B(_04128_),
    .A_N(_07455_));
 sg13g2_a221oi_1 _38045_ (.B2(_07454_),
    .C1(_04127_),
    .B1(_04806_),
    .A1(_04130_),
    .Y(_07457_),
    .A2(_04131_));
 sg13g2_or3_1 _38046_ (.A(_04137_),
    .B(_04811_),
    .C(_07457_),
    .X(_07458_));
 sg13g2_o21ai_1 _38047_ (.B1(_04137_),
    .Y(_07459_),
    .A1(_04811_),
    .A2(_07457_));
 sg13g2_and2_1 _38048_ (.A(net6340),
    .B(_07459_),
    .X(_07460_));
 sg13g2_a22oi_1 _38049_ (.Y(_07461_),
    .B1(_07458_),
    .B2(_07460_),
    .A2(_07451_),
    .A1(net6249));
 sg13g2_nor2_1 _38050_ (.A(net5865),
    .B(_07461_),
    .Y(_07462_));
 sg13g2_xnor2_1 _38051_ (.Y(_07463_),
    .A(net5865),
    .B(_07461_));
 sg13g2_inv_1 _38052_ (.Y(_07464_),
    .A(_07463_));
 sg13g2_a21o_1 _38053_ (.A2(_07459_),
    .A1(_04807_),
    .B1(_04134_),
    .X(_07465_));
 sg13g2_nand3_1 _38054_ (.B(_04807_),
    .C(_07459_),
    .A(_04134_),
    .Y(_07466_));
 sg13g2_nand3_1 _38055_ (.B(_07465_),
    .C(_07466_),
    .A(net6340),
    .Y(_07467_));
 sg13g2_nand3_1 _38056_ (.B(_04136_),
    .C(_07449_),
    .A(_04134_),
    .Y(_07468_));
 sg13g2_a21oi_1 _38057_ (.A1(_04136_),
    .A2(_07449_),
    .Y(_07469_),
    .B1(_04134_));
 sg13g2_nand2_1 _38058_ (.Y(_07470_),
    .A(net7375),
    .B(_07468_));
 sg13g2_a21oi_1 _38059_ (.A1(net7223),
    .A2(\u_inv.d_next[55] ),
    .Y(_07471_),
    .B1(net6340));
 sg13g2_o21ai_1 _38060_ (.B1(_07471_),
    .Y(_07472_),
    .A1(_07469_),
    .A2(_07470_));
 sg13g2_and2_1 _38061_ (.A(_07467_),
    .B(_07472_),
    .X(_07473_));
 sg13g2_a21oi_1 _38062_ (.A1(_07467_),
    .A2(_07472_),
    .Y(_07474_),
    .B1(net5815));
 sg13g2_and3_1 _38063_ (.X(_07475_),
    .A(net5815),
    .B(_07467_),
    .C(_07472_));
 sg13g2_nor2_1 _38064_ (.A(_07474_),
    .B(_07475_),
    .Y(_07476_));
 sg13g2_nor3_1 _38065_ (.A(_07463_),
    .B(_07474_),
    .C(_07475_),
    .Y(_07477_));
 sg13g2_a21oi_1 _38066_ (.A1(_04809_),
    .A2(_07456_),
    .Y(_07478_),
    .B1(_04132_));
 sg13g2_nand3_1 _38067_ (.B(_04809_),
    .C(_07456_),
    .A(_04132_),
    .Y(_07479_));
 sg13g2_nor2_1 _38068_ (.A(net6249),
    .B(_07478_),
    .Y(_07480_));
 sg13g2_nor2_1 _38069_ (.A(_04128_),
    .B(_07366_),
    .Y(_07481_));
 sg13g2_nor2_1 _38070_ (.A(_04126_),
    .B(_07481_),
    .Y(_07482_));
 sg13g2_o21ai_1 _38071_ (.B1(net7375),
    .Y(_07483_),
    .A1(_04132_),
    .A2(_07482_));
 sg13g2_a21oi_1 _38072_ (.A1(_04132_),
    .A2(_07482_),
    .Y(_07484_),
    .B1(_07483_));
 sg13g2_nand2_1 _38073_ (.Y(_07485_),
    .A(net7223),
    .B(\u_inv.d_next[53] ));
 sg13g2_nor2_1 _38074_ (.A(net6340),
    .B(_07484_),
    .Y(_07486_));
 sg13g2_a22oi_1 _38075_ (.Y(_07487_),
    .B1(_07485_),
    .B2(_07486_),
    .A2(_07480_),
    .A1(_07479_));
 sg13g2_nor2_1 _38076_ (.A(net5815),
    .B(_07487_),
    .Y(_07488_));
 sg13g2_xnor2_1 _38077_ (.Y(_07489_),
    .A(net5860),
    .B(_07487_));
 sg13g2_xnor2_1 _38078_ (.Y(_07490_),
    .A(_04127_),
    .B(_07455_));
 sg13g2_a21oi_1 _38079_ (.A1(_04128_),
    .A2(_07366_),
    .Y(_07491_),
    .B1(net7223));
 sg13g2_nand2b_1 _38080_ (.Y(_07492_),
    .B(_07491_),
    .A_N(_07481_));
 sg13g2_a21oi_1 _38081_ (.A1(net7223),
    .A2(\u_inv.d_next[52] ),
    .Y(_07493_),
    .B1(net6340));
 sg13g2_a22oi_1 _38082_ (.Y(_07494_),
    .B1(_07492_),
    .B2(_07493_),
    .A2(_07490_),
    .A1(net6340));
 sg13g2_nand2_1 _38083_ (.Y(_07495_),
    .A(net5815),
    .B(_07494_));
 sg13g2_xnor2_1 _38084_ (.Y(_07496_),
    .A(net5860),
    .B(_07494_));
 sg13g2_xnor2_1 _38085_ (.Y(_07497_),
    .A(_04145_),
    .B(_07453_));
 sg13g2_nand3_1 _38086_ (.B(_04168_),
    .C(_07365_),
    .A(_04145_),
    .Y(_07498_));
 sg13g2_a21oi_1 _38087_ (.A1(_04168_),
    .A2(_07365_),
    .Y(_07499_),
    .B1(_04145_));
 sg13g2_nand3b_1 _38088_ (.B(net7373),
    .C(_07498_),
    .Y(_07500_),
    .A_N(_07499_));
 sg13g2_a21oi_1 _38089_ (.A1(net7221),
    .A2(net7298),
    .Y(_07501_),
    .B1(net6335));
 sg13g2_a22oi_1 _38090_ (.Y(_07502_),
    .B1(_07500_),
    .B2(_07501_),
    .A2(_07497_),
    .A1(net6335));
 sg13g2_and2_1 _38091_ (.A(net5811),
    .B(_07502_),
    .X(_07503_));
 sg13g2_xnor2_1 _38092_ (.Y(_07504_),
    .A(net5811),
    .B(_07502_));
 sg13g2_o21ai_1 _38093_ (.B1(_04142_),
    .Y(_07505_),
    .A1(_04143_),
    .A2(_07499_));
 sg13g2_nor3_1 _38094_ (.A(_04142_),
    .B(_04143_),
    .C(_07499_),
    .Y(_07506_));
 sg13g2_nand2_1 _38095_ (.Y(_07507_),
    .A(net7375),
    .B(_07505_));
 sg13g2_a21oi_1 _38096_ (.A1(net7223),
    .A2(\u_inv.d_next[51] ),
    .Y(_07508_),
    .B1(net6336));
 sg13g2_o21ai_1 _38097_ (.B1(_07508_),
    .Y(_07509_),
    .A1(_07506_),
    .A2(_07507_));
 sg13g2_a21oi_1 _38098_ (.A1(_04145_),
    .A2(_07453_),
    .Y(_07510_),
    .B1(_04804_));
 sg13g2_and2_1 _38099_ (.A(_04141_),
    .B(_07510_),
    .X(_07511_));
 sg13g2_o21ai_1 _38100_ (.B1(net6336),
    .Y(_07512_),
    .A1(_04141_),
    .A2(_07510_));
 sg13g2_o21ai_1 _38101_ (.B1(_07509_),
    .Y(_07513_),
    .A1(_07511_),
    .A2(_07512_));
 sg13g2_nor2_1 _38102_ (.A(net5860),
    .B(_07513_),
    .Y(_07514_));
 sg13g2_xnor2_1 _38103_ (.Y(_07515_),
    .A(net5811),
    .B(_07513_));
 sg13g2_nor2b_1 _38104_ (.A(_07504_),
    .B_N(_07515_),
    .Y(_07516_));
 sg13g2_a21oi_1 _38105_ (.A1(_04149_),
    .A2(_07364_),
    .Y(_07517_),
    .B1(_04146_));
 sg13g2_nand2_1 _38106_ (.Y(_07518_),
    .A(_04148_),
    .B(_07517_));
 sg13g2_nor2_1 _38107_ (.A(net7221),
    .B(_04166_),
    .Y(_07519_));
 sg13g2_nand3_1 _38108_ (.B(_07518_),
    .C(_07519_),
    .A(_07365_),
    .Y(_07520_));
 sg13g2_nand2_1 _38109_ (.Y(_07521_),
    .A(net7221),
    .B(\u_inv.d_next[49] ));
 sg13g2_a21oi_1 _38110_ (.A1(_07520_),
    .A2(_07521_),
    .Y(_07522_),
    .B1(net6335));
 sg13g2_or2_1 _38111_ (.X(_07523_),
    .B(_04956_),
    .A(_04149_));
 sg13g2_nand2_1 _38112_ (.Y(_07524_),
    .A(_04798_),
    .B(_07523_));
 sg13g2_xnor2_1 _38113_ (.Y(_07525_),
    .A(_04146_),
    .B(_07524_));
 sg13g2_a21oi_2 _38114_ (.B1(_07522_),
    .Y(_07526_),
    .A2(_07525_),
    .A1(net6335));
 sg13g2_nand2_1 _38115_ (.Y(_07527_),
    .A(net5860),
    .B(_07526_));
 sg13g2_xnor2_1 _38116_ (.Y(_07528_),
    .A(net5811),
    .B(_07526_));
 sg13g2_xnor2_1 _38117_ (.Y(_07529_),
    .A(_04149_),
    .B(_07364_));
 sg13g2_nor2_1 _38118_ (.A(net7367),
    .B(\u_inv.d_next[48] ),
    .Y(_07530_));
 sg13g2_a21oi_1 _38119_ (.A1(net7373),
    .A2(_07529_),
    .Y(_07531_),
    .B1(_07530_));
 sg13g2_a21oi_1 _38120_ (.A1(_04149_),
    .A2(_04956_),
    .Y(_07532_),
    .B1(net6247));
 sg13g2_a22oi_1 _38121_ (.Y(_07533_),
    .B1(_07532_),
    .B2(_07523_),
    .A2(_07531_),
    .A1(net6247));
 sg13g2_nor2_1 _38122_ (.A(net5861),
    .B(_07533_),
    .Y(_07534_));
 sg13g2_xnor2_1 _38123_ (.Y(_07535_),
    .A(net5810),
    .B(_07533_));
 sg13g2_inv_1 _38124_ (.Y(_07536_),
    .A(_07535_));
 sg13g2_and3_1 _38125_ (.X(_07537_),
    .A(_07516_),
    .B(_07528_),
    .C(_07535_));
 sg13g2_inv_1 _38126_ (.Y(_07538_),
    .A(_07537_));
 sg13g2_nand4_1 _38127_ (.B(_07489_),
    .C(_07496_),
    .A(_07477_),
    .Y(_07539_),
    .D(_07537_));
 sg13g2_nor4_1 _38128_ (.A(_07407_),
    .B(_07427_),
    .C(_07444_),
    .D(_07539_),
    .Y(_07540_));
 sg13g2_o21ai_1 _38129_ (.B1(_04952_),
    .Y(_07541_),
    .A1(_04947_),
    .A2(_04949_));
 sg13g2_and2_1 _38130_ (.A(_04844_),
    .B(_07541_),
    .X(_07542_));
 sg13g2_a21oi_1 _38131_ (.A1(_04844_),
    .A2(_07541_),
    .Y(_07543_),
    .B1(_04819_));
 sg13g2_nand2b_1 _38132_ (.Y(_07544_),
    .B(_04847_),
    .A_N(_07543_));
 sg13g2_o21ai_1 _38133_ (.B1(_04822_),
    .Y(_07545_),
    .A1(_04848_),
    .A2(_07543_));
 sg13g2_and2_1 _38134_ (.A(_04858_),
    .B(_07545_),
    .X(_07546_));
 sg13g2_a221oi_1 _38135_ (.B2(_07545_),
    .C1(_04179_),
    .B1(_04858_),
    .A1(_04180_),
    .Y(_07547_),
    .A2(_04182_));
 sg13g2_o21ai_1 _38136_ (.B1(_04189_),
    .Y(_07548_),
    .A1(_04851_),
    .A2(_07547_));
 sg13g2_or3_1 _38137_ (.A(_04189_),
    .B(_04851_),
    .C(_07547_),
    .X(_07549_));
 sg13g2_nand2_1 _38138_ (.Y(_07550_),
    .A(_07548_),
    .B(_07549_));
 sg13g2_nand2_1 _38139_ (.Y(_07551_),
    .A(_04367_),
    .B(_04380_));
 sg13g2_a21oi_1 _38140_ (.A1(_04367_),
    .A2(_04380_),
    .Y(_07552_),
    .B1(_04200_));
 sg13g2_nand2b_1 _38141_ (.Y(_07553_),
    .B(_07552_),
    .A_N(_04195_));
 sg13g2_and2_1 _38142_ (.A(_04391_),
    .B(_07553_),
    .X(_07554_));
 sg13g2_o21ai_1 _38143_ (.B1(_04383_),
    .Y(_07555_),
    .A1(_04184_),
    .A2(_07554_));
 sg13g2_xnor2_1 _38144_ (.Y(_07556_),
    .A(_04189_),
    .B(_07555_));
 sg13g2_nand2_1 _38145_ (.Y(_07557_),
    .A(net7221),
    .B(\u_inv.d_next[46] ));
 sg13g2_a21oi_1 _38146_ (.A1(net7373),
    .A2(_07556_),
    .Y(_07558_),
    .B1(net6335));
 sg13g2_a22oi_1 _38147_ (.Y(_07559_),
    .B1(_07557_),
    .B2(_07558_),
    .A2(_07550_),
    .A1(net6335));
 sg13g2_nand2_1 _38148_ (.Y(_07560_),
    .A(net5810),
    .B(_07559_));
 sg13g2_xnor2_1 _38149_ (.Y(_07561_),
    .A(net5860),
    .B(_07559_));
 sg13g2_xnor2_1 _38150_ (.Y(_07562_),
    .A(net5810),
    .B(_07559_));
 sg13g2_a21o_1 _38151_ (.A2(_07548_),
    .A1(_04853_),
    .B1(_04185_),
    .X(_07563_));
 sg13g2_nand3_1 _38152_ (.B(_04853_),
    .C(_07548_),
    .A(_04185_),
    .Y(_07564_));
 sg13g2_nand3_1 _38153_ (.B(_07563_),
    .C(_07564_),
    .A(net6335),
    .Y(_07565_));
 sg13g2_a21oi_1 _38154_ (.A1(_04186_),
    .A2(_07555_),
    .Y(_07566_),
    .B1(_04187_));
 sg13g2_o21ai_1 _38155_ (.B1(net7373),
    .Y(_07567_),
    .A1(_04185_),
    .A2(_07566_));
 sg13g2_a21oi_1 _38156_ (.A1(_04185_),
    .A2(_07566_),
    .Y(_07568_),
    .B1(_07567_));
 sg13g2_o21ai_1 _38157_ (.B1(net6247),
    .Y(_07569_),
    .A1(net7374),
    .A2(_18165_));
 sg13g2_o21ai_1 _38158_ (.B1(_07565_),
    .Y(_07570_),
    .A1(_07568_),
    .A2(_07569_));
 sg13g2_nand2b_1 _38159_ (.Y(_07571_),
    .B(net5810),
    .A_N(_07570_));
 sg13g2_xnor2_1 _38160_ (.Y(_07572_),
    .A(net5810),
    .B(_07570_));
 sg13g2_o21ai_1 _38161_ (.B1(_04849_),
    .Y(_07573_),
    .A1(_04179_),
    .A2(_07546_));
 sg13g2_and2_1 _38162_ (.A(_04183_),
    .B(_07573_),
    .X(_07574_));
 sg13g2_o21ai_1 _38163_ (.B1(net6336),
    .Y(_07575_),
    .A1(_04183_),
    .A2(_07573_));
 sg13g2_nor2b_1 _38164_ (.A(_07554_),
    .B_N(_04179_),
    .Y(_07576_));
 sg13g2_a21o_1 _38165_ (.A2(\u_inv.d_reg[44] ),
    .A1(\u_inv.d_next[44] ),
    .B1(_07576_),
    .X(_07577_));
 sg13g2_and2_1 _38166_ (.A(_04183_),
    .B(_07577_),
    .X(_07578_));
 sg13g2_o21ai_1 _38167_ (.B1(net7374),
    .Y(_07579_),
    .A1(_04183_),
    .A2(_07577_));
 sg13g2_a21oi_1 _38168_ (.A1(net7221),
    .A2(\u_inv.d_next[45] ),
    .Y(_07580_),
    .B1(net6336));
 sg13g2_o21ai_1 _38169_ (.B1(_07580_),
    .Y(_07581_),
    .A1(_07578_),
    .A2(_07579_));
 sg13g2_o21ai_1 _38170_ (.B1(_07581_),
    .Y(_07582_),
    .A1(_07574_),
    .A2(_07575_));
 sg13g2_nor2_1 _38171_ (.A(net5860),
    .B(_07582_),
    .Y(_07583_));
 sg13g2_and2_1 _38172_ (.A(net5860),
    .B(_07582_),
    .X(_07584_));
 sg13g2_xnor2_1 _38173_ (.Y(_07585_),
    .A(net5810),
    .B(_07582_));
 sg13g2_xor2_1 _38174_ (.B(_07554_),
    .A(_04179_),
    .X(_07586_));
 sg13g2_o21ai_1 _38175_ (.B1(net6247),
    .Y(_07587_),
    .A1(net7373),
    .A2(\u_inv.d_next[44] ));
 sg13g2_a21o_1 _38176_ (.A2(_07586_),
    .A1(net7373),
    .B1(_07587_),
    .X(_07588_));
 sg13g2_xnor2_1 _38177_ (.Y(_07589_),
    .A(_04179_),
    .B(_07546_));
 sg13g2_o21ai_1 _38178_ (.B1(_07588_),
    .Y(_07590_),
    .A1(net6247),
    .A2(_07589_));
 sg13g2_nand2_1 _38179_ (.Y(_07591_),
    .A(net5810),
    .B(_07590_));
 sg13g2_xnor2_1 _38180_ (.Y(_07592_),
    .A(net5810),
    .B(_07590_));
 sg13g2_inv_1 _38181_ (.Y(_07593_),
    .A(_07592_));
 sg13g2_and2_1 _38182_ (.A(_07585_),
    .B(_07593_),
    .X(_07594_));
 sg13g2_a21oi_1 _38183_ (.A1(_04194_),
    .A2(_07544_),
    .Y(_07595_),
    .B1(_04855_));
 sg13g2_or2_1 _38184_ (.X(_07596_),
    .B(_07595_),
    .A(_04191_));
 sg13g2_a21oi_1 _38185_ (.A1(_04191_),
    .A2(_07595_),
    .Y(_07597_),
    .B1(net6242));
 sg13g2_o21ai_1 _38186_ (.B1(_04193_),
    .Y(_07598_),
    .A1(_04388_),
    .A2(_07552_));
 sg13g2_nand3_1 _38187_ (.B(_04192_),
    .C(_07598_),
    .A(_04191_),
    .Y(_07599_));
 sg13g2_a21oi_1 _38188_ (.A1(_04192_),
    .A2(_07598_),
    .Y(_07600_),
    .B1(_04191_));
 sg13g2_nor2_1 _38189_ (.A(net7219),
    .B(_07600_),
    .Y(_07601_));
 sg13g2_a221oi_1 _38190_ (.B2(_07601_),
    .C1(net6331),
    .B1(_07599_),
    .A1(net7219),
    .Y(_07602_),
    .A2(\u_inv.d_next[43] ));
 sg13g2_a21o_2 _38191_ (.A2(_07597_),
    .A1(_07596_),
    .B1(_07602_),
    .X(_07603_));
 sg13g2_nor2_1 _38192_ (.A(net5860),
    .B(_07603_),
    .Y(_07604_));
 sg13g2_xnor2_1 _38193_ (.Y(_07605_),
    .A(net5859),
    .B(_07603_));
 sg13g2_or3_1 _38194_ (.A(_04193_),
    .B(_04388_),
    .C(_07552_),
    .X(_07606_));
 sg13g2_nand3_1 _38195_ (.B(_07598_),
    .C(_07606_),
    .A(net7367),
    .Y(_07607_));
 sg13g2_xnor2_1 _38196_ (.Y(_07608_),
    .A(_04194_),
    .B(_07544_));
 sg13g2_a21oi_1 _38197_ (.A1(net7219),
    .A2(\u_inv.d_next[42] ),
    .Y(_07609_),
    .B1(net6331));
 sg13g2_a22oi_1 _38198_ (.Y(_07610_),
    .B1(_07609_),
    .B2(_07607_),
    .A2(_07608_),
    .A1(net6331));
 sg13g2_nand2_1 _38199_ (.Y(_07611_),
    .A(net5809),
    .B(_07610_));
 sg13g2_xnor2_1 _38200_ (.Y(_07612_),
    .A(net5812),
    .B(_07610_));
 sg13g2_or2_1 _38201_ (.X(_07613_),
    .B(_07612_),
    .A(_07605_));
 sg13g2_inv_1 _38202_ (.Y(_07614_),
    .A(_07613_));
 sg13g2_xnor2_1 _38203_ (.Y(_07615_),
    .A(_04199_),
    .B(_07551_));
 sg13g2_o21ai_1 _38204_ (.B1(net6242),
    .Y(_07616_),
    .A1(net7373),
    .A2(\u_inv.d_next[40] ));
 sg13g2_a21oi_1 _38205_ (.A1(net7373),
    .A2(_07615_),
    .Y(_07617_),
    .B1(_07616_));
 sg13g2_o21ai_1 _38206_ (.B1(net6331),
    .Y(_07618_),
    .A1(_04199_),
    .A2(_07542_));
 sg13g2_a21oi_1 _38207_ (.A1(_04199_),
    .A2(_07542_),
    .Y(_07619_),
    .B1(_07618_));
 sg13g2_nor2_2 _38208_ (.A(_07617_),
    .B(_07619_),
    .Y(_07620_));
 sg13g2_nor2_1 _38209_ (.A(net5859),
    .B(_07620_),
    .Y(_07621_));
 sg13g2_xnor2_1 _38210_ (.Y(_07622_),
    .A(net5812),
    .B(_07620_));
 sg13g2_o21ai_1 _38211_ (.B1(_04845_),
    .Y(_07623_),
    .A1(_04199_),
    .A2(_07542_));
 sg13g2_a21oi_1 _38212_ (.A1(_04197_),
    .A2(_07623_),
    .Y(_07624_),
    .B1(net6247));
 sg13g2_o21ai_1 _38213_ (.B1(_07624_),
    .Y(_07625_),
    .A1(_04197_),
    .A2(_07623_));
 sg13g2_a21o_1 _38214_ (.A2(_07551_),
    .A1(_04199_),
    .B1(_04198_),
    .X(_07626_));
 sg13g2_a21oi_1 _38215_ (.A1(_04197_),
    .A2(_07626_),
    .Y(_07627_),
    .B1(net7221));
 sg13g2_o21ai_1 _38216_ (.B1(_07627_),
    .Y(_07628_),
    .A1(_04197_),
    .A2(_07626_));
 sg13g2_a21oi_1 _38217_ (.A1(net7221),
    .A2(\u_inv.d_next[41] ),
    .Y(_07629_),
    .B1(net6335));
 sg13g2_nand2_1 _38218_ (.Y(_07630_),
    .A(_07628_),
    .B(_07629_));
 sg13g2_nand2_1 _38219_ (.Y(_07631_),
    .A(_07625_),
    .B(_07630_));
 sg13g2_xnor2_1 _38220_ (.Y(_07632_),
    .A(net5812),
    .B(_07631_));
 sg13g2_and2_1 _38221_ (.A(_07622_),
    .B(_07632_),
    .X(_07633_));
 sg13g2_nor2b_1 _38222_ (.A(_07613_),
    .B_N(_07633_),
    .Y(_07634_));
 sg13g2_nand4_1 _38223_ (.B(_07572_),
    .C(_07594_),
    .A(_07561_),
    .Y(_07635_),
    .D(_07634_));
 sg13g2_and2_1 _38224_ (.A(_04365_),
    .B(_04951_),
    .X(_07636_));
 sg13g2_a221oi_1 _38225_ (.B2(_04950_),
    .C1(_04362_),
    .B1(_04946_),
    .A1(_04363_),
    .Y(_07637_),
    .A2(_04364_));
 sg13g2_o21ai_1 _38226_ (.B1(_04828_),
    .Y(_07638_),
    .A1(_04831_),
    .A2(_07637_));
 sg13g2_nand2_2 _38227_ (.Y(_07639_),
    .A(_04833_),
    .B(_07638_));
 sg13g2_a21oi_1 _38228_ (.A1(_04826_),
    .A2(_07639_),
    .Y(_07640_),
    .B1(_04841_));
 sg13g2_xnor2_1 _38229_ (.Y(_07641_),
    .A(_04352_),
    .B(_07640_));
 sg13g2_or3_1 _38230_ (.A(_04340_),
    .B(net6995),
    .C(_04365_),
    .X(_07642_));
 sg13g2_o21ai_1 _38231_ (.B1(_04373_),
    .Y(_07643_),
    .A1(_04360_),
    .A2(_07642_));
 sg13g2_a21oi_1 _38232_ (.A1(_04346_),
    .A2(_07643_),
    .Y(_07644_),
    .B1(_04376_));
 sg13g2_nand2b_1 _38233_ (.Y(_07645_),
    .B(_04352_),
    .A_N(_07644_));
 sg13g2_a21oi_1 _38234_ (.A1(_04353_),
    .A2(_07644_),
    .Y(_07646_),
    .B1(net7211));
 sg13g2_nand2_1 _38235_ (.Y(_07647_),
    .A(_07645_),
    .B(_07646_));
 sg13g2_a21oi_1 _38236_ (.A1(net7213),
    .A2(\u_inv.d_next[38] ),
    .Y(_07648_),
    .B1(net6322));
 sg13g2_a22oi_1 _38237_ (.Y(_07649_),
    .B1(_07647_),
    .B2(_07648_),
    .A2(_07641_),
    .A1(net6322));
 sg13g2_and2_1 _38238_ (.A(net5809),
    .B(_07649_),
    .X(_07650_));
 sg13g2_xnor2_1 _38239_ (.Y(_07651_),
    .A(net5809),
    .B(_07649_));
 sg13g2_o21ai_1 _38240_ (.B1(_04837_),
    .Y(_07652_),
    .A1(_04352_),
    .A2(_07640_));
 sg13g2_and2_1 _38241_ (.A(_04350_),
    .B(_07652_),
    .X(_07653_));
 sg13g2_o21ai_1 _38242_ (.B1(net6322),
    .Y(_07654_),
    .A1(_04350_),
    .A2(_07652_));
 sg13g2_nand3_1 _38243_ (.B(_04351_),
    .C(_07645_),
    .A(_04349_),
    .Y(_07655_));
 sg13g2_a21oi_1 _38244_ (.A1(_04351_),
    .A2(_07645_),
    .Y(_07656_),
    .B1(_04349_));
 sg13g2_nand2_1 _38245_ (.Y(_07657_),
    .A(net7367),
    .B(_07655_));
 sg13g2_a21oi_1 _38246_ (.A1(net7219),
    .A2(\u_inv.d_next[39] ),
    .Y(_07658_),
    .B1(net6322));
 sg13g2_o21ai_1 _38247_ (.B1(_07658_),
    .Y(_07659_),
    .A1(_07656_),
    .A2(_07657_));
 sg13g2_o21ai_1 _38248_ (.B1(_07659_),
    .Y(_07660_),
    .A1(_07653_),
    .A2(_07654_));
 sg13g2_nor2_1 _38249_ (.A(net5859),
    .B(_07660_),
    .Y(_07661_));
 sg13g2_xnor2_1 _38250_ (.Y(_07662_),
    .A(net5859),
    .B(_07660_));
 sg13g2_nor2_1 _38251_ (.A(_07651_),
    .B(_07662_),
    .Y(_07663_));
 sg13g2_nand2_1 _38252_ (.Y(_07664_),
    .A(_04344_),
    .B(_07643_));
 sg13g2_xnor2_1 _38253_ (.Y(_07665_),
    .A(_04344_),
    .B(_07643_));
 sg13g2_o21ai_1 _38254_ (.B1(net6237),
    .Y(_07666_),
    .A1(net7360),
    .A2(\u_inv.d_next[36] ));
 sg13g2_a21o_1 _38255_ (.A2(_07665_),
    .A1(net7361),
    .B1(_07666_),
    .X(_07667_));
 sg13g2_xnor2_1 _38256_ (.Y(_07668_),
    .A(_04345_),
    .B(_07639_));
 sg13g2_o21ai_1 _38257_ (.B1(_07667_),
    .Y(_07669_),
    .A1(net6238),
    .A2(_07668_));
 sg13g2_inv_1 _38258_ (.Y(_07670_),
    .A(_07669_));
 sg13g2_nand3_1 _38259_ (.B(_04343_),
    .C(_07664_),
    .A(_04342_),
    .Y(_07671_));
 sg13g2_a21oi_1 _38260_ (.A1(_04343_),
    .A2(_07664_),
    .Y(_07672_),
    .B1(_04342_));
 sg13g2_nor2_1 _38261_ (.A(net7211),
    .B(_07672_),
    .Y(_07673_));
 sg13g2_a221oi_1 _38262_ (.B2(_07673_),
    .C1(net6322),
    .B1(_07671_),
    .A1(net7213),
    .Y(_07674_),
    .A2(\u_inv.d_next[37] ));
 sg13g2_a21oi_1 _38263_ (.A1(_04345_),
    .A2(_07639_),
    .Y(_07675_),
    .B1(_04839_));
 sg13g2_xor2_1 _38264_ (.B(_07675_),
    .A(_04342_),
    .X(_07676_));
 sg13g2_a21o_2 _38265_ (.A2(_07676_),
    .A1(net6322),
    .B1(_07674_),
    .X(_07677_));
 sg13g2_a21oi_1 _38266_ (.A1(_07670_),
    .A2(_07677_),
    .Y(_07678_),
    .B1(net5858));
 sg13g2_xnor2_1 _38267_ (.Y(_07679_),
    .A(net5858),
    .B(_07670_));
 sg13g2_nand2_1 _38268_ (.Y(_07680_),
    .A(net5858),
    .B(_07677_));
 sg13g2_xnor2_1 _38269_ (.Y(_07681_),
    .A(net5858),
    .B(_07677_));
 sg13g2_or2_1 _38270_ (.X(_07682_),
    .B(_07681_),
    .A(_07679_));
 sg13g2_a21oi_1 _38271_ (.A1(_04370_),
    .A2(_07642_),
    .Y(_07683_),
    .B1(_04358_));
 sg13g2_nand3_1 _38272_ (.B(_04370_),
    .C(_07642_),
    .A(_04358_),
    .Y(_07684_));
 sg13g2_nand2b_1 _38273_ (.Y(_07685_),
    .B(_07684_),
    .A_N(_07683_));
 sg13g2_a21oi_1 _38274_ (.A1(net7361),
    .A2(_07685_),
    .Y(_07686_),
    .B1(net6322));
 sg13g2_o21ai_1 _38275_ (.B1(_07686_),
    .Y(_07687_),
    .A1(net7361),
    .A2(\u_inv.d_next[34] ));
 sg13g2_nor3_1 _38276_ (.A(_04358_),
    .B(_04831_),
    .C(_07637_),
    .Y(_07688_));
 sg13g2_o21ai_1 _38277_ (.B1(_04358_),
    .Y(_07689_),
    .A1(_04831_),
    .A2(_07637_));
 sg13g2_nand2_1 _38278_ (.Y(_07690_),
    .A(net6322),
    .B(_07689_));
 sg13g2_o21ai_1 _38279_ (.B1(_07687_),
    .Y(_07691_),
    .A1(_07688_),
    .A2(_07690_));
 sg13g2_and2_1 _38280_ (.A(net5809),
    .B(_07691_),
    .X(_07692_));
 sg13g2_xnor2_1 _38281_ (.Y(_07693_),
    .A(net5809),
    .B(_07691_));
 sg13g2_nor2b_1 _38282_ (.A(_04832_),
    .B_N(_07689_),
    .Y(_07694_));
 sg13g2_a21oi_1 _38283_ (.A1(_04357_),
    .A2(_07694_),
    .Y(_07695_),
    .B1(net6237));
 sg13g2_o21ai_1 _38284_ (.B1(_07695_),
    .Y(_07696_),
    .A1(_04357_),
    .A2(_07694_));
 sg13g2_a21oi_1 _38285_ (.A1(\u_inv.d_next[34] ),
    .A2(\u_inv.d_reg[34] ),
    .Y(_07697_),
    .B1(_07683_));
 sg13g2_xnor2_1 _38286_ (.Y(_07698_),
    .A(_04357_),
    .B(_07697_));
 sg13g2_nor2b_1 _38287_ (.A(net7361),
    .B_N(\u_inv.d_next[35] ),
    .Y(_07699_));
 sg13g2_o21ai_1 _38288_ (.B1(net6237),
    .Y(_07700_),
    .A1(net7211),
    .A2(_07698_));
 sg13g2_o21ai_1 _38289_ (.B1(_07696_),
    .Y(_07701_),
    .A1(_07699_),
    .A2(_07700_));
 sg13g2_nor2_1 _38290_ (.A(net5858),
    .B(_07701_),
    .Y(_07702_));
 sg13g2_xnor2_1 _38291_ (.Y(_07703_),
    .A(net5858),
    .B(_07701_));
 sg13g2_nor2_1 _38292_ (.A(_07693_),
    .B(_07703_),
    .Y(_07704_));
 sg13g2_nor2_1 _38293_ (.A(_04829_),
    .B(_07636_),
    .Y(_07705_));
 sg13g2_o21ai_1 _38294_ (.B1(net6323),
    .Y(_07706_),
    .A1(net6995),
    .A2(_07705_));
 sg13g2_a21oi_1 _38295_ (.A1(net6995),
    .A2(_07705_),
    .Y(_07707_),
    .B1(_07706_));
 sg13g2_and2_1 _38296_ (.A(net6995),
    .B(_04363_),
    .X(_07708_));
 sg13g2_o21ai_1 _38297_ (.B1(_07708_),
    .Y(_07709_),
    .A1(_04340_),
    .A2(_04365_));
 sg13g2_nand2_1 _38298_ (.Y(_07710_),
    .A(net7361),
    .B(_07642_));
 sg13g2_nor2_1 _38299_ (.A(_04368_),
    .B(_07710_),
    .Y(_07711_));
 sg13g2_a22oi_1 _38300_ (.Y(_07712_),
    .B1(_07709_),
    .B2(_07711_),
    .A2(\u_inv.d_next[33] ),
    .A1(net7211));
 sg13g2_a21oi_2 _38301_ (.B1(_07707_),
    .Y(_07713_),
    .A2(_07712_),
    .A1(net6238));
 sg13g2_o21ai_1 _38302_ (.B1(net7361),
    .Y(_07714_),
    .A1(_04340_),
    .A2(_04365_));
 sg13g2_a21oi_1 _38303_ (.A1(_04340_),
    .A2(_04365_),
    .Y(_07715_),
    .B1(_07714_));
 sg13g2_a21oi_1 _38304_ (.A1(net7211),
    .A2(\u_inv.d_next[32] ),
    .Y(_07716_),
    .B1(_07715_));
 sg13g2_nor2_1 _38305_ (.A(net6238),
    .B(_07636_),
    .Y(_07717_));
 sg13g2_o21ai_1 _38306_ (.B1(_07717_),
    .Y(_07718_),
    .A1(_04365_),
    .A2(_04951_));
 sg13g2_o21ai_1 _38307_ (.B1(_07718_),
    .Y(_07719_),
    .A1(net6323),
    .A2(_07716_));
 sg13g2_o21ai_1 _38308_ (.B1(_07713_),
    .Y(_07720_),
    .A1(net5809),
    .A2(_07719_));
 sg13g2_or3_1 _38309_ (.A(_07693_),
    .B(_07703_),
    .C(_07720_),
    .X(_07721_));
 sg13g2_nor2_1 _38310_ (.A(_07692_),
    .B(_07702_),
    .Y(_07722_));
 sg13g2_nand2_1 _38311_ (.Y(_07723_),
    .A(_07721_),
    .B(_07722_));
 sg13g2_inv_1 _38312_ (.Y(_07724_),
    .A(_07723_));
 sg13g2_a21oi_1 _38313_ (.A1(_07721_),
    .A2(_07722_),
    .Y(_07725_),
    .B1(_07682_));
 sg13g2_o21ai_1 _38314_ (.B1(_07663_),
    .Y(_07726_),
    .A1(_07678_),
    .A2(_07725_));
 sg13g2_nor2_1 _38315_ (.A(_07650_),
    .B(_07661_),
    .Y(_07727_));
 sg13g2_a21oi_2 _38316_ (.B1(_07635_),
    .Y(_07728_),
    .A2(_07727_),
    .A1(_07726_));
 sg13g2_a21oi_1 _38317_ (.A1(_07620_),
    .A2(_07631_),
    .Y(_07729_),
    .B1(net5859));
 sg13g2_inv_1 _38318_ (.Y(_07730_),
    .A(_07729_));
 sg13g2_nor2b_1 _38319_ (.A(_07604_),
    .B_N(_07611_),
    .Y(_07731_));
 sg13g2_o21ai_1 _38320_ (.B1(_07731_),
    .Y(_07732_),
    .A1(_07613_),
    .A2(_07730_));
 sg13g2_nand4_1 _38321_ (.B(_07572_),
    .C(_07594_),
    .A(_07561_),
    .Y(_07733_),
    .D(_07732_));
 sg13g2_nor2b_1 _38322_ (.A(_07583_),
    .B_N(_07591_),
    .Y(_07734_));
 sg13g2_nand3b_1 _38323_ (.B(_07572_),
    .C(_07561_),
    .Y(_07735_),
    .A_N(_07734_));
 sg13g2_nand4_1 _38324_ (.B(_07571_),
    .C(_07733_),
    .A(_07560_),
    .Y(_07736_),
    .D(_07735_));
 sg13g2_nor2_2 _38325_ (.A(_07728_),
    .B(_07736_),
    .Y(_07737_));
 sg13g2_o21ai_1 _38326_ (.B1(_07540_),
    .Y(_07738_),
    .A1(_07728_),
    .A2(_07736_));
 sg13g2_o21ai_1 _38327_ (.B1(net5816),
    .Y(_07739_),
    .A1(_07433_),
    .A2(_07441_));
 sg13g2_nor3_1 _38328_ (.A(_07418_),
    .B(_07426_),
    .C(_07739_),
    .Y(_07740_));
 sg13g2_a21oi_1 _38329_ (.A1(_07417_),
    .A2(_07424_),
    .Y(_07741_),
    .B1(net5865));
 sg13g2_nor2_1 _38330_ (.A(_07740_),
    .B(_07741_),
    .Y(_07742_));
 sg13g2_nor2_1 _38331_ (.A(_07407_),
    .B(_07742_),
    .Y(_07743_));
 sg13g2_o21ai_1 _38332_ (.B1(net5817),
    .Y(_07744_),
    .A1(_07395_),
    .A2(_07402_));
 sg13g2_nor3_1 _38333_ (.A(_07379_),
    .B(_07389_),
    .C(_07744_),
    .Y(_07745_));
 sg13g2_nand2_1 _38334_ (.Y(_07746_),
    .A(_07378_),
    .B(_07388_));
 sg13g2_nor3_1 _38335_ (.A(_07743_),
    .B(_07745_),
    .C(_07746_),
    .Y(_07747_));
 sg13g2_a21oi_1 _38336_ (.A1(_07526_),
    .A2(_07533_),
    .Y(_07748_),
    .B1(net5861));
 sg13g2_or2_1 _38337_ (.X(_07749_),
    .B(_07514_),
    .A(_07503_));
 sg13g2_a21o_1 _38338_ (.A2(_07748_),
    .A1(_07516_),
    .B1(_07749_),
    .X(_07750_));
 sg13g2_nand4_1 _38339_ (.B(_07489_),
    .C(_07496_),
    .A(_07477_),
    .Y(_07751_),
    .D(_07750_));
 sg13g2_o21ai_1 _38340_ (.B1(net5815),
    .Y(_07752_),
    .A1(_07487_),
    .A2(_07494_));
 sg13g2_nand2b_1 _38341_ (.Y(_07753_),
    .B(_07477_),
    .A_N(_07752_));
 sg13g2_nor2_1 _38342_ (.A(_07462_),
    .B(_07475_),
    .Y(_07754_));
 sg13g2_nand3_1 _38343_ (.B(_07753_),
    .C(_07754_),
    .A(_07751_),
    .Y(_07755_));
 sg13g2_nand2_1 _38344_ (.Y(_07756_),
    .A(_07446_),
    .B(_07755_));
 sg13g2_and3_2 _38345_ (.X(_07757_),
    .A(_07738_),
    .B(_07747_),
    .C(_07756_));
 sg13g2_nand3_1 _38346_ (.B(_07747_),
    .C(_07756_),
    .A(_07738_),
    .Y(_07758_));
 sg13g2_nor2b_2 _38347_ (.A(_04325_),
    .B_N(_04335_),
    .Y(_07759_));
 sg13g2_nor2_1 _38348_ (.A(_04218_),
    .B(_07759_),
    .Y(_07760_));
 sg13g2_nand2b_1 _38349_ (.Y(_07761_),
    .B(_04219_),
    .A_N(_07759_));
 sg13g2_o21ai_1 _38350_ (.B1(_04233_),
    .Y(_07762_),
    .A1(_04220_),
    .A2(_07759_));
 sg13g2_a21oi_1 _38351_ (.A1(_04205_),
    .A2(_07762_),
    .Y(_07763_),
    .B1(_04223_));
 sg13g2_nor2_1 _38352_ (.A(_04208_),
    .B(_07763_),
    .Y(_07764_));
 sg13g2_xnor2_1 _38353_ (.Y(_07765_),
    .A(_04208_),
    .B(_07763_));
 sg13g2_o21ai_1 _38354_ (.B1(net6233),
    .Y(_07766_),
    .A1(net7355),
    .A2(\u_inv.d_next[30] ));
 sg13g2_a21oi_1 _38355_ (.A1(net7356),
    .A2(_07765_),
    .Y(_07767_),
    .B1(_07766_));
 sg13g2_nand2_1 _38356_ (.Y(_07768_),
    .A(_04930_),
    .B(_04944_));
 sg13g2_a21oi_1 _38357_ (.A1(_04930_),
    .A2(_04944_),
    .Y(_07769_),
    .B1(_04868_));
 sg13g2_o21ai_1 _38358_ (.B1(_04214_),
    .Y(_07770_),
    .A1(_04878_),
    .A2(_07769_));
 sg13g2_a22oi_1 _38359_ (.Y(_07771_),
    .B1(_04880_),
    .B2(_07770_),
    .A2(\u_inv.d_reg[27] ),
    .A1(_18177_));
 sg13g2_a221oi_1 _38360_ (.B2(_07770_),
    .C1(_04864_),
    .B1(_04880_),
    .A1(_18177_),
    .Y(_07772_),
    .A2(\u_inv.d_reg[27] ));
 sg13g2_nor3_1 _38361_ (.A(_04208_),
    .B(_04872_),
    .C(_07772_),
    .Y(_07773_));
 sg13g2_o21ai_1 _38362_ (.B1(_04208_),
    .Y(_07774_),
    .A1(_04872_),
    .A2(_07772_));
 sg13g2_nor2b_1 _38363_ (.A(_07773_),
    .B_N(_07774_),
    .Y(_07775_));
 sg13g2_a21oi_2 _38364_ (.B1(_07767_),
    .Y(_07776_),
    .A2(_07775_),
    .A1(net6318));
 sg13g2_nor2_1 _38365_ (.A(net5853),
    .B(_07776_),
    .Y(_07777_));
 sg13g2_nand2_1 _38366_ (.Y(_07778_),
    .A(net5853),
    .B(_07776_));
 sg13g2_nand2b_1 _38367_ (.Y(_07779_),
    .B(_07778_),
    .A_N(_07777_));
 sg13g2_a21o_1 _38368_ (.A2(_07774_),
    .A1(_04873_),
    .B1(_04206_),
    .X(_07780_));
 sg13g2_nand3_1 _38369_ (.B(_04873_),
    .C(_07774_),
    .A(_04206_),
    .Y(_07781_));
 sg13g2_nand3_1 _38370_ (.B(_07780_),
    .C(_07781_),
    .A(net6318),
    .Y(_07782_));
 sg13g2_a21oi_1 _38371_ (.A1(\u_inv.d_next[30] ),
    .A2(\u_inv.d_reg[30] ),
    .Y(_07783_),
    .B1(_07764_));
 sg13g2_o21ai_1 _38372_ (.B1(net7355),
    .Y(_07784_),
    .A1(_04206_),
    .A2(_07783_));
 sg13g2_a21oi_1 _38373_ (.A1(_04206_),
    .A2(_07783_),
    .Y(_07785_),
    .B1(_07784_));
 sg13g2_o21ai_1 _38374_ (.B1(net6233),
    .Y(_07786_),
    .A1(net7355),
    .A2(_18174_));
 sg13g2_o21ai_1 _38375_ (.B1(_07782_),
    .Y(_07787_),
    .A1(_07785_),
    .A2(_07786_));
 sg13g2_xnor2_1 _38376_ (.Y(_07788_),
    .A(net5803),
    .B(_07787_));
 sg13g2_nand2b_1 _38377_ (.Y(_07789_),
    .B(_07788_),
    .A_N(_07779_));
 sg13g2_xnor2_1 _38378_ (.Y(_07790_),
    .A(_04218_),
    .B(_07759_));
 sg13g2_a21oi_1 _38379_ (.A1(net7344),
    .A2(_07790_),
    .Y(_07791_),
    .B1(net6308));
 sg13g2_o21ai_1 _38380_ (.B1(_07791_),
    .Y(_07792_),
    .A1(net7344),
    .A2(\u_inv.d_next[24] ));
 sg13g2_xnor2_1 _38381_ (.Y(_07793_),
    .A(_04218_),
    .B(_07768_));
 sg13g2_o21ai_1 _38382_ (.B1(_07792_),
    .Y(_07794_),
    .A1(net6225),
    .A2(_07793_));
 sg13g2_and2_1 _38383_ (.A(net5802),
    .B(_07794_),
    .X(_07795_));
 sg13g2_a21oi_1 _38384_ (.A1(\u_inv.d_next[24] ),
    .A2(\u_inv.d_reg[24] ),
    .Y(_07796_),
    .B1(_07760_));
 sg13g2_o21ai_1 _38385_ (.B1(net7344),
    .Y(_07797_),
    .A1(_04217_),
    .A2(_07796_));
 sg13g2_a21oi_1 _38386_ (.A1(_04217_),
    .A2(_07796_),
    .Y(_07798_),
    .B1(_07797_));
 sg13g2_a21oi_1 _38387_ (.A1(net7203),
    .A2(\u_inv.d_next[25] ),
    .Y(_07799_),
    .B1(net6308));
 sg13g2_nand2b_1 _38388_ (.Y(_07800_),
    .B(_07799_),
    .A_N(_07798_));
 sg13g2_a21oi_1 _38389_ (.A1(_04218_),
    .A2(_07768_),
    .Y(_07801_),
    .B1(_04876_));
 sg13g2_xnor2_1 _38390_ (.Y(_07802_),
    .A(_04217_),
    .B(_07801_));
 sg13g2_o21ai_1 _38391_ (.B1(_07800_),
    .Y(_07803_),
    .A1(net6226),
    .A2(_07802_));
 sg13g2_nor2_1 _38392_ (.A(net5854),
    .B(_07803_),
    .Y(_07804_));
 sg13g2_or2_1 _38393_ (.X(_07805_),
    .B(_07804_),
    .A(_07795_));
 sg13g2_inv_1 _38394_ (.Y(_07806_),
    .A(_07805_));
 sg13g2_xnor2_1 _38395_ (.Y(_07807_),
    .A(_04204_),
    .B(_07771_));
 sg13g2_nand2b_1 _38396_ (.Y(_07808_),
    .B(_07762_),
    .A_N(_04204_));
 sg13g2_nand2b_1 _38397_ (.Y(_07809_),
    .B(_04204_),
    .A_N(_07762_));
 sg13g2_nand3_1 _38398_ (.B(_07808_),
    .C(_07809_),
    .A(net7355),
    .Y(_07810_));
 sg13g2_a21oi_1 _38399_ (.A1(net7213),
    .A2(\u_inv.d_next[28] ),
    .Y(_07811_),
    .B1(net6319));
 sg13g2_a22oi_1 _38400_ (.Y(_07812_),
    .B1(_07810_),
    .B2(_07811_),
    .A2(_07807_),
    .A1(net6319));
 sg13g2_nand2_1 _38401_ (.Y(_07813_),
    .A(net5802),
    .B(_07812_));
 sg13g2_xnor2_1 _38402_ (.Y(_07814_),
    .A(net5802),
    .B(_07812_));
 sg13g2_inv_1 _38403_ (.Y(_07815_),
    .A(_07814_));
 sg13g2_a21oi_1 _38404_ (.A1(_04204_),
    .A2(_07771_),
    .Y(_07816_),
    .B1(_04870_));
 sg13g2_and2_1 _38405_ (.A(_04203_),
    .B(_07816_),
    .X(_07817_));
 sg13g2_o21ai_1 _38406_ (.B1(net6319),
    .Y(_07818_),
    .A1(_04203_),
    .A2(_07816_));
 sg13g2_o21ai_1 _38407_ (.B1(_07808_),
    .Y(_07819_),
    .A1(_18176_),
    .A2(_18586_));
 sg13g2_xnor2_1 _38408_ (.Y(_07820_),
    .A(_04203_),
    .B(_07819_));
 sg13g2_a21oi_1 _38409_ (.A1(net7355),
    .A2(_07820_),
    .Y(_07821_),
    .B1(net6319));
 sg13g2_o21ai_1 _38410_ (.B1(_07821_),
    .Y(_07822_),
    .A1(net7355),
    .A2(_18175_));
 sg13g2_o21ai_1 _38411_ (.B1(_07822_),
    .Y(_07823_),
    .A1(_07817_),
    .A2(_07818_));
 sg13g2_nor2_1 _38412_ (.A(net5853),
    .B(_07823_),
    .Y(_07824_));
 sg13g2_xnor2_1 _38413_ (.Y(_07825_),
    .A(net5853),
    .B(_07823_));
 sg13g2_nor2_1 _38414_ (.A(_07814_),
    .B(_07825_),
    .Y(_07826_));
 sg13g2_a21o_1 _38415_ (.A2(_07761_),
    .A1(_04229_),
    .B1(_04214_),
    .X(_07827_));
 sg13g2_a21oi_1 _38416_ (.A1(_04213_),
    .A2(_07827_),
    .Y(_07828_),
    .B1(_04212_));
 sg13g2_nand3_1 _38417_ (.B(_04213_),
    .C(_07827_),
    .A(_04212_),
    .Y(_07829_));
 sg13g2_nand2_1 _38418_ (.Y(_07830_),
    .A(net7355),
    .B(_07829_));
 sg13g2_a21oi_1 _38419_ (.A1(net7213),
    .A2(\u_inv.d_next[27] ),
    .Y(_07831_),
    .B1(net6319));
 sg13g2_o21ai_1 _38420_ (.B1(_07831_),
    .Y(_07832_),
    .A1(_07828_),
    .A2(_07830_));
 sg13g2_nand2_1 _38421_ (.Y(_07833_),
    .A(_04879_),
    .B(_07770_));
 sg13g2_xor2_1 _38422_ (.B(_07833_),
    .A(_04212_),
    .X(_07834_));
 sg13g2_o21ai_1 _38423_ (.B1(_07832_),
    .Y(_07835_),
    .A1(net6233),
    .A2(_07834_));
 sg13g2_xnor2_1 _38424_ (.Y(_07836_),
    .A(net5853),
    .B(_07835_));
 sg13g2_nand3_1 _38425_ (.B(_04229_),
    .C(_07761_),
    .A(_04214_),
    .Y(_07837_));
 sg13g2_a21oi_1 _38426_ (.A1(_07827_),
    .A2(_07837_),
    .Y(_07838_),
    .B1(net7213));
 sg13g2_o21ai_1 _38427_ (.B1(net6233),
    .Y(_07839_),
    .A1(net7355),
    .A2(\u_inv.d_next[26] ));
 sg13g2_nor2_1 _38428_ (.A(_07838_),
    .B(_07839_),
    .Y(_07840_));
 sg13g2_nor3_1 _38429_ (.A(_04214_),
    .B(_04878_),
    .C(_07769_),
    .Y(_07841_));
 sg13g2_nand3b_1 _38430_ (.B(net6308),
    .C(_07770_),
    .Y(_07842_),
    .A_N(_07841_));
 sg13g2_nor2b_2 _38431_ (.A(_07840_),
    .B_N(_07842_),
    .Y(_07843_));
 sg13g2_nor2_1 _38432_ (.A(net5854),
    .B(_07843_),
    .Y(_07844_));
 sg13g2_xnor2_1 _38433_ (.Y(_07845_),
    .A(net5802),
    .B(_07843_));
 sg13g2_xnor2_1 _38434_ (.Y(_07846_),
    .A(net5854),
    .B(_07843_));
 sg13g2_nor2_1 _38435_ (.A(_07836_),
    .B(_07846_),
    .Y(_07847_));
 sg13g2_inv_1 _38436_ (.Y(_07848_),
    .A(_07847_));
 sg13g2_nor4_1 _38437_ (.A(_07814_),
    .B(_07825_),
    .C(_07836_),
    .D(_07846_),
    .Y(_07849_));
 sg13g2_a21oi_1 _38438_ (.A1(net5803),
    .A2(_07812_),
    .Y(_07850_),
    .B1(_07824_));
 sg13g2_o21ai_1 _38439_ (.B1(_07813_),
    .Y(_07851_),
    .A1(net5853),
    .A2(_07823_));
 sg13g2_a21oi_1 _38440_ (.A1(_07835_),
    .A2(_07843_),
    .Y(_07852_),
    .B1(net5853));
 sg13g2_a221oi_1 _38441_ (.B2(_07826_),
    .C1(_07851_),
    .B1(_07852_),
    .A1(_07805_),
    .Y(_07853_),
    .A2(_07849_));
 sg13g2_a21o_1 _38442_ (.A2(_07787_),
    .A1(_07776_),
    .B1(net5853),
    .X(_07854_));
 sg13g2_o21ai_1 _38443_ (.B1(_07854_),
    .Y(_07855_),
    .A1(_07789_),
    .A2(_07853_));
 sg13g2_xnor2_1 _38444_ (.Y(_07856_),
    .A(net5803),
    .B(_07803_));
 sg13g2_xnor2_1 _38445_ (.Y(_07857_),
    .A(net5854),
    .B(_07794_));
 sg13g2_nand3_1 _38446_ (.B(_07856_),
    .C(_07857_),
    .A(_07849_),
    .Y(_07858_));
 sg13g2_or2_1 _38447_ (.X(_07859_),
    .B(_07858_),
    .A(_07789_));
 sg13g2_nand2b_2 _38448_ (.Y(_07860_),
    .B(_07859_),
    .A_N(_07855_));
 sg13g2_o21ai_1 _38449_ (.B1(_04928_),
    .Y(_07861_),
    .A1(_04918_),
    .A2(_04921_));
 sg13g2_nand2_1 _38450_ (.Y(_07862_),
    .A(_04932_),
    .B(_07861_));
 sg13g2_a21oi_1 _38451_ (.A1(_04932_),
    .A2(_07861_),
    .Y(_07863_),
    .B1(_04927_));
 sg13g2_o21ai_1 _38452_ (.B1(_04299_),
    .Y(_07864_),
    .A1(_04934_),
    .A2(_07863_));
 sg13g2_a21oi_1 _38453_ (.A1(_04937_),
    .A2(_07864_),
    .Y(_07865_),
    .B1(_04301_));
 sg13g2_nor2_1 _38454_ (.A(_04939_),
    .B(_07865_),
    .Y(_07866_));
 sg13g2_o21ai_1 _38455_ (.B1(_04309_),
    .Y(_07867_),
    .A1(_04939_),
    .A2(_07865_));
 sg13g2_nand3_1 _38456_ (.B(_04935_),
    .C(_07867_),
    .A(_04305_),
    .Y(_07868_));
 sg13g2_a21oi_1 _38457_ (.A1(_04935_),
    .A2(_07867_),
    .Y(_07869_),
    .B1(_04305_));
 sg13g2_nor2_1 _38458_ (.A(net6225),
    .B(_07869_),
    .Y(_07870_));
 sg13g2_nand2_1 _38459_ (.Y(_07871_),
    .A(_04297_),
    .B(_04321_));
 sg13g2_nor2_2 _38460_ (.A(_04314_),
    .B(_07871_),
    .Y(_07872_));
 sg13g2_a21oi_2 _38461_ (.B1(_04330_),
    .Y(_07873_),
    .A2(_07872_),
    .A1(_04323_));
 sg13g2_o21ai_1 _38462_ (.B1(_04332_),
    .Y(_07874_),
    .A1(_04302_),
    .A2(_07873_));
 sg13g2_nand2_1 _38463_ (.Y(_07875_),
    .A(_04308_),
    .B(_07874_));
 sg13g2_nand3_1 _38464_ (.B(_04307_),
    .C(_07875_),
    .A(_04305_),
    .Y(_07876_));
 sg13g2_a21oi_1 _38465_ (.A1(_04307_),
    .A2(_07875_),
    .Y(_07877_),
    .B1(_04305_));
 sg13g2_nor2_1 _38466_ (.A(net7203),
    .B(_07877_),
    .Y(_07878_));
 sg13g2_a221oi_1 _38467_ (.B2(_07878_),
    .C1(net6309),
    .B1(_07876_),
    .A1(net7203),
    .Y(_07879_),
    .A2(\u_inv.d_next[23] ));
 sg13g2_a21o_2 _38468_ (.A2(_07870_),
    .A1(_07868_),
    .B1(_07879_),
    .X(_07880_));
 sg13g2_xnor2_1 _38469_ (.Y(_07881_),
    .A(net5802),
    .B(_07880_));
 sg13g2_xnor2_1 _38470_ (.Y(_07882_),
    .A(_04308_),
    .B(_07866_));
 sg13g2_nand2b_1 _38471_ (.Y(_07883_),
    .B(_04309_),
    .A_N(_07874_));
 sg13g2_nand3_1 _38472_ (.B(_07875_),
    .C(_07883_),
    .A(net7343),
    .Y(_07884_));
 sg13g2_a21oi_1 _38473_ (.A1(net7203),
    .A2(\u_inv.d_next[22] ),
    .Y(_07885_),
    .B1(net6309));
 sg13g2_a22oi_1 _38474_ (.Y(_07886_),
    .B1(_07884_),
    .B2(_07885_),
    .A2(_07882_),
    .A1(net6309));
 sg13g2_nand2_1 _38475_ (.Y(_07887_),
    .A(net5802),
    .B(_07886_));
 sg13g2_xnor2_1 _38476_ (.Y(_07888_),
    .A(net5854),
    .B(_07886_));
 sg13g2_nand2_1 _38477_ (.Y(_07889_),
    .A(_07881_),
    .B(_07888_));
 sg13g2_xnor2_1 _38478_ (.Y(_07890_),
    .A(_04299_),
    .B(_07873_));
 sg13g2_nor2_1 _38479_ (.A(net7344),
    .B(\u_inv.d_next[20] ),
    .Y(_07891_));
 sg13g2_a21oi_1 _38480_ (.A1(net7345),
    .A2(_07890_),
    .Y(_07892_),
    .B1(_07891_));
 sg13g2_nor3_1 _38481_ (.A(_04299_),
    .B(_04934_),
    .C(_07863_),
    .Y(_07893_));
 sg13g2_nor2_1 _38482_ (.A(net6226),
    .B(_07893_),
    .Y(_07894_));
 sg13g2_a22oi_1 _38483_ (.Y(_07895_),
    .B1(_07894_),
    .B2(_07864_),
    .A2(_07892_),
    .A1(net6226));
 sg13g2_nor2_1 _38484_ (.A(net5848),
    .B(_07895_),
    .Y(_07896_));
 sg13g2_o21ai_1 _38485_ (.B1(_04298_),
    .Y(_07897_),
    .A1(_04299_),
    .A2(_07873_));
 sg13g2_o21ai_1 _38486_ (.B1(net7345),
    .Y(_07898_),
    .A1(_04301_),
    .A2(_07897_));
 sg13g2_a21oi_1 _38487_ (.A1(_04301_),
    .A2(_07897_),
    .Y(_07899_),
    .B1(_07898_));
 sg13g2_a21oi_1 _38488_ (.A1(net7204),
    .A2(\u_inv.d_next[21] ),
    .Y(_07900_),
    .B1(_07899_));
 sg13g2_nand3_1 _38489_ (.B(_04937_),
    .C(_07864_),
    .A(_04301_),
    .Y(_07901_));
 sg13g2_nand3b_1 _38490_ (.B(_07901_),
    .C(net6310),
    .Y(_07902_),
    .A_N(_07865_));
 sg13g2_o21ai_1 _38491_ (.B1(_07902_),
    .Y(_07903_),
    .A1(net6310),
    .A2(_07900_));
 sg13g2_a21oi_1 _38492_ (.A1(net5802),
    .A2(_07903_),
    .Y(_07904_),
    .B1(_07896_));
 sg13g2_xnor2_1 _38493_ (.Y(_07905_),
    .A(net5794),
    .B(_07895_));
 sg13g2_or2_1 _38494_ (.X(_07906_),
    .B(_07903_),
    .A(net5802));
 sg13g2_xnor2_1 _38495_ (.Y(_07907_),
    .A(net5848),
    .B(_07903_));
 sg13g2_and2_1 _38496_ (.A(_07905_),
    .B(_07907_),
    .X(_07908_));
 sg13g2_nor3_1 _38497_ (.A(_04319_),
    .B(_04328_),
    .C(_07872_),
    .Y(_07909_));
 sg13g2_o21ai_1 _38498_ (.B1(_04319_),
    .Y(_07910_),
    .A1(_04328_),
    .A2(_07872_));
 sg13g2_nand2b_1 _38499_ (.Y(_07911_),
    .B(_07910_),
    .A_N(_07909_));
 sg13g2_o21ai_1 _38500_ (.B1(net6226),
    .Y(_07912_),
    .A1(net7344),
    .A2(net7299));
 sg13g2_a21o_1 _38501_ (.A2(_07911_),
    .A1(net7344),
    .B1(_07912_),
    .X(_07913_));
 sg13g2_a21oi_1 _38502_ (.A1(_04932_),
    .A2(_07861_),
    .Y(_07914_),
    .B1(_04319_));
 sg13g2_o21ai_1 _38503_ (.B1(net6308),
    .Y(_07915_),
    .A1(_04318_),
    .A2(_07862_));
 sg13g2_o21ai_1 _38504_ (.B1(_07913_),
    .Y(_07916_),
    .A1(_07914_),
    .A2(_07915_));
 sg13g2_nand2_1 _38505_ (.Y(_07917_),
    .A(net5794),
    .B(_07916_));
 sg13g2_xnor2_1 _38506_ (.Y(_07918_),
    .A(net5794),
    .B(_07916_));
 sg13g2_a21oi_1 _38507_ (.A1(net7299),
    .A2(_18596_),
    .Y(_07919_),
    .B1(_07914_));
 sg13g2_o21ai_1 _38508_ (.B1(net6308),
    .Y(_07920_),
    .A1(_04311_),
    .A2(_07919_));
 sg13g2_a21oi_1 _38509_ (.A1(_04311_),
    .A2(_07919_),
    .Y(_07921_),
    .B1(_07920_));
 sg13g2_a21oi_1 _38510_ (.A1(_04316_),
    .A2(_07910_),
    .Y(_07922_),
    .B1(_04311_));
 sg13g2_nand3_1 _38511_ (.B(_04316_),
    .C(_07910_),
    .A(_04311_),
    .Y(_07923_));
 sg13g2_nor2_1 _38512_ (.A(net7203),
    .B(_07922_),
    .Y(_07924_));
 sg13g2_a221oi_1 _38513_ (.B2(_07924_),
    .C1(net6308),
    .B1(_07923_),
    .A1(net7203),
    .Y(_07925_),
    .A2(\u_inv.d_next[19] ));
 sg13g2_or2_1 _38514_ (.X(_07926_),
    .B(_07925_),
    .A(_07921_));
 sg13g2_xnor2_1 _38515_ (.Y(_07927_),
    .A(net5848),
    .B(_07926_));
 sg13g2_nor2_1 _38516_ (.A(_04321_),
    .B(_04923_),
    .Y(_07928_));
 sg13g2_or2_1 _38517_ (.X(_07929_),
    .B(_07928_),
    .A(_04931_));
 sg13g2_o21ai_1 _38518_ (.B1(net6308),
    .Y(_07930_),
    .A1(_04315_),
    .A2(_07929_));
 sg13g2_a21oi_1 _38519_ (.A1(_04315_),
    .A2(_07929_),
    .Y(_07931_),
    .B1(_07930_));
 sg13g2_nand3b_1 _38520_ (.B(_07871_),
    .C(_04314_),
    .Y(_07932_),
    .A_N(_04320_));
 sg13g2_a21oi_1 _38521_ (.A1(_04315_),
    .A2(_04320_),
    .Y(_07933_),
    .B1(net7203));
 sg13g2_nand3b_1 _38522_ (.B(_07932_),
    .C(_07933_),
    .Y(_07934_),
    .A_N(_07872_));
 sg13g2_a21oi_1 _38523_ (.A1(net7209),
    .A2(\u_inv.d_next[17] ),
    .Y(_07935_),
    .B1(net6308));
 sg13g2_a21oi_2 _38524_ (.B1(_07931_),
    .Y(_07936_),
    .A2(_07935_),
    .A1(_07934_));
 sg13g2_nand2_1 _38525_ (.Y(_07937_),
    .A(_04321_),
    .B(_04923_));
 sg13g2_nor2_1 _38526_ (.A(net6226),
    .B(_07928_),
    .Y(_07938_));
 sg13g2_xnor2_1 _38527_ (.Y(_07939_),
    .A(_04297_),
    .B(_04321_));
 sg13g2_nor2_1 _38528_ (.A(net7344),
    .B(\u_inv.d_next[16] ),
    .Y(_07940_));
 sg13g2_a21oi_1 _38529_ (.A1(net7344),
    .A2(_07939_),
    .Y(_07941_),
    .B1(_07940_));
 sg13g2_a22oi_1 _38530_ (.Y(_07942_),
    .B1(_07941_),
    .B2(net6226),
    .A2(_07938_),
    .A1(_07937_));
 sg13g2_inv_1 _38531_ (.Y(_07943_),
    .A(_07942_));
 sg13g2_o21ai_1 _38532_ (.B1(net5794),
    .Y(_07944_),
    .A1(_07936_),
    .A2(_07943_));
 sg13g2_nor3_1 _38533_ (.A(_07918_),
    .B(_07927_),
    .C(_07944_),
    .Y(_07945_));
 sg13g2_o21ai_1 _38534_ (.B1(_07917_),
    .Y(_07946_),
    .A1(net5848),
    .A2(_07926_));
 sg13g2_or2_1 _38535_ (.X(_07947_),
    .B(_07946_),
    .A(_07945_));
 sg13g2_o21ai_1 _38536_ (.B1(_07908_),
    .Y(_07948_),
    .A1(_07945_),
    .A2(_07946_));
 sg13g2_a21oi_1 _38537_ (.A1(_07904_),
    .A2(_07948_),
    .Y(_07949_),
    .B1(_07889_));
 sg13g2_o21ai_1 _38538_ (.B1(_07887_),
    .Y(_07950_),
    .A1(net5854),
    .A2(_07880_));
 sg13g2_nor2_1 _38539_ (.A(_07949_),
    .B(_07950_),
    .Y(_07951_));
 sg13g2_nor3_1 _38540_ (.A(_07855_),
    .B(_07949_),
    .C(_07950_),
    .Y(_07952_));
 sg13g2_nand3_1 _38541_ (.B(_04907_),
    .C(_04908_),
    .A(_04281_),
    .Y(_07953_));
 sg13g2_nor2_1 _38542_ (.A(_04277_),
    .B(_04286_),
    .Y(_07954_));
 sg13g2_nor2b_1 _38543_ (.A(_07954_),
    .B_N(_04281_),
    .Y(_07955_));
 sg13g2_and2_1 _38544_ (.A(net6298),
    .B(_04909_),
    .X(_07956_));
 sg13g2_xor2_1 _38545_ (.B(_07954_),
    .A(_04281_),
    .X(_07957_));
 sg13g2_o21ai_1 _38546_ (.B1(net6218),
    .Y(_07958_),
    .A1(net7331),
    .A2(\u_inv.d_next[6] ));
 sg13g2_a21oi_1 _38547_ (.A1(net7331),
    .A2(_07957_),
    .Y(_07959_),
    .B1(_07958_));
 sg13g2_a21o_2 _38548_ (.A2(_07956_),
    .A1(_07953_),
    .B1(_07959_),
    .X(_07960_));
 sg13g2_xnor2_1 _38549_ (.Y(_07961_),
    .A(net5795),
    .B(_07960_));
 sg13g2_nor2_1 _38550_ (.A(_04280_),
    .B(_07955_),
    .Y(_07962_));
 sg13g2_o21ai_1 _38551_ (.B1(net7330),
    .Y(_07963_),
    .A1(_04279_),
    .A2(_07962_));
 sg13g2_a21oi_1 _38552_ (.A1(_04279_),
    .A2(_07962_),
    .Y(_07964_),
    .B1(_07963_));
 sg13g2_a21oi_1 _38553_ (.A1(net7196),
    .A2(\u_inv.d_next[7] ),
    .Y(_07965_),
    .B1(net6299));
 sg13g2_nand2b_1 _38554_ (.Y(_07966_),
    .B(_07965_),
    .A_N(_07964_));
 sg13g2_nor2b_1 _38555_ (.A(_04897_),
    .B_N(_04909_),
    .Y(_07967_));
 sg13g2_xnor2_1 _38556_ (.Y(_07968_),
    .A(_04279_),
    .B(_07967_));
 sg13g2_o21ai_1 _38557_ (.B1(_07966_),
    .Y(_07969_),
    .A1(net6218),
    .A2(_07968_));
 sg13g2_nor2_1 _38558_ (.A(net5795),
    .B(_07969_),
    .Y(_07970_));
 sg13g2_xnor2_1 _38559_ (.Y(_07971_),
    .A(net5846),
    .B(_07969_));
 sg13g2_and2_1 _38560_ (.A(_07961_),
    .B(_07971_),
    .X(_07972_));
 sg13g2_nand3_1 _38561_ (.B(_04273_),
    .C(_04276_),
    .A(_04269_),
    .Y(_07973_));
 sg13g2_o21ai_1 _38562_ (.B1(net7331),
    .Y(_07974_),
    .A1(_04269_),
    .A2(_04273_));
 sg13g2_nor2_1 _38563_ (.A(_04277_),
    .B(_07974_),
    .Y(_07975_));
 sg13g2_o21ai_1 _38564_ (.B1(net6299),
    .Y(_07976_),
    .A1(_04269_),
    .A2(_04906_));
 sg13g2_a21oi_1 _38565_ (.A1(_04269_),
    .A2(_04906_),
    .Y(_07977_),
    .B1(_07976_));
 sg13g2_a221oi_1 _38566_ (.B2(_07975_),
    .C1(net6299),
    .B1(_07973_),
    .A1(net7196),
    .Y(_07978_),
    .A2(\u_inv.d_next[5] ));
 sg13g2_nor2_2 _38567_ (.A(_07977_),
    .B(_07978_),
    .Y(_07979_));
 sg13g2_xnor2_1 _38568_ (.Y(_07980_),
    .A(net5793),
    .B(_07979_));
 sg13g2_xnor2_1 _38569_ (.Y(_07981_),
    .A(_04271_),
    .B(_04901_));
 sg13g2_o21ai_1 _38570_ (.B1(net6218),
    .Y(_07982_),
    .A1(net7330),
    .A2(\u_inv.d_next[3] ));
 sg13g2_a21oi_1 _38571_ (.A1(net7330),
    .A2(_07981_),
    .Y(_07983_),
    .B1(_07982_));
 sg13g2_xnor2_1 _38572_ (.Y(_07984_),
    .A(_04901_),
    .B(_04903_));
 sg13g2_or2_1 _38573_ (.X(_07985_),
    .B(_07984_),
    .A(net6218));
 sg13g2_nor2b_2 _38574_ (.A(_07983_),
    .B_N(_07985_),
    .Y(_07986_));
 sg13g2_inv_1 _38575_ (.Y(_07987_),
    .A(_07986_));
 sg13g2_nor2_1 _38576_ (.A(net5845),
    .B(_07986_),
    .Y(_07988_));
 sg13g2_nand2_1 _38577_ (.Y(_07989_),
    .A(net5793),
    .B(_07987_));
 sg13g2_a221oi_1 _38578_ (.B2(_05341_),
    .C1(_07987_),
    .B1(_05340_),
    .A1(_04590_),
    .Y(_07990_),
    .A2(_04592_));
 sg13g2_nand3_1 _38579_ (.B(net6757),
    .C(_05349_),
    .A(_03351_),
    .Y(_07991_));
 sg13g2_inv_1 _38580_ (.Y(_07992_),
    .A(_07991_));
 sg13g2_nor2_1 _38581_ (.A(_03351_),
    .B(_05349_),
    .Y(_07993_));
 sg13g2_a221oi_1 _38582_ (.B2(net6801),
    .C1(_04593_),
    .B1(_07993_),
    .A1(_05340_),
    .Y(_07994_),
    .A2(_05341_));
 sg13g2_or2_1 _38583_ (.X(_07995_),
    .B(_07994_),
    .A(_07992_));
 sg13g2_or3_1 _38584_ (.A(_07990_),
    .B(_07992_),
    .C(_07994_),
    .X(_07996_));
 sg13g2_and2_1 _38585_ (.A(_07989_),
    .B(_07996_),
    .X(_07997_));
 sg13g2_xnor2_1 _38586_ (.Y(_07998_),
    .A(_04275_),
    .B(_04904_));
 sg13g2_o21ai_1 _38587_ (.B1(_04275_),
    .Y(_07999_),
    .A1(_04270_),
    .A2(_04272_));
 sg13g2_nand3_1 _38588_ (.B(_04276_),
    .C(_07999_),
    .A(net7331),
    .Y(_08000_));
 sg13g2_nand2_1 _38589_ (.Y(_08001_),
    .A(net7197),
    .B(\u_inv.d_next[4] ));
 sg13g2_a21oi_1 _38590_ (.A1(_08000_),
    .A2(_08001_),
    .Y(_08002_),
    .B1(net6299));
 sg13g2_a21oi_2 _38591_ (.B1(_08002_),
    .Y(_08003_),
    .A2(_07998_),
    .A1(net6299));
 sg13g2_nand2_1 _38592_ (.Y(_08004_),
    .A(net5845),
    .B(_08003_));
 sg13g2_nand2b_1 _38593_ (.Y(_08005_),
    .B(net5793),
    .A_N(_08003_));
 sg13g2_nor2_1 _38594_ (.A(net5793),
    .B(_08003_),
    .Y(_08006_));
 sg13g2_nand2_1 _38595_ (.Y(_08007_),
    .A(_08004_),
    .B(_08005_));
 sg13g2_nor2b_1 _38596_ (.A(_07997_),
    .B_N(_08007_),
    .Y(_08008_));
 sg13g2_a221oi_1 _38597_ (.B2(_08005_),
    .C1(_07980_),
    .B1(_08004_),
    .A1(_07989_),
    .Y(_08009_),
    .A2(_07996_));
 sg13g2_and2_1 _38598_ (.A(_07979_),
    .B(_08004_),
    .X(_08010_));
 sg13g2_nor2_1 _38599_ (.A(_08009_),
    .B(_08010_),
    .Y(_08011_));
 sg13g2_o21ai_1 _38600_ (.B1(_07972_),
    .Y(_08012_),
    .A1(_08009_),
    .A2(_08010_));
 sg13g2_a21oi_1 _38601_ (.A1(net5846),
    .A2(_07960_),
    .Y(_08013_),
    .B1(_07970_));
 sg13g2_nand2_1 _38602_ (.Y(_08014_),
    .A(_08012_),
    .B(_08013_));
 sg13g2_a21oi_1 _38603_ (.A1(_04912_),
    .A2(_04913_),
    .Y(_08015_),
    .B1(_04916_));
 sg13g2_nor2_1 _38604_ (.A(_04259_),
    .B(_08015_),
    .Y(_08016_));
 sg13g2_xnor2_1 _38605_ (.Y(_08017_),
    .A(_04260_),
    .B(_08015_));
 sg13g2_nor2_1 _38606_ (.A(_04258_),
    .B(_04292_),
    .Y(_08018_));
 sg13g2_nor2_1 _38607_ (.A(_04260_),
    .B(_08018_),
    .Y(_08019_));
 sg13g2_or2_1 _38608_ (.X(_08020_),
    .B(\u_inv.d_next[10] ),
    .A(net7341));
 sg13g2_xnor2_1 _38609_ (.Y(_08021_),
    .A(_04260_),
    .B(_08018_));
 sg13g2_a21oi_1 _38610_ (.A1(net7341),
    .A2(_08021_),
    .Y(_08022_),
    .B1(net6310));
 sg13g2_a22oi_1 _38611_ (.Y(_08023_),
    .B1(_08020_),
    .B2(_08022_),
    .A2(_08017_),
    .A1(net6310));
 sg13g2_nor2_1 _38612_ (.A(net5846),
    .B(_08023_),
    .Y(_08024_));
 sg13g2_xnor2_1 _38613_ (.Y(_08025_),
    .A(net5846),
    .B(_08023_));
 sg13g2_nor2_1 _38614_ (.A(_04254_),
    .B(_08019_),
    .Y(_08026_));
 sg13g2_and2_1 _38615_ (.A(_04253_),
    .B(_08026_),
    .X(_08027_));
 sg13g2_o21ai_1 _38616_ (.B1(net7339),
    .Y(_08028_),
    .A1(_04253_),
    .A2(_08026_));
 sg13g2_a21oi_1 _38617_ (.A1(net7204),
    .A2(\u_inv.d_next[11] ),
    .Y(_08029_),
    .B1(net6307));
 sg13g2_o21ai_1 _38618_ (.B1(_08029_),
    .Y(_08030_),
    .A1(_08027_),
    .A2(_08028_));
 sg13g2_nor2_1 _38619_ (.A(_04894_),
    .B(_08016_),
    .Y(_08031_));
 sg13g2_xnor2_1 _38620_ (.Y(_08032_),
    .A(_04253_),
    .B(_08031_));
 sg13g2_o21ai_1 _38621_ (.B1(_08030_),
    .Y(_08033_),
    .A1(net6224),
    .A2(_08032_));
 sg13g2_xnor2_1 _38622_ (.Y(_08034_),
    .A(net5846),
    .B(_08033_));
 sg13g2_nor2_1 _38623_ (.A(_08025_),
    .B(_08034_),
    .Y(_08035_));
 sg13g2_a21oi_1 _38624_ (.A1(_04290_),
    .A2(_04912_),
    .Y(_08036_),
    .B1(_04914_));
 sg13g2_o21ai_1 _38625_ (.B1(net6307),
    .Y(_08037_),
    .A1(_04255_),
    .A2(_08036_));
 sg13g2_a21oi_1 _38626_ (.A1(_04255_),
    .A2(_08036_),
    .Y(_08038_),
    .B1(_08037_));
 sg13g2_nand3_1 _38627_ (.B(_04256_),
    .C(_04291_),
    .A(_04255_),
    .Y(_08039_));
 sg13g2_o21ai_1 _38628_ (.B1(net7341),
    .Y(_08040_),
    .A1(_04255_),
    .A2(_04256_));
 sg13g2_nor2_1 _38629_ (.A(_04292_),
    .B(_08040_),
    .Y(_08041_));
 sg13g2_a221oi_1 _38630_ (.B2(_08041_),
    .C1(net6307),
    .B1(_08039_),
    .A1(net7204),
    .Y(_08042_),
    .A2(\u_inv.d_next[9] ));
 sg13g2_nor2_2 _38631_ (.A(_08038_),
    .B(_08042_),
    .Y(_08043_));
 sg13g2_nand2_1 _38632_ (.Y(_08044_),
    .A(net5847),
    .B(_08043_));
 sg13g2_nor2_1 _38633_ (.A(net5847),
    .B(_08043_),
    .Y(_08045_));
 sg13g2_xnor2_1 _38634_ (.Y(_08046_),
    .A(net5795),
    .B(_08043_));
 sg13g2_xor2_1 _38635_ (.B(_04912_),
    .A(_04290_),
    .X(_08047_));
 sg13g2_xnor2_1 _38636_ (.Y(_08048_),
    .A(_04289_),
    .B(_04290_));
 sg13g2_o21ai_1 _38637_ (.B1(net6224),
    .Y(_08049_),
    .A1(net7341),
    .A2(\u_inv.d_next[8] ));
 sg13g2_a21oi_1 _38638_ (.A1(net7341),
    .A2(_08048_),
    .Y(_08050_),
    .B1(_08049_));
 sg13g2_a21oi_1 _38639_ (.A1(net6307),
    .A2(_08047_),
    .Y(_08051_),
    .B1(_08050_));
 sg13g2_or2_1 _38640_ (.X(_08052_),
    .B(_08051_),
    .A(net5795));
 sg13g2_xnor2_1 _38641_ (.Y(_08053_),
    .A(net5846),
    .B(_08051_));
 sg13g2_nand3_1 _38642_ (.B(_08046_),
    .C(_08053_),
    .A(_08035_),
    .Y(_08054_));
 sg13g2_a21oi_2 _38643_ (.B1(_08054_),
    .Y(_08055_),
    .A2(_08013_),
    .A1(_08012_));
 sg13g2_o21ai_1 _38644_ (.B1(_04895_),
    .Y(_08056_),
    .A1(_04886_),
    .A2(_08015_));
 sg13g2_a21oi_1 _38645_ (.A1(_04884_),
    .A2(_08056_),
    .Y(_08057_),
    .B1(_04889_));
 sg13g2_a21oi_1 _38646_ (.A1(_04890_),
    .A2(_08057_),
    .Y(_08058_),
    .B1(_04244_));
 sg13g2_a21oi_1 _38647_ (.A1(\u_inv.d_next[14] ),
    .A2(_18600_),
    .Y(_08059_),
    .B1(_08058_));
 sg13g2_o21ai_1 _38648_ (.B1(net6307),
    .Y(_08060_),
    .A1(_04248_),
    .A2(_08059_));
 sg13g2_a21oi_1 _38649_ (.A1(_04248_),
    .A2(_08059_),
    .Y(_08061_),
    .B1(_08060_));
 sg13g2_a21oi_2 _38650_ (.B1(_04262_),
    .Y(_08062_),
    .A2(_04293_),
    .A1(_04292_));
 sg13g2_nor2_1 _38651_ (.A(_04241_),
    .B(_08062_),
    .Y(_08063_));
 sg13g2_nor2_1 _38652_ (.A(_04263_),
    .B(_08063_),
    .Y(_08064_));
 sg13g2_o21ai_1 _38653_ (.B1(_04244_),
    .Y(_08065_),
    .A1(_04263_),
    .A2(_08063_));
 sg13g2_a21oi_1 _38654_ (.A1(_04243_),
    .A2(_08065_),
    .Y(_08066_),
    .B1(_04248_));
 sg13g2_nand3_1 _38655_ (.B(_04248_),
    .C(_08065_),
    .A(_04243_),
    .Y(_08067_));
 sg13g2_nor2_1 _38656_ (.A(net7204),
    .B(_08066_),
    .Y(_08068_));
 sg13g2_a221oi_1 _38657_ (.B2(_08068_),
    .C1(net6307),
    .B1(_08067_),
    .A1(net7204),
    .Y(_08069_),
    .A2(\u_inv.d_next[15] ));
 sg13g2_or2_1 _38658_ (.X(_08070_),
    .B(_08069_),
    .A(_08061_));
 sg13g2_xnor2_1 _38659_ (.Y(_08071_),
    .A(net5848),
    .B(_08070_));
 sg13g2_xnor2_1 _38660_ (.Y(_08072_),
    .A(_04245_),
    .B(_08064_));
 sg13g2_nor2_1 _38661_ (.A(net7341),
    .B(\u_inv.d_next[14] ),
    .Y(_08073_));
 sg13g2_a21oi_1 _38662_ (.A1(net7341),
    .A2(_08072_),
    .Y(_08074_),
    .B1(_08073_));
 sg13g2_nand3_1 _38663_ (.B(_04890_),
    .C(_08057_),
    .A(_04244_),
    .Y(_08075_));
 sg13g2_nor2_1 _38664_ (.A(net6224),
    .B(_08058_),
    .Y(_08076_));
 sg13g2_a22oi_1 _38665_ (.Y(_08077_),
    .B1(_08075_),
    .B2(_08076_),
    .A2(_08074_),
    .A1(net6224));
 sg13g2_or2_1 _38666_ (.X(_08078_),
    .B(_08077_),
    .A(net5848));
 sg13g2_inv_1 _38667_ (.Y(_08079_),
    .A(_08078_));
 sg13g2_xnor2_1 _38668_ (.Y(_08080_),
    .A(net5794),
    .B(_08077_));
 sg13g2_nor2b_1 _38669_ (.A(_08071_),
    .B_N(_08080_),
    .Y(_08081_));
 sg13g2_a21oi_1 _38670_ (.A1(_04240_),
    .A2(_08056_),
    .Y(_08082_),
    .B1(net6224));
 sg13g2_or2_1 _38671_ (.X(_08083_),
    .B(_08056_),
    .A(_04240_));
 sg13g2_xnor2_1 _38672_ (.Y(_08084_),
    .A(_04240_),
    .B(_08062_));
 sg13g2_nor2_1 _38673_ (.A(net7341),
    .B(\u_inv.d_next[12] ),
    .Y(_08085_));
 sg13g2_a21oi_1 _38674_ (.A1(net7342),
    .A2(_08084_),
    .Y(_08086_),
    .B1(_08085_));
 sg13g2_a22oi_1 _38675_ (.Y(_08087_),
    .B1(_08086_),
    .B2(net6227),
    .A2(_08083_),
    .A1(_08082_));
 sg13g2_or2_1 _38676_ (.X(_08088_),
    .B(_08087_),
    .A(net5846));
 sg13g2_xnor2_1 _38677_ (.Y(_08089_),
    .A(net5795),
    .B(_08087_));
 sg13g2_nor2_1 _38678_ (.A(net6227),
    .B(_08057_),
    .Y(_08090_));
 sg13g2_and2_1 _38679_ (.A(_04237_),
    .B(_04888_),
    .X(_08091_));
 sg13g2_o21ai_1 _38680_ (.B1(_04238_),
    .Y(_08092_),
    .A1(_04240_),
    .A2(_08062_));
 sg13g2_o21ai_1 _38681_ (.B1(net7342),
    .Y(_08093_),
    .A1(_04237_),
    .A2(_08092_));
 sg13g2_a21o_1 _38682_ (.A2(_08092_),
    .A1(_04237_),
    .B1(_08093_),
    .X(_08094_));
 sg13g2_a21oi_1 _38683_ (.A1(net7204),
    .A2(\u_inv.d_next[13] ),
    .Y(_08095_),
    .B1(net6310));
 sg13g2_a221oi_1 _38684_ (.B2(_08095_),
    .C1(_08090_),
    .B1(_08094_),
    .A1(_08082_),
    .Y(_08096_),
    .A2(_08091_));
 sg13g2_nand2_1 _38685_ (.Y(_08097_),
    .A(net5794),
    .B(_08096_));
 sg13g2_nand2b_1 _38686_ (.Y(_08098_),
    .B(net5848),
    .A_N(_08096_));
 sg13g2_xnor2_1 _38687_ (.Y(_08099_),
    .A(net5846),
    .B(_08096_));
 sg13g2_nand2_1 _38688_ (.Y(_08100_),
    .A(_08089_),
    .B(_08099_));
 sg13g2_inv_1 _38689_ (.Y(_08101_),
    .A(_08100_));
 sg13g2_and2_1 _38690_ (.A(_08081_),
    .B(_08101_),
    .X(_08102_));
 sg13g2_and2_1 _38691_ (.A(_08088_),
    .B(_08097_),
    .X(_08103_));
 sg13g2_inv_1 _38692_ (.Y(_08104_),
    .A(_08103_));
 sg13g2_nand2_1 _38693_ (.Y(_08105_),
    .A(_08044_),
    .B(_08052_));
 sg13g2_a21oi_1 _38694_ (.A1(_08023_),
    .A2(_08033_),
    .Y(_08106_),
    .B1(net5847));
 sg13g2_a21o_1 _38695_ (.A2(_08105_),
    .A1(_08035_),
    .B1(_08106_),
    .X(_08107_));
 sg13g2_a21o_1 _38696_ (.A2(_08107_),
    .A1(_08101_),
    .B1(_08104_),
    .X(_08108_));
 sg13g2_o21ai_1 _38697_ (.B1(_08078_),
    .Y(_08109_),
    .A1(net5848),
    .A2(_08070_));
 sg13g2_a221oi_1 _38698_ (.B2(_08081_),
    .C1(_08109_),
    .B1(_08108_),
    .A1(_08055_),
    .Y(_08110_),
    .A2(_08102_));
 sg13g2_nor2_1 _38699_ (.A(net5795),
    .B(_07936_),
    .Y(_08111_));
 sg13g2_xnor2_1 _38700_ (.Y(_08112_),
    .A(net5794),
    .B(_07936_));
 sg13g2_xnor2_1 _38701_ (.Y(_08113_),
    .A(net5852),
    .B(_07943_));
 sg13g2_nand2b_1 _38702_ (.Y(_08114_),
    .B(_08113_),
    .A_N(_08112_));
 sg13g2_nor3_1 _38703_ (.A(_07918_),
    .B(_07927_),
    .C(_08114_),
    .Y(_08115_));
 sg13g2_nand4_1 _38704_ (.B(_07888_),
    .C(_07908_),
    .A(_07881_),
    .Y(_08116_),
    .D(_08115_));
 sg13g2_o21ai_1 _38705_ (.B1(_07952_),
    .Y(_08117_),
    .A1(_08116_),
    .A2(_08110_));
 sg13g2_nand2_1 _38706_ (.Y(_08118_),
    .A(_07860_),
    .B(net1083));
 sg13g2_nand2_1 _38707_ (.Y(_08119_),
    .A(net5858),
    .B(_07719_));
 sg13g2_xnor2_1 _38708_ (.Y(_08120_),
    .A(net5858),
    .B(_07719_));
 sg13g2_xnor2_1 _38709_ (.Y(_08121_),
    .A(net5809),
    .B(_07713_));
 sg13g2_nor2_1 _38710_ (.A(_08120_),
    .B(_08121_),
    .Y(_08122_));
 sg13g2_nand2_1 _38711_ (.Y(_08123_),
    .A(_07663_),
    .B(_08122_));
 sg13g2_nor4_1 _38712_ (.A(_07682_),
    .B(_07693_),
    .C(_07703_),
    .D(_08123_),
    .Y(_08124_));
 sg13g2_nor2b_2 _38713_ (.A(_07635_),
    .B_N(_08124_),
    .Y(_08125_));
 sg13g2_nand3_1 _38714_ (.B(net1083),
    .C(_08125_),
    .A(_07860_),
    .Y(_08126_));
 sg13g2_and4_1 _38715_ (.A(_07540_),
    .B(_07860_),
    .C(net1083),
    .D(_08125_),
    .X(_08127_));
 sg13g2_nand4_1 _38716_ (.B(_07860_),
    .C(net1083),
    .A(_07540_),
    .Y(_08128_),
    .D(_08125_));
 sg13g2_nor2_2 _38717_ (.A(_07758_),
    .B(_08127_),
    .Y(_08129_));
 sg13g2_nand2b_1 _38718_ (.Y(_08130_),
    .B(net5874),
    .A_N(_07319_));
 sg13g2_xnor2_1 _38719_ (.Y(_08131_),
    .A(net5831),
    .B(_07319_));
 sg13g2_xnor2_1 _38720_ (.Y(_08132_),
    .A(net5874),
    .B(_07324_));
 sg13g2_or3_1 _38721_ (.A(_07311_),
    .B(_08131_),
    .C(_08132_),
    .X(_08133_));
 sg13g2_inv_2 _38722_ (.Y(_08134_),
    .A(_08133_));
 sg13g2_and4_1 _38723_ (.A(_07199_),
    .B(_07218_),
    .C(_07238_),
    .D(_08134_),
    .X(_08135_));
 sg13g2_nand2_1 _38724_ (.Y(_08136_),
    .A(_07290_),
    .B(_08135_));
 sg13g2_and4_1 _38725_ (.A(_07046_),
    .B(_07139_),
    .C(_07290_),
    .D(_08135_),
    .X(_08137_));
 sg13g2_o21ai_1 _38726_ (.B1(_08137_),
    .Y(_08138_),
    .A1(_08127_),
    .A2(_07758_));
 sg13g2_nand2_1 _38727_ (.Y(_08139_),
    .A(_07358_),
    .B(net1097));
 sg13g2_o21ai_1 _38728_ (.B1(_05088_),
    .Y(_08140_),
    .A1(_04964_),
    .A2(_05030_));
 sg13g2_a21oi_1 _38729_ (.A1(_04995_),
    .A2(_08140_),
    .Y(_08141_),
    .B1(_05144_));
 sg13g2_a21o_1 _38730_ (.A2(_08140_),
    .A1(_04995_),
    .B1(_05144_),
    .X(_08142_));
 sg13g2_a21o_2 _38731_ (.A2(_08142_),
    .A1(_04979_),
    .B1(_05103_),
    .X(_08143_));
 sg13g2_a21oi_1 _38732_ (.A1(_04971_),
    .A2(_08143_),
    .Y(_08144_),
    .B1(_05105_));
 sg13g2_nand3_1 _38733_ (.B(_04971_),
    .C(_08143_),
    .A(_04970_),
    .Y(_08145_));
 sg13g2_a21o_1 _38734_ (.A2(_08145_),
    .A1(_05108_),
    .B1(_04968_),
    .X(_08146_));
 sg13g2_nand3_1 _38735_ (.B(_05112_),
    .C(_08146_),
    .A(_03813_),
    .Y(_08147_));
 sg13g2_a21o_1 _38736_ (.A2(_08146_),
    .A1(_05112_),
    .B1(_03813_),
    .X(_08148_));
 sg13g2_a21oi_1 _38737_ (.A1(_08147_),
    .A2(_08148_),
    .Y(_08149_),
    .B1(net6258));
 sg13g2_nor2b_1 _38738_ (.A(_04409_),
    .B_N(_04408_),
    .Y(_08150_));
 sg13g2_and2_1 _38739_ (.A(_04408_),
    .B(_04410_),
    .X(_08151_));
 sg13g2_nand4_1 _38740_ (.B(_03930_),
    .C(_04408_),
    .A(_03914_),
    .Y(_08152_),
    .D(_04410_));
 sg13g2_nand2_1 _38741_ (.Y(_08153_),
    .A(_03936_),
    .B(_08152_));
 sg13g2_a21oi_2 _38742_ (.B1(_03950_),
    .Y(_08154_),
    .A2(_04412_),
    .A1(_04408_));
 sg13g2_or2_1 _38743_ (.X(_08155_),
    .B(_08154_),
    .A(_03953_));
 sg13g2_o21ai_1 _38744_ (.B1(_03873_),
    .Y(_08156_),
    .A1(_03955_),
    .A2(_08154_));
 sg13g2_a21oi_2 _38745_ (.B1(_03830_),
    .Y(_08157_),
    .A2(_08156_),
    .A1(_03876_));
 sg13g2_o21ai_1 _38746_ (.B1(_03833_),
    .Y(_08158_),
    .A1(_03824_),
    .A2(_08157_));
 sg13g2_a21oi_1 _38747_ (.A1(_03818_),
    .A2(_08158_),
    .Y(_08159_),
    .B1(_03836_));
 sg13g2_nand2b_1 _38748_ (.Y(_08160_),
    .B(_03813_),
    .A_N(_08159_));
 sg13g2_xnor2_1 _38749_ (.Y(_08161_),
    .A(_03813_),
    .B(_08159_));
 sg13g2_nand2_1 _38750_ (.Y(_08162_),
    .A(net7230),
    .B(\u_inv.d_next[126] ));
 sg13g2_a21oi_1 _38751_ (.A1(net7390),
    .A2(_08161_),
    .Y(_08163_),
    .B1(net6349));
 sg13g2_a21oi_2 _38752_ (.B1(_08149_),
    .Y(_08164_),
    .A2(_08163_),
    .A1(_08162_));
 sg13g2_xnor2_1 _38753_ (.Y(_08165_),
    .A(net5818),
    .B(_08164_));
 sg13g2_nand3_1 _38754_ (.B(_03812_),
    .C(_08160_),
    .A(_03811_),
    .Y(_08166_));
 sg13g2_a21o_1 _38755_ (.A2(_08160_),
    .A1(_03812_),
    .B1(_03811_),
    .X(_08167_));
 sg13g2_nand3_1 _38756_ (.B(_08166_),
    .C(_08167_),
    .A(net7391),
    .Y(_08168_));
 sg13g2_nand2_1 _38757_ (.Y(_08169_),
    .A(net7230),
    .B(\u_inv.d_next[127] ));
 sg13g2_nand3_1 _38758_ (.B(_08168_),
    .C(_08169_),
    .A(net6258),
    .Y(_08170_));
 sg13g2_nand3_1 _38759_ (.B(_05113_),
    .C(_08148_),
    .A(_03811_),
    .Y(_08171_));
 sg13g2_a21o_1 _38760_ (.A2(_08148_),
    .A1(_05113_),
    .B1(_03811_),
    .X(_08172_));
 sg13g2_nand3_1 _38761_ (.B(_08171_),
    .C(_08172_),
    .A(net6349),
    .Y(_08173_));
 sg13g2_and3_2 _38762_ (.X(_08174_),
    .A(net5818),
    .B(_08170_),
    .C(_08173_));
 sg13g2_a21oi_1 _38763_ (.A1(_08170_),
    .A2(_08173_),
    .Y(_08175_),
    .B1(net5819));
 sg13g2_or2_1 _38764_ (.X(_08176_),
    .B(_08175_),
    .A(_08174_));
 sg13g2_nor3_1 _38765_ (.A(_08165_),
    .B(_08174_),
    .C(_08175_),
    .Y(_08177_));
 sg13g2_a21oi_1 _38766_ (.A1(_03817_),
    .A2(_08158_),
    .Y(_08178_),
    .B1(_03816_));
 sg13g2_o21ai_1 _38767_ (.B1(net7390),
    .Y(_08179_),
    .A1(_03815_),
    .A2(_08178_));
 sg13g2_a21o_1 _38768_ (.A2(_08178_),
    .A1(_03815_),
    .B1(_08179_),
    .X(_08180_));
 sg13g2_nand2_1 _38769_ (.Y(_08181_),
    .A(net7235),
    .B(\u_inv.d_next[125] ));
 sg13g2_nand3_1 _38770_ (.B(_08180_),
    .C(_08181_),
    .A(net6258),
    .Y(_08182_));
 sg13g2_a21o_1 _38771_ (.A2(_08145_),
    .A1(_05108_),
    .B1(_03817_),
    .X(_08183_));
 sg13g2_nand3_1 _38772_ (.B(_05109_),
    .C(_08183_),
    .A(_03815_),
    .Y(_08184_));
 sg13g2_a21oi_1 _38773_ (.A1(_05109_),
    .A2(_08183_),
    .Y(_08185_),
    .B1(_03815_));
 sg13g2_nand3b_1 _38774_ (.B(net6349),
    .C(_08184_),
    .Y(_08186_),
    .A_N(_08185_));
 sg13g2_nand3_1 _38775_ (.B(_08182_),
    .C(_08186_),
    .A(net5818),
    .Y(_08187_));
 sg13g2_a21o_1 _38776_ (.A2(_08186_),
    .A1(_08182_),
    .B1(net5818),
    .X(_08188_));
 sg13g2_nand2_1 _38777_ (.Y(_08189_),
    .A(_08187_),
    .B(_08188_));
 sg13g2_nand3_1 _38778_ (.B(_05108_),
    .C(_08145_),
    .A(_03817_),
    .Y(_08190_));
 sg13g2_and2_1 _38779_ (.A(_08183_),
    .B(_08190_),
    .X(_08191_));
 sg13g2_xnor2_1 _38780_ (.Y(_08192_),
    .A(_03817_),
    .B(_08158_));
 sg13g2_o21ai_1 _38781_ (.B1(net6258),
    .Y(_08193_),
    .A1(net7390),
    .A2(\u_inv.d_next[124] ));
 sg13g2_a21oi_1 _38782_ (.A1(net7390),
    .A2(_08192_),
    .Y(_08194_),
    .B1(_08193_));
 sg13g2_a21oi_1 _38783_ (.A1(net6349),
    .A2(_08191_),
    .Y(_08195_),
    .B1(_08194_));
 sg13g2_or2_1 _38784_ (.X(_08196_),
    .B(_08195_),
    .A(net5866));
 sg13g2_xnor2_1 _38785_ (.Y(_08197_),
    .A(net5818),
    .B(_08195_));
 sg13g2_nor2b_1 _38786_ (.A(_08189_),
    .B_N(_08197_),
    .Y(_08198_));
 sg13g2_nand3_1 _38787_ (.B(_08188_),
    .C(_08197_),
    .A(_08187_),
    .Y(_08199_));
 sg13g2_nor4_1 _38788_ (.A(_08165_),
    .B(_08174_),
    .C(_08175_),
    .D(_08199_),
    .Y(_08200_));
 sg13g2_o21ai_1 _38789_ (.B1(_03821_),
    .Y(_08201_),
    .A1(_03822_),
    .A2(_08157_));
 sg13g2_a21oi_1 _38790_ (.A1(_03820_),
    .A2(_08201_),
    .Y(_08202_),
    .B1(net7230));
 sg13g2_o21ai_1 _38791_ (.B1(_08202_),
    .Y(_08203_),
    .A1(_03820_),
    .A2(_08201_));
 sg13g2_a21oi_1 _38792_ (.A1(net7230),
    .A2(\u_inv.d_next[123] ),
    .Y(_08204_),
    .B1(net6349));
 sg13g2_nand2_1 _38793_ (.Y(_08205_),
    .A(_08203_),
    .B(_08204_));
 sg13g2_o21ai_1 _38794_ (.B1(_05106_),
    .Y(_08206_),
    .A1(_03823_),
    .A2(_08144_));
 sg13g2_xnor2_1 _38795_ (.Y(_08207_),
    .A(_03820_),
    .B(_08206_));
 sg13g2_o21ai_1 _38796_ (.B1(_08205_),
    .Y(_08208_),
    .A1(net6258),
    .A2(_08207_));
 sg13g2_xnor2_1 _38797_ (.Y(_08209_),
    .A(net5868),
    .B(_08208_));
 sg13g2_xor2_1 _38798_ (.B(_08144_),
    .A(_03823_),
    .X(_08210_));
 sg13g2_xor2_1 _38799_ (.B(_08157_),
    .A(_03823_),
    .X(_08211_));
 sg13g2_o21ai_1 _38800_ (.B1(net6248),
    .Y(_08212_),
    .A1(net7376),
    .A2(\u_inv.d_next[122] ));
 sg13g2_a21oi_1 _38801_ (.A1(net7390),
    .A2(_08211_),
    .Y(_08213_),
    .B1(_08212_));
 sg13g2_a21oi_1 _38802_ (.A1(net6349),
    .A2(_08210_),
    .Y(_08214_),
    .B1(_08213_));
 sg13g2_or2_1 _38803_ (.X(_08215_),
    .B(_08214_),
    .A(net5868));
 sg13g2_xnor2_1 _38804_ (.Y(_08216_),
    .A(net5826),
    .B(_08214_));
 sg13g2_inv_1 _38805_ (.Y(_08217_),
    .A(_08216_));
 sg13g2_nor2_1 _38806_ (.A(_08209_),
    .B(_08217_),
    .Y(_08218_));
 sg13g2_a21oi_1 _38807_ (.A1(_03874_),
    .A2(_08143_),
    .Y(_08219_),
    .B1(_05104_));
 sg13g2_o21ai_1 _38808_ (.B1(net6355),
    .Y(_08220_),
    .A1(_03827_),
    .A2(_08219_));
 sg13g2_a21oi_1 _38809_ (.A1(_03827_),
    .A2(_08219_),
    .Y(_08221_),
    .B1(_08220_));
 sg13g2_nand2_1 _38810_ (.Y(_08222_),
    .A(_03875_),
    .B(_08156_));
 sg13g2_and2_1 _38811_ (.A(_03828_),
    .B(_08222_),
    .X(_08223_));
 sg13g2_o21ai_1 _38812_ (.B1(net7390),
    .Y(_08224_),
    .A1(_03827_),
    .A2(_08223_));
 sg13g2_a21o_1 _38813_ (.A2(_08223_),
    .A1(_03827_),
    .B1(_08224_),
    .X(_08225_));
 sg13g2_a21oi_1 _38814_ (.A1(net7230),
    .A2(\u_inv.d_next[121] ),
    .Y(_08226_),
    .B1(net6349));
 sg13g2_a21oi_1 _38815_ (.A1(_08225_),
    .A2(_08226_),
    .Y(_08227_),
    .B1(_08221_));
 sg13g2_nand2_1 _38816_ (.Y(_08228_),
    .A(net5826),
    .B(_08227_));
 sg13g2_xnor2_1 _38817_ (.Y(_08229_),
    .A(net5818),
    .B(_08227_));
 sg13g2_xnor2_1 _38818_ (.Y(_08230_),
    .A(_03874_),
    .B(_08143_));
 sg13g2_xnor2_1 _38819_ (.Y(_08231_),
    .A(_03875_),
    .B(_08156_));
 sg13g2_o21ai_1 _38820_ (.B1(net6258),
    .Y(_08232_),
    .A1(net7390),
    .A2(\u_inv.d_next[120] ));
 sg13g2_a21o_1 _38821_ (.A2(_08231_),
    .A1(net7390),
    .B1(_08232_),
    .X(_08233_));
 sg13g2_o21ai_1 _38822_ (.B1(_08233_),
    .Y(_08234_),
    .A1(net6258),
    .A2(_08230_));
 sg13g2_nand2_1 _38823_ (.Y(_08235_),
    .A(net5826),
    .B(_08234_));
 sg13g2_xnor2_1 _38824_ (.Y(_08236_),
    .A(net5868),
    .B(_08234_));
 sg13g2_nand2b_1 _38825_ (.Y(_08237_),
    .B(_08236_),
    .A_N(_08229_));
 sg13g2_inv_1 _38826_ (.Y(_08238_),
    .A(_08237_));
 sg13g2_nand2_1 _38827_ (.Y(_08239_),
    .A(_08218_),
    .B(_08238_));
 sg13g2_nand3_1 _38828_ (.B(_08218_),
    .C(_08238_),
    .A(_08200_),
    .Y(_08240_));
 sg13g2_nor3_1 _38829_ (.A(_03859_),
    .B(_03951_),
    .C(_08141_),
    .Y(_08241_));
 sg13g2_nor2_1 _38830_ (.A(_05090_),
    .B(_08241_),
    .Y(_08242_));
 sg13g2_o21ai_1 _38831_ (.B1(_04977_),
    .Y(_08243_),
    .A1(_05090_),
    .A2(_08241_));
 sg13g2_nand2_1 _38832_ (.Y(_08244_),
    .A(_05094_),
    .B(_08243_));
 sg13g2_a21oi_1 _38833_ (.A1(_05094_),
    .A2(_08243_),
    .Y(_08245_),
    .B1(_04974_));
 sg13g2_nor2_1 _38834_ (.A(_05101_),
    .B(_08245_),
    .Y(_08246_));
 sg13g2_o21ai_1 _38835_ (.B1(_03846_),
    .Y(_08247_),
    .A1(_05101_),
    .A2(_08245_));
 sg13g2_xnor2_1 _38836_ (.Y(_08248_),
    .A(_03845_),
    .B(_08246_));
 sg13g2_o21ai_1 _38837_ (.B1(_03867_),
    .Y(_08249_),
    .A1(_03954_),
    .A2(_08154_));
 sg13g2_nand2_1 _38838_ (.Y(_08250_),
    .A(_03852_),
    .B(_08249_));
 sg13g2_a21oi_1 _38839_ (.A1(_03853_),
    .A2(_08249_),
    .Y(_08251_),
    .B1(_03870_));
 sg13g2_nand2b_1 _38840_ (.Y(_08252_),
    .B(_03845_),
    .A_N(_08251_));
 sg13g2_a21oi_1 _38841_ (.A1(_03846_),
    .A2(_08251_),
    .Y(_08253_),
    .B1(net7232));
 sg13g2_a221oi_1 _38842_ (.B2(_08253_),
    .C1(net6353),
    .B1(_08252_),
    .A1(net7232),
    .Y(_08254_),
    .A2(\u_inv.d_next[118] ));
 sg13g2_a21o_2 _38843_ (.A2(_08248_),
    .A1(net6354),
    .B1(_08254_),
    .X(_08255_));
 sg13g2_nand2b_1 _38844_ (.Y(_08256_),
    .B(net5825),
    .A_N(_08255_));
 sg13g2_xnor2_1 _38845_ (.Y(_08257_),
    .A(net5868),
    .B(_08255_));
 sg13g2_inv_1 _38846_ (.Y(_08258_),
    .A(_08257_));
 sg13g2_a21oi_1 _38847_ (.A1(_05096_),
    .A2(_08247_),
    .Y(_08259_),
    .B1(_03843_));
 sg13g2_nand3_1 _38848_ (.B(_05096_),
    .C(_08247_),
    .A(_03843_),
    .Y(_08260_));
 sg13g2_nand3b_1 _38849_ (.B(_08260_),
    .C(net6353),
    .Y(_08261_),
    .A_N(_08259_));
 sg13g2_a21oi_1 _38850_ (.A1(_03844_),
    .A2(_08252_),
    .Y(_08262_),
    .B1(_03843_));
 sg13g2_nand3_1 _38851_ (.B(_03844_),
    .C(_08252_),
    .A(_03843_),
    .Y(_08263_));
 sg13g2_nor2_1 _38852_ (.A(net7233),
    .B(_08262_),
    .Y(_08264_));
 sg13g2_a21oi_1 _38853_ (.A1(_08263_),
    .A2(_08264_),
    .Y(_08265_),
    .B1(net6353));
 sg13g2_o21ai_1 _38854_ (.B1(_08265_),
    .Y(_08266_),
    .A1(net7392),
    .A2(_18139_));
 sg13g2_nand2_1 _38855_ (.Y(_08267_),
    .A(_08261_),
    .B(_08266_));
 sg13g2_and3_1 _38856_ (.X(_08268_),
    .A(net5825),
    .B(_08261_),
    .C(_08266_));
 sg13g2_a21oi_1 _38857_ (.A1(_08261_),
    .A2(_08266_),
    .Y(_08269_),
    .B1(net5825));
 sg13g2_nor2_1 _38858_ (.A(_08268_),
    .B(_08269_),
    .Y(_08270_));
 sg13g2_nor3_1 _38859_ (.A(_08257_),
    .B(_08268_),
    .C(_08269_),
    .Y(_08271_));
 sg13g2_a21oi_1 _38860_ (.A1(_05094_),
    .A2(_08243_),
    .Y(_08272_),
    .B1(_03852_));
 sg13g2_o21ai_1 _38861_ (.B1(_03850_),
    .Y(_08273_),
    .A1(_05099_),
    .A2(_08272_));
 sg13g2_nand3b_1 _38862_ (.B(_03849_),
    .C(_05100_),
    .Y(_08274_),
    .A_N(_08272_));
 sg13g2_and3_2 _38863_ (.X(_08275_),
    .A(net6353),
    .B(_08273_),
    .C(_08274_));
 sg13g2_and2_1 _38864_ (.A(_03851_),
    .B(_08250_),
    .X(_08276_));
 sg13g2_o21ai_1 _38865_ (.B1(net7392),
    .Y(_08277_),
    .A1(_03849_),
    .A2(_08276_));
 sg13g2_a21oi_1 _38866_ (.A1(_03849_),
    .A2(_08276_),
    .Y(_08278_),
    .B1(_08277_));
 sg13g2_a21oi_1 _38867_ (.A1(net7232),
    .A2(\u_inv.d_next[117] ),
    .Y(_08279_),
    .B1(net6354));
 sg13g2_nand2b_1 _38868_ (.Y(_08280_),
    .B(_08279_),
    .A_N(_08278_));
 sg13g2_inv_2 _38869_ (.Y(_08281_),
    .A(_08280_));
 sg13g2_nor2_1 _38870_ (.A(_08275_),
    .B(_08281_),
    .Y(_08282_));
 sg13g2_or3_1 _38871_ (.A(net5868),
    .B(_08275_),
    .C(_08281_),
    .X(_08283_));
 sg13g2_o21ai_1 _38872_ (.B1(net5868),
    .Y(_08284_),
    .A1(_08275_),
    .A2(_08281_));
 sg13g2_o21ai_1 _38873_ (.B1(net5826),
    .Y(_08285_),
    .A1(_08275_),
    .A2(_08281_));
 sg13g2_nand2_1 _38874_ (.Y(_08286_),
    .A(net5869),
    .B(_08282_));
 sg13g2_nand2_1 _38875_ (.Y(_08287_),
    .A(_08283_),
    .B(_08284_));
 sg13g2_xnor2_1 _38876_ (.Y(_08288_),
    .A(_03852_),
    .B(_08249_));
 sg13g2_o21ai_1 _38877_ (.B1(net6257),
    .Y(_08289_),
    .A1(net7392),
    .A2(\u_inv.d_next[116] ));
 sg13g2_a21oi_1 _38878_ (.A1(net7392),
    .A2(_08288_),
    .Y(_08290_),
    .B1(_08289_));
 sg13g2_xnor2_1 _38879_ (.Y(_08291_),
    .A(_03852_),
    .B(_08244_));
 sg13g2_a21oi_2 _38880_ (.B1(_08290_),
    .Y(_08292_),
    .A2(_08291_),
    .A1(net6354));
 sg13g2_nor2_1 _38881_ (.A(net5869),
    .B(_08292_),
    .Y(_08293_));
 sg13g2_xnor2_1 _38882_ (.Y(_08294_),
    .A(net5869),
    .B(_08292_));
 sg13g2_nand3b_1 _38883_ (.B(_08284_),
    .C(_08283_),
    .Y(_08295_),
    .A_N(_08294_));
 sg13g2_nor4_1 _38884_ (.A(_08257_),
    .B(_08268_),
    .C(_08269_),
    .D(_08295_),
    .Y(_08296_));
 sg13g2_o21ai_1 _38885_ (.B1(_03864_),
    .Y(_08297_),
    .A1(_05090_),
    .A2(_08241_));
 sg13g2_xnor2_1 _38886_ (.Y(_08298_),
    .A(_03864_),
    .B(_08242_));
 sg13g2_a21oi_1 _38887_ (.A1(_03862_),
    .A2(_08155_),
    .Y(_08299_),
    .B1(_03864_));
 sg13g2_nand3_1 _38888_ (.B(_03864_),
    .C(_08155_),
    .A(_03862_),
    .Y(_08300_));
 sg13g2_nand2_1 _38889_ (.Y(_08301_),
    .A(net7392),
    .B(_08300_));
 sg13g2_a21oi_1 _38890_ (.A1(net7232),
    .A2(\u_inv.d_next[114] ),
    .Y(_08302_),
    .B1(net6354));
 sg13g2_o21ai_1 _38891_ (.B1(_08302_),
    .Y(_08303_),
    .A1(_08299_),
    .A2(_08301_));
 sg13g2_o21ai_1 _38892_ (.B1(_08303_),
    .Y(_08304_),
    .A1(net6257),
    .A2(_08298_));
 sg13g2_nor2_1 _38893_ (.A(net5870),
    .B(_08304_),
    .Y(_08305_));
 sg13g2_xnor2_1 _38894_ (.Y(_08306_),
    .A(net5825),
    .B(_08304_));
 sg13g2_inv_1 _38895_ (.Y(_08307_),
    .A(_08306_));
 sg13g2_a21oi_1 _38896_ (.A1(\u_inv.d_next[114] ),
    .A2(\u_inv.d_reg[114] ),
    .Y(_08308_),
    .B1(_08299_));
 sg13g2_or2_1 _38897_ (.X(_08309_),
    .B(_08308_),
    .A(_03855_));
 sg13g2_a21oi_1 _38898_ (.A1(_03855_),
    .A2(_08308_),
    .Y(_08310_),
    .B1(net7233));
 sg13g2_a221oi_1 _38899_ (.B2(_08310_),
    .C1(net6354),
    .B1(_08309_),
    .A1(net7233),
    .Y(_08311_),
    .A2(\u_inv.d_next[115] ));
 sg13g2_nand2b_1 _38900_ (.Y(_08312_),
    .B(_08297_),
    .A_N(_05092_));
 sg13g2_xnor2_1 _38901_ (.Y(_08313_),
    .A(_03855_),
    .B(_08312_));
 sg13g2_a21o_1 _38902_ (.A2(_08313_),
    .A1(net6354),
    .B1(_08311_),
    .X(_08314_));
 sg13g2_nor2_1 _38903_ (.A(net5870),
    .B(_08314_),
    .Y(_08315_));
 sg13g2_xnor2_1 _38904_ (.Y(_08316_),
    .A(net5870),
    .B(_08314_));
 sg13g2_o21ai_1 _38905_ (.B1(_05089_),
    .Y(_08317_),
    .A1(_03951_),
    .A2(_08141_));
 sg13g2_or2_1 _38906_ (.X(_08318_),
    .B(_08317_),
    .A(_03859_));
 sg13g2_a21oi_1 _38907_ (.A1(_03859_),
    .A2(_08317_),
    .Y(_08319_),
    .B1(net6259));
 sg13g2_nor2b_1 _38908_ (.A(_03859_),
    .B_N(_03856_),
    .Y(_08320_));
 sg13g2_o21ai_1 _38909_ (.B1(_08320_),
    .Y(_08321_),
    .A1(_03952_),
    .A2(_08154_));
 sg13g2_nand4_1 _38910_ (.B(_03860_),
    .C(_08155_),
    .A(net7392),
    .Y(_08322_),
    .D(_08321_));
 sg13g2_a21oi_1 _38911_ (.A1(net7233),
    .A2(\u_inv.d_next[113] ),
    .Y(_08323_),
    .B1(net6354));
 sg13g2_a22oi_1 _38912_ (.Y(_08324_),
    .B1(_08322_),
    .B2(_08323_),
    .A2(_08319_),
    .A1(_08318_));
 sg13g2_xnor2_1 _38913_ (.Y(_08325_),
    .A(net5825),
    .B(_08324_));
 sg13g2_xnor2_1 _38914_ (.Y(_08326_),
    .A(_03952_),
    .B(_08154_));
 sg13g2_o21ai_1 _38915_ (.B1(net6259),
    .Y(_08327_),
    .A1(net7394),
    .A2(\u_inv.d_next[112] ));
 sg13g2_a21o_1 _38916_ (.A2(_08326_),
    .A1(net7394),
    .B1(_08327_),
    .X(_08328_));
 sg13g2_xnor2_1 _38917_ (.Y(_08329_),
    .A(_03951_),
    .B(_08141_));
 sg13g2_o21ai_1 _38918_ (.B1(_08328_),
    .Y(_08330_),
    .A1(net6259),
    .A2(_08329_));
 sg13g2_nand2_1 _38919_ (.Y(_08331_),
    .A(net5830),
    .B(_08330_));
 sg13g2_xnor2_1 _38920_ (.Y(_08332_),
    .A(net5830),
    .B(_08330_));
 sg13g2_inv_1 _38921_ (.Y(_08333_),
    .A(_08332_));
 sg13g2_nor4_1 _38922_ (.A(_08307_),
    .B(_08316_),
    .C(_08325_),
    .D(_08332_),
    .Y(_08334_));
 sg13g2_and2_1 _38923_ (.A(_08296_),
    .B(_08334_),
    .X(_08335_));
 sg13g2_nor2b_1 _38924_ (.A(_08240_),
    .B_N(_08335_),
    .Y(_08336_));
 sg13g2_a21oi_1 _38925_ (.A1(_03936_),
    .A2(_08152_),
    .Y(_08337_),
    .B1(_03899_));
 sg13g2_a21oi_1 _38926_ (.A1(_03936_),
    .A2(_08152_),
    .Y(_08338_),
    .B1(_03900_));
 sg13g2_or3_1 _38927_ (.A(_03894_),
    .B(_03938_),
    .C(_08338_),
    .X(_08339_));
 sg13g2_o21ai_1 _38928_ (.B1(_03894_),
    .Y(_08340_),
    .A1(_03938_),
    .A2(_08338_));
 sg13g2_nand3_1 _38929_ (.B(_08339_),
    .C(_08340_),
    .A(net7409),
    .Y(_08341_));
 sg13g2_nand2_1 _38930_ (.Y(_08342_),
    .A(net7242),
    .B(\u_inv.d_next[106] ));
 sg13g2_a21oi_1 _38931_ (.A1(_08341_),
    .A2(_08342_),
    .Y(_08343_),
    .B1(net6367));
 sg13g2_and2_1 _38932_ (.A(_04409_),
    .B(_08140_),
    .X(_08344_));
 sg13g2_nand3b_1 _38933_ (.B(_04993_),
    .C(_08140_),
    .Y(_08345_),
    .A_N(_04992_));
 sg13g2_nand2_1 _38934_ (.Y(_08346_),
    .A(_05131_),
    .B(_08345_));
 sg13g2_a21oi_2 _38935_ (.B1(_04987_),
    .Y(_08347_),
    .A2(_08345_),
    .A1(_05131_));
 sg13g2_nor3_1 _38936_ (.A(_03893_),
    .B(_05134_),
    .C(_08347_),
    .Y(_08348_));
 sg13g2_o21ai_1 _38937_ (.B1(_03893_),
    .Y(_08349_),
    .A1(_05134_),
    .A2(_08347_));
 sg13g2_nor2b_1 _38938_ (.A(_08348_),
    .B_N(_08349_),
    .Y(_08350_));
 sg13g2_a21oi_1 _38939_ (.A1(net6367),
    .A2(_08350_),
    .Y(_08351_),
    .B1(_08343_));
 sg13g2_or2_1 _38940_ (.X(_08352_),
    .B(_08351_),
    .A(net5876));
 sg13g2_xnor2_1 _38941_ (.Y(_08353_),
    .A(net5876),
    .B(_08351_));
 sg13g2_a21o_1 _38942_ (.A2(_08349_),
    .A1(_05135_),
    .B1(_03891_),
    .X(_08354_));
 sg13g2_nand3_1 _38943_ (.B(_05135_),
    .C(_08349_),
    .A(_03891_),
    .Y(_08355_));
 sg13g2_nand3_1 _38944_ (.B(_08354_),
    .C(_08355_),
    .A(net6367),
    .Y(_08356_));
 sg13g2_o21ai_1 _38945_ (.B1(_08340_),
    .Y(_08357_),
    .A1(_18144_),
    .A2(_18508_));
 sg13g2_xnor2_1 _38946_ (.Y(_08358_),
    .A(_03892_),
    .B(_08357_));
 sg13g2_a21oi_1 _38947_ (.A1(net7242),
    .A2(\u_inv.d_next[107] ),
    .Y(_08359_),
    .B1(net6367));
 sg13g2_o21ai_1 _38948_ (.B1(_08359_),
    .Y(_08360_),
    .A1(net7242),
    .A2(_08358_));
 sg13g2_nand2_1 _38949_ (.Y(_08361_),
    .A(_08356_),
    .B(_08360_));
 sg13g2_xnor2_1 _38950_ (.Y(_08362_),
    .A(net5876),
    .B(_08361_));
 sg13g2_or3_1 _38951_ (.A(_03896_),
    .B(_03897_),
    .C(_08337_),
    .X(_08363_));
 sg13g2_o21ai_1 _38952_ (.B1(_03896_),
    .Y(_08364_),
    .A1(_03897_),
    .A2(_08337_));
 sg13g2_nand3_1 _38953_ (.B(_08363_),
    .C(_08364_),
    .A(net7409),
    .Y(_08365_));
 sg13g2_a21oi_1 _38954_ (.A1(net7242),
    .A2(\u_inv.d_next[105] ),
    .Y(_08366_),
    .B1(net6367));
 sg13g2_a21oi_1 _38955_ (.A1(_03899_),
    .A2(_08346_),
    .Y(_08367_),
    .B1(_05132_));
 sg13g2_xnor2_1 _38956_ (.Y(_08368_),
    .A(_03896_),
    .B(_08367_));
 sg13g2_a22oi_1 _38957_ (.Y(_08369_),
    .B1(_08368_),
    .B2(net6367),
    .A2(_08366_),
    .A1(_08365_));
 sg13g2_xnor2_1 _38958_ (.Y(_08370_),
    .A(net5876),
    .B(_08369_));
 sg13g2_xnor2_1 _38959_ (.Y(_08371_),
    .A(_03899_),
    .B(_08346_));
 sg13g2_o21ai_1 _38960_ (.B1(net7409),
    .Y(_08372_),
    .A1(_03898_),
    .A2(_08153_));
 sg13g2_or2_1 _38961_ (.X(_08373_),
    .B(_08372_),
    .A(_08337_));
 sg13g2_a21oi_1 _38962_ (.A1(net7241),
    .A2(\u_inv.d_next[104] ),
    .Y(_08374_),
    .B1(net6366));
 sg13g2_a22oi_1 _38963_ (.Y(_08375_),
    .B1(_08373_),
    .B2(_08374_),
    .A2(_08371_),
    .A1(net6366));
 sg13g2_and2_1 _38964_ (.A(net5832),
    .B(_08375_),
    .X(_08376_));
 sg13g2_xnor2_1 _38965_ (.Y(_08377_),
    .A(net5876),
    .B(_08375_));
 sg13g2_nand2_1 _38966_ (.Y(_08378_),
    .A(_08370_),
    .B(_08377_));
 sg13g2_nor3_2 _38967_ (.A(_08353_),
    .B(_08362_),
    .C(_08378_),
    .Y(_08379_));
 sg13g2_a21oi_1 _38968_ (.A1(_03895_),
    .A2(_08338_),
    .Y(_08380_),
    .B1(_03942_));
 sg13g2_nor2_1 _38969_ (.A(_03884_),
    .B(_08380_),
    .Y(_08381_));
 sg13g2_nor3_1 _38970_ (.A(_03884_),
    .B(_03887_),
    .C(_08380_),
    .Y(_08382_));
 sg13g2_nor2_1 _38971_ (.A(_03945_),
    .B(_08382_),
    .Y(_08383_));
 sg13g2_o21ai_1 _38972_ (.B1(_03880_),
    .Y(_08384_),
    .A1(_03945_),
    .A2(_08382_));
 sg13g2_xor2_1 _38973_ (.B(_08383_),
    .A(_03880_),
    .X(_08385_));
 sg13g2_o21ai_1 _38974_ (.B1(net6268),
    .Y(_08386_),
    .A1(net7409),
    .A2(\u_inv.d_next[110] ));
 sg13g2_a21oi_1 _38975_ (.A1(net7409),
    .A2(_08385_),
    .Y(_08387_),
    .B1(_08386_));
 sg13g2_a21oi_1 _38976_ (.A1(_04985_),
    .A2(_08347_),
    .Y(_08388_),
    .B1(_05137_));
 sg13g2_a21o_1 _38977_ (.A2(_08347_),
    .A1(_04985_),
    .B1(_05137_),
    .X(_08389_));
 sg13g2_a21oi_1 _38978_ (.A1(_04983_),
    .A2(_08389_),
    .Y(_08390_),
    .B1(_05139_));
 sg13g2_xor2_1 _38979_ (.B(_08390_),
    .A(_03880_),
    .X(_08391_));
 sg13g2_a21oi_2 _38980_ (.B1(_08387_),
    .Y(_08392_),
    .A2(_08391_),
    .A1(net6366));
 sg13g2_or2_1 _38981_ (.X(_08393_),
    .B(_08392_),
    .A(net5876));
 sg13g2_xnor2_1 _38982_ (.Y(_08394_),
    .A(net5833),
    .B(_08392_));
 sg13g2_xnor2_1 _38983_ (.Y(_08395_),
    .A(net5876),
    .B(_08392_));
 sg13g2_o21ai_1 _38984_ (.B1(_05141_),
    .Y(_08396_),
    .A1(_03880_),
    .A2(_08390_));
 sg13g2_nand2b_1 _38985_ (.Y(_08397_),
    .B(_03878_),
    .A_N(_08396_));
 sg13g2_a21oi_1 _38986_ (.A1(_03877_),
    .A2(_08396_),
    .Y(_08398_),
    .B1(net6269));
 sg13g2_nand3_1 _38987_ (.B(_03879_),
    .C(_08384_),
    .A(_03878_),
    .Y(_08399_));
 sg13g2_a21o_1 _38988_ (.A2(_08384_),
    .A1(_03879_),
    .B1(_03878_),
    .X(_08400_));
 sg13g2_nand3_1 _38989_ (.B(_08399_),
    .C(_08400_),
    .A(net7409),
    .Y(_08401_));
 sg13g2_a21oi_1 _38990_ (.A1(net7241),
    .A2(\u_inv.d_next[111] ),
    .Y(_08402_),
    .B1(net6366));
 sg13g2_a22oi_1 _38991_ (.Y(_08403_),
    .B1(_08401_),
    .B2(_08402_),
    .A2(_08398_),
    .A1(_08397_));
 sg13g2_nand2_1 _38992_ (.Y(_08404_),
    .A(net5832),
    .B(_08403_));
 sg13g2_xnor2_1 _38993_ (.Y(_08405_),
    .A(net5876),
    .B(_08403_));
 sg13g2_and2_1 _38994_ (.A(_08394_),
    .B(_08405_),
    .X(_08406_));
 sg13g2_o21ai_1 _38995_ (.B1(_05138_),
    .Y(_08407_),
    .A1(_03883_),
    .A2(_08388_));
 sg13g2_or2_1 _38996_ (.X(_08408_),
    .B(_08407_),
    .A(_03888_));
 sg13g2_a21oi_1 _38997_ (.A1(_03888_),
    .A2(_08407_),
    .Y(_08409_),
    .B1(net6269));
 sg13g2_nand2_1 _38998_ (.Y(_08410_),
    .A(_03882_),
    .B(_03887_));
 sg13g2_nor2_1 _38999_ (.A(_08381_),
    .B(_08410_),
    .Y(_08411_));
 sg13g2_nor4_1 _39000_ (.A(net7241),
    .B(_03943_),
    .C(_08382_),
    .D(_08411_),
    .Y(_08412_));
 sg13g2_a21oi_1 _39001_ (.A1(net7241),
    .A2(\u_inv.d_next[109] ),
    .Y(_08413_),
    .B1(_08412_));
 sg13g2_a22oi_1 _39002_ (.Y(_08414_),
    .B1(_08413_),
    .B2(net6269),
    .A2(_08409_),
    .A1(_08408_));
 sg13g2_nand2_1 _39003_ (.Y(_08415_),
    .A(net5832),
    .B(_08414_));
 sg13g2_xnor2_1 _39004_ (.Y(_08416_),
    .A(net5832),
    .B(_08414_));
 sg13g2_nand2_1 _39005_ (.Y(_08417_),
    .A(_03884_),
    .B(_08380_));
 sg13g2_nor2_1 _39006_ (.A(net7242),
    .B(_08381_),
    .Y(_08418_));
 sg13g2_xnor2_1 _39007_ (.Y(_08419_),
    .A(_03883_),
    .B(_08388_));
 sg13g2_a221oi_1 _39008_ (.B2(_08418_),
    .C1(net6366),
    .B1(_08417_),
    .A1(net7242),
    .Y(_08420_),
    .A2(\u_inv.d_next[108] ));
 sg13g2_a21oi_1 _39009_ (.A1(net6367),
    .A2(_08419_),
    .Y(_08421_),
    .B1(_08420_));
 sg13g2_nand2_1 _39010_ (.Y(_08422_),
    .A(net5832),
    .B(_08421_));
 sg13g2_xnor2_1 _39011_ (.Y(_08423_),
    .A(net5832),
    .B(_08421_));
 sg13g2_nor2_1 _39012_ (.A(_08416_),
    .B(_08423_),
    .Y(_08424_));
 sg13g2_and3_1 _39013_ (.X(_08425_),
    .A(_08394_),
    .B(_08405_),
    .C(_08424_));
 sg13g2_nand4_1 _39014_ (.B(_08394_),
    .C(_08405_),
    .A(_08379_),
    .Y(_08426_),
    .D(_08424_));
 sg13g2_a21oi_2 _39015_ (.B1(_03932_),
    .Y(_08427_),
    .A2(_08151_),
    .A1(_03930_));
 sg13g2_nor2_1 _39016_ (.A(_03909_),
    .B(_08427_),
    .Y(_08428_));
 sg13g2_nor2_1 _39017_ (.A(_03933_),
    .B(_08428_),
    .Y(_08429_));
 sg13g2_nor2_1 _39018_ (.A(_03911_),
    .B(_08429_),
    .Y(_08430_));
 sg13g2_a21oi_1 _39019_ (.A1(_03911_),
    .A2(_08429_),
    .Y(_08431_),
    .B1(net7241));
 sg13g2_nand2b_1 _39020_ (.Y(_08432_),
    .B(_08431_),
    .A_N(_08430_));
 sg13g2_a21oi_2 _39021_ (.B1(_05119_),
    .Y(_08433_),
    .A2(_08140_),
    .A1(_04993_));
 sg13g2_o21ai_1 _39022_ (.B1(_05129_),
    .Y(_08434_),
    .A1(_04991_),
    .A2(_08433_));
 sg13g2_a21oi_1 _39023_ (.A1(_03904_),
    .A2(_08434_),
    .Y(_08435_),
    .B1(_05121_));
 sg13g2_o21ai_1 _39024_ (.B1(_05123_),
    .Y(_08436_),
    .A1(_03907_),
    .A2(_08435_));
 sg13g2_xnor2_1 _39025_ (.Y(_08437_),
    .A(_03911_),
    .B(_08436_));
 sg13g2_a21oi_1 _39026_ (.A1(net7241),
    .A2(\u_inv.d_next[102] ),
    .Y(_08438_),
    .B1(net6366));
 sg13g2_a22oi_1 _39027_ (.Y(_08439_),
    .B1(_08438_),
    .B2(_08432_),
    .A2(_08437_),
    .A1(net6366));
 sg13g2_nand2_1 _39028_ (.Y(_08440_),
    .A(net5830),
    .B(_08439_));
 sg13g2_xnor2_1 _39029_ (.Y(_08441_),
    .A(net5830),
    .B(_08439_));
 sg13g2_inv_1 _39030_ (.Y(_08442_),
    .A(_08441_));
 sg13g2_a21oi_1 _39031_ (.A1(_03911_),
    .A2(_08436_),
    .Y(_08443_),
    .B1(_05125_));
 sg13g2_or2_1 _39032_ (.X(_08444_),
    .B(_08443_),
    .A(_03913_));
 sg13g2_a21oi_1 _39033_ (.A1(_03913_),
    .A2(_08443_),
    .Y(_08445_),
    .B1(net6269));
 sg13g2_a21oi_1 _39034_ (.A1(\u_inv.d_next[102] ),
    .A2(\u_inv.d_reg[102] ),
    .Y(_08446_),
    .B1(_08430_));
 sg13g2_a21oi_1 _39035_ (.A1(_03913_),
    .A2(_08446_),
    .Y(_08447_),
    .B1(net7241));
 sg13g2_o21ai_1 _39036_ (.B1(_08447_),
    .Y(_08448_),
    .A1(_03913_),
    .A2(_08446_));
 sg13g2_a21oi_1 _39037_ (.A1(net7241),
    .A2(\u_inv.d_next[103] ),
    .Y(_08449_),
    .B1(net6366));
 sg13g2_a22oi_1 _39038_ (.Y(_08450_),
    .B1(_08448_),
    .B2(_08449_),
    .A2(_08445_),
    .A1(_08444_));
 sg13g2_nand2_1 _39039_ (.Y(_08451_),
    .A(net5830),
    .B(_08450_));
 sg13g2_xnor2_1 _39040_ (.Y(_08452_),
    .A(net5830),
    .B(_08450_));
 sg13g2_nor2_1 _39041_ (.A(_08441_),
    .B(_08452_),
    .Y(_08453_));
 sg13g2_o21ai_1 _39042_ (.B1(_03903_),
    .Y(_08454_),
    .A1(_03904_),
    .A2(_08427_));
 sg13g2_o21ai_1 _39043_ (.B1(net7405),
    .Y(_08455_),
    .A1(_03907_),
    .A2(_08454_));
 sg13g2_a21oi_1 _39044_ (.A1(_03907_),
    .A2(_08454_),
    .Y(_08456_),
    .B1(_08455_));
 sg13g2_a21oi_1 _39045_ (.A1(net7239),
    .A2(\u_inv.d_next[101] ),
    .Y(_08457_),
    .B1(_08456_));
 sg13g2_xnor2_1 _39046_ (.Y(_08458_),
    .A(_03907_),
    .B(_08435_));
 sg13g2_mux2_1 _39047_ (.A0(_08457_),
    .A1(_08458_),
    .S(net6362),
    .X(_08459_));
 sg13g2_xnor2_1 _39048_ (.Y(_08460_),
    .A(net5875),
    .B(_08459_));
 sg13g2_xnor2_1 _39049_ (.Y(_08461_),
    .A(_03904_),
    .B(_08427_));
 sg13g2_o21ai_1 _39050_ (.B1(net6267),
    .Y(_08462_),
    .A1(net7405),
    .A2(\u_inv.d_next[100] ));
 sg13g2_a21oi_1 _39051_ (.A1(net7405),
    .A2(_08461_),
    .Y(_08463_),
    .B1(_08462_));
 sg13g2_xor2_1 _39052_ (.B(_08434_),
    .A(_03904_),
    .X(_08464_));
 sg13g2_a21oi_1 _39053_ (.A1(net6362),
    .A2(_08464_),
    .Y(_08465_),
    .B1(_08463_));
 sg13g2_or2_1 _39054_ (.X(_08466_),
    .B(_08465_),
    .A(net5875));
 sg13g2_xnor2_1 _39055_ (.Y(_08467_),
    .A(net5875),
    .B(_08465_));
 sg13g2_nor4_1 _39056_ (.A(_08441_),
    .B(_08452_),
    .C(_08460_),
    .D(_08467_),
    .Y(_08468_));
 sg13g2_or4_1 _39057_ (.A(_08441_),
    .B(_08452_),
    .C(_08460_),
    .D(_08467_),
    .X(_08469_));
 sg13g2_a21oi_1 _39058_ (.A1(_03919_),
    .A2(_03920_),
    .Y(_08470_),
    .B1(_08433_));
 sg13g2_o21ai_1 _39059_ (.B1(_03918_),
    .Y(_08471_),
    .A1(_05128_),
    .A2(_08470_));
 sg13g2_nor3_1 _39060_ (.A(_03918_),
    .B(_05128_),
    .C(_08470_),
    .Y(_08472_));
 sg13g2_nand2_1 _39061_ (.Y(_08473_),
    .A(net6363),
    .B(_08471_));
 sg13g2_nor2_1 _39062_ (.A(_03927_),
    .B(_08151_),
    .Y(_08474_));
 sg13g2_o21ai_1 _39063_ (.B1(_03919_),
    .Y(_08475_),
    .A1(_03929_),
    .A2(_08474_));
 sg13g2_a21oi_1 _39064_ (.A1(_03918_),
    .A2(_08475_),
    .Y(_08476_),
    .B1(net7239));
 sg13g2_o21ai_1 _39065_ (.B1(_08476_),
    .Y(_08477_),
    .A1(_03918_),
    .A2(_08475_));
 sg13g2_a21oi_1 _39066_ (.A1(net7239),
    .A2(\u_inv.d_next[99] ),
    .Y(_08478_),
    .B1(net6363));
 sg13g2_nand2_1 _39067_ (.Y(_08479_),
    .A(_08477_),
    .B(_08478_));
 sg13g2_o21ai_1 _39068_ (.B1(_08479_),
    .Y(_08480_),
    .A1(_08472_),
    .A2(_08473_));
 sg13g2_xnor2_1 _39069_ (.Y(_08481_),
    .A(net5874),
    .B(_08480_));
 sg13g2_xnor2_1 _39070_ (.Y(_08482_),
    .A(_03929_),
    .B(_08474_));
 sg13g2_o21ai_1 _39071_ (.B1(net6270),
    .Y(_08483_),
    .A1(net7406),
    .A2(\u_inv.d_next[98] ));
 sg13g2_a21oi_1 _39072_ (.A1(net7406),
    .A2(_08482_),
    .Y(_08484_),
    .B1(_08483_));
 sg13g2_xnor2_1 _39073_ (.Y(_08485_),
    .A(_03929_),
    .B(_08433_));
 sg13g2_a21oi_2 _39074_ (.B1(_08484_),
    .Y(_08486_),
    .A2(_08485_),
    .A1(net6363));
 sg13g2_or2_1 _39075_ (.X(_08487_),
    .B(_08486_),
    .A(net5874));
 sg13g2_xnor2_1 _39076_ (.Y(_08488_),
    .A(net5831),
    .B(_08486_));
 sg13g2_inv_1 _39077_ (.Y(_08489_),
    .A(_08488_));
 sg13g2_nor2_1 _39078_ (.A(_08481_),
    .B(_08489_),
    .Y(_08490_));
 sg13g2_nand2b_1 _39079_ (.Y(_08491_),
    .B(_04409_),
    .A_N(_04408_));
 sg13g2_nand3b_1 _39080_ (.B(_08491_),
    .C(net7406),
    .Y(_08492_),
    .A_N(_08150_));
 sg13g2_xnor2_1 _39081_ (.Y(_08493_),
    .A(_04409_),
    .B(_08140_));
 sg13g2_a21oi_1 _39082_ (.A1(net7239),
    .A2(\u_inv.d_next[96] ),
    .Y(_08494_),
    .B1(net6363));
 sg13g2_a22oi_1 _39083_ (.Y(_08495_),
    .B1(_08494_),
    .B2(_08492_),
    .A2(_08493_),
    .A1(net6363));
 sg13g2_and2_1 _39084_ (.A(net5830),
    .B(_08495_),
    .X(_08496_));
 sg13g2_xnor2_1 _39085_ (.Y(_08497_),
    .A(net5875),
    .B(_08495_));
 sg13g2_inv_1 _39086_ (.Y(_08498_),
    .A(_08497_));
 sg13g2_o21ai_1 _39087_ (.B1(_03924_),
    .Y(_08499_),
    .A1(_05117_),
    .A2(_08344_));
 sg13g2_nor3_1 _39088_ (.A(_03924_),
    .B(_05117_),
    .C(_08344_),
    .Y(_08500_));
 sg13g2_nor2_1 _39089_ (.A(net6270),
    .B(_08500_),
    .Y(_08501_));
 sg13g2_nor2_1 _39090_ (.A(_03924_),
    .B(_08150_),
    .Y(_08502_));
 sg13g2_o21ai_1 _39091_ (.B1(net7406),
    .Y(_08503_),
    .A1(_03923_),
    .A2(_03925_));
 sg13g2_a221oi_1 _39092_ (.B2(_03925_),
    .C1(_08503_),
    .B1(_08502_),
    .A1(_04408_),
    .Y(_08504_),
    .A2(_04410_));
 sg13g2_a21oi_1 _39093_ (.A1(net7239),
    .A2(\u_inv.d_next[97] ),
    .Y(_08505_),
    .B1(_08504_));
 sg13g2_a22oi_1 _39094_ (.Y(_08506_),
    .B1(_08505_),
    .B2(net6270),
    .A2(_08501_),
    .A1(_08499_));
 sg13g2_xnor2_1 _39095_ (.Y(_08507_),
    .A(net5831),
    .B(_08506_));
 sg13g2_nor2_1 _39096_ (.A(_08498_),
    .B(_08507_),
    .Y(_08508_));
 sg13g2_inv_1 _39097_ (.Y(_08509_),
    .A(_08508_));
 sg13g2_nand2_1 _39098_ (.Y(_08510_),
    .A(_08490_),
    .B(_08508_));
 sg13g2_nor3_2 _39099_ (.A(_08426_),
    .B(_08469_),
    .C(_08510_),
    .Y(_08511_));
 sg13g2_inv_1 _39100_ (.Y(_08512_),
    .A(_08511_));
 sg13g2_nand3b_1 _39101_ (.B(_08335_),
    .C(_08511_),
    .Y(_08513_),
    .A_N(_08240_));
 sg13g2_a21oi_2 _39102_ (.B1(_08513_),
    .Y(_08514_),
    .A2(net1097),
    .A1(_07358_));
 sg13g2_o21ai_1 _39103_ (.B1(_08466_),
    .Y(_08515_),
    .A1(net5875),
    .A2(_08459_));
 sg13g2_nand2_1 _39104_ (.Y(_08516_),
    .A(_08440_),
    .B(_08451_));
 sg13g2_a21oi_1 _39105_ (.A1(_08453_),
    .A2(_08515_),
    .Y(_08517_),
    .B1(_08516_));
 sg13g2_a21o_1 _39106_ (.A2(_08506_),
    .A1(net5831),
    .B1(_08496_),
    .X(_08518_));
 sg13g2_o21ai_1 _39107_ (.B1(_08487_),
    .Y(_08519_),
    .A1(net5874),
    .A2(_08480_));
 sg13g2_a21o_2 _39108_ (.A2(_08518_),
    .A1(_08490_),
    .B1(_08519_),
    .X(_08520_));
 sg13g2_a221oi_1 _39109_ (.B2(_08468_),
    .C1(_08516_),
    .B1(_08520_),
    .A1(_08453_),
    .Y(_08521_),
    .A2(_08515_));
 sg13g2_nand2_1 _39110_ (.Y(_08522_),
    .A(_08415_),
    .B(_08422_));
 sg13g2_nand2_1 _39111_ (.Y(_08523_),
    .A(_08393_),
    .B(_08404_));
 sg13g2_a21oi_1 _39112_ (.A1(net5832),
    .A2(_08369_),
    .Y(_08524_),
    .B1(_08376_));
 sg13g2_nor3_1 _39113_ (.A(_08353_),
    .B(_08362_),
    .C(_08524_),
    .Y(_08525_));
 sg13g2_o21ai_1 _39114_ (.B1(_08352_),
    .Y(_08526_),
    .A1(net5877),
    .A2(_08361_));
 sg13g2_or2_1 _39115_ (.X(_08527_),
    .B(_08526_),
    .A(_08525_));
 sg13g2_a221oi_1 _39116_ (.B2(_08425_),
    .C1(_08523_),
    .B1(_08527_),
    .A1(_08406_),
    .Y(_08528_),
    .A2(_08522_));
 sg13g2_o21ai_1 _39117_ (.B1(_08528_),
    .Y(_08529_),
    .A1(_08426_),
    .A2(_08521_));
 sg13g2_nand2_1 _39118_ (.Y(_08530_),
    .A(_08228_),
    .B(_08235_));
 sg13g2_o21ai_1 _39119_ (.B1(_08215_),
    .Y(_08531_),
    .A1(net5868),
    .A2(_08208_));
 sg13g2_a21o_2 _39120_ (.A2(_08530_),
    .A1(_08218_),
    .B1(_08531_),
    .X(_08532_));
 sg13g2_and2_1 _39121_ (.A(_08187_),
    .B(_08196_),
    .X(_08533_));
 sg13g2_nand2_1 _39122_ (.Y(_08534_),
    .A(_08187_),
    .B(_08196_));
 sg13g2_a21o_1 _39123_ (.A2(_08164_),
    .A1(net5818),
    .B1(_08174_),
    .X(_08535_));
 sg13g2_a221oi_1 _39124_ (.B2(_08177_),
    .C1(_08535_),
    .B1(_08534_),
    .A1(_08200_),
    .Y(_08536_),
    .A2(_08532_));
 sg13g2_o21ai_1 _39125_ (.B1(net5830),
    .Y(_08537_),
    .A1(_08324_),
    .A2(_08330_));
 sg13g2_nor3_1 _39126_ (.A(_08307_),
    .B(_08316_),
    .C(_08537_),
    .Y(_08538_));
 sg13g2_nor3_1 _39127_ (.A(_08305_),
    .B(_08315_),
    .C(_08538_),
    .Y(_08539_));
 sg13g2_or3_1 _39128_ (.A(_08305_),
    .B(_08315_),
    .C(_08538_),
    .X(_08540_));
 sg13g2_o21ai_1 _39129_ (.B1(_08283_),
    .Y(_08541_),
    .A1(net5869),
    .A2(_08292_));
 sg13g2_o21ai_1 _39130_ (.B1(_08256_),
    .Y(_08542_),
    .A1(net5868),
    .A2(_08267_));
 sg13g2_a221oi_1 _39131_ (.B2(_08271_),
    .C1(_08542_),
    .B1(_08541_),
    .A1(_08296_),
    .Y(_08543_),
    .A2(_08540_));
 sg13g2_o21ai_1 _39132_ (.B1(_08536_),
    .Y(_08544_),
    .A1(_08240_),
    .A2(_08543_));
 sg13g2_a21o_2 _39133_ (.A2(_08529_),
    .A1(_08336_),
    .B1(_08544_),
    .X(_08545_));
 sg13g2_nor2_1 _39134_ (.A(net1086),
    .B(_08545_),
    .Y(_08546_));
 sg13g2_xnor2_1 _39135_ (.Y(_08547_),
    .A(net5819),
    .B(_06784_));
 sg13g2_xnor2_1 _39136_ (.Y(_08548_),
    .A(net5866),
    .B(_06789_));
 sg13g2_nand3b_1 _39137_ (.B(_06776_),
    .C(_08548_),
    .Y(_08549_),
    .A_N(_06769_));
 sg13g2_nor2_1 _39138_ (.A(_08547_),
    .B(_08549_),
    .Y(_08550_));
 sg13g2_or2_1 _39139_ (.X(_08551_),
    .B(_08549_),
    .A(_08547_));
 sg13g2_or3_1 _39140_ (.A(_06730_),
    .B(_06739_),
    .C(_06759_),
    .X(_08552_));
 sg13g2_nor4_2 _39141_ (.A(_06864_),
    .B(_06892_),
    .C(_08551_),
    .Y(_08553_),
    .D(_08552_));
 sg13g2_nand2_2 _39142_ (.Y(_08554_),
    .A(_06715_),
    .B(_08553_));
 sg13g2_inv_1 _39143_ (.Y(_08555_),
    .A(_08554_));
 sg13g2_nor4_1 _39144_ (.A(_06348_),
    .B(_06442_),
    .C(_06947_),
    .D(_08554_),
    .Y(_08556_));
 sg13g2_o21ai_1 _39145_ (.B1(_08556_),
    .Y(_08557_),
    .A1(_08545_),
    .A2(net1086));
 sg13g2_xnor2_1 _39146_ (.Y(_08558_),
    .A(net5791),
    .B(_06078_));
 sg13g2_inv_1 _39147_ (.Y(_08559_),
    .A(_08558_));
 sg13g2_xnor2_1 _39148_ (.Y(_08560_),
    .A(net5842),
    .B(_06087_));
 sg13g2_or3_1 _39149_ (.A(_06072_),
    .B(_08559_),
    .C(_08560_),
    .X(_08561_));
 sg13g2_nor2_2 _39150_ (.A(_06050_),
    .B(_08561_),
    .Y(_08562_));
 sg13g2_inv_1 _39151_ (.Y(_08563_),
    .A(_08562_));
 sg13g2_nand2_1 _39152_ (.Y(_08564_),
    .A(_06010_),
    .B(_08562_));
 sg13g2_nand3b_1 _39153_ (.B(_06010_),
    .C(_08562_),
    .Y(_08565_),
    .A_N(_05915_));
 sg13g2_or2_1 _39154_ (.X(_08566_),
    .B(_08565_),
    .A(_05722_));
 sg13g2_a21o_2 _39155_ (.A2(net1077),
    .A1(_06950_),
    .B1(_08566_),
    .X(_08567_));
 sg13g2_xnor2_1 _39156_ (.Y(_08568_),
    .A(_03356_),
    .B(_04589_));
 sg13g2_a21o_1 _39157_ (.A2(_08568_),
    .A1(net7327),
    .B1(_04591_),
    .X(_08569_));
 sg13g2_nor3_1 _39158_ (.A(_03355_),
    .B(_05337_),
    .C(_05339_),
    .Y(_08570_));
 sg13g2_nand2_1 _39159_ (.Y(_08571_),
    .A(net6300),
    .B(_05340_));
 sg13g2_o21ai_1 _39160_ (.B1(_08569_),
    .Y(_08572_),
    .A1(_08570_),
    .A2(_08571_));
 sg13g2_inv_1 _39161_ (.Y(_08573_),
    .A(_08572_));
 sg13g2_xnor2_1 _39162_ (.Y(_08574_),
    .A(net5839),
    .B(_08572_));
 sg13g2_a21oi_2 _39163_ (.B1(_08574_),
    .Y(_08575_),
    .A2(_08567_),
    .A1(_06165_));
 sg13g2_a21oi_1 _39164_ (.A1(net6790),
    .A2(_08573_),
    .Y(_08576_),
    .B1(net5786));
 sg13g2_a21oi_2 _39165_ (.B1(_08576_),
    .Y(_08577_),
    .A2(_08575_),
    .A1(net6790));
 sg13g2_a21o_2 _39166_ (.A2(_08575_),
    .A1(net6790),
    .B1(_08576_),
    .X(_08578_));
 sg13g2_nand2_1 _39167_ (.Y(_08579_),
    .A(net5748),
    .B(net5580));
 sg13g2_xor2_1 _39168_ (.B(_05350_),
    .A(_03351_),
    .X(_08580_));
 sg13g2_nor2_1 _39169_ (.A(_03351_),
    .B(_08579_),
    .Y(_08581_));
 sg13g2_a21o_2 _39170_ (.A2(_08580_),
    .A1(_08579_),
    .B1(_08581_),
    .X(_08582_));
 sg13g2_a21oi_1 _39171_ (.A1(_08579_),
    .A2(_08580_),
    .Y(_08583_),
    .B1(_08581_));
 sg13g2_nor2_1 _39172_ (.A(net5739),
    .B(net5572),
    .Y(_08584_));
 sg13g2_a21oi_1 _39173_ (.A1(_06372_),
    .A2(_06377_),
    .Y(_08585_),
    .B1(net6798));
 sg13g2_o21ai_1 _39174_ (.B1(_08555_),
    .Y(_08586_),
    .A1(net1086),
    .A2(_08545_));
 sg13g2_nand2_1 _39175_ (.Y(_08587_),
    .A(_06911_),
    .B(_08586_));
 sg13g2_a21oi_2 _39176_ (.B1(_06348_),
    .Y(_08588_),
    .A2(_08586_),
    .A1(_06911_));
 sg13g2_nor2_1 _39177_ (.A(_06945_),
    .B(_08588_),
    .Y(_08589_));
 sg13g2_o21ai_1 _39178_ (.B1(_06946_),
    .Y(_08590_),
    .A1(_06945_),
    .A2(_08588_));
 sg13g2_and2_1 _39179_ (.A(_06919_),
    .B(_08590_),
    .X(_08591_));
 sg13g2_a21oi_1 _39180_ (.A1(_06919_),
    .A2(_08590_),
    .Y(_08592_),
    .B1(_06439_));
 sg13g2_a21oi_1 _39181_ (.A1(_06919_),
    .A2(_08590_),
    .Y(_08593_),
    .B1(_06441_));
 sg13g2_nor2_1 _39182_ (.A(_06923_),
    .B(_08593_),
    .Y(_08594_));
 sg13g2_o21ai_1 _39183_ (.B1(_06399_),
    .Y(_08595_),
    .A1(_06923_),
    .A2(_08593_));
 sg13g2_or2_1 _39184_ (.X(_08596_),
    .B(_08595_),
    .A(_06392_));
 sg13g2_a21oi_1 _39185_ (.A1(_06926_),
    .A2(_08596_),
    .Y(_08597_),
    .B1(_06369_));
 sg13g2_nor2_1 _39186_ (.A(_06368_),
    .B(_08597_),
    .Y(_08598_));
 sg13g2_xor2_1 _39187_ (.B(_08598_),
    .A(_06380_),
    .X(_08599_));
 sg13g2_a21oi_2 _39188_ (.B1(_08585_),
    .Y(_08600_),
    .A2(_08599_),
    .A1(net6799));
 sg13g2_and2_1 _39189_ (.A(net5627),
    .B(_08600_),
    .X(_08601_));
 sg13g2_xnor2_1 _39190_ (.Y(_08602_),
    .A(net5578),
    .B(_08600_));
 sg13g2_xnor2_1 _39191_ (.Y(_08603_),
    .A(net5628),
    .B(_08600_));
 sg13g2_nand3_1 _39192_ (.B(net1077),
    .C(_08559_),
    .A(_06950_),
    .Y(_08604_));
 sg13g2_a21o_2 _39193_ (.A2(net1077),
    .A1(_06950_),
    .B1(_08559_),
    .X(_08605_));
 sg13g2_a21oi_1 _39194_ (.A1(_08604_),
    .A2(_08605_),
    .Y(_08606_),
    .B1(net6755));
 sg13g2_a21o_2 _39195_ (.A2(_06078_),
    .A1(net6755),
    .B1(_08606_),
    .X(_08607_));
 sg13g2_inv_1 _39196_ (.Y(_08608_),
    .A(_08607_));
 sg13g2_nor2_1 _39197_ (.A(net5578),
    .B(_08607_),
    .Y(_08609_));
 sg13g2_xnor2_1 _39198_ (.Y(_08610_),
    .A(net5628),
    .B(_08607_));
 sg13g2_inv_1 _39199_ (.Y(_08611_),
    .A(_08610_));
 sg13g2_nor2_1 _39200_ (.A(net6798),
    .B(_06389_),
    .Y(_08612_));
 sg13g2_nand2b_1 _39201_ (.Y(_08613_),
    .B(_08595_),
    .A_N(_06398_));
 sg13g2_xor2_1 _39202_ (.B(_08613_),
    .A(_06392_),
    .X(_08614_));
 sg13g2_a21oi_2 _39203_ (.B1(_08612_),
    .Y(_08615_),
    .A2(_08614_),
    .A1(net6799));
 sg13g2_xnor2_1 _39204_ (.Y(_08616_),
    .A(net5627),
    .B(_08615_));
 sg13g2_nand2_1 _39205_ (.Y(_08617_),
    .A(net6756),
    .B(_06367_));
 sg13g2_nand3_1 _39206_ (.B(_06926_),
    .C(_08596_),
    .A(_06369_),
    .Y(_08618_));
 sg13g2_nand2b_1 _39207_ (.Y(_08619_),
    .B(_08618_),
    .A_N(_08597_));
 sg13g2_o21ai_1 _39208_ (.B1(_08617_),
    .Y(_08620_),
    .A1(net6756),
    .A2(_08619_));
 sg13g2_xnor2_1 _39209_ (.Y(_08621_),
    .A(net5578),
    .B(_08620_));
 sg13g2_nor2b_1 _39210_ (.A(_08616_),
    .B_N(_08621_),
    .Y(_08622_));
 sg13g2_inv_1 _39211_ (.Y(_08623_),
    .A(_08622_));
 sg13g2_nor2_1 _39212_ (.A(net6799),
    .B(_06410_),
    .Y(_08624_));
 sg13g2_o21ai_1 _39213_ (.B1(_06419_),
    .Y(_08625_),
    .A1(_06921_),
    .A2(_08592_));
 sg13g2_nand2_1 _39214_ (.Y(_08626_),
    .A(_06418_),
    .B(_08625_));
 sg13g2_xor2_1 _39215_ (.B(_08626_),
    .A(_06412_),
    .X(_08627_));
 sg13g2_a21oi_2 _39216_ (.B1(_08624_),
    .Y(_08628_),
    .A2(_08627_),
    .A1(net6799));
 sg13g2_nand2_1 _39217_ (.Y(_08629_),
    .A(net5629),
    .B(_08628_));
 sg13g2_xnor2_1 _39218_ (.Y(_08630_),
    .A(net5629),
    .B(_08628_));
 sg13g2_nand2_1 _39219_ (.Y(_08631_),
    .A(net6755),
    .B(_06397_));
 sg13g2_xnor2_1 _39220_ (.Y(_08632_),
    .A(_06399_),
    .B(_08594_));
 sg13g2_o21ai_1 _39221_ (.B1(_08631_),
    .Y(_08633_),
    .A1(net6755),
    .A2(_08632_));
 sg13g2_inv_1 _39222_ (.Y(_08634_),
    .A(_08633_));
 sg13g2_xnor2_1 _39223_ (.Y(_08635_),
    .A(net5629),
    .B(_08633_));
 sg13g2_inv_1 _39224_ (.Y(_08636_),
    .A(_08635_));
 sg13g2_nor2_1 _39225_ (.A(_08630_),
    .B(_08636_),
    .Y(_08637_));
 sg13g2_or3_1 _39226_ (.A(_06419_),
    .B(_06921_),
    .C(_08592_),
    .X(_08638_));
 sg13g2_a21oi_1 _39227_ (.A1(_08625_),
    .A2(_08638_),
    .Y(_08639_),
    .B1(net6763));
 sg13g2_a21o_2 _39228_ (.A2(_06417_),
    .A1(net6763),
    .B1(_08639_),
    .X(_08640_));
 sg13g2_xnor2_1 _39229_ (.Y(_08641_),
    .A(net5578),
    .B(_08640_));
 sg13g2_inv_1 _39230_ (.Y(_08642_),
    .A(_08641_));
 sg13g2_nor2_1 _39231_ (.A(net6798),
    .B(_06428_),
    .Y(_08643_));
 sg13g2_o21ai_1 _39232_ (.B1(_06436_),
    .Y(_08644_),
    .A1(_06437_),
    .A2(_08591_));
 sg13g2_xnor2_1 _39233_ (.Y(_08645_),
    .A(_06430_),
    .B(_08644_));
 sg13g2_a21oi_2 _39234_ (.B1(_08643_),
    .Y(_08646_),
    .A2(_08645_),
    .A1(net6798));
 sg13g2_nand2_1 _39235_ (.Y(_08647_),
    .A(net5628),
    .B(_08646_));
 sg13g2_xnor2_1 _39236_ (.Y(_08648_),
    .A(net5628),
    .B(_08646_));
 sg13g2_nor4_1 _39237_ (.A(_08630_),
    .B(_08636_),
    .C(_08641_),
    .D(_08648_),
    .Y(_08649_));
 sg13g2_nand4_1 _39238_ (.B(_08610_),
    .C(_08622_),
    .A(_08602_),
    .Y(_08650_),
    .D(_08649_));
 sg13g2_nand2_1 _39239_ (.Y(_08651_),
    .A(net6763),
    .B(_06435_));
 sg13g2_xor2_1 _39240_ (.B(_08591_),
    .A(_06438_),
    .X(_08652_));
 sg13g2_o21ai_1 _39241_ (.B1(_08651_),
    .Y(_08653_),
    .A1(net6763),
    .A2(_08652_));
 sg13g2_nand2_1 _39242_ (.Y(_08654_),
    .A(net5629),
    .B(_08653_));
 sg13g2_xnor2_1 _39243_ (.Y(_08655_),
    .A(net5579),
    .B(_08653_));
 sg13g2_inv_1 _39244_ (.Y(_08656_),
    .A(_08655_));
 sg13g2_nor2_1 _39245_ (.A(net6804),
    .B(_06457_),
    .Y(_08657_));
 sg13g2_o21ai_1 _39246_ (.B1(_06524_),
    .Y(_08658_),
    .A1(_06945_),
    .A2(_08588_));
 sg13g2_o21ai_1 _39247_ (.B1(_06916_),
    .Y(_08659_),
    .A1(_06506_),
    .A2(_08658_));
 sg13g2_nand2b_1 _39248_ (.Y(_08660_),
    .B(_08659_),
    .A_N(_06475_));
 sg13g2_a21oi_1 _39249_ (.A1(_06486_),
    .A2(_08659_),
    .Y(_08661_),
    .B1(_06918_));
 sg13g2_o21ai_1 _39250_ (.B1(_06465_),
    .Y(_08662_),
    .A1(_06466_),
    .A2(_08661_));
 sg13g2_xor2_1 _39251_ (.B(_08662_),
    .A(_06459_),
    .X(_08663_));
 sg13g2_a21oi_2 _39252_ (.B1(_08657_),
    .Y(_08664_),
    .A2(_08663_),
    .A1(net6804));
 sg13g2_nand2_1 _39253_ (.Y(_08665_),
    .A(net5629),
    .B(_08664_));
 sg13g2_xnor2_1 _39254_ (.Y(_08666_),
    .A(net5629),
    .B(_08664_));
 sg13g2_or2_1 _39255_ (.X(_08667_),
    .B(_08666_),
    .A(_08656_));
 sg13g2_o21ai_1 _39256_ (.B1(net6804),
    .Y(_08668_),
    .A1(_06466_),
    .A2(_08661_));
 sg13g2_a21oi_1 _39257_ (.A1(_06466_),
    .A2(_08661_),
    .Y(_08669_),
    .B1(_08668_));
 sg13g2_a21oi_2 _39258_ (.B1(_08669_),
    .Y(_08670_),
    .A2(_06464_),
    .A1(net6763));
 sg13g2_xnor2_1 _39259_ (.Y(_08671_),
    .A(net5579),
    .B(_08670_));
 sg13g2_inv_1 _39260_ (.Y(_08672_),
    .A(_08671_));
 sg13g2_nor2_1 _39261_ (.A(net6804),
    .B(_06483_),
    .Y(_08673_));
 sg13g2_nand2_1 _39262_ (.Y(_08674_),
    .A(_06474_),
    .B(_08660_));
 sg13g2_xor2_1 _39263_ (.B(_08674_),
    .A(_06485_),
    .X(_08675_));
 sg13g2_a21oi_2 _39264_ (.B1(_08673_),
    .Y(_08676_),
    .A2(_08675_),
    .A1(net6804));
 sg13g2_nand2_1 _39265_ (.Y(_08677_),
    .A(net5628),
    .B(_08676_));
 sg13g2_xnor2_1 _39266_ (.Y(_08678_),
    .A(net5638),
    .B(_08676_));
 sg13g2_nor2_1 _39267_ (.A(net6805),
    .B(_06503_),
    .Y(_08679_));
 sg13g2_a21o_1 _39268_ (.A2(_08658_),
    .A1(_06913_),
    .B1(_06495_),
    .X(_08680_));
 sg13g2_nand2_1 _39269_ (.Y(_08681_),
    .A(_06494_),
    .B(_08680_));
 sg13g2_xnor2_1 _39270_ (.Y(_08682_),
    .A(_06504_),
    .B(_08681_));
 sg13g2_a21oi_2 _39271_ (.B1(_08679_),
    .Y(_08683_),
    .A2(_08682_),
    .A1(net6805));
 sg13g2_and2_1 _39272_ (.A(net5639),
    .B(_08683_),
    .X(_08684_));
 sg13g2_xnor2_1 _39273_ (.Y(_08685_),
    .A(net5639),
    .B(_08683_));
 sg13g2_nor2_1 _39274_ (.A(net6804),
    .B(_06473_),
    .Y(_08686_));
 sg13g2_xor2_1 _39275_ (.B(_08659_),
    .A(_06475_),
    .X(_08687_));
 sg13g2_a21oi_2 _39276_ (.B1(_08686_),
    .Y(_08688_),
    .A2(_08687_),
    .A1(net6804));
 sg13g2_xnor2_1 _39277_ (.Y(_08689_),
    .A(net5639),
    .B(_08688_));
 sg13g2_nor2_1 _39278_ (.A(_08685_),
    .B(_08689_),
    .Y(_08690_));
 sg13g2_nand2_1 _39279_ (.Y(_08691_),
    .A(net6763),
    .B(_06493_));
 sg13g2_nand3_1 _39280_ (.B(_06913_),
    .C(_08658_),
    .A(_06495_),
    .Y(_08692_));
 sg13g2_nand3_1 _39281_ (.B(_08680_),
    .C(_08692_),
    .A(net6805),
    .Y(_08693_));
 sg13g2_nand2_2 _39282_ (.Y(_08694_),
    .A(_08691_),
    .B(_08693_));
 sg13g2_inv_1 _39283_ (.Y(_08695_),
    .A(_08694_));
 sg13g2_xnor2_1 _39284_ (.Y(_08696_),
    .A(net5581),
    .B(_08694_));
 sg13g2_o21ai_1 _39285_ (.B1(_06512_),
    .Y(_08697_),
    .A1(_06513_),
    .A2(_08589_));
 sg13g2_xnor2_1 _39286_ (.Y(_08698_),
    .A(_06523_),
    .B(_08697_));
 sg13g2_nor2_1 _39287_ (.A(net6805),
    .B(_06521_),
    .Y(_08699_));
 sg13g2_a21oi_2 _39288_ (.B1(_08699_),
    .Y(_08700_),
    .A2(_08698_),
    .A1(net6805));
 sg13g2_inv_1 _39289_ (.Y(_08701_),
    .A(_08700_));
 sg13g2_xnor2_1 _39290_ (.Y(_08702_),
    .A(net5638),
    .B(_08700_));
 sg13g2_nand3_1 _39291_ (.B(_08696_),
    .C(_08702_),
    .A(_08690_),
    .Y(_08703_));
 sg13g2_inv_1 _39292_ (.Y(_08704_),
    .A(_08703_));
 sg13g2_nor4_1 _39293_ (.A(_08667_),
    .B(_08671_),
    .C(_08678_),
    .D(_08703_),
    .Y(_08705_));
 sg13g2_inv_1 _39294_ (.Y(_08706_),
    .A(_08705_));
 sg13g2_a21oi_1 _39295_ (.A1(_06911_),
    .A2(_08586_),
    .Y(_08707_),
    .B1(_06258_));
 sg13g2_nor2_1 _39296_ (.A(_06936_),
    .B(_08707_),
    .Y(_08708_));
 sg13g2_nor2_1 _39297_ (.A(_06345_),
    .B(_08708_),
    .Y(_08709_));
 sg13g2_o21ai_1 _39298_ (.B1(_06346_),
    .Y(_08710_),
    .A1(_06936_),
    .A2(_08707_));
 sg13g2_o21ai_1 _39299_ (.B1(_06347_),
    .Y(_08711_),
    .A1(_06936_),
    .A2(_08707_));
 sg13g2_a21o_1 _39300_ (.A2(_08711_),
    .A1(_06943_),
    .B1(_06293_),
    .X(_08712_));
 sg13g2_a221oi_1 _39301_ (.B2(_08711_),
    .C1(_06293_),
    .B1(_06943_),
    .A1(_06303_),
    .Y(_08713_),
    .A2(_06304_));
 sg13g2_o21ai_1 _39302_ (.B1(_06275_),
    .Y(_08714_),
    .A1(_06938_),
    .A2(_08713_));
 sg13g2_nand3_1 _39303_ (.B(_06284_),
    .C(_08714_),
    .A(_06273_),
    .Y(_08715_));
 sg13g2_a21o_1 _39304_ (.A2(_08714_),
    .A1(_06273_),
    .B1(_06284_),
    .X(_08716_));
 sg13g2_a21oi_1 _39305_ (.A1(_08715_),
    .A2(_08716_),
    .Y(_08717_),
    .B1(net6761));
 sg13g2_a21oi_2 _39306_ (.B1(_08717_),
    .Y(_08718_),
    .A2(_06283_),
    .A1(net6761));
 sg13g2_nand2_1 _39307_ (.Y(_08719_),
    .A(net5636),
    .B(_08718_));
 sg13g2_xnor2_1 _39308_ (.Y(_08720_),
    .A(net5636),
    .B(_08718_));
 sg13g2_nand2_1 _39309_ (.Y(_08721_),
    .A(net6763),
    .B(_06511_));
 sg13g2_xnor2_1 _39310_ (.Y(_08722_),
    .A(_06513_),
    .B(_08589_));
 sg13g2_o21ai_1 _39311_ (.B1(_08721_),
    .Y(_08723_),
    .A1(net6763),
    .A2(_08722_));
 sg13g2_nand2_1 _39312_ (.Y(_08724_),
    .A(net5636),
    .B(_08723_));
 sg13g2_xnor2_1 _39313_ (.Y(_08725_),
    .A(net5636),
    .B(_08723_));
 sg13g2_nor2_1 _39314_ (.A(_08720_),
    .B(_08725_),
    .Y(_08726_));
 sg13g2_nand2_1 _39315_ (.Y(_08727_),
    .A(_06292_),
    .B(_08712_));
 sg13g2_nor2_1 _39316_ (.A(net6807),
    .B(_06301_),
    .Y(_08728_));
 sg13g2_xnor2_1 _39317_ (.Y(_08729_),
    .A(_06305_),
    .B(_08727_));
 sg13g2_a21oi_2 _39318_ (.B1(_08728_),
    .Y(_08730_),
    .A2(_08729_),
    .A1(net6808));
 sg13g2_xnor2_1 _39319_ (.Y(_08731_),
    .A(net5584),
    .B(_08730_));
 sg13g2_inv_1 _39320_ (.Y(_08732_),
    .A(_08731_));
 sg13g2_nand2_1 _39321_ (.Y(_08733_),
    .A(net6761),
    .B(_06272_));
 sg13g2_nor3_1 _39322_ (.A(_06275_),
    .B(_06938_),
    .C(_08713_),
    .Y(_08734_));
 sg13g2_nand2_1 _39323_ (.Y(_08735_),
    .A(net6804),
    .B(_08714_));
 sg13g2_o21ai_1 _39324_ (.B1(_08733_),
    .Y(_08736_),
    .A1(_08734_),
    .A2(_08735_));
 sg13g2_xnor2_1 _39325_ (.Y(_08737_),
    .A(net5584),
    .B(_08736_));
 sg13g2_nand2_1 _39326_ (.Y(_08738_),
    .A(_08731_),
    .B(_08737_));
 sg13g2_nor3_1 _39327_ (.A(_08720_),
    .B(_08725_),
    .C(_08738_),
    .Y(_08739_));
 sg13g2_nand2_1 _39328_ (.Y(_08740_),
    .A(net6761),
    .B(_06291_));
 sg13g2_nand3_1 _39329_ (.B(_06943_),
    .C(_08711_),
    .A(_06293_),
    .Y(_08741_));
 sg13g2_nand3_1 _39330_ (.B(_08712_),
    .C(_08741_),
    .A(net6807),
    .Y(_08742_));
 sg13g2_nand2_2 _39331_ (.Y(_08743_),
    .A(_08740_),
    .B(_08742_));
 sg13g2_xnor2_1 _39332_ (.Y(_08744_),
    .A(net5636),
    .B(_08743_));
 sg13g2_nand2_1 _39333_ (.Y(_08745_),
    .A(net6761),
    .B(_06317_));
 sg13g2_a21oi_1 _39334_ (.A1(_06941_),
    .A2(_08710_),
    .Y(_08746_),
    .B1(_06326_));
 sg13g2_nor2_1 _39335_ (.A(_06325_),
    .B(_08746_),
    .Y(_08747_));
 sg13g2_xnor2_1 _39336_ (.Y(_08748_),
    .A(_06318_),
    .B(_08747_));
 sg13g2_o21ai_1 _39337_ (.B1(_08745_),
    .Y(_08749_),
    .A1(net6761),
    .A2(_08748_));
 sg13g2_xnor2_1 _39338_ (.Y(_08750_),
    .A(net5637),
    .B(_08749_));
 sg13g2_nand3_1 _39339_ (.B(_06941_),
    .C(_08710_),
    .A(_06326_),
    .Y(_08751_));
 sg13g2_nand3b_1 _39340_ (.B(_08751_),
    .C(net6806),
    .Y(_08752_),
    .A_N(_08746_));
 sg13g2_o21ai_1 _39341_ (.B1(_08752_),
    .Y(_08753_),
    .A1(net6806),
    .A2(_06324_));
 sg13g2_inv_1 _39342_ (.Y(_08754_),
    .A(_08753_));
 sg13g2_xnor2_1 _39343_ (.Y(_08755_),
    .A(net5637),
    .B(_08753_));
 sg13g2_nor2_1 _39344_ (.A(net6806),
    .B(_06335_),
    .Y(_08756_));
 sg13g2_nor2_1 _39345_ (.A(_06344_),
    .B(_08709_),
    .Y(_08757_));
 sg13g2_xnor2_1 _39346_ (.Y(_08758_),
    .A(_06337_),
    .B(_08757_));
 sg13g2_a21oi_2 _39347_ (.B1(_08756_),
    .Y(_08759_),
    .A2(_08758_),
    .A1(net6806));
 sg13g2_xnor2_1 _39348_ (.Y(_08760_),
    .A(net5637),
    .B(_08759_));
 sg13g2_inv_1 _39349_ (.Y(_08761_),
    .A(_08760_));
 sg13g2_nor4_2 _39350_ (.A(_08744_),
    .B(_08750_),
    .C(_08755_),
    .Y(_08762_),
    .D(_08761_));
 sg13g2_nand2_1 _39351_ (.Y(_08763_),
    .A(_08739_),
    .B(_08762_));
 sg13g2_nand2_1 _39352_ (.Y(_08764_),
    .A(net6761),
    .B(_06343_));
 sg13g2_xnor2_1 _39353_ (.Y(_08765_),
    .A(_06345_),
    .B(_08708_));
 sg13g2_o21ai_1 _39354_ (.B1(_08764_),
    .Y(_08766_),
    .A1(net6761),
    .A2(_08765_));
 sg13g2_and2_1 _39355_ (.A(net5641),
    .B(_08766_),
    .X(_08767_));
 sg13g2_xnor2_1 _39356_ (.Y(_08768_),
    .A(net5641),
    .B(_08766_));
 sg13g2_nor2_1 _39357_ (.A(net6806),
    .B(_06193_),
    .Y(_08769_));
 sg13g2_a21oi_1 _39358_ (.A1(_06911_),
    .A2(_08586_),
    .Y(_08770_),
    .B1(_06221_));
 sg13g2_a21oi_2 _39359_ (.B1(_06931_),
    .Y(_08771_),
    .A2(_08770_),
    .A1(_06254_));
 sg13g2_nor2_1 _39360_ (.A(_06212_),
    .B(_08771_),
    .Y(_08772_));
 sg13g2_o21ai_1 _39361_ (.B1(_06211_),
    .Y(_08773_),
    .A1(_06212_),
    .A2(_08771_));
 sg13g2_a21oi_1 _39362_ (.A1(_06206_),
    .A2(_08772_),
    .Y(_08774_),
    .B1(_06934_));
 sg13g2_o21ai_1 _39363_ (.B1(_06184_),
    .Y(_08775_),
    .A1(_06185_),
    .A2(_08774_));
 sg13g2_xor2_1 _39364_ (.B(_08775_),
    .A(_06195_),
    .X(_08776_));
 sg13g2_a21oi_2 _39365_ (.B1(_08769_),
    .Y(_08777_),
    .A2(_08776_),
    .A1(net6806));
 sg13g2_and2_1 _39366_ (.A(net5641),
    .B(_08777_),
    .X(_08778_));
 sg13g2_xnor2_1 _39367_ (.Y(_08779_),
    .A(net5582),
    .B(_08777_));
 sg13g2_xnor2_1 _39368_ (.Y(_08780_),
    .A(net5641),
    .B(_08777_));
 sg13g2_nand2_1 _39369_ (.Y(_08781_),
    .A(net6762),
    .B(_06183_));
 sg13g2_xnor2_1 _39370_ (.Y(_08782_),
    .A(_06185_),
    .B(_08774_));
 sg13g2_o21ai_1 _39371_ (.B1(_08781_),
    .Y(_08783_),
    .A1(net6762),
    .A2(_08782_));
 sg13g2_inv_1 _39372_ (.Y(_08784_),
    .A(_08783_));
 sg13g2_xnor2_1 _39373_ (.Y(_08785_),
    .A(net5582),
    .B(_08783_));
 sg13g2_nor2_1 _39374_ (.A(net6806),
    .B(_06204_),
    .Y(_08786_));
 sg13g2_xnor2_1 _39375_ (.Y(_08787_),
    .A(_06206_),
    .B(_08773_));
 sg13g2_a21oi_2 _39376_ (.B1(_08786_),
    .Y(_08788_),
    .A2(_08787_),
    .A1(net6806));
 sg13g2_nand2_1 _39377_ (.Y(_08789_),
    .A(net5640),
    .B(_08788_));
 sg13g2_xnor2_1 _39378_ (.Y(_08790_),
    .A(net5582),
    .B(_08788_));
 sg13g2_nand2_1 _39379_ (.Y(_08791_),
    .A(_08785_),
    .B(_08790_));
 sg13g2_nand2_1 _39380_ (.Y(_08792_),
    .A(net6762),
    .B(_06210_));
 sg13g2_xnor2_1 _39381_ (.Y(_08793_),
    .A(_06212_),
    .B(_08771_));
 sg13g2_o21ai_1 _39382_ (.B1(_08792_),
    .Y(_08794_),
    .A1(net6762),
    .A2(_08793_));
 sg13g2_and2_1 _39383_ (.A(net5641),
    .B(_08794_),
    .X(_08795_));
 sg13g2_xnor2_1 _39384_ (.Y(_08796_),
    .A(net5640),
    .B(_08794_));
 sg13g2_nor2_1 _39385_ (.A(net6807),
    .B(_06240_),
    .Y(_08797_));
 sg13g2_a21oi_1 _39386_ (.A1(_06256_),
    .A2(_08587_),
    .Y(_08798_),
    .B1(_06929_));
 sg13g2_o21ai_1 _39387_ (.B1(_06230_),
    .Y(_08799_),
    .A1(_06232_),
    .A2(_08798_));
 sg13g2_xnor2_1 _39388_ (.Y(_08800_),
    .A(_06242_),
    .B(_08799_));
 sg13g2_a21oi_2 _39389_ (.B1(_08797_),
    .Y(_08801_),
    .A2(_08800_),
    .A1(net6807));
 sg13g2_and2_1 _39390_ (.A(net5640),
    .B(_08801_),
    .X(_08802_));
 sg13g2_xnor2_1 _39391_ (.Y(_08803_),
    .A(net5640),
    .B(_08801_));
 sg13g2_o21ai_1 _39392_ (.B1(net6807),
    .Y(_08804_),
    .A1(_06232_),
    .A2(_08798_));
 sg13g2_a21o_1 _39393_ (.A2(_08798_),
    .A1(_06232_),
    .B1(_08804_),
    .X(_08805_));
 sg13g2_o21ai_1 _39394_ (.B1(_08805_),
    .Y(_08806_),
    .A1(net6807),
    .A2(_06229_));
 sg13g2_inv_1 _39395_ (.Y(_08807_),
    .A(_08806_));
 sg13g2_nor2_1 _39396_ (.A(net6807),
    .B(_06252_),
    .Y(_08808_));
 sg13g2_nor2_1 _39397_ (.A(_06220_),
    .B(_08770_),
    .Y(_08809_));
 sg13g2_xnor2_1 _39398_ (.Y(_08810_),
    .A(_06253_),
    .B(_08809_));
 sg13g2_a21oi_2 _39399_ (.B1(_08808_),
    .Y(_08811_),
    .A2(_08810_),
    .A1(net6808));
 sg13g2_and2_1 _39400_ (.A(net5640),
    .B(_08811_),
    .X(_08812_));
 sg13g2_a21oi_1 _39401_ (.A1(net5640),
    .A2(_08806_),
    .Y(_08813_),
    .B1(_08812_));
 sg13g2_nor3_1 _39402_ (.A(_08796_),
    .B(_08803_),
    .C(_08813_),
    .Y(_08814_));
 sg13g2_nor3_1 _39403_ (.A(_08795_),
    .B(_08802_),
    .C(_08814_),
    .Y(_08815_));
 sg13g2_or3_1 _39404_ (.A(_08795_),
    .B(_08802_),
    .C(_08814_),
    .X(_08816_));
 sg13g2_nor4_1 _39405_ (.A(_08768_),
    .B(_08780_),
    .C(_08791_),
    .D(_08815_),
    .Y(_08817_));
 sg13g2_o21ai_1 _39406_ (.B1(net5641),
    .Y(_08818_),
    .A1(_08783_),
    .A2(_08788_));
 sg13g2_nor3_1 _39407_ (.A(_08768_),
    .B(_08780_),
    .C(_08818_),
    .Y(_08819_));
 sg13g2_nor4_1 _39408_ (.A(_08767_),
    .B(_08778_),
    .C(_08817_),
    .D(_08819_),
    .Y(_08820_));
 sg13g2_or4_1 _39409_ (.A(_08767_),
    .B(_08778_),
    .C(_08817_),
    .D(_08819_),
    .X(_08821_));
 sg13g2_a21o_1 _39410_ (.A2(_08759_),
    .A1(_08754_),
    .B1(net5581),
    .X(_08822_));
 sg13g2_nor3_1 _39411_ (.A(_08744_),
    .B(_08750_),
    .C(_08822_),
    .Y(_08823_));
 sg13g2_o21ai_1 _39412_ (.B1(net5636),
    .Y(_08824_),
    .A1(_08743_),
    .A2(_08749_));
 sg13g2_nor2b_1 _39413_ (.A(_08823_),
    .B_N(_08824_),
    .Y(_08825_));
 sg13g2_nand2b_1 _39414_ (.Y(_08826_),
    .B(_08824_),
    .A_N(_08823_));
 sg13g2_o21ai_1 _39415_ (.B1(net5636),
    .Y(_08827_),
    .A1(_08730_),
    .A2(_08736_));
 sg13g2_inv_1 _39416_ (.Y(_08828_),
    .A(_08827_));
 sg13g2_nand2_1 _39417_ (.Y(_08829_),
    .A(_08719_),
    .B(_08724_));
 sg13g2_a221oi_1 _39418_ (.B2(_08726_),
    .C1(_08829_),
    .B1(_08828_),
    .A1(_08739_),
    .Y(_08830_),
    .A2(_08826_));
 sg13g2_o21ai_1 _39419_ (.B1(_08830_),
    .Y(_08831_),
    .A1(_08763_),
    .A2(_08820_));
 sg13g2_nand3b_1 _39420_ (.B(_08705_),
    .C(_08831_),
    .Y(_08832_),
    .A_N(_08650_));
 sg13g2_o21ai_1 _39421_ (.B1(net5639),
    .Y(_08833_),
    .A1(_08694_),
    .A2(_08701_));
 sg13g2_a21oi_1 _39422_ (.A1(_08695_),
    .A2(_08700_),
    .Y(_08834_),
    .B1(net5581));
 sg13g2_a221oi_1 _39423_ (.B2(_08834_),
    .C1(_08684_),
    .B1(_08690_),
    .A1(net5639),
    .Y(_08835_),
    .A2(_08688_));
 sg13g2_nor4_1 _39424_ (.A(_08667_),
    .B(_08671_),
    .C(_08678_),
    .D(_08835_),
    .Y(_08836_));
 sg13g2_nand2_1 _39425_ (.Y(_08837_),
    .A(_08654_),
    .B(_08665_));
 sg13g2_o21ai_1 _39426_ (.B1(_08677_),
    .Y(_08838_),
    .A1(net5579),
    .A2(_08670_));
 sg13g2_nor2b_1 _39427_ (.A(_08667_),
    .B_N(_08838_),
    .Y(_08839_));
 sg13g2_nor3_1 _39428_ (.A(_08836_),
    .B(_08837_),
    .C(_08839_),
    .Y(_08840_));
 sg13g2_or2_1 _39429_ (.X(_08841_),
    .B(_08840_),
    .A(_08650_));
 sg13g2_o21ai_1 _39430_ (.B1(_08647_),
    .Y(_08842_),
    .A1(net5578),
    .A2(_08640_));
 sg13g2_a22oi_1 _39431_ (.Y(_08843_),
    .B1(_08637_),
    .B2(_08842_),
    .A2(_08634_),
    .A1(net5628));
 sg13g2_nand2_1 _39432_ (.Y(_08844_),
    .A(_08629_),
    .B(_08843_));
 sg13g2_nand4_1 _39433_ (.B(_08610_),
    .C(_08622_),
    .A(_08602_),
    .Y(_08845_),
    .D(_08844_));
 sg13g2_o21ai_1 _39434_ (.B1(net5627),
    .Y(_08846_),
    .A1(_08615_),
    .A2(_08620_));
 sg13g2_nor3_1 _39435_ (.A(_08603_),
    .B(_08611_),
    .C(_08846_),
    .Y(_08847_));
 sg13g2_nor3_1 _39436_ (.A(_08601_),
    .B(_08609_),
    .C(_08847_),
    .Y(_08848_));
 sg13g2_and4_1 _39437_ (.A(_08832_),
    .B(_08841_),
    .C(_08845_),
    .D(_08848_),
    .X(_08849_));
 sg13g2_xnor2_1 _39438_ (.Y(_08850_),
    .A(net5640),
    .B(_08811_));
 sg13g2_xnor2_1 _39439_ (.Y(_08851_),
    .A(net5640),
    .B(_08806_));
 sg13g2_nor4_1 _39440_ (.A(_08796_),
    .B(_08803_),
    .C(_08850_),
    .D(_08851_),
    .Y(_08852_));
 sg13g2_inv_1 _39441_ (.Y(_08853_),
    .A(_08852_));
 sg13g2_nor4_1 _39442_ (.A(_08768_),
    .B(_08780_),
    .C(_08791_),
    .D(_08853_),
    .Y(_08854_));
 sg13g2_inv_1 _39443_ (.Y(_08855_),
    .A(_08854_));
 sg13g2_nand3_1 _39444_ (.B(_08762_),
    .C(_08854_),
    .A(_08739_),
    .Y(_08856_));
 sg13g2_or3_1 _39445_ (.A(_08650_),
    .B(_08706_),
    .C(_08856_),
    .X(_08857_));
 sg13g2_a21oi_1 _39446_ (.A1(_07166_),
    .A2(_07171_),
    .Y(_08858_),
    .B1(net6828));
 sg13g2_a21oi_1 _39447_ (.A1(_07757_),
    .A2(_08128_),
    .Y(_08859_),
    .B1(_08133_));
 sg13g2_o21ai_1 _39448_ (.B1(_08134_),
    .Y(_08860_),
    .A1(_07758_),
    .A2(_08127_));
 sg13g2_a21oi_2 _39449_ (.B1(_07291_),
    .Y(_08861_),
    .A2(_08860_),
    .A1(_07330_));
 sg13g2_nor2_2 _39450_ (.A(_07287_),
    .B(_08861_),
    .Y(_08862_));
 sg13g2_o21ai_1 _39451_ (.B1(_07218_),
    .Y(_08863_),
    .A1(_07287_),
    .A2(_08861_));
 sg13g2_o21ai_1 _39452_ (.B1(_07339_),
    .Y(_08864_),
    .A1(_07239_),
    .A2(_08863_));
 sg13g2_a21oi_1 _39453_ (.A1(_07197_),
    .A2(_08864_),
    .Y(_08865_),
    .B1(_07334_));
 sg13g2_o21ai_1 _39454_ (.B1(_07162_),
    .Y(_08866_),
    .A1(_07163_),
    .A2(_08865_));
 sg13g2_xor2_1 _39455_ (.B(_08866_),
    .A(_07174_),
    .X(_08867_));
 sg13g2_a21oi_2 _39456_ (.B1(_08858_),
    .Y(_08868_),
    .A2(_08867_),
    .A1(net6828));
 sg13g2_and2_1 _39457_ (.A(net5679),
    .B(_08868_),
    .X(_08869_));
 sg13g2_xnor2_1 _39458_ (.Y(_08870_),
    .A(net5604),
    .B(_08868_));
 sg13g2_a21oi_1 _39459_ (.A1(_07757_),
    .A2(_08128_),
    .Y(_08871_),
    .B1(_08136_));
 sg13g2_a21o_1 _39460_ (.A2(_08128_),
    .A1(_07757_),
    .B1(_08136_),
    .X(_08872_));
 sg13g2_nor3_1 _39461_ (.A(_07127_),
    .B(_07343_),
    .C(_08871_),
    .Y(_08873_));
 sg13g2_a21oi_1 _39462_ (.A1(_07342_),
    .A2(_08872_),
    .Y(_08874_),
    .B1(_07128_));
 sg13g2_nor3_1 _39463_ (.A(net6778),
    .B(_08873_),
    .C(_08874_),
    .Y(_08875_));
 sg13g2_a21o_2 _39464_ (.A2(_07125_),
    .A1(net6778),
    .B1(_08875_),
    .X(_08876_));
 sg13g2_xnor2_1 _39465_ (.Y(_08877_),
    .A(net5679),
    .B(_08876_));
 sg13g2_inv_1 _39466_ (.Y(_08878_),
    .A(_08877_));
 sg13g2_and2_1 _39467_ (.A(_08870_),
    .B(_08878_),
    .X(_08879_));
 sg13g2_nand2_1 _39468_ (.Y(_08880_),
    .A(net6785),
    .B(_07193_));
 sg13g2_a21oi_1 _39469_ (.A1(_07184_),
    .A2(_08864_),
    .Y(_08881_),
    .B1(_07183_));
 sg13g2_xnor2_1 _39470_ (.Y(_08882_),
    .A(_07196_),
    .B(_08881_));
 sg13g2_o21ai_1 _39471_ (.B1(_08880_),
    .Y(_08883_),
    .A1(net6785),
    .A2(_08882_));
 sg13g2_nor2_1 _39472_ (.A(net5604),
    .B(_08883_),
    .Y(_08884_));
 sg13g2_xnor2_1 _39473_ (.Y(_08885_),
    .A(net5599),
    .B(_08883_));
 sg13g2_nand2_1 _39474_ (.Y(_08886_),
    .A(net6785),
    .B(_07161_));
 sg13g2_xnor2_1 _39475_ (.Y(_08887_),
    .A(_07163_),
    .B(_08865_));
 sg13g2_o21ai_1 _39476_ (.B1(_08886_),
    .Y(_08888_),
    .A1(net6785),
    .A2(_08887_));
 sg13g2_nand2_1 _39477_ (.Y(_08889_),
    .A(net5679),
    .B(_08888_));
 sg13g2_nand2b_1 _39478_ (.Y(_08890_),
    .B(net5604),
    .A_N(_08888_));
 sg13g2_inv_1 _39479_ (.Y(_08891_),
    .A(_08890_));
 sg13g2_xnor2_1 _39480_ (.Y(_08892_),
    .A(net5604),
    .B(_08888_));
 sg13g2_nor2b_1 _39481_ (.A(_08885_),
    .B_N(_08892_),
    .Y(_08893_));
 sg13g2_a21o_1 _39482_ (.A2(_08863_),
    .A1(_07336_),
    .B1(_07237_),
    .X(_08894_));
 sg13g2_nor2b_1 _39483_ (.A(_07236_),
    .B_N(_08894_),
    .Y(_08895_));
 sg13g2_xnor2_1 _39484_ (.Y(_08896_),
    .A(_07229_),
    .B(_08895_));
 sg13g2_mux2_1 _39485_ (.A0(_07228_),
    .A1(_08896_),
    .S(net6829),
    .X(_08897_));
 sg13g2_inv_1 _39486_ (.Y(_08898_),
    .A(_08897_));
 sg13g2_nor2_1 _39487_ (.A(net5599),
    .B(_08897_),
    .Y(_08899_));
 sg13g2_xnor2_1 _39488_ (.Y(_08900_),
    .A(net5599),
    .B(_08897_));
 sg13g2_inv_1 _39489_ (.Y(_08901_),
    .A(_08900_));
 sg13g2_nor2_1 _39490_ (.A(net6828),
    .B(_07182_),
    .Y(_08902_));
 sg13g2_xor2_1 _39491_ (.B(_08864_),
    .A(_07184_),
    .X(_08903_));
 sg13g2_a21oi_2 _39492_ (.B1(_08902_),
    .Y(_08904_),
    .A2(_08903_),
    .A1(net6828));
 sg13g2_xnor2_1 _39493_ (.Y(_08905_),
    .A(net5600),
    .B(_08904_));
 sg13g2_nand3_1 _39494_ (.B(_07336_),
    .C(_08863_),
    .A(_07237_),
    .Y(_08906_));
 sg13g2_nand3_1 _39495_ (.B(_08894_),
    .C(_08906_),
    .A(net6829),
    .Y(_08907_));
 sg13g2_o21ai_1 _39496_ (.B1(_08907_),
    .Y(_08908_),
    .A1(net6829),
    .A2(_07235_));
 sg13g2_nand2b_1 _39497_ (.Y(_08909_),
    .B(net5599),
    .A_N(_08908_));
 sg13g2_inv_1 _39498_ (.Y(_08910_),
    .A(_08909_));
 sg13g2_xnor2_1 _39499_ (.Y(_08911_),
    .A(net5673),
    .B(_08908_));
 sg13g2_nor2_1 _39500_ (.A(net6828),
    .B(_07208_),
    .Y(_08912_));
 sg13g2_o21ai_1 _39501_ (.B1(_07216_),
    .Y(_08913_),
    .A1(_07217_),
    .A2(_08862_));
 sg13g2_xor2_1 _39502_ (.B(_08913_),
    .A(_07209_),
    .X(_08914_));
 sg13g2_a21oi_2 _39503_ (.B1(_08912_),
    .Y(_08915_),
    .A2(_08914_),
    .A1(net6828));
 sg13g2_nand2_1 _39504_ (.Y(_08916_),
    .A(net5673),
    .B(_08915_));
 sg13g2_xnor2_1 _39505_ (.Y(_08917_),
    .A(net5673),
    .B(_08915_));
 sg13g2_inv_1 _39506_ (.Y(_08918_),
    .A(_08917_));
 sg13g2_nor4_1 _39507_ (.A(_08900_),
    .B(_08905_),
    .C(_08911_),
    .D(_08917_),
    .Y(_08919_));
 sg13g2_nand4_1 _39508_ (.B(_08878_),
    .C(_08893_),
    .A(_08870_),
    .Y(_08920_),
    .D(_08919_));
 sg13g2_a21oi_1 _39509_ (.A1(_07247_),
    .A2(_07255_),
    .Y(_08921_),
    .B1(net6829));
 sg13g2_o21ai_1 _39510_ (.B1(_07289_),
    .Y(_08922_),
    .A1(_07331_),
    .A2(_08859_));
 sg13g2_a22oi_1 _39511_ (.Y(_08923_),
    .B1(_07285_),
    .B2(_08922_),
    .A2(_07279_),
    .A1(net5872));
 sg13g2_a221oi_1 _39512_ (.B2(_08922_),
    .C1(_07267_),
    .B1(_07285_),
    .A1(net5872),
    .Y(_08924_),
    .A2(_07279_));
 sg13g2_nor2_1 _39513_ (.A(_07266_),
    .B(_08924_),
    .Y(_08925_));
 sg13g2_xor2_1 _39514_ (.B(_08925_),
    .A(_07258_),
    .X(_08926_));
 sg13g2_a21o_2 _39515_ (.A2(_08926_),
    .A1(net6829),
    .B1(_08921_),
    .X(_08927_));
 sg13g2_inv_1 _39516_ (.Y(_08928_),
    .A(_08927_));
 sg13g2_nor2_1 _39517_ (.A(net5600),
    .B(_08927_),
    .Y(_08929_));
 sg13g2_xnor2_1 _39518_ (.Y(_08930_),
    .A(net5600),
    .B(_08927_));
 sg13g2_inv_1 _39519_ (.Y(_08931_),
    .A(_08930_));
 sg13g2_o21ai_1 _39520_ (.B1(net6828),
    .Y(_08932_),
    .A1(_07217_),
    .A2(_08862_));
 sg13g2_a21o_1 _39521_ (.A2(_08862_),
    .A1(_07217_),
    .B1(_08932_),
    .X(_08933_));
 sg13g2_o21ai_1 _39522_ (.B1(_08933_),
    .Y(_08934_),
    .A1(net6828),
    .A2(_07214_));
 sg13g2_nand2_1 _39523_ (.Y(_08935_),
    .A(net5672),
    .B(_08934_));
 sg13g2_xnor2_1 _39524_ (.Y(_08936_),
    .A(net5672),
    .B(_08934_));
 sg13g2_nor2_1 _39525_ (.A(net6785),
    .B(_08924_),
    .Y(_08937_));
 sg13g2_o21ai_1 _39526_ (.B1(_08937_),
    .Y(_08938_),
    .A1(_07268_),
    .A2(_08923_));
 sg13g2_o21ai_1 _39527_ (.B1(_08938_),
    .Y(_08939_),
    .A1(net6829),
    .A2(_07265_));
 sg13g2_nor2_1 _39528_ (.A(net5672),
    .B(_08939_),
    .Y(_08940_));
 sg13g2_xnor2_1 _39529_ (.Y(_08941_),
    .A(net5672),
    .B(_08939_));
 sg13g2_nand2_1 _39530_ (.Y(_08942_),
    .A(net6785),
    .B(_07278_));
 sg13g2_o21ai_1 _39531_ (.B1(_08922_),
    .Y(_08943_),
    .A1(net5872),
    .A2(_07284_));
 sg13g2_xnor2_1 _39532_ (.Y(_08944_),
    .A(_07288_),
    .B(_08943_));
 sg13g2_o21ai_1 _39533_ (.B1(_08942_),
    .Y(_08945_),
    .A1(net6785),
    .A2(_08944_));
 sg13g2_nand2_1 _39534_ (.Y(_08946_),
    .A(net5672),
    .B(_08945_));
 sg13g2_xnor2_1 _39535_ (.Y(_08947_),
    .A(net5672),
    .B(_08945_));
 sg13g2_inv_1 _39536_ (.Y(_08948_),
    .A(_08947_));
 sg13g2_nor4_1 _39537_ (.A(_08930_),
    .B(_08936_),
    .C(_08941_),
    .D(_08947_),
    .Y(_08949_));
 sg13g2_o21ai_1 _39538_ (.B1(_07327_),
    .Y(_08950_),
    .A1(_08129_),
    .A2(_08132_));
 sg13g2_and3_1 _39539_ (.X(_08951_),
    .A(_07301_),
    .B(_08130_),
    .C(_08950_));
 sg13g2_o21ai_1 _39540_ (.B1(_07310_),
    .Y(_08952_),
    .A1(_07300_),
    .A2(_08951_));
 sg13g2_or3_1 _39541_ (.A(_07300_),
    .B(_07310_),
    .C(_08951_),
    .X(_08953_));
 sg13g2_a21oi_1 _39542_ (.A1(_08952_),
    .A2(_08953_),
    .Y(_08954_),
    .B1(net6783));
 sg13g2_a21oi_2 _39543_ (.B1(_08954_),
    .Y(_08955_),
    .A2(_07309_),
    .A1(net6783));
 sg13g2_nand2_1 _39544_ (.Y(_08956_),
    .A(net5674),
    .B(_08955_));
 sg13g2_xnor2_1 _39545_ (.Y(_08957_),
    .A(net5675),
    .B(_08955_));
 sg13g2_nor2_1 _39546_ (.A(net6830),
    .B(_07284_),
    .Y(_08958_));
 sg13g2_nand3b_1 _39547_ (.B(_07330_),
    .C(_08860_),
    .Y(_08959_),
    .A_N(_07289_));
 sg13g2_and2_1 _39548_ (.A(_08922_),
    .B(_08959_),
    .X(_08960_));
 sg13g2_a21oi_2 _39549_ (.B1(_08958_),
    .Y(_08961_),
    .A2(_08960_),
    .A1(net6830));
 sg13g2_nor2_1 _39550_ (.A(net5599),
    .B(_08961_),
    .Y(_08962_));
 sg13g2_xnor2_1 _39551_ (.Y(_08963_),
    .A(net5674),
    .B(_08961_));
 sg13g2_nand2b_1 _39552_ (.Y(_08964_),
    .B(_08963_),
    .A_N(_08957_));
 sg13g2_nor2_1 _39553_ (.A(net6832),
    .B(_07299_),
    .Y(_08965_));
 sg13g2_a21oi_1 _39554_ (.A1(_08130_),
    .A2(_08950_),
    .Y(_08966_),
    .B1(_07301_));
 sg13g2_nor3_1 _39555_ (.A(net6783),
    .B(_08951_),
    .C(_08966_),
    .Y(_08967_));
 sg13g2_or2_1 _39556_ (.X(_08968_),
    .B(_08967_),
    .A(_08965_));
 sg13g2_nand2_1 _39557_ (.Y(_08969_),
    .A(net5675),
    .B(_08968_));
 sg13g2_nor2_1 _39558_ (.A(net6832),
    .B(_07319_),
    .Y(_08970_));
 sg13g2_o21ai_1 _39559_ (.B1(_07326_),
    .Y(_08971_),
    .A1(_08129_),
    .A2(_08132_));
 sg13g2_xor2_1 _39560_ (.B(_08971_),
    .A(_08131_),
    .X(_08972_));
 sg13g2_a21oi_2 _39561_ (.B1(_08970_),
    .Y(_08973_),
    .A2(_08972_),
    .A1(net6832));
 sg13g2_and2_1 _39562_ (.A(net5675),
    .B(_08973_),
    .X(_08974_));
 sg13g2_o21ai_1 _39563_ (.B1(net5675),
    .Y(_08975_),
    .A1(_08968_),
    .A2(_08973_));
 sg13g2_a21oi_1 _39564_ (.A1(net5672),
    .A2(_08955_),
    .Y(_08976_),
    .B1(_08962_));
 sg13g2_o21ai_1 _39565_ (.B1(_08976_),
    .Y(_08977_),
    .A1(_08964_),
    .A2(_08975_));
 sg13g2_o21ai_1 _39566_ (.B1(net5672),
    .Y(_08978_),
    .A1(_08939_),
    .A2(_08945_));
 sg13g2_or3_1 _39567_ (.A(_08930_),
    .B(_08936_),
    .C(_08978_),
    .X(_08979_));
 sg13g2_nand3b_1 _39568_ (.B(_08935_),
    .C(_08979_),
    .Y(_08980_),
    .A_N(_08929_));
 sg13g2_a21o_2 _39569_ (.A2(_08977_),
    .A1(_08949_),
    .B1(_08980_),
    .X(_08981_));
 sg13g2_nand2b_1 _39570_ (.Y(_08982_),
    .B(_08981_),
    .A_N(_08920_));
 sg13g2_o21ai_1 _39571_ (.B1(net5673),
    .Y(_08983_),
    .A1(_08908_),
    .A2(_08915_));
 sg13g2_nor3_1 _39572_ (.A(_08900_),
    .B(_08905_),
    .C(_08983_),
    .Y(_08984_));
 sg13g2_a21oi_1 _39573_ (.A1(_08897_),
    .A2(_08904_),
    .Y(_08985_),
    .B1(net5600));
 sg13g2_nor2_1 _39574_ (.A(_08984_),
    .B(_08985_),
    .Y(_08986_));
 sg13g2_nand3b_1 _39575_ (.B(_08893_),
    .C(_08879_),
    .Y(_08987_),
    .A_N(_08986_));
 sg13g2_nand2b_1 _39576_ (.Y(_08988_),
    .B(_08889_),
    .A_N(_08884_));
 sg13g2_a221oi_1 _39577_ (.B2(_08988_),
    .C1(_08869_),
    .B1(_08879_),
    .A1(net5679),
    .Y(_08989_),
    .A2(_08876_));
 sg13g2_nand3_1 _39578_ (.B(_08987_),
    .C(_08989_),
    .A(_08982_),
    .Y(_08990_));
 sg13g2_nor2_1 _39579_ (.A(net6825),
    .B(_06975_),
    .Y(_08991_));
 sg13g2_o21ai_1 _39580_ (.B1(_07138_),
    .Y(_08992_),
    .A1(_07343_),
    .A2(_08871_));
 sg13g2_a21oi_2 _39581_ (.B1(_07140_),
    .Y(_08993_),
    .A2(_08872_),
    .A1(_07342_));
 sg13g2_nor2_1 _39582_ (.A(_07357_),
    .B(_08993_),
    .Y(_08994_));
 sg13g2_o21ai_1 _39583_ (.B1(_07045_),
    .Y(_08995_),
    .A1(_07357_),
    .A2(_08993_));
 sg13g2_nand2b_2 _39584_ (.Y(_08996_),
    .B(_08995_),
    .A_N(_07347_));
 sg13g2_nand2_1 _39585_ (.Y(_08997_),
    .A(_07002_),
    .B(_08996_));
 sg13g2_a21oi_1 _39586_ (.A1(_07003_),
    .A2(_08996_),
    .Y(_08998_),
    .B1(_07349_));
 sg13g2_o21ai_1 _39587_ (.B1(_06982_),
    .Y(_08999_),
    .A1(_06983_),
    .A2(_08998_));
 sg13g2_xor2_1 _39588_ (.B(_08999_),
    .A(_06976_),
    .X(_09000_));
 sg13g2_a21oi_2 _39589_ (.B1(_08991_),
    .Y(_09001_),
    .A2(_09000_),
    .A1(net6826));
 sg13g2_nand2_1 _39590_ (.Y(_09002_),
    .A(net5675),
    .B(_09001_));
 sg13g2_xnor2_1 _39591_ (.Y(_09003_),
    .A(net5675),
    .B(_09001_));
 sg13g2_xnor2_1 _39592_ (.Y(_09004_),
    .A(_08139_),
    .B(_08497_));
 sg13g2_nand2_1 _39593_ (.Y(_09005_),
    .A(net6831),
    .B(_09004_));
 sg13g2_o21ai_1 _39594_ (.B1(_09005_),
    .Y(_09006_),
    .A1(net6831),
    .A2(_08495_));
 sg13g2_xnor2_1 _39595_ (.Y(_09007_),
    .A(net5603),
    .B(_09006_));
 sg13g2_nor2_1 _39596_ (.A(_09003_),
    .B(_09007_),
    .Y(_09008_));
 sg13g2_nand2_1 _39597_ (.Y(_09009_),
    .A(net6780),
    .B(_06981_));
 sg13g2_xnor2_1 _39598_ (.Y(_09010_),
    .A(_06983_),
    .B(_08998_));
 sg13g2_o21ai_1 _39599_ (.B1(_09009_),
    .Y(_09011_),
    .A1(net6780),
    .A2(_09010_));
 sg13g2_nand2b_1 _39600_ (.Y(_09012_),
    .B(net5597),
    .A_N(_09011_));
 sg13g2_xnor2_1 _39601_ (.Y(_09013_),
    .A(net5597),
    .B(_09011_));
 sg13g2_inv_2 _39602_ (.Y(_09014_),
    .A(_09013_));
 sg13g2_nor2_1 _39603_ (.A(net6825),
    .B(_06993_),
    .Y(_09015_));
 sg13g2_nand2_1 _39604_ (.Y(_09016_),
    .A(_07001_),
    .B(_08997_));
 sg13g2_xor2_1 _39605_ (.B(_09016_),
    .A(_06995_),
    .X(_09017_));
 sg13g2_a21oi_2 _39606_ (.B1(_09015_),
    .Y(_09018_),
    .A2(_09017_),
    .A1(net6826));
 sg13g2_and2_1 _39607_ (.A(net5668),
    .B(_09018_),
    .X(_09019_));
 sg13g2_xnor2_1 _39608_ (.Y(_09020_),
    .A(net5667),
    .B(_09018_));
 sg13g2_nor4_2 _39609_ (.A(_09003_),
    .B(_09007_),
    .C(_09014_),
    .Y(_09021_),
    .D(_09020_));
 sg13g2_nor2_1 _39610_ (.A(net6825),
    .B(_07000_),
    .Y(_09022_));
 sg13g2_xnor2_1 _39611_ (.Y(_09023_),
    .A(_07002_),
    .B(_08996_));
 sg13g2_a21oi_2 _39612_ (.B1(_09022_),
    .Y(_09024_),
    .A2(_09023_),
    .A1(net6825));
 sg13g2_and2_1 _39613_ (.A(net5668),
    .B(_09024_),
    .X(_09025_));
 sg13g2_xnor2_1 _39614_ (.Y(_09026_),
    .A(net5667),
    .B(_09024_));
 sg13g2_and2_1 _39615_ (.A(net6779),
    .B(_07022_),
    .X(_09027_));
 sg13g2_o21ai_1 _39616_ (.B1(_07043_),
    .Y(_09028_),
    .A1(_07357_),
    .A2(_08993_));
 sg13g2_nand2_1 _39617_ (.Y(_09029_),
    .A(_07042_),
    .B(_09028_));
 sg13g2_a21o_1 _39618_ (.A2(_09028_),
    .A1(_07345_),
    .B1(_07034_),
    .X(_09030_));
 sg13g2_o21ai_1 _39619_ (.B1(_07011_),
    .Y(_09031_),
    .A1(_07013_),
    .A2(_09030_));
 sg13g2_xnor2_1 _39620_ (.Y(_09032_),
    .A(_07024_),
    .B(_09031_));
 sg13g2_a21oi_2 _39621_ (.B1(_09027_),
    .Y(_09033_),
    .A2(_09032_),
    .A1(net6825));
 sg13g2_and2_1 _39622_ (.A(net5667),
    .B(_09033_),
    .X(_09034_));
 sg13g2_xnor2_1 _39623_ (.Y(_09035_),
    .A(net5597),
    .B(_09033_));
 sg13g2_xnor2_1 _39624_ (.Y(_09036_),
    .A(net5667),
    .B(_09033_));
 sg13g2_nand2_1 _39625_ (.Y(_09037_),
    .A(net6779),
    .B(_07010_));
 sg13g2_xnor2_1 _39626_ (.Y(_09038_),
    .A(_07013_),
    .B(_09030_));
 sg13g2_o21ai_1 _39627_ (.B1(_09037_),
    .Y(_09039_),
    .A1(net6780),
    .A2(_09038_));
 sg13g2_nand2b_1 _39628_ (.Y(_09040_),
    .B(net5597),
    .A_N(_09039_));
 sg13g2_inv_1 _39629_ (.Y(_09041_),
    .A(_09040_));
 sg13g2_xnor2_1 _39630_ (.Y(_09042_),
    .A(net5667),
    .B(_09039_));
 sg13g2_nor2_1 _39631_ (.A(net6825),
    .B(_07032_),
    .Y(_09043_));
 sg13g2_xnor2_1 _39632_ (.Y(_09044_),
    .A(_07036_),
    .B(_09029_));
 sg13g2_a21oi_2 _39633_ (.B1(_09043_),
    .Y(_09045_),
    .A2(_09044_),
    .A1(net6825));
 sg13g2_nand2_1 _39634_ (.Y(_09046_),
    .A(net5667),
    .B(_09045_));
 sg13g2_xnor2_1 _39635_ (.Y(_09047_),
    .A(net5667),
    .B(_09045_));
 sg13g2_inv_1 _39636_ (.Y(_09048_),
    .A(_09047_));
 sg13g2_nor4_2 _39637_ (.A(_09026_),
    .B(_09036_),
    .C(_09042_),
    .Y(_09049_),
    .D(_09047_));
 sg13g2_nand2_1 _39638_ (.Y(_09050_),
    .A(_09021_),
    .B(_09049_));
 sg13g2_a21oi_1 _39639_ (.A1(_07354_),
    .A2(_08992_),
    .Y(_09051_),
    .B1(_07098_));
 sg13g2_a21oi_1 _39640_ (.A1(net5821),
    .A2(_07096_),
    .Y(_09052_),
    .B1(_09051_));
 sg13g2_a221oi_1 _39641_ (.B2(_08992_),
    .C1(_07098_),
    .B1(_07354_),
    .A1(_07090_),
    .Y(_09053_),
    .A2(_07091_));
 sg13g2_o21ai_1 _39642_ (.B1(_07064_),
    .Y(_09054_),
    .A1(_07355_),
    .A2(_09053_));
 sg13g2_nand3_1 _39643_ (.B(_07077_),
    .C(_09054_),
    .A(_07063_),
    .Y(_09055_));
 sg13g2_a21o_1 _39644_ (.A2(_09054_),
    .A1(_07063_),
    .B1(_07077_),
    .X(_09056_));
 sg13g2_a21oi_1 _39645_ (.A1(_09055_),
    .A2(_09056_),
    .Y(_09057_),
    .B1(net6778));
 sg13g2_a21oi_2 _39646_ (.B1(_09057_),
    .Y(_09058_),
    .A2(_07074_),
    .A1(net6778));
 sg13g2_nand2_1 _39647_ (.Y(_09059_),
    .A(net5671),
    .B(_09058_));
 sg13g2_xnor2_1 _39648_ (.Y(_09060_),
    .A(net5671),
    .B(_09058_));
 sg13g2_xnor2_1 _39649_ (.Y(_09061_),
    .A(_07043_),
    .B(_08994_));
 sg13g2_mux2_1 _39650_ (.A0(_07041_),
    .A1(_09061_),
    .S(net6825),
    .X(_09062_));
 sg13g2_nand2_1 _39651_ (.Y(_09063_),
    .A(net5671),
    .B(_09062_));
 sg13g2_xnor2_1 _39652_ (.Y(_09064_),
    .A(net5598),
    .B(_09062_));
 sg13g2_inv_1 _39653_ (.Y(_09065_),
    .A(_09064_));
 sg13g2_nor2_1 _39654_ (.A(_09060_),
    .B(_09065_),
    .Y(_09066_));
 sg13g2_nand2_1 _39655_ (.Y(_09067_),
    .A(net6778),
    .B(_07062_));
 sg13g2_nor3_1 _39656_ (.A(_07064_),
    .B(_07355_),
    .C(_09053_),
    .Y(_09068_));
 sg13g2_nand2_1 _39657_ (.Y(_09069_),
    .A(net6827),
    .B(_09054_));
 sg13g2_o21ai_1 _39658_ (.B1(_09067_),
    .Y(_09070_),
    .A1(_09068_),
    .A2(_09069_));
 sg13g2_and2_1 _39659_ (.A(net5671),
    .B(_09070_),
    .X(_09071_));
 sg13g2_nand2b_1 _39660_ (.Y(_09072_),
    .B(net5598),
    .A_N(_09070_));
 sg13g2_nand2b_1 _39661_ (.Y(_09073_),
    .B(_09072_),
    .A_N(_09071_));
 sg13g2_a21oi_1 _39662_ (.A1(_07082_),
    .A2(_07088_),
    .Y(_09074_),
    .B1(net6827));
 sg13g2_xnor2_1 _39663_ (.Y(_09075_),
    .A(_07092_),
    .B(_09052_));
 sg13g2_a21oi_2 _39664_ (.B1(_09074_),
    .Y(_09076_),
    .A2(_09075_),
    .A1(net6827));
 sg13g2_xnor2_1 _39665_ (.Y(_09077_),
    .A(net5671),
    .B(_09076_));
 sg13g2_nor4_1 _39666_ (.A(_09060_),
    .B(_09065_),
    .C(_09073_),
    .D(_09077_),
    .Y(_09078_));
 sg13g2_inv_1 _39667_ (.Y(_09079_),
    .A(_09078_));
 sg13g2_nand2_1 _39668_ (.Y(_09080_),
    .A(net6781),
    .B(_07096_));
 sg13g2_nand3_1 _39669_ (.B(_07354_),
    .C(_08992_),
    .A(_07098_),
    .Y(_09081_));
 sg13g2_nand2_1 _39670_ (.Y(_09082_),
    .A(net6827),
    .B(_09081_));
 sg13g2_o21ai_1 _39671_ (.B1(_09080_),
    .Y(_09083_),
    .A1(_09051_),
    .A2(_09082_));
 sg13g2_xnor2_1 _39672_ (.Y(_09084_),
    .A(net5599),
    .B(_09083_));
 sg13g2_nand2_1 _39673_ (.Y(_09085_),
    .A(net6778),
    .B(_07110_));
 sg13g2_nor2_1 _39674_ (.A(_07126_),
    .B(_08874_),
    .Y(_09086_));
 sg13g2_a21oi_1 _39675_ (.A1(_07137_),
    .A2(_08874_),
    .Y(_09087_),
    .B1(_07352_));
 sg13g2_o21ai_1 _39676_ (.B1(_07118_),
    .Y(_09088_),
    .A1(_07119_),
    .A2(_09087_));
 sg13g2_xnor2_1 _39677_ (.Y(_09089_),
    .A(_07111_),
    .B(_09088_));
 sg13g2_o21ai_1 _39678_ (.B1(_09085_),
    .Y(_09090_),
    .A1(net6778),
    .A2(_09089_));
 sg13g2_nor2_1 _39679_ (.A(net5599),
    .B(_09090_),
    .Y(_09091_));
 sg13g2_xnor2_1 _39680_ (.Y(_09092_),
    .A(net5674),
    .B(_09090_));
 sg13g2_and2_1 _39681_ (.A(_09084_),
    .B(_09092_),
    .X(_09093_));
 sg13g2_xor2_1 _39682_ (.B(_09087_),
    .A(_07119_),
    .X(_09094_));
 sg13g2_nor2_1 _39683_ (.A(net6781),
    .B(_09094_),
    .Y(_09095_));
 sg13g2_a21oi_2 _39684_ (.B1(_09095_),
    .Y(_09096_),
    .A2(_07117_),
    .A1(net6778));
 sg13g2_or2_1 _39685_ (.X(_09097_),
    .B(_09096_),
    .A(net5674));
 sg13g2_inv_1 _39686_ (.Y(_09098_),
    .A(_09097_));
 sg13g2_xnor2_1 _39687_ (.Y(_09099_),
    .A(net5674),
    .B(_09096_));
 sg13g2_xnor2_1 _39688_ (.Y(_09100_),
    .A(_07137_),
    .B(_09086_));
 sg13g2_mux2_1 _39689_ (.A0(_07136_),
    .A1(_09100_),
    .S(net6827),
    .X(_09101_));
 sg13g2_nand2_1 _39690_ (.Y(_09102_),
    .A(net5674),
    .B(_09101_));
 sg13g2_xnor2_1 _39691_ (.Y(_09103_),
    .A(net5599),
    .B(_09101_));
 sg13g2_nand2_1 _39692_ (.Y(_09104_),
    .A(_09093_),
    .B(_09103_));
 sg13g2_nor2_1 _39693_ (.A(_09099_),
    .B(_09104_),
    .Y(_09105_));
 sg13g2_nor4_1 _39694_ (.A(_09050_),
    .B(_09079_),
    .C(_09099_),
    .D(_09104_),
    .Y(_09106_));
 sg13g2_o21ai_1 _39695_ (.B1(net5667),
    .Y(_09107_),
    .A1(_09039_),
    .A2(_09045_));
 sg13g2_nor3_1 _39696_ (.A(_09026_),
    .B(_09036_),
    .C(_09107_),
    .Y(_09108_));
 sg13g2_nor3_1 _39697_ (.A(_09025_),
    .B(_09034_),
    .C(_09108_),
    .Y(_09109_));
 sg13g2_or3_1 _39698_ (.A(_09025_),
    .B(_09034_),
    .C(_09108_),
    .X(_09110_));
 sg13g2_a21o_1 _39699_ (.A2(_09011_),
    .A1(net5675),
    .B1(_09019_),
    .X(_09111_));
 sg13g2_o21ai_1 _39700_ (.B1(_09002_),
    .Y(_09112_),
    .A1(net5603),
    .A2(_09006_));
 sg13g2_a221oi_1 _39701_ (.B2(_09008_),
    .C1(_09112_),
    .B1(_09111_),
    .A1(_09021_),
    .Y(_09113_),
    .A2(_09110_));
 sg13g2_a21o_1 _39702_ (.A2(_09076_),
    .A1(net5671),
    .B1(_09071_),
    .X(_09114_));
 sg13g2_nand2_1 _39703_ (.Y(_09115_),
    .A(_09059_),
    .B(_09063_));
 sg13g2_a21o_2 _39704_ (.A2(_09114_),
    .A1(_09066_),
    .B1(_09115_),
    .X(_09116_));
 sg13g2_o21ai_1 _39705_ (.B1(net5674),
    .Y(_09117_),
    .A1(_09096_),
    .A2(_09101_));
 sg13g2_inv_1 _39706_ (.Y(_09118_),
    .A(_09117_));
 sg13g2_a221oi_1 _39707_ (.B2(_09118_),
    .C1(_09091_),
    .B1(_09093_),
    .A1(net5674),
    .Y(_09119_),
    .A2(_09083_));
 sg13g2_inv_1 _39708_ (.Y(_09120_),
    .A(_09119_));
 sg13g2_a21oi_1 _39709_ (.A1(_09078_),
    .A2(_09120_),
    .Y(_09121_),
    .B1(_09116_));
 sg13g2_o21ai_1 _39710_ (.B1(_09113_),
    .Y(_09122_),
    .A1(_09050_),
    .A2(_09121_));
 sg13g2_nand4_1 _39711_ (.B(_09049_),
    .C(_09078_),
    .A(_09021_),
    .Y(_09123_),
    .D(_09105_));
 sg13g2_a21oi_2 _39712_ (.B1(_09122_),
    .Y(_09124_),
    .A2(_09106_),
    .A1(_08990_));
 sg13g2_nor2_1 _39713_ (.A(net6802),
    .B(_08051_),
    .Y(_09125_));
 sg13g2_nand2_1 _39714_ (.Y(_09126_),
    .A(_08014_),
    .B(_08053_));
 sg13g2_xor2_1 _39715_ (.B(_08053_),
    .A(_08014_),
    .X(_09127_));
 sg13g2_a21oi_2 _39716_ (.B1(_09125_),
    .Y(_09128_),
    .A2(_09127_),
    .A1(net6802));
 sg13g2_inv_1 _39717_ (.Y(_09129_),
    .A(_09128_));
 sg13g2_xnor2_1 _39718_ (.Y(_09130_),
    .A(net5622),
    .B(_09128_));
 sg13g2_nand2_1 _39719_ (.Y(_09131_),
    .A(net6760),
    .B(_07969_));
 sg13g2_nor2b_1 _39720_ (.A(_08011_),
    .B_N(_07961_),
    .Y(_09132_));
 sg13g2_a21o_1 _39721_ (.A2(_07960_),
    .A1(net5845),
    .B1(_09132_),
    .X(_09133_));
 sg13g2_xor2_1 _39722_ (.B(_09133_),
    .A(_07971_),
    .X(_09134_));
 sg13g2_o21ai_1 _39723_ (.B1(_09131_),
    .Y(_09135_),
    .A1(net6760),
    .A2(_09134_));
 sg13g2_nor2_1 _39724_ (.A(net5622),
    .B(_09135_),
    .Y(_09136_));
 sg13g2_xnor2_1 _39725_ (.Y(_09137_),
    .A(net5622),
    .B(_09135_));
 sg13g2_nor2_1 _39726_ (.A(_09130_),
    .B(_09137_),
    .Y(_09138_));
 sg13g2_xor2_1 _39727_ (.B(_08011_),
    .A(_07961_),
    .X(_09139_));
 sg13g2_nor2_1 _39728_ (.A(net6757),
    .B(_09139_),
    .Y(_09140_));
 sg13g2_a21oi_2 _39729_ (.B1(_09140_),
    .Y(_09141_),
    .A2(_07960_),
    .A1(net6760));
 sg13g2_nand2_1 _39730_ (.Y(_09142_),
    .A(net5580),
    .B(_09141_));
 sg13g2_xnor2_1 _39731_ (.Y(_09143_),
    .A(net5580),
    .B(_09141_));
 sg13g2_or2_1 _39732_ (.X(_09144_),
    .B(_07990_),
    .A(_07988_));
 sg13g2_a21oi_1 _39733_ (.A1(_07995_),
    .A2(_09144_),
    .Y(_09145_),
    .B1(net6757));
 sg13g2_o21ai_1 _39734_ (.B1(_09145_),
    .Y(_09146_),
    .A1(_07988_),
    .A2(_07996_));
 sg13g2_o21ai_1 _39735_ (.B1(_09146_),
    .Y(_09147_),
    .A1(net6801),
    .A2(_07986_));
 sg13g2_nand2_1 _39736_ (.Y(_09148_),
    .A(net5748),
    .B(_09147_));
 sg13g2_nor2_1 _39737_ (.A(_03351_),
    .B(_09148_),
    .Y(_09149_));
 sg13g2_nand2_1 _39738_ (.Y(_09150_),
    .A(net5699),
    .B(_08580_));
 sg13g2_o21ai_1 _39739_ (.B1(_09150_),
    .Y(_09151_),
    .A1(net5622),
    .A2(_09149_));
 sg13g2_xnor2_1 _39740_ (.Y(_09152_),
    .A(_07997_),
    .B(_08007_));
 sg13g2_nand2_1 _39741_ (.Y(_09153_),
    .A(net6801),
    .B(_09152_));
 sg13g2_o21ai_1 _39742_ (.B1(_09153_),
    .Y(_09154_),
    .A1(net6801),
    .A2(_08003_));
 sg13g2_xnor2_1 _39743_ (.Y(_09155_),
    .A(net5580),
    .B(_09154_));
 sg13g2_xnor2_1 _39744_ (.Y(_09156_),
    .A(net5622),
    .B(_09154_));
 sg13g2_nand2b_1 _39745_ (.Y(_09157_),
    .B(_09155_),
    .A_N(_09151_));
 sg13g2_nand2_1 _39746_ (.Y(_09158_),
    .A(net5622),
    .B(_09147_));
 sg13g2_o21ai_1 _39747_ (.B1(net5622),
    .Y(_09159_),
    .A1(_09147_),
    .A2(_09154_));
 sg13g2_o21ai_1 _39748_ (.B1(_09159_),
    .Y(_09160_),
    .A1(_09151_),
    .A2(_09156_));
 sg13g2_nor2_1 _39749_ (.A(_08006_),
    .B(_08008_),
    .Y(_09161_));
 sg13g2_xor2_1 _39750_ (.B(_09161_),
    .A(_07980_),
    .X(_09162_));
 sg13g2_mux2_1 _39751_ (.A0(_07979_),
    .A1(_09162_),
    .S(net6801),
    .X(_09163_));
 sg13g2_nor2_1 _39752_ (.A(net5622),
    .B(_09163_),
    .Y(_09164_));
 sg13g2_xnor2_1 _39753_ (.Y(_09165_),
    .A(net5580),
    .B(_09163_));
 sg13g2_a21oi_1 _39754_ (.A1(_09157_),
    .A2(_09159_),
    .Y(_09166_),
    .B1(_09165_));
 sg13g2_nor4_1 _39755_ (.A(_09130_),
    .B(_09137_),
    .C(_09143_),
    .D(_09165_),
    .Y(_09167_));
 sg13g2_a21oi_1 _39756_ (.A1(_09128_),
    .A2(_09135_),
    .Y(_09168_),
    .B1(net5630));
 sg13g2_nor2_1 _39757_ (.A(_09141_),
    .B(_09164_),
    .Y(_09169_));
 sg13g2_a22oi_1 _39758_ (.Y(_09170_),
    .B1(_09169_),
    .B2(_09138_),
    .A2(_09167_),
    .A1(_09160_));
 sg13g2_a221oi_1 _39759_ (.B2(_09138_),
    .C1(_09168_),
    .B1(_09169_),
    .A1(_09160_),
    .Y(_09171_),
    .A2(_09167_));
 sg13g2_nand2b_2 _39760_ (.Y(_09172_),
    .B(_09170_),
    .A_N(_09168_));
 sg13g2_nand2b_1 _39761_ (.Y(_09173_),
    .B(_08110_),
    .A_N(_08113_));
 sg13g2_nor2b_1 _39762_ (.A(_08110_),
    .B_N(_08113_),
    .Y(_09174_));
 sg13g2_nand3b_1 _39763_ (.B(net6803),
    .C(_09173_),
    .Y(_09175_),
    .A_N(_09174_));
 sg13g2_o21ai_1 _39764_ (.B1(_09175_),
    .Y(_09176_),
    .A1(net6803),
    .A2(_07942_));
 sg13g2_nand2_1 _39765_ (.Y(_09177_),
    .A(net5633),
    .B(_09176_));
 sg13g2_xnor2_1 _39766_ (.Y(_09178_),
    .A(net5631),
    .B(_09176_));
 sg13g2_nand2_1 _39767_ (.Y(_09179_),
    .A(net6759),
    .B(_08070_));
 sg13g2_o21ai_1 _39768_ (.B1(_08089_),
    .Y(_09180_),
    .A1(_08055_),
    .A2(_08107_));
 sg13g2_nand2_1 _39769_ (.Y(_09181_),
    .A(_08103_),
    .B(_09180_));
 sg13g2_and3_1 _39770_ (.X(_09182_),
    .A(_08080_),
    .B(_08098_),
    .C(_09181_));
 sg13g2_nor2_1 _39771_ (.A(_08079_),
    .B(_09182_),
    .Y(_09183_));
 sg13g2_xor2_1 _39772_ (.B(_09183_),
    .A(_08071_),
    .X(_09184_));
 sg13g2_o21ai_1 _39773_ (.B1(_09179_),
    .Y(_09185_),
    .A1(net6759),
    .A2(_09184_));
 sg13g2_inv_2 _39774_ (.Y(_09186_),
    .A(_09185_));
 sg13g2_nand2_1 _39775_ (.Y(_09187_),
    .A(net5631),
    .B(_09186_));
 sg13g2_xnor2_1 _39776_ (.Y(_09188_),
    .A(net5631),
    .B(_09186_));
 sg13g2_nor2_1 _39777_ (.A(_09178_),
    .B(_09188_),
    .Y(_09189_));
 sg13g2_nand2_1 _39778_ (.Y(_09190_),
    .A(_08088_),
    .B(_09180_));
 sg13g2_xor2_1 _39779_ (.B(_09190_),
    .A(_08099_),
    .X(_09191_));
 sg13g2_mux2_1 _39780_ (.A0(_08096_),
    .A1(_09191_),
    .S(net6802),
    .X(_09192_));
 sg13g2_nand2_1 _39781_ (.Y(_09193_),
    .A(net5631),
    .B(_09192_));
 sg13g2_xnor2_1 _39782_ (.Y(_09194_),
    .A(net5631),
    .B(_09192_));
 sg13g2_nor2_1 _39783_ (.A(net6803),
    .B(_08077_),
    .Y(_09195_));
 sg13g2_a21oi_1 _39784_ (.A1(_08098_),
    .A2(_09181_),
    .Y(_09196_),
    .B1(_08080_));
 sg13g2_nor3_1 _39785_ (.A(net6759),
    .B(_09182_),
    .C(_09196_),
    .Y(_09197_));
 sg13g2_nor2_2 _39786_ (.A(_09195_),
    .B(_09197_),
    .Y(_09198_));
 sg13g2_inv_1 _39787_ (.Y(_09199_),
    .A(_09198_));
 sg13g2_nand2_1 _39788_ (.Y(_09200_),
    .A(net5631),
    .B(_09199_));
 sg13g2_xnor2_1 _39789_ (.Y(_09201_),
    .A(net5585),
    .B(_09198_));
 sg13g2_nor4_1 _39790_ (.A(_09178_),
    .B(_09188_),
    .C(_09194_),
    .D(_09201_),
    .Y(_09202_));
 sg13g2_a21oi_1 _39791_ (.A1(_08014_),
    .A2(_08053_),
    .Y(_09203_),
    .B1(_08105_));
 sg13g2_nor2_1 _39792_ (.A(_08045_),
    .B(_09203_),
    .Y(_09204_));
 sg13g2_nor3_1 _39793_ (.A(_08025_),
    .B(_08045_),
    .C(_09203_),
    .Y(_09205_));
 sg13g2_nor2_1 _39794_ (.A(_08024_),
    .B(_09205_),
    .Y(_09206_));
 sg13g2_xor2_1 _39795_ (.B(_09206_),
    .A(_08034_),
    .X(_09207_));
 sg13g2_nor2_1 _39796_ (.A(net6760),
    .B(_09207_),
    .Y(_09208_));
 sg13g2_a21oi_2 _39797_ (.B1(_09208_),
    .Y(_09209_),
    .A2(_08033_),
    .A1(net6760));
 sg13g2_nand2_1 _39798_ (.Y(_09210_),
    .A(net5631),
    .B(_09209_));
 sg13g2_xnor2_1 _39799_ (.Y(_09211_),
    .A(net5585),
    .B(_09209_));
 sg13g2_or2_1 _39800_ (.X(_09212_),
    .B(_08087_),
    .A(net6802));
 sg13g2_nor3_1 _39801_ (.A(_08055_),
    .B(_08089_),
    .C(_08107_),
    .Y(_09213_));
 sg13g2_nand2_1 _39802_ (.Y(_09214_),
    .A(net6802),
    .B(_09180_));
 sg13g2_o21ai_1 _39803_ (.B1(_09212_),
    .Y(_09215_),
    .A1(_09213_),
    .A2(_09214_));
 sg13g2_nand2_1 _39804_ (.Y(_09216_),
    .A(net5631),
    .B(_09215_));
 sg13g2_xnor2_1 _39805_ (.Y(_09217_),
    .A(net5585),
    .B(_09215_));
 sg13g2_nor2_1 _39806_ (.A(net6802),
    .B(_08023_),
    .Y(_09218_));
 sg13g2_xnor2_1 _39807_ (.Y(_09219_),
    .A(_08025_),
    .B(_09204_));
 sg13g2_a21oi_2 _39808_ (.B1(_09218_),
    .Y(_09220_),
    .A2(_09219_),
    .A1(net6802));
 sg13g2_inv_1 _39809_ (.Y(_09221_),
    .A(_09220_));
 sg13g2_nor2_1 _39810_ (.A(net5632),
    .B(_09220_),
    .Y(_09222_));
 sg13g2_xnor2_1 _39811_ (.Y(_09223_),
    .A(net5585),
    .B(_09220_));
 sg13g2_nand2_1 _39812_ (.Y(_09224_),
    .A(_08052_),
    .B(_09126_));
 sg13g2_xnor2_1 _39813_ (.Y(_09225_),
    .A(_08046_),
    .B(_09224_));
 sg13g2_nand2_1 _39814_ (.Y(_09226_),
    .A(net6802),
    .B(_09225_));
 sg13g2_o21ai_1 _39815_ (.B1(_09226_),
    .Y(_09227_),
    .A1(net6803),
    .A2(_08043_));
 sg13g2_inv_2 _39816_ (.Y(_09228_),
    .A(_09227_));
 sg13g2_nor2_1 _39817_ (.A(net5632),
    .B(_09227_),
    .Y(_09229_));
 sg13g2_xnor2_1 _39818_ (.Y(_09230_),
    .A(net5632),
    .B(_09228_));
 sg13g2_and4_1 _39819_ (.A(_09211_),
    .B(_09217_),
    .C(_09223_),
    .D(_09230_),
    .X(_09231_));
 sg13g2_nand3b_1 _39820_ (.B(_09202_),
    .C(_09231_),
    .Y(_09232_),
    .A_N(_09171_));
 sg13g2_a21oi_1 _39821_ (.A1(_09220_),
    .A2(_09227_),
    .Y(_09233_),
    .B1(net5632));
 sg13g2_nand3_1 _39822_ (.B(_09217_),
    .C(_09233_),
    .A(_09211_),
    .Y(_09234_));
 sg13g2_nand3_1 _39823_ (.B(_09216_),
    .C(_09234_),
    .A(_09210_),
    .Y(_09235_));
 sg13g2_nand2_1 _39824_ (.Y(_09236_),
    .A(_09193_),
    .B(_09200_));
 sg13g2_nand2_1 _39825_ (.Y(_09237_),
    .A(_09177_),
    .B(_09187_));
 sg13g2_a221oi_1 _39826_ (.B2(_09189_),
    .C1(_09237_),
    .B1(_09236_),
    .A1(_09202_),
    .Y(_09238_),
    .A2(_09235_));
 sg13g2_nand2_1 _39827_ (.Y(_09239_),
    .A(_09232_),
    .B(_09238_));
 sg13g2_o21ai_1 _39828_ (.B1(_07951_),
    .Y(_09240_),
    .A1(_08110_),
    .A2(_08116_));
 sg13g2_nand3_1 _39829_ (.B(_07857_),
    .C(_09240_),
    .A(_07856_),
    .Y(_09241_));
 sg13g2_nand2_1 _39830_ (.Y(_09242_),
    .A(_07806_),
    .B(_09241_));
 sg13g2_a21oi_1 _39831_ (.A1(_07845_),
    .A2(_09242_),
    .Y(_09243_),
    .B1(_07844_));
 sg13g2_xor2_1 _39832_ (.B(_09243_),
    .A(_07836_),
    .X(_09244_));
 sg13g2_nor2_1 _39833_ (.A(net6809),
    .B(_07835_),
    .Y(_09245_));
 sg13g2_a21oi_2 _39834_ (.B1(_09245_),
    .Y(_09246_),
    .A2(_09244_),
    .A1(net6809));
 sg13g2_nand2b_1 _39835_ (.Y(_09247_),
    .B(net5644),
    .A_N(_09246_));
 sg13g2_xnor2_1 _39836_ (.Y(_09248_),
    .A(net5644),
    .B(_09246_));
 sg13g2_xnor2_1 _39837_ (.Y(_09249_),
    .A(net5586),
    .B(_09246_));
 sg13g2_nand2_1 _39838_ (.Y(_09250_),
    .A(net6765),
    .B(_07812_));
 sg13g2_a21oi_1 _39839_ (.A1(_07806_),
    .A2(_09241_),
    .Y(_09251_),
    .B1(_07848_));
 sg13g2_nor3_1 _39840_ (.A(_07815_),
    .B(_07852_),
    .C(_09251_),
    .Y(_09252_));
 sg13g2_o21ai_1 _39841_ (.B1(_07815_),
    .Y(_09253_),
    .A1(_07852_),
    .A2(_09251_));
 sg13g2_nand2_1 _39842_ (.Y(_09254_),
    .A(net6809),
    .B(_09253_));
 sg13g2_o21ai_1 _39843_ (.B1(_09250_),
    .Y(_09255_),
    .A1(_09252_),
    .A2(_09254_));
 sg13g2_nand2_1 _39844_ (.Y(_09256_),
    .A(net5645),
    .B(_09255_));
 sg13g2_xnor2_1 _39845_ (.Y(_09257_),
    .A(net5586),
    .B(_09255_));
 sg13g2_xnor2_1 _39846_ (.Y(_09258_),
    .A(net5644),
    .B(_09255_));
 sg13g2_a21oi_1 _39847_ (.A1(_07845_),
    .A2(_09242_),
    .Y(_09259_),
    .B1(net6766));
 sg13g2_o21ai_1 _39848_ (.B1(_09259_),
    .Y(_09260_),
    .A1(_07845_),
    .A2(_09242_));
 sg13g2_o21ai_1 _39849_ (.B1(_09260_),
    .Y(_09261_),
    .A1(net6809),
    .A2(_07843_));
 sg13g2_nor2_1 _39850_ (.A(net5644),
    .B(_09261_),
    .Y(_09262_));
 sg13g2_xnor2_1 _39851_ (.Y(_09263_),
    .A(net5586),
    .B(_09261_));
 sg13g2_a21o_1 _39852_ (.A2(_09240_),
    .A1(_07857_),
    .B1(_07795_),
    .X(_09264_));
 sg13g2_nand2_1 _39853_ (.Y(_09265_),
    .A(net6765),
    .B(_07803_));
 sg13g2_xor2_1 _39854_ (.B(_09264_),
    .A(_07856_),
    .X(_09266_));
 sg13g2_o21ai_1 _39855_ (.B1(_09265_),
    .Y(_09267_),
    .A1(net6766),
    .A2(_09266_));
 sg13g2_inv_1 _39856_ (.Y(_09268_),
    .A(_09267_));
 sg13g2_xnor2_1 _39857_ (.Y(_09269_),
    .A(net5644),
    .B(_09267_));
 sg13g2_and4_1 _39858_ (.A(_09248_),
    .B(_09257_),
    .C(_09263_),
    .D(_09269_),
    .X(_09270_));
 sg13g2_nor2_1 _39859_ (.A(net6809),
    .B(_07719_),
    .Y(_09271_));
 sg13g2_xnor2_1 _39860_ (.Y(_09272_),
    .A(_08118_),
    .B(_08120_));
 sg13g2_a21oi_2 _39861_ (.B1(_09271_),
    .Y(_09273_),
    .A2(_09272_),
    .A1(net6809));
 sg13g2_nand2_1 _39862_ (.Y(_09274_),
    .A(net5644),
    .B(_09273_));
 sg13g2_xnor2_1 _39863_ (.Y(_09275_),
    .A(net5644),
    .B(_09273_));
 sg13g2_nand2_1 _39864_ (.Y(_09276_),
    .A(net6767),
    .B(_07787_));
 sg13g2_a22oi_1 _39865_ (.Y(_09277_),
    .B1(_07850_),
    .B2(_09253_),
    .A2(_07823_),
    .A1(net5854));
 sg13g2_a21oi_1 _39866_ (.A1(_07778_),
    .A2(_09277_),
    .Y(_09278_),
    .B1(_07777_));
 sg13g2_xnor2_1 _39867_ (.Y(_09279_),
    .A(_07788_),
    .B(_09278_));
 sg13g2_o21ai_1 _39868_ (.B1(_09276_),
    .Y(_09280_),
    .A1(net6767),
    .A2(_09279_));
 sg13g2_or2_1 _39869_ (.X(_09281_),
    .B(_09280_),
    .A(net5586));
 sg13g2_inv_1 _39870_ (.Y(_09282_),
    .A(_09281_));
 sg13g2_xnor2_1 _39871_ (.Y(_09283_),
    .A(net5586),
    .B(_09280_));
 sg13g2_inv_1 _39872_ (.Y(_09284_),
    .A(_09283_));
 sg13g2_nor2_1 _39873_ (.A(_09275_),
    .B(_09283_),
    .Y(_09285_));
 sg13g2_nor2_1 _39874_ (.A(net6809),
    .B(_07776_),
    .Y(_09286_));
 sg13g2_xnor2_1 _39875_ (.Y(_09287_),
    .A(_07779_),
    .B(_09277_));
 sg13g2_a21oi_2 _39876_ (.B1(_09286_),
    .Y(_09288_),
    .A2(_09287_),
    .A1(net6809));
 sg13g2_inv_2 _39877_ (.Y(_09289_),
    .A(_09288_));
 sg13g2_nand2_1 _39878_ (.Y(_09290_),
    .A(net5645),
    .B(_09289_));
 sg13g2_xnor2_1 _39879_ (.Y(_09291_),
    .A(net5586),
    .B(_09288_));
 sg13g2_nand2_1 _39880_ (.Y(_09292_),
    .A(_07813_),
    .B(_09253_));
 sg13g2_xnor2_1 _39881_ (.Y(_09293_),
    .A(_07825_),
    .B(_09292_));
 sg13g2_nor2_1 _39882_ (.A(net6766),
    .B(_09293_),
    .Y(_09294_));
 sg13g2_a21oi_2 _39883_ (.B1(_09294_),
    .Y(_09295_),
    .A2(_07823_),
    .A1(net6766));
 sg13g2_nand2_1 _39884_ (.Y(_09296_),
    .A(net5645),
    .B(_09295_));
 sg13g2_xnor2_1 _39885_ (.Y(_09297_),
    .A(net5645),
    .B(_09295_));
 sg13g2_nor4_1 _39886_ (.A(_09275_),
    .B(_09283_),
    .C(_09291_),
    .D(_09297_),
    .Y(_09298_));
 sg13g2_and2_1 _39887_ (.A(_09270_),
    .B(_09298_),
    .X(_09299_));
 sg13g2_nand2_1 _39888_ (.Y(_09300_),
    .A(net6765),
    .B(_07794_));
 sg13g2_xnor2_1 _39889_ (.Y(_09301_),
    .A(_07857_),
    .B(_09240_));
 sg13g2_o21ai_1 _39890_ (.B1(_09300_),
    .Y(_09302_),
    .A1(net6765),
    .A2(_09301_));
 sg13g2_nand2_1 _39891_ (.Y(_09303_),
    .A(net5634),
    .B(_09302_));
 sg13g2_xnor2_1 _39892_ (.Y(_09304_),
    .A(net5585),
    .B(_09302_));
 sg13g2_nor2b_1 _39893_ (.A(_08110_),
    .B_N(_08115_),
    .Y(_09305_));
 sg13g2_o21ai_1 _39894_ (.B1(_07905_),
    .Y(_09306_),
    .A1(_07947_),
    .A2(_09305_));
 sg13g2_nand2_1 _39895_ (.Y(_09307_),
    .A(_07904_),
    .B(_09306_));
 sg13g2_nand3_1 _39896_ (.B(_07906_),
    .C(_09307_),
    .A(_07888_),
    .Y(_09308_));
 sg13g2_nand2_1 _39897_ (.Y(_09309_),
    .A(_07887_),
    .B(_09308_));
 sg13g2_xor2_1 _39898_ (.B(_09309_),
    .A(_07881_),
    .X(_09310_));
 sg13g2_nor2_1 _39899_ (.A(net6765),
    .B(_09310_),
    .Y(_09311_));
 sg13g2_a21oi_2 _39900_ (.B1(_09311_),
    .Y(_09312_),
    .A2(_07880_),
    .A1(net6765));
 sg13g2_nand2_1 _39901_ (.Y(_09313_),
    .A(net5634),
    .B(_09312_));
 sg13g2_xnor2_1 _39902_ (.Y(_09314_),
    .A(net5585),
    .B(_09312_));
 sg13g2_nand2_1 _39903_ (.Y(_09315_),
    .A(_09304_),
    .B(_09314_));
 sg13g2_a21o_1 _39904_ (.A2(_09307_),
    .A1(_07906_),
    .B1(_07888_),
    .X(_09316_));
 sg13g2_and2_1 _39905_ (.A(_09308_),
    .B(_09316_),
    .X(_09317_));
 sg13g2_mux2_1 _39906_ (.A0(_07886_),
    .A1(_09317_),
    .S(net6803),
    .X(_09318_));
 sg13g2_and2_1 _39907_ (.A(net5634),
    .B(_09318_),
    .X(_09319_));
 sg13g2_nor2_1 _39908_ (.A(net5634),
    .B(_09318_),
    .Y(_09320_));
 sg13g2_nor2_1 _39909_ (.A(_09319_),
    .B(_09320_),
    .Y(_09321_));
 sg13g2_nand2_1 _39910_ (.Y(_09322_),
    .A(net6765),
    .B(_07903_));
 sg13g2_nand2b_1 _39911_ (.Y(_09323_),
    .B(_09306_),
    .A_N(_07896_));
 sg13g2_xnor2_1 _39912_ (.Y(_09324_),
    .A(_07907_),
    .B(_09323_));
 sg13g2_o21ai_1 _39913_ (.B1(_09322_),
    .Y(_09325_),
    .A1(net6765),
    .A2(_09324_));
 sg13g2_nand2_1 _39914_ (.Y(_09326_),
    .A(net5634),
    .B(_09325_));
 sg13g2_xnor2_1 _39915_ (.Y(_09327_),
    .A(net5634),
    .B(_09325_));
 sg13g2_nor4_1 _39916_ (.A(_09315_),
    .B(_09319_),
    .C(_09320_),
    .D(_09327_),
    .Y(_09328_));
 sg13g2_or3_1 _39917_ (.A(_07905_),
    .B(_07947_),
    .C(_09305_),
    .X(_09329_));
 sg13g2_a21oi_1 _39918_ (.A1(_09306_),
    .A2(_09329_),
    .Y(_09330_),
    .B1(net6759));
 sg13g2_a21oi_2 _39919_ (.B1(_09330_),
    .Y(_09331_),
    .A2(_07895_),
    .A1(net6759));
 sg13g2_xnor2_1 _39920_ (.Y(_09332_),
    .A(net5633),
    .B(_09331_));
 sg13g2_nor2b_1 _39921_ (.A(_09174_),
    .B_N(_07944_),
    .Y(_09333_));
 sg13g2_nor2_1 _39922_ (.A(_08111_),
    .B(_09333_),
    .Y(_09334_));
 sg13g2_nand2b_1 _39923_ (.Y(_09335_),
    .B(_09334_),
    .A_N(_07918_));
 sg13g2_nand2_1 _39924_ (.Y(_09336_),
    .A(_07917_),
    .B(_09335_));
 sg13g2_xnor2_1 _39925_ (.Y(_09337_),
    .A(_07927_),
    .B(_09336_));
 sg13g2_nor2_1 _39926_ (.A(net6759),
    .B(_09337_),
    .Y(_09338_));
 sg13g2_a21oi_2 _39927_ (.B1(_09338_),
    .Y(_09339_),
    .A2(_07926_),
    .A1(net6759));
 sg13g2_xnor2_1 _39928_ (.Y(_09340_),
    .A(net5633),
    .B(_09339_));
 sg13g2_nand2_1 _39929_ (.Y(_09341_),
    .A(net6759),
    .B(_07916_));
 sg13g2_xor2_1 _39930_ (.B(_09334_),
    .A(_07918_),
    .X(_09342_));
 sg13g2_o21ai_1 _39931_ (.B1(_09341_),
    .Y(_09343_),
    .A1(net6760),
    .A2(_09342_));
 sg13g2_nand2_1 _39932_ (.Y(_09344_),
    .A(net5633),
    .B(_09343_));
 sg13g2_xnor2_1 _39933_ (.Y(_09345_),
    .A(net5633),
    .B(_09343_));
 sg13g2_nor2_1 _39934_ (.A(net6803),
    .B(_07936_),
    .Y(_09346_));
 sg13g2_a21oi_1 _39935_ (.A1(net5794),
    .A2(_07943_),
    .Y(_09347_),
    .B1(_09174_));
 sg13g2_xnor2_1 _39936_ (.Y(_09348_),
    .A(_08112_),
    .B(_09347_));
 sg13g2_a21oi_2 _39937_ (.B1(_09346_),
    .Y(_09349_),
    .A2(_09348_),
    .A1(net6803));
 sg13g2_xnor2_1 _39938_ (.Y(_09350_),
    .A(net5633),
    .B(_09349_));
 sg13g2_nor4_1 _39939_ (.A(_09332_),
    .B(_09340_),
    .C(_09345_),
    .D(_09350_),
    .Y(_09351_));
 sg13g2_nand2_1 _39940_ (.Y(_09352_),
    .A(_09328_),
    .B(_09351_));
 sg13g2_nand3_1 _39941_ (.B(_09328_),
    .C(_09351_),
    .A(_09299_),
    .Y(_09353_));
 sg13g2_a21oi_2 _39942_ (.B1(_09353_),
    .Y(_09354_),
    .A2(_09238_),
    .A1(_09232_));
 sg13g2_o21ai_1 _39943_ (.B1(net5633),
    .Y(_09355_),
    .A1(_09343_),
    .A2(_09349_));
 sg13g2_nor3_1 _39944_ (.A(_09332_),
    .B(_09340_),
    .C(_09355_),
    .Y(_09356_));
 sg13g2_o21ai_1 _39945_ (.B1(net5634),
    .Y(_09357_),
    .A1(_09331_),
    .A2(_09339_));
 sg13g2_nand2b_1 _39946_ (.Y(_09358_),
    .B(_09357_),
    .A_N(_09356_));
 sg13g2_inv_1 _39947_ (.Y(_09359_),
    .A(_09358_));
 sg13g2_o21ai_1 _39948_ (.B1(net5634),
    .Y(_09360_),
    .A1(_09318_),
    .A2(_09325_));
 sg13g2_nand3b_1 _39949_ (.B(_09314_),
    .C(_09304_),
    .Y(_09361_),
    .A_N(_09360_));
 sg13g2_nand3_1 _39950_ (.B(_09313_),
    .C(_09361_),
    .A(_09303_),
    .Y(_09362_));
 sg13g2_a21o_1 _39951_ (.A2(_09358_),
    .A1(_09328_),
    .B1(_09362_),
    .X(_09363_));
 sg13g2_nand2_1 _39952_ (.Y(_09364_),
    .A(_09290_),
    .B(_09296_));
 sg13g2_o21ai_1 _39953_ (.B1(net5644),
    .Y(_09365_),
    .A1(_09261_),
    .A2(_09268_));
 sg13g2_nor3_1 _39954_ (.A(_09249_),
    .B(_09258_),
    .C(_09365_),
    .Y(_09366_));
 sg13g2_nand2_1 _39955_ (.Y(_09367_),
    .A(_09247_),
    .B(_09256_));
 sg13g2_or2_1 _39956_ (.X(_09368_),
    .B(_09367_),
    .A(_09366_));
 sg13g2_o21ai_1 _39957_ (.B1(_09298_),
    .Y(_09369_),
    .A1(_09366_),
    .A2(_09367_));
 sg13g2_a21oi_1 _39958_ (.A1(_09285_),
    .A2(_09364_),
    .Y(_09370_),
    .B1(_09282_));
 sg13g2_nand3_1 _39959_ (.B(_09369_),
    .C(_09370_),
    .A(_09274_),
    .Y(_09371_));
 sg13g2_a21o_2 _39960_ (.A2(_09363_),
    .A1(_09299_),
    .B1(_09371_),
    .X(_09372_));
 sg13g2_nor2_1 _39961_ (.A(_09354_),
    .B(_09372_),
    .Y(_09373_));
 sg13g2_a21oi_1 _39962_ (.A1(_07737_),
    .A2(_08126_),
    .Y(_09374_),
    .B1(_07539_));
 sg13g2_nor2_1 _39963_ (.A(_07755_),
    .B(_09374_),
    .Y(_09375_));
 sg13g2_nor2b_1 _39964_ (.A(_09375_),
    .B_N(_07434_),
    .Y(_09376_));
 sg13g2_o21ai_1 _39965_ (.B1(_07445_),
    .Y(_09377_),
    .A1(_07755_),
    .A2(_09374_));
 sg13g2_o21ai_1 _39966_ (.B1(_07742_),
    .Y(_09378_),
    .A1(_07427_),
    .A2(_09377_));
 sg13g2_a21oi_1 _39967_ (.A1(_07405_),
    .A2(_09378_),
    .Y(_09379_),
    .B1(_07404_));
 sg13g2_nand3_1 _39968_ (.B(_07405_),
    .C(_09378_),
    .A(_07396_),
    .Y(_09380_));
 sg13g2_a21o_1 _39969_ (.A2(_09380_),
    .A1(_07744_),
    .B1(_07379_),
    .X(_09381_));
 sg13g2_a21oi_1 _39970_ (.A1(_07378_),
    .A2(_09381_),
    .Y(_09382_),
    .B1(_07389_));
 sg13g2_and3_1 _39971_ (.X(_09383_),
    .A(_07378_),
    .B(_07389_),
    .C(_09381_));
 sg13g2_nor2_1 _39972_ (.A(net6821),
    .B(_07387_),
    .Y(_09384_));
 sg13g2_inv_1 _39973_ (.Y(_09385_),
    .A(_09384_));
 sg13g2_o21ai_1 _39974_ (.B1(net6821),
    .Y(_09386_),
    .A1(_09382_),
    .A2(_09383_));
 sg13g2_and2_1 _39975_ (.A(_09385_),
    .B(_09386_),
    .X(_09387_));
 sg13g2_and3_2 _39976_ (.X(_09388_),
    .A(net5666),
    .B(_09385_),
    .C(_09386_));
 sg13g2_nand2_1 _39977_ (.Y(_09389_),
    .A(net5664),
    .B(_09387_));
 sg13g2_a21oi_2 _39978_ (.B1(net5666),
    .Y(_09390_),
    .A2(_09386_),
    .A1(_09385_));
 sg13g2_nor2_1 _39979_ (.A(_09388_),
    .B(_09390_),
    .Y(_09391_));
 sg13g2_a21oi_1 _39980_ (.A1(_08129_),
    .A2(_08132_),
    .Y(_09392_),
    .B1(net6785));
 sg13g2_o21ai_1 _39981_ (.B1(_09392_),
    .Y(_09393_),
    .A1(_08129_),
    .A2(_08132_));
 sg13g2_o21ai_1 _39982_ (.B1(_09393_),
    .Y(_09394_),
    .A1(net6830),
    .A2(_07324_));
 sg13g2_xnor2_1 _39983_ (.Y(_09395_),
    .A(net5666),
    .B(_09394_));
 sg13g2_nor3_1 _39984_ (.A(_09388_),
    .B(_09390_),
    .C(_09395_),
    .Y(_09396_));
 sg13g2_nor2_1 _39985_ (.A(net6821),
    .B(_07395_),
    .Y(_09397_));
 sg13g2_xor2_1 _39986_ (.B(_09379_),
    .A(_07396_),
    .X(_09398_));
 sg13g2_a21oi_2 _39987_ (.B1(_09397_),
    .Y(_09399_),
    .A2(_09398_),
    .A1(net6821));
 sg13g2_and2_1 _39988_ (.A(net5664),
    .B(_09399_),
    .X(_09400_));
 sg13g2_xnor2_1 _39989_ (.Y(_09401_),
    .A(net5664),
    .B(_09399_));
 sg13g2_nand3_1 _39990_ (.B(_07744_),
    .C(_09380_),
    .A(_07379_),
    .Y(_09402_));
 sg13g2_a21o_1 _39991_ (.A2(_09402_),
    .A1(_09381_),
    .B1(net6776),
    .X(_09403_));
 sg13g2_nand2b_1 _39992_ (.Y(_09404_),
    .B(net6775),
    .A_N(_07377_));
 sg13g2_nand2_1 _39993_ (.Y(_09405_),
    .A(_09403_),
    .B(_09404_));
 sg13g2_nand3_1 _39994_ (.B(_09403_),
    .C(_09404_),
    .A(net5664),
    .Y(_09406_));
 sg13g2_a21o_1 _39995_ (.A2(_09404_),
    .A1(_09403_),
    .B1(net5664),
    .X(_09407_));
 sg13g2_and2_1 _39996_ (.A(_09406_),
    .B(_09407_),
    .X(_09408_));
 sg13g2_nand3b_1 _39997_ (.B(_09406_),
    .C(_09407_),
    .Y(_09409_),
    .A_N(_09401_));
 sg13g2_nor4_1 _39998_ (.A(_09388_),
    .B(_09390_),
    .C(_09395_),
    .D(_09409_),
    .Y(_09410_));
 sg13g2_nand2_1 _39999_ (.Y(_09411_),
    .A(net6776),
    .B(_07417_));
 sg13g2_a21oi_1 _40000_ (.A1(_07739_),
    .A2(_09377_),
    .Y(_09412_),
    .B1(_07426_));
 sg13g2_nor2_1 _40001_ (.A(_07425_),
    .B(_09412_),
    .Y(_09413_));
 sg13g2_xor2_1 _40002_ (.B(_09413_),
    .A(_07418_),
    .X(_09414_));
 sg13g2_o21ai_1 _40003_ (.B1(_09411_),
    .Y(_09415_),
    .A1(net6776),
    .A2(_09414_));
 sg13g2_inv_1 _40004_ (.Y(_09416_),
    .A(_09415_));
 sg13g2_or2_1 _40005_ (.X(_09417_),
    .B(_09415_),
    .A(net5595));
 sg13g2_xnor2_1 _40006_ (.Y(_09418_),
    .A(net5595),
    .B(_09415_));
 sg13g2_nand2_1 _40007_ (.Y(_09419_),
    .A(net6776),
    .B(_07402_));
 sg13g2_xnor2_1 _40008_ (.Y(_09420_),
    .A(_07405_),
    .B(_09378_));
 sg13g2_o21ai_1 _40009_ (.B1(_09419_),
    .Y(_09421_),
    .A1(net6776),
    .A2(_09420_));
 sg13g2_nand2_1 _40010_ (.Y(_09422_),
    .A(net5664),
    .B(_09421_));
 sg13g2_xnor2_1 _40011_ (.Y(_09423_),
    .A(net5595),
    .B(_09421_));
 sg13g2_nor2b_1 _40012_ (.A(_09418_),
    .B_N(_09423_),
    .Y(_09424_));
 sg13g2_nand3_1 _40013_ (.B(_07739_),
    .C(_09377_),
    .A(_07426_),
    .Y(_09425_));
 sg13g2_nand3b_1 _40014_ (.B(_09425_),
    .C(net6823),
    .Y(_09426_),
    .A_N(_09412_));
 sg13g2_o21ai_1 _40015_ (.B1(_09426_),
    .Y(_09427_),
    .A1(net6823),
    .A2(_07424_));
 sg13g2_nor2_1 _40016_ (.A(net5666),
    .B(_09427_),
    .Y(_09428_));
 sg13g2_xnor2_1 _40017_ (.Y(_09429_),
    .A(net5595),
    .B(_09427_));
 sg13g2_a21o_1 _40018_ (.A2(_07433_),
    .A1(net5815),
    .B1(_09376_),
    .X(_09430_));
 sg13g2_nor2_1 _40019_ (.A(net6821),
    .B(_07441_),
    .Y(_09431_));
 sg13g2_xnor2_1 _40020_ (.Y(_09432_),
    .A(_07443_),
    .B(_09430_));
 sg13g2_a21oi_2 _40021_ (.B1(_09431_),
    .Y(_09433_),
    .A2(_09432_),
    .A1(net6821));
 sg13g2_nand2_1 _40022_ (.Y(_09434_),
    .A(net5666),
    .B(_09433_));
 sg13g2_xnor2_1 _40023_ (.Y(_09435_),
    .A(net5595),
    .B(_09433_));
 sg13g2_and3_1 _40024_ (.X(_09436_),
    .A(_09424_),
    .B(_09429_),
    .C(_09435_));
 sg13g2_nand2_1 _40025_ (.Y(_09437_),
    .A(_09410_),
    .B(_09436_));
 sg13g2_a21oi_1 _40026_ (.A1(_07737_),
    .A2(_08126_),
    .Y(_09438_),
    .B1(_07538_));
 sg13g2_nor2_1 _40027_ (.A(_07750_),
    .B(_09438_),
    .Y(_09439_));
 sg13g2_o21ai_1 _40028_ (.B1(_07496_),
    .Y(_09440_),
    .A1(_07750_),
    .A2(_09438_));
 sg13g2_nand2_1 _40029_ (.Y(_09441_),
    .A(_07495_),
    .B(_09440_));
 sg13g2_a21oi_1 _40030_ (.A1(_07752_),
    .A2(_09440_),
    .Y(_09442_),
    .B1(_07488_));
 sg13g2_a21oi_1 _40031_ (.A1(_07464_),
    .A2(_09442_),
    .Y(_09443_),
    .B1(_07462_));
 sg13g2_xnor2_1 _40032_ (.Y(_09444_),
    .A(_07476_),
    .B(_09443_));
 sg13g2_mux2_1 _40033_ (.A0(_07473_),
    .A1(_09444_),
    .S(net6821),
    .X(_09445_));
 sg13g2_nand2_1 _40034_ (.Y(_09446_),
    .A(net5657),
    .B(_09445_));
 sg13g2_xnor2_1 _40035_ (.Y(_09447_),
    .A(net5655),
    .B(_09445_));
 sg13g2_nand2_1 _40036_ (.Y(_09448_),
    .A(net6776),
    .B(_07433_));
 sg13g2_xor2_1 _40037_ (.B(_09375_),
    .A(_07434_),
    .X(_09449_));
 sg13g2_o21ai_1 _40038_ (.B1(_09448_),
    .Y(_09450_),
    .A1(net6776),
    .A2(_09449_));
 sg13g2_nand2_1 _40039_ (.Y(_09451_),
    .A(net5655),
    .B(_09450_));
 sg13g2_xnor2_1 _40040_ (.Y(_09452_),
    .A(net5655),
    .B(_09450_));
 sg13g2_a21oi_1 _40041_ (.A1(_07464_),
    .A2(_09442_),
    .Y(_09453_),
    .B1(net6776));
 sg13g2_o21ai_1 _40042_ (.B1(_09453_),
    .Y(_09454_),
    .A1(_07464_),
    .A2(_09442_));
 sg13g2_o21ai_1 _40043_ (.B1(_09454_),
    .Y(_09455_),
    .A1(net6821),
    .A2(_07461_));
 sg13g2_xnor2_1 _40044_ (.Y(_09456_),
    .A(net5655),
    .B(_09455_));
 sg13g2_xor2_1 _40045_ (.B(_09441_),
    .A(_07489_),
    .X(_09457_));
 sg13g2_mux2_1 _40046_ (.A0(_07487_),
    .A1(_09457_),
    .S(net6816),
    .X(_09458_));
 sg13g2_nand2_1 _40047_ (.Y(_09459_),
    .A(net5655),
    .B(_09458_));
 sg13g2_xnor2_1 _40048_ (.Y(_09460_),
    .A(net5655),
    .B(_09458_));
 sg13g2_nor4_1 _40049_ (.A(_09447_),
    .B(_09452_),
    .C(_09456_),
    .D(_09460_),
    .Y(_09461_));
 sg13g2_a21oi_1 _40050_ (.A1(_07737_),
    .A2(_08126_),
    .Y(_09462_),
    .B1(_07536_));
 sg13g2_o21ai_1 _40051_ (.B1(_07527_),
    .Y(_09463_),
    .A1(_07748_),
    .A2(_09462_));
 sg13g2_nor2_1 _40052_ (.A(_07504_),
    .B(_09463_),
    .Y(_09464_));
 sg13g2_o21ai_1 _40053_ (.B1(_07515_),
    .Y(_09465_),
    .A1(_07503_),
    .A2(_09464_));
 sg13g2_or3_1 _40054_ (.A(_07503_),
    .B(_07515_),
    .C(_09464_),
    .X(_09466_));
 sg13g2_nand3_1 _40055_ (.B(_09465_),
    .C(_09466_),
    .A(net6816),
    .Y(_09467_));
 sg13g2_o21ai_1 _40056_ (.B1(_09467_),
    .Y(_09468_),
    .A1(net6816),
    .A2(_07513_));
 sg13g2_nand2_1 _40057_ (.Y(_09469_),
    .A(net5656),
    .B(_09468_));
 sg13g2_xnor2_1 _40058_ (.Y(_09470_),
    .A(net5594),
    .B(_09468_));
 sg13g2_xnor2_1 _40059_ (.Y(_09471_),
    .A(net5656),
    .B(_09468_));
 sg13g2_nand2_1 _40060_ (.Y(_09472_),
    .A(net6772),
    .B(_07494_));
 sg13g2_xor2_1 _40061_ (.B(_09439_),
    .A(_07496_),
    .X(_09473_));
 sg13g2_o21ai_1 _40062_ (.B1(_09472_),
    .Y(_09474_),
    .A1(net6772),
    .A2(_09473_));
 sg13g2_nand2_1 _40063_ (.Y(_09475_),
    .A(net5657),
    .B(_09474_));
 sg13g2_xnor2_1 _40064_ (.Y(_09476_),
    .A(net5594),
    .B(_09474_));
 sg13g2_xnor2_1 _40065_ (.Y(_09477_),
    .A(net5656),
    .B(_09474_));
 sg13g2_nand2_1 _40066_ (.Y(_09478_),
    .A(net6772),
    .B(_07502_));
 sg13g2_xnor2_1 _40067_ (.Y(_09479_),
    .A(_07504_),
    .B(_09463_));
 sg13g2_o21ai_1 _40068_ (.B1(_09478_),
    .Y(_09480_),
    .A1(net6773),
    .A2(_09479_));
 sg13g2_nor2_1 _40069_ (.A(net5656),
    .B(_09480_),
    .Y(_09481_));
 sg13g2_xnor2_1 _40070_ (.Y(_09482_),
    .A(net5594),
    .B(_09480_));
 sg13g2_nor2_1 _40071_ (.A(net6816),
    .B(_07526_),
    .Y(_09483_));
 sg13g2_nor2_1 _40072_ (.A(_07534_),
    .B(_09462_),
    .Y(_09484_));
 sg13g2_xnor2_1 _40073_ (.Y(_09485_),
    .A(_07528_),
    .B(_09484_));
 sg13g2_a21oi_2 _40074_ (.B1(_09483_),
    .Y(_09486_),
    .A2(_09485_),
    .A1(net6816));
 sg13g2_inv_2 _40075_ (.Y(_09487_),
    .A(_09486_));
 sg13g2_nand2_1 _40076_ (.Y(_09488_),
    .A(net5656),
    .B(_09487_));
 sg13g2_xnor2_1 _40077_ (.Y(_09489_),
    .A(net5656),
    .B(_09486_));
 sg13g2_and4_1 _40078_ (.A(_09470_),
    .B(_09476_),
    .C(_09482_),
    .D(_09489_),
    .X(_09490_));
 sg13g2_inv_1 _40079_ (.Y(_09491_),
    .A(_09490_));
 sg13g2_and2_1 _40080_ (.A(_09461_),
    .B(_09490_),
    .X(_09492_));
 sg13g2_inv_1 _40081_ (.Y(_09493_),
    .A(_09492_));
 sg13g2_and3_2 _40082_ (.X(_09494_),
    .A(_09410_),
    .B(_09436_),
    .C(_09492_));
 sg13g2_and2_1 _40083_ (.A(net6771),
    .B(_07603_),
    .X(_09495_));
 sg13g2_nand3_1 _40084_ (.B(net1083),
    .C(_08124_),
    .A(_07860_),
    .Y(_09496_));
 sg13g2_nand3_1 _40085_ (.B(_07727_),
    .C(_09496_),
    .A(_07726_),
    .Y(_09497_));
 sg13g2_a21oi_1 _40086_ (.A1(_07633_),
    .A2(_09497_),
    .Y(_09498_),
    .B1(_07729_));
 sg13g2_o21ai_1 _40087_ (.B1(_07611_),
    .Y(_09499_),
    .A1(_07612_),
    .A2(_09498_));
 sg13g2_xor2_1 _40088_ (.B(_09499_),
    .A(_07605_),
    .X(_09500_));
 sg13g2_a21oi_2 _40089_ (.B1(_09495_),
    .Y(_09501_),
    .A2(_09500_),
    .A1(net6817));
 sg13g2_nand2_1 _40090_ (.Y(_09502_),
    .A(net5652),
    .B(_09501_));
 sg13g2_inv_1 _40091_ (.Y(_09503_),
    .A(_09502_));
 sg13g2_xnor2_1 _40092_ (.Y(_09504_),
    .A(net5591),
    .B(_09501_));
 sg13g2_nand2_1 _40093_ (.Y(_09505_),
    .A(net6772),
    .B(_07590_));
 sg13g2_and4_1 _40094_ (.A(_07614_),
    .B(_07622_),
    .C(_07632_),
    .D(_09497_),
    .X(_09506_));
 sg13g2_nor2_1 _40095_ (.A(_07732_),
    .B(_09506_),
    .Y(_09507_));
 sg13g2_o21ai_1 _40096_ (.B1(_07593_),
    .Y(_09508_),
    .A1(_07732_),
    .A2(_09506_));
 sg13g2_xnor2_1 _40097_ (.Y(_09509_),
    .A(_07592_),
    .B(_09507_));
 sg13g2_o21ai_1 _40098_ (.B1(_09505_),
    .Y(_09510_),
    .A1(net6772),
    .A2(_09509_));
 sg13g2_xnor2_1 _40099_ (.Y(_09511_),
    .A(net5591),
    .B(_09510_));
 sg13g2_nand2_1 _40100_ (.Y(_09512_),
    .A(_09504_),
    .B(_09511_));
 sg13g2_nand2_1 _40101_ (.Y(_09513_),
    .A(net6771),
    .B(_07610_));
 sg13g2_xnor2_1 _40102_ (.Y(_09514_),
    .A(_07612_),
    .B(_09498_));
 sg13g2_o21ai_1 _40103_ (.B1(_09513_),
    .Y(_09515_),
    .A1(net6771),
    .A2(_09514_));
 sg13g2_nor2_1 _40104_ (.A(net5653),
    .B(_09515_),
    .Y(_09516_));
 sg13g2_nand2_1 _40105_ (.Y(_09517_),
    .A(net5653),
    .B(_09515_));
 sg13g2_xnor2_1 _40106_ (.Y(_09518_),
    .A(net5591),
    .B(_09515_));
 sg13g2_a21oi_1 _40107_ (.A1(_07622_),
    .A2(_09497_),
    .Y(_09519_),
    .B1(_07621_));
 sg13g2_a21oi_1 _40108_ (.A1(_07625_),
    .A2(_07630_),
    .Y(_09520_),
    .B1(net6817));
 sg13g2_xor2_1 _40109_ (.B(_09519_),
    .A(_07632_),
    .X(_09521_));
 sg13g2_a21oi_2 _40110_ (.B1(_09520_),
    .Y(_09522_),
    .A2(_09521_),
    .A1(net6817));
 sg13g2_and2_1 _40111_ (.A(net5653),
    .B(_09522_),
    .X(_09523_));
 sg13g2_xnor2_1 _40112_ (.Y(_09524_),
    .A(net5591),
    .B(_09522_));
 sg13g2_and4_1 _40113_ (.A(_09504_),
    .B(_09511_),
    .C(_09518_),
    .D(_09524_),
    .X(_09525_));
 sg13g2_inv_1 _40114_ (.Y(_09526_),
    .A(_09525_));
 sg13g2_nor2_1 _40115_ (.A(net6816),
    .B(_07533_),
    .Y(_09527_));
 sg13g2_nand3_1 _40116_ (.B(_07737_),
    .C(_08126_),
    .A(_07536_),
    .Y(_09528_));
 sg13g2_nor2b_1 _40117_ (.A(_09462_),
    .B_N(_09528_),
    .Y(_09529_));
 sg13g2_a21oi_2 _40118_ (.B1(_09527_),
    .Y(_09530_),
    .A2(_09529_),
    .A1(net6820));
 sg13g2_inv_1 _40119_ (.Y(_09531_),
    .A(_09530_));
 sg13g2_xnor2_1 _40120_ (.Y(_09532_),
    .A(net5653),
    .B(_09530_));
 sg13g2_and2_1 _40121_ (.A(net6772),
    .B(_07570_),
    .X(_09533_));
 sg13g2_nand2_1 _40122_ (.Y(_09534_),
    .A(_07591_),
    .B(_09508_));
 sg13g2_a21o_1 _40123_ (.A2(_09508_),
    .A1(_07734_),
    .B1(_07584_),
    .X(_09535_));
 sg13g2_o21ai_1 _40124_ (.B1(_07560_),
    .Y(_09536_),
    .A1(_07562_),
    .A2(_09535_));
 sg13g2_xnor2_1 _40125_ (.Y(_09537_),
    .A(_07572_),
    .B(_09536_));
 sg13g2_a21oi_2 _40126_ (.B1(_09533_),
    .Y(_09538_),
    .A2(_09537_),
    .A1(net6816));
 sg13g2_and2_1 _40127_ (.A(net5653),
    .B(_09538_),
    .X(_09539_));
 sg13g2_xnor2_1 _40128_ (.Y(_09540_),
    .A(net5591),
    .B(_09538_));
 sg13g2_and2_1 _40129_ (.A(_09532_),
    .B(_09540_),
    .X(_09541_));
 sg13g2_nand2_1 _40130_ (.Y(_09542_),
    .A(net6772),
    .B(_07559_));
 sg13g2_xnor2_1 _40131_ (.Y(_09543_),
    .A(_07562_),
    .B(_09535_));
 sg13g2_o21ai_1 _40132_ (.B1(_09542_),
    .Y(_09544_),
    .A1(net6772),
    .A2(_09543_));
 sg13g2_nor2_1 _40133_ (.A(net5653),
    .B(_09544_),
    .Y(_09545_));
 sg13g2_xnor2_1 _40134_ (.Y(_09546_),
    .A(net5653),
    .B(_09544_));
 sg13g2_xor2_1 _40135_ (.B(_09534_),
    .A(_07585_),
    .X(_09547_));
 sg13g2_nor2_1 _40136_ (.A(net6817),
    .B(_07582_),
    .Y(_09548_));
 sg13g2_a21oi_1 _40137_ (.A1(net6816),
    .A2(_09547_),
    .Y(_09549_),
    .B1(_09548_));
 sg13g2_inv_2 _40138_ (.Y(_09550_),
    .A(_09549_));
 sg13g2_nand2_1 _40139_ (.Y(_09551_),
    .A(net5654),
    .B(_09550_));
 sg13g2_xnor2_1 _40140_ (.Y(_09552_),
    .A(net5591),
    .B(_09549_));
 sg13g2_inv_1 _40141_ (.Y(_09553_),
    .A(_09552_));
 sg13g2_nor2_1 _40142_ (.A(_09546_),
    .B(_09552_),
    .Y(_09554_));
 sg13g2_nand4_1 _40143_ (.B(_09532_),
    .C(_09540_),
    .A(_09525_),
    .Y(_09555_),
    .D(_09554_));
 sg13g2_a21oi_1 _40144_ (.A1(_07622_),
    .A2(_09497_),
    .Y(_09556_),
    .B1(net6771));
 sg13g2_o21ai_1 _40145_ (.B1(_09556_),
    .Y(_09557_),
    .A1(_07622_),
    .A2(_09497_));
 sg13g2_o21ai_1 _40146_ (.B1(_09557_),
    .Y(_09558_),
    .A1(net6817),
    .A2(_07620_));
 sg13g2_xnor2_1 _40147_ (.Y(_09559_),
    .A(net5591),
    .B(_09558_));
 sg13g2_and2_1 _40148_ (.A(net6770),
    .B(_07660_),
    .X(_09560_));
 sg13g2_nand3_1 _40149_ (.B(net1083),
    .C(_08122_),
    .A(_07860_),
    .Y(_09561_));
 sg13g2_nand4_1 _40150_ (.B(_07860_),
    .C(net1083),
    .A(_07704_),
    .Y(_09562_),
    .D(_08122_));
 sg13g2_a21oi_1 _40151_ (.A1(_07724_),
    .A2(_09562_),
    .Y(_09563_),
    .B1(_07679_));
 sg13g2_o21ai_1 _40152_ (.B1(_07680_),
    .Y(_09564_),
    .A1(_07678_),
    .A2(_09563_));
 sg13g2_nor2_1 _40153_ (.A(_07651_),
    .B(_09564_),
    .Y(_09565_));
 sg13g2_nor2_1 _40154_ (.A(_07650_),
    .B(_09565_),
    .Y(_09566_));
 sg13g2_xnor2_1 _40155_ (.Y(_09567_),
    .A(_07662_),
    .B(_09566_));
 sg13g2_a21oi_2 _40156_ (.B1(_09560_),
    .Y(_09568_),
    .A2(_09567_),
    .A1(net6817));
 sg13g2_nand2_1 _40157_ (.Y(_09569_),
    .A(net5652),
    .B(_09568_));
 sg13g2_xnor2_1 _40158_ (.Y(_09570_),
    .A(net5591),
    .B(_09568_));
 sg13g2_inv_1 _40159_ (.Y(_09571_),
    .A(_09570_));
 sg13g2_nand2_1 _40160_ (.Y(_09572_),
    .A(_07651_),
    .B(_09564_));
 sg13g2_nor2_1 _40161_ (.A(net6770),
    .B(_09565_),
    .Y(_09573_));
 sg13g2_a22oi_1 _40162_ (.Y(_09574_),
    .B1(_09572_),
    .B2(_09573_),
    .A2(_07649_),
    .A1(net6770));
 sg13g2_inv_2 _40163_ (.Y(_09575_),
    .A(_09574_));
 sg13g2_nand2_1 _40164_ (.Y(_09576_),
    .A(net5652),
    .B(_09575_));
 sg13g2_nor2_1 _40165_ (.A(net5652),
    .B(_09575_),
    .Y(_09577_));
 sg13g2_xnor2_1 _40166_ (.Y(_09578_),
    .A(net5652),
    .B(_09574_));
 sg13g2_nand2_1 _40167_ (.Y(_09579_),
    .A(net6771),
    .B(_07677_));
 sg13g2_a21oi_1 _40168_ (.A1(net5809),
    .A2(_07669_),
    .Y(_09580_),
    .B1(_09563_));
 sg13g2_xor2_1 _40169_ (.B(_09580_),
    .A(_07681_),
    .X(_09581_));
 sg13g2_o21ai_1 _40170_ (.B1(_09579_),
    .Y(_09582_),
    .A1(net6770),
    .A2(_09581_));
 sg13g2_inv_4 _40171_ (.A(_09582_),
    .Y(_09583_));
 sg13g2_nand2_1 _40172_ (.Y(_09584_),
    .A(net5652),
    .B(_09583_));
 sg13g2_xnor2_1 _40173_ (.Y(_09585_),
    .A(net5586),
    .B(_09583_));
 sg13g2_and4_1 _40174_ (.A(_09559_),
    .B(_09570_),
    .C(_09578_),
    .D(_09585_),
    .X(_09586_));
 sg13g2_a21oi_1 _40175_ (.A1(_07720_),
    .A2(_09561_),
    .Y(_09587_),
    .B1(_07693_));
 sg13g2_nor2_1 _40176_ (.A(_07692_),
    .B(_09587_),
    .Y(_09588_));
 sg13g2_xor2_1 _40177_ (.B(_09588_),
    .A(_07703_),
    .X(_09589_));
 sg13g2_nor2_1 _40178_ (.A(net6770),
    .B(_09589_),
    .Y(_09590_));
 sg13g2_a21oi_2 _40179_ (.B1(_09590_),
    .Y(_09591_),
    .A2(_07701_),
    .A1(net6770));
 sg13g2_xnor2_1 _40180_ (.Y(_09592_),
    .A(net5646),
    .B(_09591_));
 sg13g2_nand3_1 _40181_ (.B(_07724_),
    .C(_09562_),
    .A(_07679_),
    .Y(_09593_));
 sg13g2_nand3b_1 _40182_ (.B(_09593_),
    .C(net6817),
    .Y(_09594_),
    .A_N(_09563_));
 sg13g2_o21ai_1 _40183_ (.B1(_09594_),
    .Y(_09595_),
    .A1(net6817),
    .A2(_07670_));
 sg13g2_and2_1 _40184_ (.A(net5646),
    .B(_09595_),
    .X(_09596_));
 sg13g2_xnor2_1 _40185_ (.Y(_09597_),
    .A(net5647),
    .B(_09595_));
 sg13g2_o21ai_1 _40186_ (.B1(_08119_),
    .Y(_09598_),
    .A1(_08118_),
    .A2(_08120_));
 sg13g2_xor2_1 _40187_ (.B(_09598_),
    .A(_08121_),
    .X(_09599_));
 sg13g2_nand2_1 _40188_ (.Y(_09600_),
    .A(net6814),
    .B(_09599_));
 sg13g2_o21ai_1 _40189_ (.B1(_09600_),
    .Y(_09601_),
    .A1(net6814),
    .A2(_07713_));
 sg13g2_inv_2 _40190_ (.Y(_09602_),
    .A(_09601_));
 sg13g2_xnor2_1 _40191_ (.Y(_09603_),
    .A(net5589),
    .B(_09602_));
 sg13g2_nand2_1 _40192_ (.Y(_09604_),
    .A(net6770),
    .B(_07691_));
 sg13g2_nand3_1 _40193_ (.B(_07720_),
    .C(_09561_),
    .A(_07693_),
    .Y(_09605_));
 sg13g2_nand2b_1 _40194_ (.Y(_09606_),
    .B(_09605_),
    .A_N(_09587_));
 sg13g2_o21ai_1 _40195_ (.B1(_09604_),
    .Y(_09607_),
    .A1(net6770),
    .A2(_09606_));
 sg13g2_nor2_1 _40196_ (.A(net5646),
    .B(_09607_),
    .Y(_09608_));
 sg13g2_xnor2_1 _40197_ (.Y(_09609_),
    .A(net5646),
    .B(_09607_));
 sg13g2_nor4_1 _40198_ (.A(_09592_),
    .B(_09597_),
    .C(_09603_),
    .D(_09609_),
    .Y(_09610_));
 sg13g2_and2_1 _40199_ (.A(_09586_),
    .B(_09610_),
    .X(_09611_));
 sg13g2_nor2b_1 _40200_ (.A(_09555_),
    .B_N(_09611_),
    .Y(_09612_));
 sg13g2_and2_1 _40201_ (.A(_09494_),
    .B(_09612_),
    .X(_09613_));
 sg13g2_o21ai_1 _40202_ (.B1(_09613_),
    .Y(_09614_),
    .A1(_09372_),
    .A2(_09354_));
 sg13g2_o21ai_1 _40203_ (.B1(_09607_),
    .Y(_09615_),
    .A1(net5646),
    .A2(_09602_));
 sg13g2_nor3_1 _40204_ (.A(_09592_),
    .B(_09597_),
    .C(_09615_),
    .Y(_09616_));
 sg13g2_a21o_1 _40205_ (.A2(_09591_),
    .A1(net5646),
    .B1(_09596_),
    .X(_09617_));
 sg13g2_nor2_1 _40206_ (.A(_09616_),
    .B(_09617_),
    .Y(_09618_));
 sg13g2_o21ai_1 _40207_ (.B1(_09586_),
    .Y(_09619_),
    .A1(_09616_),
    .A2(_09617_));
 sg13g2_o21ai_1 _40208_ (.B1(net5652),
    .Y(_09620_),
    .A1(_09575_),
    .A2(_09583_));
 sg13g2_nand3b_1 _40209_ (.B(_09570_),
    .C(_09559_),
    .Y(_09621_),
    .A_N(_09620_));
 sg13g2_o21ai_1 _40210_ (.B1(net5652),
    .Y(_09622_),
    .A1(_09558_),
    .A2(_09568_));
 sg13g2_and2_1 _40211_ (.A(_09621_),
    .B(_09622_),
    .X(_09623_));
 sg13g2_and2_1 _40212_ (.A(_09619_),
    .B(_09623_),
    .X(_09624_));
 sg13g2_a21o_1 _40213_ (.A2(_09623_),
    .A1(_09619_),
    .B1(_09555_),
    .X(_09625_));
 sg13g2_o21ai_1 _40214_ (.B1(net5654),
    .Y(_09626_),
    .A1(_09544_),
    .A2(_09550_));
 sg13g2_inv_1 _40215_ (.Y(_09627_),
    .A(_09626_));
 sg13g2_a221oi_1 _40216_ (.B2(_09627_),
    .C1(_09539_),
    .B1(_09541_),
    .A1(net5656),
    .Y(_09628_),
    .A2(_09531_));
 sg13g2_o21ai_1 _40217_ (.B1(net5654),
    .Y(_09629_),
    .A1(_09515_),
    .A2(_09522_));
 sg13g2_o21ai_1 _40218_ (.B1(net5654),
    .Y(_09630_),
    .A1(_09501_),
    .A2(_09510_));
 sg13g2_o21ai_1 _40219_ (.B1(_09630_),
    .Y(_09631_),
    .A1(_09512_),
    .A2(_09629_));
 sg13g2_nand3_1 _40220_ (.B(_09554_),
    .C(_09631_),
    .A(_09541_),
    .Y(_09632_));
 sg13g2_and3_2 _40221_ (.X(_09633_),
    .A(_09625_),
    .B(_09628_),
    .C(_09632_));
 sg13g2_nand3_1 _40222_ (.B(_09628_),
    .C(_09632_),
    .A(_09625_),
    .Y(_09634_));
 sg13g2_o21ai_1 _40223_ (.B1(net5666),
    .Y(_09635_),
    .A1(_09427_),
    .A2(_09433_));
 sg13g2_inv_1 _40224_ (.Y(_09636_),
    .A(_09635_));
 sg13g2_nand2_1 _40225_ (.Y(_09637_),
    .A(_09417_),
    .B(_09422_));
 sg13g2_a21o_1 _40226_ (.A2(_09636_),
    .A1(_09424_),
    .B1(_09637_),
    .X(_09638_));
 sg13g2_inv_1 _40227_ (.Y(_09639_),
    .A(_09638_));
 sg13g2_nand2b_1 _40228_ (.Y(_09640_),
    .B(_09406_),
    .A_N(_09400_));
 sg13g2_a21o_1 _40229_ (.A2(_09394_),
    .A1(net5664),
    .B1(_09388_),
    .X(_09641_));
 sg13g2_a221oi_1 _40230_ (.B2(_09396_),
    .C1(_09641_),
    .B1(_09640_),
    .A1(_09410_),
    .Y(_09642_),
    .A2(_09638_));
 sg13g2_o21ai_1 _40231_ (.B1(net5656),
    .Y(_09643_),
    .A1(_09480_),
    .A2(_09487_));
 sg13g2_nor3_1 _40232_ (.A(_09471_),
    .B(_09477_),
    .C(_09643_),
    .Y(_09644_));
 sg13g2_nand2_1 _40233_ (.Y(_09645_),
    .A(_09469_),
    .B(_09475_));
 sg13g2_o21ai_1 _40234_ (.B1(_09461_),
    .Y(_09646_),
    .A1(_09644_),
    .A2(_09645_));
 sg13g2_o21ai_1 _40235_ (.B1(net5655),
    .Y(_09647_),
    .A1(_09455_),
    .A2(_09458_));
 sg13g2_or3_1 _40236_ (.A(_09447_),
    .B(_09452_),
    .C(_09647_),
    .X(_09648_));
 sg13g2_and4_1 _40237_ (.A(_09446_),
    .B(_09451_),
    .C(_09646_),
    .D(_09648_),
    .X(_09649_));
 sg13g2_nand4_1 _40238_ (.B(_09451_),
    .C(_09646_),
    .A(_09446_),
    .Y(_09650_),
    .D(_09648_));
 sg13g2_o21ai_1 _40239_ (.B1(_09642_),
    .Y(_09651_),
    .A1(_09437_),
    .A2(_09649_));
 sg13g2_a21oi_2 _40240_ (.B1(_09651_),
    .Y(_09652_),
    .A2(_09634_),
    .A1(_09494_));
 sg13g2_nand2b_1 _40241_ (.Y(_09653_),
    .B(net5603),
    .A_N(_08968_));
 sg13g2_nand2_1 _40242_ (.Y(_09654_),
    .A(_08969_),
    .B(_09653_));
 sg13g2_xnor2_1 _40243_ (.Y(_09655_),
    .A(net5675),
    .B(_08973_));
 sg13g2_nor3_1 _40244_ (.A(_08964_),
    .B(_09654_),
    .C(_09655_),
    .Y(_09656_));
 sg13g2_inv_1 _40245_ (.Y(_09657_),
    .A(_09656_));
 sg13g2_nand2_1 _40246_ (.Y(_09658_),
    .A(_08949_),
    .B(_09656_));
 sg13g2_or2_1 _40247_ (.X(_09659_),
    .B(_09658_),
    .A(_08920_));
 sg13g2_or2_1 _40248_ (.X(_09660_),
    .B(_09659_),
    .A(_09123_));
 sg13g2_a21o_2 _40249_ (.A2(_09652_),
    .A1(net1066),
    .B1(_09660_),
    .X(_09661_));
 sg13g2_nand2_2 _40250_ (.Y(_09662_),
    .A(_09124_),
    .B(_09661_));
 sg13g2_nand2_1 _40251_ (.Y(_09663_),
    .A(net6779),
    .B(_08208_));
 sg13g2_a21oi_2 _40252_ (.B1(_08512_),
    .Y(_09664_),
    .A2(net1098),
    .A1(_07358_));
 sg13g2_o21ai_1 _40253_ (.B1(_08335_),
    .Y(_09665_),
    .A1(_08529_),
    .A2(_09664_));
 sg13g2_nand2_1 _40254_ (.Y(_09666_),
    .A(_08543_),
    .B(_09665_));
 sg13g2_nand2_1 _40255_ (.Y(_09667_),
    .A(_08236_),
    .B(_09666_));
 sg13g2_a21oi_1 _40256_ (.A1(_08238_),
    .A2(_09666_),
    .Y(_09668_),
    .B1(_08530_));
 sg13g2_o21ai_1 _40257_ (.B1(_08215_),
    .Y(_09669_),
    .A1(_08217_),
    .A2(_09668_));
 sg13g2_xnor2_1 _40258_ (.Y(_09670_),
    .A(_08209_),
    .B(_09669_));
 sg13g2_o21ai_1 _40259_ (.B1(_09663_),
    .Y(_09671_),
    .A1(net6779),
    .A2(_09670_));
 sg13g2_inv_2 _40260_ (.Y(_09672_),
    .A(_09671_));
 sg13g2_nand2_1 _40261_ (.Y(_09673_),
    .A(net5670),
    .B(_09672_));
 sg13g2_xnor2_1 _40262_ (.Y(_09674_),
    .A(net5596),
    .B(_09671_));
 sg13g2_a21oi_1 _40263_ (.A1(_08543_),
    .A2(_09665_),
    .Y(_09675_),
    .B1(_08239_));
 sg13g2_o21ai_1 _40264_ (.B1(_08197_),
    .Y(_09676_),
    .A1(_08532_),
    .A2(_09675_));
 sg13g2_or3_1 _40265_ (.A(_08197_),
    .B(_08532_),
    .C(_09675_),
    .X(_09677_));
 sg13g2_nand3_1 _40266_ (.B(_09676_),
    .C(_09677_),
    .A(net6822),
    .Y(_09678_));
 sg13g2_o21ai_1 _40267_ (.B1(_09678_),
    .Y(_09679_),
    .A1(net6822),
    .A2(_08195_));
 sg13g2_xnor2_1 _40268_ (.Y(_09680_),
    .A(net5596),
    .B(_09679_));
 sg13g2_nor2b_1 _40269_ (.A(_09674_),
    .B_N(_09680_),
    .Y(_09681_));
 sg13g2_or2_1 _40270_ (.X(_09682_),
    .B(_08214_),
    .A(net6822));
 sg13g2_xnor2_1 _40271_ (.Y(_09683_),
    .A(_08217_),
    .B(_09668_));
 sg13g2_o21ai_1 _40272_ (.B1(_09682_),
    .Y(_09684_),
    .A1(net6779),
    .A2(_09683_));
 sg13g2_nand2b_1 _40273_ (.Y(_09685_),
    .B(net5596),
    .A_N(_09684_));
 sg13g2_xnor2_1 _40274_ (.Y(_09686_),
    .A(net5596),
    .B(_09684_));
 sg13g2_nand2_1 _40275_ (.Y(_09687_),
    .A(_08235_),
    .B(_09667_));
 sg13g2_nor2_1 _40276_ (.A(net6822),
    .B(_08227_),
    .Y(_09688_));
 sg13g2_xor2_1 _40277_ (.B(_09687_),
    .A(_08229_),
    .X(_09689_));
 sg13g2_a21oi_2 _40278_ (.B1(_09688_),
    .Y(_09690_),
    .A2(_09689_),
    .A1(net6824));
 sg13g2_and2_1 _40279_ (.A(net5670),
    .B(_09690_),
    .X(_09691_));
 sg13g2_xnor2_1 _40280_ (.Y(_09692_),
    .A(net5596),
    .B(_09690_));
 sg13g2_inv_1 _40281_ (.Y(_09693_),
    .A(_09692_));
 sg13g2_and3_2 _40282_ (.X(_09694_),
    .A(_09681_),
    .B(_09686_),
    .C(_09692_));
 sg13g2_o21ai_1 _40283_ (.B1(_08198_),
    .Y(_09695_),
    .A1(_08532_),
    .A2(_09675_));
 sg13g2_a21oi_1 _40284_ (.A1(_08533_),
    .A2(_09695_),
    .Y(_09696_),
    .B1(_08165_));
 sg13g2_a21oi_1 _40285_ (.A1(net5818),
    .A2(_08164_),
    .Y(_09697_),
    .B1(_09696_));
 sg13g2_xnor2_1 _40286_ (.Y(_09698_),
    .A(_08176_),
    .B(_09697_));
 sg13g2_a21oi_1 _40287_ (.A1(_08170_),
    .A2(_08173_),
    .Y(_09699_),
    .B1(net6822));
 sg13g2_a21o_2 _40288_ (.A2(_09698_),
    .A1(net6823),
    .B1(_09699_),
    .X(_09700_));
 sg13g2_nor2_1 _40289_ (.A(net5595),
    .B(_09700_),
    .Y(_09701_));
 sg13g2_xnor2_1 _40290_ (.Y(_09702_),
    .A(net5665),
    .B(_09700_));
 sg13g2_nand2_1 _40291_ (.Y(_09703_),
    .A(net6775),
    .B(_06789_));
 sg13g2_o21ai_1 _40292_ (.B1(_08548_),
    .Y(_09704_),
    .A1(net1086),
    .A2(_08545_));
 sg13g2_xor2_1 _40293_ (.B(_08548_),
    .A(_08546_),
    .X(_09705_));
 sg13g2_o21ai_1 _40294_ (.B1(_09703_),
    .Y(_09706_),
    .A1(net6775),
    .A2(_09705_));
 sg13g2_xnor2_1 _40295_ (.Y(_09707_),
    .A(net5607),
    .B(_09706_));
 sg13g2_and2_1 _40296_ (.A(_09702_),
    .B(_09707_),
    .X(_09708_));
 sg13g2_a21oi_1 _40297_ (.A1(_08182_),
    .A2(_08186_),
    .Y(_09709_),
    .B1(net6822));
 sg13g2_nand2_1 _40298_ (.Y(_09710_),
    .A(_08196_),
    .B(_09676_));
 sg13g2_xor2_1 _40299_ (.B(_09710_),
    .A(_08189_),
    .X(_09711_));
 sg13g2_a21oi_2 _40300_ (.B1(_09709_),
    .Y(_09712_),
    .A2(_09711_),
    .A1(net6823));
 sg13g2_nand2_1 _40301_ (.Y(_09713_),
    .A(net5665),
    .B(_09712_));
 sg13g2_xnor2_1 _40302_ (.Y(_09714_),
    .A(net5665),
    .B(_09712_));
 sg13g2_and3_1 _40303_ (.X(_09715_),
    .A(_08165_),
    .B(_08533_),
    .C(_09695_));
 sg13g2_nor3_1 _40304_ (.A(net6775),
    .B(_09696_),
    .C(_09715_),
    .Y(_09716_));
 sg13g2_a21o_2 _40305_ (.A2(_08164_),
    .A1(net6777),
    .B1(_09716_),
    .X(_09717_));
 sg13g2_nand2_1 _40306_ (.Y(_09718_),
    .A(net5665),
    .B(_09717_));
 sg13g2_xnor2_1 _40307_ (.Y(_09719_),
    .A(net5595),
    .B(_09717_));
 sg13g2_nor2b_1 _40308_ (.A(_09714_),
    .B_N(_09719_),
    .Y(_09720_));
 sg13g2_and3_2 _40309_ (.X(_09721_),
    .A(_09702_),
    .B(_09707_),
    .C(_09720_));
 sg13g2_nand2_1 _40310_ (.Y(_09722_),
    .A(net6779),
    .B(_08234_));
 sg13g2_xnor2_1 _40311_ (.Y(_09723_),
    .A(_08236_),
    .B(_09666_));
 sg13g2_o21ai_1 _40312_ (.B1(_09722_),
    .Y(_09724_),
    .A1(net6779),
    .A2(_09723_));
 sg13g2_xnor2_1 _40313_ (.Y(_09725_),
    .A(net5597),
    .B(_09724_));
 sg13g2_inv_1 _40314_ (.Y(_09726_),
    .A(_09725_));
 sg13g2_o21ai_1 _40315_ (.B1(_08334_),
    .Y(_09727_),
    .A1(_08529_),
    .A2(_09664_));
 sg13g2_a21oi_1 _40316_ (.A1(_08539_),
    .A2(_09727_),
    .Y(_09728_),
    .B1(_08294_));
 sg13g2_nor2_1 _40317_ (.A(_08293_),
    .B(_09728_),
    .Y(_09729_));
 sg13g2_a221oi_1 _40318_ (.B2(_09727_),
    .C1(_08294_),
    .B1(_08539_),
    .A1(_08285_),
    .Y(_09730_),
    .A2(_08286_));
 sg13g2_o21ai_1 _40319_ (.B1(_08258_),
    .Y(_09731_),
    .A1(_08541_),
    .A2(_09730_));
 sg13g2_nand2_1 _40320_ (.Y(_09732_),
    .A(_08256_),
    .B(_09731_));
 sg13g2_xor2_1 _40321_ (.B(_09732_),
    .A(_08270_),
    .X(_09733_));
 sg13g2_nor2_1 _40322_ (.A(net6824),
    .B(_08267_),
    .Y(_09734_));
 sg13g2_a21oi_1 _40323_ (.A1(net6824),
    .A2(_09733_),
    .Y(_09735_),
    .B1(_09734_));
 sg13g2_inv_2 _40324_ (.Y(_09736_),
    .A(_09735_));
 sg13g2_nand2_1 _40325_ (.Y(_09737_),
    .A(net5670),
    .B(_09736_));
 sg13g2_xnor2_1 _40326_ (.Y(_09738_),
    .A(net5596),
    .B(_09735_));
 sg13g2_or2_1 _40327_ (.X(_09739_),
    .B(_09738_),
    .A(_09726_));
 sg13g2_nor2_1 _40328_ (.A(net6824),
    .B(_08282_),
    .Y(_09740_));
 sg13g2_xnor2_1 _40329_ (.Y(_09741_),
    .A(_08287_),
    .B(_09729_));
 sg13g2_a21oi_2 _40330_ (.B1(_09740_),
    .Y(_09742_),
    .A2(_09741_),
    .A1(net6824));
 sg13g2_and2_1 _40331_ (.A(net5670),
    .B(_09742_),
    .X(_09743_));
 sg13g2_xnor2_1 _40332_ (.Y(_09744_),
    .A(net5670),
    .B(_09742_));
 sg13g2_nor2_1 _40333_ (.A(net6824),
    .B(_08255_),
    .Y(_09745_));
 sg13g2_or3_1 _40334_ (.A(_08258_),
    .B(_08541_),
    .C(_09730_),
    .X(_09746_));
 sg13g2_nand3_1 _40335_ (.B(_09731_),
    .C(_09746_),
    .A(net6824),
    .Y(_09747_));
 sg13g2_nor2b_2 _40336_ (.A(_09745_),
    .B_N(_09747_),
    .Y(_09748_));
 sg13g2_nor2_1 _40337_ (.A(net5596),
    .B(_09748_),
    .Y(_09749_));
 sg13g2_nand2_1 _40338_ (.Y(_09750_),
    .A(net5596),
    .B(_09748_));
 sg13g2_nand2b_2 _40339_ (.Y(_09751_),
    .B(_09750_),
    .A_N(_09749_));
 sg13g2_nand3_1 _40340_ (.B(_08539_),
    .C(_09727_),
    .A(_08294_),
    .Y(_09752_));
 sg13g2_nand3b_1 _40341_ (.B(_09752_),
    .C(net6827),
    .Y(_09753_),
    .A_N(_09728_));
 sg13g2_o21ai_1 _40342_ (.B1(_09753_),
    .Y(_09754_),
    .A1(net6824),
    .A2(_08292_));
 sg13g2_xnor2_1 _40343_ (.Y(_09755_),
    .A(net5597),
    .B(_09754_));
 sg13g2_o21ai_1 _40344_ (.B1(_08333_),
    .Y(_09756_),
    .A1(_08529_),
    .A2(_09664_));
 sg13g2_nand2_1 _40345_ (.Y(_09757_),
    .A(_08331_),
    .B(_09756_));
 sg13g2_o21ai_1 _40346_ (.B1(_08537_),
    .Y(_09758_),
    .A1(_08325_),
    .A2(_09756_));
 sg13g2_a21oi_1 _40347_ (.A1(_08306_),
    .A2(_09758_),
    .Y(_09759_),
    .B1(_08305_));
 sg13g2_and2_1 _40348_ (.A(net6779),
    .B(_08314_),
    .X(_09760_));
 sg13g2_xnor2_1 _40349_ (.Y(_09761_),
    .A(_08316_),
    .B(_09759_));
 sg13g2_a21oi_2 _40350_ (.B1(_09760_),
    .Y(_09762_),
    .A2(_09761_),
    .A1(net6826));
 sg13g2_and2_1 _40351_ (.A(net5669),
    .B(_09762_),
    .X(_09763_));
 sg13g2_xnor2_1 _40352_ (.Y(_09764_),
    .A(net5597),
    .B(_09762_));
 sg13g2_a21oi_1 _40353_ (.A1(_08306_),
    .A2(_09758_),
    .Y(_09765_),
    .B1(net6780));
 sg13g2_o21ai_1 _40354_ (.B1(_09765_),
    .Y(_09766_),
    .A1(_08306_),
    .A2(_09758_));
 sg13g2_o21ai_1 _40355_ (.B1(_09766_),
    .Y(_09767_),
    .A1(net6826),
    .A2(_08304_));
 sg13g2_nor2_1 _40356_ (.A(net5669),
    .B(_09767_),
    .Y(_09768_));
 sg13g2_xnor2_1 _40357_ (.Y(_09769_),
    .A(net5598),
    .B(_09767_));
 sg13g2_nor2_1 _40358_ (.A(net6826),
    .B(_08324_),
    .Y(_09770_));
 sg13g2_xor2_1 _40359_ (.B(_09757_),
    .A(_08325_),
    .X(_09771_));
 sg13g2_a21oi_2 _40360_ (.B1(_09770_),
    .Y(_09772_),
    .A2(_09771_),
    .A1(net6831));
 sg13g2_nand2_1 _40361_ (.Y(_09773_),
    .A(net5669),
    .B(_09772_));
 sg13g2_xnor2_1 _40362_ (.Y(_09774_),
    .A(net5669),
    .B(_09772_));
 sg13g2_inv_1 _40363_ (.Y(_09775_),
    .A(_09774_));
 sg13g2_nand4_1 _40364_ (.B(_09764_),
    .C(_09769_),
    .A(_09755_),
    .Y(_09776_),
    .D(_09775_));
 sg13g2_inv_1 _40365_ (.Y(_09777_),
    .A(_09776_));
 sg13g2_nor4_1 _40366_ (.A(_09739_),
    .B(_09744_),
    .C(_09751_),
    .D(_09776_),
    .Y(_09778_));
 sg13g2_nand3_1 _40367_ (.B(_09721_),
    .C(_09778_),
    .A(_09694_),
    .Y(_09779_));
 sg13g2_nand2_1 _40368_ (.Y(_09780_),
    .A(net6784),
    .B(_08421_));
 sg13g2_a21oi_1 _40369_ (.A1(_07358_),
    .A2(net1097),
    .Y(_09781_),
    .B1(_08509_));
 sg13g2_a21oi_2 _40370_ (.B1(_08520_),
    .Y(_09782_),
    .A2(_09781_),
    .A1(_08490_));
 sg13g2_o21ai_1 _40371_ (.B1(_08517_),
    .Y(_09783_),
    .A1(_08469_),
    .A2(_09782_));
 sg13g2_a21oi_1 _40372_ (.A1(_08379_),
    .A2(_09783_),
    .Y(_09784_),
    .B1(_08527_));
 sg13g2_a21o_1 _40373_ (.A2(_09783_),
    .A1(_08379_),
    .B1(_08527_),
    .X(_09785_));
 sg13g2_xnor2_1 _40374_ (.Y(_09786_),
    .A(_08423_),
    .B(_09784_));
 sg13g2_o21ai_1 _40375_ (.B1(_09780_),
    .Y(_09787_),
    .A1(net6784),
    .A2(_09786_));
 sg13g2_xnor2_1 _40376_ (.Y(_09788_),
    .A(net5604),
    .B(_09787_));
 sg13g2_a21oi_1 _40377_ (.A1(_08377_),
    .A2(_09783_),
    .Y(_09789_),
    .B1(_08376_));
 sg13g2_nand3_1 _40378_ (.B(_08377_),
    .C(_09783_),
    .A(_08370_),
    .Y(_09790_));
 sg13g2_a21o_1 _40379_ (.A2(_09790_),
    .A1(_08524_),
    .B1(_08353_),
    .X(_09791_));
 sg13g2_and3_1 _40380_ (.X(_09792_),
    .A(_08352_),
    .B(_08362_),
    .C(_09791_));
 sg13g2_a21oi_1 _40381_ (.A1(_08352_),
    .A2(_09791_),
    .Y(_09793_),
    .B1(_08362_));
 sg13g2_nand3_1 _40382_ (.B(_08356_),
    .C(_08360_),
    .A(net6784),
    .Y(_09794_));
 sg13g2_inv_1 _40383_ (.Y(_09795_),
    .A(_09794_));
 sg13g2_nor3_1 _40384_ (.A(net6784),
    .B(_09792_),
    .C(_09793_),
    .Y(_09796_));
 sg13g2_or2_1 _40385_ (.X(_09797_),
    .B(_09796_),
    .A(_09795_));
 sg13g2_o21ai_1 _40386_ (.B1(net5677),
    .Y(_09798_),
    .A1(_09795_),
    .A2(_09796_));
 sg13g2_or3_1 _40387_ (.A(net5677),
    .B(_09795_),
    .C(_09796_),
    .X(_09799_));
 sg13g2_nand2_1 _40388_ (.Y(_09800_),
    .A(_09798_),
    .B(_09799_));
 sg13g2_nand3_1 _40389_ (.B(_09798_),
    .C(_09799_),
    .A(_09788_),
    .Y(_09801_));
 sg13g2_nand3_1 _40390_ (.B(_08524_),
    .C(_09790_),
    .A(_08353_),
    .Y(_09802_));
 sg13g2_a21o_1 _40391_ (.A2(_09802_),
    .A1(_09791_),
    .B1(net6784),
    .X(_09803_));
 sg13g2_nand2_1 _40392_ (.Y(_09804_),
    .A(net6784),
    .B(_08351_));
 sg13g2_nand2_1 _40393_ (.Y(_09805_),
    .A(_09803_),
    .B(_09804_));
 sg13g2_inv_1 _40394_ (.Y(_09806_),
    .A(_09805_));
 sg13g2_and3_2 _40395_ (.X(_09807_),
    .A(net5677),
    .B(_09803_),
    .C(_09804_));
 sg13g2_a21oi_1 _40396_ (.A1(_09803_),
    .A2(_09804_),
    .Y(_09808_),
    .B1(net5677));
 sg13g2_nand2_1 _40397_ (.Y(_09809_),
    .A(net5604),
    .B(_09805_));
 sg13g2_or2_1 _40398_ (.X(_09810_),
    .B(_09808_),
    .A(_09807_));
 sg13g2_xor2_1 _40399_ (.B(_09789_),
    .A(_08370_),
    .X(_09811_));
 sg13g2_nand2_1 _40400_ (.Y(_09812_),
    .A(net6786),
    .B(_08369_));
 sg13g2_o21ai_1 _40401_ (.B1(_09812_),
    .Y(_09813_),
    .A1(net6784),
    .A2(_09811_));
 sg13g2_nand2_1 _40402_ (.Y(_09814_),
    .A(net5677),
    .B(_09813_));
 sg13g2_xnor2_1 _40403_ (.Y(_09815_),
    .A(net5677),
    .B(_09813_));
 sg13g2_nor3_1 _40404_ (.A(_09807_),
    .B(_09808_),
    .C(_09815_),
    .Y(_09816_));
 sg13g2_nand4_1 _40405_ (.B(_09798_),
    .C(_09799_),
    .A(_09788_),
    .Y(_09817_),
    .D(_09816_));
 sg13g2_nor3_1 _40406_ (.A(_08333_),
    .B(_08529_),
    .C(_09664_),
    .Y(_09818_));
 sg13g2_nand2_1 _40407_ (.Y(_09819_),
    .A(net6831),
    .B(_09756_));
 sg13g2_nor2_1 _40408_ (.A(_09818_),
    .B(_09819_),
    .Y(_09820_));
 sg13g2_a21oi_2 _40409_ (.B1(_09820_),
    .Y(_09821_),
    .A2(_08330_),
    .A1(net6783));
 sg13g2_nor2_1 _40410_ (.A(net5605),
    .B(_09821_),
    .Y(_09822_));
 sg13g2_xnor2_1 _40411_ (.Y(_09823_),
    .A(net5605),
    .B(_09821_));
 sg13g2_nor2_1 _40412_ (.A(net6833),
    .B(_08403_),
    .Y(_09824_));
 sg13g2_a21oi_1 _40413_ (.A1(_08424_),
    .A2(_09785_),
    .Y(_09825_),
    .B1(_08522_));
 sg13g2_o21ai_1 _40414_ (.B1(_08393_),
    .Y(_09826_),
    .A1(_08395_),
    .A2(_09825_));
 sg13g2_xnor2_1 _40415_ (.Y(_09827_),
    .A(_08405_),
    .B(_09826_));
 sg13g2_a21oi_2 _40416_ (.B1(_09824_),
    .Y(_09828_),
    .A2(_09827_),
    .A1(net6834));
 sg13g2_and2_1 _40417_ (.A(net5678),
    .B(_09828_),
    .X(_09829_));
 sg13g2_xnor2_1 _40418_ (.Y(_09830_),
    .A(net5678),
    .B(_09828_));
 sg13g2_nor2_1 _40419_ (.A(net6833),
    .B(_08392_),
    .Y(_09831_));
 sg13g2_xnor2_1 _40420_ (.Y(_09832_),
    .A(_08394_),
    .B(_09825_));
 sg13g2_a21oi_2 _40421_ (.B1(_09831_),
    .Y(_09833_),
    .A2(_09832_),
    .A1(net6833));
 sg13g2_nor2_1 _40422_ (.A(net5604),
    .B(_09833_),
    .Y(_09834_));
 sg13g2_xnor2_1 _40423_ (.Y(_09835_),
    .A(net5604),
    .B(_09833_));
 sg13g2_o21ai_1 _40424_ (.B1(_08422_),
    .Y(_09836_),
    .A1(_08423_),
    .A2(_09784_));
 sg13g2_nor2_1 _40425_ (.A(net6833),
    .B(_08414_),
    .Y(_09837_));
 sg13g2_xor2_1 _40426_ (.B(_09836_),
    .A(_08416_),
    .X(_09838_));
 sg13g2_a21oi_2 _40427_ (.B1(_09837_),
    .Y(_09839_),
    .A2(_09838_),
    .A1(net6833));
 sg13g2_and2_1 _40428_ (.A(net5677),
    .B(_09839_),
    .X(_09840_));
 sg13g2_xnor2_1 _40429_ (.Y(_09841_),
    .A(net5677),
    .B(_09839_));
 sg13g2_inv_1 _40430_ (.Y(_09842_),
    .A(_09841_));
 sg13g2_or2_1 _40431_ (.X(_09843_),
    .B(_09841_),
    .A(_09835_));
 sg13g2_nor3_1 _40432_ (.A(_09823_),
    .B(_09830_),
    .C(_09843_),
    .Y(_09844_));
 sg13g2_nor4_1 _40433_ (.A(_09817_),
    .B(_09823_),
    .C(_09830_),
    .D(_09843_),
    .Y(_09845_));
 sg13g2_nor2_1 _40434_ (.A(net6833),
    .B(_08375_),
    .Y(_09846_));
 sg13g2_xnor2_1 _40435_ (.Y(_09847_),
    .A(_08377_),
    .B(_09783_));
 sg13g2_a21oi_2 _40436_ (.B1(_09846_),
    .Y(_09848_),
    .A2(_09847_),
    .A1(net6833));
 sg13g2_xnor2_1 _40437_ (.Y(_09849_),
    .A(net5601),
    .B(_09848_));
 sg13g2_and2_1 _40438_ (.A(net6782),
    .B(_08450_),
    .X(_09850_));
 sg13g2_o21ai_1 _40439_ (.B1(_08466_),
    .Y(_09851_),
    .A1(_08467_),
    .A2(_09782_));
 sg13g2_nor3_1 _40440_ (.A(_08460_),
    .B(_08467_),
    .C(_09782_),
    .Y(_09852_));
 sg13g2_o21ai_1 _40441_ (.B1(_08442_),
    .Y(_09853_),
    .A1(_08515_),
    .A2(_09852_));
 sg13g2_nand2_1 _40442_ (.Y(_09854_),
    .A(_08440_),
    .B(_09853_));
 sg13g2_xnor2_1 _40443_ (.Y(_09855_),
    .A(_08452_),
    .B(_09854_));
 sg13g2_a21oi_1 _40444_ (.A1(net6831),
    .A2(_09855_),
    .Y(_09856_),
    .B1(_09850_));
 sg13g2_inv_1 _40445_ (.Y(_09857_),
    .A(_09856_));
 sg13g2_nor2_1 _40446_ (.A(net5602),
    .B(_09856_),
    .Y(_09858_));
 sg13g2_xnor2_1 _40447_ (.Y(_09859_),
    .A(net5676),
    .B(_09856_));
 sg13g2_nand2_1 _40448_ (.Y(_09860_),
    .A(net6782),
    .B(_08439_));
 sg13g2_nor3_1 _40449_ (.A(_08442_),
    .B(_08515_),
    .C(_09852_),
    .Y(_09861_));
 sg13g2_nand2_1 _40450_ (.Y(_09862_),
    .A(net6831),
    .B(_09853_));
 sg13g2_o21ai_1 _40451_ (.B1(_09860_),
    .Y(_09863_),
    .A1(_09861_),
    .A2(_09862_));
 sg13g2_and2_1 _40452_ (.A(net5676),
    .B(_09863_),
    .X(_09864_));
 sg13g2_nand2b_1 _40453_ (.Y(_09865_),
    .B(net5602),
    .A_N(_09863_));
 sg13g2_xnor2_1 _40454_ (.Y(_09866_),
    .A(net5602),
    .B(_09863_));
 sg13g2_xnor2_1 _40455_ (.Y(_09867_),
    .A(_08460_),
    .B(_09851_));
 sg13g2_nor2_1 _40456_ (.A(net6782),
    .B(_09867_),
    .Y(_09868_));
 sg13g2_a21oi_2 _40457_ (.B1(_09868_),
    .Y(_09869_),
    .A2(_08459_),
    .A1(net6782));
 sg13g2_nand2_1 _40458_ (.Y(_09870_),
    .A(net5676),
    .B(_09869_));
 sg13g2_xnor2_1 _40459_ (.Y(_09871_),
    .A(net5602),
    .B(_09869_));
 sg13g2_inv_1 _40460_ (.Y(_09872_),
    .A(_09871_));
 sg13g2_and2_1 _40461_ (.A(_09866_),
    .B(_09871_),
    .X(_09873_));
 sg13g2_nor2_1 _40462_ (.A(_08518_),
    .B(_09781_),
    .Y(_09874_));
 sg13g2_o21ai_1 _40463_ (.B1(_08487_),
    .Y(_09875_),
    .A1(_08489_),
    .A2(_09874_));
 sg13g2_nand2_1 _40464_ (.Y(_09876_),
    .A(net6783),
    .B(_08480_));
 sg13g2_xnor2_1 _40465_ (.Y(_09877_),
    .A(_08481_),
    .B(_09875_));
 sg13g2_o21ai_1 _40466_ (.B1(_09876_),
    .Y(_09878_),
    .A1(net6782),
    .A2(_09877_));
 sg13g2_inv_1 _40467_ (.Y(_09879_),
    .A(_09878_));
 sg13g2_nor2_1 _40468_ (.A(net5601),
    .B(_09878_),
    .Y(_09880_));
 sg13g2_nand2_1 _40469_ (.Y(_09881_),
    .A(net5601),
    .B(_09878_));
 sg13g2_xnor2_1 _40470_ (.Y(_09882_),
    .A(net5601),
    .B(_09878_));
 sg13g2_or2_1 _40471_ (.X(_09883_),
    .B(_08465_),
    .A(net6832));
 sg13g2_xnor2_1 _40472_ (.Y(_09884_),
    .A(_08467_),
    .B(_09782_));
 sg13g2_o21ai_1 _40473_ (.B1(_09883_),
    .Y(_09885_),
    .A1(net6782),
    .A2(_09884_));
 sg13g2_xnor2_1 _40474_ (.Y(_09886_),
    .A(net5601),
    .B(_09885_));
 sg13g2_nand2b_1 _40475_ (.Y(_09887_),
    .B(_09886_),
    .A_N(_09882_));
 sg13g2_xnor2_1 _40476_ (.Y(_09888_),
    .A(_08488_),
    .B(_09874_));
 sg13g2_nor2_1 _40477_ (.A(net6782),
    .B(_09888_),
    .Y(_09889_));
 sg13g2_a21oi_2 _40478_ (.B1(_09889_),
    .Y(_09890_),
    .A2(_08486_),
    .A1(net6782));
 sg13g2_inv_1 _40479_ (.Y(_09891_),
    .A(_09890_));
 sg13g2_xnor2_1 _40480_ (.Y(_09892_),
    .A(net5601),
    .B(_09890_));
 sg13g2_nor2_1 _40481_ (.A(net6831),
    .B(_08506_),
    .Y(_09893_));
 sg13g2_a21oi_1 _40482_ (.A1(_08139_),
    .A2(_08497_),
    .Y(_09894_),
    .B1(_08496_));
 sg13g2_xnor2_1 _40483_ (.Y(_09895_),
    .A(_08507_),
    .B(_09894_));
 sg13g2_a21oi_2 _40484_ (.B1(_09893_),
    .Y(_09896_),
    .A2(_09895_),
    .A1(net6831));
 sg13g2_nand2_1 _40485_ (.Y(_09897_),
    .A(net5676),
    .B(_09896_));
 sg13g2_xnor2_1 _40486_ (.Y(_09898_),
    .A(net5601),
    .B(_09896_));
 sg13g2_xnor2_1 _40487_ (.Y(_09899_),
    .A(net5676),
    .B(_09896_));
 sg13g2_nand2_1 _40488_ (.Y(_09900_),
    .A(_09892_),
    .B(_09898_));
 sg13g2_nor2_1 _40489_ (.A(_09887_),
    .B(_09900_),
    .Y(_09901_));
 sg13g2_and4_1 _40490_ (.A(_09849_),
    .B(_09859_),
    .C(_09873_),
    .D(_09901_),
    .X(_09902_));
 sg13g2_and2_1 _40491_ (.A(_09845_),
    .B(_09902_),
    .X(_09903_));
 sg13g2_inv_1 _40492_ (.Y(_09904_),
    .A(_09903_));
 sg13g2_nand2b_1 _40493_ (.Y(_09905_),
    .B(_09903_),
    .A_N(_09779_));
 sg13g2_a21oi_2 _40494_ (.B1(_09905_),
    .Y(_09906_),
    .A2(_09661_),
    .A1(_09124_));
 sg13g2_a21o_2 _40495_ (.A2(_09661_),
    .A1(_09124_),
    .B1(_09905_),
    .X(_09907_));
 sg13g2_o21ai_1 _40496_ (.B1(net5676),
    .Y(_09908_),
    .A1(_09890_),
    .A2(_09896_));
 sg13g2_a21oi_1 _40497_ (.A1(net5676),
    .A2(_09885_),
    .Y(_09909_),
    .B1(_09880_));
 sg13g2_o21ai_1 _40498_ (.B1(_09909_),
    .Y(_09910_),
    .A1(_09887_),
    .A2(_09908_));
 sg13g2_nand4_1 _40499_ (.B(_09859_),
    .C(_09873_),
    .A(_09849_),
    .Y(_09911_),
    .D(_09910_));
 sg13g2_nand2b_1 _40500_ (.Y(_09912_),
    .B(_09870_),
    .A_N(_09864_));
 sg13g2_nand3_1 _40501_ (.B(_09859_),
    .C(_09912_),
    .A(_09849_),
    .Y(_09913_));
 sg13g2_a21oi_1 _40502_ (.A1(net5676),
    .A2(_09848_),
    .Y(_09914_),
    .B1(_09858_));
 sg13g2_nand3_1 _40503_ (.B(_09913_),
    .C(_09914_),
    .A(_09911_),
    .Y(_09915_));
 sg13g2_nor2_1 _40504_ (.A(_09834_),
    .B(_09840_),
    .Y(_09916_));
 sg13g2_nor3_1 _40505_ (.A(_09823_),
    .B(_09830_),
    .C(_09916_),
    .Y(_09917_));
 sg13g2_nor3_2 _40506_ (.A(_09822_),
    .B(_09829_),
    .C(_09917_),
    .Y(_09918_));
 sg13g2_nor2b_1 _40507_ (.A(_09807_),
    .B_N(_09814_),
    .Y(_09919_));
 sg13g2_nor2_1 _40508_ (.A(_09801_),
    .B(_09919_),
    .Y(_09920_));
 sg13g2_o21ai_1 _40509_ (.B1(net5678),
    .Y(_09921_),
    .A1(_09787_),
    .A2(_09797_));
 sg13g2_nor2b_1 _40510_ (.A(_09920_),
    .B_N(_09921_),
    .Y(_09922_));
 sg13g2_o21ai_1 _40511_ (.B1(_09921_),
    .Y(_09923_),
    .A1(_09801_),
    .A2(_09919_));
 sg13g2_a22oi_1 _40512_ (.Y(_09924_),
    .B1(_09923_),
    .B2(_09844_),
    .A2(_09915_),
    .A1(_09845_));
 sg13g2_nand2_2 _40513_ (.Y(_09925_),
    .A(_09918_),
    .B(_09924_));
 sg13g2_a21o_2 _40514_ (.A2(_09924_),
    .A1(_09918_),
    .B1(_09779_),
    .X(_09926_));
 sg13g2_o21ai_1 _40515_ (.B1(net5669),
    .Y(_09927_),
    .A1(_09767_),
    .A2(_09772_));
 sg13g2_nand3b_1 _40516_ (.B(_09764_),
    .C(_09755_),
    .Y(_09928_),
    .A_N(_09927_));
 sg13g2_o21ai_1 _40517_ (.B1(net5669),
    .Y(_09929_),
    .A1(_09754_),
    .A2(_09762_));
 sg13g2_and2_1 _40518_ (.A(_09928_),
    .B(_09929_),
    .X(_09930_));
 sg13g2_nor4_1 _40519_ (.A(_09739_),
    .B(_09744_),
    .C(_09751_),
    .D(_09930_),
    .Y(_09931_));
 sg13g2_o21ai_1 _40520_ (.B1(net5670),
    .Y(_09932_),
    .A1(_09724_),
    .A2(_09736_));
 sg13g2_nor2_1 _40521_ (.A(_09743_),
    .B(_09749_),
    .Y(_09933_));
 sg13g2_or2_1 _40522_ (.X(_09934_),
    .B(_09749_),
    .A(_09743_));
 sg13g2_o21ai_1 _40523_ (.B1(_09932_),
    .Y(_09935_),
    .A1(_09739_),
    .A2(_09933_));
 sg13g2_nor2_2 _40524_ (.A(_09931_),
    .B(_09935_),
    .Y(_09936_));
 sg13g2_nand3b_1 _40525_ (.B(_09721_),
    .C(_09694_),
    .Y(_09937_),
    .A_N(_09936_));
 sg13g2_nand2_1 _40526_ (.Y(_09938_),
    .A(_09713_),
    .B(_09718_));
 sg13g2_a221oi_1 _40527_ (.B2(_09938_),
    .C1(_09701_),
    .B1(_09708_),
    .A1(net5665),
    .Y(_09939_),
    .A2(_09706_));
 sg13g2_a21o_1 _40528_ (.A2(_09684_),
    .A1(net5670),
    .B1(_09691_),
    .X(_09940_));
 sg13g2_a22oi_1 _40529_ (.Y(_09941_),
    .B1(_09681_),
    .B2(_09940_),
    .A2(_09679_),
    .A1(net5670));
 sg13g2_nand2_2 _40530_ (.Y(_09942_),
    .A(_09673_),
    .B(_09941_));
 sg13g2_nand2_1 _40531_ (.Y(_09943_),
    .A(_09721_),
    .B(_09942_));
 sg13g2_and4_1 _40532_ (.A(_09926_),
    .B(_09937_),
    .C(_09939_),
    .D(_09943_),
    .X(_09944_));
 sg13g2_nand4_1 _40533_ (.B(_09937_),
    .C(_09939_),
    .A(_09926_),
    .Y(_09945_),
    .D(_09943_));
 sg13g2_nand2_1 _40534_ (.Y(_09946_),
    .A(net6768),
    .B(_06644_));
 sg13g2_o21ai_1 _40535_ (.B1(_08553_),
    .Y(_09947_),
    .A1(net1086),
    .A2(_08545_));
 sg13g2_nand2_2 _40536_ (.Y(_09948_),
    .A(_06893_),
    .B(_09947_));
 sg13g2_a21oi_1 _40537_ (.A1(_06893_),
    .A2(_09947_),
    .Y(_09949_),
    .B1(_06614_));
 sg13g2_nor2_1 _40538_ (.A(_06909_),
    .B(_09949_),
    .Y(_09950_));
 sg13g2_o21ai_1 _40539_ (.B1(_06712_),
    .Y(_09951_),
    .A1(_06909_),
    .A2(_09949_));
 sg13g2_o21ai_1 _40540_ (.B1(_06898_),
    .Y(_09952_),
    .A1(_06693_),
    .A2(_09951_));
 sg13g2_a21oi_1 _40541_ (.A1(_06672_),
    .A2(_09952_),
    .Y(_09953_),
    .B1(_06899_));
 sg13g2_o21ai_1 _40542_ (.B1(_06633_),
    .Y(_09954_),
    .A1(_06635_),
    .A2(_09953_));
 sg13g2_xnor2_1 _40543_ (.Y(_09955_),
    .A(_06647_),
    .B(_09954_));
 sg13g2_o21ai_1 _40544_ (.B1(_09946_),
    .Y(_09956_),
    .A1(net6768),
    .A2(_09955_));
 sg13g2_inv_2 _40545_ (.Y(_09957_),
    .A(_09956_));
 sg13g2_nand2_1 _40546_ (.Y(_09958_),
    .A(net5642),
    .B(_09957_));
 sg13g2_xnor2_1 _40547_ (.Y(_09959_),
    .A(net5583),
    .B(_09956_));
 sg13g2_nor2_1 _40548_ (.A(net6807),
    .B(_06219_),
    .Y(_09960_));
 sg13g2_xnor2_1 _40549_ (.Y(_09961_),
    .A(_06221_),
    .B(_08587_));
 sg13g2_a21oi_2 _40550_ (.B1(_09960_),
    .Y(_09962_),
    .A2(_09961_),
    .A1(net6808));
 sg13g2_inv_1 _40551_ (.Y(_09963_),
    .A(_09962_));
 sg13g2_xnor2_1 _40552_ (.Y(_09964_),
    .A(net5582),
    .B(_09962_));
 sg13g2_nor2_1 _40553_ (.A(_09959_),
    .B(_09964_),
    .Y(_09965_));
 sg13g2_nor2_1 _40554_ (.A(net6810),
    .B(_06632_),
    .Y(_09966_));
 sg13g2_xnor2_1 _40555_ (.Y(_09967_),
    .A(_06634_),
    .B(_09953_));
 sg13g2_a21o_2 _40556_ (.A2(_09967_),
    .A1(net6810),
    .B1(_09966_),
    .X(_09968_));
 sg13g2_xnor2_1 _40557_ (.Y(_09969_),
    .A(net5583),
    .B(_09968_));
 sg13g2_nand2_1 _40558_ (.Y(_09970_),
    .A(net6768),
    .B(_06660_));
 sg13g2_a21oi_1 _40559_ (.A1(_06671_),
    .A2(_09952_),
    .Y(_09971_),
    .B1(_06669_));
 sg13g2_xor2_1 _40560_ (.B(_09971_),
    .A(_06661_),
    .X(_09972_));
 sg13g2_o21ai_1 _40561_ (.B1(_09970_),
    .Y(_09973_),
    .A1(net6768),
    .A2(_09972_));
 sg13g2_nor2_1 _40562_ (.A(net5583),
    .B(_09973_),
    .Y(_09974_));
 sg13g2_nand2_1 _40563_ (.Y(_09975_),
    .A(net5583),
    .B(_09973_));
 sg13g2_nand2b_1 _40564_ (.Y(_09976_),
    .B(_09975_),
    .A_N(_09974_));
 sg13g2_nand3b_1 _40565_ (.B(_09975_),
    .C(_09969_),
    .Y(_09977_),
    .A_N(_09974_));
 sg13g2_nor3_1 _40566_ (.A(_09959_),
    .B(_09964_),
    .C(_09977_),
    .Y(_09978_));
 sg13g2_nor2_1 _40567_ (.A(net6810),
    .B(_06684_),
    .Y(_09979_));
 sg13g2_a21o_1 _40568_ (.A2(_09951_),
    .A1(_06895_),
    .B1(_06692_),
    .X(_09980_));
 sg13g2_nand2_1 _40569_ (.Y(_09981_),
    .A(_06691_),
    .B(_09980_));
 sg13g2_xor2_1 _40570_ (.B(_09981_),
    .A(_06685_),
    .X(_09982_));
 sg13g2_a21oi_2 _40571_ (.B1(_09979_),
    .Y(_09983_),
    .A2(_09982_),
    .A1(net6811));
 sg13g2_and2_1 _40572_ (.A(net5650),
    .B(_09983_),
    .X(_09984_));
 sg13g2_xnor2_1 _40573_ (.Y(_09985_),
    .A(net5587),
    .B(_09983_));
 sg13g2_inv_1 _40574_ (.Y(_09986_),
    .A(_09985_));
 sg13g2_nor2_1 _40575_ (.A(net6810),
    .B(_06668_),
    .Y(_09987_));
 sg13g2_xnor2_1 _40576_ (.Y(_09988_),
    .A(_06670_),
    .B(_09952_));
 sg13g2_a21oi_1 _40577_ (.A1(net6810),
    .A2(_09988_),
    .Y(_09989_),
    .B1(_09987_));
 sg13g2_inv_2 _40578_ (.Y(_09990_),
    .A(_09989_));
 sg13g2_xnor2_1 _40579_ (.Y(_09991_),
    .A(net5650),
    .B(_09989_));
 sg13g2_nand2_1 _40580_ (.Y(_09992_),
    .A(_09985_),
    .B(_09991_));
 sg13g2_o21ai_1 _40581_ (.B1(_06700_),
    .Y(_09993_),
    .A1(_06702_),
    .A2(_09950_));
 sg13g2_xor2_1 _40582_ (.B(_09993_),
    .A(_06711_),
    .X(_09994_));
 sg13g2_nor2_1 _40583_ (.A(net6811),
    .B(_06709_),
    .Y(_09995_));
 sg13g2_a21oi_2 _40584_ (.B1(_09995_),
    .Y(_09996_),
    .A2(_09994_),
    .A1(net6810));
 sg13g2_inv_1 _40585_ (.Y(_09997_),
    .A(_09996_));
 sg13g2_xnor2_1 _40586_ (.Y(_09998_),
    .A(net5650),
    .B(_09996_));
 sg13g2_nand3_1 _40587_ (.B(_06895_),
    .C(_09951_),
    .A(_06692_),
    .Y(_09999_));
 sg13g2_and2_1 _40588_ (.A(net6811),
    .B(_09980_),
    .X(_10000_));
 sg13g2_a22oi_1 _40589_ (.Y(_10001_),
    .B1(_09999_),
    .B2(_10000_),
    .A2(_06690_),
    .A1(net6768));
 sg13g2_xnor2_1 _40590_ (.Y(_10002_),
    .A(net5587),
    .B(_10001_));
 sg13g2_inv_1 _40591_ (.Y(_10003_),
    .A(_10002_));
 sg13g2_nand4_1 _40592_ (.B(_09991_),
    .C(_09998_),
    .A(_09985_),
    .Y(_10004_),
    .D(_10003_));
 sg13g2_inv_1 _40593_ (.Y(_10005_),
    .A(_10004_));
 sg13g2_nor4_2 _40594_ (.A(_09959_),
    .B(_09964_),
    .C(_09977_),
    .Y(_10006_),
    .D(_10004_));
 sg13g2_nand2_1 _40595_ (.Y(_10007_),
    .A(_06611_),
    .B(_09948_));
 sg13g2_and3_1 _40596_ (.X(_10008_),
    .A(_06603_),
    .B(_06611_),
    .C(_09948_));
 sg13g2_a21oi_1 _40597_ (.A1(_06893_),
    .A2(_09947_),
    .Y(_10009_),
    .B1(_06612_));
 sg13g2_nor2_1 _40598_ (.A(_06904_),
    .B(_10009_),
    .Y(_10010_));
 sg13g2_o21ai_1 _40599_ (.B1(_06566_),
    .Y(_10011_),
    .A1(_06904_),
    .A2(_10009_));
 sg13g2_nand2_1 _40600_ (.Y(_10012_),
    .A(_06564_),
    .B(_10011_));
 sg13g2_o21ai_1 _40601_ (.B1(_06907_),
    .Y(_10013_),
    .A1(_06574_),
    .A2(_10011_));
 sg13g2_a21oi_1 _40602_ (.A1(_06555_),
    .A2(_10013_),
    .Y(_10014_),
    .B1(_06554_));
 sg13g2_xnor2_1 _40603_ (.Y(_10015_),
    .A(_06547_),
    .B(_10014_));
 sg13g2_mux2_1 _40604_ (.A0(_06546_),
    .A1(_10015_),
    .S(net6810),
    .X(_10016_));
 sg13g2_xnor2_1 _40605_ (.Y(_10017_),
    .A(net5648),
    .B(_10016_));
 sg13g2_nand2_1 _40606_ (.Y(_10018_),
    .A(net6768),
    .B(_06699_));
 sg13g2_xnor2_1 _40607_ (.Y(_10019_),
    .A(_06702_),
    .B(_09950_));
 sg13g2_o21ai_1 _40608_ (.B1(_10018_),
    .Y(_10020_),
    .A1(net6768),
    .A2(_10019_));
 sg13g2_xnor2_1 _40609_ (.Y(_10021_),
    .A(net5650),
    .B(_10020_));
 sg13g2_nor2_1 _40610_ (.A(net6810),
    .B(_06553_),
    .Y(_10022_));
 sg13g2_xor2_1 _40611_ (.B(_10013_),
    .A(_06555_),
    .X(_10023_));
 sg13g2_a21oi_2 _40612_ (.B1(_10022_),
    .Y(_10024_),
    .A2(_10023_),
    .A1(net6813));
 sg13g2_xnor2_1 _40613_ (.Y(_10025_),
    .A(net5587),
    .B(_10024_));
 sg13g2_xor2_1 _40614_ (.B(_10012_),
    .A(_06574_),
    .X(_10026_));
 sg13g2_nand2_1 _40615_ (.Y(_10027_),
    .A(net6812),
    .B(_10026_));
 sg13g2_o21ai_1 _40616_ (.B1(_10027_),
    .Y(_10028_),
    .A1(net6813),
    .A2(_06573_));
 sg13g2_inv_1 _40617_ (.Y(_10029_),
    .A(_10028_));
 sg13g2_xnor2_1 _40618_ (.Y(_10030_),
    .A(net5588),
    .B(_10028_));
 sg13g2_inv_1 _40619_ (.Y(_10031_),
    .A(_10030_));
 sg13g2_or4_1 _40620_ (.A(_10017_),
    .B(_10021_),
    .C(_10025_),
    .D(_10030_),
    .X(_10032_));
 sg13g2_inv_1 _40621_ (.Y(_10033_),
    .A(_10032_));
 sg13g2_nand2_1 _40622_ (.Y(_10034_),
    .A(net6769),
    .B(_06563_));
 sg13g2_xnor2_1 _40623_ (.Y(_10035_),
    .A(_06565_),
    .B(_10010_));
 sg13g2_o21ai_1 _40624_ (.B1(_10034_),
    .Y(_10036_),
    .A1(net6769),
    .A2(_10035_));
 sg13g2_xnor2_1 _40625_ (.Y(_10037_),
    .A(net5648),
    .B(_10036_));
 sg13g2_nor2_1 _40626_ (.A(net6812),
    .B(_06585_),
    .Y(_10038_));
 sg13g2_o21ai_1 _40627_ (.B1(_06594_),
    .Y(_10039_),
    .A1(_06902_),
    .A2(_10008_));
 sg13g2_nand2_1 _40628_ (.Y(_10040_),
    .A(_06593_),
    .B(_10039_));
 sg13g2_xnor2_1 _40629_ (.Y(_10041_),
    .A(_06587_),
    .B(_10040_));
 sg13g2_a21oi_2 _40630_ (.B1(_10038_),
    .Y(_10042_),
    .A2(_10041_),
    .A1(net6812));
 sg13g2_and2_1 _40631_ (.A(net5648),
    .B(_10042_),
    .X(_10043_));
 sg13g2_xnor2_1 _40632_ (.Y(_10044_),
    .A(net5648),
    .B(_10042_));
 sg13g2_nand2_1 _40633_ (.Y(_10045_),
    .A(net6768),
    .B(_06592_));
 sg13g2_nor3_1 _40634_ (.A(_06594_),
    .B(_06902_),
    .C(_10008_),
    .Y(_10046_));
 sg13g2_nand2_1 _40635_ (.Y(_10047_),
    .A(net6812),
    .B(_10039_));
 sg13g2_o21ai_1 _40636_ (.B1(_10045_),
    .Y(_10048_),
    .A1(_10046_),
    .A2(_10047_));
 sg13g2_inv_1 _40637_ (.Y(_10049_),
    .A(_10048_));
 sg13g2_nor2_1 _40638_ (.A(net5649),
    .B(_10048_),
    .Y(_10050_));
 sg13g2_xnor2_1 _40639_ (.Y(_10051_),
    .A(net5649),
    .B(_10048_));
 sg13g2_nor2_1 _40640_ (.A(net6812),
    .B(_06601_),
    .Y(_10052_));
 sg13g2_nand2_1 _40641_ (.Y(_10053_),
    .A(_06610_),
    .B(_10007_));
 sg13g2_xnor2_1 _40642_ (.Y(_10054_),
    .A(_06603_),
    .B(_10053_));
 sg13g2_a21oi_2 _40643_ (.B1(_10052_),
    .Y(_10055_),
    .A2(_10054_),
    .A1(net6812));
 sg13g2_nand2_1 _40644_ (.Y(_10056_),
    .A(net5648),
    .B(_10055_));
 sg13g2_xnor2_1 _40645_ (.Y(_10057_),
    .A(net5649),
    .B(_10055_));
 sg13g2_inv_1 _40646_ (.Y(_10058_),
    .A(_10057_));
 sg13g2_nor4_1 _40647_ (.A(_10037_),
    .B(_10044_),
    .C(_10051_),
    .D(_10057_),
    .Y(_10059_));
 sg13g2_inv_1 _40648_ (.Y(_10060_),
    .A(_10059_));
 sg13g2_nor2b_1 _40649_ (.A(_10032_),
    .B_N(_10059_),
    .Y(_10061_));
 sg13g2_inv_1 _40650_ (.Y(_10062_),
    .A(_10061_));
 sg13g2_nand2_1 _40651_ (.Y(_10063_),
    .A(_10006_),
    .B(_10061_));
 sg13g2_xnor2_1 _40652_ (.Y(_10064_),
    .A(_06611_),
    .B(_09948_));
 sg13g2_nand2_1 _40653_ (.Y(_10065_),
    .A(net6812),
    .B(_10064_));
 sg13g2_o21ai_1 _40654_ (.B1(_10065_),
    .Y(_10066_),
    .A1(net6812),
    .A2(_06609_));
 sg13g2_nor2_1 _40655_ (.A(net5592),
    .B(_10066_),
    .Y(_10067_));
 sg13g2_xnor2_1 _40656_ (.Y(_10068_),
    .A(net5658),
    .B(_10066_));
 sg13g2_inv_1 _40657_ (.Y(_10069_),
    .A(_10068_));
 sg13g2_nor2_1 _40658_ (.A(net6819),
    .B(_06821_),
    .Y(_10070_));
 sg13g2_o21ai_1 _40659_ (.B1(_08550_),
    .Y(_10071_),
    .A1(net1086),
    .A2(_08545_));
 sg13g2_o21ai_1 _40660_ (.B1(_06795_),
    .Y(_10072_),
    .A1(_08552_),
    .A2(_10071_));
 sg13g2_nand2_1 _40661_ (.Y(_10073_),
    .A(_06870_),
    .B(_10072_));
 sg13g2_nand4_1 _40662_ (.B(_06862_),
    .C(_06881_),
    .A(_06855_),
    .Y(_10074_),
    .D(_10072_));
 sg13g2_a21oi_1 _40663_ (.A1(_06887_),
    .A2(_10074_),
    .Y(_10075_),
    .B1(_06841_));
 sg13g2_a21oi_1 _40664_ (.A1(_06887_),
    .A2(_10074_),
    .Y(_10076_),
    .B1(_06843_));
 sg13g2_o21ai_1 _40665_ (.B1(_06813_),
    .Y(_10077_),
    .A1(_06889_),
    .A2(_10076_));
 sg13g2_nand2_1 _40666_ (.Y(_10078_),
    .A(_06812_),
    .B(_10077_));
 sg13g2_xnor2_1 _40667_ (.Y(_10079_),
    .A(_06823_),
    .B(_10078_));
 sg13g2_a21oi_2 _40668_ (.B1(_10070_),
    .Y(_10080_),
    .A2(_10079_),
    .A1(net6819));
 sg13g2_and2_1 _40669_ (.A(net5658),
    .B(_10080_),
    .X(_10081_));
 sg13g2_xnor2_1 _40670_ (.Y(_10082_),
    .A(net5592),
    .B(_10080_));
 sg13g2_xnor2_1 _40671_ (.Y(_10083_),
    .A(net5658),
    .B(_10080_));
 sg13g2_or3_1 _40672_ (.A(_06813_),
    .B(_06889_),
    .C(_10076_),
    .X(_10084_));
 sg13g2_and2_1 _40673_ (.A(net6819),
    .B(_10077_),
    .X(_10085_));
 sg13g2_a22oi_1 _40674_ (.Y(_10086_),
    .B1(_10084_),
    .B2(_10085_),
    .A2(_06811_),
    .A1(net6774));
 sg13g2_inv_1 _40675_ (.Y(_10087_),
    .A(_10086_));
 sg13g2_xnor2_1 _40676_ (.Y(_10088_),
    .A(net5592),
    .B(_10086_));
 sg13g2_a21oi_1 _40677_ (.A1(net5813),
    .A2(_06838_),
    .Y(_10089_),
    .B1(_10075_));
 sg13g2_xor2_1 _40678_ (.B(_10089_),
    .A(_06833_),
    .X(_10090_));
 sg13g2_nand2_1 _40679_ (.Y(_10091_),
    .A(net6774),
    .B(_06831_));
 sg13g2_o21ai_1 _40680_ (.B1(_10091_),
    .Y(_10092_),
    .A1(net6774),
    .A2(_10090_));
 sg13g2_nand2_1 _40681_ (.Y(_10093_),
    .A(net5658),
    .B(_10092_));
 sg13g2_xnor2_1 _40682_ (.Y(_10094_),
    .A(net5658),
    .B(_10092_));
 sg13g2_inv_1 _40683_ (.Y(_10095_),
    .A(_10094_));
 sg13g2_nor2_1 _40684_ (.A(_10088_),
    .B(_10094_),
    .Y(_10096_));
 sg13g2_nor4_1 _40685_ (.A(_10069_),
    .B(_10083_),
    .C(_10088_),
    .D(_10094_),
    .Y(_10097_));
 sg13g2_nand2_1 _40686_ (.Y(_10098_),
    .A(net6774),
    .B(_06853_));
 sg13g2_a21oi_1 _40687_ (.A1(_06881_),
    .A2(_10072_),
    .Y(_10099_),
    .B1(_06884_));
 sg13g2_o21ai_1 _40688_ (.B1(_06861_),
    .Y(_10100_),
    .A1(_06863_),
    .A2(_10099_));
 sg13g2_xnor2_1 _40689_ (.Y(_10101_),
    .A(_06855_),
    .B(_10100_));
 sg13g2_o21ai_1 _40690_ (.B1(_10098_),
    .Y(_10102_),
    .A1(net6774),
    .A2(_10101_));
 sg13g2_xnor2_1 _40691_ (.Y(_10103_),
    .A(net5658),
    .B(_10102_));
 sg13g2_nand2_1 _40692_ (.Y(_10104_),
    .A(net6774),
    .B(_06838_));
 sg13g2_nand3_1 _40693_ (.B(_06887_),
    .C(_10074_),
    .A(_06841_),
    .Y(_10105_));
 sg13g2_nand2b_1 _40694_ (.Y(_10106_),
    .B(_10105_),
    .A_N(_10075_));
 sg13g2_o21ai_1 _40695_ (.B1(_10104_),
    .Y(_10107_),
    .A1(net6774),
    .A2(_10106_));
 sg13g2_xnor2_1 _40696_ (.Y(_10108_),
    .A(net5592),
    .B(_10107_));
 sg13g2_nor2b_1 _40697_ (.A(_10103_),
    .B_N(_10108_),
    .Y(_10109_));
 sg13g2_nor2_1 _40698_ (.A(net6819),
    .B(_06860_),
    .Y(_10110_));
 sg13g2_xnor2_1 _40699_ (.Y(_10111_),
    .A(_06862_),
    .B(_10099_));
 sg13g2_a21oi_2 _40700_ (.B1(_10110_),
    .Y(_10112_),
    .A2(_10111_),
    .A1(net6819));
 sg13g2_inv_1 _40701_ (.Y(_10113_),
    .A(_10112_));
 sg13g2_xnor2_1 _40702_ (.Y(_10114_),
    .A(net5659),
    .B(_10112_));
 sg13g2_nor2_1 _40703_ (.A(net6819),
    .B(_06879_),
    .Y(_10115_));
 sg13g2_nand2_1 _40704_ (.Y(_10116_),
    .A(_06869_),
    .B(_10073_));
 sg13g2_xor2_1 _40705_ (.B(_10116_),
    .A(_06880_),
    .X(_10117_));
 sg13g2_a21oi_2 _40706_ (.B1(_10115_),
    .Y(_10118_),
    .A2(_10117_),
    .A1(net6818));
 sg13g2_nor2_1 _40707_ (.A(net5592),
    .B(_10118_),
    .Y(_10119_));
 sg13g2_xnor2_1 _40708_ (.Y(_10120_),
    .A(net5658),
    .B(_10118_));
 sg13g2_and3_1 _40709_ (.X(_10121_),
    .A(_10109_),
    .B(_10114_),
    .C(_10120_));
 sg13g2_inv_1 _40710_ (.Y(_10122_),
    .A(_10121_));
 sg13g2_and4_1 _40711_ (.A(_10068_),
    .B(_10082_),
    .C(_10096_),
    .D(_10121_),
    .X(_10123_));
 sg13g2_nor2_1 _40712_ (.A(net6818),
    .B(_06738_),
    .Y(_10124_));
 sg13g2_a21o_1 _40713_ (.A2(_10071_),
    .A1(_06793_),
    .B1(_06757_),
    .X(_10125_));
 sg13g2_a22oi_1 _40714_ (.Y(_10126_),
    .B1(_06756_),
    .B2(_10125_),
    .A2(_06755_),
    .A1(net5862));
 sg13g2_a21oi_1 _40715_ (.A1(_06729_),
    .A2(_10126_),
    .Y(_10127_),
    .B1(_06728_));
 sg13g2_xnor2_1 _40716_ (.Y(_10128_),
    .A(_06739_),
    .B(_10127_));
 sg13g2_a21oi_2 _40717_ (.B1(_10124_),
    .Y(_10129_),
    .A2(_10128_),
    .A1(net6818));
 sg13g2_and2_1 _40718_ (.A(net5660),
    .B(_10129_),
    .X(_10130_));
 sg13g2_nand2_1 _40719_ (.Y(_10131_),
    .A(net5660),
    .B(_10129_));
 sg13g2_xnor2_1 _40720_ (.Y(_10132_),
    .A(net5660),
    .B(_10129_));
 sg13g2_nand2_1 _40721_ (.Y(_10133_),
    .A(net6777),
    .B(_06868_));
 sg13g2_xnor2_1 _40722_ (.Y(_10134_),
    .A(_06870_),
    .B(_10072_));
 sg13g2_o21ai_1 _40723_ (.B1(_10133_),
    .Y(_10135_),
    .A1(net6774),
    .A2(_10134_));
 sg13g2_and2_1 _40724_ (.A(net5660),
    .B(_10135_),
    .X(_10136_));
 sg13g2_xnor2_1 _40725_ (.Y(_10137_),
    .A(net5660),
    .B(_10135_));
 sg13g2_nor2_1 _40726_ (.A(net6818),
    .B(_06727_),
    .Y(_10138_));
 sg13g2_xnor2_1 _40727_ (.Y(_10139_),
    .A(_06730_),
    .B(_10126_));
 sg13g2_a21oi_2 _40728_ (.B1(_10138_),
    .Y(_10140_),
    .A2(_10139_),
    .A1(net6818));
 sg13g2_nor2_1 _40729_ (.A(net5593),
    .B(_10140_),
    .Y(_10141_));
 sg13g2_nand2_1 _40730_ (.Y(_10142_),
    .A(net5593),
    .B(_10140_));
 sg13g2_xnor2_1 _40731_ (.Y(_10143_),
    .A(net5593),
    .B(_10140_));
 sg13g2_nor2_1 _40732_ (.A(net6818),
    .B(_06754_),
    .Y(_10144_));
 sg13g2_o21ai_1 _40733_ (.B1(_10125_),
    .Y(_10145_),
    .A1(net5862),
    .A2(_06745_));
 sg13g2_xor2_1 _40734_ (.B(_10145_),
    .A(_06758_),
    .X(_10146_));
 sg13g2_a21oi_2 _40735_ (.B1(_10144_),
    .Y(_10147_),
    .A2(_10146_),
    .A1(net6818));
 sg13g2_xnor2_1 _40736_ (.Y(_10148_),
    .A(net5660),
    .B(_10147_));
 sg13g2_or2_1 _40737_ (.X(_10149_),
    .B(_10148_),
    .A(_10143_));
 sg13g2_nor3_1 _40738_ (.A(_10132_),
    .B(_10137_),
    .C(_10149_),
    .Y(_10150_));
 sg13g2_nand2_1 _40739_ (.Y(_10151_),
    .A(_06790_),
    .B(_09704_));
 sg13g2_a22oi_1 _40740_ (.Y(_10152_),
    .B1(_06791_),
    .B2(_09704_),
    .A2(_06785_),
    .A1(net5866));
 sg13g2_a221oi_1 _40741_ (.B2(_09704_),
    .C1(_06777_),
    .B1(_06791_),
    .A1(net5866),
    .Y(_10153_),
    .A2(_06785_));
 sg13g2_or3_1 _40742_ (.A(_06769_),
    .B(_06775_),
    .C(_10153_),
    .X(_10154_));
 sg13g2_o21ai_1 _40743_ (.B1(_06769_),
    .Y(_10155_),
    .A1(_06775_),
    .A2(_10153_));
 sg13g2_nand2b_1 _40744_ (.Y(_10156_),
    .B(net6775),
    .A_N(_06767_));
 sg13g2_a21o_2 _40745_ (.A2(_10155_),
    .A1(_10154_),
    .B1(net6775),
    .X(_10157_));
 sg13g2_and2_1 _40746_ (.A(_10156_),
    .B(_10157_),
    .X(_10158_));
 sg13g2_inv_1 _40747_ (.Y(_10159_),
    .A(_10158_));
 sg13g2_a21oi_2 _40748_ (.B1(net5593),
    .Y(_10160_),
    .A2(_10157_),
    .A1(_10156_));
 sg13g2_and3_1 _40749_ (.X(_10161_),
    .A(net5593),
    .B(_10156_),
    .C(_10157_));
 sg13g2_nor2_1 _40750_ (.A(_10160_),
    .B(_10161_),
    .Y(_10162_));
 sg13g2_inv_2 _40751_ (.Y(_10163_),
    .A(_10162_));
 sg13g2_nand3_1 _40752_ (.B(_06793_),
    .C(_10071_),
    .A(_06757_),
    .Y(_10164_));
 sg13g2_nand3_1 _40753_ (.B(_10125_),
    .C(_10164_),
    .A(net6818),
    .Y(_10165_));
 sg13g2_o21ai_1 _40754_ (.B1(_10165_),
    .Y(_10166_),
    .A1(net6819),
    .A2(_06745_));
 sg13g2_xnor2_1 _40755_ (.Y(_10167_),
    .A(net5661),
    .B(_10166_));
 sg13g2_nand2_1 _40756_ (.Y(_10168_),
    .A(net6775),
    .B(_06774_));
 sg13g2_xnor2_1 _40757_ (.Y(_10169_),
    .A(_06776_),
    .B(_10152_));
 sg13g2_o21ai_1 _40758_ (.B1(_10168_),
    .Y(_10170_),
    .A1(net6775),
    .A2(_10169_));
 sg13g2_inv_1 _40759_ (.Y(_10171_),
    .A(_10170_));
 sg13g2_xnor2_1 _40760_ (.Y(_10172_),
    .A(net5661),
    .B(_10170_));
 sg13g2_nor2_1 _40761_ (.A(net6822),
    .B(_06784_),
    .Y(_10173_));
 sg13g2_xor2_1 _40762_ (.B(_10151_),
    .A(_08547_),
    .X(_10174_));
 sg13g2_a21oi_2 _40763_ (.B1(_10173_),
    .Y(_10175_),
    .A2(_10174_),
    .A1(net6822));
 sg13g2_nand2_1 _40764_ (.Y(_10176_),
    .A(net5664),
    .B(_10175_));
 sg13g2_xnor2_1 _40765_ (.Y(_10177_),
    .A(net5665),
    .B(_10175_));
 sg13g2_nor4_2 _40766_ (.A(_10163_),
    .B(_10167_),
    .C(_10172_),
    .Y(_10178_),
    .D(_10177_));
 sg13g2_and2_1 _40767_ (.A(_10150_),
    .B(_10178_),
    .X(_10179_));
 sg13g2_nand2_1 _40768_ (.Y(_10180_),
    .A(_10150_),
    .B(_10178_));
 sg13g2_and2_1 _40769_ (.A(_10123_),
    .B(_10179_),
    .X(_10181_));
 sg13g2_inv_1 _40770_ (.Y(_10182_),
    .A(_10181_));
 sg13g2_nor2b_1 _40771_ (.A(_10063_),
    .B_N(_10181_),
    .Y(_10183_));
 sg13g2_o21ai_1 _40772_ (.B1(_10183_),
    .Y(_10184_),
    .A1(_09945_),
    .A2(_09906_));
 sg13g2_o21ai_1 _40773_ (.B1(net5661),
    .Y(_10185_),
    .A1(_10170_),
    .A2(_10175_));
 sg13g2_nor4_1 _40774_ (.A(_10160_),
    .B(_10161_),
    .C(_10167_),
    .D(_10185_),
    .Y(_10186_));
 sg13g2_a21oi_1 _40775_ (.A1(net5661),
    .A2(_10166_),
    .Y(_10187_),
    .B1(_10160_));
 sg13g2_nor2b_2 _40776_ (.A(_10186_),
    .B_N(_10187_),
    .Y(_10188_));
 sg13g2_nor4_1 _40777_ (.A(_10132_),
    .B(_10137_),
    .C(_10149_),
    .D(_10188_),
    .Y(_10189_));
 sg13g2_a21oi_1 _40778_ (.A1(net5660),
    .A2(_10147_),
    .Y(_10190_),
    .B1(_10141_));
 sg13g2_inv_1 _40779_ (.Y(_10191_),
    .A(_10190_));
 sg13g2_nor3_1 _40780_ (.A(_10132_),
    .B(_10137_),
    .C(_10190_),
    .Y(_10192_));
 sg13g2_nor4_1 _40781_ (.A(_10130_),
    .B(_10136_),
    .C(_10189_),
    .D(_10192_),
    .Y(_10193_));
 sg13g2_inv_1 _40782_ (.Y(_10194_),
    .A(_10193_));
 sg13g2_o21ai_1 _40783_ (.B1(net5658),
    .Y(_10195_),
    .A1(_10087_),
    .A2(_10092_));
 sg13g2_nor3_1 _40784_ (.A(_10069_),
    .B(_10083_),
    .C(_10195_),
    .Y(_10196_));
 sg13g2_nor3_1 _40785_ (.A(_10067_),
    .B(_10081_),
    .C(_10196_),
    .Y(_10197_));
 sg13g2_a21oi_1 _40786_ (.A1(net5659),
    .A2(_10113_),
    .Y(_10198_),
    .B1(_10119_));
 sg13g2_nand2b_1 _40787_ (.Y(_10199_),
    .B(_10109_),
    .A_N(_10198_));
 sg13g2_o21ai_1 _40788_ (.B1(net5659),
    .Y(_10200_),
    .A1(_10102_),
    .A2(_10107_));
 sg13g2_nand2_1 _40789_ (.Y(_10201_),
    .A(_10199_),
    .B(_10200_));
 sg13g2_a22oi_1 _40790_ (.Y(_10202_),
    .B1(_10201_),
    .B2(_10097_),
    .A2(_10194_),
    .A1(_10123_));
 sg13g2_and2_1 _40791_ (.A(_10197_),
    .B(_10202_),
    .X(_10203_));
 sg13g2_nand2_1 _40792_ (.Y(_10204_),
    .A(_10197_),
    .B(_10202_));
 sg13g2_a21o_2 _40793_ (.A2(_10202_),
    .A1(_10197_),
    .B1(_10063_),
    .X(_10205_));
 sg13g2_o21ai_1 _40794_ (.B1(net5649),
    .Y(_10206_),
    .A1(_10048_),
    .A2(_10055_));
 sg13g2_nor3_1 _40795_ (.A(_10037_),
    .B(_10044_),
    .C(_10206_),
    .Y(_10207_));
 sg13g2_o21ai_1 _40796_ (.B1(net5648),
    .Y(_10208_),
    .A1(_10036_),
    .A2(_10042_));
 sg13g2_nand2b_1 _40797_ (.Y(_10209_),
    .B(_10208_),
    .A_N(_10207_));
 sg13g2_a21o_1 _40798_ (.A2(_10028_),
    .A1(_10024_),
    .B1(net5588),
    .X(_10210_));
 sg13g2_nor3_1 _40799_ (.A(_10017_),
    .B(_10021_),
    .C(_10210_),
    .Y(_10211_));
 sg13g2_o21ai_1 _40800_ (.B1(net5648),
    .Y(_10212_),
    .A1(_10016_),
    .A2(_10020_));
 sg13g2_nand2b_1 _40801_ (.Y(_10213_),
    .B(_10212_),
    .A_N(_10211_));
 sg13g2_a21o_2 _40802_ (.A2(_10209_),
    .A1(_10033_),
    .B1(_10213_),
    .X(_10214_));
 sg13g2_nand2_1 _40803_ (.Y(_10215_),
    .A(_10006_),
    .B(_10214_));
 sg13g2_a21o_1 _40804_ (.A2(_10001_),
    .A1(_09996_),
    .B1(net5587),
    .X(_10216_));
 sg13g2_o21ai_1 _40805_ (.B1(net5650),
    .Y(_10217_),
    .A1(_09983_),
    .A2(_09990_));
 sg13g2_o21ai_1 _40806_ (.B1(_10217_),
    .Y(_10218_),
    .A1(_09992_),
    .A2(_10216_));
 sg13g2_inv_1 _40807_ (.Y(_10219_),
    .A(_10218_));
 sg13g2_a21o_1 _40808_ (.A2(_09968_),
    .A1(net5642),
    .B1(_09974_),
    .X(_10220_));
 sg13g2_a21oi_1 _40809_ (.A1(_09956_),
    .A2(_09962_),
    .Y(_10221_),
    .B1(net5582));
 sg13g2_a221oi_1 _40810_ (.B2(_09965_),
    .C1(_10221_),
    .B1(_10220_),
    .A1(_09978_),
    .Y(_10222_),
    .A2(_10218_));
 sg13g2_and3_2 _40811_ (.X(_10223_),
    .A(_10205_),
    .B(_10215_),
    .C(_10222_));
 sg13g2_a21o_2 _40812_ (.A2(_10223_),
    .A1(net1094),
    .B1(_08857_),
    .X(_10224_));
 sg13g2_a21o_2 _40813_ (.A2(net1078),
    .A1(_06950_),
    .B1(_08565_),
    .X(_10225_));
 sg13g2_nand2_1 _40814_ (.Y(_10226_),
    .A(_06120_),
    .B(_10225_));
 sg13g2_a21oi_1 _40815_ (.A1(_06120_),
    .A2(_10225_),
    .Y(_10227_),
    .B1(_06164_));
 sg13g2_a21o_1 _40816_ (.A2(_10225_),
    .A1(_06120_),
    .B1(_06164_),
    .X(_10228_));
 sg13g2_nand2_1 _40817_ (.Y(_10229_),
    .A(_06160_),
    .B(_10228_));
 sg13g2_o21ai_1 _40818_ (.B1(_06163_),
    .Y(_10230_),
    .A1(_06161_),
    .A2(_10227_));
 sg13g2_and2_1 _40819_ (.A(_06130_),
    .B(_10230_),
    .X(_10231_));
 sg13g2_a21oi_1 _40820_ (.A1(_06130_),
    .A2(_10230_),
    .Y(_10232_),
    .B1(_05454_));
 sg13g2_o21ai_1 _40821_ (.B1(_05426_),
    .Y(_10233_),
    .A1(_06132_),
    .A2(_10232_));
 sg13g2_a21oi_1 _40822_ (.A1(_05424_),
    .A2(_10233_),
    .Y(_10234_),
    .B1(_05435_));
 sg13g2_and3_1 _40823_ (.X(_10235_),
    .A(_05424_),
    .B(_05435_),
    .C(_10233_));
 sg13g2_or2_1 _40824_ (.X(_10236_),
    .B(_05434_),
    .A(net6788));
 sg13g2_o21ai_1 _40825_ (.B1(net6788),
    .Y(_10237_),
    .A1(_10234_),
    .A2(_10235_));
 sg13g2_nand2_2 _40826_ (.Y(_10238_),
    .A(_10236_),
    .B(_10237_));
 sg13g2_and3_2 _40827_ (.X(_10239_),
    .A(net5610),
    .B(_10236_),
    .C(_10237_));
 sg13g2_a21oi_1 _40828_ (.A1(_10236_),
    .A2(_10237_),
    .Y(_10240_),
    .B1(net5609));
 sg13g2_nor2_1 _40829_ (.A(_10239_),
    .B(_10240_),
    .Y(_10241_));
 sg13g2_or2_1 _40830_ (.X(_10242_),
    .B(_10240_),
    .A(_10239_));
 sg13g2_a21oi_2 _40831_ (.B1(_05456_),
    .Y(_10243_),
    .A2(_10230_),
    .A1(_06130_));
 sg13g2_or3_1 _40832_ (.A(_05412_),
    .B(_06135_),
    .C(_10243_),
    .X(_10244_));
 sg13g2_o21ai_1 _40833_ (.B1(_05412_),
    .Y(_10245_),
    .A1(_06135_),
    .A2(_10243_));
 sg13g2_nand3_1 _40834_ (.B(_10244_),
    .C(_10245_),
    .A(net6788),
    .Y(_10246_));
 sg13g2_o21ai_1 _40835_ (.B1(_10246_),
    .Y(_10247_),
    .A1(net6788),
    .A2(_05409_));
 sg13g2_nand2_1 _40836_ (.Y(_10248_),
    .A(net5609),
    .B(_10247_));
 sg13g2_xnor2_1 _40837_ (.Y(_10249_),
    .A(net5609),
    .B(_10247_));
 sg13g2_nand2_1 _40838_ (.Y(_10250_),
    .A(net6746),
    .B(_05423_));
 sg13g2_nor3_1 _40839_ (.A(_05426_),
    .B(_06132_),
    .C(_10232_),
    .Y(_10251_));
 sg13g2_nand2_1 _40840_ (.Y(_10252_),
    .A(net6788),
    .B(_10233_));
 sg13g2_o21ai_1 _40841_ (.B1(_10250_),
    .Y(_10253_),
    .A1(_10251_),
    .A2(_10252_));
 sg13g2_nand2_1 _40842_ (.Y(_10254_),
    .A(net5609),
    .B(_10253_));
 sg13g2_xnor2_1 _40843_ (.Y(_10255_),
    .A(net5609),
    .B(_10253_));
 sg13g2_nor2_1 _40844_ (.A(net6788),
    .B(_05444_),
    .Y(_10256_));
 sg13g2_o21ai_1 _40845_ (.B1(_05451_),
    .Y(_10257_),
    .A1(_05453_),
    .A2(_10231_));
 sg13g2_xor2_1 _40846_ (.B(_10257_),
    .A(_05446_),
    .X(_10258_));
 sg13g2_a21oi_2 _40847_ (.B1(_10256_),
    .Y(_10259_),
    .A2(_10258_),
    .A1(net6789));
 sg13g2_nand2_1 _40848_ (.Y(_10260_),
    .A(net5609),
    .B(_10259_));
 sg13g2_xnor2_1 _40849_ (.Y(_10261_),
    .A(net5609),
    .B(_10259_));
 sg13g2_nor4_1 _40850_ (.A(_10242_),
    .B(_10249_),
    .C(_10255_),
    .D(_10261_),
    .Y(_10262_));
 sg13g2_nor2_1 _40851_ (.A(net6790),
    .B(_08572_),
    .Y(_10263_));
 sg13g2_and3_1 _40852_ (.X(_10264_),
    .A(_06165_),
    .B(_08567_),
    .C(_08574_));
 sg13g2_o21ai_1 _40853_ (.B1(net6790),
    .Y(_10265_),
    .A1(_08575_),
    .A2(_10264_));
 sg13g2_nor2b_2 _40854_ (.A(_10263_),
    .B_N(_10265_),
    .Y(_10266_));
 sg13g2_xnor2_1 _40855_ (.Y(_10267_),
    .A(net5608),
    .B(_10266_));
 sg13g2_o21ai_1 _40856_ (.B1(net6746),
    .Y(_10268_),
    .A1(_05385_),
    .A2(_05389_));
 sg13g2_o21ai_1 _40857_ (.B1(_05413_),
    .Y(_10269_),
    .A1(_06135_),
    .A2(_10243_));
 sg13g2_a21o_1 _40858_ (.A2(_10269_),
    .A1(_06137_),
    .B1(_05380_),
    .X(_10270_));
 sg13g2_nand3_1 _40859_ (.B(_05394_),
    .C(_10270_),
    .A(_05379_),
    .Y(_10271_));
 sg13g2_a21o_1 _40860_ (.A2(_10270_),
    .A1(_05379_),
    .B1(_05394_),
    .X(_10272_));
 sg13g2_nand3_1 _40861_ (.B(_10271_),
    .C(_10272_),
    .A(net6788),
    .Y(_10273_));
 sg13g2_nand2_1 _40862_ (.Y(_10274_),
    .A(_10268_),
    .B(_10273_));
 sg13g2_and3_2 _40863_ (.X(_10275_),
    .A(net5608),
    .B(_10268_),
    .C(_10273_));
 sg13g2_a21oi_1 _40864_ (.A1(_10268_),
    .A2(_10273_),
    .Y(_10276_),
    .B1(net5608));
 sg13g2_or2_1 _40865_ (.X(_10277_),
    .B(_10276_),
    .A(_10275_));
 sg13g2_nor2_1 _40866_ (.A(_10267_),
    .B(_10277_),
    .Y(_10278_));
 sg13g2_o21ai_1 _40867_ (.B1(net6746),
    .Y(_10279_),
    .A1(_05398_),
    .A2(_05402_));
 sg13g2_nand4_1 _40868_ (.B(_05404_),
    .C(_05411_),
    .A(_05403_),
    .Y(_10280_),
    .D(_10245_));
 sg13g2_a22oi_1 _40869_ (.Y(_10281_),
    .B1(_05411_),
    .B2(_10245_),
    .A2(_05404_),
    .A1(_05403_));
 sg13g2_nand3b_1 _40870_ (.B(net6788),
    .C(_10280_),
    .Y(_10282_),
    .A_N(_10281_));
 sg13g2_nand2_1 _40871_ (.Y(_10283_),
    .A(_10279_),
    .B(_10282_));
 sg13g2_inv_2 _40872_ (.Y(_10284_),
    .A(_10283_));
 sg13g2_nand3_1 _40873_ (.B(_10279_),
    .C(_10282_),
    .A(net5608),
    .Y(_10285_));
 sg13g2_a21o_1 _40874_ (.A2(_10282_),
    .A1(_10279_),
    .B1(net5608),
    .X(_10286_));
 sg13g2_nand2_1 _40875_ (.Y(_10287_),
    .A(_10285_),
    .B(_10286_));
 sg13g2_nand3_1 _40876_ (.B(_06137_),
    .C(_10269_),
    .A(_05380_),
    .Y(_10288_));
 sg13g2_nand2_1 _40877_ (.Y(_10289_),
    .A(net6746),
    .B(_05378_));
 sg13g2_inv_1 _40878_ (.Y(_10290_),
    .A(_10289_));
 sg13g2_a21oi_1 _40879_ (.A1(_10270_),
    .A2(_10288_),
    .Y(_10291_),
    .B1(net6746));
 sg13g2_or2_1 _40880_ (.X(_10292_),
    .B(_10291_),
    .A(_10290_));
 sg13g2_o21ai_1 _40881_ (.B1(net5576),
    .Y(_10293_),
    .A1(_10290_),
    .A2(_10291_));
 sg13g2_nand3b_1 _40882_ (.B(net5608),
    .C(_10289_),
    .Y(_10294_),
    .A_N(_10291_));
 sg13g2_and2_1 _40883_ (.A(_10293_),
    .B(_10294_),
    .X(_10295_));
 sg13g2_nand4_1 _40884_ (.B(_10286_),
    .C(_10293_),
    .A(_10285_),
    .Y(_10296_),
    .D(_10294_));
 sg13g2_nor4_1 _40885_ (.A(_10267_),
    .B(_10275_),
    .C(_10276_),
    .D(_10296_),
    .Y(_10297_));
 sg13g2_nand2_2 _40886_ (.Y(_10298_),
    .A(_10262_),
    .B(_10297_));
 sg13g2_nand2_1 _40887_ (.Y(_10299_),
    .A(net6750),
    .B(_05522_));
 sg13g2_o21ai_1 _40888_ (.B1(_05540_),
    .Y(_10300_),
    .A1(_06161_),
    .A2(_10227_));
 sg13g2_a21oi_1 _40889_ (.A1(_06160_),
    .A2(_10228_),
    .Y(_10301_),
    .B1(_05542_));
 sg13g2_o21ai_1 _40890_ (.B1(_05513_),
    .Y(_10302_),
    .A1(_06122_),
    .A2(_10301_));
 sg13g2_and3_1 _40891_ (.X(_10303_),
    .A(_05512_),
    .B(_05523_),
    .C(_10302_));
 sg13g2_a21oi_1 _40892_ (.A1(_05512_),
    .A2(_10302_),
    .Y(_10304_),
    .B1(_05523_));
 sg13g2_o21ai_1 _40893_ (.B1(net6793),
    .Y(_10305_),
    .A1(_10303_),
    .A2(_10304_));
 sg13g2_nand2_1 _40894_ (.Y(_10306_),
    .A(_10299_),
    .B(_10305_));
 sg13g2_inv_1 _40895_ (.Y(_10307_),
    .A(_10306_));
 sg13g2_and3_2 _40896_ (.X(_10308_),
    .A(net5612),
    .B(_10299_),
    .C(_10305_));
 sg13g2_a21oi_1 _40897_ (.A1(_10299_),
    .A2(_10305_),
    .Y(_10309_),
    .B1(net5612));
 sg13g2_nand2_1 _40898_ (.Y(_10310_),
    .A(net5576),
    .B(_10306_));
 sg13g2_or2_1 _40899_ (.X(_10311_),
    .B(_10309_),
    .A(_10308_));
 sg13g2_nand2_1 _40900_ (.Y(_10312_),
    .A(net6746),
    .B(_05490_));
 sg13g2_a21oi_2 _40901_ (.B1(_06124_),
    .Y(_10313_),
    .A2(_10301_),
    .A1(_05524_));
 sg13g2_xnor2_1 _40902_ (.Y(_10314_),
    .A(_05492_),
    .B(_10313_));
 sg13g2_o21ai_1 _40903_ (.B1(_10312_),
    .Y(_10315_),
    .A1(net6758),
    .A2(_10314_));
 sg13g2_xnor2_1 _40904_ (.Y(_10316_),
    .A(net5612),
    .B(_10315_));
 sg13g2_or3_1 _40905_ (.A(_05513_),
    .B(_06122_),
    .C(_10301_),
    .X(_10317_));
 sg13g2_nand3_1 _40906_ (.B(_10302_),
    .C(_10317_),
    .A(net6793),
    .Y(_10318_));
 sg13g2_o21ai_1 _40907_ (.B1(_10318_),
    .Y(_10319_),
    .A1(net6793),
    .A2(_05511_));
 sg13g2_nor2_1 _40908_ (.A(net5612),
    .B(_10319_),
    .Y(_10320_));
 sg13g2_xnor2_1 _40909_ (.Y(_10321_),
    .A(net5576),
    .B(_10319_));
 sg13g2_nor2_1 _40910_ (.A(net6793),
    .B(_05531_),
    .Y(_10322_));
 sg13g2_nand2_1 _40911_ (.Y(_10323_),
    .A(_05539_),
    .B(_10300_));
 sg13g2_xor2_1 _40912_ (.B(_10323_),
    .A(_05533_),
    .X(_10324_));
 sg13g2_a21oi_2 _40913_ (.B1(_10322_),
    .Y(_10325_),
    .A2(_10324_),
    .A1(net6793));
 sg13g2_nand2_1 _40914_ (.Y(_10326_),
    .A(net5617),
    .B(_10325_));
 sg13g2_xnor2_1 _40915_ (.Y(_10327_),
    .A(net5573),
    .B(_10325_));
 sg13g2_nand2_1 _40916_ (.Y(_10328_),
    .A(_10321_),
    .B(_10327_));
 sg13g2_nor3_1 _40917_ (.A(_10311_),
    .B(_10316_),
    .C(_10328_),
    .Y(_10329_));
 sg13g2_nand2_1 _40918_ (.Y(_10330_),
    .A(net6746),
    .B(_05450_));
 sg13g2_xnor2_1 _40919_ (.Y(_10331_),
    .A(_05453_),
    .B(_10231_));
 sg13g2_o21ai_1 _40920_ (.B1(_10330_),
    .Y(_10332_),
    .A1(net6746),
    .A2(_10331_));
 sg13g2_nand2_1 _40921_ (.Y(_10333_),
    .A(net5611),
    .B(_10332_));
 sg13g2_xnor2_1 _40922_ (.Y(_10334_),
    .A(net5611),
    .B(_10332_));
 sg13g2_nor2_1 _40923_ (.A(net6789),
    .B(_05483_),
    .Y(_10335_));
 sg13g2_o21ai_1 _40924_ (.B1(_06126_),
    .Y(_10336_),
    .A1(_05502_),
    .A2(_10313_));
 sg13g2_a21oi_1 _40925_ (.A1(_05474_),
    .A2(_10336_),
    .Y(_10337_),
    .B1(_05473_));
 sg13g2_xnor2_1 _40926_ (.Y(_10338_),
    .A(_05484_),
    .B(_10337_));
 sg13g2_a21oi_2 _40927_ (.B1(_10335_),
    .Y(_10339_),
    .A2(_10338_),
    .A1(net6789));
 sg13g2_nand2_1 _40928_ (.Y(_10340_),
    .A(net5611),
    .B(_10339_));
 sg13g2_xnor2_1 _40929_ (.Y(_10341_),
    .A(net5611),
    .B(_10339_));
 sg13g2_nor2_1 _40930_ (.A(net6789),
    .B(_05500_),
    .Y(_10342_));
 sg13g2_o21ai_1 _40931_ (.B1(_05491_),
    .Y(_10343_),
    .A1(_05492_),
    .A2(_10313_));
 sg13g2_xor2_1 _40932_ (.B(_10343_),
    .A(_05501_),
    .X(_10344_));
 sg13g2_a21oi_2 _40933_ (.B1(_10342_),
    .Y(_10345_),
    .A2(_10344_),
    .A1(net6789));
 sg13g2_nand2_1 _40934_ (.Y(_10346_),
    .A(net5611),
    .B(_10345_));
 sg13g2_xnor2_1 _40935_ (.Y(_10347_),
    .A(net5576),
    .B(_10345_));
 sg13g2_inv_2 _40936_ (.Y(_10348_),
    .A(_10347_));
 sg13g2_nor2_1 _40937_ (.A(net6789),
    .B(_05471_),
    .Y(_10349_));
 sg13g2_xnor2_1 _40938_ (.Y(_10350_),
    .A(_05474_),
    .B(_10336_));
 sg13g2_a21oi_2 _40939_ (.B1(_10349_),
    .Y(_10351_),
    .A2(_10350_),
    .A1(net6789));
 sg13g2_xnor2_1 _40940_ (.Y(_10352_),
    .A(net5611),
    .B(_10351_));
 sg13g2_nor4_1 _40941_ (.A(_10334_),
    .B(_10341_),
    .C(_10348_),
    .D(_10352_),
    .Y(_10353_));
 sg13g2_nand2_1 _40942_ (.Y(_10354_),
    .A(_10329_),
    .B(_10353_));
 sg13g2_nor2_2 _40943_ (.A(_10298_),
    .B(_10354_),
    .Y(_10355_));
 sg13g2_nand2_1 _40944_ (.Y(_10356_),
    .A(net6750),
    .B(_05568_));
 sg13g2_and2_1 _40945_ (.A(_05720_),
    .B(_10226_),
    .X(_10357_));
 sg13g2_o21ai_1 _40946_ (.B1(_05600_),
    .Y(_10358_),
    .A1(_06157_),
    .A2(_10357_));
 sg13g2_o21ai_1 _40947_ (.B1(_05611_),
    .Y(_10359_),
    .A1(_06157_),
    .A2(_10357_));
 sg13g2_o21ai_1 _40948_ (.B1(_06143_),
    .Y(_10360_),
    .A1(_05629_),
    .A2(_10359_));
 sg13g2_a21oi_1 _40949_ (.A1(_05591_),
    .A2(_10360_),
    .Y(_10361_),
    .B1(_06146_));
 sg13g2_o21ai_1 _40950_ (.B1(_05559_),
    .Y(_10362_),
    .A1(_05560_),
    .A2(_10361_));
 sg13g2_xor2_1 _40951_ (.B(_10362_),
    .A(_05569_),
    .X(_10363_));
 sg13g2_o21ai_1 _40952_ (.B1(_10356_),
    .Y(_10364_),
    .A1(net6750),
    .A2(_10363_));
 sg13g2_and2_1 _40953_ (.A(net5617),
    .B(_10364_),
    .X(_10365_));
 sg13g2_xnor2_1 _40954_ (.Y(_10366_),
    .A(net5573),
    .B(_10364_));
 sg13g2_nand2_1 _40955_ (.Y(_10367_),
    .A(net6750),
    .B(_05538_));
 sg13g2_xnor2_1 _40956_ (.Y(_10368_),
    .A(_05540_),
    .B(_10229_));
 sg13g2_o21ai_1 _40957_ (.B1(_10367_),
    .Y(_10369_),
    .A1(net6750),
    .A2(_10368_));
 sg13g2_xnor2_1 _40958_ (.Y(_10370_),
    .A(net5573),
    .B(_10369_));
 sg13g2_nand2_1 _40959_ (.Y(_10371_),
    .A(net6749),
    .B(_05588_));
 sg13g2_a21oi_1 _40960_ (.A1(_05580_),
    .A2(_10360_),
    .Y(_10372_),
    .B1(_05578_));
 sg13g2_xnor2_1 _40961_ (.Y(_10373_),
    .A(_05589_),
    .B(_10372_));
 sg13g2_o21ai_1 _40962_ (.B1(_10371_),
    .Y(_10374_),
    .A1(net6750),
    .A2(_10373_));
 sg13g2_nand2_1 _40963_ (.Y(_10375_),
    .A(net5617),
    .B(_10374_));
 sg13g2_xnor2_1 _40964_ (.Y(_10376_),
    .A(net5617),
    .B(_10374_));
 sg13g2_inv_1 _40965_ (.Y(_10377_),
    .A(_10376_));
 sg13g2_nand2_1 _40966_ (.Y(_10378_),
    .A(net6750),
    .B(_05558_));
 sg13g2_xnor2_1 _40967_ (.Y(_10379_),
    .A(_05560_),
    .B(_10361_));
 sg13g2_o21ai_1 _40968_ (.B1(_10378_),
    .Y(_10380_),
    .A1(net6750),
    .A2(_10379_));
 sg13g2_nor2_1 _40969_ (.A(net5617),
    .B(_10380_),
    .Y(_10381_));
 sg13g2_xnor2_1 _40970_ (.Y(_10382_),
    .A(net5573),
    .B(_10380_));
 sg13g2_nand4_1 _40971_ (.B(_10370_),
    .C(_10377_),
    .A(_10366_),
    .Y(_10383_),
    .D(_10382_));
 sg13g2_nand2_1 _40972_ (.Y(_10384_),
    .A(net6749),
    .B(_05627_));
 sg13g2_a21o_1 _40973_ (.A2(_10359_),
    .A1(_06140_),
    .B1(_05619_),
    .X(_10385_));
 sg13g2_a21oi_1 _40974_ (.A1(_05618_),
    .A2(_10385_),
    .Y(_10386_),
    .B1(_05628_));
 sg13g2_nand3_1 _40975_ (.B(_05628_),
    .C(_10385_),
    .A(_05618_),
    .Y(_10387_));
 sg13g2_nand2_1 _40976_ (.Y(_10388_),
    .A(net6791),
    .B(_10387_));
 sg13g2_o21ai_1 _40977_ (.B1(_10384_),
    .Y(_10389_),
    .A1(_10386_),
    .A2(_10388_));
 sg13g2_and2_1 _40978_ (.A(net5615),
    .B(_10389_),
    .X(_10390_));
 sg13g2_xnor2_1 _40979_ (.Y(_10391_),
    .A(net5571),
    .B(_10389_));
 sg13g2_nor2_1 _40980_ (.A(net6791),
    .B(_05576_),
    .Y(_10392_));
 sg13g2_xnor2_1 _40981_ (.Y(_10393_),
    .A(_05580_),
    .B(_10360_));
 sg13g2_a21oi_2 _40982_ (.B1(_10392_),
    .Y(_10394_),
    .A2(_10393_),
    .A1(net6791));
 sg13g2_xnor2_1 _40983_ (.Y(_10395_),
    .A(net5571),
    .B(_10394_));
 sg13g2_nand2_1 _40984_ (.Y(_10396_),
    .A(_10391_),
    .B(_10395_));
 sg13g2_nand3_1 _40985_ (.B(_06140_),
    .C(_10359_),
    .A(_05619_),
    .Y(_10397_));
 sg13g2_and3_1 _40986_ (.X(_10398_),
    .A(net6791),
    .B(_10385_),
    .C(_10397_));
 sg13g2_a21oi_2 _40987_ (.B1(_10398_),
    .Y(_10399_),
    .A2(_05617_),
    .A1(net6749));
 sg13g2_inv_1 _40988_ (.Y(_10400_),
    .A(_10399_));
 sg13g2_xnor2_1 _40989_ (.Y(_10401_),
    .A(net5615),
    .B(_10399_));
 sg13g2_nor2_1 _40990_ (.A(net6791),
    .B(_05608_),
    .Y(_10402_));
 sg13g2_nand2_1 _40991_ (.Y(_10403_),
    .A(_05599_),
    .B(_10358_));
 sg13g2_xnor2_1 _40992_ (.Y(_10404_),
    .A(_05610_),
    .B(_10403_));
 sg13g2_a21oi_2 _40993_ (.B1(_10402_),
    .Y(_10405_),
    .A2(_10404_),
    .A1(net6791));
 sg13g2_nand2_1 _40994_ (.Y(_10406_),
    .A(net5615),
    .B(_10405_));
 sg13g2_xnor2_1 _40995_ (.Y(_10407_),
    .A(net5571),
    .B(_10405_));
 sg13g2_nand4_1 _40996_ (.B(_10395_),
    .C(_10401_),
    .A(_10391_),
    .Y(_10408_),
    .D(_10407_));
 sg13g2_nand2_1 _40997_ (.Y(_10409_),
    .A(_05717_),
    .B(_10226_));
 sg13g2_a21oi_1 _40998_ (.A1(_06120_),
    .A2(_10225_),
    .Y(_10410_),
    .B1(_05719_));
 sg13g2_a21oi_1 _40999_ (.A1(_05701_),
    .A2(_10410_),
    .Y(_10411_),
    .B1(_06151_));
 sg13g2_o21ai_1 _41000_ (.B1(_05667_),
    .Y(_10412_),
    .A1(_05669_),
    .A2(_10411_));
 sg13g2_nand3b_1 _41001_ (.B(_05680_),
    .C(_05668_),
    .Y(_10413_),
    .A_N(_10411_));
 sg13g2_a21oi_1 _41002_ (.A1(_06154_),
    .A2(_10413_),
    .Y(_10414_),
    .B1(_05657_));
 sg13g2_or3_1 _41003_ (.A(_05650_),
    .B(_05656_),
    .C(_10414_),
    .X(_10415_));
 sg13g2_o21ai_1 _41004_ (.B1(_05650_),
    .Y(_10416_),
    .A1(_05656_),
    .A2(_10414_));
 sg13g2_nand3_1 _41005_ (.B(_05640_),
    .C(_05647_),
    .A(net6748),
    .Y(_10417_));
 sg13g2_a21o_1 _41006_ (.A2(_10416_),
    .A1(_10415_),
    .B1(net6747),
    .X(_10418_));
 sg13g2_nand2_2 _41007_ (.Y(_10419_),
    .A(_10417_),
    .B(_10418_));
 sg13g2_a21oi_1 _41008_ (.A1(_10417_),
    .A2(_10418_),
    .Y(_10420_),
    .B1(net5571));
 sg13g2_xnor2_1 _41009_ (.Y(_10421_),
    .A(net5614),
    .B(_10419_));
 sg13g2_or3_1 _41010_ (.A(_05600_),
    .B(_06157_),
    .C(_10357_),
    .X(_10422_));
 sg13g2_nand3_1 _41011_ (.B(_10358_),
    .C(_10422_),
    .A(net6791),
    .Y(_10423_));
 sg13g2_o21ai_1 _41012_ (.B1(_10423_),
    .Y(_10424_),
    .A1(net6792),
    .A2(_05598_));
 sg13g2_xnor2_1 _41013_ (.Y(_10425_),
    .A(net5614),
    .B(_10424_));
 sg13g2_nor2_1 _41014_ (.A(_10421_),
    .B(_10425_),
    .Y(_10426_));
 sg13g2_nand3_1 _41015_ (.B(_05674_),
    .C(_05677_),
    .A(net6748),
    .Y(_10427_));
 sg13g2_xnor2_1 _41016_ (.Y(_10428_),
    .A(_05680_),
    .B(_10412_));
 sg13g2_o21ai_1 _41017_ (.B1(_10427_),
    .Y(_10429_),
    .A1(net6747),
    .A2(_10428_));
 sg13g2_and2_1 _41018_ (.A(net5614),
    .B(_10429_),
    .X(_10430_));
 sg13g2_xnor2_1 _41019_ (.Y(_10431_),
    .A(net5572),
    .B(_10429_));
 sg13g2_inv_1 _41020_ (.Y(_10432_),
    .A(_10431_));
 sg13g2_and3_1 _41021_ (.X(_10433_),
    .A(_05657_),
    .B(_06154_),
    .C(_10413_));
 sg13g2_o21ai_1 _41022_ (.B1(net6791),
    .Y(_10434_),
    .A1(_10414_),
    .A2(_10433_));
 sg13g2_or2_1 _41023_ (.X(_10435_),
    .B(_05655_),
    .A(net6792));
 sg13g2_and2_1 _41024_ (.A(_10434_),
    .B(_10435_),
    .X(_10436_));
 sg13g2_nand3_1 _41025_ (.B(_10434_),
    .C(_10435_),
    .A(net5614),
    .Y(_10437_));
 sg13g2_a21o_1 _41026_ (.A2(_10435_),
    .A1(_10434_),
    .B1(net5614),
    .X(_10438_));
 sg13g2_and2_1 _41027_ (.A(_10437_),
    .B(_10438_),
    .X(_10439_));
 sg13g2_nand2_1 _41028_ (.Y(_10440_),
    .A(_10431_),
    .B(_10439_));
 sg13g2_nor3_1 _41029_ (.A(_10421_),
    .B(_10425_),
    .C(_10440_),
    .Y(_10441_));
 sg13g2_nand2_1 _41030_ (.Y(_10442_),
    .A(net6747),
    .B(_05666_));
 sg13g2_xnor2_1 _41031_ (.Y(_10443_),
    .A(_05669_),
    .B(_10411_));
 sg13g2_o21ai_1 _41032_ (.B1(_10442_),
    .Y(_10444_),
    .A1(net6747),
    .A2(_10443_));
 sg13g2_xnor2_1 _41033_ (.Y(_10445_),
    .A(net5572),
    .B(_10444_));
 sg13g2_nor2_1 _41034_ (.A(net6792),
    .B(_05699_),
    .Y(_10446_));
 sg13g2_nor2_1 _41035_ (.A(_06148_),
    .B(_10410_),
    .Y(_10447_));
 sg13g2_o21ai_1 _41036_ (.B1(_05689_),
    .Y(_10448_),
    .A1(_05691_),
    .A2(_10447_));
 sg13g2_xnor2_1 _41037_ (.Y(_10449_),
    .A(_05700_),
    .B(_10448_));
 sg13g2_a21oi_2 _41038_ (.B1(_10446_),
    .Y(_10450_),
    .A2(_10449_),
    .A1(net6792));
 sg13g2_and2_1 _41039_ (.A(net5614),
    .B(_10450_),
    .X(_10451_));
 sg13g2_xnor2_1 _41040_ (.Y(_10452_),
    .A(net5572),
    .B(_10450_));
 sg13g2_and2_1 _41041_ (.A(_10445_),
    .B(_10452_),
    .X(_10453_));
 sg13g2_nand2_1 _41042_ (.Y(_10454_),
    .A(_10445_),
    .B(_10452_));
 sg13g2_nand2_1 _41043_ (.Y(_10455_),
    .A(net6748),
    .B(_05688_));
 sg13g2_xnor2_1 _41044_ (.Y(_10456_),
    .A(_05691_),
    .B(_10447_));
 sg13g2_o21ai_1 _41045_ (.B1(_10455_),
    .Y(_10457_),
    .A1(net6748),
    .A2(_10456_));
 sg13g2_inv_1 _41046_ (.Y(_10458_),
    .A(_10457_));
 sg13g2_xnor2_1 _41047_ (.Y(_10459_),
    .A(net5571),
    .B(_10457_));
 sg13g2_nand2_1 _41048_ (.Y(_10460_),
    .A(net6747),
    .B(_05708_));
 sg13g2_nand2_1 _41049_ (.Y(_10461_),
    .A(_05716_),
    .B(_10409_));
 sg13g2_xor2_1 _41050_ (.B(_10461_),
    .A(_05710_),
    .X(_10462_));
 sg13g2_o21ai_1 _41051_ (.B1(_10460_),
    .Y(_10463_),
    .A1(net6747),
    .A2(_10462_));
 sg13g2_and2_1 _41052_ (.A(net5615),
    .B(_10463_),
    .X(_10464_));
 sg13g2_xnor2_1 _41053_ (.Y(_10465_),
    .A(net5571),
    .B(_10463_));
 sg13g2_nand3_1 _41054_ (.B(_10459_),
    .C(_10465_),
    .A(_10453_),
    .Y(_10466_));
 sg13g2_nor4_1 _41055_ (.A(_10421_),
    .B(_10425_),
    .C(_10440_),
    .D(_10466_),
    .Y(_10467_));
 sg13g2_nand4_1 _41056_ (.B(_10453_),
    .C(_10459_),
    .A(_10441_),
    .Y(_10468_),
    .D(_10465_));
 sg13g2_nor3_2 _41057_ (.A(_10383_),
    .B(_10408_),
    .C(_10468_),
    .Y(_10469_));
 sg13g2_and2_1 _41058_ (.A(_10355_),
    .B(_10469_),
    .X(_10470_));
 sg13g2_a21oi_1 _41059_ (.A1(_06950_),
    .A2(net1077),
    .Y(_10471_),
    .B1(_08561_));
 sg13g2_o21ai_1 _41060_ (.B1(_06049_),
    .Y(_10472_),
    .A1(_06090_),
    .A2(_10471_));
 sg13g2_nand2_1 _41061_ (.Y(_10473_),
    .A(_06048_),
    .B(_10472_));
 sg13g2_a22oi_1 _41062_ (.Y(_10474_),
    .B1(_06092_),
    .B2(_10472_),
    .A2(_06041_),
    .A1(net5841));
 sg13g2_a221oi_1 _41063_ (.B2(_10472_),
    .C1(_06019_),
    .B1(_06092_),
    .A1(net5842),
    .Y(_10475_),
    .A2(_06041_));
 sg13g2_o21ai_1 _41064_ (.B1(_06030_),
    .Y(_10476_),
    .A1(_06018_),
    .A2(_10475_));
 sg13g2_or3_1 _41065_ (.A(_06018_),
    .B(_06030_),
    .C(_10475_),
    .X(_10477_));
 sg13g2_a21oi_1 _41066_ (.A1(_10476_),
    .A2(_10477_),
    .Y(_10478_),
    .B1(net6753));
 sg13g2_a21oi_2 _41067_ (.B1(_10478_),
    .Y(_10479_),
    .A2(_06028_),
    .A1(net6753));
 sg13g2_and2_1 _41068_ (.A(net5623),
    .B(_10479_),
    .X(_10480_));
 sg13g2_inv_1 _41069_ (.Y(_10481_),
    .A(_10480_));
 sg13g2_xnor2_1 _41070_ (.Y(_10482_),
    .A(net5623),
    .B(_10479_));
 sg13g2_nand2_1 _41071_ (.Y(_10483_),
    .A(net6753),
    .B(_05993_));
 sg13g2_a21oi_1 _41072_ (.A1(_06950_),
    .A2(net1078),
    .Y(_10484_),
    .B1(_08563_));
 sg13g2_nor2_1 _41073_ (.A(_06094_),
    .B(_10484_),
    .Y(_10485_));
 sg13g2_o21ai_1 _41074_ (.B1(_05995_),
    .Y(_10486_),
    .A1(_06094_),
    .A2(_10484_));
 sg13g2_xnor2_1 _41075_ (.Y(_10487_),
    .A(_05995_),
    .B(_10485_));
 sg13g2_o21ai_1 _41076_ (.B1(_10483_),
    .Y(_10488_),
    .A1(net6753),
    .A2(_10487_));
 sg13g2_inv_1 _41077_ (.Y(_10489_),
    .A(_10488_));
 sg13g2_nor2_1 _41078_ (.A(net5577),
    .B(_10488_),
    .Y(_10490_));
 sg13g2_xnor2_1 _41079_ (.Y(_10491_),
    .A(net5577),
    .B(_10488_));
 sg13g2_nand2_1 _41080_ (.Y(_10492_),
    .A(net6753),
    .B(_06017_));
 sg13g2_xnor2_1 _41081_ (.Y(_10493_),
    .A(_06020_),
    .B(_10474_));
 sg13g2_o21ai_1 _41082_ (.B1(_10492_),
    .Y(_10494_),
    .A1(net6753),
    .A2(_10493_));
 sg13g2_nand2b_1 _41083_ (.Y(_10495_),
    .B(net5577),
    .A_N(_10494_));
 sg13g2_xnor2_1 _41084_ (.Y(_10496_),
    .A(net5626),
    .B(_10494_));
 sg13g2_nor2_1 _41085_ (.A(net6797),
    .B(_06040_),
    .Y(_10497_));
 sg13g2_xnor2_1 _41086_ (.Y(_10498_),
    .A(_06042_),
    .B(_10473_));
 sg13g2_a21oi_2 _41087_ (.B1(_10497_),
    .Y(_10499_),
    .A2(_10498_),
    .A1(net6796));
 sg13g2_xnor2_1 _41088_ (.Y(_10500_),
    .A(net5626),
    .B(_10499_));
 sg13g2_or2_1 _41089_ (.X(_10501_),
    .B(_10500_),
    .A(_10496_));
 sg13g2_nand2_1 _41090_ (.Y(_10502_),
    .A(net6755),
    .B(_06047_));
 sg13g2_nor3_1 _41091_ (.A(_06049_),
    .B(_06090_),
    .C(_10471_),
    .Y(_10503_));
 sg13g2_nand2_1 _41092_ (.Y(_10504_),
    .A(net6798),
    .B(_10472_));
 sg13g2_o21ai_1 _41093_ (.B1(_10502_),
    .Y(_10505_),
    .A1(_10503_),
    .A2(_10504_));
 sg13g2_xnor2_1 _41094_ (.Y(_10506_),
    .A(net5577),
    .B(_10505_));
 sg13g2_xnor2_1 _41095_ (.Y(_10507_),
    .A(net5626),
    .B(_10505_));
 sg13g2_nor2_1 _41096_ (.A(net6798),
    .B(_06070_),
    .Y(_10508_));
 sg13g2_inv_1 _41097_ (.Y(_10509_),
    .A(_10508_));
 sg13g2_nor2b_1 _41098_ (.A(_06079_),
    .B_N(_08605_),
    .Y(_10510_));
 sg13g2_a22oi_1 _41099_ (.Y(_10511_),
    .B1(_06088_),
    .B2(_08605_),
    .A2(_06087_),
    .A1(net5842));
 sg13g2_a221oi_1 _41100_ (.B2(_08605_),
    .C1(_06062_),
    .B1(_06088_),
    .A1(net5842),
    .Y(_10512_),
    .A2(_06087_));
 sg13g2_or3_1 _41101_ (.A(_06060_),
    .B(_06071_),
    .C(_10512_),
    .X(_10513_));
 sg13g2_o21ai_1 _41102_ (.B1(_06071_),
    .Y(_10514_),
    .A1(_06060_),
    .A2(_10512_));
 sg13g2_a21o_1 _41103_ (.A2(_10514_),
    .A1(_10513_),
    .B1(net6755),
    .X(_10515_));
 sg13g2_and2_1 _41104_ (.A(_10509_),
    .B(_10515_),
    .X(_10516_));
 sg13g2_and3_2 _41105_ (.X(_10517_),
    .A(net5626),
    .B(_10509_),
    .C(_10515_));
 sg13g2_a21oi_1 _41106_ (.A1(_10509_),
    .A2(_10515_),
    .Y(_10518_),
    .B1(net5626));
 sg13g2_or2_1 _41107_ (.X(_10519_),
    .B(_10518_),
    .A(_10517_));
 sg13g2_inv_1 _41108_ (.Y(_10520_),
    .A(_10519_));
 sg13g2_nor3_1 _41109_ (.A(_10507_),
    .B(_10517_),
    .C(_10518_),
    .Y(_10521_));
 sg13g2_a21oi_1 _41110_ (.A1(_06082_),
    .A2(_06086_),
    .Y(_10522_),
    .B1(net6798));
 sg13g2_xnor2_1 _41111_ (.Y(_10523_),
    .A(_08560_),
    .B(_10510_));
 sg13g2_a21oi_2 _41112_ (.B1(_10522_),
    .Y(_10524_),
    .A2(_10523_),
    .A1(net6798));
 sg13g2_nand2_1 _41113_ (.Y(_10525_),
    .A(net5627),
    .B(_10524_));
 sg13g2_xnor2_1 _41114_ (.Y(_10526_),
    .A(net5627),
    .B(_10524_));
 sg13g2_nand2b_1 _41115_ (.Y(_10527_),
    .B(net6755),
    .A_N(_06059_));
 sg13g2_xnor2_1 _41116_ (.Y(_10528_),
    .A(_06061_),
    .B(_10511_));
 sg13g2_o21ai_1 _41117_ (.B1(_10527_),
    .Y(_10529_),
    .A1(net6755),
    .A2(_10528_));
 sg13g2_inv_1 _41118_ (.Y(_10530_),
    .A(_10529_));
 sg13g2_xnor2_1 _41119_ (.Y(_10531_),
    .A(net5627),
    .B(_10529_));
 sg13g2_nor2_1 _41120_ (.A(_10526_),
    .B(_10531_),
    .Y(_10532_));
 sg13g2_nand2_1 _41121_ (.Y(_10533_),
    .A(_10521_),
    .B(_10532_));
 sg13g2_or4_1 _41122_ (.A(_10482_),
    .B(_10491_),
    .C(_10501_),
    .D(_10533_),
    .X(_10534_));
 sg13g2_nor2_1 _41123_ (.A(net6797),
    .B(_05986_),
    .Y(_10535_));
 sg13g2_o21ai_1 _41124_ (.B1(_06008_),
    .Y(_10536_),
    .A1(_06094_),
    .A2(_10484_));
 sg13g2_nand2_1 _41125_ (.Y(_10537_),
    .A(_06096_),
    .B(_10536_));
 sg13g2_a21oi_1 _41126_ (.A1(_05978_),
    .A2(_10537_),
    .Y(_10538_),
    .B1(_05977_));
 sg13g2_xor2_1 _41127_ (.B(_10538_),
    .A(_05987_),
    .X(_10539_));
 sg13g2_a21oi_2 _41128_ (.B1(_10535_),
    .Y(_10540_),
    .A2(_10539_),
    .A1(net6797));
 sg13g2_xnor2_1 _41129_ (.Y(_10541_),
    .A(net5624),
    .B(_10540_));
 sg13g2_nor2_1 _41130_ (.A(net6797),
    .B(_05965_),
    .Y(_10542_));
 sg13g2_o21ai_1 _41131_ (.B1(_06099_),
    .Y(_10543_),
    .A1(_05988_),
    .A2(_10536_));
 sg13g2_xor2_1 _41132_ (.B(_10543_),
    .A(_05967_),
    .X(_10544_));
 sg13g2_a21oi_1 _41133_ (.A1(net6797),
    .A2(_10544_),
    .Y(_10545_),
    .B1(_10542_));
 sg13g2_inv_1 _41134_ (.Y(_10546_),
    .A(_10545_));
 sg13g2_xnor2_1 _41135_ (.Y(_10547_),
    .A(net5624),
    .B(_10545_));
 sg13g2_inv_1 _41136_ (.Y(_10548_),
    .A(_10547_));
 sg13g2_nand2b_1 _41137_ (.Y(_10549_),
    .B(_10547_),
    .A_N(_10541_));
 sg13g2_nand2_1 _41138_ (.Y(_10550_),
    .A(net6754),
    .B(_05976_));
 sg13g2_xnor2_1 _41139_ (.Y(_10551_),
    .A(_05978_),
    .B(_10537_));
 sg13g2_o21ai_1 _41140_ (.B1(_10550_),
    .Y(_10552_),
    .A1(net6754),
    .A2(_10551_));
 sg13g2_inv_1 _41141_ (.Y(_10553_),
    .A(_10552_));
 sg13g2_xnor2_1 _41142_ (.Y(_10554_),
    .A(net5625),
    .B(_10552_));
 sg13g2_nor2_1 _41143_ (.A(net6797),
    .B(_06003_),
    .Y(_10555_));
 sg13g2_nand2_1 _41144_ (.Y(_10556_),
    .A(_05994_),
    .B(_10486_));
 sg13g2_xnor2_1 _41145_ (.Y(_10557_),
    .A(_06006_),
    .B(_10556_));
 sg13g2_a21oi_2 _41146_ (.B1(_10555_),
    .Y(_10558_),
    .A2(_10557_),
    .A1(net6797));
 sg13g2_nand2_1 _41147_ (.Y(_10559_),
    .A(net5625),
    .B(_10558_));
 sg13g2_xnor2_1 _41148_ (.Y(_10560_),
    .A(net5625),
    .B(_10558_));
 sg13g2_inv_1 _41149_ (.Y(_10561_),
    .A(_10560_));
 sg13g2_nor4_1 _41150_ (.A(_10541_),
    .B(_10548_),
    .C(_10554_),
    .D(_10560_),
    .Y(_10562_));
 sg13g2_inv_1 _41151_ (.Y(_10563_),
    .A(_10562_));
 sg13g2_nand2_1 _41152_ (.Y(_10564_),
    .A(net6756),
    .B(_05907_));
 sg13g2_a21oi_2 _41153_ (.B1(_08564_),
    .Y(_10565_),
    .A2(net1078),
    .A1(_06950_));
 sg13g2_nor2_1 _41154_ (.A(_06103_),
    .B(_10565_),
    .Y(_10566_));
 sg13g2_o21ai_1 _41155_ (.B1(_05909_),
    .Y(_10567_),
    .A1(_06103_),
    .A2(_10565_));
 sg13g2_xor2_1 _41156_ (.B(_10566_),
    .A(_05909_),
    .X(_10568_));
 sg13g2_o21ai_1 _41157_ (.B1(_10564_),
    .Y(_10569_),
    .A1(net6756),
    .A2(_10568_));
 sg13g2_xnor2_1 _41158_ (.Y(_10570_),
    .A(net5623),
    .B(_10569_));
 sg13g2_a21oi_1 _41159_ (.A1(_05939_),
    .A2(_05942_),
    .Y(_10571_),
    .B1(net6796));
 sg13g2_a21oi_1 _41160_ (.A1(_05968_),
    .A2(_10543_),
    .Y(_10572_),
    .B1(_06101_));
 sg13g2_o21ai_1 _41161_ (.B1(_05933_),
    .Y(_10573_),
    .A1(_05934_),
    .A2(_10572_));
 sg13g2_xnor2_1 _41162_ (.Y(_10574_),
    .A(_05946_),
    .B(_10573_));
 sg13g2_a21oi_2 _41163_ (.B1(_10571_),
    .Y(_10575_),
    .A2(_10574_),
    .A1(net6796));
 sg13g2_and2_1 _41164_ (.A(net5623),
    .B(_10575_),
    .X(_10576_));
 sg13g2_xnor2_1 _41165_ (.Y(_10577_),
    .A(net5623),
    .B(_10575_));
 sg13g2_nand3_1 _41166_ (.B(_05952_),
    .C(_05956_),
    .A(net6753),
    .Y(_10578_));
 sg13g2_a21oi_1 _41167_ (.A1(_05967_),
    .A2(_10543_),
    .Y(_10579_),
    .B1(_05966_));
 sg13g2_xnor2_1 _41168_ (.Y(_10580_),
    .A(_05959_),
    .B(_10579_));
 sg13g2_o21ai_1 _41169_ (.B1(_10578_),
    .Y(_10581_),
    .A1(net6753),
    .A2(_10580_));
 sg13g2_nand2_1 _41170_ (.Y(_10582_),
    .A(net5623),
    .B(_10581_));
 sg13g2_xnor2_1 _41171_ (.Y(_10583_),
    .A(net5577),
    .B(_10581_));
 sg13g2_xnor2_1 _41172_ (.Y(_10584_),
    .A(_05934_),
    .B(_10572_));
 sg13g2_mux2_1 _41173_ (.A0(_05932_),
    .A1(_10584_),
    .S(net6796),
    .X(_10585_));
 sg13g2_inv_1 _41174_ (.Y(_10586_),
    .A(_10585_));
 sg13g2_xnor2_1 _41175_ (.Y(_10587_),
    .A(net5623),
    .B(_10585_));
 sg13g2_nand2_1 _41176_ (.Y(_10588_),
    .A(_10583_),
    .B(_10587_));
 sg13g2_or3_1 _41177_ (.A(_10570_),
    .B(_10577_),
    .C(_10588_),
    .X(_10589_));
 sg13g2_or3_1 _41178_ (.A(_10534_),
    .B(_10563_),
    .C(_10589_),
    .X(_10590_));
 sg13g2_nand2_1 _41179_ (.Y(_10591_),
    .A(net6747),
    .B(_05715_));
 sg13g2_xnor2_1 _41180_ (.Y(_10592_),
    .A(_05717_),
    .B(_10226_));
 sg13g2_o21ai_1 _41181_ (.B1(_10591_),
    .Y(_10593_),
    .A1(net6747),
    .A2(_10592_));
 sg13g2_xnor2_1 _41182_ (.Y(_10594_),
    .A(net5616),
    .B(_10593_));
 sg13g2_inv_1 _41183_ (.Y(_10595_),
    .A(_10594_));
 sg13g2_nor2_1 _41184_ (.A(net6794),
    .B(_05749_),
    .Y(_10596_));
 sg13g2_o21ai_1 _41185_ (.B1(_05914_),
    .Y(_10597_),
    .A1(_06103_),
    .A2(_10565_));
 sg13g2_nand2_1 _41186_ (.Y(_10598_),
    .A(_06117_),
    .B(_10597_));
 sg13g2_nand2_1 _41187_ (.Y(_10599_),
    .A(_05801_),
    .B(_10598_));
 sg13g2_a21oi_2 _41188_ (.B1(_05813_),
    .Y(_10600_),
    .A2(_10597_),
    .A1(_06117_));
 sg13g2_a21oi_1 _41189_ (.A1(_05792_),
    .A2(_10600_),
    .Y(_10601_),
    .B1(_06107_));
 sg13g2_a21o_1 _41190_ (.A2(_10600_),
    .A1(_05792_),
    .B1(_06107_),
    .X(_10602_));
 sg13g2_a21oi_1 _41191_ (.A1(_05770_),
    .A2(_10602_),
    .Y(_10603_),
    .B1(_06109_));
 sg13g2_o21ai_1 _41192_ (.B1(_05741_),
    .Y(_10604_),
    .A1(_05742_),
    .A2(_10603_));
 sg13g2_xnor2_1 _41193_ (.Y(_10605_),
    .A(_05750_),
    .B(_10604_));
 sg13g2_a21oi_2 _41194_ (.B1(_10596_),
    .Y(_10606_),
    .A2(_10605_),
    .A1(net6795));
 sg13g2_nand2_1 _41195_ (.Y(_10607_),
    .A(net5616),
    .B(_10606_));
 sg13g2_xnor2_1 _41196_ (.Y(_10608_),
    .A(net5572),
    .B(_10606_));
 sg13g2_xnor2_1 _41197_ (.Y(_10609_),
    .A(net5616),
    .B(_10606_));
 sg13g2_nor2_1 _41198_ (.A(net6795),
    .B(_05760_),
    .Y(_10610_));
 sg13g2_o21ai_1 _41199_ (.B1(_05768_),
    .Y(_10611_),
    .A1(_05769_),
    .A2(_10601_));
 sg13g2_xor2_1 _41200_ (.B(_10611_),
    .A(_05762_),
    .X(_10612_));
 sg13g2_a21oi_2 _41201_ (.B1(_10610_),
    .Y(_10613_),
    .A2(_10612_),
    .A1(net6794));
 sg13g2_xnor2_1 _41202_ (.Y(_10614_),
    .A(net5616),
    .B(_10613_));
 sg13g2_nand2_1 _41203_ (.Y(_10615_),
    .A(net6751),
    .B(_05740_));
 sg13g2_xnor2_1 _41204_ (.Y(_10616_),
    .A(_05742_),
    .B(_10603_));
 sg13g2_o21ai_1 _41205_ (.B1(_10615_),
    .Y(_10617_),
    .A1(net6751),
    .A2(_10616_));
 sg13g2_nand2b_1 _41206_ (.Y(_10618_),
    .B(net5572),
    .A_N(_10617_));
 sg13g2_xnor2_1 _41207_ (.Y(_10619_),
    .A(net5572),
    .B(_10617_));
 sg13g2_nor2b_1 _41208_ (.A(_10614_),
    .B_N(_10619_),
    .Y(_10620_));
 sg13g2_nand3_1 _41209_ (.B(_10608_),
    .C(_10620_),
    .A(_10595_),
    .Y(_10621_));
 sg13g2_o21ai_1 _41210_ (.B1(_05791_),
    .Y(_10622_),
    .A1(_06105_),
    .A2(_10600_));
 sg13g2_nand2_1 _41211_ (.Y(_10623_),
    .A(_05790_),
    .B(_10622_));
 sg13g2_nor2_1 _41212_ (.A(net6794),
    .B(_05781_),
    .Y(_10624_));
 sg13g2_xnor2_1 _41213_ (.Y(_10625_),
    .A(_05783_),
    .B(_10623_));
 sg13g2_a21oi_2 _41214_ (.B1(_10624_),
    .Y(_10626_),
    .A2(_10625_),
    .A1(net6794));
 sg13g2_and2_1 _41215_ (.A(net5620),
    .B(_10626_),
    .X(_10627_));
 sg13g2_nor2_1 _41216_ (.A(net5620),
    .B(_10626_),
    .Y(_10628_));
 sg13g2_xnor2_1 _41217_ (.Y(_10629_),
    .A(net5574),
    .B(_10626_));
 sg13g2_nand2_1 _41218_ (.Y(_10630_),
    .A(net6752),
    .B(_05767_));
 sg13g2_xnor2_1 _41219_ (.Y(_10631_),
    .A(_05769_),
    .B(_10601_));
 sg13g2_o21ai_1 _41220_ (.B1(_10630_),
    .Y(_10632_),
    .A1(net6752),
    .A2(_10631_));
 sg13g2_xnor2_1 _41221_ (.Y(_10633_),
    .A(net5620),
    .B(_10632_));
 sg13g2_inv_1 _41222_ (.Y(_10634_),
    .A(_10633_));
 sg13g2_a21oi_1 _41223_ (.A1(_05800_),
    .A2(_10599_),
    .Y(_10635_),
    .B1(_05811_));
 sg13g2_and3_1 _41224_ (.X(_10636_),
    .A(_05800_),
    .B(_05811_),
    .C(_10599_));
 sg13g2_o21ai_1 _41225_ (.B1(net6794),
    .Y(_10637_),
    .A1(_10635_),
    .A2(_10636_));
 sg13g2_o21ai_1 _41226_ (.B1(_10637_),
    .Y(_10638_),
    .A1(net6794),
    .A2(_05809_));
 sg13g2_xnor2_1 _41227_ (.Y(_10639_),
    .A(net5620),
    .B(_10638_));
 sg13g2_or3_1 _41228_ (.A(_05791_),
    .B(_06105_),
    .C(_10600_),
    .X(_10640_));
 sg13g2_a21oi_1 _41229_ (.A1(_10622_),
    .A2(_10640_),
    .Y(_10641_),
    .B1(net6751));
 sg13g2_a21oi_2 _41230_ (.B1(_10641_),
    .Y(_10642_),
    .A2(_05789_),
    .A1(net6751));
 sg13g2_inv_1 _41231_ (.Y(_10643_),
    .A(_10642_));
 sg13g2_xnor2_1 _41232_ (.Y(_10644_),
    .A(net5620),
    .B(_10642_));
 sg13g2_inv_1 _41233_ (.Y(_10645_),
    .A(_10644_));
 sg13g2_and4_1 _41234_ (.A(_10629_),
    .B(_10634_),
    .C(_10639_),
    .D(_10645_),
    .X(_10646_));
 sg13g2_and4_1 _41235_ (.A(_10595_),
    .B(_10608_),
    .C(_10620_),
    .D(_10646_),
    .X(_10647_));
 sg13g2_o21ai_1 _41236_ (.B1(_05912_),
    .Y(_10648_),
    .A1(_06103_),
    .A2(_10565_));
 sg13g2_nand2_1 _41237_ (.Y(_10649_),
    .A(_06113_),
    .B(_10648_));
 sg13g2_nand2_1 _41238_ (.Y(_10650_),
    .A(_05871_),
    .B(_10649_));
 sg13g2_nand2_1 _41239_ (.Y(_10651_),
    .A(_05870_),
    .B(_10650_));
 sg13g2_a221oi_1 _41240_ (.B2(_10648_),
    .C1(_05872_),
    .B1(_06113_),
    .A1(_05861_),
    .Y(_10652_),
    .A2(_05862_));
 sg13g2_nor2_1 _41241_ (.A(_06115_),
    .B(_10652_),
    .Y(_10653_));
 sg13g2_o21ai_1 _41242_ (.B1(_05836_),
    .Y(_10654_),
    .A1(_06115_),
    .A2(_10652_));
 sg13g2_a21oi_1 _41243_ (.A1(_05834_),
    .A2(_10654_),
    .Y(_10655_),
    .B1(_05848_));
 sg13g2_and3_1 _41244_ (.X(_10656_),
    .A(_05834_),
    .B(_05848_),
    .C(_10654_));
 sg13g2_nor3_1 _41245_ (.A(net6751),
    .B(_10655_),
    .C(_10656_),
    .Y(_10657_));
 sg13g2_a21oi_2 _41246_ (.B1(_10657_),
    .Y(_10658_),
    .A2(_05845_),
    .A1(net6751));
 sg13g2_xnor2_1 _41247_ (.Y(_10659_),
    .A(net5619),
    .B(_10658_));
 sg13g2_nand2_1 _41248_ (.Y(_10660_),
    .A(net6751),
    .B(_05799_));
 sg13g2_xnor2_1 _41249_ (.Y(_10661_),
    .A(_05801_),
    .B(_10598_));
 sg13g2_o21ai_1 _41250_ (.B1(_10660_),
    .Y(_10662_),
    .A1(net6751),
    .A2(_10661_));
 sg13g2_xnor2_1 _41251_ (.Y(_10663_),
    .A(net5574),
    .B(_10662_));
 sg13g2_nor2b_1 _41252_ (.A(_10659_),
    .B_N(_10663_),
    .Y(_10664_));
 sg13g2_nand2b_1 _41253_ (.Y(_10665_),
    .B(_10663_),
    .A_N(_10659_));
 sg13g2_nor2_1 _41254_ (.A(net6794),
    .B(_05833_),
    .Y(_10666_));
 sg13g2_xnor2_1 _41255_ (.Y(_10667_),
    .A(_05836_),
    .B(_10653_));
 sg13g2_a21oi_2 _41256_ (.B1(_10666_),
    .Y(_10668_),
    .A2(_10667_),
    .A1(net6794));
 sg13g2_nor2_1 _41257_ (.A(net5574),
    .B(_10668_),
    .Y(_10669_));
 sg13g2_xnor2_1 _41258_ (.Y(_10670_),
    .A(net5618),
    .B(_10668_));
 sg13g2_xnor2_1 _41259_ (.Y(_10671_),
    .A(_05863_),
    .B(_10651_));
 sg13g2_nor2_1 _41260_ (.A(net6754),
    .B(_10671_),
    .Y(_10672_));
 sg13g2_a21oi_2 _41261_ (.B1(_10672_),
    .Y(_10673_),
    .A2(_05858_),
    .A1(net6754));
 sg13g2_nand2_1 _41262_ (.Y(_10674_),
    .A(net5618),
    .B(_10673_));
 sg13g2_xnor2_1 _41263_ (.Y(_10675_),
    .A(net5574),
    .B(_10673_));
 sg13g2_and3_1 _41264_ (.X(_10676_),
    .A(_10664_),
    .B(_10670_),
    .C(_10675_));
 sg13g2_nand2_1 _41265_ (.Y(_10677_),
    .A(net6754),
    .B(_05869_));
 sg13g2_xnor2_1 _41266_ (.Y(_10678_),
    .A(_05871_),
    .B(_10649_));
 sg13g2_o21ai_1 _41267_ (.B1(_10677_),
    .Y(_10679_),
    .A1(net6754),
    .A2(_10678_));
 sg13g2_xnor2_1 _41268_ (.Y(_10680_),
    .A(net5618),
    .B(_10679_));
 sg13g2_nor2_1 _41269_ (.A(net6796),
    .B(_05892_),
    .Y(_10681_));
 sg13g2_o21ai_1 _41270_ (.B1(_06111_),
    .Y(_10682_),
    .A1(_05902_),
    .A2(_10567_));
 sg13g2_a21oi_1 _41271_ (.A1(_05883_),
    .A2(_10682_),
    .Y(_10683_),
    .B1(_05881_));
 sg13g2_xnor2_1 _41272_ (.Y(_10684_),
    .A(_05894_),
    .B(_10683_));
 sg13g2_a21oi_2 _41273_ (.B1(_10681_),
    .Y(_10685_),
    .A2(_10684_),
    .A1(net6796));
 sg13g2_and2_1 _41274_ (.A(net5619),
    .B(_10685_),
    .X(_10686_));
 sg13g2_xnor2_1 _41275_ (.Y(_10687_),
    .A(net5618),
    .B(_10685_));
 sg13g2_nor2_1 _41276_ (.A(_10680_),
    .B(_10687_),
    .Y(_10688_));
 sg13g2_inv_1 _41277_ (.Y(_10689_),
    .A(_10688_));
 sg13g2_nor2_1 _41278_ (.A(net6796),
    .B(_05880_),
    .Y(_10690_));
 sg13g2_xnor2_1 _41279_ (.Y(_10691_),
    .A(_05884_),
    .B(_10682_));
 sg13g2_a21oi_2 _41280_ (.B1(_10690_),
    .Y(_10692_),
    .A2(_10691_),
    .A1(net6796));
 sg13g2_inv_2 _41281_ (.Y(_10693_),
    .A(_10692_));
 sg13g2_xnor2_1 _41282_ (.Y(_10694_),
    .A(net5618),
    .B(_10692_));
 sg13g2_nand2_1 _41283_ (.Y(_10695_),
    .A(_05908_),
    .B(_10567_));
 sg13g2_xnor2_1 _41284_ (.Y(_10696_),
    .A(_05902_),
    .B(_10695_));
 sg13g2_mux2_1 _41285_ (.A0(_05901_),
    .A1(_10696_),
    .S(net6800),
    .X(_10697_));
 sg13g2_nand2_1 _41286_ (.Y(_10698_),
    .A(net5618),
    .B(_10697_));
 sg13g2_xnor2_1 _41287_ (.Y(_10699_),
    .A(net5574),
    .B(_10697_));
 sg13g2_and3_1 _41288_ (.X(_10700_),
    .A(_10688_),
    .B(_10694_),
    .C(_10699_));
 sg13g2_inv_1 _41289_ (.Y(_10701_),
    .A(_10700_));
 sg13g2_and4_1 _41290_ (.A(_10664_),
    .B(_10670_),
    .C(_10675_),
    .D(_10700_),
    .X(_10702_));
 sg13g2_inv_1 _41291_ (.Y(_10703_),
    .A(_10702_));
 sg13g2_and2_1 _41292_ (.A(_10647_),
    .B(_10702_),
    .X(_10704_));
 sg13g2_nor2b_1 _41293_ (.A(_10590_),
    .B_N(_10704_),
    .Y(_10705_));
 sg13g2_inv_1 _41294_ (.Y(_10706_),
    .A(_10705_));
 sg13g2_nand3_1 _41295_ (.B(_10469_),
    .C(_10705_),
    .A(_10355_),
    .Y(_10707_));
 sg13g2_a21o_1 _41296_ (.A2(net5475),
    .A1(net5476),
    .B1(_10707_),
    .X(_10708_));
 sg13g2_o21ai_1 _41297_ (.B1(net5627),
    .Y(_10709_),
    .A1(_10524_),
    .A2(_10529_));
 sg13g2_o21ai_1 _41298_ (.B1(_10525_),
    .Y(_10710_),
    .A1(net5578),
    .A2(_10530_));
 sg13g2_a221oi_1 _41299_ (.B2(_10710_),
    .C1(_10517_),
    .B1(_10521_),
    .A1(net5625),
    .Y(_10711_),
    .A2(_10505_));
 sg13g2_nor4_1 _41300_ (.A(_10482_),
    .B(_10491_),
    .C(_10501_),
    .D(_10711_),
    .Y(_10712_));
 sg13g2_o21ai_1 _41301_ (.B1(net5626),
    .Y(_10713_),
    .A1(_10494_),
    .A2(_10499_));
 sg13g2_inv_1 _41302_ (.Y(_10714_),
    .A(_10713_));
 sg13g2_nor3_1 _41303_ (.A(_10482_),
    .B(_10491_),
    .C(_10713_),
    .Y(_10715_));
 sg13g2_nor4_1 _41304_ (.A(_10480_),
    .B(_10490_),
    .C(_10712_),
    .D(_10715_),
    .Y(_10716_));
 sg13g2_inv_1 _41305_ (.Y(_10717_),
    .A(_10716_));
 sg13g2_nor3_1 _41306_ (.A(_10563_),
    .B(_10589_),
    .C(_10716_),
    .Y(_10718_));
 sg13g2_o21ai_1 _41307_ (.B1(_10582_),
    .Y(_10719_),
    .A1(net5580),
    .A2(_10585_));
 sg13g2_inv_1 _41308_ (.Y(_10720_),
    .A(_10719_));
 sg13g2_nor3_1 _41309_ (.A(_10570_),
    .B(_10577_),
    .C(_10720_),
    .Y(_10721_));
 sg13g2_a21o_1 _41310_ (.A2(_10569_),
    .A1(net5623),
    .B1(_10576_),
    .X(_10722_));
 sg13g2_o21ai_1 _41311_ (.B1(_10559_),
    .Y(_10723_),
    .A1(net5577),
    .A2(_10553_));
 sg13g2_inv_1 _41312_ (.Y(_10724_),
    .A(_10723_));
 sg13g2_o21ai_1 _41313_ (.B1(net5624),
    .Y(_10725_),
    .A1(_10540_),
    .A2(_10546_));
 sg13g2_o21ai_1 _41314_ (.B1(_10725_),
    .Y(_10726_),
    .A1(_10549_),
    .A2(_10724_));
 sg13g2_nor2b_1 _41315_ (.A(_10589_),
    .B_N(_10726_),
    .Y(_10727_));
 sg13g2_nor4_2 _41316_ (.A(_10718_),
    .B(_10721_),
    .C(_10722_),
    .Y(_10728_),
    .D(_10727_));
 sg13g2_inv_1 _41317_ (.Y(_10729_),
    .A(_10728_));
 sg13g2_nand2b_1 _41318_ (.Y(_10730_),
    .B(_10704_),
    .A_N(_10728_));
 sg13g2_a21o_1 _41319_ (.A2(_10643_),
    .A1(_10638_),
    .B1(net5574),
    .X(_10731_));
 sg13g2_nor4_1 _41320_ (.A(_10627_),
    .B(_10628_),
    .C(_10633_),
    .D(_10731_),
    .Y(_10732_));
 sg13g2_o21ai_1 _41321_ (.B1(net5620),
    .Y(_10733_),
    .A1(_10626_),
    .A2(_10632_));
 sg13g2_nor2b_1 _41322_ (.A(_10732_),
    .B_N(_10733_),
    .Y(_10734_));
 sg13g2_nor2_1 _41323_ (.A(_10621_),
    .B(_10734_),
    .Y(_10735_));
 sg13g2_o21ai_1 _41324_ (.B1(net5616),
    .Y(_10736_),
    .A1(_10613_),
    .A2(_10617_));
 sg13g2_inv_1 _41325_ (.Y(_10737_),
    .A(_10736_));
 sg13g2_nor3_1 _41326_ (.A(_10594_),
    .B(_10609_),
    .C(_10736_),
    .Y(_10738_));
 sg13g2_o21ai_1 _41327_ (.B1(net5616),
    .Y(_10739_),
    .A1(_10593_),
    .A2(_10606_));
 sg13g2_nand2b_1 _41328_ (.Y(_10740_),
    .B(_10739_),
    .A_N(_10738_));
 sg13g2_nor2_1 _41329_ (.A(_10735_),
    .B(_10740_),
    .Y(_10741_));
 sg13g2_o21ai_1 _41330_ (.B1(net5618),
    .Y(_10742_),
    .A1(_10693_),
    .A2(_10697_));
 sg13g2_o21ai_1 _41331_ (.B1(net5619),
    .Y(_10743_),
    .A1(_10679_),
    .A2(_10685_));
 sg13g2_o21ai_1 _41332_ (.B1(_10743_),
    .Y(_10744_),
    .A1(_10689_),
    .A2(_10742_));
 sg13g2_a21oi_1 _41333_ (.A1(net5618),
    .A2(_10673_),
    .Y(_10745_),
    .B1(_10669_));
 sg13g2_o21ai_1 _41334_ (.B1(net5619),
    .Y(_10746_),
    .A1(_10658_),
    .A2(_10662_));
 sg13g2_o21ai_1 _41335_ (.B1(_10746_),
    .Y(_10747_),
    .A1(_10665_),
    .A2(_10745_));
 sg13g2_a21o_2 _41336_ (.A2(_10744_),
    .A1(_10676_),
    .B1(_10747_),
    .X(_10748_));
 sg13g2_nand2_1 _41337_ (.Y(_10749_),
    .A(_10647_),
    .B(_10748_));
 sg13g2_nand3_1 _41338_ (.B(_10741_),
    .C(_10749_),
    .A(_10730_),
    .Y(_10750_));
 sg13g2_o21ai_1 _41339_ (.B1(net5614),
    .Y(_10751_),
    .A1(_10457_),
    .A2(_10463_));
 sg13g2_nor2_1 _41340_ (.A(_10454_),
    .B(_10751_),
    .Y(_10752_));
 sg13g2_o21ai_1 _41341_ (.B1(net5615),
    .Y(_10753_),
    .A1(_10444_),
    .A2(_10450_));
 sg13g2_nor2b_1 _41342_ (.A(_10752_),
    .B_N(_10753_),
    .Y(_10754_));
 sg13g2_o21ai_1 _41343_ (.B1(_10753_),
    .Y(_10755_),
    .A1(_10454_),
    .A2(_10751_));
 sg13g2_nand2b_1 _41344_ (.Y(_10756_),
    .B(_10437_),
    .A_N(_10430_));
 sg13g2_a21o_1 _41345_ (.A2(_10424_),
    .A1(net5614),
    .B1(_10420_),
    .X(_10757_));
 sg13g2_a221oi_1 _41346_ (.B2(_10426_),
    .C1(_10757_),
    .B1(_10756_),
    .A1(_10441_),
    .Y(_10758_),
    .A2(_10755_));
 sg13g2_inv_1 _41347_ (.Y(_10759_),
    .A(_10758_));
 sg13g2_or3_1 _41348_ (.A(_10383_),
    .B(_10408_),
    .C(_10758_),
    .X(_10760_));
 sg13g2_o21ai_1 _41349_ (.B1(net5615),
    .Y(_10761_),
    .A1(_10400_),
    .A2(_10405_));
 sg13g2_o21ai_1 _41350_ (.B1(net5615),
    .Y(_10762_),
    .A1(_10389_),
    .A2(_10394_));
 sg13g2_o21ai_1 _41351_ (.B1(_10762_),
    .Y(_10763_),
    .A1(_10396_),
    .A2(_10761_));
 sg13g2_nand2b_1 _41352_ (.Y(_10764_),
    .B(_10763_),
    .A_N(_10383_));
 sg13g2_o21ai_1 _41353_ (.B1(net5617),
    .Y(_10765_),
    .A1(_10374_),
    .A2(_10380_));
 sg13g2_nand3b_1 _41354_ (.B(_10370_),
    .C(_10366_),
    .Y(_10766_),
    .A_N(_10765_));
 sg13g2_o21ai_1 _41355_ (.B1(net5617),
    .Y(_10767_),
    .A1(_10364_),
    .A2(_10369_));
 sg13g2_nand4_1 _41356_ (.B(_10764_),
    .C(_10766_),
    .A(_10760_),
    .Y(_10768_),
    .D(_10767_));
 sg13g2_o21ai_1 _41357_ (.B1(net5612),
    .Y(_10769_),
    .A1(_10319_),
    .A2(_10325_));
 sg13g2_nor4_1 _41358_ (.A(_10308_),
    .B(_10309_),
    .C(_10316_),
    .D(_10769_),
    .Y(_10770_));
 sg13g2_a21oi_1 _41359_ (.A1(net5612),
    .A2(_10315_),
    .Y(_10771_),
    .B1(_10770_));
 sg13g2_nand2b_1 _41360_ (.Y(_10772_),
    .B(_10771_),
    .A_N(_10308_));
 sg13g2_o21ai_1 _41361_ (.B1(net5611),
    .Y(_10773_),
    .A1(_10345_),
    .A2(_10351_));
 sg13g2_nor3_1 _41362_ (.A(_10334_),
    .B(_10341_),
    .C(_10773_),
    .Y(_10774_));
 sg13g2_a21oi_1 _41363_ (.A1(_10353_),
    .A2(_10772_),
    .Y(_10775_),
    .B1(_10774_));
 sg13g2_and3_1 _41364_ (.X(_10776_),
    .A(_10333_),
    .B(_10340_),
    .C(_10775_));
 sg13g2_o21ai_1 _41365_ (.B1(net5610),
    .Y(_10777_),
    .A1(_10253_),
    .A2(_10259_));
 sg13g2_or4_1 _41366_ (.A(_10239_),
    .B(_10240_),
    .C(_10249_),
    .D(_10777_),
    .X(_10778_));
 sg13g2_nand2_1 _41367_ (.Y(_10779_),
    .A(_10248_),
    .B(_10778_));
 sg13g2_nor2_1 _41368_ (.A(_10239_),
    .B(_10779_),
    .Y(_10780_));
 sg13g2_or2_1 _41369_ (.X(_10781_),
    .B(_10779_),
    .A(_10239_));
 sg13g2_nand2_1 _41370_ (.Y(_10782_),
    .A(_10285_),
    .B(_10294_));
 sg13g2_a21oi_1 _41371_ (.A1(net5608),
    .A2(_10266_),
    .Y(_10783_),
    .B1(net5683));
 sg13g2_nand2b_1 _41372_ (.Y(_10784_),
    .B(_10783_),
    .A_N(_10275_));
 sg13g2_a221oi_1 _41373_ (.B2(_10278_),
    .C1(_10784_),
    .B1(_10782_),
    .A1(_10297_),
    .Y(_10785_),
    .A2(_10781_));
 sg13g2_o21ai_1 _41374_ (.B1(_10785_),
    .Y(_10786_),
    .A1(_10298_),
    .A2(_10776_));
 sg13g2_a221oi_1 _41375_ (.B2(_10355_),
    .C1(_10786_),
    .B1(_10768_),
    .A1(_10470_),
    .Y(_10787_),
    .A2(_10750_));
 sg13g2_a22oi_1 _41376_ (.Y(_10788_),
    .B1(_10708_),
    .B2(_10787_),
    .A2(net5616),
    .A1(net5688));
 sg13g2_a21o_2 _41377_ (.A2(_10787_),
    .A1(_10708_),
    .B1(_08584_),
    .X(_10789_));
 sg13g2_xnor2_1 _41378_ (.Y(_10790_),
    .A(_08581_),
    .B(_09147_));
 sg13g2_inv_1 _41379_ (.Y(_10791_),
    .A(_10790_));
 sg13g2_o21ai_1 _41380_ (.B1(_10790_),
    .Y(_10792_),
    .A1(net5556),
    .A2(net5390));
 sg13g2_nand3_1 _41381_ (.B(_09147_),
    .C(net5445),
    .A(net5495),
    .Y(_10793_));
 sg13g2_nand3_1 _41382_ (.B(_10792_),
    .C(_10793_),
    .A(net5943),
    .Y(_10794_));
 sg13g2_a22oi_1 _41383_ (.Y(_10795_),
    .B1(net5495),
    .B2(net5892),
    .A2(net5748),
    .A1(net5977));
 sg13g2_nand2_1 _41384_ (.Y(_10796_),
    .A(_10794_),
    .B(_10795_));
 sg13g2_a21oi_1 _41385_ (.A1(net5260),
    .A2(_10796_),
    .Y(_10797_),
    .B1(net6842));
 sg13g2_o21ai_1 _41386_ (.B1(_10797_),
    .Y(_10798_),
    .A1(net5257),
    .A2(net5699));
 sg13g2_o21ai_1 _41387_ (.B1(_10798_),
    .Y(_10799_),
    .A1(net2703),
    .A2(net6487));
 sg13g2_inv_1 _41388_ (.Y(_00737_),
    .A(_10799_));
 sg13g2_nand2_1 _41389_ (.Y(_10800_),
    .A(net1680),
    .B(net6403));
 sg13g2_nand2_1 _41390_ (.Y(_10801_),
    .A(_09151_),
    .B(_09158_));
 sg13g2_xnor2_1 _41391_ (.Y(_10802_),
    .A(_09155_),
    .B(_10801_));
 sg13g2_nor2_1 _41392_ (.A(net5699),
    .B(_10802_),
    .Y(_10803_));
 sg13g2_a21oi_1 _41393_ (.A1(net5699),
    .A2(_09154_),
    .Y(_10804_),
    .B1(_10803_));
 sg13g2_inv_2 _41394_ (.Y(_10805_),
    .A(_10804_));
 sg13g2_xnor2_1 _41395_ (.Y(_10806_),
    .A(_10793_),
    .B(_10805_));
 sg13g2_nor2_1 _41396_ (.A(net5241),
    .B(_08580_),
    .Y(_10807_));
 sg13g2_a221oi_1 _41397_ (.B2(net5225),
    .C1(_10807_),
    .B1(_10806_),
    .A1(net5203),
    .Y(_10808_),
    .A2(_10791_));
 sg13g2_o21ai_1 _41398_ (.B1(_10800_),
    .Y(_00738_),
    .A1(net6842),
    .A2(_10808_));
 sg13g2_nand2_1 _41399_ (.Y(_10809_),
    .A(net5699),
    .B(_09163_));
 sg13g2_xor2_1 _41400_ (.B(_09165_),
    .A(_09160_),
    .X(_10810_));
 sg13g2_o21ai_1 _41401_ (.B1(_10809_),
    .Y(_10811_),
    .A1(net5699),
    .A2(_10810_));
 sg13g2_nand2_1 _41402_ (.Y(_10812_),
    .A(net5383),
    .B(_10811_));
 sg13g2_nor2_1 _41403_ (.A(net5383),
    .B(_10811_),
    .Y(_10813_));
 sg13g2_xnor2_1 _41404_ (.Y(_10814_),
    .A(net5383),
    .B(_10811_));
 sg13g2_nor3_1 _41405_ (.A(net5556),
    .B(_10790_),
    .C(_10804_),
    .Y(_10815_));
 sg13g2_nor3_1 _41406_ (.A(net5495),
    .B(_10791_),
    .C(_10805_),
    .Y(_10816_));
 sg13g2_inv_1 _41407_ (.Y(_10817_),
    .A(_10816_));
 sg13g2_o21ai_1 _41408_ (.B1(_10817_),
    .Y(_10818_),
    .A1(net5383),
    .A2(_10815_));
 sg13g2_xnor2_1 _41409_ (.Y(_10819_),
    .A(_10814_),
    .B(_10818_));
 sg13g2_o21ai_1 _41410_ (.B1(net5943),
    .Y(_10820_),
    .A1(net5495),
    .A2(_10811_));
 sg13g2_a21oi_1 _41411_ (.A1(net5495),
    .A2(_10819_),
    .Y(_10821_),
    .B1(_10820_));
 sg13g2_a221oi_1 _41412_ (.B2(net5892),
    .C1(_10821_),
    .B1(_10805_),
    .A1(net5977),
    .Y(_10822_),
    .A2(_09147_));
 sg13g2_o21ai_1 _41413_ (.B1(net6875),
    .Y(_10823_),
    .A1(net5260),
    .A2(_09147_));
 sg13g2_a21oi_1 _41414_ (.A1(net5260),
    .A2(_10822_),
    .Y(_10824_),
    .B1(_10823_));
 sg13g2_a21o_1 _41415_ (.A2(net6403),
    .A1(net2514),
    .B1(_10824_),
    .X(_00739_));
 sg13g2_a21o_1 _41416_ (.A2(_09163_),
    .A1(net5580),
    .B1(_09166_),
    .X(_10825_));
 sg13g2_xnor2_1 _41417_ (.Y(_10826_),
    .A(_09143_),
    .B(_10825_));
 sg13g2_nand2_1 _41418_ (.Y(_10827_),
    .A(net5748),
    .B(_10826_));
 sg13g2_o21ai_1 _41419_ (.B1(_10827_),
    .Y(_10828_),
    .A1(net5748),
    .A2(_09141_));
 sg13g2_inv_1 _41420_ (.Y(_10829_),
    .A(_10828_));
 sg13g2_xnor2_1 _41421_ (.Y(_10830_),
    .A(net5445),
    .B(_10829_));
 sg13g2_a21oi_2 _41422_ (.B1(_10813_),
    .Y(_10831_),
    .A2(_10818_),
    .A1(_10812_));
 sg13g2_nand2_1 _41423_ (.Y(_10832_),
    .A(_10830_),
    .B(_10831_));
 sg13g2_xor2_1 _41424_ (.B(_10831_),
    .A(_10830_),
    .X(_10833_));
 sg13g2_nor2_1 _41425_ (.A(net5556),
    .B(_10833_),
    .Y(_10834_));
 sg13g2_a21oi_1 _41426_ (.A1(net5556),
    .A2(_10829_),
    .Y(_10835_),
    .B1(_10834_));
 sg13g2_a22oi_1 _41427_ (.Y(_10836_),
    .B1(_10835_),
    .B2(net5225),
    .A2(_10811_),
    .A1(net5203));
 sg13g2_a22oi_1 _41428_ (.Y(_10837_),
    .B1(net5097),
    .B2(_09154_),
    .A2(net6403),
    .A1(net2974));
 sg13g2_o21ai_1 _41429_ (.B1(_10837_),
    .Y(_00740_),
    .A1(net6842),
    .A2(_10836_));
 sg13g2_o21ai_1 _41430_ (.B1(_10832_),
    .Y(_10838_),
    .A1(net5383),
    .A2(_10829_));
 sg13g2_o21ai_1 _41431_ (.B1(_09142_),
    .Y(_10839_),
    .A1(_09166_),
    .A2(_09169_));
 sg13g2_nor2_1 _41432_ (.A(_09137_),
    .B(_10839_),
    .Y(_10840_));
 sg13g2_a21oi_1 _41433_ (.A1(_09137_),
    .A2(_10839_),
    .Y(_10841_),
    .B1(net5699));
 sg13g2_nand2b_1 _41434_ (.Y(_10842_),
    .B(_10841_),
    .A_N(_10840_));
 sg13g2_o21ai_1 _41435_ (.B1(_10842_),
    .Y(_10843_),
    .A1(net5748),
    .A2(_09135_));
 sg13g2_xnor2_1 _41436_ (.Y(_10844_),
    .A(net5445),
    .B(_10843_));
 sg13g2_xnor2_1 _41437_ (.Y(_10845_),
    .A(net5383),
    .B(_10843_));
 sg13g2_o21ai_1 _41438_ (.B1(net5495),
    .Y(_10846_),
    .A1(_10838_),
    .A2(_10845_));
 sg13g2_a21oi_1 _41439_ (.A1(_10838_),
    .A2(_10845_),
    .Y(_10847_),
    .B1(_10846_));
 sg13g2_o21ai_1 _41440_ (.B1(net5943),
    .Y(_10848_),
    .A1(net5495),
    .A2(_10843_));
 sg13g2_nor2_1 _41441_ (.A(_10847_),
    .B(_10848_),
    .Y(_10849_));
 sg13g2_a221oi_1 _41442_ (.B2(net5892),
    .C1(_10849_),
    .B1(_10828_),
    .A1(net5977),
    .Y(_10850_),
    .A2(_09163_));
 sg13g2_o21ai_1 _41443_ (.B1(net6875),
    .Y(_10851_),
    .A1(net5260),
    .A2(_09163_));
 sg13g2_a21oi_1 _41444_ (.A1(net5260),
    .A2(_10850_),
    .Y(_10852_),
    .B1(_10851_));
 sg13g2_a21o_1 _41445_ (.A2(net6403),
    .A1(net2819),
    .B1(_10852_),
    .X(_00741_));
 sg13g2_nor2_1 _41446_ (.A(net5748),
    .B(_09128_),
    .Y(_10853_));
 sg13g2_nor2_1 _41447_ (.A(_09136_),
    .B(_10840_),
    .Y(_10854_));
 sg13g2_xor2_1 _41448_ (.B(_10854_),
    .A(_09130_),
    .X(_10855_));
 sg13g2_a21oi_2 _41449_ (.B1(_10853_),
    .Y(_10856_),
    .A2(_10855_),
    .A1(net5748));
 sg13g2_nand2b_1 _41450_ (.Y(_10857_),
    .B(net5445),
    .A_N(_10856_));
 sg13g2_xnor2_1 _41451_ (.Y(_10858_),
    .A(net5383),
    .B(_10856_));
 sg13g2_o21ai_1 _41452_ (.B1(_10843_),
    .Y(_10859_),
    .A1(net5383),
    .A2(_10828_));
 sg13g2_o21ai_1 _41453_ (.B1(_10859_),
    .Y(_10860_),
    .A1(_10832_),
    .A2(_10845_));
 sg13g2_nand2b_1 _41454_ (.Y(_10861_),
    .B(_10860_),
    .A_N(_10858_));
 sg13g2_xnor2_1 _41455_ (.Y(_10862_),
    .A(_10858_),
    .B(_10860_));
 sg13g2_nor2_1 _41456_ (.A(net5556),
    .B(_10862_),
    .Y(_10863_));
 sg13g2_a21oi_1 _41457_ (.A1(net5556),
    .A2(_10856_),
    .Y(_10864_),
    .B1(_10863_));
 sg13g2_a22oi_1 _41458_ (.Y(_10865_),
    .B1(_10864_),
    .B2(net5225),
    .A2(_10843_),
    .A1(net5203));
 sg13g2_nor2_1 _41459_ (.A(net6842),
    .B(_10865_),
    .Y(_10866_));
 sg13g2_a21oi_1 _41460_ (.A1(net2464),
    .A2(net6403),
    .Y(_10867_),
    .B1(_10866_));
 sg13g2_o21ai_1 _41461_ (.B1(_10867_),
    .Y(_00742_),
    .A1(net5066),
    .A2(_09141_));
 sg13g2_nand2_1 _41462_ (.Y(_10868_),
    .A(net5700),
    .B(_09227_));
 sg13g2_xnor2_1 _41463_ (.Y(_10869_),
    .A(_09171_),
    .B(_09230_));
 sg13g2_o21ai_1 _41464_ (.B1(_10868_),
    .Y(_10870_),
    .A1(net5700),
    .A2(_10869_));
 sg13g2_inv_2 _41465_ (.Y(_10871_),
    .A(_10870_));
 sg13g2_nand2_1 _41466_ (.Y(_10872_),
    .A(net5445),
    .B(_10871_));
 sg13g2_xnor2_1 _41467_ (.Y(_10873_),
    .A(net5390),
    .B(_10871_));
 sg13g2_nand2_1 _41468_ (.Y(_10874_),
    .A(_10857_),
    .B(_10861_));
 sg13g2_xor2_1 _41469_ (.B(_10874_),
    .A(_10873_),
    .X(_10875_));
 sg13g2_a21oi_1 _41470_ (.A1(net5559),
    .A2(_10870_),
    .Y(_10876_),
    .B1(net5923));
 sg13g2_o21ai_1 _41471_ (.B1(_10876_),
    .Y(_10877_),
    .A1(net5556),
    .A2(_10875_));
 sg13g2_nand2b_1 _41472_ (.Y(_10878_),
    .B(net5977),
    .A_N(_09135_));
 sg13g2_nand2b_1 _41473_ (.Y(_10879_),
    .B(net5892),
    .A_N(_10856_));
 sg13g2_nand4_1 _41474_ (.B(_10877_),
    .C(_10878_),
    .A(net5260),
    .Y(_10880_),
    .D(_10879_));
 sg13g2_nor2b_1 _41475_ (.A(net5260),
    .B_N(_09135_),
    .Y(_10881_));
 sg13g2_nor2_1 _41476_ (.A(net6842),
    .B(_10881_),
    .Y(_10882_));
 sg13g2_a22oi_1 _41477_ (.Y(_10883_),
    .B1(_10880_),
    .B2(_10882_),
    .A2(net6403),
    .A1(net2805));
 sg13g2_inv_1 _41478_ (.Y(_00743_),
    .A(_10883_));
 sg13g2_a21oi_1 _41479_ (.A1(_09172_),
    .A2(_09230_),
    .Y(_10884_),
    .B1(_09229_));
 sg13g2_a21oi_1 _41480_ (.A1(net5632),
    .A2(_09220_),
    .Y(_10885_),
    .B1(_10884_));
 sg13g2_xnor2_1 _41481_ (.Y(_10886_),
    .A(_09223_),
    .B(_10884_));
 sg13g2_nand2_1 _41482_ (.Y(_10887_),
    .A(net5750),
    .B(_10886_));
 sg13g2_o21ai_1 _41483_ (.B1(_10887_),
    .Y(_10888_),
    .A1(net5750),
    .A2(_09220_));
 sg13g2_nor2_1 _41484_ (.A(net5499),
    .B(_10888_),
    .Y(_10889_));
 sg13g2_nand2_1 _41485_ (.Y(_10890_),
    .A(net5446),
    .B(_10888_));
 sg13g2_xnor2_1 _41486_ (.Y(_10891_),
    .A(net5446),
    .B(_10888_));
 sg13g2_nor2b_1 _41487_ (.A(_10858_),
    .B_N(_10873_),
    .Y(_10892_));
 sg13g2_nand4_1 _41488_ (.B(_10831_),
    .C(_10844_),
    .A(_10830_),
    .Y(_10893_),
    .D(_10892_));
 sg13g2_nand2b_1 _41489_ (.Y(_10894_),
    .B(_10892_),
    .A_N(_10859_));
 sg13g2_nand4_1 _41490_ (.B(_10872_),
    .C(_10893_),
    .A(_10857_),
    .Y(_10895_),
    .D(_10894_));
 sg13g2_nand2b_1 _41491_ (.Y(_10896_),
    .B(_10895_),
    .A_N(_10891_));
 sg13g2_xor2_1 _41492_ (.B(_10895_),
    .A(_10891_),
    .X(_10897_));
 sg13g2_a21oi_1 _41493_ (.A1(net5499),
    .A2(_10897_),
    .Y(_10898_),
    .B1(_10889_));
 sg13g2_a22oi_1 _41494_ (.Y(_10899_),
    .B1(_10898_),
    .B2(net5225),
    .A2(_10871_),
    .A1(net5203));
 sg13g2_a22oi_1 _41495_ (.Y(_10900_),
    .B1(net5097),
    .B2(_09129_),
    .A2(net6411),
    .A1(net2736));
 sg13g2_o21ai_1 _41496_ (.B1(_10900_),
    .Y(_00744_),
    .A1(net6842),
    .A2(_10899_));
 sg13g2_and2_1 _41497_ (.A(_10890_),
    .B(_10896_),
    .X(_10901_));
 sg13g2_nor2_1 _41498_ (.A(net5750),
    .B(_09209_),
    .Y(_10902_));
 sg13g2_o21ai_1 _41499_ (.B1(_09211_),
    .Y(_10903_),
    .A1(_09222_),
    .A2(_10885_));
 sg13g2_or3_1 _41500_ (.A(_09211_),
    .B(_09222_),
    .C(_10885_),
    .X(_10904_));
 sg13g2_nand2_1 _41501_ (.Y(_10905_),
    .A(_10903_),
    .B(_10904_));
 sg13g2_a21oi_2 _41502_ (.B1(_10902_),
    .Y(_10906_),
    .A2(_10905_),
    .A1(net5750));
 sg13g2_nor2_1 _41503_ (.A(net5446),
    .B(_10906_),
    .Y(_10907_));
 sg13g2_xnor2_1 _41504_ (.Y(_10908_),
    .A(net5446),
    .B(_10906_));
 sg13g2_xnor2_1 _41505_ (.Y(_10909_),
    .A(_10901_),
    .B(_10908_));
 sg13g2_o21ai_1 _41506_ (.B1(net5947),
    .Y(_10910_),
    .A1(net5499),
    .A2(_10906_));
 sg13g2_a21oi_1 _41507_ (.A1(net5499),
    .A2(_10909_),
    .Y(_10911_),
    .B1(_10910_));
 sg13g2_a221oi_1 _41508_ (.B2(net5897),
    .C1(_10911_),
    .B1(_10888_),
    .A1(net5981),
    .Y(_10912_),
    .A2(_09228_));
 sg13g2_o21ai_1 _41509_ (.B1(net6875),
    .Y(_10913_),
    .A1(net5258),
    .A2(_09228_));
 sg13g2_a21oi_1 _41510_ (.A1(net5258),
    .A2(_10912_),
    .Y(_10914_),
    .B1(_10913_));
 sg13g2_a21o_1 _41511_ (.A2(net6411),
    .A1(net1823),
    .B1(_10914_),
    .X(_00745_));
 sg13g2_nand2_1 _41512_ (.Y(_10915_),
    .A(_09210_),
    .B(_10903_));
 sg13g2_xnor2_1 _41513_ (.Y(_10916_),
    .A(_09217_),
    .B(_10915_));
 sg13g2_nand2_1 _41514_ (.Y(_10917_),
    .A(net5700),
    .B(_09215_));
 sg13g2_o21ai_1 _41515_ (.B1(_10917_),
    .Y(_10918_),
    .A1(net5700),
    .A2(_10916_));
 sg13g2_nand2_1 _41516_ (.Y(_10919_),
    .A(net5392),
    .B(_10918_));
 sg13g2_xnor2_1 _41517_ (.Y(_10920_),
    .A(net5446),
    .B(_10918_));
 sg13g2_inv_1 _41518_ (.Y(_10921_),
    .A(_10920_));
 sg13g2_o21ai_1 _41519_ (.B1(net5446),
    .Y(_10922_),
    .A1(_10888_),
    .A2(_10906_));
 sg13g2_a21o_1 _41520_ (.A2(_10922_),
    .A1(_10896_),
    .B1(_10907_),
    .X(_10923_));
 sg13g2_xnor2_1 _41521_ (.Y(_10924_),
    .A(_10921_),
    .B(_10923_));
 sg13g2_a21oi_1 _41522_ (.A1(net5497),
    .A2(_10924_),
    .Y(_10925_),
    .B1(net5924));
 sg13g2_o21ai_1 _41523_ (.B1(_10925_),
    .Y(_10926_),
    .A1(net5497),
    .A2(_10918_));
 sg13g2_a22oi_1 _41524_ (.Y(_10927_),
    .B1(_10906_),
    .B2(net5897),
    .A2(_09221_),
    .A1(net5981));
 sg13g2_nand3_1 _41525_ (.B(_10926_),
    .C(_10927_),
    .A(net5258),
    .Y(_10928_));
 sg13g2_nor2_1 _41526_ (.A(net5259),
    .B(_09221_),
    .Y(_10929_));
 sg13g2_nor2_1 _41527_ (.A(net6845),
    .B(_10929_),
    .Y(_10930_));
 sg13g2_a22oi_1 _41528_ (.Y(_10931_),
    .B1(_10928_),
    .B2(_10930_),
    .A2(net6411),
    .A1(net3145));
 sg13g2_inv_1 _41529_ (.Y(_00746_),
    .A(_10931_));
 sg13g2_nand2_1 _41530_ (.Y(_10932_),
    .A(net5700),
    .B(_09192_));
 sg13g2_a21oi_1 _41531_ (.A1(_09172_),
    .A2(_09231_),
    .Y(_10933_),
    .B1(_09235_));
 sg13g2_xnor2_1 _41532_ (.Y(_10934_),
    .A(_09194_),
    .B(_10933_));
 sg13g2_o21ai_1 _41533_ (.B1(_10932_),
    .Y(_10935_),
    .A1(net5700),
    .A2(_10934_));
 sg13g2_xnor2_1 _41534_ (.Y(_10936_),
    .A(net5447),
    .B(_10935_));
 sg13g2_o21ai_1 _41535_ (.B1(_10919_),
    .Y(_10937_),
    .A1(_10921_),
    .A2(_10923_));
 sg13g2_xnor2_1 _41536_ (.Y(_10938_),
    .A(_10936_),
    .B(_10937_));
 sg13g2_o21ai_1 _41537_ (.B1(net5947),
    .Y(_10939_),
    .A1(net5497),
    .A2(_10935_));
 sg13g2_a21oi_1 _41538_ (.A1(net5497),
    .A2(_10938_),
    .Y(_10940_),
    .B1(_10939_));
 sg13g2_a221oi_1 _41539_ (.B2(net5897),
    .C1(_10940_),
    .B1(_10918_),
    .A1(net5981),
    .Y(_10941_),
    .A2(_09209_));
 sg13g2_o21ai_1 _41540_ (.B1(net6875),
    .Y(_10942_),
    .A1(net5258),
    .A2(_09209_));
 sg13g2_a21oi_1 _41541_ (.A1(net5258),
    .A2(_10941_),
    .Y(_10943_),
    .B1(_10942_));
 sg13g2_a21o_1 _41542_ (.A2(net6411),
    .A1(net2977),
    .B1(_10943_),
    .X(_00747_));
 sg13g2_o21ai_1 _41543_ (.B1(_09193_),
    .Y(_10944_),
    .A1(_09194_),
    .A2(_10933_));
 sg13g2_xnor2_1 _41544_ (.Y(_10945_),
    .A(_09201_),
    .B(_10944_));
 sg13g2_o21ai_1 _41545_ (.B1(_10944_),
    .Y(_10946_),
    .A1(net5632),
    .A2(_09199_));
 sg13g2_nor2_1 _41546_ (.A(net5750),
    .B(_09198_),
    .Y(_10947_));
 sg13g2_a21oi_1 _41547_ (.A1(net5750),
    .A2(_10945_),
    .Y(_10948_),
    .B1(_10947_));
 sg13g2_a21o_1 _41548_ (.A2(_10945_),
    .A1(net5750),
    .B1(_10947_),
    .X(_10949_));
 sg13g2_xnor2_1 _41549_ (.Y(_10950_),
    .A(net5392),
    .B(_10948_));
 sg13g2_nand2_1 _41550_ (.Y(_10951_),
    .A(_10920_),
    .B(_10936_));
 sg13g2_nor3_1 _41551_ (.A(_10891_),
    .B(_10908_),
    .C(_10951_),
    .Y(_10952_));
 sg13g2_nand2_1 _41552_ (.Y(_10953_),
    .A(_10895_),
    .B(_10952_));
 sg13g2_nand3b_1 _41553_ (.B(_10936_),
    .C(_10920_),
    .Y(_10954_),
    .A_N(_10922_));
 sg13g2_o21ai_1 _41554_ (.B1(net5392),
    .Y(_10955_),
    .A1(_10918_),
    .A2(_10935_));
 sg13g2_and2_1 _41555_ (.A(_10954_),
    .B(_10955_),
    .X(_10956_));
 sg13g2_nand2_1 _41556_ (.Y(_10957_),
    .A(_10953_),
    .B(_10956_));
 sg13g2_nand2_1 _41557_ (.Y(_10958_),
    .A(_10950_),
    .B(_10957_));
 sg13g2_xnor2_1 _41558_ (.Y(_10959_),
    .A(_10950_),
    .B(_10957_));
 sg13g2_o21ai_1 _41559_ (.B1(net5947),
    .Y(_10960_),
    .A1(net5497),
    .A2(_10949_));
 sg13g2_a21oi_1 _41560_ (.A1(net5497),
    .A2(_10959_),
    .Y(_10961_),
    .B1(_10960_));
 sg13g2_a221oi_1 _41561_ (.B2(net5897),
    .C1(_10961_),
    .B1(_10935_),
    .A1(net5981),
    .Y(_10962_),
    .A2(_09215_));
 sg13g2_o21ai_1 _41562_ (.B1(net6878),
    .Y(_10963_),
    .A1(net5259),
    .A2(_09215_));
 sg13g2_a21oi_1 _41563_ (.A1(net5259),
    .A2(_10962_),
    .Y(_10964_),
    .B1(_10963_));
 sg13g2_a21o_1 _41564_ (.A2(net6410),
    .A1(net1389),
    .B1(_10964_),
    .X(_00748_));
 sg13g2_o21ai_1 _41565_ (.B1(_10958_),
    .Y(_10965_),
    .A1(net5446),
    .A2(_10948_));
 sg13g2_a21o_1 _41566_ (.A2(_10946_),
    .A1(_09200_),
    .B1(_09188_),
    .X(_10966_));
 sg13g2_nand3_1 _41567_ (.B(_09200_),
    .C(_10946_),
    .A(_09188_),
    .Y(_10967_));
 sg13g2_a21oi_1 _41568_ (.A1(_10966_),
    .A2(_10967_),
    .Y(_10968_),
    .B1(net5702));
 sg13g2_a21oi_2 _41569_ (.B1(_10968_),
    .Y(_10969_),
    .A2(_09185_),
    .A1(net5702));
 sg13g2_xnor2_1 _41570_ (.Y(_10970_),
    .A(net5447),
    .B(_10969_));
 sg13g2_xnor2_1 _41571_ (.Y(_10971_),
    .A(_10965_),
    .B(_10970_));
 sg13g2_o21ai_1 _41572_ (.B1(net5947),
    .Y(_10972_),
    .A1(net5498),
    .A2(_10969_));
 sg13g2_a21oi_1 _41573_ (.A1(net5497),
    .A2(_10971_),
    .Y(_10973_),
    .B1(_10972_));
 sg13g2_a221oi_1 _41574_ (.B2(net5897),
    .C1(_10973_),
    .B1(_10949_),
    .A1(net5982),
    .Y(_10974_),
    .A2(_09192_));
 sg13g2_o21ai_1 _41575_ (.B1(net6878),
    .Y(_10975_),
    .A1(net5258),
    .A2(_09192_));
 sg13g2_a21oi_1 _41576_ (.A1(net5259),
    .A2(_10974_),
    .Y(_10976_),
    .B1(_10975_));
 sg13g2_a21o_1 _41577_ (.A2(net6411),
    .A1(net2807),
    .B1(_10976_),
    .X(_00749_));
 sg13g2_nand2_1 _41578_ (.Y(_10977_),
    .A(net2482),
    .B(net6410));
 sg13g2_nor2_1 _41579_ (.A(net5241),
    .B(_09198_),
    .Y(_10978_));
 sg13g2_nand2_1 _41580_ (.Y(_10979_),
    .A(net5700),
    .B(_09176_));
 sg13g2_nand2_1 _41581_ (.Y(_10980_),
    .A(_09187_),
    .B(_10966_));
 sg13g2_xor2_1 _41582_ (.B(_10980_),
    .A(_09178_),
    .X(_10981_));
 sg13g2_o21ai_1 _41583_ (.B1(_10979_),
    .Y(_10982_),
    .A1(net5700),
    .A2(_10981_));
 sg13g2_nor2_1 _41584_ (.A(net5498),
    .B(_10982_),
    .Y(_10983_));
 sg13g2_nand2_1 _41585_ (.Y(_10984_),
    .A(net5392),
    .B(_10982_));
 sg13g2_xnor2_1 _41586_ (.Y(_10985_),
    .A(net5446),
    .B(_10982_));
 sg13g2_inv_1 _41587_ (.Y(_10986_),
    .A(_10985_));
 sg13g2_o21ai_1 _41588_ (.B1(net5392),
    .Y(_10987_),
    .A1(_10949_),
    .A2(_10969_));
 sg13g2_nand2_1 _41589_ (.Y(_10988_),
    .A(_10958_),
    .B(_10987_));
 sg13g2_o21ai_1 _41590_ (.B1(_10988_),
    .Y(_10989_),
    .A1(net5392),
    .A2(_10969_));
 sg13g2_xnor2_1 _41591_ (.Y(_10990_),
    .A(_10986_),
    .B(_10989_));
 sg13g2_a21oi_1 _41592_ (.A1(net5498),
    .A2(_10990_),
    .Y(_10991_),
    .B1(_10983_));
 sg13g2_a221oi_1 _41593_ (.B2(net5226),
    .C1(_10978_),
    .B1(_10991_),
    .A1(net5205),
    .Y(_10992_),
    .A2(_10969_));
 sg13g2_o21ai_1 _41594_ (.B1(_10977_),
    .Y(_00750_),
    .A1(net6845),
    .A2(_10992_));
 sg13g2_nor2_1 _41595_ (.A(net5751),
    .B(_09349_),
    .Y(_10993_));
 sg13g2_a21oi_1 _41596_ (.A1(_09232_),
    .A2(_09238_),
    .Y(_10994_),
    .B1(_09350_));
 sg13g2_xor2_1 _41597_ (.B(_09350_),
    .A(_09239_),
    .X(_10995_));
 sg13g2_a21oi_2 _41598_ (.B1(_10993_),
    .Y(_10996_),
    .A2(_10995_),
    .A1(net5751));
 sg13g2_nand2_1 _41599_ (.Y(_10997_),
    .A(net5392),
    .B(_10996_));
 sg13g2_xnor2_1 _41600_ (.Y(_10998_),
    .A(net5392),
    .B(_10996_));
 sg13g2_o21ai_1 _41601_ (.B1(_10984_),
    .Y(_10999_),
    .A1(_10986_),
    .A2(_10989_));
 sg13g2_xor2_1 _41602_ (.B(_10999_),
    .A(_10998_),
    .X(_11000_));
 sg13g2_o21ai_1 _41603_ (.B1(net5947),
    .Y(_11001_),
    .A1(net5498),
    .A2(_10996_));
 sg13g2_a21oi_1 _41604_ (.A1(net5497),
    .A2(_11000_),
    .Y(_11002_),
    .B1(_11001_));
 sg13g2_a221oi_1 _41605_ (.B2(net5897),
    .C1(_11002_),
    .B1(_10982_),
    .A1(net5981),
    .Y(_11003_),
    .A2(_09186_));
 sg13g2_a21oi_1 _41606_ (.A1(net5258),
    .A2(_11003_),
    .Y(_11004_),
    .B1(net6845));
 sg13g2_o21ai_1 _41607_ (.B1(_11004_),
    .Y(_11005_),
    .A1(net5258),
    .A2(_09186_));
 sg13g2_o21ai_1 _41608_ (.B1(_11005_),
    .Y(_00751_),
    .A1(_18179_),
    .A2(net6488));
 sg13g2_nand2_1 _41609_ (.Y(_11006_),
    .A(net5701),
    .B(_09343_));
 sg13g2_a21o_1 _41610_ (.A2(_09349_),
    .A1(net5635),
    .B1(_10994_),
    .X(_11007_));
 sg13g2_xor2_1 _41611_ (.B(_11007_),
    .A(_09345_),
    .X(_11008_));
 sg13g2_o21ai_1 _41612_ (.B1(_11007_),
    .Y(_11009_),
    .A1(net5633),
    .A2(_09343_));
 sg13g2_o21ai_1 _41613_ (.B1(_11006_),
    .Y(_11010_),
    .A1(net5701),
    .A2(_11008_));
 sg13g2_inv_1 _41614_ (.Y(_11011_),
    .A(_11010_));
 sg13g2_nor2_1 _41615_ (.A(net5501),
    .B(_11010_),
    .Y(_11012_));
 sg13g2_xnor2_1 _41616_ (.Y(_11013_),
    .A(net5393),
    .B(_11011_));
 sg13g2_nor2_1 _41617_ (.A(_10986_),
    .B(_10998_),
    .Y(_11014_));
 sg13g2_nand2_1 _41618_ (.Y(_11015_),
    .A(_10950_),
    .B(_10970_));
 sg13g2_inv_1 _41619_ (.Y(_11016_),
    .A(_11015_));
 sg13g2_nand4_1 _41620_ (.B(_10952_),
    .C(_11014_),
    .A(_10895_),
    .Y(_11017_),
    .D(_11016_));
 sg13g2_o21ai_1 _41621_ (.B1(_10987_),
    .Y(_11018_),
    .A1(_10956_),
    .A2(_11015_));
 sg13g2_nand2_1 _41622_ (.Y(_11019_),
    .A(_10984_),
    .B(_10997_));
 sg13g2_a21oi_1 _41623_ (.A1(_11014_),
    .A2(_11018_),
    .Y(_11020_),
    .B1(_11019_));
 sg13g2_nand2_2 _41624_ (.Y(_11021_),
    .A(_11017_),
    .B(_11020_));
 sg13g2_nand2_1 _41625_ (.Y(_11022_),
    .A(_11013_),
    .B(_11021_));
 sg13g2_xnor2_1 _41626_ (.Y(_11023_),
    .A(_11013_),
    .B(_11021_));
 sg13g2_a21oi_1 _41627_ (.A1(net5501),
    .A2(_11023_),
    .Y(_11024_),
    .B1(_11012_));
 sg13g2_a22oi_1 _41628_ (.Y(_11025_),
    .B1(_11024_),
    .B2(net5226),
    .A2(_10996_),
    .A1(net5205));
 sg13g2_a22oi_1 _41629_ (.Y(_11026_),
    .B1(net5098),
    .B2(_09176_),
    .A2(net6412),
    .A1(net2797));
 sg13g2_o21ai_1 _41630_ (.B1(_11026_),
    .Y(_00752_),
    .A1(net6845),
    .A2(_11025_));
 sg13g2_o21ai_1 _41631_ (.B1(_11022_),
    .Y(_11027_),
    .A1(net5447),
    .A2(_11011_));
 sg13g2_a21oi_1 _41632_ (.A1(_09344_),
    .A2(_11009_),
    .Y(_11028_),
    .B1(_09340_));
 sg13g2_and3_1 _41633_ (.X(_11029_),
    .A(_09340_),
    .B(_09344_),
    .C(_11009_));
 sg13g2_nor3_1 _41634_ (.A(net5701),
    .B(_11028_),
    .C(_11029_),
    .Y(_11030_));
 sg13g2_a21o_2 _41635_ (.A2(_09339_),
    .A1(net5701),
    .B1(_11030_),
    .X(_11031_));
 sg13g2_inv_1 _41636_ (.Y(_11032_),
    .A(_11031_));
 sg13g2_xnor2_1 _41637_ (.Y(_11033_),
    .A(net5393),
    .B(_11031_));
 sg13g2_xor2_1 _41638_ (.B(_11033_),
    .A(_11027_),
    .X(_11034_));
 sg13g2_o21ai_1 _41639_ (.B1(net5951),
    .Y(_11035_),
    .A1(net5501),
    .A2(_11031_));
 sg13g2_a21oi_1 _41640_ (.A1(net5501),
    .A2(_11034_),
    .Y(_11036_),
    .B1(_11035_));
 sg13g2_a221oi_1 _41641_ (.B2(net5897),
    .C1(_11036_),
    .B1(_11010_),
    .A1(net5981),
    .Y(_11037_),
    .A2(_09349_));
 sg13g2_o21ai_1 _41642_ (.B1(net6878),
    .Y(_11038_),
    .A1(net5267),
    .A2(_09349_));
 sg13g2_a21oi_1 _41643_ (.A1(net5270),
    .A2(_11037_),
    .Y(_11039_),
    .B1(_11038_));
 sg13g2_a21o_1 _41644_ (.A2(net6412),
    .A1(net3078),
    .B1(_11039_),
    .X(_00753_));
 sg13g2_nand2_1 _41645_ (.Y(_11040_),
    .A(net2968),
    .B(net6412));
 sg13g2_a21oi_1 _41646_ (.A1(net5635),
    .A2(_09339_),
    .Y(_11041_),
    .B1(_11028_));
 sg13g2_xor2_1 _41647_ (.B(_11041_),
    .A(_09332_),
    .X(_11042_));
 sg13g2_mux2_1 _41648_ (.A0(_09331_),
    .A1(_11042_),
    .S(net5751),
    .X(_11043_));
 sg13g2_nand2_1 _41649_ (.Y(_11044_),
    .A(net5391),
    .B(_11043_));
 sg13g2_nor2_1 _41650_ (.A(net5391),
    .B(_11043_),
    .Y(_11045_));
 sg13g2_xnor2_1 _41651_ (.Y(_11046_),
    .A(net5447),
    .B(_11043_));
 sg13g2_a21oi_1 _41652_ (.A1(_11011_),
    .A2(_11032_),
    .Y(_11047_),
    .B1(net5447));
 sg13g2_nand2b_1 _41653_ (.Y(_11048_),
    .B(_11022_),
    .A_N(_11047_));
 sg13g2_o21ai_1 _41654_ (.B1(_11048_),
    .Y(_11049_),
    .A1(net5393),
    .A2(_11031_));
 sg13g2_xor2_1 _41655_ (.B(_11049_),
    .A(_11046_),
    .X(_11050_));
 sg13g2_nand2_1 _41656_ (.Y(_11051_),
    .A(net5510),
    .B(_11050_));
 sg13g2_o21ai_1 _41657_ (.B1(_11051_),
    .Y(_11052_),
    .A1(net5501),
    .A2(_11043_));
 sg13g2_nor2_1 _41658_ (.A(net5151),
    .B(_11052_),
    .Y(_11053_));
 sg13g2_a221oi_1 _41659_ (.B2(net5205),
    .C1(_11053_),
    .B1(_11031_),
    .A1(net5159),
    .Y(_11054_),
    .A2(_09343_));
 sg13g2_o21ai_1 _41660_ (.B1(_11040_),
    .Y(_00754_),
    .A1(net6845),
    .A2(_11054_));
 sg13g2_nand2_1 _41661_ (.Y(_11055_),
    .A(net5701),
    .B(_09325_));
 sg13g2_nand2_1 _41662_ (.Y(_11056_),
    .A(_09239_),
    .B(_09351_));
 sg13g2_a21o_1 _41663_ (.A2(_11056_),
    .A1(_09359_),
    .B1(_09327_),
    .X(_11057_));
 sg13g2_nand3_1 _41664_ (.B(_09359_),
    .C(_11056_),
    .A(_09327_),
    .Y(_11058_));
 sg13g2_nand3_1 _41665_ (.B(_11057_),
    .C(_11058_),
    .A(net5750),
    .Y(_11059_));
 sg13g2_nand2_2 _41666_ (.Y(_11060_),
    .A(_11055_),
    .B(_11059_));
 sg13g2_xnor2_1 _41667_ (.Y(_11061_),
    .A(net5447),
    .B(_11060_));
 sg13g2_o21ai_1 _41668_ (.B1(_11044_),
    .Y(_11062_),
    .A1(_11045_),
    .A2(_11049_));
 sg13g2_xnor2_1 _41669_ (.Y(_11063_),
    .A(_11061_),
    .B(_11062_));
 sg13g2_o21ai_1 _41670_ (.B1(net5947),
    .Y(_11064_),
    .A1(net5500),
    .A2(_11060_));
 sg13g2_a21oi_1 _41671_ (.A1(net5500),
    .A2(_11063_),
    .Y(_11065_),
    .B1(_11064_));
 sg13g2_a221oi_1 _41672_ (.B2(net5898),
    .C1(_11065_),
    .B1(_11043_),
    .A1(net5982),
    .Y(_11066_),
    .A2(_09339_));
 sg13g2_o21ai_1 _41673_ (.B1(net6878),
    .Y(_11067_),
    .A1(net5267),
    .A2(_09339_));
 sg13g2_a21oi_1 _41674_ (.A1(net5267),
    .A2(_11066_),
    .Y(_11068_),
    .B1(_11067_));
 sg13g2_a21o_1 _41675_ (.A2(net6412),
    .A1(net2381),
    .B1(_11068_),
    .X(_00755_));
 sg13g2_nand2_1 _41676_ (.Y(_11069_),
    .A(net5701),
    .B(_09318_));
 sg13g2_nand2_1 _41677_ (.Y(_11070_),
    .A(_09326_),
    .B(_11057_));
 sg13g2_xnor2_1 _41678_ (.Y(_11071_),
    .A(_09321_),
    .B(_11070_));
 sg13g2_o21ai_1 _41679_ (.B1(_11069_),
    .Y(_11072_),
    .A1(net5702),
    .A2(_11071_));
 sg13g2_nor2_1 _41680_ (.A(net5500),
    .B(_11072_),
    .Y(_11073_));
 sg13g2_nand2_1 _41681_ (.Y(_11074_),
    .A(net5391),
    .B(_11072_));
 sg13g2_xnor2_1 _41682_ (.Y(_11075_),
    .A(net5447),
    .B(_11072_));
 sg13g2_nand3_1 _41683_ (.B(_11047_),
    .C(_11061_),
    .A(_11046_),
    .Y(_11076_));
 sg13g2_o21ai_1 _41684_ (.B1(net5391),
    .Y(_11077_),
    .A1(_11043_),
    .A2(_11060_));
 sg13g2_nand2_1 _41685_ (.Y(_11078_),
    .A(_11076_),
    .B(_11077_));
 sg13g2_nand3_1 _41686_ (.B(_11046_),
    .C(_11061_),
    .A(_11013_),
    .Y(_11079_));
 sg13g2_nor2_1 _41687_ (.A(_11033_),
    .B(_11079_),
    .Y(_11080_));
 sg13g2_a21oi_1 _41688_ (.A1(_11021_),
    .A2(_11080_),
    .Y(_11081_),
    .B1(_11078_));
 sg13g2_nand2b_1 _41689_ (.Y(_11082_),
    .B(_11075_),
    .A_N(_11081_));
 sg13g2_xor2_1 _41690_ (.B(_11081_),
    .A(_11075_),
    .X(_11083_));
 sg13g2_a21oi_1 _41691_ (.A1(net5500),
    .A2(_11083_),
    .Y(_11084_),
    .B1(_11073_));
 sg13g2_a22oi_1 _41692_ (.Y(_11085_),
    .B1(_11084_),
    .B2(net5226),
    .A2(_11060_),
    .A1(net5205));
 sg13g2_a22oi_1 _41693_ (.Y(_11086_),
    .B1(net5098),
    .B2(_09331_),
    .A2(net6412),
    .A1(net3383));
 sg13g2_o21ai_1 _41694_ (.B1(_11086_),
    .Y(_00756_),
    .A1(net6845),
    .A2(_11085_));
 sg13g2_nand2_1 _41695_ (.Y(_11087_),
    .A(_11074_),
    .B(_11082_));
 sg13g2_nor2_1 _41696_ (.A(net5751),
    .B(_09312_),
    .Y(_11088_));
 sg13g2_a21oi_1 _41697_ (.A1(_09360_),
    .A2(_11057_),
    .Y(_11089_),
    .B1(_09320_));
 sg13g2_nand2_1 _41698_ (.Y(_11090_),
    .A(_09314_),
    .B(_11089_));
 sg13g2_xnor2_1 _41699_ (.Y(_11091_),
    .A(_09314_),
    .B(_11089_));
 sg13g2_a21oi_2 _41700_ (.B1(_11088_),
    .Y(_11092_),
    .A2(_11091_),
    .A1(net5751));
 sg13g2_nand2b_1 _41701_ (.Y(_11093_),
    .B(net5452),
    .A_N(_11092_));
 sg13g2_nand2_1 _41702_ (.Y(_11094_),
    .A(net5391),
    .B(_11092_));
 sg13g2_xnor2_1 _41703_ (.Y(_11095_),
    .A(net5452),
    .B(_11092_));
 sg13g2_xnor2_1 _41704_ (.Y(_11096_),
    .A(_11087_),
    .B(_11095_));
 sg13g2_o21ai_1 _41705_ (.B1(net5948),
    .Y(_11097_),
    .A1(net5500),
    .A2(_11092_));
 sg13g2_a21oi_1 _41706_ (.A1(net5500),
    .A2(_11096_),
    .Y(_11098_),
    .B1(_11097_));
 sg13g2_a221oi_1 _41707_ (.B2(net5898),
    .C1(_11098_),
    .B1(_11072_),
    .A1(net5982),
    .Y(_11099_),
    .A2(_09325_));
 sg13g2_o21ai_1 _41708_ (.B1(net6878),
    .Y(_11100_),
    .A1(net5267),
    .A2(_09325_));
 sg13g2_a21oi_1 _41709_ (.A1(net5267),
    .A2(_11099_),
    .Y(_11101_),
    .B1(_11100_));
 sg13g2_a21o_1 _41710_ (.A2(net6412),
    .A1(net3293),
    .B1(_11101_),
    .X(_00757_));
 sg13g2_nand2_1 _41711_ (.Y(_11102_),
    .A(net5701),
    .B(_09302_));
 sg13g2_nand2_1 _41712_ (.Y(_11103_),
    .A(_09313_),
    .B(_11090_));
 sg13g2_xnor2_1 _41713_ (.Y(_11104_),
    .A(_09304_),
    .B(_11103_));
 sg13g2_o21ai_1 _41714_ (.B1(_11102_),
    .Y(_11105_),
    .A1(net5701),
    .A2(_11104_));
 sg13g2_nand2_1 _41715_ (.Y(_11106_),
    .A(net5391),
    .B(_11105_));
 sg13g2_xnor2_1 _41716_ (.Y(_11107_),
    .A(net5452),
    .B(_11105_));
 sg13g2_nand2_1 _41717_ (.Y(_11108_),
    .A(_11074_),
    .B(_11094_));
 sg13g2_nand2b_1 _41718_ (.Y(_11109_),
    .B(_11082_),
    .A_N(_11108_));
 sg13g2_nand3_1 _41719_ (.B(_11107_),
    .C(_11109_),
    .A(_11093_),
    .Y(_11110_));
 sg13g2_a21o_1 _41720_ (.A2(_11109_),
    .A1(_11093_),
    .B1(_11107_),
    .X(_11111_));
 sg13g2_and2_1 _41721_ (.A(_11110_),
    .B(_11111_),
    .X(_11112_));
 sg13g2_mux2_1 _41722_ (.A0(_11105_),
    .A1(_11112_),
    .S(net5500),
    .X(_11113_));
 sg13g2_a22oi_1 _41723_ (.Y(_11114_),
    .B1(_11113_),
    .B2(net5226),
    .A2(_11092_),
    .A1(net5205));
 sg13g2_a22oi_1 _41724_ (.Y(_11115_),
    .B1(net5098),
    .B2(_09318_),
    .A2(net6413),
    .A1(net3080));
 sg13g2_o21ai_1 _41725_ (.B1(_11115_),
    .Y(_00758_),
    .A1(net6846),
    .A2(_11114_));
 sg13g2_nor2_1 _41726_ (.A(net5754),
    .B(_09267_),
    .Y(_11116_));
 sg13g2_a21oi_1 _41727_ (.A1(_09232_),
    .A2(_09238_),
    .Y(_11117_),
    .B1(_09352_));
 sg13g2_or2_1 _41728_ (.X(_11118_),
    .B(_11117_),
    .A(_09363_));
 sg13g2_nand2_1 _41729_ (.Y(_11119_),
    .A(_09269_),
    .B(_11118_));
 sg13g2_xor2_1 _41730_ (.B(_11118_),
    .A(_09269_),
    .X(_11120_));
 sg13g2_a21oi_1 _41731_ (.A1(net5751),
    .A2(_11120_),
    .Y(_11121_),
    .B1(_11116_));
 sg13g2_a21o_1 _41732_ (.A2(_11120_),
    .A1(net5751),
    .B1(_11116_),
    .X(_11122_));
 sg13g2_xnor2_1 _41733_ (.Y(_11123_),
    .A(net5391),
    .B(_11121_));
 sg13g2_nand2_1 _41734_ (.Y(_11124_),
    .A(_11106_),
    .B(_11110_));
 sg13g2_xnor2_1 _41735_ (.Y(_11125_),
    .A(_11123_),
    .B(_11124_));
 sg13g2_o21ai_1 _41736_ (.B1(net5948),
    .Y(_11126_),
    .A1(net5500),
    .A2(_11122_));
 sg13g2_a21oi_1 _41737_ (.A1(net5501),
    .A2(_11125_),
    .Y(_11127_),
    .B1(_11126_));
 sg13g2_a221oi_1 _41738_ (.B2(net5898),
    .C1(_11127_),
    .B1(_11105_),
    .A1(net5982),
    .Y(_11128_),
    .A2(_09312_));
 sg13g2_o21ai_1 _41739_ (.B1(net6878),
    .Y(_11129_),
    .A1(net5267),
    .A2(_09312_));
 sg13g2_a21oi_1 _41740_ (.A1(net5267),
    .A2(_11128_),
    .Y(_11130_),
    .B1(_11129_));
 sg13g2_a21o_1 _41741_ (.A2(net6413),
    .A1(net3210),
    .B1(_11130_),
    .X(_00759_));
 sg13g2_nand2_1 _41742_ (.Y(_11131_),
    .A(net5710),
    .B(_09261_));
 sg13g2_o21ai_1 _41743_ (.B1(_11119_),
    .Y(_11132_),
    .A1(net5586),
    .A2(_09267_));
 sg13g2_xnor2_1 _41744_ (.Y(_11133_),
    .A(_09263_),
    .B(_11132_));
 sg13g2_o21ai_1 _41745_ (.B1(_11131_),
    .Y(_11134_),
    .A1(net5710),
    .A2(_11133_));
 sg13g2_inv_1 _41746_ (.Y(_11135_),
    .A(_11134_));
 sg13g2_nor2_1 _41747_ (.A(net5511),
    .B(_11134_),
    .Y(_11136_));
 sg13g2_xnor2_1 _41748_ (.Y(_11137_),
    .A(net5404),
    .B(_11135_));
 sg13g2_and2_1 _41749_ (.A(_11107_),
    .B(_11123_),
    .X(_11138_));
 sg13g2_nand2_1 _41750_ (.Y(_11139_),
    .A(_11075_),
    .B(_11095_));
 sg13g2_a21oi_1 _41751_ (.A1(_11076_),
    .A2(_11077_),
    .Y(_11140_),
    .B1(_11139_));
 sg13g2_o21ai_1 _41752_ (.B1(_11138_),
    .Y(_11141_),
    .A1(_11108_),
    .A2(_11140_));
 sg13g2_o21ai_1 _41753_ (.B1(net5391),
    .Y(_11142_),
    .A1(_11105_),
    .A2(_11122_));
 sg13g2_nand2_2 _41754_ (.Y(_11143_),
    .A(_11141_),
    .B(_11142_));
 sg13g2_and4_1 _41755_ (.A(_11075_),
    .B(_11080_),
    .C(_11095_),
    .D(_11138_),
    .X(_11144_));
 sg13g2_a21oi_2 _41756_ (.B1(_11143_),
    .Y(_11145_),
    .A2(_11144_),
    .A1(_11021_));
 sg13g2_nand2b_1 _41757_ (.Y(_11146_),
    .B(_11137_),
    .A_N(_11145_));
 sg13g2_xor2_1 _41758_ (.B(_11145_),
    .A(_11137_),
    .X(_11147_));
 sg13g2_a21oi_1 _41759_ (.A1(net5511),
    .A2(_11147_),
    .Y(_11148_),
    .B1(_11136_));
 sg13g2_a22oi_1 _41760_ (.Y(_11149_),
    .B1(_11148_),
    .B2(net5226),
    .A2(_09302_),
    .A1(net5159));
 sg13g2_o21ai_1 _41761_ (.B1(_11149_),
    .Y(_11150_),
    .A1(net5121),
    .A2(_11121_));
 sg13g2_a22oi_1 _41762_ (.Y(_11151_),
    .B1(net6878),
    .B2(_11150_),
    .A2(net6413),
    .A1(net3142));
 sg13g2_inv_1 _41763_ (.Y(_00760_),
    .A(_11151_));
 sg13g2_nand2_1 _41764_ (.Y(_11152_),
    .A(net2537),
    .B(net6412));
 sg13g2_o21ai_1 _41765_ (.B1(_11146_),
    .Y(_11153_),
    .A1(net5453),
    .A2(_11135_));
 sg13g2_nor2_1 _41766_ (.A(net5754),
    .B(_09246_),
    .Y(_11154_));
 sg13g2_a21o_1 _41767_ (.A2(_11119_),
    .A1(_09365_),
    .B1(_09262_),
    .X(_11155_));
 sg13g2_xnor2_1 _41768_ (.Y(_11156_),
    .A(_09248_),
    .B(_11155_));
 sg13g2_a21oi_2 _41769_ (.B1(_11154_),
    .Y(_11157_),
    .A2(_11156_),
    .A1(net5754));
 sg13g2_inv_1 _41770_ (.Y(_11158_),
    .A(_11157_));
 sg13g2_xnor2_1 _41771_ (.Y(_11159_),
    .A(net5404),
    .B(_11157_));
 sg13g2_xnor2_1 _41772_ (.Y(_11160_),
    .A(_11153_),
    .B(_11159_));
 sg13g2_nand2_1 _41773_ (.Y(_11161_),
    .A(net5511),
    .B(_11160_));
 sg13g2_a21oi_1 _41774_ (.A1(net5560),
    .A2(_11157_),
    .Y(_11162_),
    .B1(net5924));
 sg13g2_a22oi_1 _41775_ (.Y(_11163_),
    .B1(_11161_),
    .B2(_11162_),
    .A2(_11134_),
    .A1(net5898));
 sg13g2_o21ai_1 _41776_ (.B1(_11163_),
    .Y(_11164_),
    .A1(net6004),
    .A2(_09267_));
 sg13g2_a21oi_2 _41777_ (.B1(_11164_),
    .Y(_11165_),
    .A2(net5316),
    .A1(net5320));
 sg13g2_o21ai_1 _41778_ (.B1(net6878),
    .Y(_11166_),
    .A1(net5267),
    .A2(_09268_));
 sg13g2_o21ai_1 _41779_ (.B1(_11152_),
    .Y(_00761_),
    .A1(_11165_),
    .A2(_11166_));
 sg13g2_o21ai_1 _41780_ (.B1(_09247_),
    .Y(_11167_),
    .A1(_09249_),
    .A2(_11155_));
 sg13g2_xnor2_1 _41781_ (.Y(_11168_),
    .A(_09257_),
    .B(_11167_));
 sg13g2_nor2_1 _41782_ (.A(net5754),
    .B(_09255_),
    .Y(_11169_));
 sg13g2_a21oi_2 _41783_ (.B1(_11169_),
    .Y(_11170_),
    .A2(_11168_),
    .A1(net5754));
 sg13g2_nor2_1 _41784_ (.A(net5511),
    .B(_11170_),
    .Y(_11171_));
 sg13g2_xnor2_1 _41785_ (.Y(_11172_),
    .A(net5404),
    .B(_11170_));
 sg13g2_o21ai_1 _41786_ (.B1(net5401),
    .Y(_11173_),
    .A1(_11134_),
    .A2(_11158_));
 sg13g2_a21oi_1 _41787_ (.A1(_11135_),
    .A2(_11157_),
    .Y(_11174_),
    .B1(net5453));
 sg13g2_a22oi_1 _41788_ (.Y(_11175_),
    .B1(_11173_),
    .B2(_11146_),
    .A2(_11157_),
    .A1(net5453));
 sg13g2_nor2b_1 _41789_ (.A(_11172_),
    .B_N(_11175_),
    .Y(_11176_));
 sg13g2_xor2_1 _41790_ (.B(_11175_),
    .A(_11172_),
    .X(_11177_));
 sg13g2_a21oi_1 _41791_ (.A1(net5511),
    .A2(_11177_),
    .Y(_11178_),
    .B1(_11171_));
 sg13g2_a22oi_1 _41792_ (.Y(_11179_),
    .B1(_11178_),
    .B2(net5226),
    .A2(_11158_),
    .A1(net5205));
 sg13g2_a22oi_1 _41793_ (.Y(_11180_),
    .B1(net5098),
    .B2(_09261_),
    .A2(net6422),
    .A1(net2948));
 sg13g2_o21ai_1 _41794_ (.B1(_11180_),
    .Y(_00762_),
    .A1(net6845),
    .A2(_11179_));
 sg13g2_nor2b_1 _41795_ (.A(net5268),
    .B_N(_09246_),
    .Y(_11181_));
 sg13g2_nand2_1 _41796_ (.Y(_11182_),
    .A(net5710),
    .B(_09295_));
 sg13g2_a21oi_1 _41797_ (.A1(_09270_),
    .A2(_11118_),
    .Y(_11183_),
    .B1(_09368_));
 sg13g2_xnor2_1 _41798_ (.Y(_11184_),
    .A(_09297_),
    .B(_11183_));
 sg13g2_o21ai_1 _41799_ (.B1(_11182_),
    .Y(_11185_),
    .A1(net5710),
    .A2(_11184_));
 sg13g2_xnor2_1 _41800_ (.Y(_11186_),
    .A(net5453),
    .B(_11185_));
 sg13g2_a21o_1 _41801_ (.A2(_11170_),
    .A1(net5401),
    .B1(_11176_),
    .X(_11187_));
 sg13g2_xnor2_1 _41802_ (.Y(_11188_),
    .A(_11186_),
    .B(_11187_));
 sg13g2_o21ai_1 _41803_ (.B1(net5950),
    .Y(_11189_),
    .A1(net5511),
    .A2(_11185_));
 sg13g2_a21oi_1 _41804_ (.A1(net5511),
    .A2(_11188_),
    .Y(_11190_),
    .B1(_11189_));
 sg13g2_a21oi_1 _41805_ (.A1(net5898),
    .A2(_11170_),
    .Y(_11191_),
    .B1(_11190_));
 sg13g2_o21ai_1 _41806_ (.B1(_11191_),
    .Y(_11192_),
    .A1(net6005),
    .A2(_09246_));
 sg13g2_nor2b_1 _41807_ (.A(_11192_),
    .B_N(net5269),
    .Y(_11193_));
 sg13g2_nor3_1 _41808_ (.A(net6845),
    .B(_11181_),
    .C(_11193_),
    .Y(_11194_));
 sg13g2_a21o_1 _41809_ (.A2(net6412),
    .A1(net3133),
    .B1(_11194_),
    .X(_00763_));
 sg13g2_o21ai_1 _41810_ (.B1(_09296_),
    .Y(_11195_),
    .A1(_09297_),
    .A2(_11183_));
 sg13g2_o21ai_1 _41811_ (.B1(_11195_),
    .Y(_11196_),
    .A1(net5645),
    .A2(_09289_));
 sg13g2_xnor2_1 _41812_ (.Y(_11197_),
    .A(_09291_),
    .B(_11195_));
 sg13g2_nand2_1 _41813_ (.Y(_11198_),
    .A(net5754),
    .B(_11197_));
 sg13g2_o21ai_1 _41814_ (.B1(_11198_),
    .Y(_11199_),
    .A1(net5754),
    .A2(_09288_));
 sg13g2_nand2_1 _41815_ (.Y(_11200_),
    .A(net5401),
    .B(_11199_));
 sg13g2_xnor2_1 _41816_ (.Y(_11201_),
    .A(net5453),
    .B(_11199_));
 sg13g2_nor2b_1 _41817_ (.A(_11172_),
    .B_N(_11186_),
    .Y(_11202_));
 sg13g2_nand3b_1 _41818_ (.B(_11174_),
    .C(_11186_),
    .Y(_11203_),
    .A_N(_11172_));
 sg13g2_o21ai_1 _41819_ (.B1(net5401),
    .Y(_11204_),
    .A1(_11170_),
    .A2(_11185_));
 sg13g2_nand2_1 _41820_ (.Y(_11205_),
    .A(_11203_),
    .B(_11204_));
 sg13g2_nand3_1 _41821_ (.B(_11159_),
    .C(_11202_),
    .A(_11137_),
    .Y(_11206_));
 sg13g2_nor2_1 _41822_ (.A(_11145_),
    .B(_11206_),
    .Y(_11207_));
 sg13g2_o21ai_1 _41823_ (.B1(_11201_),
    .Y(_11208_),
    .A1(_11205_),
    .A2(_11207_));
 sg13g2_or3_1 _41824_ (.A(_11201_),
    .B(_11205_),
    .C(_11207_),
    .X(_11209_));
 sg13g2_nand2_1 _41825_ (.Y(_11210_),
    .A(_11208_),
    .B(_11209_));
 sg13g2_o21ai_1 _41826_ (.B1(net5952),
    .Y(_11211_),
    .A1(net5512),
    .A2(_11199_));
 sg13g2_a21oi_1 _41827_ (.A1(net5512),
    .A2(_11210_),
    .Y(_11212_),
    .B1(_11211_));
 sg13g2_a221oi_1 _41828_ (.B2(net5898),
    .C1(_11212_),
    .B1(_11185_),
    .A1(net5982),
    .Y(_11213_),
    .A2(_09255_));
 sg13g2_a21oi_1 _41829_ (.A1(net5269),
    .A2(_11213_),
    .Y(_11214_),
    .B1(net6846));
 sg13g2_o21ai_1 _41830_ (.B1(_11214_),
    .Y(_11215_),
    .A1(net5268),
    .A2(_09255_));
 sg13g2_o21ai_1 _41831_ (.B1(_11215_),
    .Y(_00764_),
    .A1(_18177_),
    .A2(net6492));
 sg13g2_nand2_1 _41832_ (.Y(_11216_),
    .A(_09290_),
    .B(_11196_));
 sg13g2_xnor2_1 _41833_ (.Y(_11217_),
    .A(_09284_),
    .B(_11216_));
 sg13g2_nand2b_1 _41834_ (.Y(_11218_),
    .B(net5710),
    .A_N(_09280_));
 sg13g2_o21ai_1 _41835_ (.B1(_11218_),
    .Y(_11219_),
    .A1(net5710),
    .A2(_11217_));
 sg13g2_nand2_1 _41836_ (.Y(_11220_),
    .A(net5401),
    .B(_11219_));
 sg13g2_xnor2_1 _41837_ (.Y(_11221_),
    .A(net5453),
    .B(_11219_));
 sg13g2_nand2_1 _41838_ (.Y(_11222_),
    .A(_11200_),
    .B(_11208_));
 sg13g2_xnor2_1 _41839_ (.Y(_11223_),
    .A(_11221_),
    .B(_11222_));
 sg13g2_o21ai_1 _41840_ (.B1(net5952),
    .Y(_11224_),
    .A1(net5512),
    .A2(_11219_));
 sg13g2_a21oi_1 _41841_ (.A1(net5512),
    .A2(_11223_),
    .Y(_11225_),
    .B1(_11224_));
 sg13g2_a221oi_1 _41842_ (.B2(net5902),
    .C1(_11225_),
    .B1(_11199_),
    .A1(net5989),
    .Y(_11226_),
    .A2(_09295_));
 sg13g2_a21oi_1 _41843_ (.A1(net5269),
    .A2(_11226_),
    .Y(_11227_),
    .B1(net6850));
 sg13g2_o21ai_1 _41844_ (.B1(_11227_),
    .Y(_11228_),
    .A1(net5268),
    .A2(_09295_));
 sg13g2_o21ai_1 _41845_ (.B1(_11228_),
    .Y(_00765_),
    .A1(_18176_),
    .A2(net6492));
 sg13g2_a21oi_1 _41846_ (.A1(_09284_),
    .A2(_11216_),
    .Y(_11229_),
    .B1(_09282_));
 sg13g2_xor2_1 _41847_ (.B(_11229_),
    .A(_09275_),
    .X(_11230_));
 sg13g2_or2_1 _41848_ (.X(_11231_),
    .B(_09273_),
    .A(net5754));
 sg13g2_o21ai_1 _41849_ (.B1(_11231_),
    .Y(_11232_),
    .A1(net5710),
    .A2(_11230_));
 sg13g2_nand2b_1 _41850_ (.Y(_11233_),
    .B(net5401),
    .A_N(_11232_));
 sg13g2_inv_1 _41851_ (.Y(_11234_),
    .A(_11233_));
 sg13g2_xnor2_1 _41852_ (.Y(_11235_),
    .A(net5453),
    .B(_11232_));
 sg13g2_nand2_1 _41853_ (.Y(_11236_),
    .A(_11200_),
    .B(_11220_));
 sg13g2_nand2b_1 _41854_ (.Y(_11237_),
    .B(_11208_),
    .A_N(_11236_));
 sg13g2_o21ai_1 _41855_ (.B1(_11237_),
    .Y(_11238_),
    .A1(net5401),
    .A2(_11219_));
 sg13g2_xor2_1 _41856_ (.B(_11238_),
    .A(_11235_),
    .X(_11239_));
 sg13g2_a21oi_1 _41857_ (.A1(net5560),
    .A2(_11232_),
    .Y(_11240_),
    .B1(net5926));
 sg13g2_o21ai_1 _41858_ (.B1(_11240_),
    .Y(_11241_),
    .A1(net5560),
    .A2(_11239_));
 sg13g2_a22oi_1 _41859_ (.Y(_11242_),
    .B1(_11219_),
    .B2(net5902),
    .A2(_09289_),
    .A1(net5989));
 sg13g2_nand3_1 _41860_ (.B(_11241_),
    .C(_11242_),
    .A(net5268),
    .Y(_11243_));
 sg13g2_nor2_1 _41861_ (.A(net5269),
    .B(_09289_),
    .Y(_11244_));
 sg13g2_nor2_1 _41862_ (.A(net6850),
    .B(_11244_),
    .Y(_11245_));
 sg13g2_a22oi_1 _41863_ (.Y(_11246_),
    .B1(_11243_),
    .B2(_11245_),
    .A2(net6422),
    .A1(net1915));
 sg13g2_inv_1 _41864_ (.Y(_00766_),
    .A(_11246_));
 sg13g2_or2_1 _41865_ (.X(_11247_),
    .B(_09603_),
    .A(_09373_));
 sg13g2_a21oi_1 _41866_ (.A1(_09373_),
    .A2(_09603_),
    .Y(_11248_),
    .B1(net5709));
 sg13g2_nand2_1 _41867_ (.Y(_11249_),
    .A(_11247_),
    .B(_11248_));
 sg13g2_o21ai_1 _41868_ (.B1(_11249_),
    .Y(_11250_),
    .A1(net5757),
    .A2(_09601_));
 sg13g2_xnor2_1 _41869_ (.Y(_11251_),
    .A(net5453),
    .B(_11250_));
 sg13g2_o21ai_1 _41870_ (.B1(_11233_),
    .Y(_11252_),
    .A1(_11235_),
    .A2(_11238_));
 sg13g2_xnor2_1 _41871_ (.Y(_11253_),
    .A(_11251_),
    .B(_11252_));
 sg13g2_o21ai_1 _41872_ (.B1(net5952),
    .Y(_11254_),
    .A1(net5511),
    .A2(_11250_));
 sg13g2_a21oi_1 _41873_ (.A1(net5512),
    .A2(_11253_),
    .Y(_11255_),
    .B1(_11254_));
 sg13g2_nor2_1 _41874_ (.A(net6008),
    .B(_09280_),
    .Y(_11256_));
 sg13g2_nor2_1 _41875_ (.A(net5882),
    .B(_11232_),
    .Y(_11257_));
 sg13g2_nor3_1 _41876_ (.A(_11255_),
    .B(_11256_),
    .C(_11257_),
    .Y(_11258_));
 sg13g2_nand3_1 _41877_ (.B(net5317),
    .C(_09280_),
    .A(net5321),
    .Y(_11259_));
 sg13g2_a21oi_1 _41878_ (.A1(net5268),
    .A2(_11258_),
    .Y(_11260_),
    .B1(net6850));
 sg13g2_a22oi_1 _41879_ (.Y(_11261_),
    .B1(_11259_),
    .B2(_11260_),
    .A2(net6422),
    .A1(net3471));
 sg13g2_inv_1 _41880_ (.Y(_00767_),
    .A(_11261_));
 sg13g2_nand2b_1 _41881_ (.Y(_11262_),
    .B(_11251_),
    .A_N(_11235_));
 sg13g2_nand2_1 _41882_ (.Y(_11263_),
    .A(_11201_),
    .B(_11221_));
 sg13g2_nor3_1 _41883_ (.A(_11206_),
    .B(_11262_),
    .C(_11263_),
    .Y(_11264_));
 sg13g2_a21oi_1 _41884_ (.A1(_11203_),
    .A2(_11204_),
    .Y(_11265_),
    .B1(_11263_));
 sg13g2_nor2_1 _41885_ (.A(_11236_),
    .B(_11265_),
    .Y(_11266_));
 sg13g2_a21oi_1 _41886_ (.A1(net5401),
    .A2(_11250_),
    .Y(_11267_),
    .B1(_11234_));
 sg13g2_o21ai_1 _41887_ (.B1(_11267_),
    .Y(_11268_),
    .A1(_11262_),
    .A2(_11266_));
 sg13g2_nor3_1 _41888_ (.A(_11206_),
    .B(_11262_),
    .C(_11263_),
    .Y(_11269_));
 sg13g2_a21o_2 _41889_ (.A2(_11264_),
    .A1(_11143_),
    .B1(_11268_),
    .X(_11270_));
 sg13g2_nand2_1 _41890_ (.Y(_11271_),
    .A(_11144_),
    .B(_11269_));
 sg13g2_a21oi_2 _41891_ (.B1(_11271_),
    .Y(_11272_),
    .A2(_11020_),
    .A1(_11017_));
 sg13g2_or2_1 _41892_ (.X(_11273_),
    .B(_11272_),
    .A(_11270_));
 sg13g2_nand2_1 _41893_ (.Y(_11274_),
    .A(net5709),
    .B(_09607_));
 sg13g2_o21ai_1 _41894_ (.B1(_11247_),
    .Y(_11275_),
    .A1(net5646),
    .A2(_09601_));
 sg13g2_xor2_1 _41895_ (.B(_11275_),
    .A(_09609_),
    .X(_11276_));
 sg13g2_o21ai_1 _41896_ (.B1(_11274_),
    .Y(_11277_),
    .A1(net5709),
    .A2(_11276_));
 sg13g2_inv_1 _41897_ (.Y(_11278_),
    .A(_11277_));
 sg13g2_nand2_1 _41898_ (.Y(_11279_),
    .A(net5454),
    .B(_11278_));
 sg13g2_xnor2_1 _41899_ (.Y(_11280_),
    .A(net5402),
    .B(_11278_));
 sg13g2_nand2b_1 _41900_ (.Y(_11281_),
    .B(_11273_),
    .A_N(_11280_));
 sg13g2_xor2_1 _41901_ (.B(_11280_),
    .A(_11273_),
    .X(_11282_));
 sg13g2_o21ai_1 _41902_ (.B1(net5952),
    .Y(_11283_),
    .A1(net5513),
    .A2(_11277_));
 sg13g2_a21oi_1 _41903_ (.A1(net5513),
    .A2(_11282_),
    .Y(_11284_),
    .B1(_11283_));
 sg13g2_a221oi_1 _41904_ (.B2(net5902),
    .C1(_11284_),
    .B1(_11250_),
    .A1(net5989),
    .Y(_11285_),
    .A2(_09273_));
 sg13g2_a21oi_1 _41905_ (.A1(net5268),
    .A2(_11285_),
    .Y(_11286_),
    .B1(net6850));
 sg13g2_o21ai_1 _41906_ (.B1(_11286_),
    .Y(_11287_),
    .A1(net5268),
    .A2(_09273_));
 sg13g2_o21ai_1 _41907_ (.B1(_11287_),
    .Y(_00768_),
    .A1(_18174_),
    .A2(net6491));
 sg13g2_o21ai_1 _41908_ (.B1(_11281_),
    .Y(_11288_),
    .A1(net5402),
    .A2(_11278_));
 sg13g2_nand2_1 _41909_ (.Y(_11289_),
    .A(net5709),
    .B(_09591_));
 sg13g2_and2_1 _41910_ (.A(_09615_),
    .B(_11247_),
    .X(_11290_));
 sg13g2_nor2_1 _41911_ (.A(_09608_),
    .B(_11290_),
    .Y(_11291_));
 sg13g2_nor3_1 _41912_ (.A(_09592_),
    .B(_09608_),
    .C(_11290_),
    .Y(_11292_));
 sg13g2_xor2_1 _41913_ (.B(_11291_),
    .A(_09592_),
    .X(_11293_));
 sg13g2_o21ai_1 _41914_ (.B1(_11289_),
    .Y(_11294_),
    .A1(net5709),
    .A2(_11293_));
 sg13g2_xnor2_1 _41915_ (.Y(_11295_),
    .A(net5454),
    .B(_11294_));
 sg13g2_xnor2_1 _41916_ (.Y(_11296_),
    .A(_11288_),
    .B(_11295_));
 sg13g2_o21ai_1 _41917_ (.B1(net5952),
    .Y(_11297_),
    .A1(net5513),
    .A2(_11294_));
 sg13g2_a21oi_1 _41918_ (.A1(net5513),
    .A2(_11296_),
    .Y(_11298_),
    .B1(_11297_));
 sg13g2_a221oi_1 _41919_ (.B2(net5902),
    .C1(_11298_),
    .B1(_11277_),
    .A1(net5989),
    .Y(_11299_),
    .A2(_09602_));
 sg13g2_o21ai_1 _41920_ (.B1(net6880),
    .Y(_11300_),
    .A1(net5277),
    .A2(_09602_));
 sg13g2_a21oi_1 _41921_ (.A1(net5278),
    .A2(_11299_),
    .Y(_11301_),
    .B1(_11300_));
 sg13g2_a21o_1 _41922_ (.A2(net6426),
    .A1(net2100),
    .B1(_11301_),
    .X(_00769_));
 sg13g2_nand2_1 _41923_ (.Y(_11302_),
    .A(net5709),
    .B(_09595_));
 sg13g2_a21oi_1 _41924_ (.A1(net5646),
    .A2(_09591_),
    .Y(_11303_),
    .B1(_11292_));
 sg13g2_xnor2_1 _41925_ (.Y(_11304_),
    .A(_09597_),
    .B(_11303_));
 sg13g2_o21ai_1 _41926_ (.B1(_11302_),
    .Y(_11305_),
    .A1(net5709),
    .A2(_11304_));
 sg13g2_nor2_1 _41927_ (.A(net5513),
    .B(_11305_),
    .Y(_11306_));
 sg13g2_nand2_1 _41928_ (.Y(_11307_),
    .A(net5402),
    .B(_11305_));
 sg13g2_xnor2_1 _41929_ (.Y(_11308_),
    .A(net5454),
    .B(_11305_));
 sg13g2_nor2b_1 _41930_ (.A(_11281_),
    .B_N(_11295_),
    .Y(_11309_));
 sg13g2_a21o_1 _41931_ (.A2(_11294_),
    .A1(_11279_),
    .B1(_11309_),
    .X(_11310_));
 sg13g2_nand2_1 _41932_ (.Y(_11311_),
    .A(_11308_),
    .B(_11310_));
 sg13g2_xnor2_1 _41933_ (.Y(_11312_),
    .A(_11308_),
    .B(_11310_));
 sg13g2_a21oi_1 _41934_ (.A1(net5513),
    .A2(_11312_),
    .Y(_11313_),
    .B1(_11306_));
 sg13g2_a22oi_1 _41935_ (.Y(_11314_),
    .B1(_11313_),
    .B2(net5228),
    .A2(_11294_),
    .A1(net5209));
 sg13g2_a22oi_1 _41936_ (.Y(_11315_),
    .B1(net5101),
    .B2(_09607_),
    .A2(net6426),
    .A1(net3096));
 sg13g2_o21ai_1 _41937_ (.B1(_11315_),
    .Y(_00770_),
    .A1(net6850),
    .A2(_11314_));
 sg13g2_o21ai_1 _41938_ (.B1(_09610_),
    .Y(_11316_),
    .A1(_09354_),
    .A2(_09372_));
 sg13g2_nand2_1 _41939_ (.Y(_11317_),
    .A(_09618_),
    .B(_11316_));
 sg13g2_nand2_1 _41940_ (.Y(_11318_),
    .A(_09585_),
    .B(_11317_));
 sg13g2_nor2_1 _41941_ (.A(_09585_),
    .B(_11317_),
    .Y(_11319_));
 sg13g2_nor2_1 _41942_ (.A(net5709),
    .B(_11319_),
    .Y(_11320_));
 sg13g2_a22oi_1 _41943_ (.Y(_11321_),
    .B1(_11318_),
    .B2(_11320_),
    .A2(_09583_),
    .A1(net5713));
 sg13g2_inv_1 _41944_ (.Y(_11322_),
    .A(_11321_));
 sg13g2_xnor2_1 _41945_ (.Y(_11323_),
    .A(net5402),
    .B(_11321_));
 sg13g2_nand2_1 _41946_ (.Y(_11324_),
    .A(_11307_),
    .B(_11311_));
 sg13g2_xor2_1 _41947_ (.B(_11324_),
    .A(_11323_),
    .X(_11325_));
 sg13g2_a21oi_1 _41948_ (.A1(net5559),
    .A2(_11321_),
    .Y(_11326_),
    .B1(net5926));
 sg13g2_o21ai_1 _41949_ (.B1(_11326_),
    .Y(_11327_),
    .A1(net5559),
    .A2(_11325_));
 sg13g2_a22oi_1 _41950_ (.Y(_11328_),
    .B1(_11305_),
    .B2(net5902),
    .A2(_09591_),
    .A1(net5989));
 sg13g2_nand3_1 _41951_ (.B(_11327_),
    .C(_11328_),
    .A(net5277),
    .Y(_11329_));
 sg13g2_o21ai_1 _41952_ (.B1(net6880),
    .Y(_11330_),
    .A1(net5277),
    .A2(_09591_));
 sg13g2_nand2b_1 _41953_ (.Y(_11331_),
    .B(_11329_),
    .A_N(_11330_));
 sg13g2_o21ai_1 _41954_ (.B1(_11331_),
    .Y(_00771_),
    .A1(_18172_),
    .A2(net6493));
 sg13g2_nand2_1 _41955_ (.Y(_11332_),
    .A(_09584_),
    .B(_11318_));
 sg13g2_a21o_1 _41956_ (.A2(_11318_),
    .A1(_09584_),
    .B1(_09577_),
    .X(_11333_));
 sg13g2_xor2_1 _41957_ (.B(_11332_),
    .A(_09578_),
    .X(_11334_));
 sg13g2_nand2_1 _41958_ (.Y(_11335_),
    .A(net5757),
    .B(_11334_));
 sg13g2_o21ai_1 _41959_ (.B1(_11335_),
    .Y(_11336_),
    .A1(net5757),
    .A2(_09574_));
 sg13g2_nor2_1 _41960_ (.A(net5514),
    .B(_11336_),
    .Y(_11337_));
 sg13g2_xnor2_1 _41961_ (.Y(_11338_),
    .A(net5402),
    .B(_11336_));
 sg13g2_and2_1 _41962_ (.A(_11308_),
    .B(_11323_),
    .X(_11339_));
 sg13g2_and4_1 _41963_ (.A(_11279_),
    .B(_11294_),
    .C(_11308_),
    .D(_11323_),
    .X(_11340_));
 sg13g2_o21ai_1 _41964_ (.B1(_11307_),
    .Y(_11341_),
    .A1(net5454),
    .A2(_11321_));
 sg13g2_or2_1 _41965_ (.X(_11342_),
    .B(_11341_),
    .A(_11340_));
 sg13g2_a21oi_1 _41966_ (.A1(_11309_),
    .A2(_11339_),
    .Y(_11343_),
    .B1(_11342_));
 sg13g2_nor2_1 _41967_ (.A(_11338_),
    .B(_11343_),
    .Y(_11344_));
 sg13g2_xnor2_1 _41968_ (.Y(_11345_),
    .A(_11338_),
    .B(_11343_));
 sg13g2_a21oi_1 _41969_ (.A1(net5514),
    .A2(_11345_),
    .Y(_11346_),
    .B1(_11337_));
 sg13g2_a22oi_1 _41970_ (.Y(_11347_),
    .B1(_11346_),
    .B2(net5228),
    .A2(_11322_),
    .A1(net5209));
 sg13g2_a22oi_1 _41971_ (.Y(_11348_),
    .B1(net5101),
    .B2(_09595_),
    .A2(net6426),
    .A1(net2646));
 sg13g2_o21ai_1 _41972_ (.B1(_11348_),
    .Y(_00772_),
    .A1(net6858),
    .A2(_11347_));
 sg13g2_nor2_1 _41973_ (.A(net5758),
    .B(_09568_),
    .Y(_11349_));
 sg13g2_a21o_1 _41974_ (.A2(_11333_),
    .A1(_09576_),
    .B1(_09571_),
    .X(_11350_));
 sg13g2_nand3_1 _41975_ (.B(_09576_),
    .C(_11333_),
    .A(_09571_),
    .Y(_11351_));
 sg13g2_a21oi_1 _41976_ (.A1(_11350_),
    .A2(_11351_),
    .Y(_11352_),
    .B1(net5716));
 sg13g2_nor2_2 _41977_ (.A(_11349_),
    .B(_11352_),
    .Y(_11353_));
 sg13g2_xnor2_1 _41978_ (.Y(_11354_),
    .A(net5403),
    .B(_11353_));
 sg13g2_a21oi_1 _41979_ (.A1(net5403),
    .A2(_11336_),
    .Y(_11355_),
    .B1(_11344_));
 sg13g2_xnor2_1 _41980_ (.Y(_11356_),
    .A(_11354_),
    .B(_11355_));
 sg13g2_o21ai_1 _41981_ (.B1(net5953),
    .Y(_11357_),
    .A1(net5514),
    .A2(_11353_));
 sg13g2_a21oi_1 _41982_ (.A1(net5514),
    .A2(_11356_),
    .Y(_11358_),
    .B1(_11357_));
 sg13g2_a221oi_1 _41983_ (.B2(net5903),
    .C1(_11358_),
    .B1(_11336_),
    .A1(net5986),
    .Y(_11359_),
    .A2(_09583_));
 sg13g2_a21oi_1 _41984_ (.A1(net5277),
    .A2(_11359_),
    .Y(_11360_),
    .B1(net6851));
 sg13g2_o21ai_1 _41985_ (.B1(_11360_),
    .Y(_11361_),
    .A1(net5277),
    .A2(_09583_));
 sg13g2_o21ai_1 _41986_ (.B1(_11361_),
    .Y(_00773_),
    .A1(_18171_),
    .A2(net6499));
 sg13g2_nor2_1 _41987_ (.A(net5758),
    .B(_09558_),
    .Y(_11362_));
 sg13g2_nand2_1 _41988_ (.Y(_11363_),
    .A(_09569_),
    .B(_11350_));
 sg13g2_xnor2_1 _41989_ (.Y(_11364_),
    .A(_09559_),
    .B(_11363_));
 sg13g2_a21oi_2 _41990_ (.B1(_11362_),
    .Y(_11365_),
    .A2(_11364_),
    .A1(net5758));
 sg13g2_nand2_1 _41991_ (.Y(_11366_),
    .A(net5402),
    .B(_11365_));
 sg13g2_xnor2_1 _41992_ (.Y(_11367_),
    .A(net5402),
    .B(_11365_));
 sg13g2_o21ai_1 _41993_ (.B1(net5402),
    .Y(_11368_),
    .A1(_11336_),
    .A2(_11353_));
 sg13g2_o21ai_1 _41994_ (.B1(_11368_),
    .Y(_11369_),
    .A1(_11338_),
    .A2(_11343_));
 sg13g2_o21ai_1 _41995_ (.B1(_11369_),
    .Y(_11370_),
    .A1(net5403),
    .A2(_11353_));
 sg13g2_xnor2_1 _41996_ (.Y(_11371_),
    .A(_11367_),
    .B(_11370_));
 sg13g2_a21oi_1 _41997_ (.A1(net5513),
    .A2(_11371_),
    .Y(_11372_),
    .B1(net5929));
 sg13g2_o21ai_1 _41998_ (.B1(_11372_),
    .Y(_11373_),
    .A1(net5513),
    .A2(_11365_));
 sg13g2_a22oi_1 _41999_ (.Y(_11374_),
    .B1(_11353_),
    .B2(net5903),
    .A2(_09575_),
    .A1(net5986));
 sg13g2_nand3_1 _42000_ (.B(_11373_),
    .C(_11374_),
    .A(net5277),
    .Y(_11375_));
 sg13g2_nor2_1 _42001_ (.A(net5277),
    .B(_09575_),
    .Y(_11376_));
 sg13g2_nor2_1 _42002_ (.A(net6851),
    .B(_11376_),
    .Y(_11377_));
 sg13g2_a22oi_1 _42003_ (.Y(_11378_),
    .B1(_11375_),
    .B2(_11377_),
    .A2(net6429),
    .A1(net2764));
 sg13g2_inv_1 _42004_ (.Y(_00774_),
    .A(_11378_));
 sg13g2_nand2_1 _42005_ (.Y(_11379_),
    .A(net5716),
    .B(_09522_));
 sg13g2_o21ai_1 _42006_ (.B1(_09611_),
    .Y(_11380_),
    .A1(_09354_),
    .A2(_09372_));
 sg13g2_nand2_1 _42007_ (.Y(_11381_),
    .A(_09624_),
    .B(_11380_));
 sg13g2_xnor2_1 _42008_ (.Y(_11382_),
    .A(_09524_),
    .B(_11381_));
 sg13g2_o21ai_1 _42009_ (.B1(_11379_),
    .Y(_11383_),
    .A1(net5716),
    .A2(_11382_));
 sg13g2_nand2_1 _42010_ (.Y(_11384_),
    .A(net5403),
    .B(_11383_));
 sg13g2_xnor2_1 _42011_ (.Y(_11385_),
    .A(net5454),
    .B(_11383_));
 sg13g2_o21ai_1 _42012_ (.B1(_11366_),
    .Y(_11386_),
    .A1(_11367_),
    .A2(_11370_));
 sg13g2_xnor2_1 _42013_ (.Y(_11387_),
    .A(_11385_),
    .B(_11386_));
 sg13g2_o21ai_1 _42014_ (.B1(net5954),
    .Y(_11388_),
    .A1(net5514),
    .A2(_11383_));
 sg13g2_a21oi_1 _42015_ (.A1(net5514),
    .A2(_11387_),
    .Y(_11389_),
    .B1(_11388_));
 sg13g2_a221oi_1 _42016_ (.B2(net5903),
    .C1(_11389_),
    .B1(_11365_),
    .A1(net5986),
    .Y(_11390_),
    .A2(_09568_));
 sg13g2_a21oi_1 _42017_ (.A1(net5278),
    .A2(_11390_),
    .Y(_11391_),
    .B1(net6851));
 sg13g2_o21ai_1 _42018_ (.B1(_11391_),
    .Y(_11392_),
    .A1(net5278),
    .A2(_09568_));
 sg13g2_o21ai_1 _42019_ (.B1(_11392_),
    .Y(_00775_),
    .A1(_18170_),
    .A2(net6493));
 sg13g2_a21oi_1 _42020_ (.A1(_09524_),
    .A2(_11381_),
    .Y(_11393_),
    .B1(_09523_));
 sg13g2_xor2_1 _42021_ (.B(_11393_),
    .A(_09518_),
    .X(_11394_));
 sg13g2_nand2_1 _42022_ (.Y(_11395_),
    .A(net5716),
    .B(_09515_));
 sg13g2_o21ai_1 _42023_ (.B1(_11395_),
    .Y(_11396_),
    .A1(net5716),
    .A2(_11394_));
 sg13g2_nor2_1 _42024_ (.A(net5520),
    .B(_11396_),
    .Y(_11397_));
 sg13g2_nand2_1 _42025_ (.Y(_11398_),
    .A(net5413),
    .B(_11396_));
 sg13g2_xnor2_1 _42026_ (.Y(_11399_),
    .A(net5457),
    .B(_11396_));
 sg13g2_nand2b_1 _42027_ (.Y(_11400_),
    .B(_11385_),
    .A_N(_11367_));
 sg13g2_nor2_1 _42028_ (.A(_11338_),
    .B(_11354_),
    .Y(_11401_));
 sg13g2_o21ai_1 _42029_ (.B1(_11401_),
    .Y(_11402_),
    .A1(_11340_),
    .A2(_11341_));
 sg13g2_a21oi_1 _42030_ (.A1(_11368_),
    .A2(_11402_),
    .Y(_11403_),
    .B1(_11400_));
 sg13g2_nand2_1 _42031_ (.Y(_11404_),
    .A(_11366_),
    .B(_11384_));
 sg13g2_nand3b_1 _42032_ (.B(_11295_),
    .C(_11339_),
    .Y(_11405_),
    .A_N(_11280_));
 sg13g2_nor4_1 _42033_ (.A(_11338_),
    .B(_11354_),
    .C(_11400_),
    .D(_11405_),
    .Y(_11406_));
 sg13g2_and2_1 _42034_ (.A(_11273_),
    .B(_11406_),
    .X(_11407_));
 sg13g2_nor3_1 _42035_ (.A(_11403_),
    .B(_11404_),
    .C(_11407_),
    .Y(_11408_));
 sg13g2_nand2b_1 _42036_ (.Y(_11409_),
    .B(_11399_),
    .A_N(_11408_));
 sg13g2_xor2_1 _42037_ (.B(_11408_),
    .A(_11399_),
    .X(_11410_));
 sg13g2_a21oi_1 _42038_ (.A1(net5520),
    .A2(_11410_),
    .Y(_11411_),
    .B1(_11397_));
 sg13g2_a22oi_1 _42039_ (.Y(_11412_),
    .B1(_11411_),
    .B2(net5229),
    .A2(_11383_),
    .A1(net5210));
 sg13g2_a22oi_1 _42040_ (.Y(_11413_),
    .B1(net5102),
    .B2(_09558_),
    .A2(net6429),
    .A1(net3163));
 sg13g2_o21ai_1 _42041_ (.B1(_11413_),
    .Y(_00776_),
    .A1(net6851),
    .A2(_11412_));
 sg13g2_nand2_1 _42042_ (.Y(_11414_),
    .A(_11398_),
    .B(_11409_));
 sg13g2_nor2_1 _42043_ (.A(net5758),
    .B(_09501_),
    .Y(_11415_));
 sg13g2_o21ai_1 _42044_ (.B1(_09517_),
    .Y(_11416_),
    .A1(_09516_),
    .A2(_11393_));
 sg13g2_xnor2_1 _42045_ (.Y(_11417_),
    .A(_09504_),
    .B(_11416_));
 sg13g2_a21oi_2 _42046_ (.B1(_11415_),
    .Y(_11418_),
    .A2(_11417_),
    .A1(net5758));
 sg13g2_nand2b_1 _42047_ (.Y(_11419_),
    .B(net5457),
    .A_N(_11418_));
 sg13g2_xnor2_1 _42048_ (.Y(_11420_),
    .A(net5413),
    .B(_11418_));
 sg13g2_xor2_1 _42049_ (.B(_11420_),
    .A(_11414_),
    .X(_11421_));
 sg13g2_o21ai_1 _42050_ (.B1(net5954),
    .Y(_11422_),
    .A1(net5520),
    .A2(_11418_));
 sg13g2_a21oi_1 _42051_ (.A1(net5520),
    .A2(_11421_),
    .Y(_11423_),
    .B1(_11422_));
 sg13g2_a221oi_1 _42052_ (.B2(net5903),
    .C1(_11423_),
    .B1(_11396_),
    .A1(net5986),
    .Y(_11424_),
    .A2(_09522_));
 sg13g2_o21ai_1 _42053_ (.B1(net6880),
    .Y(_11425_),
    .A1(net5279),
    .A2(_09522_));
 sg13g2_a21oi_1 _42054_ (.A1(net5279),
    .A2(_11424_),
    .Y(_11426_),
    .B1(_11425_));
 sg13g2_a21o_1 _42055_ (.A2(net6429),
    .A1(net3323),
    .B1(_11426_),
    .X(_00777_));
 sg13g2_nand2_1 _42056_ (.Y(_11427_),
    .A(net5716),
    .B(_09510_));
 sg13g2_a21oi_1 _42057_ (.A1(_09504_),
    .A2(_11416_),
    .Y(_11428_),
    .B1(_09503_));
 sg13g2_xor2_1 _42058_ (.B(_11428_),
    .A(_09511_),
    .X(_11429_));
 sg13g2_o21ai_1 _42059_ (.B1(_11427_),
    .Y(_11430_),
    .A1(net5716),
    .A2(_11429_));
 sg13g2_nor2_1 _42060_ (.A(net5520),
    .B(_11430_),
    .Y(_11431_));
 sg13g2_nand2_1 _42061_ (.Y(_11432_),
    .A(net5413),
    .B(_11430_));
 sg13g2_xnor2_1 _42062_ (.Y(_11433_),
    .A(net5457),
    .B(_11430_));
 sg13g2_o21ai_1 _42063_ (.B1(net5413),
    .Y(_11434_),
    .A1(_11396_),
    .A2(_11418_));
 sg13g2_nand2_1 _42064_ (.Y(_11435_),
    .A(_11409_),
    .B(_11434_));
 sg13g2_nand3_1 _42065_ (.B(_11433_),
    .C(_11435_),
    .A(_11419_),
    .Y(_11436_));
 sg13g2_a21o_1 _42066_ (.A2(_11435_),
    .A1(_11419_),
    .B1(_11433_),
    .X(_11437_));
 sg13g2_nand2_1 _42067_ (.Y(_11438_),
    .A(_11436_),
    .B(_11437_));
 sg13g2_a21oi_1 _42068_ (.A1(net5520),
    .A2(_11438_),
    .Y(_11439_),
    .B1(_11431_));
 sg13g2_a22oi_1 _42069_ (.Y(_11440_),
    .B1(_11439_),
    .B2(net5229),
    .A2(_11418_),
    .A1(net5210));
 sg13g2_a22oi_1 _42070_ (.Y(_11441_),
    .B1(net5102),
    .B2(_09515_),
    .A2(net6429),
    .A1(net3416));
 sg13g2_o21ai_1 _42071_ (.B1(_11441_),
    .Y(_00778_),
    .A1(net6851),
    .A2(_11440_));
 sg13g2_nand2_1 _42072_ (.Y(_11442_),
    .A(net5716),
    .B(_09550_));
 sg13g2_a21oi_1 _42073_ (.A1(_09624_),
    .A2(_11380_),
    .Y(_11443_),
    .B1(_09526_));
 sg13g2_o21ai_1 _42074_ (.B1(_09553_),
    .Y(_11444_),
    .A1(_09631_),
    .A2(_11443_));
 sg13g2_or3_1 _42075_ (.A(_09553_),
    .B(_09631_),
    .C(_11443_),
    .X(_11445_));
 sg13g2_nand2_1 _42076_ (.Y(_11446_),
    .A(_11444_),
    .B(_11445_));
 sg13g2_o21ai_1 _42077_ (.B1(_11442_),
    .Y(_11447_),
    .A1(net5717),
    .A2(_11446_));
 sg13g2_xnor2_1 _42078_ (.Y(_11448_),
    .A(net5457),
    .B(_11447_));
 sg13g2_nand2_1 _42079_ (.Y(_11449_),
    .A(_11432_),
    .B(_11436_));
 sg13g2_xnor2_1 _42080_ (.Y(_11450_),
    .A(_11448_),
    .B(_11449_));
 sg13g2_o21ai_1 _42081_ (.B1(net5954),
    .Y(_11451_),
    .A1(net5520),
    .A2(_11447_));
 sg13g2_a21oi_1 _42082_ (.A1(net5520),
    .A2(_11450_),
    .Y(_11452_),
    .B1(_11451_));
 sg13g2_a221oi_1 _42083_ (.B2(net5903),
    .C1(_11452_),
    .B1(_11430_),
    .A1(net5986),
    .Y(_11453_),
    .A2(_09501_));
 sg13g2_a21oi_1 _42084_ (.A1(net5279),
    .A2(_11453_),
    .Y(_11454_),
    .B1(net6851));
 sg13g2_o21ai_1 _42085_ (.B1(_11454_),
    .Y(_11455_),
    .A1(net5279),
    .A2(_09501_));
 sg13g2_o21ai_1 _42086_ (.B1(_11455_),
    .Y(_00779_),
    .A1(_18169_),
    .A2(net6497));
 sg13g2_a21oi_1 _42087_ (.A1(_09551_),
    .A2(_11444_),
    .Y(_11456_),
    .B1(_09546_));
 sg13g2_and3_1 _42088_ (.X(_11457_),
    .A(_09546_),
    .B(_09551_),
    .C(_11444_));
 sg13g2_nor3_1 _42089_ (.A(net5717),
    .B(_11456_),
    .C(_11457_),
    .Y(_11458_));
 sg13g2_a21o_2 _42090_ (.A2(_09544_),
    .A1(net5717),
    .B1(_11458_),
    .X(_11459_));
 sg13g2_nor2_1 _42091_ (.A(net5521),
    .B(_11459_),
    .Y(_11460_));
 sg13g2_nand2_1 _42092_ (.Y(_11461_),
    .A(net5413),
    .B(_11459_));
 sg13g2_xnor2_1 _42093_ (.Y(_11462_),
    .A(net5457),
    .B(_11459_));
 sg13g2_nand2_1 _42094_ (.Y(_11463_),
    .A(_11433_),
    .B(_11448_));
 sg13g2_o21ai_1 _42095_ (.B1(net5413),
    .Y(_11464_),
    .A1(_11430_),
    .A2(_11447_));
 sg13g2_o21ai_1 _42096_ (.B1(_11464_),
    .Y(_11465_),
    .A1(_11434_),
    .A2(_11463_));
 sg13g2_nand3_1 _42097_ (.B(_11433_),
    .C(_11448_),
    .A(_11399_),
    .Y(_11466_));
 sg13g2_or2_1 _42098_ (.X(_11467_),
    .B(_11466_),
    .A(_11420_));
 sg13g2_nor2_1 _42099_ (.A(_11408_),
    .B(_11467_),
    .Y(_11468_));
 sg13g2_or2_1 _42100_ (.X(_11469_),
    .B(_11468_),
    .A(_11465_));
 sg13g2_and2_1 _42101_ (.A(_11462_),
    .B(_11469_),
    .X(_11470_));
 sg13g2_xnor2_1 _42102_ (.Y(_11471_),
    .A(_11462_),
    .B(_11469_));
 sg13g2_a21oi_1 _42103_ (.A1(net5521),
    .A2(_11471_),
    .Y(_11472_),
    .B1(_11460_));
 sg13g2_a22oi_1 _42104_ (.Y(_11473_),
    .B1(_11472_),
    .B2(net5229),
    .A2(_11447_),
    .A1(net5211));
 sg13g2_a22oi_1 _42105_ (.Y(_11474_),
    .B1(net5104),
    .B2(_09510_),
    .A2(net6439),
    .A1(net3011));
 sg13g2_o21ai_1 _42106_ (.B1(_11474_),
    .Y(_00780_),
    .A1(net6851),
    .A2(_11473_));
 sg13g2_nor2_1 _42107_ (.A(net5758),
    .B(_09538_),
    .Y(_11475_));
 sg13g2_a21oi_1 _42108_ (.A1(_09626_),
    .A2(_11444_),
    .Y(_11476_),
    .B1(_09545_));
 sg13g2_xnor2_1 _42109_ (.Y(_11477_),
    .A(_09540_),
    .B(_11476_));
 sg13g2_a21oi_2 _42110_ (.B1(_11475_),
    .Y(_11478_),
    .A2(_11477_),
    .A1(net5759));
 sg13g2_nand2_1 _42111_ (.Y(_11479_),
    .A(net5413),
    .B(_11478_));
 sg13g2_nand2b_1 _42112_ (.Y(_11480_),
    .B(net5457),
    .A_N(_11478_));
 sg13g2_nand2_1 _42113_ (.Y(_11481_),
    .A(_11479_),
    .B(_11480_));
 sg13g2_a21oi_1 _42114_ (.A1(net5413),
    .A2(_11459_),
    .Y(_11482_),
    .B1(_11470_));
 sg13g2_xnor2_1 _42115_ (.Y(_11483_),
    .A(_11481_),
    .B(_11482_));
 sg13g2_o21ai_1 _42116_ (.B1(net5953),
    .Y(_11484_),
    .A1(net5521),
    .A2(_11478_));
 sg13g2_a21oi_1 _42117_ (.A1(net5521),
    .A2(_11483_),
    .Y(_11485_),
    .B1(_11484_));
 sg13g2_a221oi_1 _42118_ (.B2(net5903),
    .C1(_11485_),
    .B1(_11459_),
    .A1(net5986),
    .Y(_11486_),
    .A2(_09550_));
 sg13g2_a21oi_1 _42119_ (.A1(net5281),
    .A2(_11486_),
    .Y(_11487_),
    .B1(net6851));
 sg13g2_o21ai_1 _42120_ (.B1(_11487_),
    .Y(_11488_),
    .A1(net5279),
    .A2(_09550_));
 sg13g2_o21ai_1 _42121_ (.B1(_11488_),
    .Y(_00781_),
    .A1(_18167_),
    .A2(net6498));
 sg13g2_nor2_1 _42122_ (.A(net5758),
    .B(_09530_),
    .Y(_11489_));
 sg13g2_a21oi_1 _42123_ (.A1(_09540_),
    .A2(_11476_),
    .Y(_11490_),
    .B1(_09539_));
 sg13g2_xnor2_1 _42124_ (.Y(_11491_),
    .A(_09532_),
    .B(_11490_));
 sg13g2_a21oi_2 _42125_ (.B1(_11489_),
    .Y(_11492_),
    .A2(_11491_),
    .A1(net5758));
 sg13g2_or2_1 _42126_ (.X(_11493_),
    .B(_11492_),
    .A(net5457));
 sg13g2_xnor2_1 _42127_ (.Y(_11494_),
    .A(net5457),
    .B(_11492_));
 sg13g2_nand2_1 _42128_ (.Y(_11495_),
    .A(_11461_),
    .B(_11479_));
 sg13g2_o21ai_1 _42129_ (.B1(_11480_),
    .Y(_11496_),
    .A1(_11470_),
    .A2(_11495_));
 sg13g2_xor2_1 _42130_ (.B(_11496_),
    .A(_11494_),
    .X(_11497_));
 sg13g2_o21ai_1 _42131_ (.B1(net5956),
    .Y(_11498_),
    .A1(net5562),
    .A2(_11497_));
 sg13g2_a21oi_1 _42132_ (.A1(net5562),
    .A2(_11492_),
    .Y(_11499_),
    .B1(_11498_));
 sg13g2_a221oi_1 _42133_ (.B2(net5903),
    .C1(_11499_),
    .B1(_11478_),
    .A1(net5986),
    .Y(_11500_),
    .A2(_09544_));
 sg13g2_a21oi_1 _42134_ (.A1(net5279),
    .A2(_11500_),
    .Y(_11501_),
    .B1(net6854));
 sg13g2_o21ai_1 _42135_ (.B1(_11501_),
    .Y(_11502_),
    .A1(net5279),
    .A2(_09544_));
 sg13g2_o21ai_1 _42136_ (.B1(_11502_),
    .Y(_00782_),
    .A1(_18166_),
    .A2(net6498));
 sg13g2_nand2_1 _42137_ (.Y(_11503_),
    .A(net2662),
    .B(net6439));
 sg13g2_nor2_1 _42138_ (.A(net5759),
    .B(_09486_),
    .Y(_11504_));
 sg13g2_o21ai_1 _42139_ (.B1(_09612_),
    .Y(_11505_),
    .A1(_09354_),
    .A2(_09372_));
 sg13g2_nand2_1 _42140_ (.Y(_11506_),
    .A(_09633_),
    .B(_11505_));
 sg13g2_nand2_1 _42141_ (.Y(_11507_),
    .A(_09489_),
    .B(_11506_));
 sg13g2_xor2_1 _42142_ (.B(_11506_),
    .A(_09489_),
    .X(_11508_));
 sg13g2_a21oi_2 _42143_ (.B1(_11504_),
    .Y(_11509_),
    .A2(_11508_),
    .A1(net5759));
 sg13g2_inv_1 _42144_ (.Y(_11510_),
    .A(_11509_));
 sg13g2_xnor2_1 _42145_ (.Y(_11511_),
    .A(net5412),
    .B(_11509_));
 sg13g2_o21ai_1 _42146_ (.B1(_11493_),
    .Y(_11512_),
    .A1(_11494_),
    .A2(_11496_));
 sg13g2_xor2_1 _42147_ (.B(_11512_),
    .A(_11511_),
    .X(_11513_));
 sg13g2_a21oi_1 _42148_ (.A1(net5562),
    .A2(_11509_),
    .Y(_11514_),
    .B1(net5927));
 sg13g2_o21ai_1 _42149_ (.B1(_11514_),
    .Y(_11515_),
    .A1(net5562),
    .A2(_11513_));
 sg13g2_nor2_1 _42150_ (.A(net5882),
    .B(_11492_),
    .Y(_11516_));
 sg13g2_a21oi_1 _42151_ (.A1(net5986),
    .A2(_09538_),
    .Y(_11517_),
    .B1(_11516_));
 sg13g2_and3_1 _42152_ (.X(_11518_),
    .A(net5279),
    .B(_11515_),
    .C(_11517_));
 sg13g2_o21ai_1 _42153_ (.B1(net6880),
    .Y(_11519_),
    .A1(net5284),
    .A2(_09538_));
 sg13g2_o21ai_1 _42154_ (.B1(_11503_),
    .Y(_00783_),
    .A1(_11518_),
    .A2(_11519_));
 sg13g2_nand2_1 _42155_ (.Y(_11520_),
    .A(net5718),
    .B(_09480_));
 sg13g2_and2_1 _42156_ (.A(_09488_),
    .B(_11507_),
    .X(_11521_));
 sg13g2_xor2_1 _42157_ (.B(_11521_),
    .A(_09482_),
    .X(_11522_));
 sg13g2_o21ai_1 _42158_ (.B1(_11520_),
    .Y(_11523_),
    .A1(net5718),
    .A2(_11522_));
 sg13g2_nor2_1 _42159_ (.A(net5525),
    .B(_11523_),
    .Y(_11524_));
 sg13g2_nand2_1 _42160_ (.Y(_11525_),
    .A(net5409),
    .B(_11523_));
 sg13g2_xnor2_1 _42161_ (.Y(_11526_),
    .A(net5409),
    .B(_11523_));
 sg13g2_nor2b_1 _42162_ (.A(_11494_),
    .B_N(_11511_),
    .Y(_11527_));
 sg13g2_and4_1 _42163_ (.A(_11462_),
    .B(_11479_),
    .C(_11480_),
    .D(_11527_),
    .X(_11528_));
 sg13g2_nor2b_1 _42164_ (.A(_11467_),
    .B_N(_11528_),
    .Y(_11529_));
 sg13g2_o21ai_1 _42165_ (.B1(_11529_),
    .Y(_11530_),
    .A1(_11403_),
    .A2(_11404_));
 sg13g2_a21oi_1 _42166_ (.A1(_11492_),
    .A2(_11509_),
    .Y(_11531_),
    .B1(net5464));
 sg13g2_a221oi_1 _42167_ (.B2(_11465_),
    .C1(_11531_),
    .B1(_11528_),
    .A1(_11495_),
    .Y(_11532_),
    .A2(_11527_));
 sg13g2_nand2_1 _42168_ (.Y(_11533_),
    .A(_11406_),
    .B(_11529_));
 sg13g2_inv_1 _42169_ (.Y(_11534_),
    .A(_11533_));
 sg13g2_o21ai_1 _42170_ (.B1(_11534_),
    .Y(_11535_),
    .A1(_11270_),
    .A2(_11272_));
 sg13g2_and3_2 _42171_ (.X(_11536_),
    .A(_11530_),
    .B(_11532_),
    .C(_11535_));
 sg13g2_or2_1 _42172_ (.X(_11537_),
    .B(_11536_),
    .A(_11526_));
 sg13g2_xnor2_1 _42173_ (.Y(_11538_),
    .A(_11526_),
    .B(_11536_));
 sg13g2_a21oi_1 _42174_ (.A1(net5525),
    .A2(_11538_),
    .Y(_11539_),
    .B1(_11524_));
 sg13g2_a22oi_1 _42175_ (.Y(_11540_),
    .B1(_11539_),
    .B2(net5229),
    .A2(_11510_),
    .A1(net5212));
 sg13g2_a22oi_1 _42176_ (.Y(_11541_),
    .B1(net5104),
    .B2(_09531_),
    .A2(net6439),
    .A1(net3045));
 sg13g2_o21ai_1 _42177_ (.B1(_11541_),
    .Y(_00784_),
    .A1(net6854),
    .A2(_11540_));
 sg13g2_nand2_1 _42178_ (.Y(_11542_),
    .A(_11525_),
    .B(_11537_));
 sg13g2_nor2_1 _42179_ (.A(net5760),
    .B(_09468_),
    .Y(_11543_));
 sg13g2_a21o_1 _42180_ (.A2(_11507_),
    .A1(_09643_),
    .B1(_09481_),
    .X(_11544_));
 sg13g2_xnor2_1 _42181_ (.Y(_11545_),
    .A(_09471_),
    .B(_11544_));
 sg13g2_a21oi_2 _42182_ (.B1(_11543_),
    .Y(_11546_),
    .A2(_11545_),
    .A1(net5760));
 sg13g2_nand2b_1 _42183_ (.Y(_11547_),
    .B(net5459),
    .A_N(_11546_));
 sg13g2_xnor2_1 _42184_ (.Y(_11548_),
    .A(net5409),
    .B(_11546_));
 sg13g2_xor2_1 _42185_ (.B(_11548_),
    .A(_11542_),
    .X(_11549_));
 sg13g2_o21ai_1 _42186_ (.B1(net5956),
    .Y(_11550_),
    .A1(net5525),
    .A2(_11546_));
 sg13g2_a21oi_1 _42187_ (.A1(net5525),
    .A2(_11549_),
    .Y(_11551_),
    .B1(_11550_));
 sg13g2_a221oi_1 _42188_ (.B2(net5905),
    .C1(_11551_),
    .B1(_11523_),
    .A1(net5990),
    .Y(_11552_),
    .A2(_09487_));
 sg13g2_o21ai_1 _42189_ (.B1(net6881),
    .Y(_11553_),
    .A1(net5281),
    .A2(_09487_));
 sg13g2_a21oi_2 _42190_ (.B1(_11553_),
    .Y(_11554_),
    .A2(_11552_),
    .A1(net5281));
 sg13g2_a21o_1 _42191_ (.A2(net6433),
    .A1(net2480),
    .B1(_11554_),
    .X(_00785_));
 sg13g2_nand2_1 _42192_ (.Y(_11555_),
    .A(net2916),
    .B(net6439));
 sg13g2_o21ai_1 _42193_ (.B1(_09469_),
    .Y(_11556_),
    .A1(_09471_),
    .A2(_11544_));
 sg13g2_nor2_1 _42194_ (.A(net5759),
    .B(_09474_),
    .Y(_11557_));
 sg13g2_xnor2_1 _42195_ (.Y(_11558_),
    .A(_09476_),
    .B(_11556_));
 sg13g2_a21oi_2 _42196_ (.B1(_11557_),
    .Y(_11559_),
    .A2(_11558_),
    .A1(net5760));
 sg13g2_nand2_1 _42197_ (.Y(_11560_),
    .A(net5409),
    .B(_11559_));
 sg13g2_xnor2_1 _42198_ (.Y(_11561_),
    .A(net5459),
    .B(_11559_));
 sg13g2_o21ai_1 _42199_ (.B1(net5409),
    .Y(_11562_),
    .A1(_11523_),
    .A2(_11546_));
 sg13g2_nand2_1 _42200_ (.Y(_11563_),
    .A(_11537_),
    .B(_11562_));
 sg13g2_nand3_1 _42201_ (.B(_11561_),
    .C(_11563_),
    .A(_11547_),
    .Y(_11564_));
 sg13g2_a21o_1 _42202_ (.A2(_11563_),
    .A1(_11547_),
    .B1(_11561_),
    .X(_11565_));
 sg13g2_a21o_1 _42203_ (.A2(_11565_),
    .A1(_11564_),
    .B1(net5562),
    .X(_11566_));
 sg13g2_o21ai_1 _42204_ (.B1(_11566_),
    .Y(_11567_),
    .A1(net5525),
    .A2(_11559_));
 sg13g2_nor2_1 _42205_ (.A(net5153),
    .B(_11567_),
    .Y(_11568_));
 sg13g2_a221oi_1 _42206_ (.B2(net5212),
    .C1(_11568_),
    .B1(_11546_),
    .A1(net5162),
    .Y(_11569_),
    .A2(_09480_));
 sg13g2_o21ai_1 _42207_ (.B1(_11555_),
    .Y(_00786_),
    .A1(net6854),
    .A2(_11569_));
 sg13g2_and2_1 _42208_ (.A(net5718),
    .B(_09458_),
    .X(_11570_));
 sg13g2_a21oi_1 _42209_ (.A1(_09633_),
    .A2(_11505_),
    .Y(_11571_),
    .B1(_09491_));
 sg13g2_nor3_1 _42210_ (.A(_09644_),
    .B(_09645_),
    .C(_11571_),
    .Y(_11572_));
 sg13g2_or2_1 _42211_ (.X(_11573_),
    .B(_11572_),
    .A(_09460_));
 sg13g2_a21oi_1 _42212_ (.A1(_09460_),
    .A2(_11572_),
    .Y(_11574_),
    .B1(net5718));
 sg13g2_a21o_2 _42213_ (.A2(_11574_),
    .A1(_11573_),
    .B1(_11570_),
    .X(_11575_));
 sg13g2_xnor2_1 _42214_ (.Y(_11576_),
    .A(net5460),
    .B(_11575_));
 sg13g2_nand2_1 _42215_ (.Y(_11577_),
    .A(_11560_),
    .B(_11564_));
 sg13g2_xnor2_1 _42216_ (.Y(_11578_),
    .A(_11576_),
    .B(_11577_));
 sg13g2_o21ai_1 _42217_ (.B1(net5956),
    .Y(_11579_),
    .A1(net5525),
    .A2(_11575_));
 sg13g2_a21oi_1 _42218_ (.A1(net5525),
    .A2(_11578_),
    .Y(_11580_),
    .B1(_11579_));
 sg13g2_a221oi_1 _42219_ (.B2(net5905),
    .C1(_11580_),
    .B1(_11559_),
    .A1(net5990),
    .Y(_11581_),
    .A2(_09468_));
 sg13g2_o21ai_1 _42220_ (.B1(net6881),
    .Y(_11582_),
    .A1(net5281),
    .A2(_09468_));
 sg13g2_a21oi_1 _42221_ (.A1(net5281),
    .A2(_11581_),
    .Y(_11583_),
    .B1(_11582_));
 sg13g2_a21o_1 _42222_ (.A2(net6439),
    .A1(net7298),
    .B1(_11583_),
    .X(_00787_));
 sg13g2_a21oi_1 _42223_ (.A1(_09459_),
    .A2(_11573_),
    .Y(_11584_),
    .B1(_09456_));
 sg13g2_and3_1 _42224_ (.X(_11585_),
    .A(_09456_),
    .B(_09459_),
    .C(_11573_));
 sg13g2_nor3_1 _42225_ (.A(net5718),
    .B(_11584_),
    .C(_11585_),
    .Y(_11586_));
 sg13g2_a21o_2 _42226_ (.A2(_09455_),
    .A1(net5721),
    .B1(_11586_),
    .X(_11587_));
 sg13g2_nor2_1 _42227_ (.A(net5525),
    .B(_11587_),
    .Y(_11588_));
 sg13g2_nand2_1 _42228_ (.Y(_11589_),
    .A(net5409),
    .B(_11587_));
 sg13g2_xnor2_1 _42229_ (.Y(_11590_),
    .A(net5459),
    .B(_11587_));
 sg13g2_nand2_1 _42230_ (.Y(_11591_),
    .A(_11561_),
    .B(_11576_));
 sg13g2_o21ai_1 _42231_ (.B1(_11560_),
    .Y(_11592_),
    .A1(_11562_),
    .A2(_11591_));
 sg13g2_a21o_1 _42232_ (.A2(_11575_),
    .A1(net5411),
    .B1(_11592_),
    .X(_11593_));
 sg13g2_nor3_1 _42233_ (.A(_11526_),
    .B(_11548_),
    .C(_11591_),
    .Y(_11594_));
 sg13g2_nand2b_1 _42234_ (.Y(_11595_),
    .B(_11594_),
    .A_N(_11536_));
 sg13g2_nand2b_2 _42235_ (.Y(_11596_),
    .B(_11595_),
    .A_N(_11593_));
 sg13g2_and2_1 _42236_ (.A(_11590_),
    .B(_11596_),
    .X(_11597_));
 sg13g2_xnor2_1 _42237_ (.Y(_11598_),
    .A(_11590_),
    .B(_11596_));
 sg13g2_a21oi_1 _42238_ (.A1(net5526),
    .A2(_11598_),
    .Y(_11599_),
    .B1(_11588_));
 sg13g2_a22oi_1 _42239_ (.Y(_11600_),
    .B1(_11599_),
    .B2(net5229),
    .A2(_11575_),
    .A1(net5212));
 sg13g2_a22oi_1 _42240_ (.Y(_11601_),
    .B1(net5104),
    .B2(_09474_),
    .A2(net6439),
    .A1(net3579));
 sg13g2_o21ai_1 _42241_ (.B1(_11601_),
    .Y(_00788_),
    .A1(net6854),
    .A2(_11600_));
 sg13g2_nand2_1 _42242_ (.Y(_11602_),
    .A(net3408),
    .B(net6441));
 sg13g2_or2_1 _42243_ (.X(_11603_),
    .B(_09445_),
    .A(net5759));
 sg13g2_o21ai_1 _42244_ (.B1(_09647_),
    .Y(_11604_),
    .A1(_09460_),
    .A2(_11572_));
 sg13g2_o21ai_1 _42245_ (.B1(_11604_),
    .Y(_11605_),
    .A1(net5655),
    .A2(_09455_));
 sg13g2_xor2_1 _42246_ (.B(_11605_),
    .A(_09447_),
    .X(_11606_));
 sg13g2_o21ai_1 _42247_ (.B1(_11603_),
    .Y(_11607_),
    .A1(net5718),
    .A2(_11606_));
 sg13g2_nand2_1 _42248_ (.Y(_11608_),
    .A(net5459),
    .B(_11607_));
 sg13g2_xnor2_1 _42249_ (.Y(_11609_),
    .A(net5459),
    .B(_11607_));
 sg13g2_a21oi_1 _42250_ (.A1(net5411),
    .A2(_11587_),
    .Y(_11610_),
    .B1(_11597_));
 sg13g2_xor2_1 _42251_ (.B(_11610_),
    .A(_11609_),
    .X(_11611_));
 sg13g2_a21oi_1 _42252_ (.A1(net5561),
    .A2(_11607_),
    .Y(_11612_),
    .B1(net5927));
 sg13g2_o21ai_1 _42253_ (.B1(_11612_),
    .Y(_11613_),
    .A1(net5561),
    .A2(_11611_));
 sg13g2_a22oi_1 _42254_ (.Y(_11614_),
    .B1(_11587_),
    .B2(net5905),
    .A2(_09458_),
    .A1(net5990));
 sg13g2_and3_1 _42255_ (.X(_11615_),
    .A(net5286),
    .B(_11613_),
    .C(_11614_));
 sg13g2_o21ai_1 _42256_ (.B1(net6881),
    .Y(_11616_),
    .A1(net5288),
    .A2(_09458_));
 sg13g2_o21ai_1 _42257_ (.B1(_11602_),
    .Y(_00789_),
    .A1(_11615_),
    .A2(_11616_));
 sg13g2_nand2_1 _42258_ (.Y(_11617_),
    .A(net5718),
    .B(_09450_));
 sg13g2_o21ai_1 _42259_ (.B1(_09446_),
    .Y(_11618_),
    .A1(_09447_),
    .A2(_11605_));
 sg13g2_xor2_1 _42260_ (.B(_11618_),
    .A(_09452_),
    .X(_11619_));
 sg13g2_o21ai_1 _42261_ (.B1(_11617_),
    .Y(_11620_),
    .A1(net5718),
    .A2(_11619_));
 sg13g2_nor2_1 _42262_ (.A(net5522),
    .B(_11620_),
    .Y(_11621_));
 sg13g2_nand2_1 _42263_ (.Y(_11622_),
    .A(net5409),
    .B(_11620_));
 sg13g2_xnor2_1 _42264_ (.Y(_11623_),
    .A(net5459),
    .B(_11620_));
 sg13g2_inv_1 _42265_ (.Y(_11624_),
    .A(_11623_));
 sg13g2_o21ai_1 _42266_ (.B1(_11589_),
    .Y(_11625_),
    .A1(net5459),
    .A2(_11607_));
 sg13g2_o21ai_1 _42267_ (.B1(_11608_),
    .Y(_11626_),
    .A1(_11597_),
    .A2(_11625_));
 sg13g2_xnor2_1 _42268_ (.Y(_11627_),
    .A(_11624_),
    .B(_11626_));
 sg13g2_a21oi_1 _42269_ (.A1(net5522),
    .A2(_11627_),
    .Y(_11628_),
    .B1(_11621_));
 sg13g2_a22oi_1 _42270_ (.Y(_11629_),
    .B1(_11628_),
    .B2(net5233),
    .A2(_09455_),
    .A1(net5162));
 sg13g2_o21ai_1 _42271_ (.B1(_11629_),
    .Y(_11630_),
    .A1(net5120),
    .A2(_11607_));
 sg13g2_a22oi_1 _42272_ (.Y(_11631_),
    .B1(net6881),
    .B2(_11630_),
    .A2(net6441),
    .A1(net3236));
 sg13g2_inv_1 _42273_ (.Y(_00790_),
    .A(_11631_));
 sg13g2_nand2_1 _42274_ (.Y(_11632_),
    .A(net5723),
    .B(_09433_));
 sg13g2_a21oi_1 _42275_ (.A1(_09633_),
    .A2(_11505_),
    .Y(_11633_),
    .B1(_09493_));
 sg13g2_o21ai_1 _42276_ (.B1(_09435_),
    .Y(_11634_),
    .A1(_09650_),
    .A2(_11633_));
 sg13g2_or3_1 _42277_ (.A(_09435_),
    .B(_09650_),
    .C(_11633_),
    .X(_11635_));
 sg13g2_nand2_1 _42278_ (.Y(_11636_),
    .A(_11634_),
    .B(_11635_));
 sg13g2_o21ai_1 _42279_ (.B1(_11632_),
    .Y(_11637_),
    .A1(net5723),
    .A2(_11636_));
 sg13g2_xnor2_1 _42280_ (.Y(_11638_),
    .A(net5459),
    .B(_11637_));
 sg13g2_o21ai_1 _42281_ (.B1(_11622_),
    .Y(_11639_),
    .A1(_11624_),
    .A2(_11626_));
 sg13g2_xnor2_1 _42282_ (.Y(_11640_),
    .A(_11638_),
    .B(_11639_));
 sg13g2_o21ai_1 _42283_ (.B1(net5956),
    .Y(_11641_),
    .A1(net5522),
    .A2(_11637_));
 sg13g2_a21oi_1 _42284_ (.A1(net5522),
    .A2(_11640_),
    .Y(_11642_),
    .B1(_11641_));
 sg13g2_a221oi_1 _42285_ (.B2(net5905),
    .C1(_11642_),
    .B1(_11620_),
    .A1(net5990),
    .Y(_11643_),
    .A2(_09445_));
 sg13g2_a21oi_1 _42286_ (.A1(net5288),
    .A2(_11643_),
    .Y(_11644_),
    .B1(net6854));
 sg13g2_o21ai_1 _42287_ (.B1(_11644_),
    .Y(_11645_),
    .A1(net5288),
    .A2(_09445_));
 sg13g2_o21ai_1 _42288_ (.B1(_11645_),
    .Y(_00791_),
    .A1(_18163_),
    .A2(net6498));
 sg13g2_nand2_1 _42289_ (.Y(_11646_),
    .A(net2483),
    .B(net6441));
 sg13g2_nand2_1 _42290_ (.Y(_11647_),
    .A(_09434_),
    .B(_11634_));
 sg13g2_xnor2_1 _42291_ (.Y(_11648_),
    .A(_09429_),
    .B(_11647_));
 sg13g2_nand2_1 _42292_ (.Y(_11649_),
    .A(net5723),
    .B(_09427_));
 sg13g2_o21ai_1 _42293_ (.B1(_11649_),
    .Y(_11650_),
    .A1(net5723),
    .A2(_11648_));
 sg13g2_inv_1 _42294_ (.Y(_11651_),
    .A(_11650_));
 sg13g2_xnor2_1 _42295_ (.Y(_11652_),
    .A(net5462),
    .B(_11651_));
 sg13g2_nand3_1 _42296_ (.B(_11625_),
    .C(_11638_),
    .A(_11623_),
    .Y(_11653_));
 sg13g2_o21ai_1 _42297_ (.B1(net5409),
    .Y(_11654_),
    .A1(_11620_),
    .A2(_11637_));
 sg13g2_nand2_1 _42298_ (.Y(_11655_),
    .A(_11653_),
    .B(_11654_));
 sg13g2_nand3_1 _42299_ (.B(_11623_),
    .C(_11638_),
    .A(_11590_),
    .Y(_11656_));
 sg13g2_nor2_1 _42300_ (.A(_11609_),
    .B(_11656_),
    .Y(_11657_));
 sg13g2_a21oi_1 _42301_ (.A1(_11593_),
    .A2(_11657_),
    .Y(_11658_),
    .B1(_11655_));
 sg13g2_a21o_1 _42302_ (.A2(_11657_),
    .A1(_11596_),
    .B1(_11655_),
    .X(_11659_));
 sg13g2_nor2b_1 _42303_ (.A(_11652_),
    .B_N(_11659_),
    .Y(_11660_));
 sg13g2_nor2b_1 _42304_ (.A(_11659_),
    .B_N(_11652_),
    .Y(_11661_));
 sg13g2_o21ai_1 _42305_ (.B1(net5528),
    .Y(_11662_),
    .A1(_11660_),
    .A2(_11661_));
 sg13g2_o21ai_1 _42306_ (.B1(_11662_),
    .Y(_11663_),
    .A1(net5528),
    .A2(_11650_));
 sg13g2_nor2_1 _42307_ (.A(net5153),
    .B(_11663_),
    .Y(_11664_));
 sg13g2_a221oi_1 _42308_ (.B2(net5214),
    .C1(_11664_),
    .B1(_11637_),
    .A1(net5162),
    .Y(_11665_),
    .A2(_09450_));
 sg13g2_o21ai_1 _42309_ (.B1(_11646_),
    .Y(_00792_),
    .A1(net6854),
    .A2(_11665_));
 sg13g2_nor2_1 _42310_ (.A(net5763),
    .B(_09416_),
    .Y(_11666_));
 sg13g2_a21oi_1 _42311_ (.A1(_09635_),
    .A2(_11634_),
    .Y(_11667_),
    .B1(_09428_));
 sg13g2_nand2b_1 _42312_ (.Y(_11668_),
    .B(_11667_),
    .A_N(_09418_));
 sg13g2_xor2_1 _42313_ (.B(_11667_),
    .A(_09418_),
    .X(_11669_));
 sg13g2_a21oi_2 _42314_ (.B1(_11666_),
    .Y(_11670_),
    .A2(_11669_),
    .A1(net5763));
 sg13g2_nand2b_1 _42315_ (.Y(_11671_),
    .B(net5462),
    .A_N(_11670_));
 sg13g2_nand2_1 _42316_ (.Y(_11672_),
    .A(net5414),
    .B(_11670_));
 sg13g2_xnor2_1 _42317_ (.Y(_11673_),
    .A(net5414),
    .B(_11670_));
 sg13g2_a21oi_1 _42318_ (.A1(net5414),
    .A2(_11650_),
    .Y(_11674_),
    .B1(_11660_));
 sg13g2_xnor2_1 _42319_ (.Y(_11675_),
    .A(_11673_),
    .B(_11674_));
 sg13g2_o21ai_1 _42320_ (.B1(net5957),
    .Y(_11676_),
    .A1(net5528),
    .A2(_11670_));
 sg13g2_a21oi_1 _42321_ (.A1(net5528),
    .A2(_11675_),
    .Y(_11677_),
    .B1(_11676_));
 sg13g2_a221oi_1 _42322_ (.B2(net5906),
    .C1(_11677_),
    .B1(_11650_),
    .A1(net5991),
    .Y(_11678_),
    .A2(_09433_));
 sg13g2_o21ai_1 _42323_ (.B1(net6882),
    .Y(_11679_),
    .A1(net5288),
    .A2(_09433_));
 sg13g2_a21oi_1 _42324_ (.A1(net5288),
    .A2(_11678_),
    .Y(_11680_),
    .B1(_11679_));
 sg13g2_a21o_1 _42325_ (.A2(net6441),
    .A1(net3583),
    .B1(_11680_),
    .X(_00793_));
 sg13g2_nand2_1 _42326_ (.Y(_11681_),
    .A(net5722),
    .B(_09421_));
 sg13g2_nand2_1 _42327_ (.Y(_11682_),
    .A(_09417_),
    .B(_11668_));
 sg13g2_xnor2_1 _42328_ (.Y(_11683_),
    .A(_09423_),
    .B(_11682_));
 sg13g2_o21ai_1 _42329_ (.B1(_11681_),
    .Y(_11684_),
    .A1(net5722),
    .A2(_11683_));
 sg13g2_nor2_1 _42330_ (.A(net5528),
    .B(_11684_),
    .Y(_11685_));
 sg13g2_nand2_1 _42331_ (.Y(_11686_),
    .A(net5414),
    .B(_11684_));
 sg13g2_xnor2_1 _42332_ (.Y(_11687_),
    .A(net5462),
    .B(_11684_));
 sg13g2_inv_1 _42333_ (.Y(_11688_),
    .A(_11687_));
 sg13g2_o21ai_1 _42334_ (.B1(_11672_),
    .Y(_11689_),
    .A1(net5462),
    .A2(_11651_));
 sg13g2_o21ai_1 _42335_ (.B1(_11671_),
    .Y(_11690_),
    .A1(_11660_),
    .A2(_11689_));
 sg13g2_xnor2_1 _42336_ (.Y(_11691_),
    .A(_11688_),
    .B(_11690_));
 sg13g2_a21oi_1 _42337_ (.A1(net5528),
    .A2(_11691_),
    .Y(_11692_),
    .B1(_11685_));
 sg13g2_a22oi_1 _42338_ (.Y(_11693_),
    .B1(_11692_),
    .B2(net5233),
    .A2(_11670_),
    .A1(net5212));
 sg13g2_a22oi_1 _42339_ (.Y(_11694_),
    .B1(net5104),
    .B2(_09427_),
    .A2(net6441),
    .A1(net3681));
 sg13g2_o21ai_1 _42340_ (.B1(_11694_),
    .Y(_00794_),
    .A1(net6856),
    .A2(_11693_));
 sg13g2_o21ai_1 _42341_ (.B1(_09436_),
    .Y(_11695_),
    .A1(_09650_),
    .A2(_11633_));
 sg13g2_a21oi_1 _42342_ (.A1(_09639_),
    .A2(_11695_),
    .Y(_11696_),
    .B1(_09401_));
 sg13g2_and3_1 _42343_ (.X(_11697_),
    .A(_09401_),
    .B(_09639_),
    .C(_11695_));
 sg13g2_nor3_1 _42344_ (.A(net5722),
    .B(_11696_),
    .C(_11697_),
    .Y(_11698_));
 sg13g2_a21oi_2 _42345_ (.B1(_11698_),
    .Y(_11699_),
    .A2(_09399_),
    .A1(net5722));
 sg13g2_or2_1 _42346_ (.X(_11700_),
    .B(_11699_),
    .A(net5462));
 sg13g2_xnor2_1 _42347_ (.Y(_11701_),
    .A(net5414),
    .B(_11699_));
 sg13g2_o21ai_1 _42348_ (.B1(_11686_),
    .Y(_11702_),
    .A1(_11688_),
    .A2(_11690_));
 sg13g2_xor2_1 _42349_ (.B(_11702_),
    .A(_11701_),
    .X(_11703_));
 sg13g2_a21oi_1 _42350_ (.A1(net5563),
    .A2(_11699_),
    .Y(_11704_),
    .B1(net5928));
 sg13g2_o21ai_1 _42351_ (.B1(_11704_),
    .Y(_11705_),
    .A1(net5563),
    .A2(_11703_));
 sg13g2_a22oi_1 _42352_ (.Y(_11706_),
    .B1(_11684_),
    .B2(net5906),
    .A2(_09416_),
    .A1(net5991));
 sg13g2_nand3_1 _42353_ (.B(_11705_),
    .C(_11706_),
    .A(net5286),
    .Y(_11707_));
 sg13g2_nor2_1 _42354_ (.A(net5287),
    .B(_09416_),
    .Y(_11708_));
 sg13g2_nor2_1 _42355_ (.A(net6856),
    .B(_11708_),
    .Y(_11709_));
 sg13g2_a22oi_1 _42356_ (.Y(_11710_),
    .B1(_11707_),
    .B2(_11709_),
    .A2(net6441),
    .A1(net2614));
 sg13g2_inv_1 _42357_ (.Y(_00795_),
    .A(_11710_));
 sg13g2_nand2_1 _42358_ (.Y(_11711_),
    .A(net2979),
    .B(net6441));
 sg13g2_nor2_1 _42359_ (.A(_09400_),
    .B(_11696_),
    .Y(_11712_));
 sg13g2_xnor2_1 _42360_ (.Y(_11713_),
    .A(_09408_),
    .B(_11712_));
 sg13g2_nand2_1 _42361_ (.Y(_11714_),
    .A(net5763),
    .B(_11713_));
 sg13g2_o21ai_1 _42362_ (.B1(_11714_),
    .Y(_11715_),
    .A1(net5763),
    .A2(_09405_));
 sg13g2_nand2_1 _42363_ (.Y(_11716_),
    .A(net5415),
    .B(_11715_));
 sg13g2_xnor2_1 _42364_ (.Y(_11717_),
    .A(net5462),
    .B(_11715_));
 sg13g2_nand3_1 _42365_ (.B(_11689_),
    .C(_11701_),
    .A(_11687_),
    .Y(_11718_));
 sg13g2_nand3_1 _42366_ (.B(_11700_),
    .C(_11718_),
    .A(_11686_),
    .Y(_11719_));
 sg13g2_nor2_1 _42367_ (.A(_11652_),
    .B(_11673_),
    .Y(_11720_));
 sg13g2_nand3_1 _42368_ (.B(_11701_),
    .C(_11720_),
    .A(_11687_),
    .Y(_11721_));
 sg13g2_inv_1 _42369_ (.Y(_11722_),
    .A(_11721_));
 sg13g2_a21oi_1 _42370_ (.A1(_11659_),
    .A2(_11722_),
    .Y(_11723_),
    .B1(_11719_));
 sg13g2_nand2b_1 _42371_ (.Y(_11724_),
    .B(_11717_),
    .A_N(_11723_));
 sg13g2_xor2_1 _42372_ (.B(_11723_),
    .A(_11717_),
    .X(_11725_));
 sg13g2_o21ai_1 _42373_ (.B1(net5957),
    .Y(_11726_),
    .A1(net5528),
    .A2(_11715_));
 sg13g2_a21o_1 _42374_ (.A2(_11725_),
    .A1(net5528),
    .B1(_11726_),
    .X(_11727_));
 sg13g2_o21ai_1 _42375_ (.B1(_11727_),
    .Y(_11728_),
    .A1(net5882),
    .A2(_11699_));
 sg13g2_a221oi_1 _42376_ (.B2(_09421_),
    .C1(_11728_),
    .B1(net5991),
    .A1(net5321),
    .Y(_11729_),
    .A2(net5317));
 sg13g2_o21ai_1 _42377_ (.B1(net6882),
    .Y(_11730_),
    .A1(net5288),
    .A2(_09421_));
 sg13g2_o21ai_1 _42378_ (.B1(_11711_),
    .Y(_00796_),
    .A1(_11729_),
    .A2(_11730_));
 sg13g2_nand2_1 _42379_ (.Y(_11731_),
    .A(_11716_),
    .B(_11724_));
 sg13g2_nor2_1 _42380_ (.A(net5763),
    .B(_09387_),
    .Y(_11732_));
 sg13g2_o21ai_1 _42381_ (.B1(_09407_),
    .Y(_11733_),
    .A1(_09640_),
    .A2(_11696_));
 sg13g2_xor2_1 _42382_ (.B(_11733_),
    .A(_09391_),
    .X(_11734_));
 sg13g2_a21oi_2 _42383_ (.B1(_11732_),
    .Y(_11735_),
    .A2(_11734_),
    .A1(net5763));
 sg13g2_nor2_1 _42384_ (.A(net5415),
    .B(_11735_),
    .Y(_11736_));
 sg13g2_xnor2_1 _42385_ (.Y(_11737_),
    .A(net5463),
    .B(_11735_));
 sg13g2_xnor2_1 _42386_ (.Y(_11738_),
    .A(_11731_),
    .B(_11737_));
 sg13g2_o21ai_1 _42387_ (.B1(net5957),
    .Y(_11739_),
    .A1(net5529),
    .A2(_11735_));
 sg13g2_a21oi_1 _42388_ (.A1(net5529),
    .A2(_11738_),
    .Y(_11740_),
    .B1(_11739_));
 sg13g2_a221oi_1 _42389_ (.B2(net5906),
    .C1(_11740_),
    .B1(_11715_),
    .A1(net5992),
    .Y(_11741_),
    .A2(_09399_));
 sg13g2_o21ai_1 _42390_ (.B1(net6882),
    .Y(_11742_),
    .A1(net5287),
    .A2(_09399_));
 sg13g2_a21oi_1 _42391_ (.A1(net5287),
    .A2(_11741_),
    .Y(_11743_),
    .B1(_11742_));
 sg13g2_a21o_1 _42392_ (.A2(net6441),
    .A1(net2120),
    .B1(_11743_),
    .X(_00797_));
 sg13g2_o21ai_1 _42393_ (.B1(_09389_),
    .Y(_11744_),
    .A1(_09390_),
    .A2(_11733_));
 sg13g2_xor2_1 _42394_ (.B(_11744_),
    .A(_09395_),
    .X(_11745_));
 sg13g2_nand2_1 _42395_ (.Y(_11746_),
    .A(net5723),
    .B(_09394_));
 sg13g2_o21ai_1 _42396_ (.B1(_11746_),
    .Y(_11747_),
    .A1(net5722),
    .A2(_11745_));
 sg13g2_nand2_1 _42397_ (.Y(_11748_),
    .A(net5414),
    .B(_11747_));
 sg13g2_inv_1 _42398_ (.Y(_11749_),
    .A(_11748_));
 sg13g2_xnor2_1 _42399_ (.Y(_11750_),
    .A(net5462),
    .B(_11747_));
 sg13g2_o21ai_1 _42400_ (.B1(net5414),
    .Y(_11751_),
    .A1(_11715_),
    .A2(_11735_));
 sg13g2_a21oi_1 _42401_ (.A1(_11724_),
    .A2(_11751_),
    .Y(_11752_),
    .B1(_11736_));
 sg13g2_xnor2_1 _42402_ (.Y(_11753_),
    .A(_11750_),
    .B(_11752_));
 sg13g2_a21oi_1 _42403_ (.A1(net5529),
    .A2(_11753_),
    .Y(_11754_),
    .B1(net5927));
 sg13g2_o21ai_1 _42404_ (.B1(_11754_),
    .Y(_11755_),
    .A1(net5529),
    .A2(_11747_));
 sg13g2_nor2_1 _42405_ (.A(net6008),
    .B(_09405_),
    .Y(_11756_));
 sg13g2_a21oi_1 _42406_ (.A1(net5906),
    .A2(_11735_),
    .Y(_11757_),
    .B1(_11756_));
 sg13g2_nand3_1 _42407_ (.B(_11755_),
    .C(_11757_),
    .A(net5287),
    .Y(_11758_));
 sg13g2_nor2b_1 _42408_ (.A(net5287),
    .B_N(_09405_),
    .Y(_11759_));
 sg13g2_nor2_1 _42409_ (.A(net6856),
    .B(_11759_),
    .Y(_11760_));
 sg13g2_a22oi_1 _42410_ (.Y(_11761_),
    .B1(_11758_),
    .B2(_11760_),
    .A2(net6444),
    .A1(net3074));
 sg13g2_inv_1 _42411_ (.Y(_00798_),
    .A(_11761_));
 sg13g2_nand2_1 _42412_ (.Y(_11762_),
    .A(net2436),
    .B(net6444));
 sg13g2_a21oi_1 _42413_ (.A1(net1067),
    .A2(_09652_),
    .Y(_11763_),
    .B1(_09655_));
 sg13g2_and3_1 _42414_ (.X(_11764_),
    .A(net1067),
    .B(_09652_),
    .C(_09655_));
 sg13g2_nor3_1 _42415_ (.A(net5732),
    .B(_11763_),
    .C(_11764_),
    .Y(_11765_));
 sg13g2_a21oi_2 _42416_ (.B1(_11765_),
    .Y(_11766_),
    .A2(_08973_),
    .A1(net5732));
 sg13g2_nor2_1 _42417_ (.A(net5462),
    .B(_11766_),
    .Y(_11767_));
 sg13g2_xnor2_1 _42418_ (.Y(_11768_),
    .A(net5414),
    .B(_11766_));
 sg13g2_a21oi_1 _42419_ (.A1(_11750_),
    .A2(_11752_),
    .Y(_11769_),
    .B1(_11749_));
 sg13g2_xnor2_1 _42420_ (.Y(_11770_),
    .A(_11768_),
    .B(_11769_));
 sg13g2_a21oi_1 _42421_ (.A1(net5563),
    .A2(_11766_),
    .Y(_11771_),
    .B1(net5927));
 sg13g2_o21ai_1 _42422_ (.B1(_11771_),
    .Y(_11772_),
    .A1(net5563),
    .A2(_11770_));
 sg13g2_a22oi_1 _42423_ (.Y(_11773_),
    .B1(_11747_),
    .B2(net5906),
    .A2(_09387_),
    .A1(net5992));
 sg13g2_and3_1 _42424_ (.X(_11774_),
    .A(net5287),
    .B(_11772_),
    .C(_11773_));
 sg13g2_o21ai_1 _42425_ (.B1(net6882),
    .Y(_11775_),
    .A1(net5287),
    .A2(_09387_));
 sg13g2_o21ai_1 _42426_ (.B1(_11762_),
    .Y(_00799_),
    .A1(_11774_),
    .A2(_11775_));
 sg13g2_nor2_1 _42427_ (.A(_08974_),
    .B(_11763_),
    .Y(_11776_));
 sg13g2_o21ai_1 _42428_ (.B1(_09653_),
    .Y(_11777_),
    .A1(_08974_),
    .A2(_11763_));
 sg13g2_xor2_1 _42429_ (.B(_11776_),
    .A(_09654_),
    .X(_11778_));
 sg13g2_mux2_1 _42430_ (.A0(_08968_),
    .A1(_11778_),
    .S(net5770),
    .X(_11779_));
 sg13g2_inv_1 _42431_ (.Y(_11780_),
    .A(_11779_));
 sg13g2_nor2_1 _42432_ (.A(net5545),
    .B(_11779_),
    .Y(_11781_));
 sg13g2_xnor2_1 _42433_ (.Y(_11782_),
    .A(net5424),
    .B(_11780_));
 sg13g2_nand2_1 _42434_ (.Y(_11783_),
    .A(_11750_),
    .B(_11768_));
 sg13g2_nand2_1 _42435_ (.Y(_11784_),
    .A(_11717_),
    .B(_11737_));
 sg13g2_nor2_1 _42436_ (.A(_11783_),
    .B(_11784_),
    .Y(_11785_));
 sg13g2_nand4_1 _42437_ (.B(_11657_),
    .C(_11722_),
    .A(_11594_),
    .Y(_11786_),
    .D(_11785_));
 sg13g2_nor2_1 _42438_ (.A(_11533_),
    .B(_11786_),
    .Y(_11787_));
 sg13g2_o21ai_1 _42439_ (.B1(_11787_),
    .Y(_11788_),
    .A1(_11272_),
    .A2(_11270_));
 sg13g2_a21oi_2 _42440_ (.B1(_11786_),
    .Y(_11789_),
    .A2(_11532_),
    .A1(_11530_));
 sg13g2_o21ai_1 _42441_ (.B1(_11748_),
    .Y(_11790_),
    .A1(_11751_),
    .A2(_11783_));
 sg13g2_a21o_1 _42442_ (.A2(_11785_),
    .A1(_11719_),
    .B1(_11790_),
    .X(_11791_));
 sg13g2_nor4_1 _42443_ (.A(_11658_),
    .B(_11721_),
    .C(_11783_),
    .D(_11784_),
    .Y(_11792_));
 sg13g2_nor4_2 _42444_ (.A(_11767_),
    .B(_11791_),
    .C(_11789_),
    .Y(_11793_),
    .D(_11792_));
 sg13g2_nand2_2 _42445_ (.Y(_11794_),
    .A(net1074),
    .B(net1144));
 sg13g2_nand2_1 _42446_ (.Y(_11795_),
    .A(_11782_),
    .B(_11794_));
 sg13g2_xnor2_1 _42447_ (.Y(_11796_),
    .A(_11782_),
    .B(_11794_));
 sg13g2_a21oi_1 _42448_ (.A1(net5545),
    .A2(_11796_),
    .Y(_11797_),
    .B1(_11781_));
 sg13g2_nand2_1 _42449_ (.Y(_11798_),
    .A(net5230),
    .B(_11797_));
 sg13g2_o21ai_1 _42450_ (.B1(_11798_),
    .Y(_11799_),
    .A1(net5120),
    .A2(_11766_));
 sg13g2_a22oi_1 _42451_ (.Y(_11800_),
    .B1(_11799_),
    .B2(net6884),
    .A2(_09394_),
    .A1(net5109));
 sg13g2_o21ai_1 _42452_ (.B1(_11800_),
    .Y(_00800_),
    .A1(_18160_),
    .A2(net6504));
 sg13g2_nand2_1 _42453_ (.Y(_11801_),
    .A(net2253),
    .B(net6470));
 sg13g2_o21ai_1 _42454_ (.B1(_11795_),
    .Y(_11802_),
    .A1(net5469),
    .A2(_11780_));
 sg13g2_a21o_1 _42455_ (.A2(_11777_),
    .A1(_08969_),
    .B1(_08957_),
    .X(_11803_));
 sg13g2_nand3_1 _42456_ (.B(_08969_),
    .C(_11777_),
    .A(_08957_),
    .Y(_11804_));
 sg13g2_and2_1 _42457_ (.A(net5770),
    .B(_11804_),
    .X(_11805_));
 sg13g2_a22oi_1 _42458_ (.Y(_11806_),
    .B1(_11803_),
    .B2(_11805_),
    .A2(_08955_),
    .A1(net5732));
 sg13g2_nand2_1 _42459_ (.Y(_11807_),
    .A(net5470),
    .B(_11806_));
 sg13g2_xnor2_1 _42460_ (.Y(_11808_),
    .A(net5424),
    .B(_11806_));
 sg13g2_xor2_1 _42461_ (.B(_11808_),
    .A(_11802_),
    .X(_11809_));
 sg13g2_a21oi_1 _42462_ (.A1(net5567),
    .A2(_11806_),
    .Y(_11810_),
    .B1(net5932));
 sg13g2_o21ai_1 _42463_ (.B1(_11810_),
    .Y(_11811_),
    .A1(net5569),
    .A2(_11809_));
 sg13g2_a22oi_1 _42464_ (.Y(_11812_),
    .B1(_11779_),
    .B2(net5912),
    .A2(_08973_),
    .A1(net5997));
 sg13g2_and3_1 _42465_ (.X(_11813_),
    .A(net5296),
    .B(_11811_),
    .C(_11812_));
 sg13g2_o21ai_1 _42466_ (.B1(net6886),
    .Y(_11814_),
    .A1(net5296),
    .A2(_08973_));
 sg13g2_o21ai_1 _42467_ (.B1(_11801_),
    .Y(_00801_),
    .A1(_11813_),
    .A2(_11814_));
 sg13g2_or2_1 _42468_ (.X(_11815_),
    .B(_08961_),
    .A(net5771));
 sg13g2_nand2_1 _42469_ (.Y(_11816_),
    .A(_08956_),
    .B(_11803_));
 sg13g2_xnor2_1 _42470_ (.Y(_11817_),
    .A(_08963_),
    .B(_11816_));
 sg13g2_o21ai_1 _42471_ (.B1(_11815_),
    .Y(_11818_),
    .A1(net5732),
    .A2(_11817_));
 sg13g2_and2_1 _42472_ (.A(net5424),
    .B(_11818_),
    .X(_11819_));
 sg13g2_xnor2_1 _42473_ (.Y(_11820_),
    .A(net5469),
    .B(_11818_));
 sg13g2_a21o_1 _42474_ (.A2(_11806_),
    .A1(_11780_),
    .B1(net5469),
    .X(_11821_));
 sg13g2_nand2_1 _42475_ (.Y(_11822_),
    .A(_11795_),
    .B(_11821_));
 sg13g2_nand3_1 _42476_ (.B(_11820_),
    .C(_11822_),
    .A(_11807_),
    .Y(_11823_));
 sg13g2_a21o_1 _42477_ (.A2(_11822_),
    .A1(_11807_),
    .B1(_11820_),
    .X(_11824_));
 sg13g2_nand2_1 _42478_ (.Y(_11825_),
    .A(_11823_),
    .B(_11824_));
 sg13g2_a21oi_1 _42479_ (.A1(net5541),
    .A2(_11825_),
    .Y(_11826_),
    .B1(net5932));
 sg13g2_o21ai_1 _42480_ (.B1(_11826_),
    .Y(_11827_),
    .A1(net5541),
    .A2(_11818_));
 sg13g2_o21ai_1 _42481_ (.B1(_11827_),
    .Y(_11828_),
    .A1(net5881),
    .A2(_11806_));
 sg13g2_a21oi_1 _42482_ (.A1(net5997),
    .A2(_08968_),
    .Y(_11829_),
    .B1(_11828_));
 sg13g2_o21ai_1 _42483_ (.B1(net6886),
    .Y(_11830_),
    .A1(net5298),
    .A2(_08968_));
 sg13g2_a21oi_1 _42484_ (.A1(net5298),
    .A2(_11829_),
    .Y(_11831_),
    .B1(_11830_));
 sg13g2_a21o_1 _42485_ (.A2(net6469),
    .A1(net2814),
    .B1(_11831_),
    .X(_00802_));
 sg13g2_and2_1 _42486_ (.A(net5728),
    .B(_08945_),
    .X(_11832_));
 sg13g2_a21oi_1 _42487_ (.A1(net1067),
    .A2(_09652_),
    .Y(_11833_),
    .B1(_09657_));
 sg13g2_nor2_1 _42488_ (.A(_08977_),
    .B(_11833_),
    .Y(_11834_));
 sg13g2_o21ai_1 _42489_ (.B1(_08948_),
    .Y(_11835_),
    .A1(_08977_),
    .A2(_11833_));
 sg13g2_a21oi_1 _42490_ (.A1(_08947_),
    .A2(_11834_),
    .Y(_11836_),
    .B1(net5728));
 sg13g2_a21o_2 _42491_ (.A2(_11836_),
    .A1(_11835_),
    .B1(_11832_),
    .X(_11837_));
 sg13g2_nand2_1 _42492_ (.Y(_11838_),
    .A(net5425),
    .B(_11837_));
 sg13g2_xnor2_1 _42493_ (.Y(_11839_),
    .A(net5470),
    .B(_11837_));
 sg13g2_nand2b_1 _42494_ (.Y(_11840_),
    .B(_11823_),
    .A_N(_11819_));
 sg13g2_xnor2_1 _42495_ (.Y(_11841_),
    .A(_11839_),
    .B(_11840_));
 sg13g2_o21ai_1 _42496_ (.B1(net5965),
    .Y(_11842_),
    .A1(net5541),
    .A2(_11837_));
 sg13g2_a21oi_1 _42497_ (.A1(net5538),
    .A2(_11841_),
    .Y(_11843_),
    .B1(_11842_));
 sg13g2_a221oi_1 _42498_ (.B2(net5912),
    .C1(_11843_),
    .B1(_11818_),
    .A1(net5997),
    .Y(_11844_),
    .A2(_08955_));
 sg13g2_a21oi_1 _42499_ (.A1(net5296),
    .A2(_11844_),
    .Y(_11845_),
    .B1(net6860));
 sg13g2_o21ai_1 _42500_ (.B1(_11845_),
    .Y(_11846_),
    .A1(net5296),
    .A2(_08955_));
 sg13g2_o21ai_1 _42501_ (.B1(_11846_),
    .Y(_00803_),
    .A1(_18159_),
    .A2(net6508));
 sg13g2_a21oi_1 _42502_ (.A1(_08946_),
    .A2(_11835_),
    .Y(_11847_),
    .B1(_08941_));
 sg13g2_and3_1 _42503_ (.X(_11848_),
    .A(_08941_),
    .B(_08946_),
    .C(_11835_));
 sg13g2_nor3_1 _42504_ (.A(net5728),
    .B(_11847_),
    .C(_11848_),
    .Y(_11849_));
 sg13g2_a21oi_2 _42505_ (.B1(_11849_),
    .Y(_11850_),
    .A2(_08939_),
    .A1(net5728));
 sg13g2_or2_1 _42506_ (.X(_11851_),
    .B(_11850_),
    .A(net5470));
 sg13g2_xnor2_1 _42507_ (.Y(_11852_),
    .A(net5425),
    .B(_11850_));
 sg13g2_inv_1 _42508_ (.Y(_11853_),
    .A(_11852_));
 sg13g2_nand3b_1 _42509_ (.B(_11839_),
    .C(_11820_),
    .Y(_11854_),
    .A_N(_11821_));
 sg13g2_nand3b_1 _42510_ (.B(_11838_),
    .C(_11854_),
    .Y(_11855_),
    .A_N(_11819_));
 sg13g2_nand4_1 _42511_ (.B(_11808_),
    .C(_11820_),
    .A(_11782_),
    .Y(_11856_),
    .D(_11839_));
 sg13g2_a21oi_2 _42512_ (.B1(_11856_),
    .Y(_11857_),
    .A2(net1144),
    .A1(net1074));
 sg13g2_o21ai_1 _42513_ (.B1(_11852_),
    .Y(_11858_),
    .A1(_11855_),
    .A2(_11857_));
 sg13g2_or3_1 _42514_ (.A(_11852_),
    .B(_11855_),
    .C(_11857_),
    .X(_11859_));
 sg13g2_a21oi_1 _42515_ (.A1(_11858_),
    .A2(_11859_),
    .Y(_11860_),
    .B1(net5567));
 sg13g2_a21oi_1 _42516_ (.A1(net5567),
    .A2(_11850_),
    .Y(_11861_),
    .B1(_11860_));
 sg13g2_a22oi_1 _42517_ (.Y(_11862_),
    .B1(_11861_),
    .B2(net5965),
    .A2(_11837_),
    .A1(net5912));
 sg13g2_o21ai_1 _42518_ (.B1(_11862_),
    .Y(_11863_),
    .A1(net6007),
    .A2(_08961_));
 sg13g2_a21oi_1 _42519_ (.A1(net5321),
    .A2(net5317),
    .Y(_11864_),
    .B1(_11863_));
 sg13g2_nor2b_1 _42520_ (.A(net5298),
    .B_N(_08961_),
    .Y(_11865_));
 sg13g2_nor3_1 _42521_ (.A(net6860),
    .B(_11864_),
    .C(_11865_),
    .Y(_11866_));
 sg13g2_a21o_1 _42522_ (.A2(net6470),
    .A1(net3199),
    .B1(_11866_),
    .X(_00804_));
 sg13g2_nand2_1 _42523_ (.Y(_11867_),
    .A(_11851_),
    .B(_11858_));
 sg13g2_nor2_1 _42524_ (.A(net5771),
    .B(_08928_),
    .Y(_11868_));
 sg13g2_a21oi_1 _42525_ (.A1(_08978_),
    .A2(_11835_),
    .Y(_11869_),
    .B1(_08940_));
 sg13g2_xnor2_1 _42526_ (.Y(_11870_),
    .A(_08931_),
    .B(_11869_));
 sg13g2_a21oi_2 _42527_ (.B1(_11868_),
    .Y(_11871_),
    .A2(_11870_),
    .A1(net5771));
 sg13g2_nand2_1 _42528_ (.Y(_11872_),
    .A(net5425),
    .B(_11871_));
 sg13g2_nand2b_1 _42529_ (.Y(_11873_),
    .B(net5470),
    .A_N(_11871_));
 sg13g2_nand2_1 _42530_ (.Y(_11874_),
    .A(_11872_),
    .B(_11873_));
 sg13g2_xor2_1 _42531_ (.B(_11874_),
    .A(_11867_),
    .X(_11875_));
 sg13g2_nor2_1 _42532_ (.A(net5537),
    .B(_11871_),
    .Y(_11876_));
 sg13g2_a21oi_1 _42533_ (.A1(net5537),
    .A2(_11875_),
    .Y(_11877_),
    .B1(_11876_));
 sg13g2_nor2_1 _42534_ (.A(net5881),
    .B(_11850_),
    .Y(_11878_));
 sg13g2_a221oi_1 _42535_ (.B2(net5965),
    .C1(_11878_),
    .B1(_11877_),
    .A1(net5997),
    .Y(_11879_),
    .A2(_08945_));
 sg13g2_o21ai_1 _42536_ (.B1(net6886),
    .Y(_11880_),
    .A1(net5294),
    .A2(_08945_));
 sg13g2_a21oi_1 _42537_ (.A1(net5294),
    .A2(_11879_),
    .Y(_11881_),
    .B1(_11880_));
 sg13g2_a21o_1 _42538_ (.A2(net6469),
    .A1(net3340),
    .B1(_11881_),
    .X(_00805_));
 sg13g2_nand2_1 _42539_ (.Y(_11882_),
    .A(net5728),
    .B(_08934_));
 sg13g2_a21oi_1 _42540_ (.A1(_08931_),
    .A2(_11869_),
    .Y(_11883_),
    .B1(_08929_));
 sg13g2_xnor2_1 _42541_ (.Y(_11884_),
    .A(_08936_),
    .B(_11883_));
 sg13g2_o21ai_1 _42542_ (.B1(_11882_),
    .Y(_11885_),
    .A1(net5728),
    .A2(_11884_));
 sg13g2_nor2_1 _42543_ (.A(net5538),
    .B(_11885_),
    .Y(_11886_));
 sg13g2_nand2_1 _42544_ (.Y(_11887_),
    .A(net5425),
    .B(_11885_));
 sg13g2_xnor2_1 _42545_ (.Y(_11888_),
    .A(net5470),
    .B(_11885_));
 sg13g2_and2_1 _42546_ (.A(_11851_),
    .B(_11872_),
    .X(_11889_));
 sg13g2_nand2_1 _42547_ (.Y(_11890_),
    .A(_11858_),
    .B(_11889_));
 sg13g2_nand3_1 _42548_ (.B(_11888_),
    .C(_11890_),
    .A(_11873_),
    .Y(_11891_));
 sg13g2_a21o_1 _42549_ (.A2(_11890_),
    .A1(_11873_),
    .B1(_11888_),
    .X(_11892_));
 sg13g2_nand2_1 _42550_ (.Y(_11893_),
    .A(_11891_),
    .B(_11892_));
 sg13g2_a21oi_1 _42551_ (.A1(net5538),
    .A2(_11893_),
    .Y(_11894_),
    .B1(_11886_));
 sg13g2_a22oi_1 _42552_ (.Y(_11895_),
    .B1(_11894_),
    .B2(net5230),
    .A2(_11871_),
    .A1(net5218));
 sg13g2_a22oi_1 _42553_ (.Y(_11896_),
    .B1(net5107),
    .B2(_08939_),
    .A2(net6469),
    .A1(net3239));
 sg13g2_o21ai_1 _42554_ (.B1(_11896_),
    .Y(_00806_),
    .A1(net6860),
    .A2(_11895_));
 sg13g2_and2_1 _42555_ (.A(net5728),
    .B(_08915_),
    .X(_11897_));
 sg13g2_a21oi_2 _42556_ (.B1(_09658_),
    .Y(_11898_),
    .A2(_09652_),
    .A1(net1067));
 sg13g2_o21ai_1 _42557_ (.B1(_08918_),
    .Y(_11899_),
    .A1(_08981_),
    .A2(_11898_));
 sg13g2_nor3_1 _42558_ (.A(_08918_),
    .B(_08981_),
    .C(_11898_),
    .Y(_11900_));
 sg13g2_nor2_1 _42559_ (.A(net5728),
    .B(_11900_),
    .Y(_11901_));
 sg13g2_a21o_2 _42560_ (.A2(_11901_),
    .A1(_11899_),
    .B1(_11897_),
    .X(_11902_));
 sg13g2_xnor2_1 _42561_ (.Y(_11903_),
    .A(net5470),
    .B(_11902_));
 sg13g2_and2_1 _42562_ (.A(_11887_),
    .B(_11891_),
    .X(_11904_));
 sg13g2_xor2_1 _42563_ (.B(_11904_),
    .A(_11903_),
    .X(_11905_));
 sg13g2_o21ai_1 _42564_ (.B1(net5966),
    .Y(_11906_),
    .A1(net5538),
    .A2(_11902_));
 sg13g2_a21oi_1 _42565_ (.A1(net5538),
    .A2(_11905_),
    .Y(_11907_),
    .B1(_11906_));
 sg13g2_a221oi_1 _42566_ (.B2(net5912),
    .C1(_11907_),
    .B1(_11885_),
    .A1(net5997),
    .Y(_11908_),
    .A2(_08928_));
 sg13g2_o21ai_1 _42567_ (.B1(net6886),
    .Y(_11909_),
    .A1(net5297),
    .A2(_08928_));
 sg13g2_a21oi_1 _42568_ (.A1(net5294),
    .A2(_11908_),
    .Y(_11910_),
    .B1(_11909_));
 sg13g2_a21oi_1 _42569_ (.A1(net1867),
    .A2(net6469),
    .Y(_11911_),
    .B1(_11910_));
 sg13g2_inv_1 _42570_ (.Y(_00807_),
    .A(_11911_));
 sg13g2_nand2_1 _42571_ (.Y(_11912_),
    .A(net2804),
    .B(net6469));
 sg13g2_nand2_1 _42572_ (.Y(_11913_),
    .A(_08916_),
    .B(_11899_));
 sg13g2_xor2_1 _42573_ (.B(_11913_),
    .A(_08911_),
    .X(_11914_));
 sg13g2_nor2_1 _42574_ (.A(net5735),
    .B(_11914_),
    .Y(_11915_));
 sg13g2_a21oi_2 _42575_ (.B1(_11915_),
    .Y(_11916_),
    .A2(_08908_),
    .A1(net5729));
 sg13g2_nor2_1 _42576_ (.A(net5473),
    .B(_11916_),
    .Y(_11917_));
 sg13g2_xnor2_1 _42577_ (.Y(_11918_),
    .A(net5425),
    .B(_11916_));
 sg13g2_nand2_1 _42578_ (.Y(_11919_),
    .A(_11888_),
    .B(_11903_));
 sg13g2_nor3_1 _42579_ (.A(_11853_),
    .B(_11874_),
    .C(_11919_),
    .Y(_11920_));
 sg13g2_o21ai_1 _42580_ (.B1(_11887_),
    .Y(_11921_),
    .A1(_11889_),
    .A2(_11919_));
 sg13g2_a221oi_1 _42581_ (.B2(_11855_),
    .C1(_11921_),
    .B1(_11920_),
    .A1(net5425),
    .Y(_11922_),
    .A2(_11902_));
 sg13g2_nand2b_1 _42582_ (.Y(_11923_),
    .B(_11920_),
    .A_N(_11856_));
 sg13g2_nand2b_1 _42583_ (.Y(_11924_),
    .B(_11794_),
    .A_N(_11923_));
 sg13g2_nand2_1 _42584_ (.Y(_11925_),
    .A(_11922_),
    .B(_11924_));
 sg13g2_and2_1 _42585_ (.A(_11918_),
    .B(_11925_),
    .X(_11926_));
 sg13g2_xnor2_1 _42586_ (.Y(_11927_),
    .A(_11918_),
    .B(_11925_));
 sg13g2_nand2_1 _42587_ (.Y(_11928_),
    .A(net5569),
    .B(_11916_));
 sg13g2_a21oi_1 _42588_ (.A1(net5537),
    .A2(_11927_),
    .Y(_11929_),
    .B1(net5932));
 sg13g2_a22oi_1 _42589_ (.Y(_11930_),
    .B1(_11902_),
    .B2(net5912),
    .A2(_08934_),
    .A1(net5998));
 sg13g2_nand2_1 _42590_ (.Y(_11931_),
    .A(net5297),
    .B(_11930_));
 sg13g2_a21oi_1 _42591_ (.A1(_11928_),
    .A2(_11929_),
    .Y(_11932_),
    .B1(_11931_));
 sg13g2_o21ai_1 _42592_ (.B1(net6886),
    .Y(_11933_),
    .A1(net5294),
    .A2(_08934_));
 sg13g2_o21ai_1 _42593_ (.B1(_11912_),
    .Y(_00808_),
    .A1(_11932_),
    .A2(_11933_));
 sg13g2_a21oi_1 _42594_ (.A1(_08983_),
    .A2(_11899_),
    .Y(_11934_),
    .B1(_08910_));
 sg13g2_xnor2_1 _42595_ (.Y(_11935_),
    .A(_08900_),
    .B(_11934_));
 sg13g2_nor2_1 _42596_ (.A(net5768),
    .B(_08897_),
    .Y(_11936_));
 sg13g2_a21o_1 _42597_ (.A2(_11935_),
    .A1(net5768),
    .B1(_11936_),
    .X(_11937_));
 sg13g2_a21oi_1 _42598_ (.A1(net5768),
    .A2(_11935_),
    .Y(_11938_),
    .B1(_11936_));
 sg13g2_nand2_1 _42599_ (.Y(_11939_),
    .A(net5471),
    .B(_11938_));
 sg13g2_xnor2_1 _42600_ (.Y(_11940_),
    .A(net5425),
    .B(_11937_));
 sg13g2_inv_1 _42601_ (.Y(_11941_),
    .A(_11940_));
 sg13g2_o21ai_1 _42602_ (.B1(_11940_),
    .Y(_11942_),
    .A1(_11917_),
    .A2(_11926_));
 sg13g2_nor3_1 _42603_ (.A(_11917_),
    .B(_11926_),
    .C(_11940_),
    .Y(_11943_));
 sg13g2_nor2_1 _42604_ (.A(net5567),
    .B(_11943_),
    .Y(_11944_));
 sg13g2_a22oi_1 _42605_ (.Y(_11945_),
    .B1(_11942_),
    .B2(_11944_),
    .A2(_11938_),
    .A1(net5567));
 sg13g2_nor2_1 _42606_ (.A(net5883),
    .B(_11916_),
    .Y(_11946_));
 sg13g2_a221oi_1 _42607_ (.B2(net5965),
    .C1(_11946_),
    .B1(_11945_),
    .A1(net5998),
    .Y(_11947_),
    .A2(_08915_));
 sg13g2_a21oi_1 _42608_ (.A1(net5297),
    .A2(_11947_),
    .Y(_11948_),
    .B1(net6860));
 sg13g2_o21ai_1 _42609_ (.B1(_11948_),
    .Y(_11949_),
    .A1(net5303),
    .A2(_08915_));
 sg13g2_o21ai_1 _42610_ (.B1(_11949_),
    .Y(_00809_),
    .A1(_18157_),
    .A2(net6508));
 sg13g2_nand2_1 _42611_ (.Y(_11950_),
    .A(net3260),
    .B(net6469));
 sg13g2_or2_1 _42612_ (.X(_11951_),
    .B(_08904_),
    .A(net5771));
 sg13g2_a21oi_1 _42613_ (.A1(_08901_),
    .A2(_11934_),
    .Y(_11952_),
    .B1(_08899_));
 sg13g2_xnor2_1 _42614_ (.Y(_11953_),
    .A(_08905_),
    .B(_11952_));
 sg13g2_o21ai_1 _42615_ (.B1(_11951_),
    .Y(_11954_),
    .A1(net5734),
    .A2(_11953_));
 sg13g2_nand2_1 _42616_ (.Y(_11955_),
    .A(net5426),
    .B(_11954_));
 sg13g2_xnor2_1 _42617_ (.Y(_11956_),
    .A(net5470),
    .B(_11954_));
 sg13g2_inv_1 _42618_ (.Y(_11957_),
    .A(_11956_));
 sg13g2_a21oi_1 _42619_ (.A1(_11916_),
    .A2(_11938_),
    .Y(_11958_),
    .B1(net5471));
 sg13g2_o21ai_1 _42620_ (.B1(_11939_),
    .Y(_11959_),
    .A1(_11926_),
    .A2(_11958_));
 sg13g2_xnor2_1 _42621_ (.Y(_11960_),
    .A(_11957_),
    .B(_11959_));
 sg13g2_nand2_1 _42622_ (.Y(_11961_),
    .A(net5541),
    .B(_11960_));
 sg13g2_o21ai_1 _42623_ (.B1(_11961_),
    .Y(_11962_),
    .A1(net5544),
    .A2(_11954_));
 sg13g2_nor2_1 _42624_ (.A(net5153),
    .B(_11962_),
    .Y(_11963_));
 sg13g2_a221oi_1 _42625_ (.B2(net5220),
    .C1(_11963_),
    .B1(_11937_),
    .A1(net5167),
    .Y(_11964_),
    .A2(_08908_));
 sg13g2_o21ai_1 _42626_ (.B1(_11950_),
    .Y(_00810_),
    .A1(net6860),
    .A2(_11964_));
 sg13g2_nor2_1 _42627_ (.A(net5768),
    .B(_08883_),
    .Y(_11965_));
 sg13g2_o21ai_1 _42628_ (.B1(_08919_),
    .Y(_11966_),
    .A1(_08981_),
    .A2(_11898_));
 sg13g2_a21oi_1 _42629_ (.A1(_08986_),
    .A2(_11966_),
    .Y(_11967_),
    .B1(_08885_));
 sg13g2_and3_1 _42630_ (.X(_11968_),
    .A(_08885_),
    .B(_08986_),
    .C(_11966_));
 sg13g2_nor3_1 _42631_ (.A(net5734),
    .B(_11967_),
    .C(_11968_),
    .Y(_11969_));
 sg13g2_nor2_1 _42632_ (.A(_11965_),
    .B(_11969_),
    .Y(_11970_));
 sg13g2_nor2_1 _42633_ (.A(net5471),
    .B(_11970_),
    .Y(_11971_));
 sg13g2_xnor2_1 _42634_ (.Y(_11972_),
    .A(net5426),
    .B(_11970_));
 sg13g2_o21ai_1 _42635_ (.B1(_11955_),
    .Y(_11973_),
    .A1(_11957_),
    .A2(_11959_));
 sg13g2_xor2_1 _42636_ (.B(_11973_),
    .A(_11972_),
    .X(_11974_));
 sg13g2_a21oi_1 _42637_ (.A1(net5568),
    .A2(_11970_),
    .Y(_11975_),
    .B1(net5933));
 sg13g2_o21ai_1 _42638_ (.B1(_11975_),
    .Y(_11976_),
    .A1(net5567),
    .A2(_11974_));
 sg13g2_a22oi_1 _42639_ (.Y(_11977_),
    .B1(_11954_),
    .B2(net5912),
    .A2(_08898_),
    .A1(net5998));
 sg13g2_nand3_1 _42640_ (.B(_11976_),
    .C(_11977_),
    .A(net5298),
    .Y(_11978_));
 sg13g2_nor2_1 _42641_ (.A(net5298),
    .B(_08898_),
    .Y(_11979_));
 sg13g2_nor2_1 _42642_ (.A(net6860),
    .B(_11979_),
    .Y(_11980_));
 sg13g2_a22oi_1 _42643_ (.Y(_11981_),
    .B1(_11978_),
    .B2(_11980_),
    .A2(net6472),
    .A1(net3477));
 sg13g2_inv_1 _42644_ (.Y(_00811_),
    .A(_11981_));
 sg13g2_nor2b_1 _42645_ (.A(net5294),
    .B_N(_08904_),
    .Y(_11982_));
 sg13g2_nor2_1 _42646_ (.A(_08884_),
    .B(_11967_),
    .Y(_11983_));
 sg13g2_xor2_1 _42647_ (.B(_11983_),
    .A(_08892_),
    .X(_11984_));
 sg13g2_nand2_1 _42648_ (.Y(_11985_),
    .A(net5734),
    .B(_08888_));
 sg13g2_o21ai_1 _42649_ (.B1(_11985_),
    .Y(_11986_),
    .A1(net5734),
    .A2(_11984_));
 sg13g2_nand2_1 _42650_ (.Y(_11987_),
    .A(net5426),
    .B(_11986_));
 sg13g2_xnor2_1 _42651_ (.Y(_11988_),
    .A(net5471),
    .B(_11986_));
 sg13g2_nand3_1 _42652_ (.B(_11958_),
    .C(_11972_),
    .A(_11956_),
    .Y(_11989_));
 sg13g2_nand2_1 _42653_ (.Y(_11990_),
    .A(_11955_),
    .B(_11989_));
 sg13g2_nor2_1 _42654_ (.A(_11971_),
    .B(_11990_),
    .Y(_11991_));
 sg13g2_or2_1 _42655_ (.X(_11992_),
    .B(_11990_),
    .A(_11971_));
 sg13g2_nand4_1 _42656_ (.B(_11941_),
    .C(_11956_),
    .A(_11918_),
    .Y(_11993_),
    .D(_11972_));
 sg13g2_a21oi_1 _42657_ (.A1(_11922_),
    .A2(_11924_),
    .Y(_11994_),
    .B1(_11993_));
 sg13g2_nor2_1 _42658_ (.A(_11992_),
    .B(_11994_),
    .Y(_11995_));
 sg13g2_o21ai_1 _42659_ (.B1(_11988_),
    .Y(_11996_),
    .A1(_11992_),
    .A2(_11994_));
 sg13g2_xor2_1 _42660_ (.B(_11995_),
    .A(_11988_),
    .X(_11997_));
 sg13g2_o21ai_1 _42661_ (.B1(net5965),
    .Y(_11998_),
    .A1(net5541),
    .A2(_11986_));
 sg13g2_a21o_1 _42662_ (.A2(_11997_),
    .A1(net5541),
    .B1(_11998_),
    .X(_11999_));
 sg13g2_or2_1 _42663_ (.X(_12000_),
    .B(_08904_),
    .A(net6007));
 sg13g2_o21ai_1 _42664_ (.B1(net5914),
    .Y(_12001_),
    .A1(_11965_),
    .A2(_11969_));
 sg13g2_nand4_1 _42665_ (.B(_11999_),
    .C(_12000_),
    .A(net5297),
    .Y(_12002_),
    .D(_12001_));
 sg13g2_nor2_1 _42666_ (.A(net6860),
    .B(_11982_),
    .Y(_12003_));
 sg13g2_a22oi_1 _42667_ (.Y(_12004_),
    .B1(_12002_),
    .B2(_12003_),
    .A2(net6470),
    .A1(net3393));
 sg13g2_inv_1 _42668_ (.Y(_00812_),
    .A(_12004_));
 sg13g2_nor2_1 _42669_ (.A(net5768),
    .B(_08868_),
    .Y(_12005_));
 sg13g2_o21ai_1 _42670_ (.B1(_08889_),
    .Y(_12006_),
    .A1(_08891_),
    .A2(_11983_));
 sg13g2_xnor2_1 _42671_ (.Y(_12007_),
    .A(_08870_),
    .B(_12006_));
 sg13g2_a21oi_2 _42672_ (.B1(_12005_),
    .Y(_12008_),
    .A2(_12007_),
    .A1(net5768));
 sg13g2_nor2_1 _42673_ (.A(net5426),
    .B(_12008_),
    .Y(_12009_));
 sg13g2_xnor2_1 _42674_ (.Y(_12010_),
    .A(net5471),
    .B(_12008_));
 sg13g2_nand2_1 _42675_ (.Y(_12011_),
    .A(_11987_),
    .B(_11996_));
 sg13g2_xnor2_1 _42676_ (.Y(_12012_),
    .A(_12010_),
    .B(_12011_));
 sg13g2_o21ai_1 _42677_ (.B1(net5965),
    .Y(_12013_),
    .A1(net5544),
    .A2(_12008_));
 sg13g2_a21oi_1 _42678_ (.A1(net5544),
    .A2(_12012_),
    .Y(_12014_),
    .B1(_12013_));
 sg13g2_nand2b_1 _42679_ (.Y(_12015_),
    .B(net5997),
    .A_N(_08883_));
 sg13g2_a21oi_1 _42680_ (.A1(net5912),
    .A2(_11986_),
    .Y(_12016_),
    .B1(_12014_));
 sg13g2_nand3_1 _42681_ (.B(_12015_),
    .C(_12016_),
    .A(net5297),
    .Y(_12017_));
 sg13g2_nand3_1 _42682_ (.B(net5318),
    .C(_08883_),
    .A(net5322),
    .Y(_12018_));
 sg13g2_nand3_1 _42683_ (.B(_12017_),
    .C(_12018_),
    .A(net6886),
    .Y(_12019_));
 sg13g2_o21ai_1 _42684_ (.B1(_12019_),
    .Y(_00813_),
    .A1(_18155_),
    .A2(net6508));
 sg13g2_and2_1 _42685_ (.A(net5734),
    .B(_08876_),
    .X(_12020_));
 sg13g2_a21oi_1 _42686_ (.A1(_08870_),
    .A2(_12006_),
    .Y(_12021_),
    .B1(_08869_));
 sg13g2_xnor2_1 _42687_ (.Y(_12022_),
    .A(_08878_),
    .B(_12021_));
 sg13g2_a21oi_2 _42688_ (.B1(_12020_),
    .Y(_12023_),
    .A2(_12022_),
    .A1(net5768));
 sg13g2_nor2_1 _42689_ (.A(net5471),
    .B(_12023_),
    .Y(_12024_));
 sg13g2_xnor2_1 _42690_ (.Y(_12025_),
    .A(net5426),
    .B(_12023_));
 sg13g2_o21ai_1 _42691_ (.B1(net5426),
    .Y(_12026_),
    .A1(_11986_),
    .A2(_12008_));
 sg13g2_a21oi_1 _42692_ (.A1(_11996_),
    .A2(_12026_),
    .Y(_12027_),
    .B1(_12009_));
 sg13g2_xor2_1 _42693_ (.B(_12027_),
    .A(_12025_),
    .X(_12028_));
 sg13g2_o21ai_1 _42694_ (.B1(net5965),
    .Y(_12029_),
    .A1(net5567),
    .A2(_12028_));
 sg13g2_a21oi_1 _42695_ (.A1(net5567),
    .A2(_12023_),
    .Y(_12030_),
    .B1(_12029_));
 sg13g2_a221oi_1 _42696_ (.B2(net5912),
    .C1(_12030_),
    .B1(_12008_),
    .A1(net5997),
    .Y(_12031_),
    .A2(_08888_));
 sg13g2_a21oi_1 _42697_ (.A1(net5297),
    .A2(_12031_),
    .Y(_12032_),
    .B1(net6861));
 sg13g2_o21ai_1 _42698_ (.B1(_12032_),
    .Y(_12033_),
    .A1(net5297),
    .A2(_08888_));
 sg13g2_o21ai_1 _42699_ (.B1(_12033_),
    .Y(_00814_),
    .A1(_18154_),
    .A2(net6506));
 sg13g2_nand2_1 _42700_ (.Y(_12034_),
    .A(net5729),
    .B(_09101_));
 sg13g2_a21oi_2 _42701_ (.B1(_09659_),
    .Y(_12035_),
    .A2(_09652_),
    .A1(net1067));
 sg13g2_nor2_1 _42702_ (.A(_08990_),
    .B(_12035_),
    .Y(_12036_));
 sg13g2_o21ai_1 _42703_ (.B1(_09103_),
    .Y(_12037_),
    .A1(_08990_),
    .A2(_12035_));
 sg13g2_xor2_1 _42704_ (.B(_12036_),
    .A(_09103_),
    .X(_12038_));
 sg13g2_o21ai_1 _42705_ (.B1(_12034_),
    .Y(_12039_),
    .A1(net5732),
    .A2(_12038_));
 sg13g2_nand2_1 _42706_ (.Y(_12040_),
    .A(net5425),
    .B(_12039_));
 sg13g2_xnor2_1 _42707_ (.Y(_12041_),
    .A(net5470),
    .B(_12039_));
 sg13g2_a21oi_1 _42708_ (.A1(_12025_),
    .A2(_12027_),
    .Y(_12042_),
    .B1(_12024_));
 sg13g2_xor2_1 _42709_ (.B(_12042_),
    .A(_12041_),
    .X(_12043_));
 sg13g2_nor2_1 _42710_ (.A(net5541),
    .B(_12039_),
    .Y(_12044_));
 sg13g2_a21oi_1 _42711_ (.A1(net5541),
    .A2(_12043_),
    .Y(_12045_),
    .B1(_12044_));
 sg13g2_nor2_1 _42712_ (.A(net5883),
    .B(_12023_),
    .Y(_12046_));
 sg13g2_a221oi_1 _42713_ (.B2(net5965),
    .C1(_12046_),
    .B1(_12045_),
    .A1(net5997),
    .Y(_12047_),
    .A2(_08868_));
 sg13g2_o21ai_1 _42714_ (.B1(net6886),
    .Y(_12048_),
    .A1(net5297),
    .A2(_08868_));
 sg13g2_a21oi_1 _42715_ (.A1(net5298),
    .A2(_12047_),
    .Y(_12049_),
    .B1(_12048_));
 sg13g2_a21o_1 _42716_ (.A2(net6469),
    .A1(net3274),
    .B1(_12049_),
    .X(_00815_));
 sg13g2_nor2_1 _42717_ (.A(net5771),
    .B(_09096_),
    .Y(_12050_));
 sg13g2_nand2_1 _42718_ (.Y(_12051_),
    .A(_09102_),
    .B(_12037_));
 sg13g2_xor2_1 _42719_ (.B(_12051_),
    .A(_09099_),
    .X(_12052_));
 sg13g2_a21oi_2 _42720_ (.B1(_12050_),
    .Y(_12053_),
    .A2(_12052_),
    .A1(net5771));
 sg13g2_nor2_1 _42721_ (.A(net5537),
    .B(_12053_),
    .Y(_12054_));
 sg13g2_nand2_1 _42722_ (.Y(_12055_),
    .A(net5430),
    .B(_12053_));
 sg13g2_xnor2_1 _42723_ (.Y(_12056_),
    .A(net5430),
    .B(_12053_));
 sg13g2_nand2_1 _42724_ (.Y(_12057_),
    .A(_12025_),
    .B(_12041_));
 sg13g2_nand2_1 _42725_ (.Y(_12058_),
    .A(_11988_),
    .B(_12010_));
 sg13g2_nor4_1 _42726_ (.A(_11922_),
    .B(_11993_),
    .C(_12057_),
    .D(_12058_),
    .Y(_12059_));
 sg13g2_nor3_1 _42727_ (.A(_11991_),
    .B(_12057_),
    .C(_12058_),
    .Y(_12060_));
 sg13g2_o21ai_1 _42728_ (.B1(_12040_),
    .Y(_12061_),
    .A1(_12026_),
    .A2(_12057_));
 sg13g2_or4_1 _42729_ (.A(_12024_),
    .B(_12059_),
    .C(_12060_),
    .D(_12061_),
    .X(_12062_));
 sg13g2_or4_1 _42730_ (.A(_11923_),
    .B(_11993_),
    .C(_12057_),
    .D(_12058_),
    .X(_12063_));
 sg13g2_inv_4 _42731_ (.A(_12063_),
    .Y(_12064_));
 sg13g2_a21oi_2 _42732_ (.B1(_12062_),
    .Y(_12065_),
    .A2(_12064_),
    .A1(_11794_));
 sg13g2_or2_1 _42733_ (.X(_12066_),
    .B(_12065_),
    .A(_12056_));
 sg13g2_xnor2_1 _42734_ (.Y(_12067_),
    .A(_12056_),
    .B(_12065_));
 sg13g2_a21oi_1 _42735_ (.A1(net5537),
    .A2(_12067_),
    .Y(_12068_),
    .B1(_12054_));
 sg13g2_a22oi_1 _42736_ (.Y(_12069_),
    .B1(_12068_),
    .B2(net5230),
    .A2(_12039_),
    .A1(net5218));
 sg13g2_a22oi_1 _42737_ (.Y(_12070_),
    .B1(net5107),
    .B2(_08876_),
    .A2(net6469),
    .A1(net2325));
 sg13g2_o21ai_1 _42738_ (.B1(_12070_),
    .Y(_00816_),
    .A1(net6860),
    .A2(_12069_));
 sg13g2_nand2_1 _42739_ (.Y(_12071_),
    .A(_12055_),
    .B(_12066_));
 sg13g2_nand2b_1 _42740_ (.Y(_12072_),
    .B(net5729),
    .A_N(_09090_));
 sg13g2_a21oi_1 _42741_ (.A1(_09117_),
    .A2(_12037_),
    .Y(_12073_),
    .B1(_09098_));
 sg13g2_xnor2_1 _42742_ (.Y(_12074_),
    .A(_09092_),
    .B(_12073_));
 sg13g2_o21ai_1 _42743_ (.B1(_12072_),
    .Y(_12075_),
    .A1(net5729),
    .A2(_12074_));
 sg13g2_or2_1 _42744_ (.X(_12076_),
    .B(_12075_),
    .A(net5430));
 sg13g2_xnor2_1 _42745_ (.Y(_12077_),
    .A(net5430),
    .B(_12075_));
 sg13g2_xor2_1 _42746_ (.B(_12077_),
    .A(_12071_),
    .X(_12078_));
 sg13g2_o21ai_1 _42747_ (.B1(net5964),
    .Y(_12079_),
    .A1(net5537),
    .A2(_12075_));
 sg13g2_a21oi_1 _42748_ (.A1(net5537),
    .A2(_12078_),
    .Y(_12080_),
    .B1(_12079_));
 sg13g2_a221oi_1 _42749_ (.B2(net5910),
    .C1(_12080_),
    .B1(_12053_),
    .A1(net5995),
    .Y(_12081_),
    .A2(_09101_));
 sg13g2_a21oi_1 _42750_ (.A1(net5294),
    .A2(_12081_),
    .Y(_12082_),
    .B1(net6862));
 sg13g2_o21ai_1 _42751_ (.B1(_12082_),
    .Y(_12083_),
    .A1(net5293),
    .A2(_09101_));
 sg13g2_o21ai_1 _42752_ (.B1(_12083_),
    .Y(_00817_),
    .A1(_18153_),
    .A2(net6508));
 sg13g2_a21oi_1 _42753_ (.A1(_09092_),
    .A2(_12073_),
    .Y(_12084_),
    .B1(_09091_));
 sg13g2_xor2_1 _42754_ (.B(_12084_),
    .A(_09084_),
    .X(_12085_));
 sg13g2_nor2_1 _42755_ (.A(net5729),
    .B(_12085_),
    .Y(_12086_));
 sg13g2_a21oi_2 _42756_ (.B1(_12086_),
    .Y(_12087_),
    .A2(_09083_),
    .A1(net5729));
 sg13g2_nor2_1 _42757_ (.A(net5473),
    .B(_12087_),
    .Y(_12088_));
 sg13g2_xnor2_1 _42758_ (.Y(_12089_),
    .A(net5430),
    .B(_12087_));
 sg13g2_o21ai_1 _42759_ (.B1(net5430),
    .Y(_12090_),
    .A1(_12053_),
    .A2(_12075_));
 sg13g2_inv_1 _42760_ (.Y(_12091_),
    .A(_12090_));
 sg13g2_nand2_1 _42761_ (.Y(_12092_),
    .A(_12066_),
    .B(_12090_));
 sg13g2_nand3_1 _42762_ (.B(_12089_),
    .C(_12092_),
    .A(_12076_),
    .Y(_12093_));
 sg13g2_a21o_1 _42763_ (.A2(_12092_),
    .A1(_12076_),
    .B1(_12089_),
    .X(_12094_));
 sg13g2_and2_1 _42764_ (.A(_12093_),
    .B(_12094_),
    .X(_12095_));
 sg13g2_o21ai_1 _42765_ (.B1(net5964),
    .Y(_12096_),
    .A1(net5569),
    .A2(_12095_));
 sg13g2_a21oi_1 _42766_ (.A1(net5569),
    .A2(_12087_),
    .Y(_12097_),
    .B1(_12096_));
 sg13g2_a221oi_1 _42767_ (.B2(net5910),
    .C1(_12097_),
    .B1(_12075_),
    .A1(net5995),
    .Y(_12098_),
    .A2(_09096_));
 sg13g2_a21oi_1 _42768_ (.A1(net5293),
    .A2(_12098_),
    .Y(_12099_),
    .B1(net6862));
 sg13g2_o21ai_1 _42769_ (.B1(_12099_),
    .Y(_12100_),
    .A1(net5293),
    .A2(_09096_));
 sg13g2_o21ai_1 _42770_ (.B1(_12100_),
    .Y(_00818_),
    .A1(_18152_),
    .A2(net6508));
 sg13g2_o21ai_1 _42771_ (.B1(_09105_),
    .Y(_12101_),
    .A1(_08990_),
    .A2(_12035_));
 sg13g2_a21oi_1 _42772_ (.A1(_09119_),
    .A2(_12101_),
    .Y(_12102_),
    .B1(_09077_));
 sg13g2_and3_1 _42773_ (.X(_12103_),
    .A(_09077_),
    .B(_09119_),
    .C(_12101_));
 sg13g2_nor3_1 _42774_ (.A(net5729),
    .B(_12102_),
    .C(_12103_),
    .Y(_12104_));
 sg13g2_a21oi_2 _42775_ (.B1(_12104_),
    .Y(_12105_),
    .A2(_09076_),
    .A1(net5729));
 sg13g2_xnor2_1 _42776_ (.Y(_12106_),
    .A(net5430),
    .B(_12105_));
 sg13g2_nor2b_1 _42777_ (.A(_12088_),
    .B_N(_12093_),
    .Y(_12107_));
 sg13g2_xnor2_1 _42778_ (.Y(_12108_),
    .A(_12106_),
    .B(_12107_));
 sg13g2_a21oi_1 _42779_ (.A1(net5569),
    .A2(_12105_),
    .Y(_12109_),
    .B1(net5932));
 sg13g2_o21ai_1 _42780_ (.B1(_12109_),
    .Y(_12110_),
    .A1(net5569),
    .A2(_12108_));
 sg13g2_nand2b_1 _42781_ (.Y(_12111_),
    .B(net5995),
    .A_N(_09090_));
 sg13g2_nand2b_1 _42782_ (.Y(_12112_),
    .B(net5910),
    .A_N(_12087_));
 sg13g2_nand4_1 _42783_ (.B(_12110_),
    .C(_12111_),
    .A(net5293),
    .Y(_12113_),
    .D(_12112_));
 sg13g2_nor2b_1 _42784_ (.A(net5294),
    .B_N(_09090_),
    .Y(_12114_));
 sg13g2_nor2_1 _42785_ (.A(net6863),
    .B(_12114_),
    .Y(_12115_));
 sg13g2_a22oi_1 _42786_ (.Y(_12116_),
    .B1(_12113_),
    .B2(_12115_),
    .A2(net6459),
    .A1(net2746));
 sg13g2_inv_1 _42787_ (.Y(_00819_),
    .A(_12116_));
 sg13g2_a21oi_1 _42788_ (.A1(net5671),
    .A2(_09076_),
    .Y(_12117_),
    .B1(_12102_));
 sg13g2_xnor2_1 _42789_ (.Y(_12118_),
    .A(_09073_),
    .B(_12117_));
 sg13g2_nand2_1 _42790_ (.Y(_12119_),
    .A(net5736),
    .B(_09070_));
 sg13g2_o21ai_1 _42791_ (.B1(_12119_),
    .Y(_12120_),
    .A1(net5736),
    .A2(_12118_));
 sg13g2_nor2_1 _42792_ (.A(net5536),
    .B(_12120_),
    .Y(_12121_));
 sg13g2_xnor2_1 _42793_ (.Y(_12122_),
    .A(net5468),
    .B(_12120_));
 sg13g2_and2_1 _42794_ (.A(_12089_),
    .B(_12106_),
    .X(_12123_));
 sg13g2_a21oi_1 _42795_ (.A1(_12087_),
    .A2(_12105_),
    .Y(_12124_),
    .B1(net5473));
 sg13g2_a21oi_1 _42796_ (.A1(_12091_),
    .A2(_12123_),
    .Y(_12125_),
    .B1(_12124_));
 sg13g2_nor2_1 _42797_ (.A(_12056_),
    .B(_12077_),
    .Y(_12126_));
 sg13g2_nand2_1 _42798_ (.Y(_12127_),
    .A(_12123_),
    .B(_12126_));
 sg13g2_o21ai_1 _42799_ (.B1(_12125_),
    .Y(_12128_),
    .A1(_12065_),
    .A2(_12127_));
 sg13g2_and2_1 _42800_ (.A(_12122_),
    .B(_12128_),
    .X(_12129_));
 sg13g2_xnor2_1 _42801_ (.Y(_12130_),
    .A(_12122_),
    .B(_12128_));
 sg13g2_a21oi_1 _42802_ (.A1(net5537),
    .A2(_12130_),
    .Y(_12131_),
    .B1(_12121_));
 sg13g2_a22oi_1 _42803_ (.Y(_12132_),
    .B1(_12131_),
    .B2(net5231),
    .A2(_09083_),
    .A1(net5166));
 sg13g2_o21ai_1 _42804_ (.B1(_12132_),
    .Y(_12133_),
    .A1(net5120),
    .A2(_12105_));
 sg13g2_a22oi_1 _42805_ (.Y(_12134_),
    .B1(net6888),
    .B2(_12133_),
    .A2(net6467),
    .A1(net3462));
 sg13g2_inv_1 _42806_ (.Y(_00820_),
    .A(_12134_));
 sg13g2_nor2_1 _42807_ (.A(net5767),
    .B(_09058_),
    .Y(_12135_));
 sg13g2_o21ai_1 _42808_ (.B1(_09072_),
    .Y(_12136_),
    .A1(_09114_),
    .A2(_12102_));
 sg13g2_xnor2_1 _42809_ (.Y(_12137_),
    .A(_09060_),
    .B(_12136_));
 sg13g2_a21oi_2 _42810_ (.B1(_12135_),
    .Y(_12138_),
    .A2(_12137_),
    .A1(net5767));
 sg13g2_nor2_1 _42811_ (.A(net5421),
    .B(_12138_),
    .Y(_12139_));
 sg13g2_nand2_1 _42812_ (.Y(_12140_),
    .A(net5421),
    .B(_12138_));
 sg13g2_nand2b_1 _42813_ (.Y(_12141_),
    .B(_12140_),
    .A_N(_12139_));
 sg13g2_a21oi_1 _42814_ (.A1(net5421),
    .A2(_12120_),
    .Y(_12142_),
    .B1(_12129_));
 sg13g2_xnor2_1 _42815_ (.Y(_12143_),
    .A(_12141_),
    .B(_12142_));
 sg13g2_o21ai_1 _42816_ (.B1(net5964),
    .Y(_12144_),
    .A1(net5536),
    .A2(_12138_));
 sg13g2_a21oi_1 _42817_ (.A1(net5536),
    .A2(_12143_),
    .Y(_12145_),
    .B1(_12144_));
 sg13g2_a221oi_1 _42818_ (.B2(net5910),
    .C1(_12145_),
    .B1(_12120_),
    .A1(net5995),
    .Y(_12146_),
    .A2(_09076_));
 sg13g2_o21ai_1 _42819_ (.B1(net6884),
    .Y(_12147_),
    .A1(net5293),
    .A2(_09076_));
 sg13g2_a21oi_1 _42820_ (.A1(net5293),
    .A2(_12146_),
    .Y(_12148_),
    .B1(_12147_));
 sg13g2_a21o_1 _42821_ (.A2(net6470),
    .A1(net3334),
    .B1(_12148_),
    .X(_00821_));
 sg13g2_nand2_1 _42822_ (.Y(_12149_),
    .A(net2119),
    .B(net6467));
 sg13g2_o21ai_1 _42823_ (.B1(_09059_),
    .Y(_12150_),
    .A1(_09060_),
    .A2(_12136_));
 sg13g2_xnor2_1 _42824_ (.Y(_12151_),
    .A(_09064_),
    .B(_12150_));
 sg13g2_nor2_1 _42825_ (.A(net5767),
    .B(_09062_),
    .Y(_12152_));
 sg13g2_a21oi_2 _42826_ (.B1(_12152_),
    .Y(_12153_),
    .A2(_12151_),
    .A1(net5767));
 sg13g2_xnor2_1 _42827_ (.Y(_12154_),
    .A(net5421),
    .B(_12153_));
 sg13g2_o21ai_1 _42828_ (.B1(net5421),
    .Y(_12155_),
    .A1(_12120_),
    .A2(_12138_));
 sg13g2_nor2b_1 _42829_ (.A(_12129_),
    .B_N(_12155_),
    .Y(_12156_));
 sg13g2_or2_1 _42830_ (.X(_12157_),
    .B(_12156_),
    .A(_12139_));
 sg13g2_nor2_1 _42831_ (.A(_12154_),
    .B(_12157_),
    .Y(_12158_));
 sg13g2_and2_1 _42832_ (.A(_12154_),
    .B(_12157_),
    .X(_12159_));
 sg13g2_o21ai_1 _42833_ (.B1(net5536),
    .Y(_12160_),
    .A1(_12158_),
    .A2(_12159_));
 sg13g2_o21ai_1 _42834_ (.B1(_12160_),
    .Y(_12161_),
    .A1(net5536),
    .A2(_12153_));
 sg13g2_nor2_1 _42835_ (.A(net5153),
    .B(_12161_),
    .Y(_12162_));
 sg13g2_a221oi_1 _42836_ (.B2(net5218),
    .C1(_12162_),
    .B1(_12138_),
    .A1(net5167),
    .Y(_12163_),
    .A2(_09070_));
 sg13g2_o21ai_1 _42837_ (.B1(_12149_),
    .Y(_00822_),
    .A1(net6864),
    .A2(_12163_));
 sg13g2_nand2_1 _42838_ (.Y(_12164_),
    .A(net5725),
    .B(_09045_));
 sg13g2_a21oi_2 _42839_ (.B1(_09079_),
    .Y(_12165_),
    .A2(_12101_),
    .A1(_09119_));
 sg13g2_o21ai_1 _42840_ (.B1(_09048_),
    .Y(_12166_),
    .A1(_09116_),
    .A2(_12165_));
 sg13g2_nor3_1 _42841_ (.A(_09048_),
    .B(_09116_),
    .C(_12165_),
    .Y(_12167_));
 sg13g2_nand3b_1 _42842_ (.B(net5765),
    .C(_12166_),
    .Y(_12168_),
    .A_N(_12167_));
 sg13g2_nand2_2 _42843_ (.Y(_12169_),
    .A(_12164_),
    .B(_12168_));
 sg13g2_xnor2_1 _42844_ (.Y(_12170_),
    .A(net5421),
    .B(_12169_));
 sg13g2_a21oi_1 _42845_ (.A1(net5421),
    .A2(_12153_),
    .Y(_12171_),
    .B1(_12158_));
 sg13g2_xnor2_1 _42846_ (.Y(_12172_),
    .A(_12170_),
    .B(_12171_));
 sg13g2_o21ai_1 _42847_ (.B1(net5964),
    .Y(_12173_),
    .A1(net5536),
    .A2(_12169_));
 sg13g2_a21oi_1 _42848_ (.A1(net5536),
    .A2(_12172_),
    .Y(_12174_),
    .B1(_12173_));
 sg13g2_a221oi_1 _42849_ (.B2(net5910),
    .C1(_12174_),
    .B1(_12153_),
    .A1(net5995),
    .Y(_12175_),
    .A2(_09058_));
 sg13g2_o21ai_1 _42850_ (.B1(net6884),
    .Y(_12176_),
    .A1(net5293),
    .A2(_09058_));
 sg13g2_a21oi_1 _42851_ (.A1(net5293),
    .A2(_12175_),
    .Y(_12177_),
    .B1(_12176_));
 sg13g2_a21o_1 _42852_ (.A2(net6467),
    .A1(net3510),
    .B1(_12177_),
    .X(_00823_));
 sg13g2_nand2_1 _42853_ (.Y(_12178_),
    .A(_09046_),
    .B(_12166_));
 sg13g2_xor2_1 _42854_ (.B(_12178_),
    .A(_09042_),
    .X(_12179_));
 sg13g2_nand2_1 _42855_ (.Y(_12180_),
    .A(net5725),
    .B(_09039_));
 sg13g2_o21ai_1 _42856_ (.B1(_12180_),
    .Y(_12181_),
    .A1(net5725),
    .A2(_12179_));
 sg13g2_nand2_1 _42857_ (.Y(_12182_),
    .A(net5418),
    .B(_12181_));
 sg13g2_xnor2_1 _42858_ (.Y(_12183_),
    .A(net5465),
    .B(_12181_));
 sg13g2_or2_1 _42859_ (.X(_12184_),
    .B(_12170_),
    .A(_12154_));
 sg13g2_nand3b_1 _42860_ (.B(_12140_),
    .C(_12122_),
    .Y(_12185_),
    .A_N(_12139_));
 sg13g2_nor3_1 _42861_ (.A(_12125_),
    .B(_12184_),
    .C(_12185_),
    .Y(_12186_));
 sg13g2_o21ai_1 _42862_ (.B1(net5421),
    .Y(_12187_),
    .A1(_12153_),
    .A2(_12169_));
 sg13g2_o21ai_1 _42863_ (.B1(_12187_),
    .Y(_12188_),
    .A1(_12155_),
    .A2(_12184_));
 sg13g2_nor2_1 _42864_ (.A(_12186_),
    .B(_12188_),
    .Y(_12189_));
 sg13g2_or3_1 _42865_ (.A(_12127_),
    .B(_12184_),
    .C(_12185_),
    .X(_12190_));
 sg13g2_o21ai_1 _42866_ (.B1(_12189_),
    .Y(_12191_),
    .A1(_12065_),
    .A2(_12190_));
 sg13g2_and2_1 _42867_ (.A(_12183_),
    .B(_12191_),
    .X(_12192_));
 sg13g2_xnor2_1 _42868_ (.Y(_12193_),
    .A(_12183_),
    .B(_12191_));
 sg13g2_o21ai_1 _42869_ (.B1(net5964),
    .Y(_12194_),
    .A1(net5534),
    .A2(_12181_));
 sg13g2_a21oi_1 _42870_ (.A1(net5534),
    .A2(_12193_),
    .Y(_12195_),
    .B1(_12194_));
 sg13g2_a221oi_1 _42871_ (.B2(net5910),
    .C1(_12195_),
    .B1(_12169_),
    .A1(net5995),
    .Y(_12196_),
    .A2(_09062_));
 sg13g2_o21ai_1 _42872_ (.B1(net6884),
    .Y(_12197_),
    .A1(net5290),
    .A2(_09062_));
 sg13g2_a21oi_1 _42873_ (.A1(net5290),
    .A2(_12196_),
    .Y(_12198_),
    .B1(_12197_));
 sg13g2_a21o_1 _42874_ (.A2(net6467),
    .A1(net3494),
    .B1(_12198_),
    .X(_00824_));
 sg13g2_a21oi_1 _42875_ (.A1(net5418),
    .A2(_12181_),
    .Y(_12199_),
    .B1(_12192_));
 sg13g2_nor2_1 _42876_ (.A(net5765),
    .B(_09033_),
    .Y(_12200_));
 sg13g2_a21oi_1 _42877_ (.A1(_09107_),
    .A2(_12166_),
    .Y(_12201_),
    .B1(_09041_));
 sg13g2_xnor2_1 _42878_ (.Y(_12202_),
    .A(_09035_),
    .B(_12201_));
 sg13g2_a21oi_2 _42879_ (.B1(_12200_),
    .Y(_12203_),
    .A2(_12202_),
    .A1(net5765));
 sg13g2_nor2_1 _42880_ (.A(net5419),
    .B(_12203_),
    .Y(_12204_));
 sg13g2_nand2b_1 _42881_ (.Y(_12205_),
    .B(net5465),
    .A_N(_12203_));
 sg13g2_nand2_1 _42882_ (.Y(_12206_),
    .A(net5418),
    .B(_12203_));
 sg13g2_nand2_1 _42883_ (.Y(_12207_),
    .A(_12205_),
    .B(_12206_));
 sg13g2_xnor2_1 _42884_ (.Y(_12208_),
    .A(_12199_),
    .B(_12207_));
 sg13g2_o21ai_1 _42885_ (.B1(net5968),
    .Y(_12209_),
    .A1(net5534),
    .A2(_12203_));
 sg13g2_a21oi_1 _42886_ (.A1(net5535),
    .A2(_12208_),
    .Y(_12210_),
    .B1(_12209_));
 sg13g2_a221oi_1 _42887_ (.B2(net5909),
    .C1(_12210_),
    .B1(_12181_),
    .A1(net5994),
    .Y(_12211_),
    .A2(_09045_));
 sg13g2_o21ai_1 _42888_ (.B1(net6884),
    .Y(_12212_),
    .A1(net5290),
    .A2(_09045_));
 sg13g2_a21oi_1 _42889_ (.A1(net5290),
    .A2(_12211_),
    .Y(_12213_),
    .B1(_12212_));
 sg13g2_a21o_1 _42890_ (.A2(net6467),
    .A1(net2538),
    .B1(_12213_),
    .X(_00825_));
 sg13g2_a21oi_1 _42891_ (.A1(_09035_),
    .A2(_12201_),
    .Y(_12214_),
    .B1(_09034_));
 sg13g2_xnor2_1 _42892_ (.Y(_12215_),
    .A(_09026_),
    .B(_12214_));
 sg13g2_nor2_1 _42893_ (.A(net5765),
    .B(_09024_),
    .Y(_12216_));
 sg13g2_a21oi_2 _42894_ (.B1(_12216_),
    .Y(_12217_),
    .A2(_12215_),
    .A1(net5765));
 sg13g2_nor2_1 _42895_ (.A(net5534),
    .B(_12217_),
    .Y(_12218_));
 sg13g2_nand2_1 _42896_ (.Y(_12219_),
    .A(net5418),
    .B(_12217_));
 sg13g2_xnor2_1 _42897_ (.Y(_12220_),
    .A(net5418),
    .B(_12217_));
 sg13g2_nand2_1 _42898_ (.Y(_12221_),
    .A(_12182_),
    .B(_12206_));
 sg13g2_nor2_1 _42899_ (.A(_12192_),
    .B(_12221_),
    .Y(_12222_));
 sg13g2_or3_1 _42900_ (.A(_12204_),
    .B(_12220_),
    .C(_12222_),
    .X(_12223_));
 sg13g2_o21ai_1 _42901_ (.B1(_12220_),
    .Y(_12224_),
    .A1(_12204_),
    .A2(_12222_));
 sg13g2_a21oi_1 _42902_ (.A1(_12223_),
    .A2(_12224_),
    .Y(_12225_),
    .B1(net5565));
 sg13g2_nor2_1 _42903_ (.A(_12218_),
    .B(_12225_),
    .Y(_12226_));
 sg13g2_a22oi_1 _42904_ (.Y(_12227_),
    .B1(_12226_),
    .B2(net5230),
    .A2(_12203_),
    .A1(net5218));
 sg13g2_a22oi_1 _42905_ (.Y(_12228_),
    .B1(net5107),
    .B2(_09039_),
    .A2(net6467),
    .A1(net3566));
 sg13g2_o21ai_1 _42906_ (.B1(_12228_),
    .Y(_00826_),
    .A1(net6862),
    .A2(_12227_));
 sg13g2_nand2_1 _42907_ (.Y(_12229_),
    .A(net2316),
    .B(net6467));
 sg13g2_o21ai_1 _42908_ (.B1(_09049_),
    .Y(_12230_),
    .A1(_09116_),
    .A2(_12165_));
 sg13g2_a21oi_1 _42909_ (.A1(_09109_),
    .A2(_12230_),
    .Y(_12231_),
    .B1(_09020_));
 sg13g2_and3_1 _42910_ (.X(_12232_),
    .A(_09020_),
    .B(_09109_),
    .C(_12230_));
 sg13g2_nor3_1 _42911_ (.A(net5725),
    .B(_12231_),
    .C(_12232_),
    .Y(_12233_));
 sg13g2_a21oi_2 _42912_ (.B1(_12233_),
    .Y(_12234_),
    .A2(_09018_),
    .A1(net5725));
 sg13g2_xnor2_1 _42913_ (.Y(_12235_),
    .A(net5418),
    .B(_12234_));
 sg13g2_nand2_1 _42914_ (.Y(_12236_),
    .A(_12219_),
    .B(_12223_));
 sg13g2_xor2_1 _42915_ (.B(_12236_),
    .A(_12235_),
    .X(_12237_));
 sg13g2_a21oi_1 _42916_ (.A1(net5565),
    .A2(_12234_),
    .Y(_12238_),
    .B1(net5931));
 sg13g2_o21ai_1 _42917_ (.B1(_12238_),
    .Y(_12239_),
    .A1(net5565),
    .A2(_12237_));
 sg13g2_a22oi_1 _42918_ (.Y(_12240_),
    .B1(_12217_),
    .B2(net5910),
    .A2(_09033_),
    .A1(net5995));
 sg13g2_and3_1 _42919_ (.X(_12241_),
    .A(net5290),
    .B(_12239_),
    .C(_12240_));
 sg13g2_o21ai_1 _42920_ (.B1(net6885),
    .Y(_12242_),
    .A1(net5296),
    .A2(_09033_));
 sg13g2_o21ai_1 _42921_ (.B1(_12229_),
    .Y(_00827_),
    .A1(_12241_),
    .A2(_12242_));
 sg13g2_nand2_1 _42922_ (.Y(_12243_),
    .A(net5725),
    .B(_09011_));
 sg13g2_a21oi_1 _42923_ (.A1(net5668),
    .A2(_09018_),
    .Y(_12244_),
    .B1(_12231_));
 sg13g2_xnor2_1 _42924_ (.Y(_12245_),
    .A(_09014_),
    .B(_12244_));
 sg13g2_o21ai_1 _42925_ (.B1(_12243_),
    .Y(_12246_),
    .A1(net5725),
    .A2(_12245_));
 sg13g2_nand2_1 _42926_ (.Y(_12247_),
    .A(net5418),
    .B(_12246_));
 sg13g2_xnor2_1 _42927_ (.Y(_12248_),
    .A(net5465),
    .B(_12246_));
 sg13g2_nor2b_1 _42928_ (.A(_12220_),
    .B_N(_12235_),
    .Y(_12249_));
 sg13g2_o21ai_1 _42929_ (.B1(_12219_),
    .Y(_12250_),
    .A1(net5465),
    .A2(_12234_));
 sg13g2_a21o_1 _42930_ (.A2(_12249_),
    .A1(_12221_),
    .B1(_12250_),
    .X(_12251_));
 sg13g2_and3_1 _42931_ (.X(_12252_),
    .A(_12183_),
    .B(_12205_),
    .C(_12206_));
 sg13g2_nand3b_1 _42932_ (.B(_12235_),
    .C(_12252_),
    .Y(_12253_),
    .A_N(_12220_));
 sg13g2_nor2b_1 _42933_ (.A(_12253_),
    .B_N(_12191_),
    .Y(_12254_));
 sg13g2_nor2_1 _42934_ (.A(_12251_),
    .B(_12254_),
    .Y(_12255_));
 sg13g2_nand2b_1 _42935_ (.Y(_12256_),
    .B(_12248_),
    .A_N(_12255_));
 sg13g2_xor2_1 _42936_ (.B(_12255_),
    .A(_12248_),
    .X(_12257_));
 sg13g2_nor2_1 _42937_ (.A(net5534),
    .B(_12246_),
    .Y(_12258_));
 sg13g2_a21oi_1 _42938_ (.A1(net5534),
    .A2(_12257_),
    .Y(_12259_),
    .B1(_12258_));
 sg13g2_nor2_1 _42939_ (.A(net5120),
    .B(_12234_),
    .Y(_12260_));
 sg13g2_nand2_1 _42940_ (.Y(_12261_),
    .A(net1638),
    .B(net6454));
 sg13g2_a221oi_1 _42941_ (.B2(net5232),
    .C1(_12260_),
    .B1(_12259_),
    .A1(net5165),
    .Y(_12262_),
    .A2(_09024_));
 sg13g2_o21ai_1 _42942_ (.B1(_12261_),
    .Y(_00828_),
    .A1(net6864),
    .A2(_12262_));
 sg13g2_nor2_1 _42943_ (.A(net5765),
    .B(_09001_),
    .Y(_12263_));
 sg13g2_o21ai_1 _42944_ (.B1(_09012_),
    .Y(_12264_),
    .A1(_09111_),
    .A2(_12231_));
 sg13g2_xnor2_1 _42945_ (.Y(_12265_),
    .A(_09003_),
    .B(_12264_));
 sg13g2_a21oi_2 _42946_ (.B1(_12263_),
    .Y(_12266_),
    .A2(_12265_),
    .A1(net5765));
 sg13g2_nor2_1 _42947_ (.A(net5419),
    .B(_12266_),
    .Y(_12267_));
 sg13g2_xnor2_1 _42948_ (.Y(_12268_),
    .A(net5465),
    .B(_12266_));
 sg13g2_nand2_1 _42949_ (.Y(_12269_),
    .A(_12247_),
    .B(_12256_));
 sg13g2_xnor2_1 _42950_ (.Y(_12270_),
    .A(_12268_),
    .B(_12269_));
 sg13g2_o21ai_1 _42951_ (.B1(net5964),
    .Y(_12271_),
    .A1(net5534),
    .A2(_12266_));
 sg13g2_a21oi_1 _42952_ (.A1(net5534),
    .A2(_12270_),
    .Y(_12272_),
    .B1(_12271_));
 sg13g2_a221oi_1 _42953_ (.B2(net5911),
    .C1(_12272_),
    .B1(_12246_),
    .A1(net5996),
    .Y(_12273_),
    .A2(_09018_));
 sg13g2_o21ai_1 _42954_ (.B1(net6884),
    .Y(_12274_),
    .A1(net5290),
    .A2(_09018_));
 sg13g2_a21oi_1 _42955_ (.A1(net5290),
    .A2(_12273_),
    .Y(_12275_),
    .B1(_12274_));
 sg13g2_a21o_1 _42956_ (.A2(net6454),
    .A1(net2475),
    .B1(_12275_),
    .X(_00829_));
 sg13g2_o21ai_1 _42957_ (.B1(_09002_),
    .Y(_12276_),
    .A1(_09003_),
    .A2(_12264_));
 sg13g2_xnor2_1 _42958_ (.Y(_12277_),
    .A(_09007_),
    .B(_12276_));
 sg13g2_nand2_1 _42959_ (.Y(_12278_),
    .A(net5732),
    .B(_09006_));
 sg13g2_o21ai_1 _42960_ (.B1(_12278_),
    .Y(_12279_),
    .A1(net5725),
    .A2(_12277_));
 sg13g2_inv_1 _42961_ (.Y(_12280_),
    .A(_12279_));
 sg13g2_xnor2_1 _42962_ (.Y(_12281_),
    .A(net5465),
    .B(_12279_));
 sg13g2_o21ai_1 _42963_ (.B1(net5419),
    .Y(_12282_),
    .A1(_12246_),
    .A2(_12266_));
 sg13g2_a21oi_1 _42964_ (.A1(_12256_),
    .A2(_12282_),
    .Y(_12283_),
    .B1(_12267_));
 sg13g2_nand2b_1 _42965_ (.Y(_12284_),
    .B(_12283_),
    .A_N(_12281_));
 sg13g2_xnor2_1 _42966_ (.Y(_12285_),
    .A(_12281_),
    .B(_12283_));
 sg13g2_o21ai_1 _42967_ (.B1(net5964),
    .Y(_12286_),
    .A1(net5565),
    .A2(_12285_));
 sg13g2_a21oi_1 _42968_ (.A1(net5565),
    .A2(_12279_),
    .Y(_12287_),
    .B1(_12286_));
 sg13g2_a221oi_1 _42969_ (.B2(net5911),
    .C1(_12287_),
    .B1(_12266_),
    .A1(net5996),
    .Y(_12288_),
    .A2(_09011_));
 sg13g2_o21ai_1 _42970_ (.B1(net6884),
    .Y(_12289_),
    .A1(net5296),
    .A2(_09011_));
 sg13g2_a21oi_1 _42971_ (.A1(net5290),
    .A2(_12288_),
    .Y(_12290_),
    .B1(_12289_));
 sg13g2_a21o_1 _42972_ (.A2(net6467),
    .A1(net3175),
    .B1(_12290_),
    .X(_00830_));
 sg13g2_nand2_1 _42973_ (.Y(_12291_),
    .A(net2083),
    .B(net6468));
 sg13g2_a21o_1 _42974_ (.A2(_09661_),
    .A1(_09124_),
    .B1(_09899_),
    .X(_12292_));
 sg13g2_nor2_1 _42975_ (.A(_09662_),
    .B(_09898_),
    .Y(_12293_));
 sg13g2_nor2_1 _42976_ (.A(net5731),
    .B(_12293_),
    .Y(_12294_));
 sg13g2_a22oi_1 _42977_ (.Y(_12295_),
    .B1(_12292_),
    .B2(_12294_),
    .A2(_09896_),
    .A1(net5731));
 sg13g2_xnor2_1 _42978_ (.Y(_12296_),
    .A(net5418),
    .B(_12295_));
 sg13g2_inv_2 _42979_ (.Y(_12297_),
    .A(_12296_));
 sg13g2_o21ai_1 _42980_ (.B1(_12284_),
    .Y(_12298_),
    .A1(net5465),
    .A2(_12279_));
 sg13g2_xnor2_1 _42981_ (.Y(_12299_),
    .A(_12297_),
    .B(_12298_));
 sg13g2_a21oi_1 _42982_ (.A1(net5565),
    .A2(_12295_),
    .Y(_12300_),
    .B1(net5932));
 sg13g2_o21ai_1 _42983_ (.B1(_12300_),
    .Y(_12301_),
    .A1(net5565),
    .A2(_12299_));
 sg13g2_a22oi_1 _42984_ (.Y(_12302_),
    .B1(_12280_),
    .B2(net5911),
    .A2(_09001_),
    .A1(net5996));
 sg13g2_and3_1 _42985_ (.X(_12303_),
    .A(net5296),
    .B(_12301_),
    .C(_12302_));
 sg13g2_o21ai_1 _42986_ (.B1(net6884),
    .Y(_12304_),
    .A1(net5296),
    .A2(_09001_));
 sg13g2_o21ai_1 _42987_ (.B1(_12291_),
    .Y(_00831_),
    .A1(_12303_),
    .A2(_12304_));
 sg13g2_nand2_1 _42988_ (.Y(_12305_),
    .A(_09897_),
    .B(_12292_));
 sg13g2_xnor2_1 _42989_ (.Y(_12306_),
    .A(_09892_),
    .B(_12305_));
 sg13g2_nand2_1 _42990_ (.Y(_12307_),
    .A(net5731),
    .B(_09890_));
 sg13g2_o21ai_1 _42991_ (.B1(_12307_),
    .Y(_12308_),
    .A1(net5731),
    .A2(_12306_));
 sg13g2_xnor2_1 _42992_ (.Y(_12309_),
    .A(net5469),
    .B(_12308_));
 sg13g2_nand2_1 _42993_ (.Y(_12310_),
    .A(_12248_),
    .B(_12268_));
 sg13g2_nor3_1 _42994_ (.A(_12281_),
    .B(_12297_),
    .C(_12310_),
    .Y(_12311_));
 sg13g2_nor4_1 _42995_ (.A(_12253_),
    .B(_12281_),
    .C(_12297_),
    .D(_12310_),
    .Y(_12312_));
 sg13g2_nor2b_1 _42996_ (.A(_12190_),
    .B_N(_12312_),
    .Y(_12313_));
 sg13g2_nand2_1 _42997_ (.Y(_12314_),
    .A(_12064_),
    .B(_12313_));
 sg13g2_a21oi_1 _42998_ (.A1(net1074),
    .A2(net1143),
    .Y(_12315_),
    .B1(_12314_));
 sg13g2_nand2_1 _42999_ (.Y(_12316_),
    .A(_12062_),
    .B(_12313_));
 sg13g2_nand2b_1 _43000_ (.Y(_12317_),
    .B(_12312_),
    .A_N(_12189_));
 sg13g2_nand2_1 _43001_ (.Y(_12318_),
    .A(_12251_),
    .B(_12311_));
 sg13g2_nor3_1 _43002_ (.A(_12281_),
    .B(_12282_),
    .C(_12297_),
    .Y(_12319_));
 sg13g2_a21oi_1 _43003_ (.A1(_12279_),
    .A2(_12295_),
    .Y(_12320_),
    .B1(net5465));
 sg13g2_nor2_1 _43004_ (.A(_12319_),
    .B(_12320_),
    .Y(_12321_));
 sg13g2_nand4_1 _43005_ (.B(_12317_),
    .C(_12318_),
    .A(_12316_),
    .Y(_12322_),
    .D(_12321_));
 sg13g2_or2_1 _43006_ (.X(_12323_),
    .B(_12322_),
    .A(_12315_));
 sg13g2_and2_1 _43007_ (.A(_12309_),
    .B(_12323_),
    .X(_12324_));
 sg13g2_xnor2_1 _43008_ (.Y(_12325_),
    .A(_12309_),
    .B(_12323_));
 sg13g2_a21oi_1 _43009_ (.A1(net5539),
    .A2(_12325_),
    .Y(_12326_),
    .B1(net5932));
 sg13g2_o21ai_1 _43010_ (.B1(_12326_),
    .Y(_12327_),
    .A1(net5539),
    .A2(_12308_));
 sg13g2_nand2b_1 _43011_ (.Y(_12328_),
    .B(net5996),
    .A_N(_09006_));
 sg13g2_nand2b_1 _43012_ (.Y(_12329_),
    .B(net5911),
    .A_N(_12295_));
 sg13g2_nand4_1 _43013_ (.B(_12327_),
    .C(_12328_),
    .A(net5295),
    .Y(_12330_),
    .D(_12329_));
 sg13g2_nor2b_1 _43014_ (.A(net5295),
    .B_N(_09006_),
    .Y(_12331_));
 sg13g2_nor2_1 _43015_ (.A(net6862),
    .B(_12331_),
    .Y(_12332_));
 sg13g2_a22oi_1 _43016_ (.Y(_12333_),
    .B1(_12330_),
    .B2(_12332_),
    .A2(net6468),
    .A1(net3723));
 sg13g2_inv_1 _43017_ (.Y(_00832_),
    .A(_12333_));
 sg13g2_a21oi_1 _43018_ (.A1(net5422),
    .A2(_12308_),
    .Y(_12334_),
    .B1(_12324_));
 sg13g2_a22oi_1 _43019_ (.Y(_12335_),
    .B1(_09908_),
    .B2(_12292_),
    .A2(_09891_),
    .A1(net5601));
 sg13g2_xnor2_1 _43020_ (.Y(_12336_),
    .A(_09882_),
    .B(_12335_));
 sg13g2_nand2_1 _43021_ (.Y(_12337_),
    .A(net5770),
    .B(_12336_));
 sg13g2_o21ai_1 _43022_ (.B1(_12337_),
    .Y(_12338_),
    .A1(net5770),
    .A2(_09878_));
 sg13g2_or2_1 _43023_ (.X(_12339_),
    .B(_12338_),
    .A(net5422));
 sg13g2_xnor2_1 _43024_ (.Y(_12340_),
    .A(net5469),
    .B(_12338_));
 sg13g2_xor2_1 _43025_ (.B(_12340_),
    .A(_12334_),
    .X(_12341_));
 sg13g2_o21ai_1 _43026_ (.B1(net5964),
    .Y(_12342_),
    .A1(net5539),
    .A2(_12338_));
 sg13g2_a21oi_1 _43027_ (.A1(net5540),
    .A2(_12341_),
    .Y(_12343_),
    .B1(_12342_));
 sg13g2_a221oi_1 _43028_ (.B2(net5911),
    .C1(_12343_),
    .B1(_12308_),
    .A1(net5996),
    .Y(_12344_),
    .A2(_09896_));
 sg13g2_o21ai_1 _43029_ (.B1(net6885),
    .Y(_12345_),
    .A1(net5302),
    .A2(_09896_));
 sg13g2_a21oi_1 _43030_ (.A1(net5295),
    .A2(_12344_),
    .Y(_12346_),
    .B1(_12345_));
 sg13g2_a21o_1 _43031_ (.A2(net6471),
    .A1(net2319),
    .B1(_12346_),
    .X(_00833_));
 sg13g2_nand2_1 _43032_ (.Y(_12347_),
    .A(net5730),
    .B(_09885_));
 sg13g2_a21oi_1 _43033_ (.A1(_09881_),
    .A2(_12335_),
    .Y(_12348_),
    .B1(_09880_));
 sg13g2_xor2_1 _43034_ (.B(_12348_),
    .A(_09886_),
    .X(_12349_));
 sg13g2_o21ai_1 _43035_ (.B1(_12347_),
    .Y(_12350_),
    .A1(net5730),
    .A2(_12349_));
 sg13g2_nand2_1 _43036_ (.Y(_12351_),
    .A(net5422),
    .B(_12350_));
 sg13g2_xnor2_1 _43037_ (.Y(_12352_),
    .A(net5469),
    .B(_12350_));
 sg13g2_o21ai_1 _43038_ (.B1(net5422),
    .Y(_12353_),
    .A1(_12308_),
    .A2(_12338_));
 sg13g2_nand2b_1 _43039_ (.Y(_12354_),
    .B(_12353_),
    .A_N(_12324_));
 sg13g2_nand3_1 _43040_ (.B(_12352_),
    .C(_12354_),
    .A(_12339_),
    .Y(_12355_));
 sg13g2_a21o_1 _43041_ (.A2(_12354_),
    .A1(_12339_),
    .B1(_12352_),
    .X(_12356_));
 sg13g2_and2_1 _43042_ (.A(_12355_),
    .B(_12356_),
    .X(_12357_));
 sg13g2_mux2_1 _43043_ (.A0(_12350_),
    .A1(_12357_),
    .S(net5539),
    .X(_12358_));
 sg13g2_a22oi_1 _43044_ (.Y(_12359_),
    .B1(_12358_),
    .B2(net5230),
    .A2(_12338_),
    .A1(net5218));
 sg13g2_a22oi_1 _43045_ (.Y(_12360_),
    .B1(net5107),
    .B2(_09890_),
    .A2(net6468),
    .A1(net3652));
 sg13g2_o21ai_1 _43046_ (.B1(_12360_),
    .Y(_00834_),
    .A1(net6862),
    .A2(_12359_));
 sg13g2_nand2_1 _43047_ (.Y(_12361_),
    .A(net5730),
    .B(_09869_));
 sg13g2_a21oi_1 _43048_ (.A1(_09662_),
    .A2(_09901_),
    .Y(_12362_),
    .B1(_09910_));
 sg13g2_xnor2_1 _43049_ (.Y(_12363_),
    .A(_09872_),
    .B(_12362_));
 sg13g2_o21ai_1 _43050_ (.B1(_12361_),
    .Y(_12364_),
    .A1(net5730),
    .A2(_12363_));
 sg13g2_xnor2_1 _43051_ (.Y(_12365_),
    .A(net5469),
    .B(_12364_));
 sg13g2_nand2_1 _43052_ (.Y(_12366_),
    .A(_12351_),
    .B(_12355_));
 sg13g2_xnor2_1 _43053_ (.Y(_12367_),
    .A(_12365_),
    .B(_12366_));
 sg13g2_o21ai_1 _43054_ (.B1(net5967),
    .Y(_12368_),
    .A1(net5539),
    .A2(_12364_));
 sg13g2_a21oi_1 _43055_ (.A1(net5539),
    .A2(_12367_),
    .Y(_12369_),
    .B1(_12368_));
 sg13g2_a221oi_1 _43056_ (.B2(net5911),
    .C1(_12369_),
    .B1(_12350_),
    .A1(net5996),
    .Y(_12370_),
    .A2(_09879_));
 sg13g2_o21ai_1 _43057_ (.B1(net6885),
    .Y(_12371_),
    .A1(net5295),
    .A2(_09879_));
 sg13g2_a21oi_1 _43058_ (.A1(net5295),
    .A2(_12370_),
    .Y(_12372_),
    .B1(_12371_));
 sg13g2_a21oi_1 _43059_ (.A1(net2972),
    .A2(net6468),
    .Y(_12373_),
    .B1(_12372_));
 sg13g2_inv_1 _43060_ (.Y(_00835_),
    .A(_12373_));
 sg13g2_o21ai_1 _43061_ (.B1(_09870_),
    .Y(_12374_),
    .A1(_09872_),
    .A2(_12362_));
 sg13g2_xnor2_1 _43062_ (.Y(_12375_),
    .A(_09866_),
    .B(_12374_));
 sg13g2_nand2_1 _43063_ (.Y(_12376_),
    .A(net5730),
    .B(_09863_));
 sg13g2_o21ai_1 _43064_ (.B1(_12376_),
    .Y(_12377_),
    .A1(net5730),
    .A2(_12375_));
 sg13g2_nor2_1 _43065_ (.A(net5540),
    .B(_12377_),
    .Y(_12378_));
 sg13g2_nand2_1 _43066_ (.Y(_12379_),
    .A(net5422),
    .B(_12377_));
 sg13g2_inv_1 _43067_ (.Y(_12380_),
    .A(_12379_));
 sg13g2_xnor2_1 _43068_ (.Y(_12381_),
    .A(net5422),
    .B(_12377_));
 sg13g2_nand2_1 _43069_ (.Y(_12382_),
    .A(_12352_),
    .B(_12365_));
 sg13g2_o21ai_1 _43070_ (.B1(net5422),
    .Y(_12383_),
    .A1(_12350_),
    .A2(_12364_));
 sg13g2_o21ai_1 _43071_ (.B1(_12383_),
    .Y(_12384_),
    .A1(_12353_),
    .A2(_12382_));
 sg13g2_and4_1 _43072_ (.A(_12309_),
    .B(_12340_),
    .C(_12352_),
    .D(_12365_),
    .X(_12385_));
 sg13g2_a21oi_1 _43073_ (.A1(_12323_),
    .A2(_12385_),
    .Y(_12386_),
    .B1(_12384_));
 sg13g2_nor2_1 _43074_ (.A(_12381_),
    .B(_12386_),
    .Y(_12387_));
 sg13g2_xnor2_1 _43075_ (.Y(_12388_),
    .A(_12381_),
    .B(_12386_));
 sg13g2_a21oi_1 _43076_ (.A1(net5540),
    .A2(_12388_),
    .Y(_12389_),
    .B1(_12378_));
 sg13g2_a22oi_1 _43077_ (.Y(_12390_),
    .B1(_12389_),
    .B2(net5231),
    .A2(_12364_),
    .A1(net5218));
 sg13g2_a22oi_1 _43078_ (.Y(_12391_),
    .B1(net5107),
    .B2(_09885_),
    .A2(net6471),
    .A1(net3664));
 sg13g2_o21ai_1 _43079_ (.B1(_12391_),
    .Y(_00836_),
    .A1(net6861),
    .A2(_12390_));
 sg13g2_a21o_1 _43080_ (.A2(_12374_),
    .A1(_09865_),
    .B1(_09864_),
    .X(_12392_));
 sg13g2_xnor2_1 _43081_ (.Y(_12393_),
    .A(_09859_),
    .B(_12392_));
 sg13g2_nand2_1 _43082_ (.Y(_12394_),
    .A(net5732),
    .B(_09857_));
 sg13g2_o21ai_1 _43083_ (.B1(_12394_),
    .Y(_12395_),
    .A1(net5730),
    .A2(_12393_));
 sg13g2_nor2_1 _43084_ (.A(net5423),
    .B(_12395_),
    .Y(_12396_));
 sg13g2_xnor2_1 _43085_ (.Y(_12397_),
    .A(net5423),
    .B(_12395_));
 sg13g2_nor2_1 _43086_ (.A(_12380_),
    .B(_12387_),
    .Y(_12398_));
 sg13g2_xnor2_1 _43087_ (.Y(_12399_),
    .A(_12397_),
    .B(_12398_));
 sg13g2_o21ai_1 _43088_ (.B1(net5966),
    .Y(_12400_),
    .A1(net5540),
    .A2(_12395_));
 sg13g2_a21oi_1 _43089_ (.A1(net5540),
    .A2(_12399_),
    .Y(_12401_),
    .B1(_12400_));
 sg13g2_a221oi_1 _43090_ (.B2(net5913),
    .C1(_12401_),
    .B1(_12377_),
    .A1(net5998),
    .Y(_12402_),
    .A2(_09869_));
 sg13g2_o21ai_1 _43091_ (.B1(net6887),
    .Y(_12403_),
    .A1(net5295),
    .A2(_09869_));
 sg13g2_a21oi_1 _43092_ (.A1(net5302),
    .A2(_12402_),
    .Y(_12404_),
    .B1(_12403_));
 sg13g2_a21o_1 _43093_ (.A2(net6471),
    .A1(net1701),
    .B1(_12404_),
    .X(_00837_));
 sg13g2_nand2_1 _43094_ (.Y(_12405_),
    .A(net5730),
    .B(_09848_));
 sg13g2_a21oi_1 _43095_ (.A1(_09859_),
    .A2(_12392_),
    .Y(_12406_),
    .B1(_09858_));
 sg13g2_xor2_1 _43096_ (.B(_12406_),
    .A(_09849_),
    .X(_12407_));
 sg13g2_o21ai_1 _43097_ (.B1(_12405_),
    .Y(_12408_),
    .A1(net5731),
    .A2(_12407_));
 sg13g2_nor2_1 _43098_ (.A(net5540),
    .B(_12408_),
    .Y(_12409_));
 sg13g2_nand2_1 _43099_ (.Y(_12410_),
    .A(net5423),
    .B(_12408_));
 sg13g2_xnor2_1 _43100_ (.Y(_12411_),
    .A(net5473),
    .B(_12408_));
 sg13g2_a21o_1 _43101_ (.A2(_12395_),
    .A1(net5423),
    .B1(_12380_),
    .X(_12412_));
 sg13g2_nor2_1 _43102_ (.A(_12387_),
    .B(_12412_),
    .Y(_12413_));
 sg13g2_nor2_1 _43103_ (.A(_12396_),
    .B(_12413_),
    .Y(_12414_));
 sg13g2_nand2_1 _43104_ (.Y(_12415_),
    .A(_12411_),
    .B(_12414_));
 sg13g2_xnor2_1 _43105_ (.Y(_12416_),
    .A(_12411_),
    .B(_12414_));
 sg13g2_a21oi_1 _43106_ (.A1(net5540),
    .A2(_12416_),
    .Y(_12417_),
    .B1(_12409_));
 sg13g2_a22oi_1 _43107_ (.Y(_12418_),
    .B1(_12417_),
    .B2(net5231),
    .A2(_12395_),
    .A1(net5218));
 sg13g2_a22oi_1 _43108_ (.Y(_12419_),
    .B1(net5107),
    .B2(_09863_),
    .A2(net6471),
    .A1(net3119));
 sg13g2_o21ai_1 _43109_ (.B1(_12419_),
    .Y(_00838_),
    .A1(net6861),
    .A2(_12418_));
 sg13g2_nand2_1 _43110_ (.Y(_12420_),
    .A(net2992),
    .B(net6471));
 sg13g2_nand2_1 _43111_ (.Y(_12421_),
    .A(net5733),
    .B(_09813_));
 sg13g2_a21oi_2 _43112_ (.B1(_09915_),
    .Y(_12422_),
    .A2(_09902_),
    .A1(_09662_));
 sg13g2_xnor2_1 _43113_ (.Y(_12423_),
    .A(_09815_),
    .B(_12422_));
 sg13g2_o21ai_1 _43114_ (.B1(_12421_),
    .Y(_12424_),
    .A1(net5733),
    .A2(_12423_));
 sg13g2_nand2_1 _43115_ (.Y(_12425_),
    .A(net5422),
    .B(_12424_));
 sg13g2_xnor2_1 _43116_ (.Y(_12426_),
    .A(net5469),
    .B(_12424_));
 sg13g2_nand2_1 _43117_ (.Y(_12427_),
    .A(_12410_),
    .B(_12415_));
 sg13g2_xnor2_1 _43118_ (.Y(_12428_),
    .A(_12426_),
    .B(_12427_));
 sg13g2_o21ai_1 _43119_ (.B1(net5967),
    .Y(_12429_),
    .A1(net5543),
    .A2(_12424_));
 sg13g2_a21oi_1 _43120_ (.A1(net5543),
    .A2(_12428_),
    .Y(_12430_),
    .B1(_12429_));
 sg13g2_a221oi_1 _43121_ (.B2(net5913),
    .C1(_12430_),
    .B1(_12408_),
    .A1(net5998),
    .Y(_12431_),
    .A2(_09857_));
 sg13g2_and2_1 _43122_ (.A(net5301),
    .B(_12431_),
    .X(_12432_));
 sg13g2_o21ai_1 _43123_ (.B1(net6887),
    .Y(_12433_),
    .A1(net5301),
    .A2(_09857_));
 sg13g2_o21ai_1 _43124_ (.B1(_12420_),
    .Y(_00839_),
    .A1(_12432_),
    .A2(_12433_));
 sg13g2_nor2_1 _43125_ (.A(net5769),
    .B(_09805_),
    .Y(_12434_));
 sg13g2_o21ai_1 _43126_ (.B1(_09814_),
    .Y(_12435_),
    .A1(_09815_),
    .A2(_12422_));
 sg13g2_xnor2_1 _43127_ (.Y(_12436_),
    .A(_09810_),
    .B(_12435_));
 sg13g2_a21oi_1 _43128_ (.A1(net5769),
    .A2(_12436_),
    .Y(_12437_),
    .B1(_12434_));
 sg13g2_a21o_2 _43129_ (.A2(_12436_),
    .A1(net5769),
    .B1(_12434_),
    .X(_12438_));
 sg13g2_xnor2_1 _43130_ (.Y(_12439_),
    .A(net5427),
    .B(_12437_));
 sg13g2_nor2_1 _43131_ (.A(_12381_),
    .B(_12397_),
    .Y(_12440_));
 sg13g2_nand4_1 _43132_ (.B(_12411_),
    .C(_12426_),
    .A(_12384_),
    .Y(_12441_),
    .D(_12440_));
 sg13g2_nand3_1 _43133_ (.B(_12412_),
    .C(_12426_),
    .A(_12411_),
    .Y(_12442_));
 sg13g2_nand4_1 _43134_ (.B(_12425_),
    .C(_12441_),
    .A(_12410_),
    .Y(_12443_),
    .D(_12442_));
 sg13g2_and4_1 _43135_ (.A(_12385_),
    .B(_12411_),
    .C(_12426_),
    .D(_12440_),
    .X(_12444_));
 sg13g2_a21oi_2 _43136_ (.B1(_12443_),
    .Y(_12445_),
    .A2(_12444_),
    .A1(_12323_));
 sg13g2_nand2b_1 _43137_ (.Y(_12446_),
    .B(_12439_),
    .A_N(_12445_));
 sg13g2_xor2_1 _43138_ (.B(_12445_),
    .A(_12439_),
    .X(_12447_));
 sg13g2_o21ai_1 _43139_ (.B1(net5967),
    .Y(_12448_),
    .A1(net5542),
    .A2(_12438_));
 sg13g2_a21oi_1 _43140_ (.A1(net5542),
    .A2(_12447_),
    .Y(_12449_),
    .B1(_12448_));
 sg13g2_a221oi_1 _43141_ (.B2(net5913),
    .C1(_12449_),
    .B1(_12424_),
    .A1(net5998),
    .Y(_12450_),
    .A2(_09848_));
 sg13g2_o21ai_1 _43142_ (.B1(net6887),
    .Y(_12451_),
    .A1(net5299),
    .A2(_09848_));
 sg13g2_a21oi_1 _43143_ (.A1(net5299),
    .A2(_12450_),
    .Y(_12452_),
    .B1(_12451_));
 sg13g2_a21o_1 _43144_ (.A2(net6472),
    .A1(net3342),
    .B1(_12452_),
    .X(_00840_));
 sg13g2_o21ai_1 _43145_ (.B1(_12446_),
    .Y(_12453_),
    .A1(net5472),
    .A2(_12437_));
 sg13g2_nor2_1 _43146_ (.A(net5769),
    .B(_09797_),
    .Y(_12454_));
 sg13g2_a21oi_1 _43147_ (.A1(_09809_),
    .A2(_12435_),
    .Y(_12455_),
    .B1(_09807_));
 sg13g2_xnor2_1 _43148_ (.Y(_12456_),
    .A(_09800_),
    .B(_12455_));
 sg13g2_a21oi_2 _43149_ (.B1(_12454_),
    .Y(_12457_),
    .A2(_12456_),
    .A1(net5769));
 sg13g2_nor2_1 _43150_ (.A(net5427),
    .B(_12457_),
    .Y(_12458_));
 sg13g2_xnor2_1 _43151_ (.Y(_12459_),
    .A(net5472),
    .B(_12457_));
 sg13g2_xnor2_1 _43152_ (.Y(_12460_),
    .A(_12453_),
    .B(_12459_));
 sg13g2_o21ai_1 _43153_ (.B1(net5966),
    .Y(_12461_),
    .A1(net5542),
    .A2(_12457_));
 sg13g2_a21oi_1 _43154_ (.A1(net5542),
    .A2(_12460_),
    .Y(_12462_),
    .B1(_12461_));
 sg13g2_a221oi_1 _43155_ (.B2(net5913),
    .C1(_12462_),
    .B1(_12438_),
    .A1(net5999),
    .Y(_12463_),
    .A2(_09813_));
 sg13g2_a21oi_1 _43156_ (.A1(net5299),
    .A2(_12463_),
    .Y(_12464_),
    .B1(net6861));
 sg13g2_o21ai_1 _43157_ (.B1(_12464_),
    .Y(_12465_),
    .A1(net5299),
    .A2(_09813_));
 sg13g2_o21ai_1 _43158_ (.B1(_12465_),
    .Y(_00841_),
    .A1(_18146_),
    .A2(net6508));
 sg13g2_nand2_1 _43159_ (.Y(_12466_),
    .A(net5733),
    .B(_09787_));
 sg13g2_o21ai_1 _43160_ (.B1(_09798_),
    .Y(_12467_),
    .A1(_09800_),
    .A2(_12455_));
 sg13g2_xnor2_1 _43161_ (.Y(_12468_),
    .A(_09788_),
    .B(_12467_));
 sg13g2_o21ai_1 _43162_ (.B1(_12466_),
    .Y(_12469_),
    .A1(net5734),
    .A2(_12468_));
 sg13g2_nor2_1 _43163_ (.A(net5542),
    .B(_12469_),
    .Y(_12470_));
 sg13g2_nand2_1 _43164_ (.Y(_12471_),
    .A(net5428),
    .B(_12469_));
 sg13g2_xnor2_1 _43165_ (.Y(_12472_),
    .A(net5472),
    .B(_12469_));
 sg13g2_o21ai_1 _43166_ (.B1(net5428),
    .Y(_12473_),
    .A1(_12438_),
    .A2(_12457_));
 sg13g2_a21oi_1 _43167_ (.A1(_12446_),
    .A2(_12473_),
    .Y(_12474_),
    .B1(_12458_));
 sg13g2_nand2_1 _43168_ (.Y(_12475_),
    .A(_12472_),
    .B(_12474_));
 sg13g2_xnor2_1 _43169_ (.Y(_12476_),
    .A(_12472_),
    .B(_12474_));
 sg13g2_a21oi_1 _43170_ (.A1(net5542),
    .A2(_12476_),
    .Y(_12477_),
    .B1(_12470_));
 sg13g2_a22oi_1 _43171_ (.Y(_12478_),
    .B1(_12477_),
    .B2(net5230),
    .A2(_12457_),
    .A1(net5220));
 sg13g2_a22oi_1 _43172_ (.Y(_12479_),
    .B1(net5109),
    .B2(_09806_),
    .A2(net6471),
    .A1(net2986));
 sg13g2_o21ai_1 _43173_ (.B1(_12479_),
    .Y(_00842_),
    .A1(net6861),
    .A2(_12478_));
 sg13g2_o21ai_1 _43174_ (.B1(_09922_),
    .Y(_12480_),
    .A1(_09817_),
    .A2(_12422_));
 sg13g2_nand2_1 _43175_ (.Y(_12481_),
    .A(_09842_),
    .B(_12480_));
 sg13g2_nor2_1 _43176_ (.A(_09842_),
    .B(_12480_),
    .Y(_12482_));
 sg13g2_nor2_1 _43177_ (.A(net5733),
    .B(_12482_),
    .Y(_12483_));
 sg13g2_a22oi_1 _43178_ (.Y(_12484_),
    .B1(_12481_),
    .B2(_12483_),
    .A2(_09839_),
    .A1(net5733));
 sg13g2_inv_1 _43179_ (.Y(_12485_),
    .A(_12484_));
 sg13g2_nand2_1 _43180_ (.Y(_12486_),
    .A(net5428),
    .B(_12485_));
 sg13g2_xnor2_1 _43181_ (.Y(_12487_),
    .A(net5428),
    .B(_12484_));
 sg13g2_nand2_1 _43182_ (.Y(_12488_),
    .A(_12471_),
    .B(_12475_));
 sg13g2_xor2_1 _43183_ (.B(_12488_),
    .A(_12487_),
    .X(_12489_));
 sg13g2_a21oi_1 _43184_ (.A1(net5568),
    .A2(_12484_),
    .Y(_12490_),
    .B1(net5932));
 sg13g2_o21ai_1 _43185_ (.B1(_12490_),
    .Y(_12491_),
    .A1(net5568),
    .A2(_12489_));
 sg13g2_a22oi_1 _43186_ (.Y(_12492_),
    .B1(_12469_),
    .B2(net5914),
    .A2(_09797_),
    .A1(net5999));
 sg13g2_nand3_1 _43187_ (.B(_12491_),
    .C(_12492_),
    .A(net5299),
    .Y(_12493_));
 sg13g2_o21ai_1 _43188_ (.B1(net6886),
    .Y(_12494_),
    .A1(net5299),
    .A2(_09797_));
 sg13g2_nand2b_1 _43189_ (.Y(_12495_),
    .B(_12493_),
    .A_N(_12494_));
 sg13g2_o21ai_1 _43190_ (.B1(_12495_),
    .Y(_00843_),
    .A1(_18144_),
    .A2(net6509));
 sg13g2_a21oi_1 _43191_ (.A1(_09842_),
    .A2(_12480_),
    .Y(_12496_),
    .B1(_09840_));
 sg13g2_xnor2_1 _43192_ (.Y(_12497_),
    .A(_09835_),
    .B(_12496_));
 sg13g2_or2_1 _43193_ (.X(_12498_),
    .B(_09833_),
    .A(net5768));
 sg13g2_o21ai_1 _43194_ (.B1(_12498_),
    .Y(_12499_),
    .A1(net5733),
    .A2(_12497_));
 sg13g2_nand2_1 _43195_ (.Y(_12500_),
    .A(net5427),
    .B(_12499_));
 sg13g2_xnor2_1 _43196_ (.Y(_12501_),
    .A(net5427),
    .B(_12499_));
 sg13g2_nand3b_1 _43197_ (.B(_12487_),
    .C(_12472_),
    .Y(_12502_),
    .A_N(_12473_));
 sg13g2_nand3_1 _43198_ (.B(_12486_),
    .C(_12502_),
    .A(_12471_),
    .Y(_12503_));
 sg13g2_and4_1 _43199_ (.A(_12439_),
    .B(_12459_),
    .C(_12472_),
    .D(_12487_),
    .X(_12504_));
 sg13g2_nand2b_1 _43200_ (.Y(_12505_),
    .B(_12504_),
    .A_N(_12445_));
 sg13g2_nand2b_1 _43201_ (.Y(_12506_),
    .B(_12505_),
    .A_N(_12503_));
 sg13g2_nand2b_1 _43202_ (.Y(_12507_),
    .B(_12506_),
    .A_N(_12501_));
 sg13g2_xor2_1 _43203_ (.B(_12506_),
    .A(_12501_),
    .X(_12508_));
 sg13g2_o21ai_1 _43204_ (.B1(net5966),
    .Y(_12509_),
    .A1(net5543),
    .A2(_12499_));
 sg13g2_a21oi_1 _43205_ (.A1(net5543),
    .A2(_12508_),
    .Y(_12510_),
    .B1(_12509_));
 sg13g2_a221oi_1 _43206_ (.B2(net5913),
    .C1(_12510_),
    .B1(_12485_),
    .A1(net5999),
    .Y(_12511_),
    .A2(_09787_));
 sg13g2_a21oi_1 _43207_ (.A1(net5300),
    .A2(_12511_),
    .Y(_12512_),
    .B1(net6861));
 sg13g2_o21ai_1 _43208_ (.B1(_12512_),
    .Y(_12513_),
    .A1(net5299),
    .A2(_09787_));
 sg13g2_o21ai_1 _43209_ (.B1(_12513_),
    .Y(_00844_),
    .A1(_18143_),
    .A2(net6508));
 sg13g2_a22oi_1 _43210_ (.Y(_12514_),
    .B1(_09916_),
    .B2(_12481_),
    .A2(_09833_),
    .A1(net5605));
 sg13g2_a221oi_1 _43211_ (.B2(_12481_),
    .C1(_09830_),
    .B1(_09916_),
    .A1(net5605),
    .Y(_12515_),
    .A2(_09833_));
 sg13g2_xnor2_1 _43212_ (.Y(_12516_),
    .A(_09830_),
    .B(_12514_));
 sg13g2_mux2_1 _43213_ (.A0(_09828_),
    .A1(_12516_),
    .S(net5769),
    .X(_12517_));
 sg13g2_nor2_1 _43214_ (.A(net5427),
    .B(_12517_),
    .Y(_12518_));
 sg13g2_nand2_1 _43215_ (.Y(_12519_),
    .A(net5427),
    .B(_12517_));
 sg13g2_xnor2_1 _43216_ (.Y(_12520_),
    .A(net5427),
    .B(_12517_));
 sg13g2_nand2_1 _43217_ (.Y(_12521_),
    .A(_12500_),
    .B(_12507_));
 sg13g2_xor2_1 _43218_ (.B(_12521_),
    .A(_12520_),
    .X(_12522_));
 sg13g2_o21ai_1 _43219_ (.B1(net5966),
    .Y(_12523_),
    .A1(net5542),
    .A2(_12517_));
 sg13g2_a21oi_1 _43220_ (.A1(net5542),
    .A2(_12522_),
    .Y(_12524_),
    .B1(_12523_));
 sg13g2_a221oi_1 _43221_ (.B2(net5913),
    .C1(_12524_),
    .B1(_12499_),
    .A1(net5999),
    .Y(_12525_),
    .A2(_09839_));
 sg13g2_o21ai_1 _43222_ (.B1(net6887),
    .Y(_12526_),
    .A1(net5300),
    .A2(_09839_));
 sg13g2_a21oi_1 _43223_ (.A1(net5300),
    .A2(_12525_),
    .Y(_12527_),
    .B1(_12526_));
 sg13g2_a21o_1 _43224_ (.A2(net6472),
    .A1(net3321),
    .B1(_12527_),
    .X(_00845_));
 sg13g2_nor2_1 _43225_ (.A(_09829_),
    .B(_12515_),
    .Y(_12528_));
 sg13g2_xor2_1 _43226_ (.B(_12528_),
    .A(_09823_),
    .X(_12529_));
 sg13g2_nand2_1 _43227_ (.Y(_12530_),
    .A(net5733),
    .B(_09821_));
 sg13g2_o21ai_1 _43228_ (.B1(_12530_),
    .Y(_12531_),
    .A1(net5733),
    .A2(_12529_));
 sg13g2_inv_1 _43229_ (.Y(_12532_),
    .A(_12531_));
 sg13g2_nor2_1 _43230_ (.A(net5472),
    .B(_12531_),
    .Y(_12533_));
 sg13g2_xnor2_1 _43231_ (.Y(_12534_),
    .A(net5472),
    .B(_12531_));
 sg13g2_nand2_1 _43232_ (.Y(_12535_),
    .A(_12500_),
    .B(_12519_));
 sg13g2_nor2b_1 _43233_ (.A(_12535_),
    .B_N(_12507_),
    .Y(_12536_));
 sg13g2_or3_1 _43234_ (.A(_12518_),
    .B(_12534_),
    .C(_12536_),
    .X(_12537_));
 sg13g2_o21ai_1 _43235_ (.B1(_12534_),
    .Y(_12538_),
    .A1(_12518_),
    .A2(_12536_));
 sg13g2_a21oi_1 _43236_ (.A1(_12537_),
    .A2(_12538_),
    .Y(_12539_),
    .B1(net5568));
 sg13g2_a21oi_1 _43237_ (.A1(net5568),
    .A2(_12531_),
    .Y(_12540_),
    .B1(_12539_));
 sg13g2_nor2_1 _43238_ (.A(net6007),
    .B(_09833_),
    .Y(_12541_));
 sg13g2_a221oi_1 _43239_ (.B2(net5966),
    .C1(_12541_),
    .B1(_12540_),
    .A1(net5913),
    .Y(_12542_),
    .A2(_12517_));
 sg13g2_nand3_1 _43240_ (.B(net5318),
    .C(_09833_),
    .A(net5322),
    .Y(_12543_));
 sg13g2_nand2_1 _43241_ (.Y(_12544_),
    .A(net6887),
    .B(_12543_));
 sg13g2_a21o_1 _43242_ (.A2(_12542_),
    .A1(net5301),
    .B1(_12544_),
    .X(_12545_));
 sg13g2_o21ai_1 _43243_ (.B1(_12545_),
    .Y(_00846_),
    .A1(_18142_),
    .A2(net6508));
 sg13g2_nand2_1 _43244_ (.Y(_12546_),
    .A(net2134),
    .B(net6471));
 sg13g2_nand2_1 _43245_ (.Y(_12547_),
    .A(net5731),
    .B(_09772_));
 sg13g2_a21oi_2 _43246_ (.B1(_09904_),
    .Y(_12548_),
    .A2(_09661_),
    .A1(_09124_));
 sg13g2_nor2_1 _43247_ (.A(_09925_),
    .B(_12548_),
    .Y(_12549_));
 sg13g2_o21ai_1 _43248_ (.B1(_09775_),
    .Y(_12550_),
    .A1(_09925_),
    .A2(_12548_));
 sg13g2_xnor2_1 _43249_ (.Y(_12551_),
    .A(_09774_),
    .B(_12549_));
 sg13g2_o21ai_1 _43250_ (.B1(_12547_),
    .Y(_12552_),
    .A1(net5731),
    .A2(_12551_));
 sg13g2_xnor2_1 _43251_ (.Y(_12553_),
    .A(net5472),
    .B(_12552_));
 sg13g2_nand2b_1 _43252_ (.Y(_12554_),
    .B(_12537_),
    .A_N(_12533_));
 sg13g2_xnor2_1 _43253_ (.Y(_12555_),
    .A(_12553_),
    .B(_12554_));
 sg13g2_o21ai_1 _43254_ (.B1(net5966),
    .Y(_12556_),
    .A1(net5543),
    .A2(_12552_));
 sg13g2_a21oi_1 _43255_ (.A1(net5543),
    .A2(_12555_),
    .Y(_12557_),
    .B1(_12556_));
 sg13g2_a22oi_1 _43256_ (.Y(_12558_),
    .B1(_12532_),
    .B2(net5913),
    .A2(_09828_),
    .A1(net5998));
 sg13g2_nand2_1 _43257_ (.Y(_12559_),
    .A(net5299),
    .B(_12558_));
 sg13g2_nor2_1 _43258_ (.A(_12557_),
    .B(_12559_),
    .Y(_12560_));
 sg13g2_o21ai_1 _43259_ (.B1(net6887),
    .Y(_12561_),
    .A1(net5300),
    .A2(_09828_));
 sg13g2_o21ai_1 _43260_ (.B1(_12546_),
    .Y(_00847_),
    .A1(_12560_),
    .A2(_12561_));
 sg13g2_nand2_1 _43261_ (.Y(_12562_),
    .A(_09773_),
    .B(_12550_));
 sg13g2_xnor2_1 _43262_ (.Y(_12563_),
    .A(_09769_),
    .B(_12562_));
 sg13g2_nand2_1 _43263_ (.Y(_12564_),
    .A(net5726),
    .B(_09767_));
 sg13g2_o21ai_1 _43264_ (.B1(_12564_),
    .Y(_12565_),
    .A1(net5726),
    .A2(_12563_));
 sg13g2_nor2_1 _43265_ (.A(net5539),
    .B(_12565_),
    .Y(_12566_));
 sg13g2_nand2_1 _43266_ (.Y(_12567_),
    .A(net5419),
    .B(_12565_));
 sg13g2_xnor2_1 _43267_ (.Y(_12568_),
    .A(net5466),
    .B(_12565_));
 sg13g2_nor2b_2 _43268_ (.A(_12534_),
    .B_N(_12553_),
    .Y(_12569_));
 sg13g2_nor2_1 _43269_ (.A(_12501_),
    .B(_12520_),
    .Y(_12570_));
 sg13g2_nand4_1 _43270_ (.B(_12504_),
    .C(_12569_),
    .A(_12443_),
    .Y(_12571_),
    .D(_12570_));
 sg13g2_a221oi_1 _43271_ (.B2(_12535_),
    .C1(_12533_),
    .B1(_12569_),
    .A1(net5427),
    .Y(_12572_),
    .A2(_12552_));
 sg13g2_nand3_1 _43272_ (.B(_12569_),
    .C(_12570_),
    .A(_12503_),
    .Y(_12573_));
 sg13g2_nand3_1 _43273_ (.B(_12572_),
    .C(_12573_),
    .A(_12571_),
    .Y(_12574_));
 sg13g2_and4_1 _43274_ (.A(_12444_),
    .B(_12504_),
    .C(_12569_),
    .D(_12570_),
    .X(_12575_));
 sg13g2_a21oi_2 _43275_ (.B1(_12574_),
    .Y(_12576_),
    .A2(_12575_),
    .A1(_12323_));
 sg13g2_nand2b_1 _43276_ (.Y(_12577_),
    .B(_12568_),
    .A_N(_12576_));
 sg13g2_xor2_1 _43277_ (.B(_12576_),
    .A(_12568_),
    .X(_12578_));
 sg13g2_a21oi_1 _43278_ (.A1(net5539),
    .A2(_12578_),
    .Y(_12579_),
    .B1(_12566_));
 sg13g2_a22oi_1 _43279_ (.Y(_12580_),
    .B1(_12579_),
    .B2(net5230),
    .A2(_12552_),
    .A1(net5218));
 sg13g2_nor2_1 _43280_ (.A(net5065),
    .B(_09821_),
    .Y(_12581_));
 sg13g2_a21oi_1 _43281_ (.A1(net3739),
    .A2(net6471),
    .Y(_12582_),
    .B1(_12581_));
 sg13g2_o21ai_1 _43282_ (.B1(_12582_),
    .Y(_00848_),
    .A1(net6862),
    .A2(_12580_));
 sg13g2_nand2_1 _43283_ (.Y(_12583_),
    .A(net3327),
    .B(net6468));
 sg13g2_nor2_1 _43284_ (.A(net5295),
    .B(_09772_),
    .Y(_12584_));
 sg13g2_nand2_1 _43285_ (.Y(_12585_),
    .A(_12567_),
    .B(_12577_));
 sg13g2_a21oi_1 _43286_ (.A1(_09927_),
    .A2(_12550_),
    .Y(_12586_),
    .B1(_09768_));
 sg13g2_xnor2_1 _43287_ (.Y(_12587_),
    .A(_09764_),
    .B(_12586_));
 sg13g2_nand2_1 _43288_ (.Y(_12588_),
    .A(net5765),
    .B(_12587_));
 sg13g2_o21ai_1 _43289_ (.B1(_12588_),
    .Y(_12589_),
    .A1(net5766),
    .A2(_09762_));
 sg13g2_nor2_1 _43290_ (.A(net5466),
    .B(_12589_),
    .Y(_12590_));
 sg13g2_xnor2_1 _43291_ (.Y(_12591_),
    .A(net5419),
    .B(_12589_));
 sg13g2_xor2_1 _43292_ (.B(_12591_),
    .A(_12585_),
    .X(_12592_));
 sg13g2_a21oi_1 _43293_ (.A1(net5565),
    .A2(_12589_),
    .Y(_12593_),
    .B1(net5932));
 sg13g2_o21ai_1 _43294_ (.B1(_12593_),
    .Y(_12594_),
    .A1(net5566),
    .A2(_12592_));
 sg13g2_a22oi_1 _43295_ (.Y(_12595_),
    .B1(_12565_),
    .B2(net5910),
    .A2(_09772_),
    .A1(net5995));
 sg13g2_nand3_1 _43296_ (.B(_12594_),
    .C(_12595_),
    .A(net5295),
    .Y(_12596_));
 sg13g2_nand2_1 _43297_ (.Y(_12597_),
    .A(net6885),
    .B(_12596_));
 sg13g2_o21ai_1 _43298_ (.B1(_12583_),
    .Y(_00849_),
    .A1(_12584_),
    .A2(_12597_));
 sg13g2_a21oi_1 _43299_ (.A1(_09764_),
    .A2(_12586_),
    .Y(_12598_),
    .B1(_09763_));
 sg13g2_xor2_1 _43300_ (.B(_12598_),
    .A(_09755_),
    .X(_12599_));
 sg13g2_nor2_1 _43301_ (.A(net5726),
    .B(_12599_),
    .Y(_12600_));
 sg13g2_a21oi_2 _43302_ (.B1(_12600_),
    .Y(_12601_),
    .A2(_09754_),
    .A1(net5726));
 sg13g2_inv_1 _43303_ (.Y(_12602_),
    .A(_12601_));
 sg13g2_nor2_1 _43304_ (.A(net5535),
    .B(_12602_),
    .Y(_12603_));
 sg13g2_nor2_1 _43305_ (.A(net5466),
    .B(_12601_),
    .Y(_12604_));
 sg13g2_xnor2_1 _43306_ (.Y(_12605_),
    .A(net5419),
    .B(_12601_));
 sg13g2_a21oi_1 _43307_ (.A1(net5419),
    .A2(_12565_),
    .Y(_12606_),
    .B1(_12590_));
 sg13g2_a22oi_1 _43308_ (.Y(_12607_),
    .B1(_12606_),
    .B2(_12577_),
    .A2(_12589_),
    .A1(net5466));
 sg13g2_xnor2_1 _43309_ (.Y(_12608_),
    .A(_12605_),
    .B(_12607_));
 sg13g2_a21oi_1 _43310_ (.A1(net5535),
    .A2(_12608_),
    .Y(_12609_),
    .B1(_12603_));
 sg13g2_a22oi_1 _43311_ (.Y(_12610_),
    .B1(_12609_),
    .B2(net5230),
    .A2(_09767_),
    .A1(net5167));
 sg13g2_o21ai_1 _43312_ (.B1(_12610_),
    .Y(_12611_),
    .A1(net5120),
    .A2(_12589_));
 sg13g2_a22oi_1 _43313_ (.Y(_12612_),
    .B1(net6885),
    .B2(_12611_),
    .A2(net6468),
    .A1(net3052));
 sg13g2_inv_1 _43314_ (.Y(_00850_),
    .A(_12612_));
 sg13g2_nand2_1 _43315_ (.Y(_12613_),
    .A(net3252),
    .B(net6468));
 sg13g2_o21ai_1 _43316_ (.B1(_09777_),
    .Y(_12614_),
    .A1(_09925_),
    .A2(_12548_));
 sg13g2_a21oi_1 _43317_ (.A1(_09930_),
    .A2(_12614_),
    .Y(_12615_),
    .B1(_09744_));
 sg13g2_nand3_1 _43318_ (.B(_09930_),
    .C(_12614_),
    .A(_09744_),
    .Y(_12616_));
 sg13g2_nand2b_1 _43319_ (.Y(_12617_),
    .B(_12616_),
    .A_N(_12615_));
 sg13g2_nor2_1 _43320_ (.A(net5726),
    .B(_12617_),
    .Y(_12618_));
 sg13g2_a21oi_2 _43321_ (.B1(_12618_),
    .Y(_12619_),
    .A2(_09742_),
    .A1(net5726));
 sg13g2_xnor2_1 _43322_ (.Y(_12620_),
    .A(net5420),
    .B(_12619_));
 sg13g2_a21oi_1 _43323_ (.A1(_12605_),
    .A2(_12607_),
    .Y(_12621_),
    .B1(_12604_));
 sg13g2_xnor2_1 _43324_ (.Y(_12622_),
    .A(_12620_),
    .B(_12621_));
 sg13g2_a21oi_1 _43325_ (.A1(net5566),
    .A2(_12619_),
    .Y(_12623_),
    .B1(net5931));
 sg13g2_o21ai_1 _43326_ (.B1(_12623_),
    .Y(_12624_),
    .A1(net5566),
    .A2(_12622_));
 sg13g2_a22oi_1 _43327_ (.Y(_12625_),
    .B1(_12602_),
    .B2(net5911),
    .A2(_09762_),
    .A1(net5996));
 sg13g2_and3_1 _43328_ (.X(_12626_),
    .A(net5291),
    .B(_12624_),
    .C(_12625_));
 sg13g2_o21ai_1 _43329_ (.B1(net6885),
    .Y(_12627_),
    .A1(net5291),
    .A2(_09762_));
 sg13g2_o21ai_1 _43330_ (.B1(_12613_),
    .Y(_00851_),
    .A1(_12626_),
    .A2(_12627_));
 sg13g2_or2_1 _43331_ (.X(_12628_),
    .B(_09748_),
    .A(net5766));
 sg13g2_nor2_1 _43332_ (.A(_09743_),
    .B(_12615_),
    .Y(_12629_));
 sg13g2_xnor2_1 _43333_ (.Y(_12630_),
    .A(_09751_),
    .B(_12629_));
 sg13g2_o21ai_1 _43334_ (.B1(_12628_),
    .Y(_12631_),
    .A1(net5727),
    .A2(_12630_));
 sg13g2_nand2_1 _43335_ (.Y(_12632_),
    .A(net5417),
    .B(_12631_));
 sg13g2_inv_1 _43336_ (.Y(_12633_),
    .A(_12632_));
 sg13g2_xnor2_1 _43337_ (.Y(_12634_),
    .A(net5467),
    .B(_12631_));
 sg13g2_inv_1 _43338_ (.Y(_12635_),
    .A(_12634_));
 sg13g2_nand3b_1 _43339_ (.B(_12620_),
    .C(_12605_),
    .Y(_12636_),
    .A_N(_12606_));
 sg13g2_a21o_1 _43340_ (.A2(_12619_),
    .A1(_12601_),
    .B1(net5466),
    .X(_12637_));
 sg13g2_and2_1 _43341_ (.A(_12636_),
    .B(_12637_),
    .X(_12638_));
 sg13g2_and4_1 _43342_ (.A(_12568_),
    .B(_12591_),
    .C(_12605_),
    .D(_12620_),
    .X(_12639_));
 sg13g2_inv_1 _43343_ (.Y(_12640_),
    .A(_12639_));
 sg13g2_o21ai_1 _43344_ (.B1(_12638_),
    .Y(_12641_),
    .A1(_12576_),
    .A2(_12640_));
 sg13g2_and2_1 _43345_ (.A(_12634_),
    .B(_12641_),
    .X(_12642_));
 sg13g2_xnor2_1 _43346_ (.Y(_12643_),
    .A(_12634_),
    .B(_12641_));
 sg13g2_nor2_1 _43347_ (.A(net5533),
    .B(_12631_),
    .Y(_12644_));
 sg13g2_a21oi_1 _43348_ (.A1(net5535),
    .A2(_12643_),
    .Y(_12645_),
    .B1(_12644_));
 sg13g2_nand2_1 _43349_ (.Y(_12646_),
    .A(net5232),
    .B(_12645_));
 sg13g2_o21ai_1 _43350_ (.B1(_12646_),
    .Y(_12647_),
    .A1(net5121),
    .A2(_12619_));
 sg13g2_a22oi_1 _43351_ (.Y(_12648_),
    .B1(_12647_),
    .B2(net6889),
    .A2(_09754_),
    .A1(net5108));
 sg13g2_o21ai_1 _43352_ (.B1(_12648_),
    .Y(_00852_),
    .A1(_18140_),
    .A2(net6504));
 sg13g2_nor2_1 _43353_ (.A(net5766),
    .B(_09736_),
    .Y(_12649_));
 sg13g2_o21ai_1 _43354_ (.B1(_09750_),
    .Y(_12650_),
    .A1(_09934_),
    .A2(_12615_));
 sg13g2_xnor2_1 _43355_ (.Y(_12651_),
    .A(_09738_),
    .B(_12650_));
 sg13g2_a21oi_2 _43356_ (.B1(_12649_),
    .Y(_12652_),
    .A2(_12651_),
    .A1(net5766));
 sg13g2_nor2_1 _43357_ (.A(net5417),
    .B(_12652_),
    .Y(_12653_));
 sg13g2_xnor2_1 _43358_ (.Y(_12654_),
    .A(net5417),
    .B(_12652_));
 sg13g2_nor2_1 _43359_ (.A(_12633_),
    .B(_12642_),
    .Y(_12655_));
 sg13g2_xnor2_1 _43360_ (.Y(_12656_),
    .A(_12654_),
    .B(_12655_));
 sg13g2_o21ai_1 _43361_ (.B1(net5968),
    .Y(_12657_),
    .A1(net5533),
    .A2(_12652_));
 sg13g2_a21oi_1 _43362_ (.A1(net5532),
    .A2(_12656_),
    .Y(_12658_),
    .B1(_12657_));
 sg13g2_a221oi_1 _43363_ (.B2(net5909),
    .C1(_12658_),
    .B1(_12631_),
    .A1(net5994),
    .Y(_12659_),
    .A2(_09742_));
 sg13g2_o21ai_1 _43364_ (.B1(net6889),
    .Y(_12660_),
    .A1(net5291),
    .A2(_09742_));
 sg13g2_a21oi_1 _43365_ (.A1(net5291),
    .A2(_12659_),
    .Y(_12661_),
    .B1(_12660_));
 sg13g2_a21o_1 _43366_ (.A2(net6454),
    .A1(net2980),
    .B1(_12661_),
    .X(_00853_));
 sg13g2_o21ai_1 _43367_ (.B1(_09737_),
    .Y(_12662_),
    .A1(_09738_),
    .A2(_12650_));
 sg13g2_xnor2_1 _43368_ (.Y(_12663_),
    .A(_09725_),
    .B(_12662_));
 sg13g2_nand2_1 _43369_ (.Y(_12664_),
    .A(net5724),
    .B(_09724_));
 sg13g2_o21ai_1 _43370_ (.B1(_12664_),
    .Y(_12665_),
    .A1(net5724),
    .A2(_12663_));
 sg13g2_nand2_1 _43371_ (.Y(_12666_),
    .A(net5420),
    .B(_12665_));
 sg13g2_xnor2_1 _43372_ (.Y(_12667_),
    .A(net5467),
    .B(_12665_));
 sg13g2_a21o_1 _43373_ (.A2(_12652_),
    .A1(net5420),
    .B1(_12633_),
    .X(_12668_));
 sg13g2_nor2_1 _43374_ (.A(_12642_),
    .B(_12668_),
    .Y(_12669_));
 sg13g2_nor2_1 _43375_ (.A(_12653_),
    .B(_12669_),
    .Y(_12670_));
 sg13g2_nand2_1 _43376_ (.Y(_12671_),
    .A(_12667_),
    .B(_12670_));
 sg13g2_xnor2_1 _43377_ (.Y(_12672_),
    .A(_12667_),
    .B(_12670_));
 sg13g2_nor2_1 _43378_ (.A(net5533),
    .B(_12665_),
    .Y(_12673_));
 sg13g2_a21oi_1 _43379_ (.A1(net5533),
    .A2(_12672_),
    .Y(_12674_),
    .B1(_12673_));
 sg13g2_a22oi_1 _43380_ (.Y(_12675_),
    .B1(_12674_),
    .B2(net5232),
    .A2(_12652_),
    .A1(net5217));
 sg13g2_nor2_1 _43381_ (.A(net6859),
    .B(_12675_),
    .Y(_12676_));
 sg13g2_a21oi_1 _43382_ (.A1(net2877),
    .A2(net6455),
    .Y(_12677_),
    .B1(_12676_));
 sg13g2_o21ai_1 _43383_ (.B1(_12677_),
    .Y(_00854_),
    .A1(_02375_),
    .A2(_09748_));
 sg13g2_nand2_1 _43384_ (.Y(_12678_),
    .A(net2361),
    .B(net6455));
 sg13g2_o21ai_1 _43385_ (.B1(_09778_),
    .Y(_12679_),
    .A1(_09925_),
    .A2(_12548_));
 sg13g2_nand2_2 _43386_ (.Y(_12680_),
    .A(_09936_),
    .B(_12679_));
 sg13g2_a21oi_1 _43387_ (.A1(_09936_),
    .A2(_12679_),
    .Y(_12681_),
    .B1(_09693_));
 sg13g2_o21ai_1 _43388_ (.B1(net5766),
    .Y(_12682_),
    .A1(_09692_),
    .A2(_12680_));
 sg13g2_nor2_1 _43389_ (.A(_12681_),
    .B(_12682_),
    .Y(_12683_));
 sg13g2_a21oi_2 _43390_ (.B1(_12683_),
    .Y(_12684_),
    .A2(_09690_),
    .A1(net5724));
 sg13g2_inv_1 _43391_ (.Y(_12685_),
    .A(_12684_));
 sg13g2_xnor2_1 _43392_ (.Y(_12686_),
    .A(net5417),
    .B(_12684_));
 sg13g2_nand2_1 _43393_ (.Y(_12687_),
    .A(_12666_),
    .B(_12671_));
 sg13g2_xor2_1 _43394_ (.B(_12687_),
    .A(_12686_),
    .X(_12688_));
 sg13g2_a21oi_1 _43395_ (.A1(net5566),
    .A2(_12684_),
    .Y(_12689_),
    .B1(net5931));
 sg13g2_o21ai_1 _43396_ (.B1(_12689_),
    .Y(_12690_),
    .A1(net5566),
    .A2(_12688_));
 sg13g2_a22oi_1 _43397_ (.Y(_12691_),
    .B1(_12665_),
    .B2(net5909),
    .A2(_09736_),
    .A1(net5994));
 sg13g2_and3_1 _43398_ (.X(_12692_),
    .A(net5291),
    .B(_12690_),
    .C(_12691_));
 sg13g2_o21ai_1 _43399_ (.B1(net6889),
    .Y(_12693_),
    .A1(net5291),
    .A2(_09736_));
 sg13g2_o21ai_1 _43400_ (.B1(_12678_),
    .Y(_00855_),
    .A1(_12692_),
    .A2(_12693_));
 sg13g2_nand2_1 _43401_ (.Y(_12694_),
    .A(net5724),
    .B(_09684_));
 sg13g2_nor2_1 _43402_ (.A(_09691_),
    .B(_12681_),
    .Y(_12695_));
 sg13g2_xor2_1 _43403_ (.B(_12695_),
    .A(_09686_),
    .X(_12696_));
 sg13g2_o21ai_1 _43404_ (.B1(_12694_),
    .Y(_12697_),
    .A1(net5724),
    .A2(_12696_));
 sg13g2_nand2_1 _43405_ (.Y(_12698_),
    .A(net5417),
    .B(_12697_));
 sg13g2_inv_1 _43406_ (.Y(_12699_),
    .A(_12698_));
 sg13g2_xnor2_1 _43407_ (.Y(_12700_),
    .A(net5467),
    .B(_12697_));
 sg13g2_nand2_1 _43408_ (.Y(_12701_),
    .A(_12667_),
    .B(_12686_));
 sg13g2_nor3_1 _43409_ (.A(_12635_),
    .B(_12654_),
    .C(_12701_),
    .Y(_12702_));
 sg13g2_nor2b_1 _43410_ (.A(_12638_),
    .B_N(_12702_),
    .Y(_12703_));
 sg13g2_nor2b_1 _43411_ (.A(_12701_),
    .B_N(_12668_),
    .Y(_12704_));
 sg13g2_o21ai_1 _43412_ (.B1(_12666_),
    .Y(_12705_),
    .A1(net5467),
    .A2(_12684_));
 sg13g2_nor3_1 _43413_ (.A(_12703_),
    .B(_12704_),
    .C(_12705_),
    .Y(_12706_));
 sg13g2_and2_1 _43414_ (.A(_12639_),
    .B(_12702_),
    .X(_12707_));
 sg13g2_inv_1 _43415_ (.Y(_12708_),
    .A(_12707_));
 sg13g2_o21ai_1 _43416_ (.B1(_12706_),
    .Y(_12709_),
    .A1(_12576_),
    .A2(_12708_));
 sg13g2_and2_1 _43417_ (.A(_12700_),
    .B(_12709_),
    .X(_12710_));
 sg13g2_xnor2_1 _43418_ (.Y(_12711_),
    .A(_12700_),
    .B(_12709_));
 sg13g2_nor2_1 _43419_ (.A(net5532),
    .B(_12697_),
    .Y(_12712_));
 sg13g2_a21oi_1 _43420_ (.A1(net5532),
    .A2(_12711_),
    .Y(_12713_),
    .B1(_12712_));
 sg13g2_a22oi_1 _43421_ (.Y(_12714_),
    .B1(_12713_),
    .B2(net5232),
    .A2(_12685_),
    .A1(net5217));
 sg13g2_a22oi_1 _43422_ (.Y(_12715_),
    .B1(net5108),
    .B2(_09724_),
    .A2(net6455),
    .A1(net2890));
 sg13g2_o21ai_1 _43423_ (.B1(_12715_),
    .Y(_00856_),
    .A1(net6859),
    .A2(_12714_));
 sg13g2_nor2_1 _43424_ (.A(net5766),
    .B(_09672_),
    .Y(_12716_));
 sg13g2_o21ai_1 _43425_ (.B1(_09685_),
    .Y(_12717_),
    .A1(_09940_),
    .A2(_12681_));
 sg13g2_xnor2_1 _43426_ (.Y(_12718_),
    .A(_09674_),
    .B(_12717_));
 sg13g2_a21oi_2 _43427_ (.B1(_12716_),
    .Y(_12719_),
    .A2(_12718_),
    .A1(net5766));
 sg13g2_nand2b_1 _43428_ (.Y(_12720_),
    .B(net5467),
    .A_N(_12719_));
 sg13g2_xnor2_1 _43429_ (.Y(_12721_),
    .A(net5467),
    .B(_12719_));
 sg13g2_nor2_1 _43430_ (.A(_12699_),
    .B(_12710_),
    .Y(_12722_));
 sg13g2_xor2_1 _43431_ (.B(_12722_),
    .A(_12721_),
    .X(_12723_));
 sg13g2_o21ai_1 _43432_ (.B1(net5961),
    .Y(_12724_),
    .A1(net5532),
    .A2(_12719_));
 sg13g2_a21oi_1 _43433_ (.A1(net5532),
    .A2(_12723_),
    .Y(_12725_),
    .B1(_12724_));
 sg13g2_a221oi_1 _43434_ (.B2(net5909),
    .C1(_12725_),
    .B1(_12697_),
    .A1(net5993),
    .Y(_12726_),
    .A2(_09690_));
 sg13g2_o21ai_1 _43435_ (.B1(net6889),
    .Y(_12727_),
    .A1(net5292),
    .A2(_09690_));
 sg13g2_a21oi_1 _43436_ (.A1(net5292),
    .A2(_12726_),
    .Y(_12728_),
    .B1(_12727_));
 sg13g2_a21o_1 _43437_ (.A2(net6454),
    .A1(net2225),
    .B1(_12728_),
    .X(_00857_));
 sg13g2_nand2_1 _43438_ (.Y(_12729_),
    .A(net5724),
    .B(_09679_));
 sg13g2_o21ai_1 _43439_ (.B1(_09673_),
    .Y(_12730_),
    .A1(_09674_),
    .A2(_12717_));
 sg13g2_xnor2_1 _43440_ (.Y(_12731_),
    .A(_09680_),
    .B(_12730_));
 sg13g2_o21ai_1 _43441_ (.B1(_12729_),
    .Y(_12732_),
    .A1(net5724),
    .A2(_12731_));
 sg13g2_nand2_1 _43442_ (.Y(_12733_),
    .A(net5417),
    .B(_12732_));
 sg13g2_xnor2_1 _43443_ (.Y(_12734_),
    .A(net5467),
    .B(_12732_));
 sg13g2_a21o_1 _43444_ (.A2(_12719_),
    .A1(net5417),
    .B1(_12699_),
    .X(_12735_));
 sg13g2_or2_1 _43445_ (.X(_12736_),
    .B(_12735_),
    .A(_12710_));
 sg13g2_nand2_1 _43446_ (.Y(_12737_),
    .A(_12720_),
    .B(_12736_));
 sg13g2_nand3_1 _43447_ (.B(_12734_),
    .C(_12736_),
    .A(_12720_),
    .Y(_12738_));
 sg13g2_xnor2_1 _43448_ (.Y(_12739_),
    .A(_12734_),
    .B(_12737_));
 sg13g2_mux2_1 _43449_ (.A0(_12732_),
    .A1(_12739_),
    .S(net5532),
    .X(_12740_));
 sg13g2_a22oi_1 _43450_ (.Y(_12741_),
    .B1(_12740_),
    .B2(net5232),
    .A2(_12719_),
    .A1(net5217));
 sg13g2_a22oi_1 _43451_ (.Y(_12742_),
    .B1(net5108),
    .B2(_09684_),
    .A2(net6454),
    .A1(net3128));
 sg13g2_o21ai_1 _43452_ (.B1(_12742_),
    .Y(_00858_),
    .A1(net6859),
    .A2(_12741_));
 sg13g2_nand2_1 _43453_ (.Y(_12743_),
    .A(net5724),
    .B(_09712_));
 sg13g2_a21oi_1 _43454_ (.A1(_09694_),
    .A2(_12680_),
    .Y(_12744_),
    .B1(_09942_));
 sg13g2_a21o_1 _43455_ (.A2(_12680_),
    .A1(_09694_),
    .B1(_09942_),
    .X(_12745_));
 sg13g2_xnor2_1 _43456_ (.Y(_12746_),
    .A(_09714_),
    .B(_12744_));
 sg13g2_o21ai_1 _43457_ (.B1(_12743_),
    .Y(_12747_),
    .A1(net5723),
    .A2(_12746_));
 sg13g2_xnor2_1 _43458_ (.Y(_12748_),
    .A(net5467),
    .B(_12747_));
 sg13g2_nand2_1 _43459_ (.Y(_12749_),
    .A(_12733_),
    .B(_12738_));
 sg13g2_xnor2_1 _43460_ (.Y(_12750_),
    .A(_12748_),
    .B(_12749_));
 sg13g2_o21ai_1 _43461_ (.B1(net5961),
    .Y(_12751_),
    .A1(net5532),
    .A2(_12747_));
 sg13g2_a21o_1 _43462_ (.A2(_12750_),
    .A1(net5532),
    .B1(_12751_),
    .X(_12752_));
 sg13g2_a22oi_1 _43463_ (.Y(_12753_),
    .B1(_12732_),
    .B2(net5909),
    .A2(_09672_),
    .A1(net5994));
 sg13g2_nand3_1 _43464_ (.B(_12752_),
    .C(_12753_),
    .A(net5289),
    .Y(_12754_));
 sg13g2_nor2_1 _43465_ (.A(net5289),
    .B(_09672_),
    .Y(_12755_));
 sg13g2_nor2_1 _43466_ (.A(net6864),
    .B(_12755_),
    .Y(_12756_));
 sg13g2_a22oi_1 _43467_ (.Y(_12757_),
    .B1(_12754_),
    .B2(_12756_),
    .A2(net6454),
    .A1(net3157));
 sg13g2_inv_1 _43468_ (.Y(_00859_),
    .A(_12757_));
 sg13g2_o21ai_1 _43469_ (.B1(_09713_),
    .Y(_12758_),
    .A1(_09714_),
    .A2(_12744_));
 sg13g2_o21ai_1 _43470_ (.B1(net5764),
    .Y(_12759_),
    .A1(_09719_),
    .A2(_12758_));
 sg13g2_a21oi_1 _43471_ (.A1(_09719_),
    .A2(_12758_),
    .Y(_12760_),
    .B1(_12759_));
 sg13g2_a21oi_2 _43472_ (.B1(_12760_),
    .Y(_12761_),
    .A2(_09717_),
    .A1(net5722));
 sg13g2_xnor2_1 _43473_ (.Y(_12762_),
    .A(net5463),
    .B(_12761_));
 sg13g2_and2_1 _43474_ (.A(_12734_),
    .B(_12748_),
    .X(_12763_));
 sg13g2_a22oi_1 _43475_ (.Y(_12764_),
    .B1(_12763_),
    .B2(_12735_),
    .A2(_12747_),
    .A1(net5417));
 sg13g2_nand2_1 _43476_ (.Y(_12765_),
    .A(_12733_),
    .B(_12764_));
 sg13g2_and3_1 _43477_ (.X(_12766_),
    .A(_12700_),
    .B(_12721_),
    .C(_12763_));
 sg13g2_nand3_1 _43478_ (.B(_12721_),
    .C(_12763_),
    .A(_12700_),
    .Y(_12767_));
 sg13g2_a21oi_1 _43479_ (.A1(_12709_),
    .A2(_12766_),
    .Y(_12768_),
    .B1(_12765_));
 sg13g2_or2_1 _43480_ (.X(_12769_),
    .B(_12768_),
    .A(_12762_));
 sg13g2_xor2_1 _43481_ (.B(_12768_),
    .A(_12762_),
    .X(_12770_));
 sg13g2_o21ai_1 _43482_ (.B1(net5961),
    .Y(_12771_),
    .A1(net5566),
    .A2(_12770_));
 sg13g2_a21oi_1 _43483_ (.A1(net5566),
    .A2(_12761_),
    .Y(_12772_),
    .B1(_12771_));
 sg13g2_a221oi_1 _43484_ (.B2(net5909),
    .C1(_12772_),
    .B1(_12747_),
    .A1(net5994),
    .Y(_12773_),
    .A2(_09679_));
 sg13g2_a21oi_1 _43485_ (.A1(net5289),
    .A2(_12773_),
    .Y(_12774_),
    .B1(net6859));
 sg13g2_o21ai_1 _43486_ (.B1(_12774_),
    .Y(_12775_),
    .A1(net5289),
    .A2(_09679_));
 sg13g2_o21ai_1 _43487_ (.B1(_12775_),
    .Y(_00860_),
    .A1(_18138_),
    .A2(net6504));
 sg13g2_nor2_1 _43488_ (.A(net5764),
    .B(_09700_),
    .Y(_12776_));
 sg13g2_a21o_1 _43489_ (.A2(_12745_),
    .A1(_09720_),
    .B1(_09938_),
    .X(_12777_));
 sg13g2_xor2_1 _43490_ (.B(_12777_),
    .A(_09702_),
    .X(_12778_));
 sg13g2_a21oi_2 _43491_ (.B1(_12776_),
    .Y(_12779_),
    .A2(_12778_),
    .A1(net5764));
 sg13g2_xnor2_1 _43492_ (.Y(_12780_),
    .A(net5463),
    .B(_12779_));
 sg13g2_o21ai_1 _43493_ (.B1(_12769_),
    .Y(_12781_),
    .A1(net5463),
    .A2(_12761_));
 sg13g2_a21oi_1 _43494_ (.A1(_12780_),
    .A2(_12781_),
    .Y(_12782_),
    .B1(net5564));
 sg13g2_o21ai_1 _43495_ (.B1(_12782_),
    .Y(_12783_),
    .A1(_12780_),
    .A2(_12781_));
 sg13g2_a21oi_1 _43496_ (.A1(net5564),
    .A2(_12779_),
    .Y(_12784_),
    .B1(net5931));
 sg13g2_nor2_1 _43497_ (.A(net5881),
    .B(_12761_),
    .Y(_12785_));
 sg13g2_a221oi_1 _43498_ (.B2(_12784_),
    .C1(_12785_),
    .B1(_12783_),
    .A1(net5993),
    .Y(_12786_),
    .A2(_09712_));
 sg13g2_o21ai_1 _43499_ (.B1(net6889),
    .Y(_12787_),
    .A1(net5289),
    .A2(_09712_));
 sg13g2_a21oi_1 _43500_ (.A1(net5289),
    .A2(_12786_),
    .Y(_12788_),
    .B1(_12787_));
 sg13g2_a21o_1 _43501_ (.A2(net6454),
    .A1(net2437),
    .B1(_12788_),
    .X(_00861_));
 sg13g2_nand2_1 _43502_ (.Y(_12789_),
    .A(net5723),
    .B(_09706_));
 sg13g2_a21oi_1 _43503_ (.A1(_09702_),
    .A2(_12777_),
    .Y(_12790_),
    .B1(_09701_));
 sg13g2_xor2_1 _43504_ (.B(_12790_),
    .A(_09707_),
    .X(_12791_));
 sg13g2_o21ai_1 _43505_ (.B1(_12789_),
    .Y(_12792_),
    .A1(net5737),
    .A2(_12791_));
 sg13g2_and2_1 _43506_ (.A(net5416),
    .B(_12792_),
    .X(_12793_));
 sg13g2_xnor2_1 _43507_ (.Y(_12794_),
    .A(net5464),
    .B(_12792_));
 sg13g2_a21o_1 _43508_ (.A2(_12779_),
    .A1(_12761_),
    .B1(net5463),
    .X(_12795_));
 sg13g2_a22oi_1 _43509_ (.Y(_12796_),
    .B1(_12795_),
    .B2(_12769_),
    .A2(_12779_),
    .A1(net5463));
 sg13g2_xnor2_1 _43510_ (.Y(_12797_),
    .A(_12794_),
    .B(_12796_));
 sg13g2_nor2_1 _43511_ (.A(net5531),
    .B(_12792_),
    .Y(_12798_));
 sg13g2_a21oi_1 _43512_ (.A1(net5531),
    .A2(_12797_),
    .Y(_12799_),
    .B1(_12798_));
 sg13g2_a22oi_1 _43513_ (.Y(_12800_),
    .B1(_12799_),
    .B2(net5232),
    .A2(_09717_),
    .A1(net5165));
 sg13g2_o21ai_1 _43514_ (.B1(_12800_),
    .Y(_12801_),
    .A1(net5120),
    .A2(_12779_));
 sg13g2_a22oi_1 _43515_ (.Y(_12802_),
    .B1(net6889),
    .B2(_12801_),
    .A2(net6456),
    .A1(net3360));
 sg13g2_inv_1 _43516_ (.Y(_00862_),
    .A(_12802_));
 sg13g2_nand2_1 _43517_ (.Y(_12803_),
    .A(net5722),
    .B(_10175_));
 sg13g2_a21o_2 _43518_ (.A2(_09944_),
    .A1(_09907_),
    .B1(_10177_),
    .X(_12804_));
 sg13g2_nand3_1 _43519_ (.B(_09944_),
    .C(_10177_),
    .A(_09907_),
    .Y(_12805_));
 sg13g2_nand3_1 _43520_ (.B(_12804_),
    .C(_12805_),
    .A(net5763),
    .Y(_12806_));
 sg13g2_nand2_2 _43521_ (.Y(_12807_),
    .A(_12803_),
    .B(_12806_));
 sg13g2_xnor2_1 _43522_ (.Y(_12808_),
    .A(net5464),
    .B(_12807_));
 sg13g2_a21oi_1 _43523_ (.A1(_12794_),
    .A2(_12796_),
    .Y(_12809_),
    .B1(_12793_));
 sg13g2_xor2_1 _43524_ (.B(_12809_),
    .A(_12808_),
    .X(_12810_));
 sg13g2_o21ai_1 _43525_ (.B1(net5961),
    .Y(_12811_),
    .A1(net5531),
    .A2(_12807_));
 sg13g2_a21oi_1 _43526_ (.A1(net5531),
    .A2(_12810_),
    .Y(_12812_),
    .B1(_12811_));
 sg13g2_nor2_1 _43527_ (.A(net6006),
    .B(_09700_),
    .Y(_12813_));
 sg13g2_a21oi_1 _43528_ (.A1(net5909),
    .A2(_12792_),
    .Y(_12814_),
    .B1(_12813_));
 sg13g2_nand2_1 _43529_ (.Y(_12815_),
    .A(net5289),
    .B(_12814_));
 sg13g2_nor2_1 _43530_ (.A(_12812_),
    .B(_12815_),
    .Y(_12816_));
 sg13g2_nor2b_1 _43531_ (.A(net5289),
    .B_N(_09700_),
    .Y(_12817_));
 sg13g2_nor3_1 _43532_ (.A(net6859),
    .B(_12816_),
    .C(_12817_),
    .Y(_12818_));
 sg13g2_a21o_1 _43533_ (.A2(net6454),
    .A1(net2401),
    .B1(_12818_),
    .X(_00863_));
 sg13g2_nand2_1 _43534_ (.Y(_12819_),
    .A(net3585),
    .B(net6443));
 sg13g2_nand2_1 _43535_ (.Y(_12820_),
    .A(net5722),
    .B(_10170_));
 sg13g2_nand2_1 _43536_ (.Y(_12821_),
    .A(_10176_),
    .B(_12804_));
 sg13g2_xor2_1 _43537_ (.B(_12821_),
    .A(_10172_),
    .X(_12822_));
 sg13g2_mux2_1 _43538_ (.A0(_10171_),
    .A1(_12822_),
    .S(net5760),
    .X(_12823_));
 sg13g2_o21ai_1 _43539_ (.B1(_12820_),
    .Y(_12824_),
    .A1(net5720),
    .A2(_12822_));
 sg13g2_nand2_1 _43540_ (.Y(_12825_),
    .A(net5563),
    .B(_12823_));
 sg13g2_nand2_1 _43541_ (.Y(_12826_),
    .A(net5415),
    .B(_12824_));
 sg13g2_xnor2_1 _43542_ (.Y(_12827_),
    .A(net5410),
    .B(_12823_));
 sg13g2_nand2_1 _43543_ (.Y(_12828_),
    .A(_12794_),
    .B(_12808_));
 sg13g2_nor3_1 _43544_ (.A(_12762_),
    .B(_12780_),
    .C(_12828_),
    .Y(_12829_));
 sg13g2_nor4_1 _43545_ (.A(_12762_),
    .B(_12767_),
    .C(_12780_),
    .D(_12828_),
    .Y(_12830_));
 sg13g2_and2_1 _43546_ (.A(_12707_),
    .B(_12830_),
    .X(_12831_));
 sg13g2_and2_1 _43547_ (.A(_12574_),
    .B(_12831_),
    .X(_12832_));
 sg13g2_nor2b_1 _43548_ (.A(_12706_),
    .B_N(_12830_),
    .Y(_12833_));
 sg13g2_and2_1 _43549_ (.A(_12765_),
    .B(_12829_),
    .X(_12834_));
 sg13g2_o21ai_1 _43550_ (.B1(net5416),
    .Y(_12835_),
    .A1(_12792_),
    .A2(_12807_));
 sg13g2_o21ai_1 _43551_ (.B1(_12835_),
    .Y(_12836_),
    .A1(_12795_),
    .A2(_12828_));
 sg13g2_nor4_2 _43552_ (.A(_12832_),
    .B(_12833_),
    .C(_12834_),
    .Y(_12837_),
    .D(_12836_));
 sg13g2_and2_1 _43553_ (.A(_12575_),
    .B(_12831_),
    .X(_12838_));
 sg13g2_o21ai_1 _43554_ (.B1(_12838_),
    .Y(_12839_),
    .A1(_12322_),
    .A2(_12315_));
 sg13g2_and2_1 _43555_ (.A(_12837_),
    .B(net1064),
    .X(_12840_));
 sg13g2_nand2b_1 _43556_ (.Y(_12841_),
    .B(_12827_),
    .A_N(_12840_));
 sg13g2_xnor2_1 _43557_ (.Y(_12842_),
    .A(_12827_),
    .B(_12840_));
 sg13g2_o21ai_1 _43558_ (.B1(_12825_),
    .Y(_12843_),
    .A1(net5563),
    .A2(_12842_));
 sg13g2_nor2_1 _43559_ (.A(net5153),
    .B(_12843_),
    .Y(_12844_));
 sg13g2_a221oi_1 _43560_ (.B2(net5212),
    .C1(_12844_),
    .B1(_12807_),
    .A1(net5162),
    .Y(_12845_),
    .A2(_09706_));
 sg13g2_o21ai_1 _43561_ (.B1(_12819_),
    .Y(_00864_),
    .A1(net6856),
    .A2(_12845_));
 sg13g2_nor2_1 _43562_ (.A(net5760),
    .B(_10158_),
    .Y(_12846_));
 sg13g2_a22oi_1 _43563_ (.Y(_12847_),
    .B1(_10185_),
    .B2(_12804_),
    .A2(_10171_),
    .A1(net5593));
 sg13g2_a221oi_1 _43564_ (.B2(_12804_),
    .C1(_10163_),
    .B1(_10185_),
    .A1(net5594),
    .Y(_12848_),
    .A2(_10171_));
 sg13g2_xnor2_1 _43565_ (.Y(_12849_),
    .A(_10163_),
    .B(_12847_));
 sg13g2_a21oi_2 _43566_ (.B1(_12846_),
    .Y(_12850_),
    .A2(_12849_),
    .A1(net5763));
 sg13g2_a21o_1 _43567_ (.A2(_12849_),
    .A1(net5764),
    .B1(_12846_),
    .X(_12851_));
 sg13g2_xnor2_1 _43568_ (.Y(_12852_),
    .A(net5410),
    .B(_12850_));
 sg13g2_nand3_1 _43569_ (.B(_12841_),
    .C(_12852_),
    .A(_12826_),
    .Y(_12853_));
 sg13g2_a21oi_1 _43570_ (.A1(_12826_),
    .A2(_12841_),
    .Y(_12854_),
    .B1(_12852_));
 sg13g2_nor2_1 _43571_ (.A(net5563),
    .B(_12854_),
    .Y(_12855_));
 sg13g2_a221oi_1 _43572_ (.B2(_12855_),
    .C1(net5927),
    .B1(_12853_),
    .A1(net5563),
    .Y(_12856_),
    .A2(_12850_));
 sg13g2_a221oi_1 _43573_ (.B2(net5905),
    .C1(_12856_),
    .B1(_12824_),
    .A1(net5991),
    .Y(_12857_),
    .A2(_10175_));
 sg13g2_a21oi_1 _43574_ (.A1(net5285),
    .A2(_12857_),
    .Y(_12858_),
    .B1(net6855));
 sg13g2_o21ai_1 _43575_ (.B1(_12858_),
    .Y(_12859_),
    .A1(net5285),
    .A2(_10175_));
 sg13g2_o21ai_1 _43576_ (.B1(_12859_),
    .Y(_00865_),
    .A1(_18136_),
    .A2(net6498));
 sg13g2_or3_1 _43577_ (.A(_10160_),
    .B(_10167_),
    .C(_12848_),
    .X(_12860_));
 sg13g2_o21ai_1 _43578_ (.B1(_10167_),
    .Y(_12861_),
    .A1(_10160_),
    .A2(_12848_));
 sg13g2_nor2_1 _43579_ (.A(net5760),
    .B(_10166_),
    .Y(_12862_));
 sg13g2_inv_1 _43580_ (.Y(_12863_),
    .A(_12862_));
 sg13g2_nand3_1 _43581_ (.B(_12860_),
    .C(_12861_),
    .A(net5762),
    .Y(_12864_));
 sg13g2_and2_1 _43582_ (.A(_12863_),
    .B(_12864_),
    .X(_12865_));
 sg13g2_nand3_1 _43583_ (.B(_12863_),
    .C(_12864_),
    .A(net5410),
    .Y(_12866_));
 sg13g2_inv_1 _43584_ (.Y(_12867_),
    .A(_12866_));
 sg13g2_a21o_1 _43585_ (.A2(_12864_),
    .A1(_12863_),
    .B1(net5410),
    .X(_12868_));
 sg13g2_and2_1 _43586_ (.A(_12866_),
    .B(_12868_),
    .X(_12869_));
 sg13g2_o21ai_1 _43587_ (.B1(net5415),
    .Y(_12870_),
    .A1(_12824_),
    .A2(_12851_));
 sg13g2_a21oi_1 _43588_ (.A1(_12823_),
    .A2(_12850_),
    .Y(_12871_),
    .B1(net5460));
 sg13g2_a22oi_1 _43589_ (.Y(_12872_),
    .B1(_12870_),
    .B2(_12841_),
    .A2(_12850_),
    .A1(net5463));
 sg13g2_xnor2_1 _43590_ (.Y(_12873_),
    .A(_12869_),
    .B(_12872_));
 sg13g2_o21ai_1 _43591_ (.B1(net5957),
    .Y(_12874_),
    .A1(net5530),
    .A2(_12865_));
 sg13g2_a21oi_1 _43592_ (.A1(net5530),
    .A2(_12873_),
    .Y(_12875_),
    .B1(_12874_));
 sg13g2_a221oi_1 _43593_ (.B2(net5905),
    .C1(_12875_),
    .B1(_12851_),
    .A1(net5990),
    .Y(_12876_),
    .A2(_10170_));
 sg13g2_o21ai_1 _43594_ (.B1(net6881),
    .Y(_12877_),
    .A1(net5285),
    .A2(_10170_));
 sg13g2_a21oi_1 _43595_ (.A1(net5285),
    .A2(_12876_),
    .Y(_12878_),
    .B1(_12877_));
 sg13g2_a21o_1 _43596_ (.A2(net6442),
    .A1(net3299),
    .B1(_12878_),
    .X(_00866_));
 sg13g2_o21ai_1 _43597_ (.B1(_10178_),
    .Y(_12879_),
    .A1(_09906_),
    .A2(_09945_));
 sg13g2_a21oi_1 _43598_ (.A1(_10188_),
    .A2(_12879_),
    .Y(_12880_),
    .B1(_10148_));
 sg13g2_and3_1 _43599_ (.X(_12881_),
    .A(_10148_),
    .B(_10188_),
    .C(_12879_));
 sg13g2_nor3_1 _43600_ (.A(net5720),
    .B(_12880_),
    .C(_12881_),
    .Y(_12882_));
 sg13g2_a21oi_1 _43601_ (.A1(net5720),
    .A2(_10147_),
    .Y(_12883_),
    .B1(_12882_));
 sg13g2_inv_1 _43602_ (.Y(_12884_),
    .A(_12883_));
 sg13g2_nand2_1 _43603_ (.Y(_12885_),
    .A(net5410),
    .B(_12884_));
 sg13g2_xnor2_1 _43604_ (.Y(_12886_),
    .A(net5411),
    .B(_12883_));
 sg13g2_a21oi_1 _43605_ (.A1(_12869_),
    .A2(_12872_),
    .Y(_12887_),
    .B1(_12867_));
 sg13g2_a21oi_1 _43606_ (.A1(_12886_),
    .A2(_12887_),
    .Y(_12888_),
    .B1(net5562));
 sg13g2_o21ai_1 _43607_ (.B1(_12888_),
    .Y(_12889_),
    .A1(_12886_),
    .A2(_12887_));
 sg13g2_a21oi_1 _43608_ (.A1(net5562),
    .A2(_12883_),
    .Y(_12890_),
    .B1(net5927));
 sg13g2_nand2_1 _43609_ (.Y(_12891_),
    .A(_12889_),
    .B(_12890_));
 sg13g2_a22oi_1 _43610_ (.Y(_12892_),
    .B1(_12865_),
    .B2(net5905),
    .A2(_10159_),
    .A1(net5990));
 sg13g2_nand3_1 _43611_ (.B(_12891_),
    .C(_12892_),
    .A(net5286),
    .Y(_12893_));
 sg13g2_nor2_1 _43612_ (.A(net5286),
    .B(_10159_),
    .Y(_12894_));
 sg13g2_nor2_1 _43613_ (.A(net6855),
    .B(_12894_),
    .Y(_12895_));
 sg13g2_a22oi_1 _43614_ (.Y(_12896_),
    .B1(_12893_),
    .B2(_12895_),
    .A2(net6442),
    .A1(net3751));
 sg13g2_inv_1 _43615_ (.Y(_00867_),
    .A(_12896_));
 sg13g2_or2_1 _43616_ (.X(_12897_),
    .B(_10140_),
    .A(net5760));
 sg13g2_a21oi_1 _43617_ (.A1(net5660),
    .A2(_10147_),
    .Y(_12898_),
    .B1(_12880_));
 sg13g2_xnor2_1 _43618_ (.Y(_12899_),
    .A(_10143_),
    .B(_12898_));
 sg13g2_o21ai_1 _43619_ (.B1(_12897_),
    .Y(_12900_),
    .A1(net5720),
    .A2(_12899_));
 sg13g2_nand2_1 _43620_ (.Y(_12901_),
    .A(net5411),
    .B(_12900_));
 sg13g2_xnor2_1 _43621_ (.Y(_12902_),
    .A(net5460),
    .B(_12900_));
 sg13g2_nand4_1 _43622_ (.B(_12868_),
    .C(_12871_),
    .A(_12866_),
    .Y(_12903_),
    .D(_12886_));
 sg13g2_nand3_1 _43623_ (.B(_12885_),
    .C(_12903_),
    .A(_12866_),
    .Y(_12904_));
 sg13g2_nand4_1 _43624_ (.B(_12852_),
    .C(_12869_),
    .A(_12827_),
    .Y(_12905_),
    .D(_12886_));
 sg13g2_nor2_1 _43625_ (.A(_12840_),
    .B(_12905_),
    .Y(_12906_));
 sg13g2_or2_1 _43626_ (.X(_12907_),
    .B(_12906_),
    .A(_12904_));
 sg13g2_nand2_1 _43627_ (.Y(_12908_),
    .A(_12902_),
    .B(_12907_));
 sg13g2_xnor2_1 _43628_ (.Y(_12909_),
    .A(_12902_),
    .B(_12907_));
 sg13g2_nor2_1 _43629_ (.A(net5526),
    .B(_12900_),
    .Y(_12910_));
 sg13g2_a21oi_1 _43630_ (.A1(net5526),
    .A2(_12909_),
    .Y(_12911_),
    .B1(_12910_));
 sg13g2_a22oi_1 _43631_ (.Y(_12912_),
    .B1(_12911_),
    .B2(net5229),
    .A2(_12884_),
    .A1(net5212));
 sg13g2_a22oi_1 _43632_ (.Y(_12913_),
    .B1(net5103),
    .B2(_10166_),
    .A2(net6440),
    .A1(net3363));
 sg13g2_o21ai_1 _43633_ (.B1(_12913_),
    .Y(_00868_),
    .A1(net6858),
    .A2(_12912_));
 sg13g2_nand2_1 _43634_ (.Y(_12914_),
    .A(_12901_),
    .B(_12908_));
 sg13g2_nor2_1 _43635_ (.A(net5762),
    .B(_10129_),
    .Y(_12915_));
 sg13g2_o21ai_1 _43636_ (.B1(_10142_),
    .Y(_12916_),
    .A1(_10191_),
    .A2(_12880_));
 sg13g2_xnor2_1 _43637_ (.Y(_12917_),
    .A(_10132_),
    .B(_12916_));
 sg13g2_a21oi_2 _43638_ (.B1(_12915_),
    .Y(_12918_),
    .A2(_12917_),
    .A1(net5760));
 sg13g2_nand2_1 _43639_ (.Y(_12919_),
    .A(net5411),
    .B(_12918_));
 sg13g2_nor2_1 _43640_ (.A(net5410),
    .B(_12918_),
    .Y(_12920_));
 sg13g2_xnor2_1 _43641_ (.Y(_12921_),
    .A(net5460),
    .B(_12918_));
 sg13g2_xnor2_1 _43642_ (.Y(_12922_),
    .A(_12914_),
    .B(_12921_));
 sg13g2_o21ai_1 _43643_ (.B1(net5956),
    .Y(_12923_),
    .A1(net5526),
    .A2(_12918_));
 sg13g2_a21oi_1 _43644_ (.A1(net5526),
    .A2(_12922_),
    .Y(_12924_),
    .B1(_12923_));
 sg13g2_a221oi_1 _43645_ (.B2(net5905),
    .C1(_12924_),
    .B1(_12900_),
    .A1(net5990),
    .Y(_12925_),
    .A2(_10147_));
 sg13g2_o21ai_1 _43646_ (.B1(net6881),
    .Y(_12926_),
    .A1(net5285),
    .A2(_10147_));
 sg13g2_a21oi_1 _43647_ (.A1(net5285),
    .A2(_12925_),
    .Y(_12927_),
    .B1(_12926_));
 sg13g2_a21o_1 _43648_ (.A2(net6439),
    .A1(net3413),
    .B1(_12927_),
    .X(_00869_));
 sg13g2_nand2_1 _43649_ (.Y(_12928_),
    .A(net3296),
    .B(net6440));
 sg13g2_nor2_1 _43650_ (.A(net5242),
    .B(_10140_),
    .Y(_12929_));
 sg13g2_nand2_1 _43651_ (.Y(_12930_),
    .A(net5720),
    .B(_10135_));
 sg13g2_o21ai_1 _43652_ (.B1(_10131_),
    .Y(_12931_),
    .A1(_10132_),
    .A2(_12916_));
 sg13g2_xor2_1 _43653_ (.B(_12931_),
    .A(_10137_),
    .X(_12932_));
 sg13g2_o21ai_1 _43654_ (.B1(_12930_),
    .Y(_12933_),
    .A1(net5720),
    .A2(_12932_));
 sg13g2_nor2_1 _43655_ (.A(net5526),
    .B(_12933_),
    .Y(_12934_));
 sg13g2_nand2_1 _43656_ (.Y(_12935_),
    .A(net5410),
    .B(_12933_));
 sg13g2_xnor2_1 _43657_ (.Y(_12936_),
    .A(net5460),
    .B(_12933_));
 sg13g2_nand2_1 _43658_ (.Y(_12937_),
    .A(_12901_),
    .B(_12919_));
 sg13g2_a21oi_1 _43659_ (.A1(_12902_),
    .A2(_12907_),
    .Y(_12938_),
    .B1(_12937_));
 sg13g2_nor2_1 _43660_ (.A(_12920_),
    .B(_12938_),
    .Y(_12939_));
 sg13g2_nand2_1 _43661_ (.Y(_12940_),
    .A(_12936_),
    .B(_12939_));
 sg13g2_xnor2_1 _43662_ (.Y(_12941_),
    .A(_12936_),
    .B(_12939_));
 sg13g2_a21oi_1 _43663_ (.A1(net5526),
    .A2(_12941_),
    .Y(_12942_),
    .B1(_12934_));
 sg13g2_a221oi_1 _43664_ (.B2(net5229),
    .C1(_12929_),
    .B1(_12942_),
    .A1(net5212),
    .Y(_12943_),
    .A2(_12918_));
 sg13g2_o21ai_1 _43665_ (.B1(_12928_),
    .Y(_00870_),
    .A1(net6854),
    .A2(_12943_));
 sg13g2_nand2_1 _43666_ (.Y(_12944_),
    .A(net3225),
    .B(net6439));
 sg13g2_nor2_1 _43667_ (.A(net5761),
    .B(_10118_),
    .Y(_12945_));
 sg13g2_a21oi_1 _43668_ (.A1(_09907_),
    .A2(_09944_),
    .Y(_12946_),
    .B1(_10180_));
 sg13g2_o21ai_1 _43669_ (.B1(_10179_),
    .Y(_12947_),
    .A1(_09906_),
    .A2(_09945_));
 sg13g2_o21ai_1 _43670_ (.B1(_10120_),
    .Y(_12948_),
    .A1(_10194_),
    .A2(_12946_));
 sg13g2_nor3_1 _43671_ (.A(_10120_),
    .B(_10194_),
    .C(_12946_),
    .Y(_12949_));
 sg13g2_nor2_1 _43672_ (.A(net5719),
    .B(_12949_),
    .Y(_12950_));
 sg13g2_a21oi_2 _43673_ (.B1(_12945_),
    .Y(_12951_),
    .A2(_12950_),
    .A1(_12948_));
 sg13g2_or2_1 _43674_ (.X(_12952_),
    .B(_12951_),
    .A(net5460));
 sg13g2_xnor2_1 _43675_ (.Y(_12953_),
    .A(net5410),
    .B(_12951_));
 sg13g2_nand2_1 _43676_ (.Y(_12954_),
    .A(_12935_),
    .B(_12940_));
 sg13g2_xor2_1 _43677_ (.B(_12954_),
    .A(_12953_),
    .X(_12955_));
 sg13g2_a21oi_1 _43678_ (.A1(net5561),
    .A2(_12951_),
    .Y(_12956_),
    .B1(net5927));
 sg13g2_o21ai_1 _43679_ (.B1(_12956_),
    .Y(_12957_),
    .A1(net5561),
    .A2(_12955_));
 sg13g2_a22oi_1 _43680_ (.Y(_12958_),
    .B1(_12933_),
    .B2(net5906),
    .A2(_10129_),
    .A1(net5991));
 sg13g2_and3_1 _43681_ (.X(_12959_),
    .A(net5281),
    .B(_12957_),
    .C(_12958_));
 sg13g2_o21ai_1 _43682_ (.B1(net6881),
    .Y(_12960_),
    .A1(net5281),
    .A2(_10129_));
 sg13g2_o21ai_1 _43683_ (.B1(_12944_),
    .Y(_00871_),
    .A1(_12959_),
    .A2(_12960_));
 sg13g2_nor2_1 _43684_ (.A(net5761),
    .B(_10112_),
    .Y(_12961_));
 sg13g2_nand2b_1 _43685_ (.Y(_12962_),
    .B(_12948_),
    .A_N(_10119_));
 sg13g2_xor2_1 _43686_ (.B(_12962_),
    .A(_10114_),
    .X(_12963_));
 sg13g2_a21oi_2 _43687_ (.B1(_12961_),
    .Y(_12964_),
    .A2(_12963_),
    .A1(net5761));
 sg13g2_nor2_1 _43688_ (.A(net5458),
    .B(_12964_),
    .Y(_12965_));
 sg13g2_xnor2_1 _43689_ (.Y(_12966_),
    .A(net5412),
    .B(_12964_));
 sg13g2_and2_1 _43690_ (.A(_12902_),
    .B(_12921_),
    .X(_12967_));
 sg13g2_nand3_1 _43691_ (.B(_12953_),
    .C(_12967_),
    .A(_12936_),
    .Y(_12968_));
 sg13g2_nand4_1 _43692_ (.B(_12936_),
    .C(_12953_),
    .A(_12904_),
    .Y(_12969_),
    .D(_12967_));
 sg13g2_nand3_1 _43693_ (.B(_12937_),
    .C(_12953_),
    .A(_12936_),
    .Y(_12970_));
 sg13g2_and4_1 _43694_ (.A(_12935_),
    .B(_12952_),
    .C(_12969_),
    .D(_12970_),
    .X(_12971_));
 sg13g2_nand4_1 _43695_ (.B(_12952_),
    .C(_12969_),
    .A(_12935_),
    .Y(_12972_),
    .D(_12970_));
 sg13g2_or2_1 _43696_ (.X(_12973_),
    .B(_12968_),
    .A(_12905_));
 sg13g2_o21ai_1 _43697_ (.B1(_12971_),
    .Y(_12974_),
    .A1(_12840_),
    .A2(_12973_));
 sg13g2_and2_1 _43698_ (.A(_12966_),
    .B(_12974_),
    .X(_12975_));
 sg13g2_xnor2_1 _43699_ (.Y(_12976_),
    .A(_12966_),
    .B(_12974_));
 sg13g2_nand2_1 _43700_ (.Y(_12977_),
    .A(net5561),
    .B(_12964_));
 sg13g2_a21oi_1 _43701_ (.A1(net5524),
    .A2(_12976_),
    .Y(_12978_),
    .B1(net5927));
 sg13g2_nor2_1 _43702_ (.A(net5882),
    .B(_12951_),
    .Y(_12979_));
 sg13g2_a221oi_1 _43703_ (.B2(_12978_),
    .C1(_12979_),
    .B1(_12977_),
    .A1(net5991),
    .Y(_12980_),
    .A2(_10135_));
 sg13g2_a21oi_1 _43704_ (.A1(net5281),
    .A2(_12980_),
    .Y(_12981_),
    .B1(net6854));
 sg13g2_o21ai_1 _43705_ (.B1(_12981_),
    .Y(_12982_),
    .A1(net5282),
    .A2(_10135_));
 sg13g2_o21ai_1 _43706_ (.B1(_12982_),
    .Y(_00872_),
    .A1(_18133_),
    .A2(net6498));
 sg13g2_nor2_1 _43707_ (.A(_12965_),
    .B(_12975_),
    .Y(_12983_));
 sg13g2_nand2_1 _43708_ (.Y(_12984_),
    .A(net5719),
    .B(_10102_));
 sg13g2_a22oi_1 _43709_ (.Y(_12985_),
    .B1(_10198_),
    .B2(_12948_),
    .A2(_10112_),
    .A1(net5592));
 sg13g2_a221oi_1 _43710_ (.B2(_12948_),
    .C1(_10103_),
    .B1(_10198_),
    .A1(net5593),
    .Y(_12986_),
    .A2(_10112_));
 sg13g2_xor2_1 _43711_ (.B(_12985_),
    .A(_10103_),
    .X(_12987_));
 sg13g2_o21ai_1 _43712_ (.B1(_12984_),
    .Y(_12988_),
    .A1(net5719),
    .A2(_12987_));
 sg13g2_or2_1 _43713_ (.X(_12989_),
    .B(_12988_),
    .A(net5412));
 sg13g2_xnor2_1 _43714_ (.Y(_12990_),
    .A(net5458),
    .B(_12988_));
 sg13g2_xor2_1 _43715_ (.B(_12990_),
    .A(_12983_),
    .X(_12991_));
 sg13g2_o21ai_1 _43716_ (.B1(net5956),
    .Y(_12992_),
    .A1(net5523),
    .A2(_12988_));
 sg13g2_a21oi_1 _43717_ (.A1(net5523),
    .A2(_12991_),
    .Y(_12993_),
    .B1(_12992_));
 sg13g2_nor2_1 _43718_ (.A(net6008),
    .B(_10118_),
    .Y(_12994_));
 sg13g2_nor2_1 _43719_ (.A(net5882),
    .B(_12964_),
    .Y(_12995_));
 sg13g2_nor3_1 _43720_ (.A(_12993_),
    .B(_12994_),
    .C(_12995_),
    .Y(_12996_));
 sg13g2_nand3_1 _43721_ (.B(net5317),
    .C(_10118_),
    .A(net5321),
    .Y(_12997_));
 sg13g2_a21oi_1 _43722_ (.A1(net5282),
    .A2(_12996_),
    .Y(_12998_),
    .B1(net6852));
 sg13g2_a22oi_1 _43723_ (.Y(_12999_),
    .B1(_12997_),
    .B2(_12998_),
    .A2(net6440),
    .A1(net2826));
 sg13g2_inv_1 _43724_ (.Y(_00873_),
    .A(_12999_));
 sg13g2_nand2_1 _43725_ (.Y(_13000_),
    .A(net5719),
    .B(_10107_));
 sg13g2_a21oi_1 _43726_ (.A1(net5659),
    .A2(_10102_),
    .Y(_13001_),
    .B1(_12986_));
 sg13g2_xor2_1 _43727_ (.B(_13001_),
    .A(_10108_),
    .X(_13002_));
 sg13g2_o21ai_1 _43728_ (.B1(_13000_),
    .Y(_13003_),
    .A1(net5719),
    .A2(_13002_));
 sg13g2_nand2_1 _43729_ (.Y(_13004_),
    .A(net5412),
    .B(_13003_));
 sg13g2_xnor2_1 _43730_ (.Y(_13005_),
    .A(net5461),
    .B(_13003_));
 sg13g2_inv_1 _43731_ (.Y(_13006_),
    .A(_13005_));
 sg13g2_a21o_1 _43732_ (.A2(_12988_),
    .A1(net5412),
    .B1(_12965_),
    .X(_13007_));
 sg13g2_o21ai_1 _43733_ (.B1(_12989_),
    .Y(_13008_),
    .A1(_12975_),
    .A2(_13007_));
 sg13g2_xnor2_1 _43734_ (.Y(_13009_),
    .A(_13006_),
    .B(_13008_));
 sg13g2_nor2_1 _43735_ (.A(net5523),
    .B(_13003_),
    .Y(_13010_));
 sg13g2_a21oi_1 _43736_ (.A1(net5524),
    .A2(_13009_),
    .Y(_13011_),
    .B1(_13010_));
 sg13g2_a22oi_1 _43737_ (.Y(_13012_),
    .B1(_13011_),
    .B2(net5228),
    .A2(_12988_),
    .A1(net5210));
 sg13g2_a22oi_1 _43738_ (.Y(_13013_),
    .B1(net5101),
    .B2(_10113_),
    .A2(net6440),
    .A1(net3307));
 sg13g2_o21ai_1 _43739_ (.B1(_13013_),
    .Y(_00874_),
    .A1(net6852),
    .A2(_13012_));
 sg13g2_nand2_1 _43740_ (.Y(_13014_),
    .A(net2082),
    .B(net6429));
 sg13g2_and2_1 _43741_ (.A(net5719),
    .B(_10092_),
    .X(_13015_));
 sg13g2_a21oi_1 _43742_ (.A1(_10193_),
    .A2(_12947_),
    .Y(_13016_),
    .B1(_10122_));
 sg13g2_nor2_1 _43743_ (.A(_10201_),
    .B(_13016_),
    .Y(_13017_));
 sg13g2_o21ai_1 _43744_ (.B1(_10095_),
    .Y(_13018_),
    .A1(_10201_),
    .A2(_13016_));
 sg13g2_a21oi_1 _43745_ (.A1(_10094_),
    .A2(_13017_),
    .Y(_13019_),
    .B1(net5720));
 sg13g2_a21o_2 _43746_ (.A2(_13019_),
    .A1(_13018_),
    .B1(_13015_),
    .X(_13020_));
 sg13g2_xnor2_1 _43747_ (.Y(_13021_),
    .A(net5461),
    .B(_13020_));
 sg13g2_o21ai_1 _43748_ (.B1(_13004_),
    .Y(_13022_),
    .A1(_13006_),
    .A2(_13008_));
 sg13g2_xnor2_1 _43749_ (.Y(_13023_),
    .A(_13021_),
    .B(_13022_));
 sg13g2_o21ai_1 _43750_ (.B1(net5953),
    .Y(_13024_),
    .A1(net5524),
    .A2(_13020_));
 sg13g2_a21oi_1 _43751_ (.A1(net5524),
    .A2(_13023_),
    .Y(_13025_),
    .B1(_13024_));
 sg13g2_a221oi_1 _43752_ (.B2(net5903),
    .C1(_13025_),
    .B1(_13003_),
    .A1(net5987),
    .Y(_13026_),
    .A2(_10102_));
 sg13g2_and2_1 _43753_ (.A(net5280),
    .B(_13026_),
    .X(_13027_));
 sg13g2_o21ai_1 _43754_ (.B1(net6880),
    .Y(_13028_),
    .A1(net5280),
    .A2(_10102_));
 sg13g2_o21ai_1 _43755_ (.B1(_13014_),
    .Y(_00875_),
    .A1(_13027_),
    .A2(_13028_));
 sg13g2_a21o_1 _43756_ (.A2(_13018_),
    .A1(_10093_),
    .B1(_10088_),
    .X(_13029_));
 sg13g2_nand3_1 _43757_ (.B(_10093_),
    .C(_13018_),
    .A(_10088_),
    .Y(_13030_));
 sg13g2_nand3_1 _43758_ (.B(_13029_),
    .C(_13030_),
    .A(net5761),
    .Y(_13031_));
 sg13g2_o21ai_1 _43759_ (.B1(_13031_),
    .Y(_13032_),
    .A1(net5761),
    .A2(_10086_));
 sg13g2_nor2_1 _43760_ (.A(net5523),
    .B(_13032_),
    .Y(_13033_));
 sg13g2_xnor2_1 _43761_ (.Y(_13034_),
    .A(net5458),
    .B(_13032_));
 sg13g2_nand3_1 _43762_ (.B(_13007_),
    .C(_13021_),
    .A(_13005_),
    .Y(_13035_));
 sg13g2_o21ai_1 _43763_ (.B1(net5412),
    .Y(_13036_),
    .A1(_13003_),
    .A2(_13020_));
 sg13g2_nand2_1 _43764_ (.Y(_13037_),
    .A(_13035_),
    .B(_13036_));
 sg13g2_nand4_1 _43765_ (.B(_12990_),
    .C(_13005_),
    .A(_12966_),
    .Y(_13038_),
    .D(_13021_));
 sg13g2_inv_1 _43766_ (.Y(_13039_),
    .A(_13038_));
 sg13g2_a21oi_1 _43767_ (.A1(_12974_),
    .A2(_13039_),
    .Y(_13040_),
    .B1(_13037_));
 sg13g2_nor2b_1 _43768_ (.A(_13040_),
    .B_N(_13034_),
    .Y(_13041_));
 sg13g2_xor2_1 _43769_ (.B(_13040_),
    .A(_13034_),
    .X(_13042_));
 sg13g2_a21oi_1 _43770_ (.A1(net5523),
    .A2(_13042_),
    .Y(_13043_),
    .B1(_13033_));
 sg13g2_a22oi_1 _43771_ (.Y(_13044_),
    .B1(_13043_),
    .B2(net5228),
    .A2(_13020_),
    .A1(net5210));
 sg13g2_a22oi_1 _43772_ (.Y(_13045_),
    .B1(net5102),
    .B2(_10107_),
    .A2(net6429),
    .A1(net3568));
 sg13g2_o21ai_1 _43773_ (.B1(_13045_),
    .Y(_00876_),
    .A1(net6852),
    .A2(_13044_));
 sg13g2_nor2_1 _43774_ (.A(net5761),
    .B(_10080_),
    .Y(_13046_));
 sg13g2_a22oi_1 _43775_ (.Y(_13047_),
    .B1(_10195_),
    .B2(_13018_),
    .A2(_10086_),
    .A1(net5592));
 sg13g2_a221oi_1 _43776_ (.B2(_13018_),
    .C1(_10083_),
    .B1(_10195_),
    .A1(net5592),
    .Y(_13048_),
    .A2(_10086_));
 sg13g2_xnor2_1 _43777_ (.Y(_13049_),
    .A(_10082_),
    .B(_13047_));
 sg13g2_a21oi_2 _43778_ (.B1(_13046_),
    .Y(_13050_),
    .A2(_13049_),
    .A1(net5761));
 sg13g2_nand2b_1 _43779_ (.Y(_13051_),
    .B(net5458),
    .A_N(_13050_));
 sg13g2_xnor2_1 _43780_ (.Y(_13052_),
    .A(net5458),
    .B(_13050_));
 sg13g2_a21oi_1 _43781_ (.A1(net5412),
    .A2(_13032_),
    .Y(_13053_),
    .B1(_13041_));
 sg13g2_xor2_1 _43782_ (.B(_13053_),
    .A(_13052_),
    .X(_13054_));
 sg13g2_o21ai_1 _43783_ (.B1(net5953),
    .Y(_13055_),
    .A1(net5523),
    .A2(_13050_));
 sg13g2_a21oi_1 _43784_ (.A1(net5523),
    .A2(_13054_),
    .Y(_13056_),
    .B1(_13055_));
 sg13g2_a221oi_1 _43785_ (.B2(net5904),
    .C1(_13056_),
    .B1(_13032_),
    .A1(net5987),
    .Y(_13057_),
    .A2(_10092_));
 sg13g2_o21ai_1 _43786_ (.B1(net6880),
    .Y(_13058_),
    .A1(net5282),
    .A2(_10092_));
 sg13g2_a21oi_1 _43787_ (.A1(net5282),
    .A2(_13057_),
    .Y(_13059_),
    .B1(_13058_));
 sg13g2_a21o_1 _43788_ (.A2(net6429),
    .A1(net2606),
    .B1(_13059_),
    .X(_00877_));
 sg13g2_or3_1 _43789_ (.A(_10068_),
    .B(_10081_),
    .C(_13048_),
    .X(_13060_));
 sg13g2_o21ai_1 _43790_ (.B1(_10068_),
    .Y(_13061_),
    .A1(_10081_),
    .A2(_13048_));
 sg13g2_and2_1 _43791_ (.A(net5719),
    .B(_10066_),
    .X(_13062_));
 sg13g2_a21oi_1 _43792_ (.A1(_13060_),
    .A2(_13061_),
    .Y(_13063_),
    .B1(net5719));
 sg13g2_or2_1 _43793_ (.X(_13064_),
    .B(_13063_),
    .A(_13062_));
 sg13g2_or3_1 _43794_ (.A(net5458),
    .B(_13062_),
    .C(_13063_),
    .X(_13065_));
 sg13g2_o21ai_1 _43795_ (.B1(net5458),
    .Y(_13066_),
    .A1(_13062_),
    .A2(_13063_));
 sg13g2_nand2_1 _43796_ (.Y(_13067_),
    .A(_13065_),
    .B(_13066_));
 sg13g2_o21ai_1 _43797_ (.B1(net5412),
    .Y(_13068_),
    .A1(_13032_),
    .A2(_13050_));
 sg13g2_inv_1 _43798_ (.Y(_13069_),
    .A(_13068_));
 sg13g2_o21ai_1 _43799_ (.B1(_13051_),
    .Y(_13070_),
    .A1(_13041_),
    .A2(_13069_));
 sg13g2_xnor2_1 _43800_ (.Y(_13071_),
    .A(_13067_),
    .B(_13070_));
 sg13g2_a21o_1 _43801_ (.A2(_13064_),
    .A1(net5561),
    .B1(net5926),
    .X(_13072_));
 sg13g2_a21oi_1 _43802_ (.A1(net5523),
    .A2(_13071_),
    .Y(_13073_),
    .B1(_13072_));
 sg13g2_a221oi_1 _43803_ (.B2(net5904),
    .C1(_13073_),
    .B1(_13050_),
    .A1(net5987),
    .Y(_13074_),
    .A2(_10087_));
 sg13g2_nand2_1 _43804_ (.Y(_13075_),
    .A(net5280),
    .B(_13074_));
 sg13g2_nor2_1 _43805_ (.A(net5283),
    .B(_10087_),
    .Y(_13076_));
 sg13g2_nor2_1 _43806_ (.A(net6852),
    .B(_13076_),
    .Y(_13077_));
 sg13g2_a22oi_1 _43807_ (.Y(_13078_),
    .B1(_13075_),
    .B2(_13077_),
    .A2(net6430),
    .A1(net3253));
 sg13g2_inv_1 _43808_ (.Y(_00878_),
    .A(_13078_));
 sg13g2_a21oi_2 _43809_ (.B1(_10182_),
    .Y(_13079_),
    .A2(_09944_),
    .A1(_09907_));
 sg13g2_o21ai_1 _43810_ (.B1(_10181_),
    .Y(_13080_),
    .A1(_09906_),
    .A2(_09945_));
 sg13g2_o21ai_1 _43811_ (.B1(_10058_),
    .Y(_13081_),
    .A1(_10204_),
    .A2(_13079_));
 sg13g2_nor3_1 _43812_ (.A(_10058_),
    .B(_10204_),
    .C(_13079_),
    .Y(_13082_));
 sg13g2_nor2_1 _43813_ (.A(net5711),
    .B(_13082_),
    .Y(_13083_));
 sg13g2_a22oi_1 _43814_ (.Y(_13084_),
    .B1(_13081_),
    .B2(_13083_),
    .A2(_10055_),
    .A1(net5711));
 sg13g2_inv_1 _43815_ (.Y(_13085_),
    .A(_13084_));
 sg13g2_xnor2_1 _43816_ (.Y(_13086_),
    .A(net5407),
    .B(_13084_));
 sg13g2_o21ai_1 _43817_ (.B1(_13065_),
    .Y(_13087_),
    .A1(_13067_),
    .A2(_13070_));
 sg13g2_xor2_1 _43818_ (.B(_13087_),
    .A(_13086_),
    .X(_13088_));
 sg13g2_a21oi_1 _43819_ (.A1(net5561),
    .A2(_13084_),
    .Y(_13089_),
    .B1(net5926));
 sg13g2_o21ai_1 _43820_ (.B1(_13089_),
    .Y(_13090_),
    .A1(net5561),
    .A2(_13088_));
 sg13g2_nor2_1 _43821_ (.A(net5882),
    .B(_13064_),
    .Y(_13091_));
 sg13g2_a21oi_1 _43822_ (.A1(net5987),
    .A2(_10080_),
    .Y(_13092_),
    .B1(_13091_));
 sg13g2_and3_1 _43823_ (.X(_13093_),
    .A(net5280),
    .B(_13090_),
    .C(_13092_));
 sg13g2_o21ai_1 _43824_ (.B1(net6880),
    .Y(_13094_),
    .A1(net5280),
    .A2(_10080_));
 sg13g2_nand2_1 _43825_ (.Y(_13095_),
    .A(net2744),
    .B(net6430));
 sg13g2_o21ai_1 _43826_ (.B1(_13095_),
    .Y(_00879_),
    .A1(_13093_),
    .A2(_13094_));
 sg13g2_and2_1 _43827_ (.A(_10056_),
    .B(_13081_),
    .X(_13096_));
 sg13g2_xnor2_1 _43828_ (.Y(_13097_),
    .A(_10051_),
    .B(_13096_));
 sg13g2_nor2_1 _43829_ (.A(net5755),
    .B(_10048_),
    .Y(_13098_));
 sg13g2_a21o_1 _43830_ (.A2(_13097_),
    .A1(net5756),
    .B1(_13098_),
    .X(_13099_));
 sg13g2_a21oi_1 _43831_ (.A1(net5756),
    .A2(_13097_),
    .Y(_13100_),
    .B1(_13098_));
 sg13g2_xnor2_1 _43832_ (.Y(_13101_),
    .A(net5407),
    .B(_13099_));
 sg13g2_nand3_1 _43833_ (.B(_13066_),
    .C(_13086_),
    .A(_13065_),
    .Y(_13102_));
 sg13g2_nand2_1 _43834_ (.Y(_13103_),
    .A(_13034_),
    .B(_13052_));
 sg13g2_nor2_1 _43835_ (.A(_13102_),
    .B(_13103_),
    .Y(_13104_));
 sg13g2_nor3_1 _43836_ (.A(_13038_),
    .B(_13102_),
    .C(_13103_),
    .Y(_13105_));
 sg13g2_nand2_1 _43837_ (.Y(_13106_),
    .A(_13039_),
    .B(_13104_));
 sg13g2_a21o_1 _43838_ (.A2(_13084_),
    .A1(_13064_),
    .B1(net5458),
    .X(_13107_));
 sg13g2_o21ai_1 _43839_ (.B1(_13107_),
    .Y(_13108_),
    .A1(_13068_),
    .A2(_13102_));
 sg13g2_a21oi_1 _43840_ (.A1(_13037_),
    .A2(_13104_),
    .Y(_13109_),
    .B1(_13108_));
 sg13g2_a221oi_1 _43841_ (.B2(_12972_),
    .C1(_13108_),
    .B1(_13105_),
    .A1(_13037_),
    .Y(_13110_),
    .A2(_13104_));
 sg13g2_o21ai_1 _43842_ (.B1(_13109_),
    .Y(_13111_),
    .A1(_12971_),
    .A2(_13106_));
 sg13g2_nor2_2 _43843_ (.A(_12973_),
    .B(_13106_),
    .Y(_13112_));
 sg13g2_inv_1 _43844_ (.Y(_13113_),
    .A(_13112_));
 sg13g2_a21oi_2 _43845_ (.B1(_13113_),
    .Y(_13114_),
    .A2(net1064),
    .A1(_12837_));
 sg13g2_nor2_1 _43846_ (.A(_13111_),
    .B(_13114_),
    .Y(_13115_));
 sg13g2_o21ai_1 _43847_ (.B1(_13101_),
    .Y(_13116_),
    .A1(_13111_),
    .A2(_13114_));
 sg13g2_xor2_1 _43848_ (.B(_13115_),
    .A(_13101_),
    .X(_13117_));
 sg13g2_nor2_1 _43849_ (.A(net5518),
    .B(_13100_),
    .Y(_13118_));
 sg13g2_a21oi_1 _43850_ (.A1(net5518),
    .A2(_13117_),
    .Y(_13119_),
    .B1(_13118_));
 sg13g2_a22oi_1 _43851_ (.Y(_13120_),
    .B1(_13119_),
    .B2(net5228),
    .A2(_13085_),
    .A1(net5210));
 sg13g2_nor2_1 _43852_ (.A(net5065),
    .B(_10066_),
    .Y(_13121_));
 sg13g2_a21oi_1 _43853_ (.A1(net3396),
    .A2(net6429),
    .Y(_13122_),
    .B1(_13121_));
 sg13g2_o21ai_1 _43854_ (.B1(_13122_),
    .Y(_00880_),
    .A1(net6852),
    .A2(_13120_));
 sg13g2_o21ai_1 _43855_ (.B1(_13116_),
    .Y(_13123_),
    .A1(net5455),
    .A2(_13099_));
 sg13g2_nor2_1 _43856_ (.A(net5755),
    .B(_10042_),
    .Y(_13124_));
 sg13g2_a21o_1 _43857_ (.A2(_13081_),
    .A1(_10206_),
    .B1(_10050_),
    .X(_13125_));
 sg13g2_a221oi_1 _43858_ (.B2(_13081_),
    .C1(_10044_),
    .B1(_10206_),
    .A1(net5587),
    .Y(_13126_),
    .A2(_10049_));
 sg13g2_xnor2_1 _43859_ (.Y(_13127_),
    .A(_10044_),
    .B(_13125_));
 sg13g2_a21oi_2 _43860_ (.B1(_13124_),
    .Y(_13128_),
    .A2(_13127_),
    .A1(net5755));
 sg13g2_nor2_1 _43861_ (.A(net5407),
    .B(_13128_),
    .Y(_13129_));
 sg13g2_xnor2_1 _43862_ (.Y(_13130_),
    .A(net5455),
    .B(_13128_));
 sg13g2_xnor2_1 _43863_ (.Y(_13131_),
    .A(_13123_),
    .B(_13130_));
 sg13g2_o21ai_1 _43864_ (.B1(net5953),
    .Y(_13132_),
    .A1(net5517),
    .A2(_13128_));
 sg13g2_a21oi_1 _43865_ (.A1(net5517),
    .A2(_13131_),
    .Y(_13133_),
    .B1(_13132_));
 sg13g2_a221oi_1 _43866_ (.B2(net5904),
    .C1(_13133_),
    .B1(_13100_),
    .A1(net5988),
    .Y(_13134_),
    .A2(_10055_));
 sg13g2_o21ai_1 _43867_ (.B1(net6880),
    .Y(_13135_),
    .A1(net5280),
    .A2(_10055_));
 sg13g2_a21oi_1 _43868_ (.A1(net5280),
    .A2(_13134_),
    .Y(_13136_),
    .B1(_13135_));
 sg13g2_a21o_1 _43869_ (.A2(net6430),
    .A1(net2726),
    .B1(_13136_),
    .X(_00881_));
 sg13g2_nand2_1 _43870_ (.Y(_13137_),
    .A(net5712),
    .B(_10036_));
 sg13g2_or3_1 _43871_ (.A(_10037_),
    .B(_10043_),
    .C(_13126_),
    .X(_13138_));
 sg13g2_o21ai_1 _43872_ (.B1(_10037_),
    .Y(_13139_),
    .A1(_10043_),
    .A2(_13126_));
 sg13g2_a21o_1 _43873_ (.A2(_13139_),
    .A1(_13138_),
    .B1(net5712),
    .X(_13140_));
 sg13g2_nand2_1 _43874_ (.Y(_13141_),
    .A(_13137_),
    .B(_13140_));
 sg13g2_a21oi_1 _43875_ (.A1(_13137_),
    .A2(_13140_),
    .Y(_13142_),
    .B1(net5455));
 sg13g2_xnor2_1 _43876_ (.Y(_13143_),
    .A(net5456),
    .B(_13141_));
 sg13g2_o21ai_1 _43877_ (.B1(net5407),
    .Y(_13144_),
    .A1(_13100_),
    .A2(_13128_));
 sg13g2_a21oi_1 _43878_ (.A1(_13116_),
    .A2(_13144_),
    .Y(_13145_),
    .B1(_13129_));
 sg13g2_xnor2_1 _43879_ (.Y(_13146_),
    .A(_13143_),
    .B(_13145_));
 sg13g2_nor2_1 _43880_ (.A(net5517),
    .B(_13141_),
    .Y(_13147_));
 sg13g2_a21oi_1 _43881_ (.A1(net5518),
    .A2(_13146_),
    .Y(_13148_),
    .B1(_13147_));
 sg13g2_a22oi_1 _43882_ (.Y(_13149_),
    .B1(_13148_),
    .B2(net5228),
    .A2(_13128_),
    .A1(net5210));
 sg13g2_a22oi_1 _43883_ (.Y(_13150_),
    .B1(net5102),
    .B2(_10048_),
    .A2(net6428),
    .A1(net2835));
 sg13g2_o21ai_1 _43884_ (.B1(_13150_),
    .Y(_00882_),
    .A1(net6853),
    .A2(_13149_));
 sg13g2_nand2_1 _43885_ (.Y(_13151_),
    .A(net2694),
    .B(net6428));
 sg13g2_a21oi_1 _43886_ (.A1(_10203_),
    .A2(_13080_),
    .Y(_13152_),
    .B1(_10060_));
 sg13g2_o21ai_1 _43887_ (.B1(_10031_),
    .Y(_13153_),
    .A1(_10209_),
    .A2(_13152_));
 sg13g2_or3_1 _43888_ (.A(_10031_),
    .B(_10209_),
    .C(_13152_),
    .X(_13154_));
 sg13g2_a21oi_1 _43889_ (.A1(_13153_),
    .A2(_13154_),
    .Y(_13155_),
    .B1(net5712));
 sg13g2_a21oi_2 _43890_ (.B1(_13155_),
    .Y(_13156_),
    .A2(_10028_),
    .A1(net5712));
 sg13g2_xnor2_1 _43891_ (.Y(_13157_),
    .A(net5456),
    .B(_13156_));
 sg13g2_a21oi_1 _43892_ (.A1(_13143_),
    .A2(_13145_),
    .Y(_13158_),
    .B1(_13142_));
 sg13g2_xor2_1 _43893_ (.B(_13158_),
    .A(_13157_),
    .X(_13159_));
 sg13g2_o21ai_1 _43894_ (.B1(net5953),
    .Y(_13160_),
    .A1(net5517),
    .A2(_13156_));
 sg13g2_a21oi_1 _43895_ (.A1(net5518),
    .A2(_13159_),
    .Y(_13161_),
    .B1(_13160_));
 sg13g2_a221oi_1 _43896_ (.B2(net5904),
    .C1(_13161_),
    .B1(_13141_),
    .A1(net5988),
    .Y(_13162_),
    .A2(_10042_));
 sg13g2_and2_1 _43897_ (.A(net5274),
    .B(_13162_),
    .X(_13163_));
 sg13g2_o21ai_1 _43898_ (.B1(net6883),
    .Y(_13164_),
    .A1(net5274),
    .A2(_10042_));
 sg13g2_o21ai_1 _43899_ (.B1(_13151_),
    .Y(_00883_),
    .A1(_13163_),
    .A2(_13164_));
 sg13g2_or2_1 _43900_ (.X(_13165_),
    .B(_10024_),
    .A(net5756));
 sg13g2_o21ai_1 _43901_ (.B1(_13153_),
    .Y(_13166_),
    .A1(net5588),
    .A2(_10028_));
 sg13g2_xor2_1 _43902_ (.B(_13166_),
    .A(_10025_),
    .X(_13167_));
 sg13g2_o21ai_1 _43903_ (.B1(_13165_),
    .Y(_13168_),
    .A1(net5712),
    .A2(_13167_));
 sg13g2_nor2_1 _43904_ (.A(net5517),
    .B(_13168_),
    .Y(_13169_));
 sg13g2_and2_1 _43905_ (.A(net5406),
    .B(_13168_),
    .X(_13170_));
 sg13g2_xnor2_1 _43906_ (.Y(_13171_),
    .A(net5455),
    .B(_13168_));
 sg13g2_nand2_1 _43907_ (.Y(_13172_),
    .A(_13143_),
    .B(_13157_));
 sg13g2_a21oi_1 _43908_ (.A1(net5407),
    .A2(_13156_),
    .Y(_13173_),
    .B1(_13142_));
 sg13g2_o21ai_1 _43909_ (.B1(_13173_),
    .Y(_13174_),
    .A1(_13144_),
    .A2(_13172_));
 sg13g2_and4_1 _43910_ (.A(_13101_),
    .B(_13130_),
    .C(_13143_),
    .D(_13157_),
    .X(_13175_));
 sg13g2_o21ai_1 _43911_ (.B1(_13175_),
    .Y(_13176_),
    .A1(_13111_),
    .A2(_13114_));
 sg13g2_nand2b_1 _43912_ (.Y(_13177_),
    .B(_13176_),
    .A_N(_13174_));
 sg13g2_and2_1 _43913_ (.A(_13171_),
    .B(_13177_),
    .X(_13178_));
 sg13g2_xnor2_1 _43914_ (.Y(_13179_),
    .A(_13171_),
    .B(_13177_));
 sg13g2_a21oi_1 _43915_ (.A1(net5517),
    .A2(_13179_),
    .Y(_13180_),
    .B1(_13169_));
 sg13g2_a22oi_1 _43916_ (.Y(_13181_),
    .B1(_13180_),
    .B2(net5228),
    .A2(_13156_),
    .A1(net5210));
 sg13g2_a22oi_1 _43917_ (.Y(_13182_),
    .B1(net5102),
    .B2(_10036_),
    .A2(net6430),
    .A1(net3625));
 sg13g2_o21ai_1 _43918_ (.B1(_13182_),
    .Y(_00884_),
    .A1(net6853),
    .A2(_13181_));
 sg13g2_nor2_1 _43919_ (.A(net5755),
    .B(_10016_),
    .Y(_13183_));
 sg13g2_a22oi_1 _43920_ (.Y(_13184_),
    .B1(_10210_),
    .B2(_13153_),
    .A2(_10024_),
    .A1(net5588));
 sg13g2_a221oi_1 _43921_ (.B2(_13153_),
    .C1(_10017_),
    .B1(_10210_),
    .A1(net5588),
    .Y(_13185_),
    .A2(_10024_));
 sg13g2_xor2_1 _43922_ (.B(_13184_),
    .A(_10017_),
    .X(_13186_));
 sg13g2_a21oi_2 _43923_ (.B1(_13183_),
    .Y(_13187_),
    .A2(_13186_),
    .A1(net5756));
 sg13g2_nor2_1 _43924_ (.A(net5406),
    .B(_13187_),
    .Y(_13188_));
 sg13g2_nand2_1 _43925_ (.Y(_13189_),
    .A(net5406),
    .B(_13187_));
 sg13g2_nand2b_1 _43926_ (.Y(_13190_),
    .B(_13189_),
    .A_N(_13188_));
 sg13g2_nor2_1 _43927_ (.A(_13170_),
    .B(_13178_),
    .Y(_13191_));
 sg13g2_xnor2_1 _43928_ (.Y(_13192_),
    .A(_13190_),
    .B(_13191_));
 sg13g2_o21ai_1 _43929_ (.B1(net5953),
    .Y(_13193_),
    .A1(net5517),
    .A2(_13187_));
 sg13g2_a21oi_1 _43930_ (.A1(net5517),
    .A2(_13192_),
    .Y(_13194_),
    .B1(_13193_));
 sg13g2_a221oi_1 _43931_ (.B2(net5904),
    .C1(_13194_),
    .B1(_13168_),
    .A1(net5988),
    .Y(_13195_),
    .A2(_10029_));
 sg13g2_nand3_1 _43932_ (.B(net5317),
    .C(_10028_),
    .A(net5321),
    .Y(_13196_));
 sg13g2_a21oi_1 _43933_ (.A1(net5280),
    .A2(_13195_),
    .Y(_13197_),
    .B1(net6853));
 sg13g2_a22oi_1 _43934_ (.Y(_13198_),
    .B1(_13196_),
    .B2(_13197_),
    .A2(net6428),
    .A1(net3366));
 sg13g2_inv_1 _43935_ (.Y(_00885_),
    .A(_13198_));
 sg13g2_nand2_1 _43936_ (.Y(_13199_),
    .A(net5711),
    .B(_10020_));
 sg13g2_a21oi_1 _43937_ (.A1(net5648),
    .A2(_10016_),
    .Y(_13200_),
    .B1(_13185_));
 sg13g2_xnor2_1 _43938_ (.Y(_13201_),
    .A(_10021_),
    .B(_13200_));
 sg13g2_o21ai_1 _43939_ (.B1(_13199_),
    .Y(_13202_),
    .A1(net5711),
    .A2(_13201_));
 sg13g2_nand2_1 _43940_ (.Y(_13203_),
    .A(net5406),
    .B(_13202_));
 sg13g2_xnor2_1 _43941_ (.Y(_13204_),
    .A(net5406),
    .B(_13202_));
 sg13g2_nand2b_1 _43942_ (.Y(_13205_),
    .B(_13189_),
    .A_N(_13170_));
 sg13g2_nor2_1 _43943_ (.A(_13178_),
    .B(_13205_),
    .Y(_13206_));
 sg13g2_or3_1 _43944_ (.A(_13188_),
    .B(_13204_),
    .C(_13206_),
    .X(_13207_));
 sg13g2_o21ai_1 _43945_ (.B1(_13204_),
    .Y(_13208_),
    .A1(_13188_),
    .A2(_13206_));
 sg13g2_and2_1 _43946_ (.A(_13207_),
    .B(_13208_),
    .X(_13209_));
 sg13g2_nor2_1 _43947_ (.A(net5516),
    .B(_13202_),
    .Y(_13210_));
 sg13g2_nor2_1 _43948_ (.A(net5929),
    .B(_13210_),
    .Y(_13211_));
 sg13g2_o21ai_1 _43949_ (.B1(_13211_),
    .Y(_13212_),
    .A1(net5559),
    .A2(_13209_));
 sg13g2_nor2_1 _43950_ (.A(net6008),
    .B(_10024_),
    .Y(_13213_));
 sg13g2_a21oi_1 _43951_ (.A1(net5904),
    .A2(_13187_),
    .Y(_13214_),
    .B1(_13213_));
 sg13g2_nand3_1 _43952_ (.B(_13212_),
    .C(_13214_),
    .A(net5274),
    .Y(_13215_));
 sg13g2_nand3_1 _43953_ (.B(net5317),
    .C(_10024_),
    .A(net5321),
    .Y(_13216_));
 sg13g2_nand3_1 _43954_ (.B(_13215_),
    .C(_13216_),
    .A(net6883),
    .Y(_13217_));
 sg13g2_o21ai_1 _43955_ (.B1(_13217_),
    .Y(_00886_),
    .A1(_18129_),
    .A2(net6499));
 sg13g2_a21oi_2 _43956_ (.B1(_10062_),
    .Y(_13218_),
    .A2(_13080_),
    .A1(_10203_));
 sg13g2_o21ai_1 _43957_ (.B1(_09998_),
    .Y(_13219_),
    .A1(_10214_),
    .A2(_13218_));
 sg13g2_nor3_1 _43958_ (.A(_09998_),
    .B(_10214_),
    .C(_13218_),
    .Y(_13220_));
 sg13g2_nand3b_1 _43959_ (.B(net5755),
    .C(_13219_),
    .Y(_13221_),
    .A_N(_13220_));
 sg13g2_o21ai_1 _43960_ (.B1(_13221_),
    .Y(_13222_),
    .A1(net5755),
    .A2(_09996_));
 sg13g2_nand2_1 _43961_ (.Y(_13223_),
    .A(net5406),
    .B(_13222_));
 sg13g2_xnor2_1 _43962_ (.Y(_13224_),
    .A(net5455),
    .B(_13222_));
 sg13g2_inv_1 _43963_ (.Y(_13225_),
    .A(_13224_));
 sg13g2_nand2_1 _43964_ (.Y(_13226_),
    .A(_13203_),
    .B(_13207_));
 sg13g2_xnor2_1 _43965_ (.Y(_13227_),
    .A(_13224_),
    .B(_13226_));
 sg13g2_o21ai_1 _43966_ (.B1(net5953),
    .Y(_13228_),
    .A1(net5516),
    .A2(_13222_));
 sg13g2_a21oi_1 _43967_ (.A1(net5516),
    .A2(_13227_),
    .Y(_13229_),
    .B1(_13228_));
 sg13g2_a22oi_1 _43968_ (.Y(_13230_),
    .B1(_13202_),
    .B2(net5904),
    .A2(_10016_),
    .A1(net5988));
 sg13g2_nand2_1 _43969_ (.Y(_13231_),
    .A(net5275),
    .B(_13230_));
 sg13g2_nor2_1 _43970_ (.A(net5274),
    .B(_10016_),
    .Y(_13232_));
 sg13g2_o21ai_1 _43971_ (.B1(net6877),
    .Y(_13233_),
    .A1(_13229_),
    .A2(_13231_));
 sg13g2_nand2_1 _43972_ (.Y(_13234_),
    .A(net2581),
    .B(net6428));
 sg13g2_o21ai_1 _43973_ (.B1(_13234_),
    .Y(_00887_),
    .A1(_13232_),
    .A2(_13233_));
 sg13g2_nand2_1 _43974_ (.Y(_13235_),
    .A(net3285),
    .B(net6428));
 sg13g2_o21ai_1 _43975_ (.B1(_13219_),
    .Y(_13236_),
    .A1(net5587),
    .A2(_09996_));
 sg13g2_xnor2_1 _43976_ (.Y(_13237_),
    .A(_10002_),
    .B(_13236_));
 sg13g2_nor2_1 _43977_ (.A(net5711),
    .B(_13237_),
    .Y(_13238_));
 sg13g2_a21oi_2 _43978_ (.B1(_13238_),
    .Y(_13239_),
    .A2(_10001_),
    .A1(net5711));
 sg13g2_and2_1 _43979_ (.A(net5405),
    .B(_13239_),
    .X(_13240_));
 sg13g2_xnor2_1 _43980_ (.Y(_13241_),
    .A(net5405),
    .B(_13239_));
 sg13g2_nor2_1 _43981_ (.A(_13204_),
    .B(_13225_),
    .Y(_13242_));
 sg13g2_nand3b_1 _43982_ (.B(_13189_),
    .C(_13171_),
    .Y(_13243_),
    .A_N(_13188_));
 sg13g2_nor3_1 _43983_ (.A(_13204_),
    .B(_13225_),
    .C(_13243_),
    .Y(_13244_));
 sg13g2_nand2_1 _43984_ (.Y(_13245_),
    .A(_13203_),
    .B(_13223_));
 sg13g2_a221oi_1 _43985_ (.B2(_13174_),
    .C1(_13245_),
    .B1(_13244_),
    .A1(_13205_),
    .Y(_13246_),
    .A2(_13242_));
 sg13g2_and2_1 _43986_ (.A(_13175_),
    .B(_13244_),
    .X(_13247_));
 sg13g2_o21ai_1 _43987_ (.B1(_13247_),
    .Y(_13248_),
    .A1(_13111_),
    .A2(_13114_));
 sg13g2_a21oi_1 _43988_ (.A1(_13246_),
    .A2(_13248_),
    .Y(_13249_),
    .B1(_13241_));
 sg13g2_nand3_1 _43989_ (.B(_13246_),
    .C(_13248_),
    .A(_13241_),
    .Y(_13250_));
 sg13g2_nand2b_1 _43990_ (.Y(_13251_),
    .B(_13250_),
    .A_N(_13249_));
 sg13g2_nand2_1 _43991_ (.Y(_13252_),
    .A(net5519),
    .B(_13251_));
 sg13g2_o21ai_1 _43992_ (.B1(_13252_),
    .Y(_13253_),
    .A1(net5516),
    .A2(_13239_));
 sg13g2_nor2_1 _43993_ (.A(net5153),
    .B(_13253_),
    .Y(_13254_));
 sg13g2_a221oi_1 _43994_ (.B2(net5210),
    .C1(_13254_),
    .B1(_13222_),
    .A1(net5163),
    .Y(_13255_),
    .A2(_10020_));
 sg13g2_o21ai_1 _43995_ (.B1(_13235_),
    .Y(_00888_),
    .A1(net6853),
    .A2(_13255_));
 sg13g2_nor2_1 _43996_ (.A(_13240_),
    .B(_13249_),
    .Y(_13256_));
 sg13g2_nand2_1 _43997_ (.Y(_13257_),
    .A(net5711),
    .B(_09983_));
 sg13g2_a22oi_1 _43998_ (.Y(_13258_),
    .B1(_10216_),
    .B2(_13219_),
    .A2(_10001_),
    .A1(net5587));
 sg13g2_a221oi_1 _43999_ (.B2(_13219_),
    .C1(_09986_),
    .B1(_10216_),
    .A1(net5587),
    .Y(_13259_),
    .A2(_10001_));
 sg13g2_o21ai_1 _44000_ (.B1(net5755),
    .Y(_13260_),
    .A1(_09985_),
    .A2(_13258_));
 sg13g2_o21ai_1 _44001_ (.B1(_13257_),
    .Y(_13261_),
    .A1(_13259_),
    .A2(_13260_));
 sg13g2_or2_1 _44002_ (.X(_13262_),
    .B(_13261_),
    .A(net5405));
 sg13g2_xnor2_1 _44003_ (.Y(_13263_),
    .A(net5405),
    .B(_13261_));
 sg13g2_xnor2_1 _44004_ (.Y(_13264_),
    .A(_13256_),
    .B(_13263_));
 sg13g2_o21ai_1 _44005_ (.B1(net5950),
    .Y(_13265_),
    .A1(net5516),
    .A2(_13261_));
 sg13g2_a21oi_1 _44006_ (.A1(net5516),
    .A2(_13264_),
    .Y(_13266_),
    .B1(_13265_));
 sg13g2_a221oi_1 _44007_ (.B2(net5900),
    .C1(_13266_),
    .B1(_13239_),
    .A1(net5984),
    .Y(_13267_),
    .A2(_09997_));
 sg13g2_o21ai_1 _44008_ (.B1(net6877),
    .Y(_13268_),
    .A1(net5274),
    .A2(_09997_));
 sg13g2_a21oi_1 _44009_ (.A1(net5274),
    .A2(_13267_),
    .Y(_13269_),
    .B1(_13268_));
 sg13g2_a21o_1 _44010_ (.A2(net6428),
    .A1(net2589),
    .B1(_13269_),
    .X(_00889_));
 sg13g2_nand2_1 _44011_ (.Y(_13270_),
    .A(net2490),
    .B(net6428));
 sg13g2_or3_1 _44012_ (.A(_09984_),
    .B(_09991_),
    .C(_13259_),
    .X(_13271_));
 sg13g2_o21ai_1 _44013_ (.B1(_09991_),
    .Y(_13272_),
    .A1(_09984_),
    .A2(_13259_));
 sg13g2_nand2_1 _44014_ (.Y(_13273_),
    .A(net5711),
    .B(_09990_));
 sg13g2_inv_1 _44015_ (.Y(_13274_),
    .A(_13273_));
 sg13g2_and3_1 _44016_ (.X(_13275_),
    .A(net5755),
    .B(_13271_),
    .C(_13272_));
 sg13g2_or2_1 _44017_ (.X(_13276_),
    .B(_13275_),
    .A(_13274_));
 sg13g2_o21ai_1 _44018_ (.B1(net5405),
    .Y(_13277_),
    .A1(_13274_),
    .A2(_13275_));
 sg13g2_nand3b_1 _44019_ (.B(net5455),
    .C(_13273_),
    .Y(_13278_),
    .A_N(_13275_));
 sg13g2_nand2_1 _44020_ (.Y(_13279_),
    .A(_13277_),
    .B(_13278_));
 sg13g2_o21ai_1 _44021_ (.B1(net5405),
    .Y(_13280_),
    .A1(_13239_),
    .A2(_13261_));
 sg13g2_a21o_1 _44022_ (.A2(_13261_),
    .A1(net5405),
    .B1(_13240_),
    .X(_13281_));
 sg13g2_o21ai_1 _44023_ (.B1(_13262_),
    .Y(_13282_),
    .A1(_13249_),
    .A2(_13281_));
 sg13g2_xnor2_1 _44024_ (.Y(_13283_),
    .A(_13279_),
    .B(_13282_));
 sg13g2_nor2_1 _44025_ (.A(net5516),
    .B(_13276_),
    .Y(_13284_));
 sg13g2_a21oi_1 _44026_ (.A1(net5516),
    .A2(_13283_),
    .Y(_13285_),
    .B1(_13284_));
 sg13g2_nor2_1 _44027_ (.A(net5242),
    .B(_10001_),
    .Y(_13286_));
 sg13g2_a221oi_1 _44028_ (.B2(net5226),
    .C1(_13286_),
    .B1(_13285_),
    .A1(net5206),
    .Y(_13287_),
    .A2(_13261_));
 sg13g2_o21ai_1 _44029_ (.B1(_13270_),
    .Y(_00890_),
    .A1(net6848),
    .A2(_13287_));
 sg13g2_o21ai_1 _44030_ (.B1(_10005_),
    .Y(_13288_),
    .A1(_10214_),
    .A2(_13218_));
 sg13g2_a21oi_1 _44031_ (.A1(_10219_),
    .A2(_13288_),
    .Y(_13289_),
    .B1(_09976_));
 sg13g2_nand3_1 _44032_ (.B(_10219_),
    .C(_13288_),
    .A(_09976_),
    .Y(_13290_));
 sg13g2_nand2b_1 _44033_ (.Y(_13291_),
    .B(_13290_),
    .A_N(_13289_));
 sg13g2_mux2_1 _44034_ (.A0(_09973_),
    .A1(_13291_),
    .S(net5753),
    .X(_13292_));
 sg13g2_inv_1 _44035_ (.Y(_13293_),
    .A(_13292_));
 sg13g2_xnor2_1 _44036_ (.Y(_13294_),
    .A(net5405),
    .B(_13292_));
 sg13g2_o21ai_1 _44037_ (.B1(_13277_),
    .Y(_13295_),
    .A1(_13279_),
    .A2(_13282_));
 sg13g2_xor2_1 _44038_ (.B(_13295_),
    .A(_13294_),
    .X(_13296_));
 sg13g2_a21oi_1 _44039_ (.A1(net5559),
    .A2(_13292_),
    .Y(_13297_),
    .B1(net5924));
 sg13g2_o21ai_1 _44040_ (.B1(_13297_),
    .Y(_13298_),
    .A1(net5559),
    .A2(_13296_));
 sg13g2_a22oi_1 _44041_ (.Y(_13299_),
    .B1(_13276_),
    .B2(net5900),
    .A2(_09983_),
    .A1(net5984));
 sg13g2_and3_1 _44042_ (.X(_13300_),
    .A(net5274),
    .B(_13298_),
    .C(_13299_));
 sg13g2_o21ai_1 _44043_ (.B1(net6877),
    .Y(_13301_),
    .A1(net5274),
    .A2(_09983_));
 sg13g2_nand2_1 _44044_ (.Y(_13302_),
    .A(net2886),
    .B(net6428));
 sg13g2_o21ai_1 _44045_ (.B1(_13302_),
    .Y(_00891_),
    .A1(_13300_),
    .A2(_13301_));
 sg13g2_nor2_1 _44046_ (.A(_09974_),
    .B(_13289_),
    .Y(_13303_));
 sg13g2_xnor2_1 _44047_ (.Y(_13304_),
    .A(_09969_),
    .B(_13303_));
 sg13g2_nand2b_1 _44048_ (.Y(_13305_),
    .B(net5708),
    .A_N(_09968_));
 sg13g2_o21ai_1 _44049_ (.B1(_13305_),
    .Y(_13306_),
    .A1(net5708),
    .A2(_13304_));
 sg13g2_or2_1 _44050_ (.X(_13307_),
    .B(_13306_),
    .A(net5450));
 sg13g2_xnor2_1 _44051_ (.Y(_13308_),
    .A(net5399),
    .B(_13306_));
 sg13g2_nand3_1 _44052_ (.B(_13278_),
    .C(_13294_),
    .A(_13277_),
    .Y(_13309_));
 sg13g2_o21ai_1 _44053_ (.B1(_13277_),
    .Y(_13310_),
    .A1(_13280_),
    .A2(_13309_));
 sg13g2_a21o_1 _44054_ (.A2(_13293_),
    .A1(net5399),
    .B1(_13310_),
    .X(_13311_));
 sg13g2_or3_1 _44055_ (.A(_13241_),
    .B(_13263_),
    .C(_13309_),
    .X(_13312_));
 sg13g2_a21oi_1 _44056_ (.A1(_13246_),
    .A2(_13248_),
    .Y(_13313_),
    .B1(_13312_));
 sg13g2_o21ai_1 _44057_ (.B1(_13308_),
    .Y(_13314_),
    .A1(_13311_),
    .A2(_13313_));
 sg13g2_or3_1 _44058_ (.A(_13308_),
    .B(_13311_),
    .C(_13313_),
    .X(_13315_));
 sg13g2_a21oi_1 _44059_ (.A1(_13314_),
    .A2(_13315_),
    .Y(_13316_),
    .B1(net5558));
 sg13g2_a21oi_1 _44060_ (.A1(net5559),
    .A2(_13306_),
    .Y(_13317_),
    .B1(_13316_));
 sg13g2_a22oi_1 _44061_ (.Y(_13318_),
    .B1(_13317_),
    .B2(net5227),
    .A2(_13293_),
    .A1(net5206));
 sg13g2_a22oi_1 _44062_ (.Y(_13319_),
    .B1(net5099),
    .B2(_09990_),
    .A2(net6416),
    .A1(net2950));
 sg13g2_o21ai_1 _44063_ (.B1(_13319_),
    .Y(_00892_),
    .A1(net6848),
    .A2(_13318_));
 sg13g2_a21oi_1 _44064_ (.A1(_09969_),
    .A2(_13289_),
    .Y(_13320_),
    .B1(_10220_));
 sg13g2_xor2_1 _44065_ (.B(_13320_),
    .A(_09959_),
    .X(_13321_));
 sg13g2_mux2_1 _44066_ (.A0(_09957_),
    .A1(_13321_),
    .S(net5753),
    .X(_13322_));
 sg13g2_inv_1 _44067_ (.Y(_13323_),
    .A(_13322_));
 sg13g2_nand2_1 _44068_ (.Y(_13324_),
    .A(net5399),
    .B(_13322_));
 sg13g2_xnor2_1 _44069_ (.Y(_13325_),
    .A(net5450),
    .B(_13322_));
 sg13g2_nand3_1 _44070_ (.B(_13314_),
    .C(_13325_),
    .A(_13307_),
    .Y(_13326_));
 sg13g2_a21oi_1 _44071_ (.A1(_13307_),
    .A2(_13314_),
    .Y(_13327_),
    .B1(_13325_));
 sg13g2_nor2_1 _44072_ (.A(net5558),
    .B(_13327_),
    .Y(_13328_));
 sg13g2_a221oi_1 _44073_ (.B2(_13328_),
    .C1(net5924),
    .B1(_13326_),
    .A1(net5558),
    .Y(_13329_),
    .A2(_13323_));
 sg13g2_nor2_1 _44074_ (.A(net6004),
    .B(_09973_),
    .Y(_13330_));
 sg13g2_nor2_1 _44075_ (.A(net5883),
    .B(_13306_),
    .Y(_13331_));
 sg13g2_nor3_1 _44076_ (.A(_13329_),
    .B(_13330_),
    .C(_13331_),
    .Y(_13332_));
 sg13g2_nand2_1 _44077_ (.Y(_13333_),
    .A(net5273),
    .B(_13332_));
 sg13g2_nor2b_1 _44078_ (.A(net5273),
    .B_N(_09973_),
    .Y(_13334_));
 sg13g2_nor2_1 _44079_ (.A(net6848),
    .B(_13334_),
    .Y(_13335_));
 sg13g2_a22oi_1 _44080_ (.Y(_13336_),
    .B1(_13333_),
    .B2(_13335_),
    .A2(net6417),
    .A1(net2669));
 sg13g2_inv_1 _44081_ (.Y(_00893_),
    .A(_13336_));
 sg13g2_nand2_1 _44082_ (.Y(_13337_),
    .A(net3220),
    .B(net6417));
 sg13g2_nand2_1 _44083_ (.Y(_13338_),
    .A(net5708),
    .B(_09962_));
 sg13g2_o21ai_1 _44084_ (.B1(_09958_),
    .Y(_13339_),
    .A1(_09959_),
    .A2(_13320_));
 sg13g2_xnor2_1 _44085_ (.Y(_13340_),
    .A(_09964_),
    .B(_13339_));
 sg13g2_o21ai_1 _44086_ (.B1(_13338_),
    .Y(_13341_),
    .A1(net5708),
    .A2(_13340_));
 sg13g2_nand2_1 _44087_ (.Y(_13342_),
    .A(net5558),
    .B(_13341_));
 sg13g2_nor2_1 _44088_ (.A(net5450),
    .B(_13341_),
    .Y(_13343_));
 sg13g2_xnor2_1 _44089_ (.Y(_13344_),
    .A(net5450),
    .B(_13341_));
 sg13g2_and2_1 _44090_ (.A(_13307_),
    .B(_13324_),
    .X(_13345_));
 sg13g2_nand2_1 _44091_ (.Y(_13346_),
    .A(_13307_),
    .B(_13324_));
 sg13g2_nand2_1 _44092_ (.Y(_13347_),
    .A(_13314_),
    .B(_13345_));
 sg13g2_o21ai_1 _44093_ (.B1(_13347_),
    .Y(_13348_),
    .A1(net5399),
    .A2(_13322_));
 sg13g2_a221oi_1 _44094_ (.B2(_13314_),
    .C1(_13344_),
    .B1(_13345_),
    .A1(net5450),
    .Y(_13349_),
    .A2(_13323_));
 sg13g2_xor2_1 _44095_ (.B(_13348_),
    .A(_13344_),
    .X(_13350_));
 sg13g2_o21ai_1 _44096_ (.B1(_13342_),
    .Y(_13351_),
    .A1(net5558),
    .A2(_13350_));
 sg13g2_nor2_1 _44097_ (.A(net5152),
    .B(_13351_),
    .Y(_13352_));
 sg13g2_a221oi_1 _44098_ (.B2(net5206),
    .C1(_13352_),
    .B1(_13322_),
    .A1(net5159),
    .Y(_13353_),
    .A2(_09968_));
 sg13g2_o21ai_1 _44099_ (.B1(_13337_),
    .Y(_00894_),
    .A1(net6848),
    .A2(_13353_));
 sg13g2_nand2_1 _44100_ (.Y(_13354_),
    .A(net5706),
    .B(_08811_));
 sg13g2_a21o_2 _44101_ (.A2(_10223_),
    .A1(net1094),
    .B1(_08850_),
    .X(_13355_));
 sg13g2_nand3_1 _44102_ (.B(net1094),
    .C(_10223_),
    .A(_08850_),
    .Y(_13356_));
 sg13g2_nand3_1 _44103_ (.B(_13355_),
    .C(_13356_),
    .A(net5753),
    .Y(_13357_));
 sg13g2_nand2_2 _44104_ (.Y(_13358_),
    .A(_13354_),
    .B(_13357_));
 sg13g2_nand2_1 _44105_ (.Y(_13359_),
    .A(net5399),
    .B(_13358_));
 sg13g2_xnor2_1 _44106_ (.Y(_13360_),
    .A(net5450),
    .B(_13358_));
 sg13g2_inv_2 _44107_ (.Y(_13361_),
    .A(_13360_));
 sg13g2_nor2_1 _44108_ (.A(_13343_),
    .B(_13349_),
    .Y(_13362_));
 sg13g2_xnor2_1 _44109_ (.Y(_13363_),
    .A(_13361_),
    .B(_13362_));
 sg13g2_o21ai_1 _44110_ (.B1(net5950),
    .Y(_13364_),
    .A1(net5509),
    .A2(_13358_));
 sg13g2_a21o_1 _44111_ (.A2(_13363_),
    .A1(net5509),
    .B1(_13364_),
    .X(_13365_));
 sg13g2_nor2_1 _44112_ (.A(net5883),
    .B(_13341_),
    .Y(_13366_));
 sg13g2_a221oi_1 _44113_ (.B2(_09957_),
    .C1(_13366_),
    .B1(net5984),
    .A1(net5320),
    .Y(_13367_),
    .A2(net5316));
 sg13g2_o21ai_1 _44114_ (.B1(net6877),
    .Y(_13368_),
    .A1(net5273),
    .A2(_09957_));
 sg13g2_a21oi_1 _44115_ (.A1(_13365_),
    .A2(_13367_),
    .Y(_13369_),
    .B1(_13368_));
 sg13g2_a21oi_1 _44116_ (.A1(net2471),
    .A2(net6417),
    .Y(_13370_),
    .B1(_13369_));
 sg13g2_inv_1 _44117_ (.Y(_00895_),
    .A(_13370_));
 sg13g2_nand2_1 _44118_ (.Y(_13371_),
    .A(net5706),
    .B(_08806_));
 sg13g2_nor2b_1 _44119_ (.A(_08812_),
    .B_N(_13355_),
    .Y(_13372_));
 sg13g2_xnor2_1 _44120_ (.Y(_13373_),
    .A(_08851_),
    .B(_13372_));
 sg13g2_o21ai_1 _44121_ (.B1(_13371_),
    .Y(_13374_),
    .A1(net5706),
    .A2(_13373_));
 sg13g2_nand2_1 _44122_ (.Y(_13375_),
    .A(net5397),
    .B(_13374_));
 sg13g2_xnor2_1 _44123_ (.Y(_13376_),
    .A(net5449),
    .B(_13374_));
 sg13g2_nor2_1 _44124_ (.A(_13344_),
    .B(_13361_),
    .Y(_13377_));
 sg13g2_nand2_1 _44125_ (.Y(_13378_),
    .A(_13308_),
    .B(_13325_));
 sg13g2_nor3_1 _44126_ (.A(_13344_),
    .B(_13361_),
    .C(_13378_),
    .Y(_13379_));
 sg13g2_nor4_1 _44127_ (.A(_13312_),
    .B(_13344_),
    .C(_13361_),
    .D(_13378_),
    .Y(_13380_));
 sg13g2_nand3b_1 _44128_ (.B(_13247_),
    .C(_13380_),
    .Y(_13381_),
    .A_N(_13110_));
 sg13g2_nand2b_1 _44129_ (.Y(_13382_),
    .B(_13380_),
    .A_N(_13246_));
 sg13g2_a221oi_1 _44130_ (.B2(_13311_),
    .C1(_13343_),
    .B1(_13379_),
    .A1(_13346_),
    .Y(_13383_),
    .A2(_13377_));
 sg13g2_nand4_1 _44131_ (.B(_13381_),
    .C(_13382_),
    .A(_13359_),
    .Y(_13384_),
    .D(_13383_));
 sg13g2_nand3_1 _44132_ (.B(_13247_),
    .C(_13380_),
    .A(_13112_),
    .Y(_13385_));
 sg13g2_a21oi_1 _44133_ (.A1(_12837_),
    .A2(net1064),
    .Y(_13386_),
    .B1(_13385_));
 sg13g2_or2_1 _44134_ (.X(_13387_),
    .B(_13386_),
    .A(_13384_));
 sg13g2_nand2_1 _44135_ (.Y(_13388_),
    .A(_13376_),
    .B(_13387_));
 sg13g2_xnor2_1 _44136_ (.Y(_13389_),
    .A(_13376_),
    .B(_13387_));
 sg13g2_nor2_1 _44137_ (.A(net5507),
    .B(_13374_),
    .Y(_13390_));
 sg13g2_a21oi_1 _44138_ (.A1(net5507),
    .A2(_13389_),
    .Y(_13391_),
    .B1(_13390_));
 sg13g2_a22oi_1 _44139_ (.Y(_13392_),
    .B1(_13391_),
    .B2(net5227),
    .A2(_13358_),
    .A1(net5207));
 sg13g2_a22oi_1 _44140_ (.Y(_13393_),
    .B1(net5098),
    .B2(_09963_),
    .A2(net6416),
    .A1(net3314));
 sg13g2_o21ai_1 _44141_ (.B1(_13393_),
    .Y(_00896_),
    .A1(net6847),
    .A2(_13392_));
 sg13g2_nand2_1 _44142_ (.Y(_13394_),
    .A(_13375_),
    .B(_13388_));
 sg13g2_nand2_1 _44143_ (.Y(_13395_),
    .A(net5706),
    .B(_08801_));
 sg13g2_a22oi_1 _44144_ (.Y(_13396_),
    .B1(_08813_),
    .B2(_13355_),
    .A2(_08807_),
    .A1(net5582));
 sg13g2_a221oi_1 _44145_ (.B2(_13355_),
    .C1(_08803_),
    .B1(_08813_),
    .A1(net5582),
    .Y(_13397_),
    .A2(_08807_));
 sg13g2_xor2_1 _44146_ (.B(_13396_),
    .A(_08803_),
    .X(_13398_));
 sg13g2_o21ai_1 _44147_ (.B1(_13395_),
    .Y(_13399_),
    .A1(net5706),
    .A2(_13398_));
 sg13g2_xnor2_1 _44148_ (.Y(_13400_),
    .A(net5398),
    .B(_13399_));
 sg13g2_xor2_1 _44149_ (.B(_13400_),
    .A(_13394_),
    .X(_13401_));
 sg13g2_o21ai_1 _44150_ (.B1(net5950),
    .Y(_13402_),
    .A1(net5508),
    .A2(_13399_));
 sg13g2_a21oi_1 _44151_ (.A1(net5508),
    .A2(_13401_),
    .Y(_13403_),
    .B1(_13402_));
 sg13g2_a221oi_1 _44152_ (.B2(net5899),
    .C1(_13403_),
    .B1(_13374_),
    .A1(net5984),
    .Y(_13404_),
    .A2(_08811_));
 sg13g2_o21ai_1 _44153_ (.B1(net6876),
    .Y(_13405_),
    .A1(net5271),
    .A2(_08811_));
 sg13g2_a21oi_1 _44154_ (.A1(net5271),
    .A2(_13404_),
    .Y(_13406_),
    .B1(_13405_));
 sg13g2_a21o_1 _44155_ (.A2(net6416),
    .A1(net3105),
    .B1(_13406_),
    .X(_00897_));
 sg13g2_nand2_1 _44156_ (.Y(_13407_),
    .A(net5706),
    .B(_08794_));
 sg13g2_or3_1 _44157_ (.A(_08796_),
    .B(_08802_),
    .C(_13397_),
    .X(_13408_));
 sg13g2_o21ai_1 _44158_ (.B1(_08796_),
    .Y(_13409_),
    .A1(_08802_),
    .A2(_13397_));
 sg13g2_a21o_1 _44159_ (.A2(_13409_),
    .A1(_13408_),
    .B1(net5707),
    .X(_13410_));
 sg13g2_nand2_1 _44160_ (.Y(_13411_),
    .A(_13407_),
    .B(_13410_));
 sg13g2_nor2_1 _44161_ (.A(net5507),
    .B(_13411_),
    .Y(_13412_));
 sg13g2_a21oi_1 _44162_ (.A1(_13407_),
    .A2(_13410_),
    .Y(_13413_),
    .B1(net5449));
 sg13g2_nand2_1 _44163_ (.Y(_13414_),
    .A(net5397),
    .B(_13411_));
 sg13g2_nand3_1 _44164_ (.B(_13407_),
    .C(_13410_),
    .A(net5449),
    .Y(_13415_));
 sg13g2_nor2b_1 _44165_ (.A(_13413_),
    .B_N(_13415_),
    .Y(_13416_));
 sg13g2_inv_1 _44166_ (.Y(_13417_),
    .A(_13416_));
 sg13g2_o21ai_1 _44167_ (.B1(net5398),
    .Y(_13418_),
    .A1(_13374_),
    .A2(_13399_));
 sg13g2_nand2_1 _44168_ (.Y(_13419_),
    .A(_13388_),
    .B(_13418_));
 sg13g2_o21ai_1 _44169_ (.B1(_13419_),
    .Y(_13420_),
    .A1(net5398),
    .A2(_13399_));
 sg13g2_xnor2_1 _44170_ (.Y(_13421_),
    .A(_13417_),
    .B(_13420_));
 sg13g2_a21oi_1 _44171_ (.A1(net5509),
    .A2(_13421_),
    .Y(_13422_),
    .B1(_13412_));
 sg13g2_a22oi_1 _44172_ (.Y(_13423_),
    .B1(_13422_),
    .B2(net5226),
    .A2(_13399_),
    .A1(net5206));
 sg13g2_a22oi_1 _44173_ (.Y(_13424_),
    .B1(net5099),
    .B2(_08806_),
    .A2(net6416),
    .A1(net2266));
 sg13g2_o21ai_1 _44174_ (.B1(_13424_),
    .Y(_00898_),
    .A1(net6847),
    .A2(_13423_));
 sg13g2_nand2_1 _44175_ (.Y(_13425_),
    .A(net2006),
    .B(net6416));
 sg13g2_nand2_1 _44176_ (.Y(_13426_),
    .A(net5707),
    .B(_08788_));
 sg13g2_a21oi_1 _44177_ (.A1(net1094),
    .A2(_10223_),
    .Y(_13427_),
    .B1(_08853_));
 sg13g2_o21ai_1 _44178_ (.B1(_08790_),
    .Y(_13428_),
    .A1(_08816_),
    .A2(_13427_));
 sg13g2_or3_1 _44179_ (.A(_08790_),
    .B(_08816_),
    .C(_13427_),
    .X(_13429_));
 sg13g2_nand2_1 _44180_ (.Y(_13430_),
    .A(_13428_),
    .B(_13429_));
 sg13g2_o21ai_1 _44181_ (.B1(_13426_),
    .Y(_13431_),
    .A1(net5707),
    .A2(_13430_));
 sg13g2_xnor2_1 _44182_ (.Y(_13432_),
    .A(net5449),
    .B(_13431_));
 sg13g2_o21ai_1 _44183_ (.B1(_13414_),
    .Y(_13433_),
    .A1(_13417_),
    .A2(_13420_));
 sg13g2_xnor2_1 _44184_ (.Y(_13434_),
    .A(_13432_),
    .B(_13433_));
 sg13g2_o21ai_1 _44185_ (.B1(net5950),
    .Y(_13435_),
    .A1(net5506),
    .A2(_13431_));
 sg13g2_a21oi_1 _44186_ (.A1(net5506),
    .A2(_13434_),
    .Y(_13436_),
    .B1(_13435_));
 sg13g2_a221oi_1 _44187_ (.B2(net5900),
    .C1(_13436_),
    .B1(_13411_),
    .A1(net5984),
    .Y(_13437_),
    .A2(_08801_));
 sg13g2_and2_1 _44188_ (.A(net5271),
    .B(_13437_),
    .X(_13438_));
 sg13g2_o21ai_1 _44189_ (.B1(net6876),
    .Y(_13439_),
    .A1(net5272),
    .A2(_08801_));
 sg13g2_o21ai_1 _44190_ (.B1(_13425_),
    .Y(_00899_),
    .A1(_13438_),
    .A2(_13439_));
 sg13g2_nand2_1 _44191_ (.Y(_13440_),
    .A(net5707),
    .B(_08783_));
 sg13g2_nand2_1 _44192_ (.Y(_13441_),
    .A(_08789_),
    .B(_13428_));
 sg13g2_xnor2_1 _44193_ (.Y(_13442_),
    .A(_08785_),
    .B(_13441_));
 sg13g2_o21ai_1 _44194_ (.B1(_13440_),
    .Y(_13443_),
    .A1(net5707),
    .A2(_13442_));
 sg13g2_nand2_1 _44195_ (.Y(_13444_),
    .A(net5397),
    .B(_13443_));
 sg13g2_xnor2_1 _44196_ (.Y(_13445_),
    .A(net5449),
    .B(_13443_));
 sg13g2_nand3b_1 _44197_ (.B(_13415_),
    .C(_13432_),
    .Y(_13446_),
    .A_N(_13413_));
 sg13g2_a21oi_1 _44198_ (.A1(net5397),
    .A2(_13431_),
    .Y(_13447_),
    .B1(_13413_));
 sg13g2_o21ai_1 _44199_ (.B1(_13447_),
    .Y(_13448_),
    .A1(_13418_),
    .A2(_13446_));
 sg13g2_nand3_1 _44200_ (.B(_13416_),
    .C(_13432_),
    .A(_13376_),
    .Y(_13449_));
 sg13g2_nor2_1 _44201_ (.A(_13400_),
    .B(_13449_),
    .Y(_13450_));
 sg13g2_a21oi_1 _44202_ (.A1(_13387_),
    .A2(_13450_),
    .Y(_13451_),
    .B1(_13448_));
 sg13g2_nand2b_1 _44203_ (.Y(_13452_),
    .B(_13445_),
    .A_N(_13451_));
 sg13g2_xor2_1 _44204_ (.B(_13451_),
    .A(_13445_),
    .X(_13453_));
 sg13g2_o21ai_1 _44205_ (.B1(net5950),
    .Y(_13454_),
    .A1(net5506),
    .A2(_13443_));
 sg13g2_a21oi_1 _44206_ (.A1(net5507),
    .A2(_13453_),
    .Y(_13455_),
    .B1(_13454_));
 sg13g2_a221oi_1 _44207_ (.B2(net5899),
    .C1(_13455_),
    .B1(_13431_),
    .A1(net5984),
    .Y(_13456_),
    .A2(_08794_));
 sg13g2_a21oi_1 _44208_ (.A1(net5272),
    .A2(_13456_),
    .Y(_13457_),
    .B1(net6847));
 sg13g2_o21ai_1 _44209_ (.B1(_13457_),
    .Y(_13458_),
    .A1(net5271),
    .A2(_08794_));
 sg13g2_o21ai_1 _44210_ (.B1(_13458_),
    .Y(_00900_),
    .A1(_18125_),
    .A2(net6489));
 sg13g2_nor2_1 _44211_ (.A(net5752),
    .B(_08777_),
    .Y(_13459_));
 sg13g2_a22oi_1 _44212_ (.Y(_13460_),
    .B1(_08818_),
    .B2(_13428_),
    .A2(_08784_),
    .A1(net5582));
 sg13g2_xnor2_1 _44213_ (.Y(_13461_),
    .A(_08779_),
    .B(_13460_));
 sg13g2_a21oi_2 _44214_ (.B1(_13459_),
    .Y(_13462_),
    .A2(_13461_),
    .A1(net5752));
 sg13g2_nor2_1 _44215_ (.A(net5397),
    .B(_13462_),
    .Y(_13463_));
 sg13g2_xnor2_1 _44216_ (.Y(_13464_),
    .A(net5449),
    .B(_13462_));
 sg13g2_and2_1 _44217_ (.A(_13444_),
    .B(_13452_),
    .X(_13465_));
 sg13g2_xor2_1 _44218_ (.B(_13465_),
    .A(_13464_),
    .X(_13466_));
 sg13g2_o21ai_1 _44219_ (.B1(net5949),
    .Y(_13467_),
    .A1(net5506),
    .A2(_13462_));
 sg13g2_a21oi_1 _44220_ (.A1(net5507),
    .A2(_13466_),
    .Y(_13468_),
    .B1(_13467_));
 sg13g2_a221oi_1 _44221_ (.B2(net5900),
    .C1(_13468_),
    .B1(_13443_),
    .A1(net5984),
    .Y(_13469_),
    .A2(_08788_));
 sg13g2_o21ai_1 _44222_ (.B1(net6876),
    .Y(_13470_),
    .A1(net5271),
    .A2(_08788_));
 sg13g2_a21oi_1 _44223_ (.A1(net5271),
    .A2(_13469_),
    .Y(_13471_),
    .B1(_13470_));
 sg13g2_a21o_1 _44224_ (.A2(net6416),
    .A1(net2712),
    .B1(_13471_),
    .X(_00901_));
 sg13g2_nand2_1 _44225_ (.Y(_13472_),
    .A(net5706),
    .B(_08766_));
 sg13g2_a21oi_1 _44226_ (.A1(_08779_),
    .A2(_13460_),
    .Y(_13473_),
    .B1(_08778_));
 sg13g2_xnor2_1 _44227_ (.Y(_13474_),
    .A(_08768_),
    .B(_13473_));
 sg13g2_o21ai_1 _44228_ (.B1(_13472_),
    .Y(_13475_),
    .A1(net5706),
    .A2(_13474_));
 sg13g2_xnor2_1 _44229_ (.Y(_13476_),
    .A(net5449),
    .B(_13475_));
 sg13g2_o21ai_1 _44230_ (.B1(net5397),
    .Y(_13477_),
    .A1(_13443_),
    .A2(_13462_));
 sg13g2_a21oi_1 _44231_ (.A1(_13452_),
    .A2(_13477_),
    .Y(_13478_),
    .B1(_13463_));
 sg13g2_and2_1 _44232_ (.A(_13476_),
    .B(_13478_),
    .X(_13479_));
 sg13g2_xnor2_1 _44233_ (.Y(_13480_),
    .A(_13476_),
    .B(_13478_));
 sg13g2_o21ai_1 _44234_ (.B1(net5949),
    .Y(_13481_),
    .A1(net5506),
    .A2(_13475_));
 sg13g2_a21oi_1 _44235_ (.A1(net5506),
    .A2(_13480_),
    .Y(_13482_),
    .B1(_13481_));
 sg13g2_a221oi_1 _44236_ (.B2(net5900),
    .C1(_13482_),
    .B1(_13462_),
    .A1(net5983),
    .Y(_13483_),
    .A2(_08783_));
 sg13g2_a21oi_1 _44237_ (.A1(net5271),
    .A2(_13483_),
    .Y(_13484_),
    .B1(net6847));
 sg13g2_o21ai_1 _44238_ (.B1(_13484_),
    .Y(_13485_),
    .A1(net5271),
    .A2(_08783_));
 sg13g2_o21ai_1 _44239_ (.B1(_13485_),
    .Y(_00902_),
    .A1(_18124_),
    .A2(net6489));
 sg13g2_a21oi_1 _44240_ (.A1(net1094),
    .A2(_10223_),
    .Y(_13486_),
    .B1(_08855_));
 sg13g2_o21ai_1 _44241_ (.B1(_08760_),
    .Y(_13487_),
    .A1(_08821_),
    .A2(_13486_));
 sg13g2_or3_1 _44242_ (.A(_08760_),
    .B(_08821_),
    .C(_13486_),
    .X(_13488_));
 sg13g2_nand3_1 _44243_ (.B(_13487_),
    .C(_13488_),
    .A(net5752),
    .Y(_13489_));
 sg13g2_o21ai_1 _44244_ (.B1(_13489_),
    .Y(_13490_),
    .A1(net5752),
    .A2(_08759_));
 sg13g2_xnor2_1 _44245_ (.Y(_13491_),
    .A(net5449),
    .B(_13490_));
 sg13g2_a21o_1 _44246_ (.A2(_13475_),
    .A1(net5397),
    .B1(_13479_),
    .X(_13492_));
 sg13g2_xnor2_1 _44247_ (.Y(_13493_),
    .A(_13491_),
    .B(_13492_));
 sg13g2_o21ai_1 _44248_ (.B1(net5950),
    .Y(_13494_),
    .A1(net5506),
    .A2(_13490_));
 sg13g2_a21oi_1 _44249_ (.A1(net5506),
    .A2(_13493_),
    .Y(_13495_),
    .B1(_13494_));
 sg13g2_a22oi_1 _44250_ (.Y(_13496_),
    .B1(_13475_),
    .B2(net5899),
    .A2(_08777_),
    .A1(net5983));
 sg13g2_nand2_1 _44251_ (.Y(_13497_),
    .A(net5272),
    .B(_13496_));
 sg13g2_nor2_1 _44252_ (.A(_13495_),
    .B(_13497_),
    .Y(_13498_));
 sg13g2_o21ai_1 _44253_ (.B1(net6876),
    .Y(_13499_),
    .A1(net5263),
    .A2(_08777_));
 sg13g2_nand2_1 _44254_ (.Y(_13500_),
    .A(net2991),
    .B(net6416));
 sg13g2_o21ai_1 _44255_ (.B1(_13500_),
    .Y(_00903_),
    .A1(_13498_),
    .A2(_13499_));
 sg13g2_nand2_1 _44256_ (.Y(_13501_),
    .A(net3181),
    .B(net6416));
 sg13g2_nor2_1 _44257_ (.A(net5752),
    .B(_08753_),
    .Y(_13502_));
 sg13g2_o21ai_1 _44258_ (.B1(_13487_),
    .Y(_13503_),
    .A1(net5581),
    .A2(_08759_));
 sg13g2_xor2_1 _44259_ (.B(_13503_),
    .A(_08755_),
    .X(_13504_));
 sg13g2_a21oi_2 _44260_ (.B1(_13502_),
    .Y(_13505_),
    .A2(_13504_),
    .A1(net5752));
 sg13g2_xnor2_1 _44261_ (.Y(_13506_),
    .A(net5448),
    .B(_13505_));
 sg13g2_and2_1 _44262_ (.A(_13445_),
    .B(_13464_),
    .X(_13507_));
 sg13g2_nand4_1 _44263_ (.B(_13476_),
    .C(_13491_),
    .A(_13448_),
    .Y(_13508_),
    .D(_13507_));
 sg13g2_nand3b_1 _44264_ (.B(_13491_),
    .C(_13476_),
    .Y(_13509_),
    .A_N(_13477_));
 sg13g2_o21ai_1 _44265_ (.B1(net5397),
    .Y(_13510_),
    .A1(_13475_),
    .A2(_13490_));
 sg13g2_nand3_1 _44266_ (.B(_13509_),
    .C(_13510_),
    .A(_13508_),
    .Y(_13511_));
 sg13g2_and4_1 _44267_ (.A(_13450_),
    .B(_13476_),
    .C(_13491_),
    .D(_13507_),
    .X(_13512_));
 sg13g2_a21oi_1 _44268_ (.A1(_13387_),
    .A2(_13512_),
    .Y(_13513_),
    .B1(_13511_));
 sg13g2_nor2b_1 _44269_ (.A(_13513_),
    .B_N(_13506_),
    .Y(_13514_));
 sg13g2_nor2b_1 _44270_ (.A(_13506_),
    .B_N(_13513_),
    .Y(_13515_));
 sg13g2_o21ai_1 _44271_ (.B1(net5503),
    .Y(_13516_),
    .A1(_13514_),
    .A2(_13515_));
 sg13g2_o21ai_1 _44272_ (.B1(_13516_),
    .Y(_13517_),
    .A1(net5503),
    .A2(_13505_));
 sg13g2_nor2_1 _44273_ (.A(net5152),
    .B(_13517_),
    .Y(_13518_));
 sg13g2_a221oi_1 _44274_ (.B2(net5206),
    .C1(_13518_),
    .B1(_13490_),
    .A1(net5159),
    .Y(_13519_),
    .A2(_08766_));
 sg13g2_o21ai_1 _44275_ (.B1(_13501_),
    .Y(_00904_),
    .A1(net6847),
    .A2(_13519_));
 sg13g2_a21oi_1 _44276_ (.A1(net5394),
    .A2(_13505_),
    .Y(_13520_),
    .B1(_13514_));
 sg13g2_nand2_1 _44277_ (.Y(_13521_),
    .A(net5703),
    .B(_08749_));
 sg13g2_a22oi_1 _44278_ (.Y(_13522_),
    .B1(_08822_),
    .B2(_13487_),
    .A2(_08754_),
    .A1(net5581));
 sg13g2_a221oi_1 _44279_ (.B2(_13487_),
    .C1(_08750_),
    .B1(_08822_),
    .A1(net5581),
    .Y(_13523_),
    .A2(_08754_));
 sg13g2_xor2_1 _44280_ (.B(_13522_),
    .A(_08750_),
    .X(_13524_));
 sg13g2_o21ai_1 _44281_ (.B1(_13521_),
    .Y(_13525_),
    .A1(net5703),
    .A2(_13524_));
 sg13g2_or2_1 _44282_ (.X(_13526_),
    .B(_13525_),
    .A(net5394));
 sg13g2_xnor2_1 _44283_ (.Y(_13527_),
    .A(net5448),
    .B(_13525_));
 sg13g2_xor2_1 _44284_ (.B(_13527_),
    .A(_13520_),
    .X(_13528_));
 sg13g2_o21ai_1 _44285_ (.B1(net5949),
    .Y(_13529_),
    .A1(net5504),
    .A2(_13525_));
 sg13g2_a21oi_1 _44286_ (.A1(net5504),
    .A2(_13528_),
    .Y(_13530_),
    .B1(_13529_));
 sg13g2_nand2_1 _44287_ (.Y(_13531_),
    .A(net5899),
    .B(_13505_));
 sg13g2_o21ai_1 _44288_ (.B1(_13531_),
    .Y(_13532_),
    .A1(net6004),
    .A2(_08759_));
 sg13g2_nor2_1 _44289_ (.A(_13530_),
    .B(_13532_),
    .Y(_13533_));
 sg13g2_nand3_1 _44290_ (.B(net5316),
    .C(_08759_),
    .A(net5320),
    .Y(_13534_));
 sg13g2_a21oi_1 _44291_ (.A1(net5264),
    .A2(_13533_),
    .Y(_13535_),
    .B1(net6847));
 sg13g2_a22oi_1 _44292_ (.Y(_13536_),
    .B1(_13534_),
    .B2(_13535_),
    .A2(net6414),
    .A1(net3058));
 sg13g2_inv_1 _44293_ (.Y(_00905_),
    .A(_13536_));
 sg13g2_nand2_1 _44294_ (.Y(_13537_),
    .A(net5703),
    .B(_08743_));
 sg13g2_a21oi_1 _44295_ (.A1(net5637),
    .A2(_08749_),
    .Y(_13538_),
    .B1(_13523_));
 sg13g2_xnor2_1 _44296_ (.Y(_13539_),
    .A(_08744_),
    .B(_13538_));
 sg13g2_o21ai_1 _44297_ (.B1(_13537_),
    .Y(_13540_),
    .A1(net5703),
    .A2(_13539_));
 sg13g2_nand2_1 _44298_ (.Y(_13541_),
    .A(net5395),
    .B(_13540_));
 sg13g2_nor2_1 _44299_ (.A(net5395),
    .B(_13540_),
    .Y(_13542_));
 sg13g2_xnor2_1 _44300_ (.Y(_13543_),
    .A(net5448),
    .B(_13540_));
 sg13g2_o21ai_1 _44301_ (.B1(net5395),
    .Y(_13544_),
    .A1(_13505_),
    .A2(_13525_));
 sg13g2_inv_1 _44302_ (.Y(_13545_),
    .A(_13544_));
 sg13g2_o21ai_1 _44303_ (.B1(_13526_),
    .Y(_13546_),
    .A1(_13514_),
    .A2(_13545_));
 sg13g2_xor2_1 _44304_ (.B(_13546_),
    .A(_13543_),
    .X(_13547_));
 sg13g2_nand2_1 _44305_ (.Y(_13548_),
    .A(net5503),
    .B(_13547_));
 sg13g2_o21ai_1 _44306_ (.B1(_13548_),
    .Y(_13549_),
    .A1(net5504),
    .A2(_13540_));
 sg13g2_a22oi_1 _44307_ (.Y(_13550_),
    .B1(_13525_),
    .B2(net5206),
    .A2(_08753_),
    .A1(net5159));
 sg13g2_o21ai_1 _44308_ (.B1(_13550_),
    .Y(_13551_),
    .A1(net5152),
    .A2(_13549_));
 sg13g2_a22oi_1 _44309_ (.Y(_13552_),
    .B1(net6876),
    .B2(_13551_),
    .A2(net6415),
    .A1(net3561));
 sg13g2_inv_1 _44310_ (.Y(_00906_),
    .A(_13552_));
 sg13g2_o21ai_1 _44311_ (.B1(_08762_),
    .Y(_13553_),
    .A1(_08821_),
    .A2(_13486_));
 sg13g2_a21oi_1 _44312_ (.A1(_08825_),
    .A2(_13553_),
    .Y(_13554_),
    .B1(_08732_));
 sg13g2_and3_1 _44313_ (.X(_13555_),
    .A(_08732_),
    .B(_08825_),
    .C(_13553_));
 sg13g2_nor3_1 _44314_ (.A(net5704),
    .B(_13554_),
    .C(_13555_),
    .Y(_13556_));
 sg13g2_a21oi_2 _44315_ (.B1(_13556_),
    .Y(_13557_),
    .A2(_08730_),
    .A1(net5704));
 sg13g2_nor2_1 _44316_ (.A(net5448),
    .B(_13557_),
    .Y(_13558_));
 sg13g2_xnor2_1 _44317_ (.Y(_13559_),
    .A(net5395),
    .B(_13557_));
 sg13g2_o21ai_1 _44318_ (.B1(_13541_),
    .Y(_13560_),
    .A1(_13542_),
    .A2(_13546_));
 sg13g2_xnor2_1 _44319_ (.Y(_13561_),
    .A(_13559_),
    .B(_13560_));
 sg13g2_nand2_1 _44320_ (.Y(_13562_),
    .A(net5503),
    .B(_13561_));
 sg13g2_a21oi_1 _44321_ (.A1(net5558),
    .A2(_13557_),
    .Y(_13563_),
    .B1(net5924));
 sg13g2_a22oi_1 _44322_ (.Y(_13564_),
    .B1(_13540_),
    .B2(net5899),
    .A2(_08749_),
    .A1(net5983));
 sg13g2_nand2_1 _44323_ (.Y(_13565_),
    .A(net5263),
    .B(_13564_));
 sg13g2_a21oi_1 _44324_ (.A1(_13562_),
    .A2(_13563_),
    .Y(_13566_),
    .B1(_13565_));
 sg13g2_o21ai_1 _44325_ (.B1(net6876),
    .Y(_13567_),
    .A1(net5263),
    .A2(_08749_));
 sg13g2_nand2_1 _44326_ (.Y(_13568_),
    .A(net2427),
    .B(net6415));
 sg13g2_o21ai_1 _44327_ (.B1(_13568_),
    .Y(_00907_),
    .A1(_13566_),
    .A2(_13567_));
 sg13g2_nand2_1 _44328_ (.Y(_13569_),
    .A(net5703),
    .B(_08736_));
 sg13g2_a21oi_1 _44329_ (.A1(net5636),
    .A2(_08730_),
    .Y(_13570_),
    .B1(_13554_));
 sg13g2_xor2_1 _44330_ (.B(_13570_),
    .A(_08737_),
    .X(_13571_));
 sg13g2_o21ai_1 _44331_ (.B1(_13569_),
    .Y(_13572_),
    .A1(net5704),
    .A2(_13571_));
 sg13g2_nand2_1 _44332_ (.Y(_13573_),
    .A(net5394),
    .B(_13572_));
 sg13g2_xnor2_1 _44333_ (.Y(_13574_),
    .A(net5448),
    .B(_13572_));
 sg13g2_nand2_1 _44334_ (.Y(_13575_),
    .A(_13543_),
    .B(_13559_));
 sg13g2_nor2_1 _44335_ (.A(_13544_),
    .B(_13575_),
    .Y(_13576_));
 sg13g2_a21oi_1 _44336_ (.A1(net5395),
    .A2(_13540_),
    .Y(_13577_),
    .B1(_13558_));
 sg13g2_nor2b_1 _44337_ (.A(_13576_),
    .B_N(_13577_),
    .Y(_13578_));
 sg13g2_o21ai_1 _44338_ (.B1(_13577_),
    .Y(_13579_),
    .A1(_13544_),
    .A2(_13575_));
 sg13g2_and4_1 _44339_ (.A(_13506_),
    .B(_13527_),
    .C(_13543_),
    .D(_13559_),
    .X(_13580_));
 sg13g2_inv_1 _44340_ (.Y(_13581_),
    .A(_13580_));
 sg13g2_o21ai_1 _44341_ (.B1(_13578_),
    .Y(_13582_),
    .A1(_13513_),
    .A2(_13581_));
 sg13g2_and2_1 _44342_ (.A(_13574_),
    .B(_13582_),
    .X(_13583_));
 sg13g2_xnor2_1 _44343_ (.Y(_13584_),
    .A(_13574_),
    .B(_13582_));
 sg13g2_nor2_1 _44344_ (.A(net5503),
    .B(_13572_),
    .Y(_13585_));
 sg13g2_a21oi_1 _44345_ (.A1(net5503),
    .A2(_13584_),
    .Y(_13586_),
    .B1(_13585_));
 sg13g2_nor2_1 _44346_ (.A(net5883),
    .B(_13557_),
    .Y(_13587_));
 sg13g2_a221oi_1 _44347_ (.B2(net5949),
    .C1(_13587_),
    .B1(_13586_),
    .A1(net5983),
    .Y(_13588_),
    .A2(_08743_));
 sg13g2_o21ai_1 _44348_ (.B1(net6876),
    .Y(_13589_),
    .A1(net5263),
    .A2(_08743_));
 sg13g2_a21oi_1 _44349_ (.A1(net5263),
    .A2(_13588_),
    .Y(_13590_),
    .B1(_13589_));
 sg13g2_a21o_1 _44350_ (.A2(net6414),
    .A1(net2196),
    .B1(_13590_),
    .X(_00908_));
 sg13g2_nand2_1 _44351_ (.Y(_13591_),
    .A(net5703),
    .B(_08718_));
 sg13g2_a21oi_1 _44352_ (.A1(_08737_),
    .A2(_13554_),
    .Y(_13592_),
    .B1(_08828_));
 sg13g2_xnor2_1 _44353_ (.Y(_13593_),
    .A(_08720_),
    .B(_13592_));
 sg13g2_o21ai_1 _44354_ (.B1(_13591_),
    .Y(_13594_),
    .A1(net5703),
    .A2(_13593_));
 sg13g2_or2_1 _44355_ (.X(_13595_),
    .B(_13594_),
    .A(net5394));
 sg13g2_nand2_1 _44356_ (.Y(_13596_),
    .A(net5394),
    .B(_13594_));
 sg13g2_xnor2_1 _44357_ (.Y(_13597_),
    .A(net5448),
    .B(_13594_));
 sg13g2_a21oi_1 _44358_ (.A1(net5394),
    .A2(_13572_),
    .Y(_13598_),
    .B1(_13583_));
 sg13g2_xor2_1 _44359_ (.B(_13598_),
    .A(_13597_),
    .X(_13599_));
 sg13g2_o21ai_1 _44360_ (.B1(net5949),
    .Y(_13600_),
    .A1(net5502),
    .A2(_13594_));
 sg13g2_a21oi_1 _44361_ (.A1(net5502),
    .A2(_13599_),
    .Y(_13601_),
    .B1(_13600_));
 sg13g2_a221oi_1 _44362_ (.B2(net5899),
    .C1(_13601_),
    .B1(_13572_),
    .A1(net5983),
    .Y(_13602_),
    .A2(_08730_));
 sg13g2_o21ai_1 _44363_ (.B1(net6876),
    .Y(_13603_),
    .A1(net5263),
    .A2(_08730_));
 sg13g2_a21oi_1 _44364_ (.A1(net5263),
    .A2(_13602_),
    .Y(_13604_),
    .B1(_13603_));
 sg13g2_a21o_1 _44365_ (.A2(net6414),
    .A1(net3065),
    .B1(_13604_),
    .X(_00909_));
 sg13g2_o21ai_1 _44366_ (.B1(_08719_),
    .Y(_13605_),
    .A1(_08720_),
    .A2(_13592_));
 sg13g2_xor2_1 _44367_ (.B(_13605_),
    .A(_08725_),
    .X(_13606_));
 sg13g2_nand2_1 _44368_ (.Y(_13607_),
    .A(net5703),
    .B(_08723_));
 sg13g2_o21ai_1 _44369_ (.B1(_13607_),
    .Y(_13608_),
    .A1(net5704),
    .A2(_13606_));
 sg13g2_nor2_1 _44370_ (.A(net5502),
    .B(_13608_),
    .Y(_13609_));
 sg13g2_nand2_1 _44371_ (.Y(_13610_),
    .A(net5394),
    .B(_13608_));
 sg13g2_xnor2_1 _44372_ (.Y(_13611_),
    .A(net5396),
    .B(_13608_));
 sg13g2_nand2_1 _44373_ (.Y(_13612_),
    .A(_13573_),
    .B(_13596_));
 sg13g2_o21ai_1 _44374_ (.B1(_13595_),
    .Y(_13613_),
    .A1(_13583_),
    .A2(_13612_));
 sg13g2_xnor2_1 _44375_ (.Y(_13614_),
    .A(_13611_),
    .B(_13613_));
 sg13g2_a21oi_1 _44376_ (.A1(net5502),
    .A2(_13614_),
    .Y(_13615_),
    .B1(_13609_));
 sg13g2_a22oi_1 _44377_ (.Y(_13616_),
    .B1(_13615_),
    .B2(net5227),
    .A2(_13594_),
    .A1(net5206));
 sg13g2_a22oi_1 _44378_ (.Y(_13617_),
    .B1(net5098),
    .B2(_08736_),
    .A2(net6414),
    .A1(net2191));
 sg13g2_o21ai_1 _44379_ (.B1(_13617_),
    .Y(_00910_),
    .A1(net6847),
    .A2(_13616_));
 sg13g2_a21oi_2 _44380_ (.B1(_08856_),
    .Y(_13618_),
    .A2(_10223_),
    .A1(net1094));
 sg13g2_o21ai_1 _44381_ (.B1(_08702_),
    .Y(_13619_),
    .A1(_08831_),
    .A2(_13618_));
 sg13g2_nor3_1 _44382_ (.A(_08702_),
    .B(_08831_),
    .C(_13618_),
    .Y(_13620_));
 sg13g2_nand3b_1 _44383_ (.B(net5752),
    .C(_13619_),
    .Y(_13621_),
    .A_N(_13620_));
 sg13g2_o21ai_1 _44384_ (.B1(_13621_),
    .Y(_13622_),
    .A1(net5752),
    .A2(_08700_));
 sg13g2_xnor2_1 _44385_ (.Y(_13623_),
    .A(net5396),
    .B(_13622_));
 sg13g2_o21ai_1 _44386_ (.B1(_13610_),
    .Y(_13624_),
    .A1(_13611_),
    .A2(_13613_));
 sg13g2_xor2_1 _44387_ (.B(_13624_),
    .A(_13623_),
    .X(_13625_));
 sg13g2_o21ai_1 _44388_ (.B1(net5949),
    .Y(_13626_),
    .A1(net5502),
    .A2(_13622_));
 sg13g2_a21oi_1 _44389_ (.A1(net5502),
    .A2(_13625_),
    .Y(_13627_),
    .B1(_13626_));
 sg13g2_a22oi_1 _44390_ (.Y(_13628_),
    .B1(_13608_),
    .B2(net5899),
    .A2(_08718_),
    .A1(net5983));
 sg13g2_nand2_1 _44391_ (.Y(_13629_),
    .A(net5263),
    .B(_13628_));
 sg13g2_nor2_1 _44392_ (.A(net5264),
    .B(_08718_),
    .Y(_13630_));
 sg13g2_o21ai_1 _44393_ (.B1(net6874),
    .Y(_13631_),
    .A1(_13627_),
    .A2(_13629_));
 sg13g2_nand2_1 _44394_ (.Y(_13632_),
    .A(net1782),
    .B(net6414));
 sg13g2_o21ai_1 _44395_ (.B1(_13632_),
    .Y(_00911_),
    .A1(_13630_),
    .A2(_13631_));
 sg13g2_o21ai_1 _44396_ (.B1(_13619_),
    .Y(_13633_),
    .A1(net5584),
    .A2(_08700_));
 sg13g2_xnor2_1 _44397_ (.Y(_13634_),
    .A(_08696_),
    .B(_13633_));
 sg13g2_nand2_1 _44398_ (.Y(_13635_),
    .A(net5705),
    .B(_08694_));
 sg13g2_o21ai_1 _44399_ (.B1(_13635_),
    .Y(_13636_),
    .A1(net5705),
    .A2(_13634_));
 sg13g2_nand2_1 _44400_ (.Y(_13637_),
    .A(net5396),
    .B(_13636_));
 sg13g2_xnor2_1 _44401_ (.Y(_13638_),
    .A(net5451),
    .B(_13636_));
 sg13g2_inv_2 _44402_ (.Y(_13639_),
    .A(_13638_));
 sg13g2_nor2_1 _44403_ (.A(_13611_),
    .B(_13623_),
    .Y(_13640_));
 sg13g2_nand2_1 _44404_ (.Y(_13641_),
    .A(_13574_),
    .B(_13597_));
 sg13g2_nor3_1 _44405_ (.A(_13611_),
    .B(_13623_),
    .C(_13641_),
    .Y(_13642_));
 sg13g2_nand3_1 _44406_ (.B(_13580_),
    .C(_13642_),
    .A(_13511_),
    .Y(_13643_));
 sg13g2_a22oi_1 _44407_ (.Y(_13644_),
    .B1(_13640_),
    .B2(_13612_),
    .A2(_13622_),
    .A1(net5394));
 sg13g2_nand2_1 _44408_ (.Y(_13645_),
    .A(_13579_),
    .B(_13642_));
 sg13g2_nand4_1 _44409_ (.B(_13643_),
    .C(_13644_),
    .A(_13610_),
    .Y(_13646_),
    .D(_13645_));
 sg13g2_inv_1 _44410_ (.Y(_13647_),
    .A(_13646_));
 sg13g2_and3_1 _44411_ (.X(_13648_),
    .A(_13512_),
    .B(_13580_),
    .C(_13642_));
 sg13g2_nand3_1 _44412_ (.B(_13580_),
    .C(_13642_),
    .A(_13512_),
    .Y(_13649_));
 sg13g2_o21ai_1 _44413_ (.B1(_13648_),
    .Y(_13650_),
    .A1(_13384_),
    .A2(_13386_));
 sg13g2_and2_1 _44414_ (.A(_13647_),
    .B(_13650_),
    .X(_13651_));
 sg13g2_xnor2_1 _44415_ (.Y(_13652_),
    .A(_13639_),
    .B(_13651_));
 sg13g2_o21ai_1 _44416_ (.B1(net5949),
    .Y(_13653_),
    .A1(net5502),
    .A2(_13636_));
 sg13g2_a21oi_1 _44417_ (.A1(net5502),
    .A2(_13652_),
    .Y(_13654_),
    .B1(_13653_));
 sg13g2_a221oi_1 _44418_ (.B2(net5899),
    .C1(_13654_),
    .B1(_13622_),
    .A1(net5983),
    .Y(_13655_),
    .A2(_08723_));
 sg13g2_a21oi_1 _44419_ (.A1(net5264),
    .A2(_13655_),
    .Y(_13656_),
    .B1(net6847));
 sg13g2_o21ai_1 _44420_ (.B1(_13656_),
    .Y(_13657_),
    .A1(net5265),
    .A2(_08723_));
 sg13g2_o21ai_1 _44421_ (.B1(_13657_),
    .Y(_00912_),
    .A1(_18122_),
    .A2(net6489));
 sg13g2_o21ai_1 _44422_ (.B1(_13637_),
    .Y(_13658_),
    .A1(_13639_),
    .A2(_13651_));
 sg13g2_nand2_1 _44423_ (.Y(_13659_),
    .A(net5705),
    .B(_08683_));
 sg13g2_a22oi_1 _44424_ (.Y(_13660_),
    .B1(_08833_),
    .B2(_13619_),
    .A2(_08695_),
    .A1(net5581));
 sg13g2_a221oi_1 _44425_ (.B2(_13619_),
    .C1(_08685_),
    .B1(_08833_),
    .A1(net5581),
    .Y(_13661_),
    .A2(_08695_));
 sg13g2_xor2_1 _44426_ (.B(_13660_),
    .A(_08685_),
    .X(_13662_));
 sg13g2_o21ai_1 _44427_ (.B1(_13659_),
    .Y(_13663_),
    .A1(net5705),
    .A2(_13662_));
 sg13g2_xnor2_1 _44428_ (.Y(_13664_),
    .A(net5451),
    .B(_13663_));
 sg13g2_xnor2_1 _44429_ (.Y(_13665_),
    .A(_13658_),
    .B(_13664_));
 sg13g2_o21ai_1 _44430_ (.B1(net5949),
    .Y(_13666_),
    .A1(net5505),
    .A2(_13663_));
 sg13g2_a21oi_1 _44431_ (.A1(net5505),
    .A2(_13665_),
    .Y(_13667_),
    .B1(_13666_));
 sg13g2_a221oi_1 _44432_ (.B2(net5894),
    .C1(_13667_),
    .B1(_13636_),
    .A1(net5983),
    .Y(_13668_),
    .A2(_08701_));
 sg13g2_o21ai_1 _44433_ (.B1(net6874),
    .Y(_13669_),
    .A1(net5265),
    .A2(_08701_));
 sg13g2_a21oi_1 _44434_ (.A1(net5265),
    .A2(_13668_),
    .Y(_13670_),
    .B1(_13669_));
 sg13g2_a21oi_1 _44435_ (.A1(net3111),
    .A2(net6414),
    .Y(_13671_),
    .B1(_13670_));
 sg13g2_inv_1 _44436_ (.Y(_00913_),
    .A(_13671_));
 sg13g2_or3_1 _44437_ (.A(_08684_),
    .B(_08689_),
    .C(_13661_),
    .X(_13672_));
 sg13g2_o21ai_1 _44438_ (.B1(_08689_),
    .Y(_13673_),
    .A1(_08684_),
    .A2(_13661_));
 sg13g2_nand2_1 _44439_ (.Y(_13674_),
    .A(net5705),
    .B(_08688_));
 sg13g2_a21o_1 _44440_ (.A2(_13673_),
    .A1(_13672_),
    .B1(net5705),
    .X(_13675_));
 sg13g2_nand2_1 _44441_ (.Y(_13676_),
    .A(_13674_),
    .B(_13675_));
 sg13g2_a21oi_1 _44442_ (.A1(_13674_),
    .A2(_13675_),
    .Y(_13677_),
    .B1(net5448));
 sg13g2_nand2_1 _44443_ (.Y(_13678_),
    .A(net5400),
    .B(_13676_));
 sg13g2_and3_2 _44444_ (.X(_13679_),
    .A(net5448),
    .B(_13674_),
    .C(_13675_));
 sg13g2_nor2_1 _44445_ (.A(_13677_),
    .B(_13679_),
    .Y(_13680_));
 sg13g2_o21ai_1 _44446_ (.B1(net5396),
    .Y(_13681_),
    .A1(_13636_),
    .A2(_13663_));
 sg13g2_o21ai_1 _44447_ (.B1(_13681_),
    .Y(_13682_),
    .A1(_13639_),
    .A2(_13651_));
 sg13g2_o21ai_1 _44448_ (.B1(_13682_),
    .Y(_13683_),
    .A1(net5396),
    .A2(_13663_));
 sg13g2_xor2_1 _44449_ (.B(_13683_),
    .A(_13680_),
    .X(_13684_));
 sg13g2_nand2_1 _44450_ (.Y(_13685_),
    .A(net5505),
    .B(_13684_));
 sg13g2_o21ai_1 _44451_ (.B1(_13685_),
    .Y(_13686_),
    .A1(net5505),
    .A2(_13676_));
 sg13g2_a22oi_1 _44452_ (.Y(_13687_),
    .B1(_13663_),
    .B2(net5206),
    .A2(_08694_),
    .A1(net5159));
 sg13g2_o21ai_1 _44453_ (.B1(_13687_),
    .Y(_13688_),
    .A1(net5152),
    .A2(_13686_));
 sg13g2_a22oi_1 _44454_ (.Y(_13689_),
    .B1(net6874),
    .B2(_13688_),
    .A2(net6414),
    .A1(net2707));
 sg13g2_inv_1 _44455_ (.Y(_00914_),
    .A(_13689_));
 sg13g2_o21ai_1 _44456_ (.B1(_08704_),
    .Y(_13690_),
    .A1(_08831_),
    .A2(_13618_));
 sg13g2_a21oi_1 _44457_ (.A1(_08835_),
    .A2(_13690_),
    .Y(_13691_),
    .B1(_08678_));
 sg13g2_and3_1 _44458_ (.X(_13692_),
    .A(_08678_),
    .B(_08835_),
    .C(_13690_));
 sg13g2_nor3_1 _44459_ (.A(net5697),
    .B(_13691_),
    .C(_13692_),
    .Y(_13693_));
 sg13g2_a21oi_2 _44460_ (.B1(_13693_),
    .Y(_13694_),
    .A2(_08676_),
    .A1(net5704));
 sg13g2_or2_1 _44461_ (.X(_13695_),
    .B(_13694_),
    .A(net5443));
 sg13g2_xnor2_1 _44462_ (.Y(_13696_),
    .A(net5443),
    .B(_13694_));
 sg13g2_o21ai_1 _44463_ (.B1(_13678_),
    .Y(_13697_),
    .A1(_13679_),
    .A2(_13683_));
 sg13g2_xnor2_1 _44464_ (.Y(_13698_),
    .A(_13696_),
    .B(_13697_));
 sg13g2_a21oi_1 _44465_ (.A1(net5558),
    .A2(_13694_),
    .Y(_13699_),
    .B1(net5923));
 sg13g2_o21ai_1 _44466_ (.B1(_13699_),
    .Y(_13700_),
    .A1(net5558),
    .A2(_13698_));
 sg13g2_a22oi_1 _44467_ (.Y(_13701_),
    .B1(_13676_),
    .B2(net5894),
    .A2(_08683_),
    .A1(net5979));
 sg13g2_and3_1 _44468_ (.X(_13702_),
    .A(net5265),
    .B(_13700_),
    .C(_13701_));
 sg13g2_o21ai_1 _44469_ (.B1(net6874),
    .Y(_13703_),
    .A1(net5265),
    .A2(_08683_));
 sg13g2_nand2_1 _44470_ (.Y(_13704_),
    .A(net2074),
    .B(net6415));
 sg13g2_o21ai_1 _44471_ (.B1(_13704_),
    .Y(_00915_),
    .A1(_13702_),
    .A2(_13703_));
 sg13g2_or2_1 _44472_ (.X(_13705_),
    .B(_08670_),
    .A(net5747));
 sg13g2_a21oi_1 _44473_ (.A1(net5638),
    .A2(_08676_),
    .Y(_13706_),
    .B1(_13691_));
 sg13g2_xnor2_1 _44474_ (.Y(_13707_),
    .A(_08671_),
    .B(_13706_));
 sg13g2_o21ai_1 _44475_ (.B1(_13705_),
    .Y(_13708_),
    .A1(net5697),
    .A2(_13707_));
 sg13g2_nor2_1 _44476_ (.A(net5493),
    .B(_13708_),
    .Y(_13709_));
 sg13g2_nand2_1 _44477_ (.Y(_13710_),
    .A(net5388),
    .B(_13708_));
 sg13g2_xnor2_1 _44478_ (.Y(_13711_),
    .A(net5388),
    .B(_13708_));
 sg13g2_or4_1 _44479_ (.A(_13677_),
    .B(_13679_),
    .C(_13681_),
    .D(_13696_),
    .X(_13712_));
 sg13g2_nand3_1 _44480_ (.B(_13695_),
    .C(_13712_),
    .A(_13678_),
    .Y(_13713_));
 sg13g2_nand2_1 _44481_ (.Y(_13714_),
    .A(_13638_),
    .B(_13664_));
 sg13g2_or4_1 _44482_ (.A(_13677_),
    .B(_13679_),
    .C(_13696_),
    .D(_13714_),
    .X(_13715_));
 sg13g2_a21oi_1 _44483_ (.A1(_13647_),
    .A2(_13650_),
    .Y(_13716_),
    .B1(_13715_));
 sg13g2_or2_1 _44484_ (.X(_13717_),
    .B(_13716_),
    .A(_13713_));
 sg13g2_nand2b_1 _44485_ (.Y(_13718_),
    .B(_13717_),
    .A_N(_13711_));
 sg13g2_xor2_1 _44486_ (.B(_13717_),
    .A(_13711_),
    .X(_13719_));
 sg13g2_a21oi_1 _44487_ (.A1(net5493),
    .A2(_13719_),
    .Y(_13720_),
    .B1(_13709_));
 sg13g2_nand2_1 _44488_ (.Y(_13721_),
    .A(net5224),
    .B(_13720_));
 sg13g2_o21ai_1 _44489_ (.B1(_13721_),
    .Y(_13722_),
    .A1(net5122),
    .A2(_13694_));
 sg13g2_a22oi_1 _44490_ (.Y(_13723_),
    .B1(_13722_),
    .B2(net6875),
    .A2(_08688_),
    .A1(net5099));
 sg13g2_o21ai_1 _44491_ (.B1(_13723_),
    .Y(_00916_),
    .A1(_18120_),
    .A2(net6489));
 sg13g2_nand2_1 _44492_ (.Y(_13724_),
    .A(net2031),
    .B(net6414));
 sg13g2_nor2_1 _44493_ (.A(net5747),
    .B(_08664_),
    .Y(_13725_));
 sg13g2_a21oi_1 _44494_ (.A1(_08672_),
    .A2(_13691_),
    .Y(_13726_),
    .B1(_08838_));
 sg13g2_xnor2_1 _44495_ (.Y(_13727_),
    .A(_08666_),
    .B(_13726_));
 sg13g2_a21oi_2 _44496_ (.B1(_13725_),
    .Y(_13728_),
    .A2(_13727_),
    .A1(net5747));
 sg13g2_inv_1 _44497_ (.Y(_13729_),
    .A(_13728_));
 sg13g2_xnor2_1 _44498_ (.Y(_13730_),
    .A(net5388),
    .B(_13728_));
 sg13g2_nand2_1 _44499_ (.Y(_13731_),
    .A(_13710_),
    .B(_13718_));
 sg13g2_xor2_1 _44500_ (.B(_13731_),
    .A(_13730_),
    .X(_13732_));
 sg13g2_o21ai_1 _44501_ (.B1(net5945),
    .Y(_13733_),
    .A1(net5494),
    .A2(_13728_));
 sg13g2_a21oi_1 _44502_ (.A1(net5493),
    .A2(_13732_),
    .Y(_13734_),
    .B1(_13733_));
 sg13g2_a221oi_1 _44503_ (.B2(net5895),
    .C1(_13734_),
    .B1(_13708_),
    .A1(net5979),
    .Y(_13735_),
    .A2(_08676_));
 sg13g2_and2_1 _44504_ (.A(net5265),
    .B(_13735_),
    .X(_13736_));
 sg13g2_o21ai_1 _44505_ (.B1(net6874),
    .Y(_13737_),
    .A1(net5265),
    .A2(_08676_));
 sg13g2_o21ai_1 _44506_ (.B1(_13724_),
    .Y(_00917_),
    .A1(_13736_),
    .A2(_13737_));
 sg13g2_nor2_1 _44507_ (.A(_18119_),
    .B(net6490),
    .Y(_13738_));
 sg13g2_nand2_1 _44508_ (.Y(_13739_),
    .A(net5698),
    .B(_08653_));
 sg13g2_o21ai_1 _44509_ (.B1(_08665_),
    .Y(_13740_),
    .A1(_08666_),
    .A2(_13726_));
 sg13g2_xnor2_1 _44510_ (.Y(_13741_),
    .A(_08655_),
    .B(_13740_));
 sg13g2_o21ai_1 _44511_ (.B1(_13739_),
    .Y(_13742_),
    .A1(net5698),
    .A2(_13741_));
 sg13g2_and2_1 _44512_ (.A(net5388),
    .B(_13742_),
    .X(_13743_));
 sg13g2_xnor2_1 _44513_ (.Y(_13744_),
    .A(net5443),
    .B(_13742_));
 sg13g2_o21ai_1 _44514_ (.B1(net5388),
    .Y(_13745_),
    .A1(_13708_),
    .A2(_13728_));
 sg13g2_a22oi_1 _44515_ (.Y(_13746_),
    .B1(_13745_),
    .B2(_13718_),
    .A2(_13729_),
    .A1(net5443));
 sg13g2_xnor2_1 _44516_ (.Y(_13747_),
    .A(_13744_),
    .B(_13746_));
 sg13g2_nor2_1 _44517_ (.A(net5494),
    .B(_13742_),
    .Y(_13748_));
 sg13g2_a21oi_1 _44518_ (.A1(net5494),
    .A2(_13747_),
    .Y(_13749_),
    .B1(_13748_));
 sg13g2_nor2_1 _44519_ (.A(net6004),
    .B(_08670_),
    .Y(_13750_));
 sg13g2_a221oi_1 _44520_ (.B2(net5945),
    .C1(_13750_),
    .B1(_13749_),
    .A1(net5894),
    .Y(_13751_),
    .A2(_13728_));
 sg13g2_nand3_1 _44521_ (.B(net5316),
    .C(_08670_),
    .A(net5320),
    .Y(_13752_));
 sg13g2_a21oi_1 _44522_ (.A1(net5262),
    .A2(_13751_),
    .Y(_13753_),
    .B1(net6843));
 sg13g2_a21o_1 _44523_ (.A2(_13753_),
    .A1(_13752_),
    .B1(_13738_),
    .X(_00918_));
 sg13g2_nand2_1 _44524_ (.Y(_13754_),
    .A(net2095),
    .B(net6415));
 sg13g2_o21ai_1 _44525_ (.B1(_08705_),
    .Y(_13755_),
    .A1(_08831_),
    .A2(_13618_));
 sg13g2_nand2_1 _44526_ (.Y(_13756_),
    .A(_08840_),
    .B(_13755_));
 sg13g2_a21oi_1 _44527_ (.A1(_08840_),
    .A2(_13755_),
    .Y(_13757_),
    .B1(_08648_));
 sg13g2_nor2b_1 _44528_ (.A(_13756_),
    .B_N(_08648_),
    .Y(_13758_));
 sg13g2_nor3_1 _44529_ (.A(net5696),
    .B(_13757_),
    .C(_13758_),
    .Y(_13759_));
 sg13g2_a21oi_1 _44530_ (.A1(net5697),
    .A2(_08646_),
    .Y(_13760_),
    .B1(_13759_));
 sg13g2_inv_1 _44531_ (.Y(_13761_),
    .A(_13760_));
 sg13g2_xnor2_1 _44532_ (.Y(_13762_),
    .A(net5389),
    .B(_13760_));
 sg13g2_a21oi_1 _44533_ (.A1(_13744_),
    .A2(_13746_),
    .Y(_13763_),
    .B1(_13743_));
 sg13g2_xnor2_1 _44534_ (.Y(_13764_),
    .A(_13762_),
    .B(_13763_));
 sg13g2_a21oi_1 _44535_ (.A1(net5553),
    .A2(_13760_),
    .Y(_13765_),
    .B1(net5922));
 sg13g2_o21ai_1 _44536_ (.B1(_13765_),
    .Y(_13766_),
    .A1(net5553),
    .A2(_13764_));
 sg13g2_a22oi_1 _44537_ (.Y(_13767_),
    .B1(_13742_),
    .B2(net5895),
    .A2(_08664_),
    .A1(net5979));
 sg13g2_and3_1 _44538_ (.X(_13768_),
    .A(net5261),
    .B(_13766_),
    .C(_13767_));
 sg13g2_o21ai_1 _44539_ (.B1(net6874),
    .Y(_13769_),
    .A1(net5262),
    .A2(_08664_));
 sg13g2_o21ai_1 _44540_ (.B1(_13754_),
    .Y(_00919_),
    .A1(_13768_),
    .A2(_13769_));
 sg13g2_a21oi_1 _44541_ (.A1(net5628),
    .A2(_08646_),
    .Y(_13770_),
    .B1(_13757_));
 sg13g2_xnor2_1 _44542_ (.Y(_13771_),
    .A(_08642_),
    .B(_13770_));
 sg13g2_nor2_1 _44543_ (.A(net5696),
    .B(_13771_),
    .Y(_13772_));
 sg13g2_a21oi_2 _44544_ (.B1(_13772_),
    .Y(_13773_),
    .A2(_08640_),
    .A1(net5697));
 sg13g2_nor2_1 _44545_ (.A(net5493),
    .B(_13773_),
    .Y(_13774_));
 sg13g2_nand2_1 _44546_ (.Y(_13775_),
    .A(net5388),
    .B(_13773_));
 sg13g2_xnor2_1 _44547_ (.Y(_13776_),
    .A(net5388),
    .B(_13773_));
 sg13g2_inv_1 _44548_ (.Y(_13777_),
    .A(_13776_));
 sg13g2_nor2_1 _44549_ (.A(_13711_),
    .B(_13730_),
    .Y(_13778_));
 sg13g2_nand3_1 _44550_ (.B(_13762_),
    .C(_13778_),
    .A(_13744_),
    .Y(_13779_));
 sg13g2_nand4_1 _44551_ (.B(_13744_),
    .C(_13762_),
    .A(_13713_),
    .Y(_13780_),
    .D(_13778_));
 sg13g2_nand3b_1 _44552_ (.B(_13762_),
    .C(_13744_),
    .Y(_13781_),
    .A_N(_13745_));
 sg13g2_o21ai_1 _44553_ (.B1(net5389),
    .Y(_13782_),
    .A1(_13742_),
    .A2(_13761_));
 sg13g2_nand3_1 _44554_ (.B(_13781_),
    .C(_13782_),
    .A(_13780_),
    .Y(_13783_));
 sg13g2_or2_1 _44555_ (.X(_13784_),
    .B(_13779_),
    .A(_13715_));
 sg13g2_a21oi_1 _44556_ (.A1(_13647_),
    .A2(_13650_),
    .Y(_13785_),
    .B1(_13784_));
 sg13g2_or2_1 _44557_ (.X(_13786_),
    .B(_13785_),
    .A(_13783_));
 sg13g2_nand2_1 _44558_ (.Y(_13787_),
    .A(_13777_),
    .B(_13786_));
 sg13g2_xnor2_1 _44559_ (.Y(_13788_),
    .A(_13777_),
    .B(_13786_));
 sg13g2_a21oi_1 _44560_ (.A1(net5494),
    .A2(_13788_),
    .Y(_13789_),
    .B1(_13774_));
 sg13g2_a22oi_1 _44561_ (.Y(_13790_),
    .B1(_13789_),
    .B2(net5224),
    .A2(_13761_),
    .A1(net5203));
 sg13g2_a22oi_1 _44562_ (.Y(_13791_),
    .B1(net5097),
    .B2(_08653_),
    .A2(net6415),
    .A1(net2654));
 sg13g2_o21ai_1 _44563_ (.B1(_13791_),
    .Y(_00920_),
    .A1(net6843),
    .A2(_13790_));
 sg13g2_nand2_1 _44564_ (.Y(_13792_),
    .A(net2314),
    .B(net6407));
 sg13g2_nor2_1 _44565_ (.A(net5746),
    .B(_08628_),
    .Y(_13793_));
 sg13g2_a21oi_1 _44566_ (.A1(_08642_),
    .A2(_13757_),
    .Y(_13794_),
    .B1(_08842_));
 sg13g2_xnor2_1 _44567_ (.Y(_13795_),
    .A(_08630_),
    .B(_13794_));
 sg13g2_a21oi_2 _44568_ (.B1(_13793_),
    .Y(_13796_),
    .A2(_13795_),
    .A1(net5746));
 sg13g2_inv_1 _44569_ (.Y(_13797_),
    .A(_13796_));
 sg13g2_xnor2_1 _44570_ (.Y(_13798_),
    .A(net5388),
    .B(_13796_));
 sg13g2_nand2_1 _44571_ (.Y(_13799_),
    .A(_13775_),
    .B(_13787_));
 sg13g2_or2_1 _44572_ (.X(_13800_),
    .B(_13799_),
    .A(_13798_));
 sg13g2_a21oi_1 _44573_ (.A1(_13798_),
    .A2(_13799_),
    .Y(_13801_),
    .B1(net5554));
 sg13g2_a221oi_1 _44574_ (.B2(_13801_),
    .C1(net5152),
    .B1(_13800_),
    .A1(net5554),
    .Y(_13802_),
    .A2(_13797_));
 sg13g2_a221oi_1 _44575_ (.B2(net5204),
    .C1(_13802_),
    .B1(_13773_),
    .A1(net5158),
    .Y(_13803_),
    .A2(_08646_));
 sg13g2_o21ai_1 _44576_ (.B1(_13792_),
    .Y(_00921_),
    .A1(net6844),
    .A2(_13803_));
 sg13g2_nand2_1 _44577_ (.Y(_13804_),
    .A(net5697),
    .B(_08633_));
 sg13g2_o21ai_1 _44578_ (.B1(_08629_),
    .Y(_13805_),
    .A1(_08630_),
    .A2(_13794_));
 sg13g2_xnor2_1 _44579_ (.Y(_13806_),
    .A(_08636_),
    .B(_13805_));
 sg13g2_o21ai_1 _44580_ (.B1(_13804_),
    .Y(_13807_),
    .A1(net5697),
    .A2(_13806_));
 sg13g2_inv_1 _44581_ (.Y(_13808_),
    .A(_13807_));
 sg13g2_nor2_1 _44582_ (.A(net5442),
    .B(_13807_),
    .Y(_13809_));
 sg13g2_nand2_1 _44583_ (.Y(_13810_),
    .A(net5442),
    .B(_13807_));
 sg13g2_xnor2_1 _44584_ (.Y(_13811_),
    .A(net5443),
    .B(_13807_));
 sg13g2_o21ai_1 _44585_ (.B1(net5390),
    .Y(_13812_),
    .A1(_13773_),
    .A2(_13796_));
 sg13g2_a22oi_1 _44586_ (.Y(_13813_),
    .B1(_13812_),
    .B2(_13787_),
    .A2(_13797_),
    .A1(net5444));
 sg13g2_xnor2_1 _44587_ (.Y(_13814_),
    .A(_13811_),
    .B(_13813_));
 sg13g2_a21oi_1 _44588_ (.A1(net5553),
    .A2(_13807_),
    .Y(_13815_),
    .B1(net5922));
 sg13g2_o21ai_1 _44589_ (.B1(_13815_),
    .Y(_13816_),
    .A1(net5554),
    .A2(_13814_));
 sg13g2_nor2_1 _44590_ (.A(net6004),
    .B(_08640_),
    .Y(_13817_));
 sg13g2_a21oi_1 _44591_ (.A1(net5894),
    .A2(_13796_),
    .Y(_13818_),
    .B1(_13817_));
 sg13g2_nand3_1 _44592_ (.B(_13816_),
    .C(_13818_),
    .A(net5261),
    .Y(_13819_));
 sg13g2_nand3_1 _44593_ (.B(net5316),
    .C(_08640_),
    .A(net5320),
    .Y(_13820_));
 sg13g2_nand3_1 _44594_ (.B(_13819_),
    .C(_13820_),
    .A(net6874),
    .Y(_13821_));
 sg13g2_o21ai_1 _44595_ (.B1(_13821_),
    .Y(_00922_),
    .A1(_18117_),
    .A2(net6490));
 sg13g2_a21oi_1 _44596_ (.A1(_08649_),
    .A2(_13756_),
    .Y(_13822_),
    .B1(_08844_));
 sg13g2_nor2_1 _44597_ (.A(_08616_),
    .B(_13822_),
    .Y(_13823_));
 sg13g2_xnor2_1 _44598_ (.Y(_13824_),
    .A(_08616_),
    .B(_13822_));
 sg13g2_nand2_1 _44599_ (.Y(_13825_),
    .A(net5746),
    .B(_13824_));
 sg13g2_o21ai_1 _44600_ (.B1(_13825_),
    .Y(_13826_),
    .A1(net5746),
    .A2(_08615_));
 sg13g2_inv_1 _44601_ (.Y(_13827_),
    .A(_13826_));
 sg13g2_xnor2_1 _44602_ (.Y(_13828_),
    .A(net5443),
    .B(_13826_));
 sg13g2_a21oi_1 _44603_ (.A1(_13810_),
    .A2(_13813_),
    .Y(_13829_),
    .B1(_13809_));
 sg13g2_xor2_1 _44604_ (.B(_13829_),
    .A(_13828_),
    .X(_13830_));
 sg13g2_a21oi_1 _44605_ (.A1(net5554),
    .A2(_13826_),
    .Y(_13831_),
    .B1(net5922));
 sg13g2_o21ai_1 _44606_ (.B1(_13831_),
    .Y(_13832_),
    .A1(net5554),
    .A2(_13830_));
 sg13g2_a22oi_1 _44607_ (.Y(_13833_),
    .B1(_13808_),
    .B2(net5894),
    .A2(_08628_),
    .A1(net5980));
 sg13g2_and3_1 _44608_ (.X(_13834_),
    .A(net5266),
    .B(_13832_),
    .C(_13833_));
 sg13g2_o21ai_1 _44609_ (.B1(net6874),
    .Y(_13835_),
    .A1(net5262),
    .A2(_08628_));
 sg13g2_nand2_1 _44610_ (.Y(_13836_),
    .A(net2440),
    .B(net6407));
 sg13g2_o21ai_1 _44611_ (.B1(_13836_),
    .Y(_00923_),
    .A1(_13834_),
    .A2(_13835_));
 sg13g2_nand2_1 _44612_ (.Y(_13837_),
    .A(net5696),
    .B(_08620_));
 sg13g2_a21oi_1 _44613_ (.A1(net5627),
    .A2(_08615_),
    .Y(_13838_),
    .B1(_13823_));
 sg13g2_xor2_1 _44614_ (.B(_13838_),
    .A(_08621_),
    .X(_13839_));
 sg13g2_o21ai_1 _44615_ (.B1(_13837_),
    .Y(_13840_),
    .A1(net5696),
    .A2(_13839_));
 sg13g2_nor2_1 _44616_ (.A(net5493),
    .B(_13840_),
    .Y(_13841_));
 sg13g2_nand2_1 _44617_ (.Y(_13842_),
    .A(net5389),
    .B(_13840_));
 sg13g2_xnor2_1 _44618_ (.Y(_13843_),
    .A(net5389),
    .B(_13840_));
 sg13g2_nor3_1 _44619_ (.A(_13811_),
    .B(_13812_),
    .C(_13828_),
    .Y(_13844_));
 sg13g2_a21oi_1 _44620_ (.A1(_13807_),
    .A2(_13826_),
    .Y(_13845_),
    .B1(net5443));
 sg13g2_or2_1 _44621_ (.X(_13846_),
    .B(_13845_),
    .A(_13844_));
 sg13g2_inv_1 _44622_ (.Y(_13847_),
    .A(_13846_));
 sg13g2_nor4_1 _44623_ (.A(_13776_),
    .B(_13798_),
    .C(_13811_),
    .D(_13828_),
    .Y(_13848_));
 sg13g2_inv_1 _44624_ (.Y(_13849_),
    .A(_13848_));
 sg13g2_o21ai_1 _44625_ (.B1(_13848_),
    .Y(_13850_),
    .A1(_13783_),
    .A2(_13785_));
 sg13g2_a21o_1 _44626_ (.A2(_13850_),
    .A1(_13847_),
    .B1(_13843_),
    .X(_13851_));
 sg13g2_nand3_1 _44627_ (.B(_13847_),
    .C(_13850_),
    .A(_13843_),
    .Y(_13852_));
 sg13g2_a21oi_1 _44628_ (.A1(_13851_),
    .A2(_13852_),
    .Y(_13853_),
    .B1(net5553));
 sg13g2_nor2_1 _44629_ (.A(_13841_),
    .B(_13853_),
    .Y(_13854_));
 sg13g2_a22oi_1 _44630_ (.Y(_13855_),
    .B1(_13854_),
    .B2(net5224),
    .A2(_13827_),
    .A1(net5204));
 sg13g2_a22oi_1 _44631_ (.Y(_13856_),
    .B1(net5097),
    .B2(_08634_),
    .A2(net6408),
    .A1(net1483));
 sg13g2_o21ai_1 _44632_ (.B1(_13856_),
    .Y(_00924_),
    .A1(net6843),
    .A2(_13855_));
 sg13g2_and2_1 _44633_ (.A(net5696),
    .B(_08600_),
    .X(_13857_));
 sg13g2_o21ai_1 _44634_ (.B1(_08846_),
    .Y(_13858_),
    .A1(_08623_),
    .A2(_13822_));
 sg13g2_xnor2_1 _44635_ (.Y(_13859_),
    .A(_08603_),
    .B(_13858_));
 sg13g2_a21oi_2 _44636_ (.B1(_13857_),
    .Y(_13860_),
    .A2(_13859_),
    .A1(net5746));
 sg13g2_nor2_1 _44637_ (.A(net5442),
    .B(_13860_),
    .Y(_13861_));
 sg13g2_xnor2_1 _44638_ (.Y(_13862_),
    .A(net5442),
    .B(_13860_));
 sg13g2_nand2_1 _44639_ (.Y(_13863_),
    .A(_13842_),
    .B(_13851_));
 sg13g2_xnor2_1 _44640_ (.Y(_13864_),
    .A(_13862_),
    .B(_13863_));
 sg13g2_a21oi_1 _44641_ (.A1(net5553),
    .A2(_13860_),
    .Y(_13865_),
    .B1(net5922));
 sg13g2_o21ai_1 _44642_ (.B1(_13865_),
    .Y(_13866_),
    .A1(net5553),
    .A2(_13864_));
 sg13g2_a22oi_1 _44643_ (.Y(_13867_),
    .B1(_13840_),
    .B2(net5894),
    .A2(_08615_),
    .A1(net5979));
 sg13g2_and3_1 _44644_ (.X(_13868_),
    .A(net5261),
    .B(_13866_),
    .C(_13867_));
 sg13g2_o21ai_1 _44645_ (.B1(net6872),
    .Y(_13869_),
    .A1(net5261),
    .A2(_08615_));
 sg13g2_nand2_1 _44646_ (.Y(_13870_),
    .A(net2687),
    .B(net6407));
 sg13g2_o21ai_1 _44647_ (.B1(_13870_),
    .Y(_00925_),
    .A1(_13868_),
    .A2(_13869_));
 sg13g2_nand2b_1 _44648_ (.Y(_13871_),
    .B(net5204),
    .A_N(_13860_));
 sg13g2_nor2_1 _44649_ (.A(net5746),
    .B(_08607_),
    .Y(_13872_));
 sg13g2_a21oi_1 _44650_ (.A1(_08602_),
    .A2(_13858_),
    .Y(_13873_),
    .B1(_08601_));
 sg13g2_xnor2_1 _44651_ (.Y(_13874_),
    .A(_08610_),
    .B(_13873_));
 sg13g2_a21oi_2 _44652_ (.B1(_13872_),
    .Y(_13875_),
    .A2(_13874_),
    .A1(net5746));
 sg13g2_inv_1 _44653_ (.Y(_13876_),
    .A(_13875_));
 sg13g2_nor2_1 _44654_ (.A(net5442),
    .B(_13875_),
    .Y(_13877_));
 sg13g2_nand2_1 _44655_ (.Y(_13878_),
    .A(net5442),
    .B(_13875_));
 sg13g2_xnor2_1 _44656_ (.Y(_13879_),
    .A(net5442),
    .B(_13875_));
 sg13g2_a21oi_1 _44657_ (.A1(net5389),
    .A2(_13840_),
    .Y(_13880_),
    .B1(_13861_));
 sg13g2_a22oi_1 _44658_ (.Y(_13881_),
    .B1(_13880_),
    .B2(_13851_),
    .A2(_13860_),
    .A1(net5442));
 sg13g2_xnor2_1 _44659_ (.Y(_13882_),
    .A(_13879_),
    .B(_13881_));
 sg13g2_o21ai_1 _44660_ (.B1(net5225),
    .Y(_13883_),
    .A1(net5553),
    .A2(_13882_));
 sg13g2_a21o_1 _44661_ (.A2(_13875_),
    .A1(net5553),
    .B1(_13883_),
    .X(_13884_));
 sg13g2_a21oi_1 _44662_ (.A1(_13871_),
    .A2(_13884_),
    .Y(_13885_),
    .B1(net6843));
 sg13g2_a22oi_1 _44663_ (.Y(_13886_),
    .B1(net5097),
    .B2(_08620_),
    .A2(net6407),
    .A1(net3754));
 sg13g2_nand2b_1 _44664_ (.Y(_00926_),
    .B(_13886_),
    .A_N(_13885_));
 sg13g2_nor2_1 _44665_ (.A(net5746),
    .B(_10524_),
    .Y(_13887_));
 sg13g2_a21o_2 _44666_ (.A2(net5475),
    .A1(net5476),
    .B1(_10526_),
    .X(_13888_));
 sg13g2_nand3_1 _44667_ (.B(net5475),
    .C(_10526_),
    .A(net5476),
    .Y(_13889_));
 sg13g2_a21oi_1 _44668_ (.A1(_13888_),
    .A2(_13889_),
    .Y(_13890_),
    .B1(net5696));
 sg13g2_nor2_2 _44669_ (.A(_13887_),
    .B(_13890_),
    .Y(_13891_));
 sg13g2_nand2_1 _44670_ (.Y(_13892_),
    .A(net5389),
    .B(_13891_));
 sg13g2_xnor2_1 _44671_ (.Y(_13893_),
    .A(net5389),
    .B(_13891_));
 sg13g2_a21oi_1 _44672_ (.A1(_13878_),
    .A2(_13881_),
    .Y(_13894_),
    .B1(_13877_));
 sg13g2_xnor2_1 _44673_ (.Y(_13895_),
    .A(_13893_),
    .B(_13894_));
 sg13g2_o21ai_1 _44674_ (.B1(net5945),
    .Y(_13896_),
    .A1(net5493),
    .A2(_13891_));
 sg13g2_a21oi_1 _44675_ (.A1(net5493),
    .A2(_13895_),
    .Y(_13897_),
    .B1(_13896_));
 sg13g2_a22oi_1 _44676_ (.Y(_13898_),
    .B1(_13876_),
    .B2(net5894),
    .A2(_08600_),
    .A1(net5980));
 sg13g2_nand2_1 _44677_ (.Y(_13899_),
    .A(net5261),
    .B(_13898_));
 sg13g2_nor2_1 _44678_ (.A(net5262),
    .B(_08600_),
    .Y(_13900_));
 sg13g2_o21ai_1 _44679_ (.B1(net6873),
    .Y(_13901_),
    .A1(_13897_),
    .A2(_13899_));
 sg13g2_nand2_1 _44680_ (.Y(_13902_),
    .A(net2548),
    .B(net6407));
 sg13g2_o21ai_1 _44681_ (.B1(_13902_),
    .Y(_00927_),
    .A1(_13900_),
    .A2(_13901_));
 sg13g2_nand2_1 _44682_ (.Y(_13903_),
    .A(net5696),
    .B(_10529_));
 sg13g2_nand2_1 _44683_ (.Y(_13904_),
    .A(_10525_),
    .B(_13888_));
 sg13g2_xor2_1 _44684_ (.B(_13904_),
    .A(_10531_),
    .X(_13905_));
 sg13g2_o21ai_1 _44685_ (.B1(_13903_),
    .Y(_13906_),
    .A1(net5696),
    .A2(_13905_));
 sg13g2_nand2_1 _44686_ (.Y(_13907_),
    .A(net5385),
    .B(_13906_));
 sg13g2_xnor2_1 _44687_ (.Y(_13908_),
    .A(net5441),
    .B(_13906_));
 sg13g2_or4_1 _44688_ (.A(_13843_),
    .B(_13862_),
    .C(_13879_),
    .D(_13893_),
    .X(_13909_));
 sg13g2_nor3_1 _44689_ (.A(_13784_),
    .B(_13849_),
    .C(_13909_),
    .Y(_13910_));
 sg13g2_nor4_1 _44690_ (.A(_13649_),
    .B(_13784_),
    .C(_13849_),
    .D(_13909_),
    .Y(_13911_));
 sg13g2_and2_1 _44691_ (.A(_13384_),
    .B(_13911_),
    .X(_13912_));
 sg13g2_nand3b_1 _44692_ (.B(_13783_),
    .C(_13848_),
    .Y(_13913_),
    .A_N(_13909_));
 sg13g2_nand2b_1 _44693_ (.Y(_13914_),
    .B(_13846_),
    .A_N(_13909_));
 sg13g2_nor3_1 _44694_ (.A(_13879_),
    .B(_13880_),
    .C(_13893_),
    .Y(_13915_));
 sg13g2_nor2_1 _44695_ (.A(_13877_),
    .B(_13915_),
    .Y(_13916_));
 sg13g2_nand4_1 _44696_ (.B(_13913_),
    .C(_13914_),
    .A(_13892_),
    .Y(_13917_),
    .D(_13916_));
 sg13g2_and2_1 _44697_ (.A(_13646_),
    .B(_13910_),
    .X(_13918_));
 sg13g2_nor3_2 _44698_ (.A(_13912_),
    .B(_13917_),
    .C(_13918_),
    .Y(_13919_));
 sg13g2_or3_1 _44699_ (.A(_13912_),
    .B(_13917_),
    .C(_13918_),
    .X(_13920_));
 sg13g2_nand2b_1 _44700_ (.Y(_13921_),
    .B(_13911_),
    .A_N(_13385_));
 sg13g2_a21oi_1 _44701_ (.A1(_12837_),
    .A2(net1064),
    .Y(_13922_),
    .B1(_13921_));
 sg13g2_a21o_2 _44702_ (.A2(net1064),
    .A1(_12837_),
    .B1(_13921_),
    .X(_13923_));
 sg13g2_nand2_2 _44703_ (.Y(_13924_),
    .A(_13919_),
    .B(_13923_));
 sg13g2_nand2_1 _44704_ (.Y(_13925_),
    .A(_13908_),
    .B(_13924_));
 sg13g2_xnor2_1 _44705_ (.Y(_13926_),
    .A(_13908_),
    .B(_13924_));
 sg13g2_o21ai_1 _44706_ (.B1(net5945),
    .Y(_13927_),
    .A1(net5491),
    .A2(_13906_));
 sg13g2_a21oi_1 _44707_ (.A1(net5493),
    .A2(_13926_),
    .Y(_13928_),
    .B1(_13927_));
 sg13g2_a221oi_1 _44708_ (.B2(net5894),
    .C1(_13928_),
    .B1(_13891_),
    .A1(net5979),
    .Y(_13929_),
    .A2(_08608_));
 sg13g2_o21ai_1 _44709_ (.B1(net6872),
    .Y(_13930_),
    .A1(net5261),
    .A2(_08608_));
 sg13g2_a21oi_1 _44710_ (.A1(net5261),
    .A2(_13929_),
    .Y(_13931_),
    .B1(_13930_));
 sg13g2_a21oi_1 _44711_ (.A1(net3539),
    .A2(net6408),
    .Y(_13932_),
    .B1(_13931_));
 sg13g2_inv_1 _44712_ (.Y(_00928_),
    .A(_13932_));
 sg13g2_nand2_1 _44713_ (.Y(_13933_),
    .A(net5695),
    .B(_10516_));
 sg13g2_a22oi_1 _44714_ (.Y(_13934_),
    .B1(_10709_),
    .B2(_13888_),
    .A2(_10530_),
    .A1(net5578));
 sg13g2_a221oi_1 _44715_ (.B2(_13888_),
    .C1(_10519_),
    .B1(_10709_),
    .A1(net5578),
    .Y(_13935_),
    .A2(_10530_));
 sg13g2_o21ai_1 _44716_ (.B1(net5745),
    .Y(_13936_),
    .A1(_10520_),
    .A2(_13934_));
 sg13g2_o21ai_1 _44717_ (.B1(_13933_),
    .Y(_13937_),
    .A1(_13935_),
    .A2(_13936_));
 sg13g2_xnor2_1 _44718_ (.Y(_13938_),
    .A(net5441),
    .B(_13937_));
 sg13g2_nand2_1 _44719_ (.Y(_13939_),
    .A(_13907_),
    .B(_13925_));
 sg13g2_xnor2_1 _44720_ (.Y(_13940_),
    .A(_13938_),
    .B(_13939_));
 sg13g2_o21ai_1 _44721_ (.B1(net5945),
    .Y(_13941_),
    .A1(net5491),
    .A2(_13937_));
 sg13g2_a21oi_1 _44722_ (.A1(net5491),
    .A2(_13940_),
    .Y(_13942_),
    .B1(_13941_));
 sg13g2_a221oi_1 _44723_ (.B2(net5893),
    .C1(_13942_),
    .B1(_13906_),
    .A1(net5978),
    .Y(_13943_),
    .A2(_10524_));
 sg13g2_o21ai_1 _44724_ (.B1(net6872),
    .Y(_13944_),
    .A1(net5262),
    .A2(_10524_));
 sg13g2_a21oi_1 _44725_ (.A1(net5262),
    .A2(_13943_),
    .Y(_13945_),
    .B1(_13944_));
 sg13g2_a21o_1 _44726_ (.A2(net6407),
    .A1(net2925),
    .B1(_13945_),
    .X(_00929_));
 sg13g2_o21ai_1 _44727_ (.B1(_10506_),
    .Y(_13946_),
    .A1(_10517_),
    .A2(_13935_));
 sg13g2_or3_1 _44728_ (.A(_10506_),
    .B(_10517_),
    .C(_13935_),
    .X(_13947_));
 sg13g2_nor2_1 _44729_ (.A(net5744),
    .B(_10505_),
    .Y(_13948_));
 sg13g2_a21oi_1 _44730_ (.A1(_13946_),
    .A2(_13947_),
    .Y(_13949_),
    .B1(net5694));
 sg13g2_nor2_1 _44731_ (.A(_13948_),
    .B(_13949_),
    .Y(_13950_));
 sg13g2_nor2_1 _44732_ (.A(net5491),
    .B(_13950_),
    .Y(_13951_));
 sg13g2_nor3_1 _44733_ (.A(net5441),
    .B(_13948_),
    .C(_13949_),
    .Y(_13952_));
 sg13g2_nand2_1 _44734_ (.Y(_13953_),
    .A(net5385),
    .B(_13950_));
 sg13g2_o21ai_1 _44735_ (.B1(net5441),
    .Y(_13954_),
    .A1(_13948_),
    .A2(_13949_));
 sg13g2_nor2b_1 _44736_ (.A(_13952_),
    .B_N(_13954_),
    .Y(_13955_));
 sg13g2_inv_1 _44737_ (.Y(_13956_),
    .A(_13955_));
 sg13g2_o21ai_1 _44738_ (.B1(net5386),
    .Y(_13957_),
    .A1(_13906_),
    .A2(_13937_));
 sg13g2_nand2_1 _44739_ (.Y(_13958_),
    .A(_13925_),
    .B(_13957_));
 sg13g2_o21ai_1 _44740_ (.B1(_13958_),
    .Y(_13959_),
    .A1(net5385),
    .A2(_13937_));
 sg13g2_xnor2_1 _44741_ (.Y(_13960_),
    .A(_13956_),
    .B(_13959_));
 sg13g2_a21oi_1 _44742_ (.A1(net5491),
    .A2(_13960_),
    .Y(_13961_),
    .B1(_13951_));
 sg13g2_a22oi_1 _44743_ (.Y(_13962_),
    .B1(_13961_),
    .B2(net5224),
    .A2(_13937_),
    .A1(net5204));
 sg13g2_a22oi_1 _44744_ (.Y(_13963_),
    .B1(net5097),
    .B2(_10529_),
    .A2(net6407),
    .A1(net3547));
 sg13g2_o21ai_1 _44745_ (.B1(_13963_),
    .Y(_00930_),
    .A1(net6843),
    .A2(_13962_));
 sg13g2_nand2_1 _44746_ (.Y(_13964_),
    .A(net2447),
    .B(net6407));
 sg13g2_a21o_1 _44747_ (.A2(net5475),
    .A1(net5476),
    .B1(_10533_),
    .X(_13965_));
 sg13g2_a21oi_1 _44748_ (.A1(_10711_),
    .A2(_13965_),
    .Y(_13966_),
    .B1(_10500_));
 sg13g2_nand3_1 _44749_ (.B(_10711_),
    .C(_13965_),
    .A(_10500_),
    .Y(_13967_));
 sg13g2_nand2b_1 _44750_ (.Y(_13968_),
    .B(_13967_),
    .A_N(_13966_));
 sg13g2_nor2_1 _44751_ (.A(net5745),
    .B(_10499_),
    .Y(_13969_));
 sg13g2_a21o_2 _44752_ (.A2(_13968_),
    .A1(net5745),
    .B1(_13969_),
    .X(_13970_));
 sg13g2_nor2_1 _44753_ (.A(net5441),
    .B(_13970_),
    .Y(_13971_));
 sg13g2_xnor2_1 _44754_ (.Y(_13972_),
    .A(net5385),
    .B(_13970_));
 sg13g2_o21ai_1 _44755_ (.B1(_13953_),
    .Y(_13973_),
    .A1(_13956_),
    .A2(_13959_));
 sg13g2_xor2_1 _44756_ (.B(_13973_),
    .A(_13972_),
    .X(_13974_));
 sg13g2_a21oi_1 _44757_ (.A1(net5555),
    .A2(_13970_),
    .Y(_13975_),
    .B1(net5922));
 sg13g2_o21ai_1 _44758_ (.B1(_13975_),
    .Y(_13976_),
    .A1(net5555),
    .A2(_13974_));
 sg13g2_a22oi_1 _44759_ (.Y(_13977_),
    .B1(_13950_),
    .B2(net5895),
    .A2(_10516_),
    .A1(net5979));
 sg13g2_and3_1 _44760_ (.X(_13978_),
    .A(net5261),
    .B(_13976_),
    .C(_13977_));
 sg13g2_o21ai_1 _44761_ (.B1(net6872),
    .Y(_13979_),
    .A1(net5262),
    .A2(_10516_));
 sg13g2_o21ai_1 _44762_ (.B1(_13964_),
    .Y(_00931_),
    .A1(_13978_),
    .A2(_13979_));
 sg13g2_a21oi_1 _44763_ (.A1(net5626),
    .A2(_10499_),
    .Y(_13980_),
    .B1(_13966_));
 sg13g2_xnor2_1 _44764_ (.Y(_13981_),
    .A(_10496_),
    .B(_13980_));
 sg13g2_nand2_1 _44765_ (.Y(_13982_),
    .A(net5695),
    .B(_10494_));
 sg13g2_o21ai_1 _44766_ (.B1(_13982_),
    .Y(_13983_),
    .A1(net5695),
    .A2(_13981_));
 sg13g2_nor2_1 _44767_ (.A(net5491),
    .B(_13983_),
    .Y(_13984_));
 sg13g2_nand2_1 _44768_ (.Y(_13985_),
    .A(net5385),
    .B(_13983_));
 sg13g2_xnor2_1 _44769_ (.Y(_13986_),
    .A(net5441),
    .B(_13983_));
 sg13g2_xnor2_1 _44770_ (.Y(_13987_),
    .A(net5385),
    .B(_13983_));
 sg13g2_nand3b_1 _44771_ (.B(_13954_),
    .C(_13972_),
    .Y(_13988_),
    .A_N(_13952_));
 sg13g2_nor2_1 _44772_ (.A(_13952_),
    .B(_13971_),
    .Y(_13989_));
 sg13g2_o21ai_1 _44773_ (.B1(_13989_),
    .Y(_13990_),
    .A1(_13957_),
    .A2(_13988_));
 sg13g2_nand4_1 _44774_ (.B(_13938_),
    .C(_13955_),
    .A(_13908_),
    .Y(_13991_),
    .D(_13972_));
 sg13g2_a21oi_1 _44775_ (.A1(_13919_),
    .A2(_13923_),
    .Y(_13992_),
    .B1(_13991_));
 sg13g2_o21ai_1 _44776_ (.B1(_13986_),
    .Y(_13993_),
    .A1(_13990_),
    .A2(_13992_));
 sg13g2_or3_1 _44777_ (.A(_13986_),
    .B(_13990_),
    .C(_13992_),
    .X(_13994_));
 sg13g2_a21oi_1 _44778_ (.A1(_13993_),
    .A2(_13994_),
    .Y(_13995_),
    .B1(net5555));
 sg13g2_nor2_1 _44779_ (.A(_13984_),
    .B(_13995_),
    .Y(_13996_));
 sg13g2_a22oi_1 _44780_ (.Y(_13997_),
    .B1(_13996_),
    .B2(net5224),
    .A2(_10505_),
    .A1(net5158));
 sg13g2_o21ai_1 _44781_ (.B1(_13997_),
    .Y(_13998_),
    .A1(net5122),
    .A2(_13970_));
 sg13g2_a22oi_1 _44782_ (.Y(_13999_),
    .B1(net6873),
    .B2(_13998_),
    .A2(net6408),
    .A1(net3389));
 sg13g2_inv_1 _44783_ (.Y(_00932_),
    .A(_13999_));
 sg13g2_nor2_1 _44784_ (.A(net5745),
    .B(_10479_),
    .Y(_14000_));
 sg13g2_o21ai_1 _44785_ (.B1(_10495_),
    .Y(_14001_),
    .A1(_10714_),
    .A2(_13966_));
 sg13g2_xnor2_1 _44786_ (.Y(_14002_),
    .A(_10482_),
    .B(_14001_));
 sg13g2_a21oi_2 _44787_ (.B1(_14000_),
    .Y(_14003_),
    .A2(_14002_),
    .A1(net5744));
 sg13g2_nor2_1 _44788_ (.A(net5384),
    .B(_14003_),
    .Y(_14004_));
 sg13g2_xnor2_1 _44789_ (.Y(_14005_),
    .A(net5384),
    .B(_14003_));
 sg13g2_nand2_1 _44790_ (.Y(_14006_),
    .A(_13985_),
    .B(_13993_));
 sg13g2_xor2_1 _44791_ (.B(_14006_),
    .A(_14005_),
    .X(_14007_));
 sg13g2_o21ai_1 _44792_ (.B1(net5944),
    .Y(_14008_),
    .A1(net5490),
    .A2(_14003_));
 sg13g2_a21oi_1 _44793_ (.A1(net5491),
    .A2(_14007_),
    .Y(_14009_),
    .B1(_14008_));
 sg13g2_a221oi_1 _44794_ (.B2(net5895),
    .C1(_14009_),
    .B1(_13983_),
    .A1(net5979),
    .Y(_14010_),
    .A2(_10499_));
 sg13g2_o21ai_1 _44795_ (.B1(net6873),
    .Y(_14011_),
    .A1(net5255),
    .A2(_10499_));
 sg13g2_a21oi_1 _44796_ (.A1(net5255),
    .A2(_14010_),
    .Y(_14012_),
    .B1(_14011_));
 sg13g2_a21o_1 _44797_ (.A2(net6408),
    .A1(net3549),
    .B1(_14012_),
    .X(_00933_));
 sg13g2_nand2_1 _44798_ (.Y(_14013_),
    .A(net3438),
    .B(net6404));
 sg13g2_nand2_1 _44799_ (.Y(_14014_),
    .A(net5693),
    .B(_10488_));
 sg13g2_o21ai_1 _44800_ (.B1(_10481_),
    .Y(_14015_),
    .A1(_10482_),
    .A2(_14001_));
 sg13g2_xnor2_1 _44801_ (.Y(_14016_),
    .A(_10491_),
    .B(_14015_));
 sg13g2_o21ai_1 _44802_ (.B1(_14014_),
    .Y(_14017_),
    .A1(net5693),
    .A2(_14016_));
 sg13g2_inv_1 _44803_ (.Y(_14018_),
    .A(_14017_));
 sg13g2_nand2_1 _44804_ (.Y(_14019_),
    .A(net5555),
    .B(_14017_));
 sg13g2_nor2_1 _44805_ (.A(net5440),
    .B(_14017_),
    .Y(_14020_));
 sg13g2_xnor2_1 _44806_ (.Y(_14021_),
    .A(net5385),
    .B(_14017_));
 sg13g2_xnor2_1 _44807_ (.Y(_14022_),
    .A(net5440),
    .B(_14017_));
 sg13g2_o21ai_1 _44808_ (.B1(net5384),
    .Y(_14023_),
    .A1(_13983_),
    .A2(_14003_));
 sg13g2_a21oi_1 _44809_ (.A1(_13993_),
    .A2(_14023_),
    .Y(_14024_),
    .B1(_14004_));
 sg13g2_xnor2_1 _44810_ (.Y(_14025_),
    .A(_14022_),
    .B(_14024_));
 sg13g2_o21ai_1 _44811_ (.B1(_14019_),
    .Y(_14026_),
    .A1(net5555),
    .A2(_14025_));
 sg13g2_nor2_1 _44812_ (.A(net5152),
    .B(_14026_),
    .Y(_14027_));
 sg13g2_a221oi_1 _44813_ (.B2(net5204),
    .C1(_14027_),
    .B1(_14003_),
    .A1(net5158),
    .Y(_14028_),
    .A2(_10494_));
 sg13g2_o21ai_1 _44814_ (.B1(_14013_),
    .Y(_00934_),
    .A1(net6843),
    .A2(_14028_));
 sg13g2_a21oi_1 _44815_ (.A1(net5476),
    .A2(net5475),
    .Y(_14029_),
    .B1(_10534_));
 sg13g2_a21o_1 _44816_ (.A2(net5475),
    .A1(net5476),
    .B1(_10534_),
    .X(_14030_));
 sg13g2_o21ai_1 _44817_ (.B1(_10561_),
    .Y(_14031_),
    .A1(_10717_),
    .A2(_14029_));
 sg13g2_nor3_1 _44818_ (.A(_10561_),
    .B(_10717_),
    .C(_14029_),
    .Y(_14032_));
 sg13g2_nor2_1 _44819_ (.A(net5693),
    .B(_14032_),
    .Y(_14033_));
 sg13g2_a22oi_1 _44820_ (.Y(_14034_),
    .B1(_14031_),
    .B2(_14033_),
    .A2(_10558_),
    .A1(net5694));
 sg13g2_xnor2_1 _44821_ (.Y(_14035_),
    .A(net5385),
    .B(_14034_));
 sg13g2_inv_1 _44822_ (.Y(_14036_),
    .A(_14035_));
 sg13g2_a21o_1 _44823_ (.A2(_14024_),
    .A1(_14021_),
    .B1(_14020_),
    .X(_14037_));
 sg13g2_xnor2_1 _44824_ (.Y(_14038_),
    .A(_14036_),
    .B(_14037_));
 sg13g2_a21oi_1 _44825_ (.A1(net5555),
    .A2(_14034_),
    .Y(_14039_),
    .B1(net5922));
 sg13g2_o21ai_1 _44826_ (.B1(_14039_),
    .Y(_14040_),
    .A1(net5555),
    .A2(_14038_));
 sg13g2_a22oi_1 _44827_ (.Y(_14041_),
    .B1(_14018_),
    .B2(net5893),
    .A2(_10479_),
    .A1(net5978));
 sg13g2_and3_1 _44828_ (.X(_14042_),
    .A(net5254),
    .B(_14040_),
    .C(_14041_));
 sg13g2_o21ai_1 _44829_ (.B1(net6873),
    .Y(_14043_),
    .A1(net5255),
    .A2(_10479_));
 sg13g2_nand2_1 _44830_ (.Y(_14044_),
    .A(net2561),
    .B(net6404));
 sg13g2_o21ai_1 _44831_ (.B1(_14044_),
    .Y(_00935_),
    .A1(_14042_),
    .A2(_14043_));
 sg13g2_nand2_1 _44832_ (.Y(_14045_),
    .A(_10559_),
    .B(_14031_));
 sg13g2_xnor2_1 _44833_ (.Y(_14046_),
    .A(_10554_),
    .B(_14045_));
 sg13g2_nand2_1 _44834_ (.Y(_14047_),
    .A(net5745),
    .B(_14046_));
 sg13g2_o21ai_1 _44835_ (.B1(_14047_),
    .Y(_14048_),
    .A1(net5744),
    .A2(_10553_));
 sg13g2_xnor2_1 _44836_ (.Y(_14049_),
    .A(net5386),
    .B(_14048_));
 sg13g2_nor2_1 _44837_ (.A(_13987_),
    .B(_14005_),
    .Y(_14050_));
 sg13g2_nand3_1 _44838_ (.B(_14035_),
    .C(_14050_),
    .A(_14021_),
    .Y(_14051_));
 sg13g2_and4_1 _44839_ (.A(_13990_),
    .B(_14021_),
    .C(_14035_),
    .D(_14050_),
    .X(_14052_));
 sg13g2_nor3_1 _44840_ (.A(_14022_),
    .B(_14023_),
    .C(_14036_),
    .Y(_14053_));
 sg13g2_nor3_1 _44841_ (.A(_14020_),
    .B(_14052_),
    .C(_14053_),
    .Y(_14054_));
 sg13g2_o21ai_1 _44842_ (.B1(_14054_),
    .Y(_14055_),
    .A1(net5441),
    .A2(_14034_));
 sg13g2_nor2_1 _44843_ (.A(_13991_),
    .B(_14051_),
    .Y(_14056_));
 sg13g2_a21oi_2 _44844_ (.B1(_14055_),
    .Y(_14057_),
    .A2(_14056_),
    .A1(_13924_));
 sg13g2_nor2_1 _44845_ (.A(_14049_),
    .B(_14057_),
    .Y(_14058_));
 sg13g2_xnor2_1 _44846_ (.Y(_14059_),
    .A(_14049_),
    .B(_14057_));
 sg13g2_nor2_1 _44847_ (.A(net5491),
    .B(_14048_),
    .Y(_14060_));
 sg13g2_a21oi_1 _44848_ (.A1(net5492),
    .A2(_14059_),
    .Y(_14061_),
    .B1(_14060_));
 sg13g2_a22oi_1 _44849_ (.Y(_14062_),
    .B1(_14061_),
    .B2(net5224),
    .A2(_10489_),
    .A1(net5158));
 sg13g2_o21ai_1 _44850_ (.B1(_14062_),
    .Y(_14063_),
    .A1(net5122),
    .A2(_14034_));
 sg13g2_a22oi_1 _44851_ (.Y(_14064_),
    .B1(net6873),
    .B2(_14063_),
    .A2(net6406),
    .A1(net3027));
 sg13g2_inv_1 _44852_ (.Y(_00936_),
    .A(_14064_));
 sg13g2_nor2_1 _44853_ (.A(net5744),
    .B(_10540_),
    .Y(_14065_));
 sg13g2_nand2_1 _44854_ (.Y(_14066_),
    .A(_10724_),
    .B(_14031_));
 sg13g2_o21ai_1 _44855_ (.B1(_14066_),
    .Y(_14067_),
    .A1(net5625),
    .A2(_10552_));
 sg13g2_a221oi_1 _44856_ (.B2(_14031_),
    .C1(_10541_),
    .B1(_10724_),
    .A1(net5577),
    .Y(_14068_),
    .A2(_10553_));
 sg13g2_xnor2_1 _44857_ (.Y(_14069_),
    .A(_10541_),
    .B(_14067_));
 sg13g2_a21oi_2 _44858_ (.B1(_14065_),
    .Y(_14070_),
    .A2(_14069_),
    .A1(net5744));
 sg13g2_nand2b_1 _44859_ (.Y(_14071_),
    .B(net5440),
    .A_N(_14070_));
 sg13g2_xnor2_1 _44860_ (.Y(_14072_),
    .A(net5386),
    .B(_14070_));
 sg13g2_a21oi_1 _44861_ (.A1(net5386),
    .A2(_14048_),
    .Y(_14073_),
    .B1(_14058_));
 sg13g2_xnor2_1 _44862_ (.Y(_14074_),
    .A(_14072_),
    .B(_14073_));
 sg13g2_o21ai_1 _44863_ (.B1(net5944),
    .Y(_14075_),
    .A1(net5489),
    .A2(_14070_));
 sg13g2_a21oi_1 _44864_ (.A1(net5492),
    .A2(_14074_),
    .Y(_14076_),
    .B1(_14075_));
 sg13g2_a221oi_1 _44865_ (.B2(net5893),
    .C1(_14076_),
    .B1(_14048_),
    .A1(net5978),
    .Y(_14077_),
    .A2(_10558_));
 sg13g2_o21ai_1 _44866_ (.B1(net6872),
    .Y(_14078_),
    .A1(net5254),
    .A2(_10558_));
 sg13g2_a21oi_1 _44867_ (.A1(net5254),
    .A2(_14077_),
    .Y(_14079_),
    .B1(_14078_));
 sg13g2_a21o_1 _44868_ (.A2(net6404),
    .A1(net2691),
    .B1(_14079_),
    .X(_00937_));
 sg13g2_nand2_1 _44869_ (.Y(_14080_),
    .A(net5693),
    .B(_10546_));
 sg13g2_a21oi_1 _44870_ (.A1(net5625),
    .A2(_10540_),
    .Y(_14081_),
    .B1(_14068_));
 sg13g2_xnor2_1 _44871_ (.Y(_14082_),
    .A(_10548_),
    .B(_14081_));
 sg13g2_o21ai_1 _44872_ (.B1(_14080_),
    .Y(_14083_),
    .A1(net5694),
    .A2(_14082_));
 sg13g2_nand2_1 _44873_ (.Y(_14084_),
    .A(net5387),
    .B(_14083_));
 sg13g2_xnor2_1 _44874_ (.Y(_14085_),
    .A(net5440),
    .B(_14083_));
 sg13g2_o21ai_1 _44875_ (.B1(net5387),
    .Y(_14086_),
    .A1(_14048_),
    .A2(_14070_));
 sg13g2_o21ai_1 _44876_ (.B1(_14086_),
    .Y(_14087_),
    .A1(_14049_),
    .A2(_14057_));
 sg13g2_nand2_1 _44877_ (.Y(_14088_),
    .A(_14071_),
    .B(_14087_));
 sg13g2_nand3_1 _44878_ (.B(_14085_),
    .C(_14087_),
    .A(_14071_),
    .Y(_14089_));
 sg13g2_xor2_1 _44879_ (.B(_14088_),
    .A(_14085_),
    .X(_14090_));
 sg13g2_o21ai_1 _44880_ (.B1(net5944),
    .Y(_14091_),
    .A1(net5489),
    .A2(_14083_));
 sg13g2_a21oi_1 _44881_ (.A1(net5490),
    .A2(_14090_),
    .Y(_14092_),
    .B1(_14091_));
 sg13g2_a221oi_1 _44882_ (.B2(net5893),
    .C1(_14092_),
    .B1(_14070_),
    .A1(net5978),
    .Y(_14093_),
    .A2(_10552_));
 sg13g2_o21ai_1 _44883_ (.B1(net6872),
    .Y(_14094_),
    .A1(net5254),
    .A2(_10552_));
 sg13g2_a21oi_1 _44884_ (.A1(net5254),
    .A2(_14093_),
    .Y(_14095_),
    .B1(_14094_));
 sg13g2_a21o_1 _44885_ (.A2(net6404),
    .A1(net2772),
    .B1(_14095_),
    .X(_00938_));
 sg13g2_nand2_1 _44886_ (.Y(_14096_),
    .A(net5694),
    .B(_10581_));
 sg13g2_a21oi_1 _44887_ (.A1(_10716_),
    .A2(_14030_),
    .Y(_14097_),
    .B1(_10563_));
 sg13g2_o21ai_1 _44888_ (.B1(_10583_),
    .Y(_14098_),
    .A1(_10726_),
    .A2(_14097_));
 sg13g2_or3_1 _44889_ (.A(_10583_),
    .B(_10726_),
    .C(_14097_),
    .X(_14099_));
 sg13g2_nand3_1 _44890_ (.B(_14098_),
    .C(_14099_),
    .A(net5744),
    .Y(_14100_));
 sg13g2_nand2_2 _44891_ (.Y(_14101_),
    .A(_14096_),
    .B(_14100_));
 sg13g2_xnor2_1 _44892_ (.Y(_14102_),
    .A(net5440),
    .B(_14101_));
 sg13g2_nand2_1 _44893_ (.Y(_14103_),
    .A(_14084_),
    .B(_14089_));
 sg13g2_xnor2_1 _44894_ (.Y(_14104_),
    .A(_14102_),
    .B(_14103_));
 sg13g2_o21ai_1 _44895_ (.B1(net5944),
    .Y(_14105_),
    .A1(net5490),
    .A2(_14101_));
 sg13g2_a21oi_1 _44896_ (.A1(net5490),
    .A2(_14104_),
    .Y(_14106_),
    .B1(_14105_));
 sg13g2_a221oi_1 _44897_ (.B2(net5893),
    .C1(_14106_),
    .B1(_14083_),
    .A1(net5978),
    .Y(_14107_),
    .A2(_10540_));
 sg13g2_and2_1 _44898_ (.A(net5254),
    .B(_14107_),
    .X(_14108_));
 sg13g2_o21ai_1 _44899_ (.B1(net6872),
    .Y(_14109_),
    .A1(net5255),
    .A2(_10540_));
 sg13g2_nand2_1 _44900_ (.Y(_14110_),
    .A(net2693),
    .B(net6404));
 sg13g2_o21ai_1 _44901_ (.B1(_14110_),
    .Y(_00939_),
    .A1(_14108_),
    .A2(_14109_));
 sg13g2_and3_1 _44902_ (.X(_14111_),
    .A(_10582_),
    .B(_10587_),
    .C(_14098_));
 sg13g2_a21oi_1 _44903_ (.A1(_10582_),
    .A2(_14098_),
    .Y(_14112_),
    .B1(_10587_));
 sg13g2_nor3_1 _44904_ (.A(net5693),
    .B(_14111_),
    .C(_14112_),
    .Y(_14113_));
 sg13g2_a21oi_2 _44905_ (.B1(_14113_),
    .Y(_14114_),
    .A2(_10585_),
    .A1(net5693));
 sg13g2_nor2_1 _44906_ (.A(net5489),
    .B(_14114_),
    .Y(_14115_));
 sg13g2_xnor2_1 _44907_ (.Y(_14116_),
    .A(net5440),
    .B(_14114_));
 sg13g2_inv_1 _44908_ (.Y(_14117_),
    .A(_14116_));
 sg13g2_nand2_1 _44909_ (.Y(_14118_),
    .A(_14085_),
    .B(_14102_));
 sg13g2_o21ai_1 _44910_ (.B1(net5387),
    .Y(_14119_),
    .A1(_14083_),
    .A2(_14101_));
 sg13g2_o21ai_1 _44911_ (.B1(_14119_),
    .Y(_14120_),
    .A1(_14086_),
    .A2(_14118_));
 sg13g2_inv_1 _44912_ (.Y(_14121_),
    .A(_14120_));
 sg13g2_nor2_1 _44913_ (.A(_14049_),
    .B(_14072_),
    .Y(_14122_));
 sg13g2_nand3_1 _44914_ (.B(_14102_),
    .C(_14122_),
    .A(_14085_),
    .Y(_14123_));
 sg13g2_o21ai_1 _44915_ (.B1(_14121_),
    .Y(_14124_),
    .A1(_14057_),
    .A2(_14123_));
 sg13g2_and2_1 _44916_ (.A(_14116_),
    .B(_14124_),
    .X(_14125_));
 sg13g2_xnor2_1 _44917_ (.Y(_14126_),
    .A(_14116_),
    .B(_14124_));
 sg13g2_a21oi_1 _44918_ (.A1(net5489),
    .A2(_14126_),
    .Y(_14127_),
    .B1(_14115_));
 sg13g2_a22oi_1 _44919_ (.Y(_14128_),
    .B1(_14127_),
    .B2(net5224),
    .A2(_14101_),
    .A1(net5204));
 sg13g2_a22oi_1 _44920_ (.Y(_14129_),
    .B1(net5099),
    .B2(_10546_),
    .A2(net6406),
    .A1(net3455));
 sg13g2_o21ai_1 _44921_ (.B1(_14129_),
    .Y(_00940_),
    .A1(net6843),
    .A2(_14128_));
 sg13g2_nor2_1 _44922_ (.A(net5744),
    .B(_10575_),
    .Y(_14130_));
 sg13g2_nand2_1 _44923_ (.Y(_14131_),
    .A(_10720_),
    .B(_14098_));
 sg13g2_o21ai_1 _44924_ (.B1(_14131_),
    .Y(_14132_),
    .A1(net5624),
    .A2(_10586_));
 sg13g2_a221oi_1 _44925_ (.B2(_14098_),
    .C1(_10577_),
    .B1(_10720_),
    .A1(net5577),
    .Y(_14133_),
    .A2(_10585_));
 sg13g2_xnor2_1 _44926_ (.Y(_14134_),
    .A(_10577_),
    .B(_14132_));
 sg13g2_a21oi_2 _44927_ (.B1(_14130_),
    .Y(_14135_),
    .A2(_14134_),
    .A1(net5744));
 sg13g2_nand2b_1 _44928_ (.Y(_14136_),
    .B(net5440),
    .A_N(_14135_));
 sg13g2_xnor2_1 _44929_ (.Y(_14137_),
    .A(net5384),
    .B(_14135_));
 sg13g2_a21oi_1 _44930_ (.A1(net5384),
    .A2(_14114_),
    .Y(_14138_),
    .B1(_14125_));
 sg13g2_xnor2_1 _44931_ (.Y(_14139_),
    .A(_14137_),
    .B(_14138_));
 sg13g2_o21ai_1 _44932_ (.B1(net5944),
    .Y(_14140_),
    .A1(net5489),
    .A2(_14135_));
 sg13g2_a21oi_1 _44933_ (.A1(net5489),
    .A2(_14139_),
    .Y(_14141_),
    .B1(_14140_));
 sg13g2_a221oi_1 _44934_ (.B2(net5893),
    .C1(_14141_),
    .B1(_14114_),
    .A1(net5978),
    .Y(_14142_),
    .A2(_10581_));
 sg13g2_and2_1 _44935_ (.A(net5253),
    .B(_14142_),
    .X(_14143_));
 sg13g2_o21ai_1 _44936_ (.B1(net6872),
    .Y(_14144_),
    .A1(net5255),
    .A2(_10581_));
 sg13g2_nand2_1 _44937_ (.Y(_14145_),
    .A(net2456),
    .B(net6404));
 sg13g2_o21ai_1 _44938_ (.B1(_14145_),
    .Y(_00941_),
    .A1(_14143_),
    .A2(_14144_));
 sg13g2_nand2_1 _44939_ (.Y(_14146_),
    .A(net5693),
    .B(_10569_));
 sg13g2_or3_1 _44940_ (.A(_10570_),
    .B(_10576_),
    .C(_14133_),
    .X(_14147_));
 sg13g2_o21ai_1 _44941_ (.B1(_10570_),
    .Y(_14148_),
    .A1(_10576_),
    .A2(_14133_));
 sg13g2_a21o_1 _44942_ (.A2(_14148_),
    .A1(_14147_),
    .B1(net5693),
    .X(_14149_));
 sg13g2_nand2_1 _44943_ (.Y(_14150_),
    .A(_14146_),
    .B(_14149_));
 sg13g2_nor2_1 _44944_ (.A(net5489),
    .B(_14150_),
    .Y(_14151_));
 sg13g2_a21oi_1 _44945_ (.A1(_14146_),
    .A2(_14149_),
    .Y(_14152_),
    .B1(net5438));
 sg13g2_nand2_1 _44946_ (.Y(_14153_),
    .A(net5384),
    .B(_14150_));
 sg13g2_nand3_1 _44947_ (.B(_14146_),
    .C(_14149_),
    .A(net5440),
    .Y(_14154_));
 sg13g2_nand2_1 _44948_ (.Y(_14155_),
    .A(_14153_),
    .B(_14154_));
 sg13g2_o21ai_1 _44949_ (.B1(net5384),
    .Y(_14156_),
    .A1(_14114_),
    .A2(_14135_));
 sg13g2_inv_1 _44950_ (.Y(_14157_),
    .A(_14156_));
 sg13g2_o21ai_1 _44951_ (.B1(_14136_),
    .Y(_14158_),
    .A1(_14125_),
    .A2(_14157_));
 sg13g2_xnor2_1 _44952_ (.Y(_14159_),
    .A(_14155_),
    .B(_14158_));
 sg13g2_a21oi_1 _44953_ (.A1(net5489),
    .A2(_14159_),
    .Y(_14160_),
    .B1(_14151_));
 sg13g2_a22oi_1 _44954_ (.Y(_14161_),
    .B1(_14160_),
    .B2(net5224),
    .A2(_14135_),
    .A1(net5204));
 sg13g2_a22oi_1 _44955_ (.Y(_14162_),
    .B1(net5099),
    .B2(_10586_),
    .A2(net6406),
    .A1(net2824));
 sg13g2_o21ai_1 _44956_ (.B1(_14162_),
    .Y(_00942_),
    .A1(net6843),
    .A2(_14161_));
 sg13g2_a21oi_2 _44957_ (.B1(_10590_),
    .Y(_14163_),
    .A2(_10224_),
    .A1(_08849_));
 sg13g2_a21o_1 _44958_ (.A2(net5475),
    .A1(net5476),
    .B1(_10590_),
    .X(_14164_));
 sg13g2_o21ai_1 _44959_ (.B1(_10699_),
    .Y(_14165_),
    .A1(_10729_),
    .A2(_14163_));
 sg13g2_nor3_1 _44960_ (.A(_10699_),
    .B(_10729_),
    .C(_14163_),
    .Y(_14166_));
 sg13g2_nor2_1 _44961_ (.A(net5690),
    .B(_14166_),
    .Y(_14167_));
 sg13g2_a22oi_1 _44962_ (.Y(_14168_),
    .B1(_14165_),
    .B2(_14167_),
    .A2(_10697_),
    .A1(net5690));
 sg13g2_inv_1 _44963_ (.Y(_14169_),
    .A(_14168_));
 sg13g2_xnor2_1 _44964_ (.Y(_14170_),
    .A(net5381),
    .B(_14168_));
 sg13g2_o21ai_1 _44965_ (.B1(_14153_),
    .Y(_14171_),
    .A1(_14155_),
    .A2(_14158_));
 sg13g2_xor2_1 _44966_ (.B(_14171_),
    .A(_14170_),
    .X(_14172_));
 sg13g2_a21oi_1 _44967_ (.A1(net5551),
    .A2(_14168_),
    .Y(_14173_),
    .B1(net5922));
 sg13g2_o21ai_1 _44968_ (.B1(_14173_),
    .Y(_14174_),
    .A1(net5555),
    .A2(_14172_));
 sg13g2_a22oi_1 _44969_ (.Y(_14175_),
    .B1(_14150_),
    .B2(net5893),
    .A2(_10575_),
    .A1(net5978));
 sg13g2_and3_1 _44970_ (.X(_14176_),
    .A(net5253),
    .B(_14174_),
    .C(_14175_));
 sg13g2_o21ai_1 _44971_ (.B1(net6868),
    .Y(_14177_),
    .A1(net5253),
    .A2(_10575_));
 sg13g2_nand2_1 _44972_ (.Y(_14178_),
    .A(net2922),
    .B(net6404));
 sg13g2_o21ai_1 _44973_ (.B1(_14178_),
    .Y(_00943_),
    .A1(_14176_),
    .A2(_14177_));
 sg13g2_nand2_1 _44974_ (.Y(_14179_),
    .A(_10698_),
    .B(_14165_));
 sg13g2_xor2_1 _44975_ (.B(_14179_),
    .A(_10694_),
    .X(_14180_));
 sg13g2_mux2_1 _44976_ (.A0(_10693_),
    .A1(_14180_),
    .S(net5742),
    .X(_14181_));
 sg13g2_nand2_1 _44977_ (.Y(_14182_),
    .A(net5382),
    .B(_14181_));
 sg13g2_xnor2_1 _44978_ (.Y(_14183_),
    .A(net5438),
    .B(_14181_));
 sg13g2_nand3b_1 _44979_ (.B(_14154_),
    .C(_14170_),
    .Y(_14184_),
    .A_N(_14152_));
 sg13g2_nor3_1 _44980_ (.A(_14117_),
    .B(_14137_),
    .C(_14184_),
    .Y(_14185_));
 sg13g2_nor2b_1 _44981_ (.A(_14123_),
    .B_N(_14185_),
    .Y(_14186_));
 sg13g2_a21oi_1 _44982_ (.A1(net5384),
    .A2(_14169_),
    .Y(_14187_),
    .B1(_14152_));
 sg13g2_o21ai_1 _44983_ (.B1(_14187_),
    .Y(_14188_),
    .A1(_14156_),
    .A2(_14184_));
 sg13g2_a22oi_1 _44984_ (.Y(_14189_),
    .B1(_14186_),
    .B2(_14055_),
    .A2(_14185_),
    .A1(_14120_));
 sg13g2_nand2b_2 _44985_ (.Y(_14190_),
    .B(_14189_),
    .A_N(_14188_));
 sg13g2_and2_1 _44986_ (.A(_14056_),
    .B(_14186_),
    .X(_14191_));
 sg13g2_inv_1 _44987_ (.Y(_14192_),
    .A(_14191_));
 sg13g2_a21oi_2 _44988_ (.B1(_14192_),
    .Y(_14193_),
    .A2(_13923_),
    .A1(_13919_));
 sg13g2_nor2_1 _44989_ (.A(_14190_),
    .B(_14193_),
    .Y(_14194_));
 sg13g2_o21ai_1 _44990_ (.B1(_14183_),
    .Y(_14195_),
    .A1(_14190_),
    .A2(_14193_));
 sg13g2_xor2_1 _44991_ (.B(_14194_),
    .A(_14183_),
    .X(_14196_));
 sg13g2_o21ai_1 _44992_ (.B1(net5944),
    .Y(_14197_),
    .A1(net5487),
    .A2(_14181_));
 sg13g2_a21oi_1 _44993_ (.A1(net5487),
    .A2(_14196_),
    .Y(_14198_),
    .B1(_14197_));
 sg13g2_a221oi_1 _44994_ (.B2(net5893),
    .C1(_14198_),
    .B1(_14169_),
    .A1(net5978),
    .Y(_14199_),
    .A2(_10569_));
 sg13g2_o21ai_1 _44995_ (.B1(net6868),
    .Y(_14200_),
    .A1(net5253),
    .A2(_10569_));
 sg13g2_a21oi_1 _44996_ (.A1(net5253),
    .A2(_14199_),
    .Y(_14201_),
    .B1(_14200_));
 sg13g2_a21o_1 _44997_ (.A2(net6404),
    .A1(net2721),
    .B1(_14201_),
    .X(_00944_));
 sg13g2_nand2_1 _44998_ (.Y(_14202_),
    .A(net5690),
    .B(_10685_));
 sg13g2_a22oi_1 _44999_ (.Y(_14203_),
    .B1(_10742_),
    .B2(_14165_),
    .A2(_10692_),
    .A1(net5575));
 sg13g2_a221oi_1 _45000_ (.B2(_14165_),
    .C1(_10687_),
    .B1(_10742_),
    .A1(net5575),
    .Y(_14204_),
    .A2(_10692_));
 sg13g2_xor2_1 _45001_ (.B(_14203_),
    .A(_10687_),
    .X(_14205_));
 sg13g2_o21ai_1 _45002_ (.B1(_14202_),
    .Y(_14206_),
    .A1(net5691),
    .A2(_14205_));
 sg13g2_nor2_1 _45003_ (.A(net5381),
    .B(_14206_),
    .Y(_14207_));
 sg13g2_xnor2_1 _45004_ (.Y(_14208_),
    .A(net5438),
    .B(_14206_));
 sg13g2_nand2_1 _45005_ (.Y(_14209_),
    .A(_14182_),
    .B(_14195_));
 sg13g2_xnor2_1 _45006_ (.Y(_14210_),
    .A(_14208_),
    .B(_14209_));
 sg13g2_o21ai_1 _45007_ (.B1(net5944),
    .Y(_14211_),
    .A1(net5487),
    .A2(_14206_));
 sg13g2_a21oi_1 _45008_ (.A1(net5487),
    .A2(_14210_),
    .Y(_14212_),
    .B1(_14211_));
 sg13g2_a221oi_1 _45009_ (.B2(net5889),
    .C1(_14212_),
    .B1(_14181_),
    .A1(net5974),
    .Y(_14213_),
    .A2(_10697_));
 sg13g2_o21ai_1 _45010_ (.B1(net6868),
    .Y(_14214_),
    .A1(net5253),
    .A2(_10697_));
 sg13g2_a21oi_1 _45011_ (.A1(net5253),
    .A2(_14213_),
    .Y(_14215_),
    .B1(_14214_));
 sg13g2_a21o_1 _45012_ (.A2(net6405),
    .A1(net3425),
    .B1(_14215_),
    .X(_00945_));
 sg13g2_or3_1 _45013_ (.A(_10680_),
    .B(_10686_),
    .C(_14204_),
    .X(_14216_));
 sg13g2_o21ai_1 _45014_ (.B1(_10680_),
    .Y(_14217_),
    .A1(_10686_),
    .A2(_14204_));
 sg13g2_a21oi_1 _45015_ (.A1(_14216_),
    .A2(_14217_),
    .Y(_14218_),
    .B1(net5691));
 sg13g2_a21oi_2 _45016_ (.B1(_14218_),
    .Y(_14219_),
    .A2(_10679_),
    .A1(net5691));
 sg13g2_inv_1 _45017_ (.Y(_14220_),
    .A(_14219_));
 sg13g2_nor2_2 _45018_ (.A(net5438),
    .B(_14219_),
    .Y(_14221_));
 sg13g2_and2_1 _45019_ (.A(net5438),
    .B(_14219_),
    .X(_14222_));
 sg13g2_nor2_1 _45020_ (.A(_14221_),
    .B(_14222_),
    .Y(_14223_));
 sg13g2_o21ai_1 _45021_ (.B1(net5381),
    .Y(_14224_),
    .A1(_14181_),
    .A2(_14206_));
 sg13g2_a21oi_1 _45022_ (.A1(_14195_),
    .A2(_14224_),
    .Y(_14225_),
    .B1(_14207_));
 sg13g2_xor2_1 _45023_ (.B(_14225_),
    .A(_14223_),
    .X(_14226_));
 sg13g2_a21oi_1 _45024_ (.A1(net5551),
    .A2(_14219_),
    .Y(_14227_),
    .B1(net5922));
 sg13g2_o21ai_1 _45025_ (.B1(_14227_),
    .Y(_14228_),
    .A1(net5551),
    .A2(_14226_));
 sg13g2_a22oi_1 _45026_ (.Y(_14229_),
    .B1(_14206_),
    .B2(net5889),
    .A2(_10693_),
    .A1(net5974));
 sg13g2_nand3_1 _45027_ (.B(_14228_),
    .C(_14229_),
    .A(net5253),
    .Y(_14230_));
 sg13g2_nor2_1 _45028_ (.A(net5254),
    .B(_10693_),
    .Y(_14231_));
 sg13g2_nor2_1 _45029_ (.A(net6838),
    .B(_14231_),
    .Y(_14232_));
 sg13g2_a22oi_1 _45030_ (.Y(_14233_),
    .B1(_14230_),
    .B2(_14232_),
    .A2(net6405),
    .A1(net3271));
 sg13g2_inv_1 _45031_ (.Y(_00946_),
    .A(_14233_));
 sg13g2_nand2_1 _45032_ (.Y(_14234_),
    .A(net2871),
    .B(net6405));
 sg13g2_nand2_1 _45033_ (.Y(_14235_),
    .A(net5690),
    .B(_10673_));
 sg13g2_a21oi_1 _45034_ (.A1(_10728_),
    .A2(_14164_),
    .Y(_14236_),
    .B1(_10701_));
 sg13g2_o21ai_1 _45035_ (.B1(_10675_),
    .Y(_14237_),
    .A1(_10744_),
    .A2(_14236_));
 sg13g2_or3_1 _45036_ (.A(_10675_),
    .B(_10744_),
    .C(_14236_),
    .X(_14238_));
 sg13g2_nand3_1 _45037_ (.B(_14237_),
    .C(_14238_),
    .A(net5742),
    .Y(_14239_));
 sg13g2_nand2_2 _45038_ (.Y(_14240_),
    .A(_14235_),
    .B(_14239_));
 sg13g2_xnor2_1 _45039_ (.Y(_14241_),
    .A(net5381),
    .B(_14240_));
 sg13g2_a21oi_1 _45040_ (.A1(_14223_),
    .A2(_14225_),
    .Y(_14242_),
    .B1(_14221_));
 sg13g2_xnor2_1 _45041_ (.Y(_14243_),
    .A(_14241_),
    .B(_14242_));
 sg13g2_o21ai_1 _45042_ (.B1(net5944),
    .Y(_14244_),
    .A1(net5487),
    .A2(_14240_));
 sg13g2_a21oi_1 _45043_ (.A1(net5487),
    .A2(_14243_),
    .Y(_14245_),
    .B1(_14244_));
 sg13g2_a221oi_1 _45044_ (.B2(net5889),
    .C1(_14245_),
    .B1(_14220_),
    .A1(net5974),
    .Y(_14246_),
    .A2(_10685_));
 sg13g2_and2_1 _45045_ (.A(net5252),
    .B(_14246_),
    .X(_14247_));
 sg13g2_o21ai_1 _45046_ (.B1(net6868),
    .Y(_14248_),
    .A1(net5252),
    .A2(_10685_));
 sg13g2_o21ai_1 _45047_ (.B1(_14234_),
    .Y(_00947_),
    .A1(_14247_),
    .A2(_14248_));
 sg13g2_nand2_1 _45048_ (.Y(_14249_),
    .A(_10674_),
    .B(_14237_));
 sg13g2_xor2_1 _45049_ (.B(_14249_),
    .A(_10670_),
    .X(_14250_));
 sg13g2_nand2_1 _45050_ (.Y(_14251_),
    .A(net5742),
    .B(_14250_));
 sg13g2_o21ai_1 _45051_ (.B1(_14251_),
    .Y(_14252_),
    .A1(net5741),
    .A2(_10668_));
 sg13g2_nor2_1 _45052_ (.A(net5487),
    .B(_14252_),
    .Y(_14253_));
 sg13g2_xnor2_1 _45053_ (.Y(_14254_),
    .A(net5438),
    .B(_14252_));
 sg13g2_nor4_1 _45054_ (.A(_14221_),
    .B(_14222_),
    .C(_14224_),
    .D(_14241_),
    .Y(_14255_));
 sg13g2_a21oi_1 _45055_ (.A1(net5381),
    .A2(_14240_),
    .Y(_14256_),
    .B1(_14221_));
 sg13g2_nor2b_1 _45056_ (.A(_14255_),
    .B_N(_14256_),
    .Y(_14257_));
 sg13g2_nand2_1 _45057_ (.Y(_14258_),
    .A(_14183_),
    .B(_14208_));
 sg13g2_nor4_1 _45058_ (.A(_14221_),
    .B(_14222_),
    .C(_14241_),
    .D(_14258_),
    .Y(_14259_));
 sg13g2_inv_1 _45059_ (.Y(_14260_),
    .A(_14259_));
 sg13g2_o21ai_1 _45060_ (.B1(_14257_),
    .Y(_14261_),
    .A1(_14194_),
    .A2(_14260_));
 sg13g2_and2_1 _45061_ (.A(_14254_),
    .B(_14261_),
    .X(_14262_));
 sg13g2_xnor2_1 _45062_ (.Y(_14263_),
    .A(_14254_),
    .B(_14261_));
 sg13g2_a21oi_1 _45063_ (.A1(net5487),
    .A2(_14263_),
    .Y(_14264_),
    .B1(_14253_));
 sg13g2_a22oi_1 _45064_ (.Y(_14265_),
    .B1(_14264_),
    .B2(net5221),
    .A2(_14240_),
    .A1(net5200));
 sg13g2_a22oi_1 _45065_ (.Y(_14266_),
    .B1(net5099),
    .B2(_10679_),
    .A2(net6405),
    .A1(net2787));
 sg13g2_o21ai_1 _45066_ (.B1(_14266_),
    .Y(_00948_),
    .A1(net6839),
    .A2(_14265_));
 sg13g2_nor2_1 _45067_ (.A(net5741),
    .B(_10658_),
    .Y(_14267_));
 sg13g2_a22oi_1 _45068_ (.Y(_14268_),
    .B1(_10745_),
    .B2(_14237_),
    .A2(_10668_),
    .A1(net5575));
 sg13g2_nor2b_1 _45069_ (.A(_10659_),
    .B_N(_14268_),
    .Y(_14269_));
 sg13g2_xor2_1 _45070_ (.B(_14268_),
    .A(_10659_),
    .X(_14270_));
 sg13g2_a21oi_2 _45071_ (.B1(_14267_),
    .Y(_14271_),
    .A2(_14270_),
    .A1(net5741));
 sg13g2_nand2b_1 _45072_ (.Y(_14272_),
    .B(net5438),
    .A_N(_14271_));
 sg13g2_nand2_1 _45073_ (.Y(_14273_),
    .A(net5379),
    .B(_14271_));
 sg13g2_nand2_1 _45074_ (.Y(_14274_),
    .A(_14272_),
    .B(_14273_));
 sg13g2_a21oi_1 _45075_ (.A1(net5381),
    .A2(_14252_),
    .Y(_14275_),
    .B1(_14262_));
 sg13g2_xnor2_1 _45076_ (.Y(_14276_),
    .A(_14274_),
    .B(_14275_));
 sg13g2_o21ai_1 _45077_ (.B1(net5940),
    .Y(_14277_),
    .A1(net5485),
    .A2(_14271_));
 sg13g2_a21oi_1 _45078_ (.A1(net5488),
    .A2(_14276_),
    .Y(_14278_),
    .B1(_14277_));
 sg13g2_a221oi_1 _45079_ (.B2(net5890),
    .C1(_14278_),
    .B1(_14252_),
    .A1(net5974),
    .Y(_14279_),
    .A2(_10673_));
 sg13g2_and2_1 _45080_ (.A(net5252),
    .B(_14279_),
    .X(_14280_));
 sg13g2_o21ai_1 _45081_ (.B1(net6869),
    .Y(_14281_),
    .A1(net5256),
    .A2(_10673_));
 sg13g2_nand2_1 _45082_ (.Y(_14282_),
    .A(net2283),
    .B(net6405));
 sg13g2_o21ai_1 _45083_ (.B1(_14282_),
    .Y(_00949_),
    .A1(_14280_),
    .A2(_14281_));
 sg13g2_nand2_1 _45084_ (.Y(_14283_),
    .A(net5690),
    .B(_10662_));
 sg13g2_a21oi_1 _45085_ (.A1(net5619),
    .A2(_10658_),
    .Y(_14284_),
    .B1(_14269_));
 sg13g2_xor2_1 _45086_ (.B(_14284_),
    .A(_10663_),
    .X(_14285_));
 sg13g2_o21ai_1 _45087_ (.B1(_14283_),
    .Y(_14286_),
    .A1(net5690),
    .A2(_14285_));
 sg13g2_nor2_1 _45088_ (.A(net5486),
    .B(_14286_),
    .Y(_14287_));
 sg13g2_and2_1 _45089_ (.A(net5380),
    .B(_14286_),
    .X(_14288_));
 sg13g2_nand2_1 _45090_ (.Y(_14289_),
    .A(net5380),
    .B(_14286_));
 sg13g2_xnor2_1 _45091_ (.Y(_14290_),
    .A(net5380),
    .B(_14286_));
 sg13g2_o21ai_1 _45092_ (.B1(net5379),
    .Y(_14291_),
    .A1(_14252_),
    .A2(_14271_));
 sg13g2_inv_1 _45093_ (.Y(_14292_),
    .A(_14291_));
 sg13g2_o21ai_1 _45094_ (.B1(_14272_),
    .Y(_14293_),
    .A1(_14262_),
    .A2(_14292_));
 sg13g2_xnor2_1 _45095_ (.Y(_14294_),
    .A(_14290_),
    .B(_14293_));
 sg13g2_a21oi_1 _45096_ (.A1(net5485),
    .A2(_14294_),
    .Y(_14295_),
    .B1(_14287_));
 sg13g2_a22oi_1 _45097_ (.Y(_14296_),
    .B1(_14295_),
    .B2(net5222),
    .A2(_14271_),
    .A1(net5201));
 sg13g2_nor2_1 _45098_ (.A(net5066),
    .B(_10668_),
    .Y(_14297_));
 sg13g2_a21oi_1 _45099_ (.A1(net3620),
    .A2(net6405),
    .Y(_14298_),
    .B1(_14297_));
 sg13g2_o21ai_1 _45100_ (.B1(_14298_),
    .Y(_00950_),
    .A1(net6839),
    .A2(_14296_));
 sg13g2_a21oi_1 _45101_ (.A1(_10728_),
    .A2(_14164_),
    .Y(_14299_),
    .B1(_10703_));
 sg13g2_o21ai_1 _45102_ (.B1(_10639_),
    .Y(_14300_),
    .A1(_10748_),
    .A2(_14299_));
 sg13g2_nor3_1 _45103_ (.A(_10639_),
    .B(_10748_),
    .C(_14299_),
    .Y(_14301_));
 sg13g2_nand3b_1 _45104_ (.B(net5741),
    .C(_14300_),
    .Y(_14302_),
    .A_N(_14301_));
 sg13g2_o21ai_1 _45105_ (.B1(_14302_),
    .Y(_14303_),
    .A1(net5741),
    .A2(_10638_));
 sg13g2_and2_1 _45106_ (.A(net5380),
    .B(_14303_),
    .X(_14304_));
 sg13g2_xnor2_1 _45107_ (.Y(_14305_),
    .A(net5380),
    .B(_14303_));
 sg13g2_o21ai_1 _45108_ (.B1(_14289_),
    .Y(_14306_),
    .A1(_14290_),
    .A2(_14293_));
 sg13g2_xor2_1 _45109_ (.B(_14306_),
    .A(_14305_),
    .X(_14307_));
 sg13g2_o21ai_1 _45110_ (.B1(net5940),
    .Y(_14308_),
    .A1(net5486),
    .A2(_14303_));
 sg13g2_a21oi_1 _45111_ (.A1(net5486),
    .A2(_14307_),
    .Y(_14309_),
    .B1(_14308_));
 sg13g2_a22oi_1 _45112_ (.Y(_14310_),
    .B1(_14286_),
    .B2(net5890),
    .A2(_10658_),
    .A1(net5975));
 sg13g2_nand2_1 _45113_ (.Y(_14311_),
    .A(net5252),
    .B(_14310_));
 sg13g2_nor2_1 _45114_ (.A(net5252),
    .B(_10658_),
    .Y(_14312_));
 sg13g2_o21ai_1 _45115_ (.B1(net6869),
    .Y(_14313_),
    .A1(_14309_),
    .A2(_14311_));
 sg13g2_nand2_1 _45116_ (.Y(_14314_),
    .A(net2920),
    .B(net6405));
 sg13g2_o21ai_1 _45117_ (.B1(_14314_),
    .Y(_00951_),
    .A1(_14312_),
    .A2(_14313_));
 sg13g2_nand2_1 _45118_ (.Y(_14315_),
    .A(net3581),
    .B(net6405));
 sg13g2_nor2_1 _45119_ (.A(net5741),
    .B(_10642_),
    .Y(_14316_));
 sg13g2_o21ai_1 _45120_ (.B1(_14300_),
    .Y(_14317_),
    .A1(net5574),
    .A2(_10638_));
 sg13g2_xnor2_1 _45121_ (.Y(_14318_),
    .A(_10645_),
    .B(_14317_));
 sg13g2_a21oi_2 _45122_ (.B1(_14316_),
    .Y(_14319_),
    .A2(_14318_),
    .A1(net5741));
 sg13g2_nand2_1 _45123_ (.Y(_14320_),
    .A(net5379),
    .B(_14319_));
 sg13g2_xnor2_1 _45124_ (.Y(_14321_),
    .A(net5379),
    .B(_14319_));
 sg13g2_inv_1 _45125_ (.Y(_14322_),
    .A(_14321_));
 sg13g2_nand3_1 _45126_ (.B(_14272_),
    .C(_14273_),
    .A(_14254_),
    .Y(_14323_));
 sg13g2_nor4_1 _45127_ (.A(_14257_),
    .B(_14290_),
    .C(_14305_),
    .D(_14323_),
    .Y(_14324_));
 sg13g2_nor3_1 _45128_ (.A(_14290_),
    .B(_14291_),
    .C(_14305_),
    .Y(_14325_));
 sg13g2_nor4_2 _45129_ (.A(_14288_),
    .B(_14304_),
    .C(_14324_),
    .Y(_14326_),
    .D(_14325_));
 sg13g2_inv_1 _45130_ (.Y(_14327_),
    .A(_14326_));
 sg13g2_or4_1 _45131_ (.A(_14260_),
    .B(_14290_),
    .C(_14305_),
    .D(_14323_),
    .X(_14328_));
 sg13g2_inv_1 _45132_ (.Y(_14329_),
    .A(_14328_));
 sg13g2_o21ai_1 _45133_ (.B1(_14329_),
    .Y(_14330_),
    .A1(_14190_),
    .A2(_14193_));
 sg13g2_a21oi_1 _45134_ (.A1(_14326_),
    .A2(_14330_),
    .Y(_14331_),
    .B1(_14321_));
 sg13g2_and3_1 _45135_ (.X(_14332_),
    .A(_14321_),
    .B(_14326_),
    .C(_14330_));
 sg13g2_o21ai_1 _45136_ (.B1(net5485),
    .Y(_14333_),
    .A1(_14331_),
    .A2(_14332_));
 sg13g2_o21ai_1 _45137_ (.B1(_14333_),
    .Y(_14334_),
    .A1(net5485),
    .A2(_14319_));
 sg13g2_nor2_1 _45138_ (.A(net5151),
    .B(_14334_),
    .Y(_14335_));
 sg13g2_a221oi_1 _45139_ (.B2(net5201),
    .C1(_14335_),
    .B1(_14303_),
    .A1(net5157),
    .Y(_14336_),
    .A2(_10662_));
 sg13g2_o21ai_1 _45140_ (.B1(_14315_),
    .Y(_00952_),
    .A1(net6839),
    .A2(_14336_));
 sg13g2_nand2_1 _45141_ (.Y(_14337_),
    .A(net5690),
    .B(_10626_));
 sg13g2_a22oi_1 _45142_ (.Y(_14338_),
    .B1(_10731_),
    .B2(_14300_),
    .A2(_10643_),
    .A1(net5574));
 sg13g2_xnor2_1 _45143_ (.Y(_14339_),
    .A(_10629_),
    .B(_14338_));
 sg13g2_o21ai_1 _45144_ (.B1(_14337_),
    .Y(_14340_),
    .A1(net5690),
    .A2(_14339_));
 sg13g2_nor2_1 _45145_ (.A(net5379),
    .B(_14340_),
    .Y(_14341_));
 sg13g2_or2_1 _45146_ (.X(_14342_),
    .B(_14340_),
    .A(net5379));
 sg13g2_nand2_1 _45147_ (.Y(_14343_),
    .A(net5379),
    .B(_14340_));
 sg13g2_nand2_1 _45148_ (.Y(_14344_),
    .A(_14342_),
    .B(_14343_));
 sg13g2_a21oi_1 _45149_ (.A1(net5379),
    .A2(_14319_),
    .Y(_14345_),
    .B1(_14331_));
 sg13g2_xnor2_1 _45150_ (.Y(_14346_),
    .A(_14344_),
    .B(_14345_));
 sg13g2_o21ai_1 _45151_ (.B1(net5940),
    .Y(_14347_),
    .A1(net5485),
    .A2(_14340_));
 sg13g2_a21oi_1 _45152_ (.A1(net5485),
    .A2(_14346_),
    .Y(_14348_),
    .B1(_14347_));
 sg13g2_nor2_1 _45153_ (.A(net6005),
    .B(_10638_),
    .Y(_14349_));
 sg13g2_a21oi_1 _45154_ (.A1(net5889),
    .A2(_14319_),
    .Y(_14350_),
    .B1(_14349_));
 sg13g2_nand2_1 _45155_ (.Y(_14351_),
    .A(net5252),
    .B(_14350_));
 sg13g2_nor2b_1 _45156_ (.A(net5252),
    .B_N(_10638_),
    .Y(_14352_));
 sg13g2_o21ai_1 _45157_ (.B1(net6869),
    .Y(_14353_),
    .A1(_14348_),
    .A2(_14351_));
 sg13g2_nand2_1 _45158_ (.Y(_14354_),
    .A(net2298),
    .B(net6396));
 sg13g2_o21ai_1 _45159_ (.B1(_14354_),
    .Y(_00953_),
    .A1(_14352_),
    .A2(_14353_));
 sg13g2_a21oi_1 _45160_ (.A1(_10629_),
    .A2(_14338_),
    .Y(_14355_),
    .B1(_10627_));
 sg13g2_xnor2_1 _45161_ (.Y(_14356_),
    .A(_10633_),
    .B(_14355_));
 sg13g2_nor2_1 _45162_ (.A(net5738),
    .B(_10632_),
    .Y(_14357_));
 sg13g2_a21oi_2 _45163_ (.B1(_14357_),
    .Y(_14358_),
    .A2(_14356_),
    .A1(net5741));
 sg13g2_nand2_1 _45164_ (.Y(_14359_),
    .A(net5377),
    .B(_14358_));
 sg13g2_inv_1 _45165_ (.Y(_14360_),
    .A(_14359_));
 sg13g2_xnor2_1 _45166_ (.Y(_14361_),
    .A(net5377),
    .B(_14358_));
 sg13g2_nand2_1 _45167_ (.Y(_14362_),
    .A(_14320_),
    .B(_14343_));
 sg13g2_nor2_1 _45168_ (.A(_14331_),
    .B(_14362_),
    .Y(_14363_));
 sg13g2_nor3_1 _45169_ (.A(_14341_),
    .B(_14361_),
    .C(_14363_),
    .Y(_14364_));
 sg13g2_o21ai_1 _45170_ (.B1(_14361_),
    .Y(_14365_),
    .A1(_14341_),
    .A2(_14363_));
 sg13g2_nand2b_1 _45171_ (.Y(_14366_),
    .B(_14365_),
    .A_N(_14364_));
 sg13g2_nor2_1 _45172_ (.A(net5485),
    .B(_14358_),
    .Y(_14367_));
 sg13g2_a21oi_1 _45173_ (.A1(net5485),
    .A2(_14366_),
    .Y(_14368_),
    .B1(_14367_));
 sg13g2_a22oi_1 _45174_ (.Y(_14369_),
    .B1(_14368_),
    .B2(net5222),
    .A2(_14340_),
    .A1(net5201));
 sg13g2_a22oi_1 _45175_ (.Y(_14370_),
    .B1(net5095),
    .B2(_10642_),
    .A2(net6397),
    .A1(net3506));
 sg13g2_o21ai_1 _45176_ (.B1(_14370_),
    .Y(_00954_),
    .A1(net6839),
    .A2(_14369_));
 sg13g2_nand2_1 _45177_ (.Y(_14371_),
    .A(net5688),
    .B(_10613_));
 sg13g2_o21ai_1 _45178_ (.B1(_10646_),
    .Y(_14372_),
    .A1(_10748_),
    .A2(_14299_));
 sg13g2_a21oi_1 _45179_ (.A1(_10734_),
    .A2(_14372_),
    .Y(_14373_),
    .B1(_10614_));
 sg13g2_nand3_1 _45180_ (.B(_10734_),
    .C(_14372_),
    .A(_10614_),
    .Y(_14374_));
 sg13g2_nand2_1 _45181_ (.Y(_14375_),
    .A(net5739),
    .B(_14374_));
 sg13g2_o21ai_1 _45182_ (.B1(_14371_),
    .Y(_14376_),
    .A1(_14373_),
    .A2(_14375_));
 sg13g2_nand2_1 _45183_ (.Y(_14377_),
    .A(net5377),
    .B(_14376_));
 sg13g2_xnor2_1 _45184_ (.Y(_14378_),
    .A(net5378),
    .B(_14376_));
 sg13g2_nor3_1 _45185_ (.A(_14360_),
    .B(_14364_),
    .C(_14378_),
    .Y(_14379_));
 sg13g2_o21ai_1 _45186_ (.B1(_14378_),
    .Y(_14380_),
    .A1(_14360_),
    .A2(_14364_));
 sg13g2_nor2_1 _45187_ (.A(net5549),
    .B(_14379_),
    .Y(_14381_));
 sg13g2_o21ai_1 _45188_ (.B1(net5940),
    .Y(_14382_),
    .A1(net5483),
    .A2(_14376_));
 sg13g2_a21oi_1 _45189_ (.A1(_14380_),
    .A2(_14381_),
    .Y(_14383_),
    .B1(_14382_));
 sg13g2_a22oi_1 _45190_ (.Y(_14384_),
    .B1(_14358_),
    .B2(net5889),
    .A2(_10626_),
    .A1(net5974));
 sg13g2_nand2_1 _45191_ (.Y(_14385_),
    .A(net5251),
    .B(_14384_));
 sg13g2_nor2_1 _45192_ (.A(_14383_),
    .B(_14385_),
    .Y(_14386_));
 sg13g2_o21ai_1 _45193_ (.B1(net6869),
    .Y(_14387_),
    .A1(net5251),
    .A2(_10626_));
 sg13g2_nand2_1 _45194_ (.Y(_14388_),
    .A(net2368),
    .B(net6396));
 sg13g2_o21ai_1 _45195_ (.B1(_14388_),
    .Y(_00955_),
    .A1(_14386_),
    .A2(_14387_));
 sg13g2_nand2_1 _45196_ (.Y(_14389_),
    .A(net5688),
    .B(_10617_));
 sg13g2_a21oi_1 _45197_ (.A1(net5621),
    .A2(_10613_),
    .Y(_14390_),
    .B1(_14373_));
 sg13g2_xor2_1 _45198_ (.B(_14390_),
    .A(_10619_),
    .X(_14391_));
 sg13g2_o21ai_1 _45199_ (.B1(_14389_),
    .Y(_14392_),
    .A1(net5688),
    .A2(_14391_));
 sg13g2_nand2_1 _45200_ (.Y(_14393_),
    .A(net5377),
    .B(_14392_));
 sg13g2_xnor2_1 _45201_ (.Y(_14394_),
    .A(net5436),
    .B(_14392_));
 sg13g2_nor2_1 _45202_ (.A(_14361_),
    .B(_14378_),
    .Y(_14395_));
 sg13g2_nand2_1 _45203_ (.Y(_14396_),
    .A(_14359_),
    .B(_14377_));
 sg13g2_a21o_1 _45204_ (.A2(_14395_),
    .A1(_14362_),
    .B1(_14396_),
    .X(_14397_));
 sg13g2_nand4_1 _45205_ (.B(_14342_),
    .C(_14343_),
    .A(_14322_),
    .Y(_14398_),
    .D(_14395_));
 sg13g2_a21oi_1 _45206_ (.A1(_14326_),
    .A2(_14330_),
    .Y(_14399_),
    .B1(_14398_));
 sg13g2_o21ai_1 _45207_ (.B1(_14394_),
    .Y(_14400_),
    .A1(_14397_),
    .A2(_14399_));
 sg13g2_or3_1 _45208_ (.A(_14394_),
    .B(_14397_),
    .C(_14399_),
    .X(_14401_));
 sg13g2_nand2_1 _45209_ (.Y(_14402_),
    .A(_14400_),
    .B(_14401_));
 sg13g2_o21ai_1 _45210_ (.B1(net5940),
    .Y(_14403_),
    .A1(net5483),
    .A2(_14392_));
 sg13g2_a21oi_1 _45211_ (.A1(net5488),
    .A2(_14402_),
    .Y(_14404_),
    .B1(_14403_));
 sg13g2_a221oi_1 _45212_ (.B2(net5889),
    .C1(_14404_),
    .B1(_14376_),
    .A1(net5974),
    .Y(_14405_),
    .A2(_10632_));
 sg13g2_o21ai_1 _45213_ (.B1(net6867),
    .Y(_14406_),
    .A1(net5251),
    .A2(_10632_));
 sg13g2_a21oi_1 _45214_ (.A1(net5251),
    .A2(_14405_),
    .Y(_14407_),
    .B1(_14406_));
 sg13g2_a21o_1 _45215_ (.A2(net6396),
    .A1(net2122),
    .B1(_14407_),
    .X(_00956_));
 sg13g2_nand2_1 _45216_ (.Y(_14408_),
    .A(_14393_),
    .B(_14400_));
 sg13g2_nor2_1 _45217_ (.A(net5739),
    .B(_10606_),
    .Y(_14409_));
 sg13g2_o21ai_1 _45218_ (.B1(_10618_),
    .Y(_14410_),
    .A1(_10737_),
    .A2(_14373_));
 sg13g2_xnor2_1 _45219_ (.Y(_14411_),
    .A(_10609_),
    .B(_14410_));
 sg13g2_a21oi_2 _45220_ (.B1(_14409_),
    .Y(_14412_),
    .A2(_14411_),
    .A1(net5739));
 sg13g2_nand2b_1 _45221_ (.Y(_14413_),
    .B(net5436),
    .A_N(_14412_));
 sg13g2_inv_1 _45222_ (.Y(_14414_),
    .A(_14413_));
 sg13g2_xnor2_1 _45223_ (.Y(_14415_),
    .A(net5436),
    .B(_14412_));
 sg13g2_xnor2_1 _45224_ (.Y(_14416_),
    .A(_14408_),
    .B(_14415_));
 sg13g2_o21ai_1 _45225_ (.B1(net5940),
    .Y(_14417_),
    .A1(net5483),
    .A2(_14412_));
 sg13g2_a21oi_1 _45226_ (.A1(net5483),
    .A2(_14416_),
    .Y(_14418_),
    .B1(_14417_));
 sg13g2_a22oi_1 _45227_ (.Y(_14419_),
    .B1(_14392_),
    .B2(net5889),
    .A2(_10613_),
    .A1(net5974));
 sg13g2_nand2_1 _45228_ (.Y(_14420_),
    .A(net5251),
    .B(_14419_));
 sg13g2_nor2_1 _45229_ (.A(net5251),
    .B(_10613_),
    .Y(_14421_));
 sg13g2_o21ai_1 _45230_ (.B1(net6867),
    .Y(_14422_),
    .A1(_14418_),
    .A2(_14420_));
 sg13g2_nand2_1 _45231_ (.Y(_14423_),
    .A(net1987),
    .B(net6396));
 sg13g2_o21ai_1 _45232_ (.B1(_14423_),
    .Y(_00957_),
    .A1(_14421_),
    .A2(_14422_));
 sg13g2_nand2_1 _45233_ (.Y(_14424_),
    .A(net5688),
    .B(_10593_));
 sg13g2_o21ai_1 _45234_ (.B1(_10607_),
    .Y(_14425_),
    .A1(_10609_),
    .A2(_14410_));
 sg13g2_xnor2_1 _45235_ (.Y(_14426_),
    .A(_10595_),
    .B(_14425_));
 sg13g2_o21ai_1 _45236_ (.B1(_14424_),
    .Y(_14427_),
    .A1(net5688),
    .A2(_14426_));
 sg13g2_nand2_1 _45237_ (.Y(_14428_),
    .A(net5377),
    .B(_14427_));
 sg13g2_inv_1 _45238_ (.Y(_14429_),
    .A(_14428_));
 sg13g2_xnor2_1 _45239_ (.Y(_14430_),
    .A(net5436),
    .B(_14427_));
 sg13g2_o21ai_1 _45240_ (.B1(net5377),
    .Y(_14431_),
    .A1(_14392_),
    .A2(_14412_));
 sg13g2_a21oi_1 _45241_ (.A1(_14400_),
    .A2(_14431_),
    .Y(_14432_),
    .B1(_14414_));
 sg13g2_xnor2_1 _45242_ (.Y(_14433_),
    .A(_14430_),
    .B(_14432_));
 sg13g2_nor2_1 _45243_ (.A(net5483),
    .B(_14427_),
    .Y(_14434_));
 sg13g2_a21oi_1 _45244_ (.A1(net5483),
    .A2(_14433_),
    .Y(_14435_),
    .B1(_14434_));
 sg13g2_a22oi_1 _45245_ (.Y(_14436_),
    .B1(_14435_),
    .B2(net5221),
    .A2(_14412_),
    .A1(net5201));
 sg13g2_a22oi_1 _45246_ (.Y(_14437_),
    .B1(net5095),
    .B2(_10617_),
    .A2(net6396),
    .A1(net2417));
 sg13g2_o21ai_1 _45247_ (.B1(_14437_),
    .Y(_00958_),
    .A1(net6839),
    .A2(_14436_));
 sg13g2_nand2_1 _45248_ (.Y(_14438_),
    .A(net2033),
    .B(net6396));
 sg13g2_nand2_1 _45249_ (.Y(_14439_),
    .A(net5688),
    .B(_10463_));
 sg13g2_a21oi_2 _45250_ (.B1(_10706_),
    .Y(_14440_),
    .A2(net5475),
    .A1(net5476));
 sg13g2_nor2_1 _45251_ (.A(_10750_),
    .B(_14440_),
    .Y(_14441_));
 sg13g2_o21ai_1 _45252_ (.B1(_10465_),
    .Y(_14442_),
    .A1(_10750_),
    .A2(_14440_));
 sg13g2_xor2_1 _45253_ (.B(_14441_),
    .A(_10465_),
    .X(_14443_));
 sg13g2_o21ai_1 _45254_ (.B1(_14439_),
    .Y(_14444_),
    .A1(net5689),
    .A2(_14443_));
 sg13g2_xnor2_1 _45255_ (.Y(_14445_),
    .A(net5436),
    .B(_14444_));
 sg13g2_a21oi_1 _45256_ (.A1(_14430_),
    .A2(_14432_),
    .Y(_14446_),
    .B1(_14429_));
 sg13g2_xor2_1 _45257_ (.B(_14446_),
    .A(_14445_),
    .X(_14447_));
 sg13g2_o21ai_1 _45258_ (.B1(net5940),
    .Y(_14448_),
    .A1(net5483),
    .A2(_14444_));
 sg13g2_a21oi_1 _45259_ (.A1(net5483),
    .A2(_14447_),
    .Y(_14449_),
    .B1(_14448_));
 sg13g2_a22oi_1 _45260_ (.Y(_14450_),
    .B1(_14427_),
    .B2(net5889),
    .A2(_10606_),
    .A1(net5974));
 sg13g2_nand2_1 _45261_ (.Y(_14451_),
    .A(net5251),
    .B(_14450_));
 sg13g2_nor2_1 _45262_ (.A(_14449_),
    .B(_14451_),
    .Y(_14452_));
 sg13g2_o21ai_1 _45263_ (.B1(net6867),
    .Y(_14453_),
    .A1(net5251),
    .A2(_10606_));
 sg13g2_o21ai_1 _45264_ (.B1(_14438_),
    .Y(_00959_),
    .A1(_14452_),
    .A2(_14453_));
 sg13g2_nand2_1 _45265_ (.Y(_14454_),
    .A(net5686),
    .B(_10457_));
 sg13g2_nor2b_1 _45266_ (.A(_10464_),
    .B_N(_14442_),
    .Y(_14455_));
 sg13g2_xor2_1 _45267_ (.B(_14455_),
    .A(_10459_),
    .X(_14456_));
 sg13g2_o21ai_1 _45268_ (.B1(_14454_),
    .Y(_14457_),
    .A1(net5687),
    .A2(_14456_));
 sg13g2_nand2_1 _45269_ (.Y(_14458_),
    .A(net5375),
    .B(_14457_));
 sg13g2_xnor2_1 _45270_ (.Y(_14459_),
    .A(net5434),
    .B(_14457_));
 sg13g2_nand4_1 _45271_ (.B(_14415_),
    .C(_14430_),
    .A(_14394_),
    .Y(_14460_),
    .D(_14445_));
 sg13g2_nor2_1 _45272_ (.A(_14398_),
    .B(_14460_),
    .Y(_14461_));
 sg13g2_nor3_2 _45273_ (.A(_14328_),
    .B(_14398_),
    .C(_14460_),
    .Y(_14462_));
 sg13g2_and2_1 _45274_ (.A(_14191_),
    .B(_14462_),
    .X(_14463_));
 sg13g2_o21ai_1 _45275_ (.B1(_14463_),
    .Y(_14464_),
    .A1(_13922_),
    .A2(_13920_));
 sg13g2_nand2b_1 _45276_ (.Y(_14465_),
    .B(_14397_),
    .A_N(_14460_));
 sg13g2_nand3b_1 _45277_ (.B(_14445_),
    .C(_14430_),
    .Y(_14466_),
    .A_N(_14431_));
 sg13g2_o21ai_1 _45278_ (.B1(net5377),
    .Y(_14467_),
    .A1(_14427_),
    .A2(_14444_));
 sg13g2_nand3_1 _45279_ (.B(_14466_),
    .C(_14467_),
    .A(_14465_),
    .Y(_14468_));
 sg13g2_a221oi_1 _45280_ (.B2(_14190_),
    .C1(_14468_),
    .B1(_14462_),
    .A1(_14327_),
    .Y(_14469_),
    .A2(_14461_));
 sg13g2_and2_1 _45281_ (.A(net1121),
    .B(_14469_),
    .X(_14470_));
 sg13g2_nor2b_1 _45282_ (.A(_14470_),
    .B_N(_14459_),
    .Y(_14471_));
 sg13g2_xor2_1 _45283_ (.B(_14470_),
    .A(_14459_),
    .X(_14472_));
 sg13g2_nand2_1 _45284_ (.Y(_14473_),
    .A(net5481),
    .B(_14472_));
 sg13g2_o21ai_1 _45285_ (.B1(_14473_),
    .Y(_14474_),
    .A1(net5481),
    .A2(_14457_));
 sg13g2_a22oi_1 _45286_ (.Y(_14475_),
    .B1(_14444_),
    .B2(net5200),
    .A2(_10593_),
    .A1(net5157));
 sg13g2_o21ai_1 _45287_ (.B1(_14475_),
    .Y(_14476_),
    .A1(net5151),
    .A2(_14474_));
 sg13g2_nand2_1 _45288_ (.Y(_14477_),
    .A(net6868),
    .B(_14476_));
 sg13g2_o21ai_1 _45289_ (.B1(_14477_),
    .Y(_00960_),
    .A1(_18108_),
    .A2(net6483));
 sg13g2_nand2_1 _45290_ (.Y(_14478_),
    .A(net5687),
    .B(_10450_));
 sg13g2_a22oi_1 _45291_ (.Y(_14479_),
    .B1(_10751_),
    .B2(_14442_),
    .A2(_10458_),
    .A1(net5571));
 sg13g2_xnor2_1 _45292_ (.Y(_14480_),
    .A(_10452_),
    .B(_14479_));
 sg13g2_o21ai_1 _45293_ (.B1(_14478_),
    .Y(_14481_),
    .A1(net5687),
    .A2(_14480_));
 sg13g2_or2_1 _45294_ (.X(_14482_),
    .B(_14481_),
    .A(net5376));
 sg13g2_nand2_1 _45295_ (.Y(_14483_),
    .A(net5376),
    .B(_14481_));
 sg13g2_and2_1 _45296_ (.A(_14482_),
    .B(_14483_),
    .X(_14484_));
 sg13g2_a21oi_1 _45297_ (.A1(net5375),
    .A2(_14457_),
    .Y(_14485_),
    .B1(_14471_));
 sg13g2_xor2_1 _45298_ (.B(_14485_),
    .A(_14484_),
    .X(_14486_));
 sg13g2_o21ai_1 _45299_ (.B1(net5939),
    .Y(_14487_),
    .A1(net5481),
    .A2(_14481_));
 sg13g2_a21oi_1 _45300_ (.A1(net5481),
    .A2(_14486_),
    .Y(_14488_),
    .B1(_14487_));
 sg13g2_a221oi_1 _45301_ (.B2(net5887),
    .C1(_14488_),
    .B1(_14457_),
    .A1(net5972),
    .Y(_14489_),
    .A2(_10463_));
 sg13g2_o21ai_1 _45302_ (.B1(net6867),
    .Y(_14490_),
    .A1(net5249),
    .A2(_10463_));
 sg13g2_a21oi_2 _45303_ (.B1(_14490_),
    .Y(_14491_),
    .A2(_14489_),
    .A1(net5249));
 sg13g2_a21o_1 _45304_ (.A2(net6387),
    .A1(net2989),
    .B1(_14491_),
    .X(_00961_));
 sg13g2_nand2_1 _45305_ (.Y(_14492_),
    .A(net2533),
    .B(net6387));
 sg13g2_a21oi_1 _45306_ (.A1(_10452_),
    .A2(_14479_),
    .Y(_14493_),
    .B1(_10451_));
 sg13g2_xnor2_1 _45307_ (.Y(_14494_),
    .A(_10445_),
    .B(_14493_));
 sg13g2_mux2_1 _45308_ (.A0(_10444_),
    .A1(_14494_),
    .S(net5738),
    .X(_14495_));
 sg13g2_nor2_1 _45309_ (.A(net5482),
    .B(_14495_),
    .Y(_14496_));
 sg13g2_nand2_1 _45310_ (.Y(_14497_),
    .A(net5376),
    .B(_14495_));
 sg13g2_xnor2_1 _45311_ (.Y(_14498_),
    .A(net5434),
    .B(_14495_));
 sg13g2_inv_1 _45312_ (.Y(_14499_),
    .A(_14498_));
 sg13g2_nand2_1 _45313_ (.Y(_14500_),
    .A(_14458_),
    .B(_14483_));
 sg13g2_o21ai_1 _45314_ (.B1(_14482_),
    .Y(_14501_),
    .A1(_14471_),
    .A2(_14500_));
 sg13g2_xnor2_1 _45315_ (.Y(_14502_),
    .A(_14498_),
    .B(_14501_));
 sg13g2_nor2_1 _45316_ (.A(net5548),
    .B(_14502_),
    .Y(_14503_));
 sg13g2_nor3_1 _45317_ (.A(net5151),
    .B(_14496_),
    .C(_14503_),
    .Y(_14504_));
 sg13g2_a221oi_1 _45318_ (.B2(net5200),
    .C1(_14504_),
    .B1(_14481_),
    .A1(net5157),
    .Y(_14505_),
    .A2(_10457_));
 sg13g2_o21ai_1 _45319_ (.B1(_14492_),
    .Y(_00962_),
    .A1(net6836),
    .A2(_14505_));
 sg13g2_or2_1 _45320_ (.X(_14506_),
    .B(_14441_),
    .A(_10466_));
 sg13g2_a21oi_1 _45321_ (.A1(_10754_),
    .A2(_14506_),
    .Y(_14507_),
    .B1(_10432_));
 sg13g2_nand3_1 _45322_ (.B(_10754_),
    .C(_14506_),
    .A(_10432_),
    .Y(_14508_));
 sg13g2_nand2_1 _45323_ (.Y(_14509_),
    .A(net5738),
    .B(_14508_));
 sg13g2_nor2_1 _45324_ (.A(_14507_),
    .B(_14509_),
    .Y(_14510_));
 sg13g2_a21oi_2 _45325_ (.B1(_14510_),
    .Y(_14511_),
    .A2(_10429_),
    .A1(net5686));
 sg13g2_xnor2_1 _45326_ (.Y(_14512_),
    .A(net5375),
    .B(_14511_));
 sg13g2_o21ai_1 _45327_ (.B1(_14497_),
    .Y(_14513_),
    .A1(_14499_),
    .A2(_14501_));
 sg13g2_xor2_1 _45328_ (.B(_14513_),
    .A(_14512_),
    .X(_14514_));
 sg13g2_a21oi_1 _45329_ (.A1(net5548),
    .A2(_14511_),
    .Y(_14515_),
    .B1(net5920));
 sg13g2_o21ai_1 _45330_ (.B1(_14515_),
    .Y(_14516_),
    .A1(net5548),
    .A2(_14514_));
 sg13g2_a22oi_1 _45331_ (.Y(_14517_),
    .B1(_14495_),
    .B2(net5888),
    .A2(_10450_),
    .A1(net5973));
 sg13g2_and3_1 _45332_ (.X(_14518_),
    .A(net5249),
    .B(_14516_),
    .C(_14517_));
 sg13g2_o21ai_1 _45333_ (.B1(net6866),
    .Y(_14519_),
    .A1(net5248),
    .A2(_10450_));
 sg13g2_nand2_1 _45334_ (.Y(_14520_),
    .A(net2591),
    .B(net6394));
 sg13g2_o21ai_1 _45335_ (.B1(_14520_),
    .Y(_00963_),
    .A1(_14518_),
    .A2(_14519_));
 sg13g2_nor2_1 _45336_ (.A(_10430_),
    .B(_14507_),
    .Y(_14521_));
 sg13g2_xor2_1 _45337_ (.B(_14521_),
    .A(_10439_),
    .X(_14522_));
 sg13g2_nand2_1 _45338_ (.Y(_14523_),
    .A(net5686),
    .B(_10436_));
 sg13g2_o21ai_1 _45339_ (.B1(_14523_),
    .Y(_14524_),
    .A1(net5686),
    .A2(_14522_));
 sg13g2_nand2_1 _45340_ (.Y(_14525_),
    .A(net5375),
    .B(_14524_));
 sg13g2_xnor2_1 _45341_ (.Y(_14526_),
    .A(net5434),
    .B(_14524_));
 sg13g2_nand3_1 _45342_ (.B(_14500_),
    .C(_14512_),
    .A(_14498_),
    .Y(_14527_));
 sg13g2_o21ai_1 _45343_ (.B1(_14497_),
    .Y(_14528_),
    .A1(net5435),
    .A2(_14511_));
 sg13g2_nor2b_1 _45344_ (.A(_14528_),
    .B_N(_14527_),
    .Y(_14529_));
 sg13g2_nand4_1 _45345_ (.B(_14484_),
    .C(_14498_),
    .A(_14459_),
    .Y(_14530_),
    .D(_14512_));
 sg13g2_o21ai_1 _45346_ (.B1(_14529_),
    .Y(_14531_),
    .A1(_14470_),
    .A2(_14530_));
 sg13g2_nand2_2 _45347_ (.Y(_14532_),
    .A(_14526_),
    .B(_14531_));
 sg13g2_xnor2_1 _45348_ (.Y(_14533_),
    .A(_14526_),
    .B(_14531_));
 sg13g2_nor2_1 _45349_ (.A(net5481),
    .B(_14524_),
    .Y(_14534_));
 sg13g2_a21oi_1 _45350_ (.A1(net5481),
    .A2(_14533_),
    .Y(_14535_),
    .B1(_14534_));
 sg13g2_a22oi_1 _45351_ (.Y(_14536_),
    .B1(_14535_),
    .B2(net5221),
    .A2(_10444_),
    .A1(net5157));
 sg13g2_o21ai_1 _45352_ (.B1(_14536_),
    .Y(_14537_),
    .A1(net5122),
    .A2(_14511_));
 sg13g2_a22oi_1 _45353_ (.Y(_14538_),
    .B1(net6866),
    .B2(_14537_),
    .A2(net6394),
    .A1(net3376));
 sg13g2_inv_1 _45354_ (.Y(_00964_),
    .A(_14538_));
 sg13g2_nand2_1 _45355_ (.Y(_14539_),
    .A(net5686),
    .B(_10419_));
 sg13g2_o21ai_1 _45356_ (.B1(_10438_),
    .Y(_14540_),
    .A1(_10756_),
    .A2(_14507_));
 sg13g2_nor2_1 _45357_ (.A(_10421_),
    .B(_14540_),
    .Y(_14541_));
 sg13g2_a21o_1 _45358_ (.A2(_14540_),
    .A1(_10421_),
    .B1(net5686),
    .X(_14542_));
 sg13g2_o21ai_1 _45359_ (.B1(_14539_),
    .Y(_14543_),
    .A1(_14541_),
    .A2(_14542_));
 sg13g2_inv_1 _45360_ (.Y(_14544_),
    .A(_14543_));
 sg13g2_xnor2_1 _45361_ (.Y(_14545_),
    .A(net5435),
    .B(_14543_));
 sg13g2_nand3_1 _45362_ (.B(_14532_),
    .C(_14545_),
    .A(_14525_),
    .Y(_14546_));
 sg13g2_a21oi_1 _45363_ (.A1(_14525_),
    .A2(_14532_),
    .Y(_14547_),
    .B1(_14545_));
 sg13g2_nor2_1 _45364_ (.A(net5549),
    .B(_14547_),
    .Y(_14548_));
 sg13g2_a221oi_1 _45365_ (.B2(_14548_),
    .C1(net5920),
    .B1(_14546_),
    .A1(net5549),
    .Y(_14549_),
    .A2(_14544_));
 sg13g2_a221oi_1 _45366_ (.B2(net5887),
    .C1(_14549_),
    .B1(_14524_),
    .A1(net5972),
    .Y(_14550_),
    .A2(_10429_));
 sg13g2_and2_1 _45367_ (.A(net5248),
    .B(_14550_),
    .X(_14551_));
 sg13g2_o21ai_1 _45368_ (.B1(net6866),
    .Y(_14552_),
    .A1(net5247),
    .A2(_10429_));
 sg13g2_nand2_1 _45369_ (.Y(_14553_),
    .A(net3231),
    .B(net6394));
 sg13g2_o21ai_1 _45370_ (.B1(_14553_),
    .Y(_00965_),
    .A1(_14551_),
    .A2(_14552_));
 sg13g2_nand2_1 _45371_ (.Y(_14554_),
    .A(net5686),
    .B(_10424_));
 sg13g2_nor2_1 _45372_ (.A(_10420_),
    .B(_14541_),
    .Y(_14555_));
 sg13g2_xnor2_1 _45373_ (.Y(_14556_),
    .A(_10425_),
    .B(_14555_));
 sg13g2_o21ai_1 _45374_ (.B1(_14554_),
    .Y(_14557_),
    .A1(net5686),
    .A2(_14556_));
 sg13g2_nor2_1 _45375_ (.A(net5481),
    .B(_14557_),
    .Y(_14558_));
 sg13g2_xnor2_1 _45376_ (.Y(_14559_),
    .A(net5435),
    .B(_14557_));
 sg13g2_inv_1 _45377_ (.Y(_14560_),
    .A(_14559_));
 sg13g2_o21ai_1 _45378_ (.B1(_14525_),
    .Y(_14561_),
    .A1(net5435),
    .A2(_14544_));
 sg13g2_inv_1 _45379_ (.Y(_14562_),
    .A(_14561_));
 sg13g2_nand2_1 _45380_ (.Y(_14563_),
    .A(_14532_),
    .B(_14562_));
 sg13g2_o21ai_1 _45381_ (.B1(_14563_),
    .Y(_14564_),
    .A1(net5375),
    .A2(_14543_));
 sg13g2_a221oi_1 _45382_ (.B2(_14532_),
    .C1(_14560_),
    .B1(_14562_),
    .A1(net5435),
    .Y(_14565_),
    .A2(_14544_));
 sg13g2_xnor2_1 _45383_ (.Y(_14566_),
    .A(_14560_),
    .B(_14564_));
 sg13g2_a21oi_1 _45384_ (.A1(net5481),
    .A2(_14566_),
    .Y(_14567_),
    .B1(_14558_));
 sg13g2_a22oi_1 _45385_ (.Y(_14568_),
    .B1(_14567_),
    .B2(net5221),
    .A2(_14543_),
    .A1(net5200));
 sg13g2_a22oi_1 _45386_ (.Y(_14569_),
    .B1(net5096),
    .B2(_10436_),
    .A2(net6394),
    .A1(net3445));
 sg13g2_o21ai_1 _45387_ (.B1(_14569_),
    .Y(_00966_),
    .A1(net6838),
    .A2(_14568_));
 sg13g2_nand2_1 _45388_ (.Y(_14570_),
    .A(net2786),
    .B(net6394));
 sg13g2_nor2_1 _45389_ (.A(_10468_),
    .B(_14441_),
    .Y(_14571_));
 sg13g2_o21ai_1 _45390_ (.B1(_10467_),
    .Y(_14572_),
    .A1(_10750_),
    .A2(_14440_));
 sg13g2_o21ai_1 _45391_ (.B1(_10407_),
    .Y(_14573_),
    .A1(_10759_),
    .A2(_14571_));
 sg13g2_nor3_1 _45392_ (.A(_10407_),
    .B(_10759_),
    .C(_14571_),
    .Y(_14574_));
 sg13g2_nor2_1 _45393_ (.A(net5687),
    .B(_14574_),
    .Y(_14575_));
 sg13g2_a22oi_1 _45394_ (.Y(_14576_),
    .B1(_14573_),
    .B2(_14575_),
    .A2(_10405_),
    .A1(net5687));
 sg13g2_inv_1 _45395_ (.Y(_14577_),
    .A(_14576_));
 sg13g2_xnor2_1 _45396_ (.Y(_14578_),
    .A(net5375),
    .B(_14576_));
 sg13g2_a21oi_1 _45397_ (.A1(net5375),
    .A2(_14557_),
    .Y(_14579_),
    .B1(_14565_));
 sg13g2_xnor2_1 _45398_ (.Y(_14580_),
    .A(_14578_),
    .B(_14579_));
 sg13g2_a21oi_1 _45399_ (.A1(net5549),
    .A2(_14576_),
    .Y(_14581_),
    .B1(net5921));
 sg13g2_o21ai_1 _45400_ (.B1(_14581_),
    .Y(_14582_),
    .A1(net5548),
    .A2(_14580_));
 sg13g2_a22oi_1 _45401_ (.Y(_14583_),
    .B1(_14557_),
    .B2(net5887),
    .A2(_10419_),
    .A1(net5972));
 sg13g2_and3_1 _45402_ (.X(_14584_),
    .A(net5248),
    .B(_14582_),
    .C(_14583_));
 sg13g2_o21ai_1 _45403_ (.B1(net6868),
    .Y(_14585_),
    .A1(net5248),
    .A2(_10419_));
 sg13g2_o21ai_1 _45404_ (.B1(_14570_),
    .Y(_00967_),
    .A1(_14584_),
    .A2(_14585_));
 sg13g2_and3_1 _45405_ (.X(_14586_),
    .A(_10401_),
    .B(_10406_),
    .C(_14573_));
 sg13g2_a21oi_1 _45406_ (.A1(_10406_),
    .A2(_14573_),
    .Y(_14587_),
    .B1(_10401_));
 sg13g2_o21ai_1 _45407_ (.B1(net5738),
    .Y(_14588_),
    .A1(_14586_),
    .A2(_14587_));
 sg13g2_o21ai_1 _45408_ (.B1(_14588_),
    .Y(_14589_),
    .A1(net5738),
    .A2(_10399_));
 sg13g2_nand2_1 _45409_ (.Y(_14590_),
    .A(net5376),
    .B(_14589_));
 sg13g2_xnor2_1 _45410_ (.Y(_14591_),
    .A(net5434),
    .B(_14589_));
 sg13g2_nand2_1 _45411_ (.Y(_14592_),
    .A(_14559_),
    .B(_14578_));
 sg13g2_nand2_1 _45412_ (.Y(_14593_),
    .A(_14526_),
    .B(_14545_));
 sg13g2_nor2_1 _45413_ (.A(_14529_),
    .B(_14593_),
    .Y(_14594_));
 sg13g2_nor2_1 _45414_ (.A(_14561_),
    .B(_14594_),
    .Y(_14595_));
 sg13g2_o21ai_1 _45415_ (.B1(net5375),
    .Y(_14596_),
    .A1(_14557_),
    .A2(_14577_));
 sg13g2_o21ai_1 _45416_ (.B1(_14596_),
    .Y(_14597_),
    .A1(_14592_),
    .A2(_14595_));
 sg13g2_nor3_1 _45417_ (.A(_14530_),
    .B(_14592_),
    .C(_14593_),
    .Y(_14598_));
 sg13g2_inv_1 _45418_ (.Y(_14599_),
    .A(_14598_));
 sg13g2_a21oi_1 _45419_ (.A1(net1121),
    .A2(_14469_),
    .Y(_14600_),
    .B1(_14599_));
 sg13g2_or2_1 _45420_ (.X(_14601_),
    .B(_14600_),
    .A(_14597_));
 sg13g2_and2_1 _45421_ (.A(_14591_),
    .B(_14601_),
    .X(_14602_));
 sg13g2_nand2_1 _45422_ (.Y(_14603_),
    .A(_14591_),
    .B(_14601_));
 sg13g2_xnor2_1 _45423_ (.Y(_14604_),
    .A(_14591_),
    .B(_14601_));
 sg13g2_o21ai_1 _45424_ (.B1(net5939),
    .Y(_14605_),
    .A1(net5482),
    .A2(_14589_));
 sg13g2_a21oi_1 _45425_ (.A1(net5482),
    .A2(_14604_),
    .Y(_14606_),
    .B1(_14605_));
 sg13g2_a221oi_1 _45426_ (.B2(net5887),
    .C1(_14606_),
    .B1(_14577_),
    .A1(net5972),
    .Y(_14607_),
    .A2(_10424_));
 sg13g2_o21ai_1 _45427_ (.B1(net6866),
    .Y(_14608_),
    .A1(net5247),
    .A2(_10424_));
 sg13g2_a21oi_1 _45428_ (.A1(net5248),
    .A2(_14607_),
    .Y(_14609_),
    .B1(_14608_));
 sg13g2_a21o_1 _45429_ (.A2(net6394),
    .A1(net3149),
    .B1(_14609_),
    .X(_00968_));
 sg13g2_nor2_1 _45430_ (.A(net5738),
    .B(_10389_),
    .Y(_14610_));
 sg13g2_a22oi_1 _45431_ (.Y(_14611_),
    .B1(_10761_),
    .B2(_14573_),
    .A2(_10399_),
    .A1(net5571));
 sg13g2_xnor2_1 _45432_ (.Y(_14612_),
    .A(_10391_),
    .B(_14611_));
 sg13g2_a21oi_1 _45433_ (.A1(net5738),
    .A2(_14612_),
    .Y(_14613_),
    .B1(_14610_));
 sg13g2_inv_1 _45434_ (.Y(_14614_),
    .A(_14613_));
 sg13g2_nand2_1 _45435_ (.Y(_14615_),
    .A(net5434),
    .B(_14614_));
 sg13g2_nand2_1 _45436_ (.Y(_14616_),
    .A(net5376),
    .B(_14613_));
 sg13g2_and2_1 _45437_ (.A(_14615_),
    .B(_14616_),
    .X(_14617_));
 sg13g2_nand3_1 _45438_ (.B(_14603_),
    .C(_14617_),
    .A(_14590_),
    .Y(_14618_));
 sg13g2_a21oi_1 _45439_ (.A1(_14590_),
    .A2(_14603_),
    .Y(_14619_),
    .B1(_14617_));
 sg13g2_nor2_1 _45440_ (.A(net5548),
    .B(_14619_),
    .Y(_14620_));
 sg13g2_a221oi_1 _45441_ (.B2(_14620_),
    .C1(net5921),
    .B1(_14618_),
    .A1(net5548),
    .Y(_14621_),
    .A2(_14614_));
 sg13g2_a221oi_1 _45442_ (.B2(net5887),
    .C1(_14621_),
    .B1(_14589_),
    .A1(net5972),
    .Y(_14622_),
    .A2(_10405_));
 sg13g2_and2_1 _45443_ (.A(net5247),
    .B(_14622_),
    .X(_14623_));
 sg13g2_o21ai_1 _45444_ (.B1(net6866),
    .Y(_14624_),
    .A1(net5247),
    .A2(_10405_));
 sg13g2_nand2_1 _45445_ (.Y(_14625_),
    .A(net3273),
    .B(net6394));
 sg13g2_o21ai_1 _45446_ (.B1(_14625_),
    .Y(_00969_),
    .A1(_14623_),
    .A2(_14624_));
 sg13g2_or2_1 _45447_ (.X(_14626_),
    .B(_10394_),
    .A(net5738));
 sg13g2_a21oi_1 _45448_ (.A1(_10391_),
    .A2(_14611_),
    .Y(_14627_),
    .B1(_10390_));
 sg13g2_xnor2_1 _45449_ (.Y(_14628_),
    .A(_10395_),
    .B(_14627_));
 sg13g2_o21ai_1 _45450_ (.B1(_14626_),
    .Y(_14629_),
    .A1(net5687),
    .A2(_14628_));
 sg13g2_nor2_1 _45451_ (.A(net5434),
    .B(_14629_),
    .Y(_14630_));
 sg13g2_xnor2_1 _45452_ (.Y(_14631_),
    .A(net5434),
    .B(_14629_));
 sg13g2_nand2_1 _45453_ (.Y(_14632_),
    .A(_14590_),
    .B(_14616_));
 sg13g2_inv_1 _45454_ (.Y(_14633_),
    .A(_14632_));
 sg13g2_o21ai_1 _45455_ (.B1(_14615_),
    .Y(_14634_),
    .A1(_14602_),
    .A2(_14632_));
 sg13g2_a221oi_1 _45456_ (.B2(_14603_),
    .C1(_14631_),
    .B1(_14633_),
    .A1(net5434),
    .Y(_14635_),
    .A2(_14614_));
 sg13g2_xor2_1 _45457_ (.B(_14634_),
    .A(_14631_),
    .X(_14636_));
 sg13g2_a21oi_1 _45458_ (.A1(net5548),
    .A2(_14629_),
    .Y(_14637_),
    .B1(net5921));
 sg13g2_o21ai_1 _45459_ (.B1(_14637_),
    .Y(_14638_),
    .A1(net5548),
    .A2(_14636_));
 sg13g2_a22oi_1 _45460_ (.Y(_14639_),
    .B1(_14613_),
    .B2(net5887),
    .A2(_10400_),
    .A1(net5972));
 sg13g2_nand3_1 _45461_ (.B(_14638_),
    .C(_14639_),
    .A(net5247),
    .Y(_14640_));
 sg13g2_nor2_1 _45462_ (.A(net5247),
    .B(_10400_),
    .Y(_14641_));
 sg13g2_nor2_1 _45463_ (.A(net6838),
    .B(_14641_),
    .Y(_14642_));
 sg13g2_a22oi_1 _45464_ (.Y(_14643_),
    .B1(_14640_),
    .B2(_14642_),
    .A2(net6395),
    .A1(net3161));
 sg13g2_inv_1 _45465_ (.Y(_00970_),
    .A(_14643_));
 sg13g2_nand2_1 _45466_ (.Y(_14644_),
    .A(net5685),
    .B(_10374_));
 sg13g2_a21oi_1 _45467_ (.A1(_10758_),
    .A2(_14572_),
    .Y(_14645_),
    .B1(_10408_));
 sg13g2_o21ai_1 _45468_ (.B1(_10377_),
    .Y(_14646_),
    .A1(_10763_),
    .A2(_14645_));
 sg13g2_or3_1 _45469_ (.A(_10377_),
    .B(_10763_),
    .C(_14645_),
    .X(_14647_));
 sg13g2_nand3_1 _45470_ (.B(_14646_),
    .C(_14647_),
    .A(net5740),
    .Y(_14648_));
 sg13g2_nand2_2 _45471_ (.Y(_14649_),
    .A(_14644_),
    .B(_14648_));
 sg13g2_nand2_1 _45472_ (.Y(_14650_),
    .A(net5374),
    .B(_14649_));
 sg13g2_xnor2_1 _45473_ (.Y(_14651_),
    .A(net5374),
    .B(_14649_));
 sg13g2_nor2_1 _45474_ (.A(_14630_),
    .B(_14635_),
    .Y(_14652_));
 sg13g2_xnor2_1 _45475_ (.Y(_14653_),
    .A(_14651_),
    .B(_14652_));
 sg13g2_o21ai_1 _45476_ (.B1(net5939),
    .Y(_14654_),
    .A1(net5484),
    .A2(_14649_));
 sg13g2_a21oi_1 _45477_ (.A1(net5484),
    .A2(_14653_),
    .Y(_14655_),
    .B1(_14654_));
 sg13g2_nor2_1 _45478_ (.A(net5880),
    .B(_14629_),
    .Y(_14656_));
 sg13g2_a21oi_1 _45479_ (.A1(net5972),
    .A2(_10389_),
    .Y(_14657_),
    .B1(_14656_));
 sg13g2_nand2_1 _45480_ (.Y(_14658_),
    .A(net5247),
    .B(_14657_));
 sg13g2_nor2_1 _45481_ (.A(net5247),
    .B(_10389_),
    .Y(_14659_));
 sg13g2_o21ai_1 _45482_ (.B1(net6868),
    .Y(_14660_),
    .A1(_14655_),
    .A2(_14658_));
 sg13g2_nand2_1 _45483_ (.Y(_14661_),
    .A(net2620),
    .B(net6394));
 sg13g2_o21ai_1 _45484_ (.B1(_14661_),
    .Y(_00971_),
    .A1(_14659_),
    .A2(_14660_));
 sg13g2_nand2_1 _45485_ (.Y(_14662_),
    .A(_10375_),
    .B(_14646_));
 sg13g2_xnor2_1 _45486_ (.Y(_14663_),
    .A(_10382_),
    .B(_14662_));
 sg13g2_nand2_1 _45487_ (.Y(_14664_),
    .A(net5685),
    .B(_10380_));
 sg13g2_o21ai_1 _45488_ (.B1(_14664_),
    .Y(_14665_),
    .A1(net5685),
    .A2(_14663_));
 sg13g2_nor2_1 _45489_ (.A(net5484),
    .B(_14665_),
    .Y(_14666_));
 sg13g2_nand2_1 _45490_ (.Y(_14667_),
    .A(net5374),
    .B(_14665_));
 sg13g2_xnor2_1 _45491_ (.Y(_14668_),
    .A(net5378),
    .B(_14665_));
 sg13g2_nor2_1 _45492_ (.A(_14631_),
    .B(_14651_),
    .Y(_14669_));
 sg13g2_a21o_1 _45493_ (.A2(_14669_),
    .A1(_14632_),
    .B1(_14630_),
    .X(_14670_));
 sg13g2_nor2b_1 _45494_ (.A(_14670_),
    .B_N(_14650_),
    .Y(_14671_));
 sg13g2_nand2b_1 _45495_ (.Y(_14672_),
    .B(_14650_),
    .A_N(_14670_));
 sg13g2_and3_1 _45496_ (.X(_14673_),
    .A(_14591_),
    .B(_14617_),
    .C(_14669_));
 sg13g2_o21ai_1 _45497_ (.B1(_14673_),
    .Y(_14674_),
    .A1(_14597_),
    .A2(_14600_));
 sg13g2_a21o_2 _45498_ (.A2(_14674_),
    .A1(_14671_),
    .B1(_14668_),
    .X(_14675_));
 sg13g2_nand3_1 _45499_ (.B(_14671_),
    .C(_14674_),
    .A(_14668_),
    .Y(_14676_));
 sg13g2_a21oi_1 _45500_ (.A1(_14675_),
    .A2(_14676_),
    .Y(_14677_),
    .B1(net5550));
 sg13g2_nor2_1 _45501_ (.A(_14666_),
    .B(_14677_),
    .Y(_14678_));
 sg13g2_a22oi_1 _45502_ (.Y(_14679_),
    .B1(_14678_),
    .B2(net5221),
    .A2(_14649_),
    .A1(net5200));
 sg13g2_a22oi_1 _45503_ (.Y(_14680_),
    .B1(net5096),
    .B2(_10394_),
    .A2(net6396),
    .A1(net3593));
 sg13g2_o21ai_1 _45504_ (.B1(_14680_),
    .Y(_00972_),
    .A1(net6838),
    .A2(_14679_));
 sg13g2_nand2_1 _45505_ (.Y(_14681_),
    .A(net5685),
    .B(_10364_));
 sg13g2_a21oi_1 _45506_ (.A1(_10765_),
    .A2(_14646_),
    .Y(_14682_),
    .B1(_10381_));
 sg13g2_xnor2_1 _45507_ (.Y(_14683_),
    .A(_10366_),
    .B(_14682_));
 sg13g2_o21ai_1 _45508_ (.B1(_14681_),
    .Y(_14684_),
    .A1(net5685),
    .A2(_14683_));
 sg13g2_inv_1 _45509_ (.Y(_14685_),
    .A(_14684_));
 sg13g2_xnor2_1 _45510_ (.Y(_14686_),
    .A(net5374),
    .B(_14684_));
 sg13g2_nand2_1 _45511_ (.Y(_14687_),
    .A(_14667_),
    .B(_14675_));
 sg13g2_xor2_1 _45512_ (.B(_14687_),
    .A(_14686_),
    .X(_14688_));
 sg13g2_o21ai_1 _45513_ (.B1(net5939),
    .Y(_14689_),
    .A1(net5484),
    .A2(_14684_));
 sg13g2_a21oi_1 _45514_ (.A1(net5484),
    .A2(_14688_),
    .Y(_14690_),
    .B1(_14689_));
 sg13g2_a22oi_1 _45515_ (.Y(_14691_),
    .B1(_14665_),
    .B2(net5887),
    .A2(_10374_),
    .A1(net5975));
 sg13g2_nand2_1 _45516_ (.Y(_14692_),
    .A(net5246),
    .B(_14691_));
 sg13g2_nor2_1 _45517_ (.A(net5246),
    .B(_10374_),
    .Y(_14693_));
 sg13g2_o21ai_1 _45518_ (.B1(net6867),
    .Y(_14694_),
    .A1(_14690_),
    .A2(_14692_));
 sg13g2_nand2_1 _45519_ (.Y(_14695_),
    .A(net2376),
    .B(net6396));
 sg13g2_o21ai_1 _45520_ (.B1(_14695_),
    .Y(_00973_),
    .A1(_14693_),
    .A2(_14694_));
 sg13g2_nand2_1 _45521_ (.Y(_14696_),
    .A(net5200),
    .B(_14684_));
 sg13g2_nand2_1 _45522_ (.Y(_14697_),
    .A(net5685),
    .B(_10369_));
 sg13g2_a21oi_1 _45523_ (.A1(_10366_),
    .A2(_14682_),
    .Y(_14698_),
    .B1(_10365_));
 sg13g2_xor2_1 _45524_ (.B(_14698_),
    .A(_10370_),
    .X(_14699_));
 sg13g2_o21ai_1 _45525_ (.B1(_14697_),
    .Y(_14700_),
    .A1(net5689),
    .A2(_14699_));
 sg13g2_xnor2_1 _45526_ (.Y(_14701_),
    .A(net5437),
    .B(_14700_));
 sg13g2_inv_1 _45527_ (.Y(_14702_),
    .A(_14701_));
 sg13g2_o21ai_1 _45528_ (.B1(net5374),
    .Y(_14703_),
    .A1(_14665_),
    .A2(_14684_));
 sg13g2_a22oi_1 _45529_ (.Y(_14704_),
    .B1(_14703_),
    .B2(_14675_),
    .A2(_14685_),
    .A1(net5437));
 sg13g2_a221oi_1 _45530_ (.B2(_14675_),
    .C1(_14702_),
    .B1(_14703_),
    .A1(net5437),
    .Y(_14705_),
    .A2(_14685_));
 sg13g2_xnor2_1 _45531_ (.Y(_14706_),
    .A(_14702_),
    .B(_14704_));
 sg13g2_nor2_1 _45532_ (.A(net5484),
    .B(_14700_),
    .Y(_14707_));
 sg13g2_o21ai_1 _45533_ (.B1(net5221),
    .Y(_14708_),
    .A1(net5550),
    .A2(_14706_));
 sg13g2_o21ai_1 _45534_ (.B1(_14696_),
    .Y(_14709_),
    .A1(_14707_),
    .A2(_14708_));
 sg13g2_a22oi_1 _45535_ (.Y(_14710_),
    .B1(_14709_),
    .B2(net6867),
    .A2(_10380_),
    .A1(net5096));
 sg13g2_o21ai_1 _45536_ (.B1(_14710_),
    .Y(_00974_),
    .A1(_18106_),
    .A2(net6483));
 sg13g2_o21ai_1 _45537_ (.B1(_10469_),
    .Y(_14711_),
    .A1(_10750_),
    .A2(_14440_));
 sg13g2_nand2b_2 _45538_ (.Y(_14712_),
    .B(_14711_),
    .A_N(_10768_));
 sg13g2_nand2_1 _45539_ (.Y(_14713_),
    .A(_10327_),
    .B(_14712_));
 sg13g2_o21ai_1 _45540_ (.B1(net5740),
    .Y(_14714_),
    .A1(_10327_),
    .A2(_14712_));
 sg13g2_nor2b_1 _45541_ (.A(_14714_),
    .B_N(_14713_),
    .Y(_14715_));
 sg13g2_a21oi_1 _45542_ (.A1(net5685),
    .A2(_10325_),
    .Y(_14716_),
    .B1(_14715_));
 sg13g2_inv_1 _45543_ (.Y(_14717_),
    .A(_14716_));
 sg13g2_xnor2_1 _45544_ (.Y(_14718_),
    .A(net5437),
    .B(_14716_));
 sg13g2_inv_1 _45545_ (.Y(_14719_),
    .A(_14718_));
 sg13g2_a21oi_1 _45546_ (.A1(net5374),
    .A2(_14700_),
    .Y(_14720_),
    .B1(_14705_));
 sg13g2_xnor2_1 _45547_ (.Y(_14721_),
    .A(_14719_),
    .B(_14720_));
 sg13g2_a21oi_1 _45548_ (.A1(net5550),
    .A2(_14716_),
    .Y(_14722_),
    .B1(net5921));
 sg13g2_o21ai_1 _45549_ (.B1(_14722_),
    .Y(_14723_),
    .A1(net5550),
    .A2(_14721_));
 sg13g2_a22oi_1 _45550_ (.Y(_14724_),
    .B1(_14700_),
    .B2(net5887),
    .A2(_10364_),
    .A1(net5972));
 sg13g2_and3_1 _45551_ (.X(_14725_),
    .A(net5246),
    .B(_14723_),
    .C(_14724_));
 sg13g2_o21ai_1 _45552_ (.B1(net6871),
    .Y(_14726_),
    .A1(net5246),
    .A2(_10364_));
 sg13g2_nand2_1 _45553_ (.Y(_14727_),
    .A(net2671),
    .B(net6395));
 sg13g2_o21ai_1 _45554_ (.B1(_14727_),
    .Y(_00975_),
    .A1(_14725_),
    .A2(_14726_));
 sg13g2_nand2_1 _45555_ (.Y(_14728_),
    .A(net2235),
    .B(net6395));
 sg13g2_nand2_1 _45556_ (.Y(_14729_),
    .A(net5684),
    .B(_10319_));
 sg13g2_nand2_1 _45557_ (.Y(_14730_),
    .A(_10326_),
    .B(_14713_));
 sg13g2_xnor2_1 _45558_ (.Y(_14731_),
    .A(_10321_),
    .B(_14730_));
 sg13g2_o21ai_1 _45559_ (.B1(_14729_),
    .Y(_14732_),
    .A1(net5685),
    .A2(_14731_));
 sg13g2_and2_1 _45560_ (.A(net5371),
    .B(_14732_),
    .X(_14733_));
 sg13g2_xnor2_1 _45561_ (.Y(_14734_),
    .A(net5432),
    .B(_14732_));
 sg13g2_xnor2_1 _45562_ (.Y(_14735_),
    .A(net5374),
    .B(_14732_));
 sg13g2_nand2_1 _45563_ (.Y(_14736_),
    .A(_14701_),
    .B(_14719_));
 sg13g2_nor3_1 _45564_ (.A(_14668_),
    .B(_14686_),
    .C(_14736_),
    .Y(_14737_));
 sg13g2_and2_1 _45565_ (.A(_14673_),
    .B(_14737_),
    .X(_14738_));
 sg13g2_nand2_1 _45566_ (.Y(_14739_),
    .A(_14598_),
    .B(_14738_));
 sg13g2_a21o_2 _45567_ (.A2(_14469_),
    .A1(net1121),
    .B1(_14739_),
    .X(_14740_));
 sg13g2_o21ai_1 _45568_ (.B1(net5374),
    .Y(_14741_),
    .A1(_14700_),
    .A2(_14717_));
 sg13g2_o21ai_1 _45569_ (.B1(_14741_),
    .Y(_14742_),
    .A1(_14703_),
    .A2(_14736_));
 sg13g2_a221oi_1 _45570_ (.B2(_14597_),
    .C1(_14742_),
    .B1(_14738_),
    .A1(_14672_),
    .Y(_14743_),
    .A2(_14737_));
 sg13g2_a21o_1 _45571_ (.A2(_14743_),
    .A1(_14740_),
    .B1(_14735_),
    .X(_14744_));
 sg13g2_nand3b_1 _45572_ (.B(_14740_),
    .C(_14743_),
    .Y(_14745_),
    .A_N(_14734_));
 sg13g2_and2_1 _45573_ (.A(_14744_),
    .B(_14745_),
    .X(_14746_));
 sg13g2_nor2_1 _45574_ (.A(net5484),
    .B(_14732_),
    .Y(_14747_));
 sg13g2_o21ai_1 _45575_ (.B1(net5939),
    .Y(_14748_),
    .A1(net5550),
    .A2(_14746_));
 sg13g2_a22oi_1 _45576_ (.Y(_14749_),
    .B1(_14717_),
    .B2(net5888),
    .A2(_10369_),
    .A1(net5973));
 sg13g2_o21ai_1 _45577_ (.B1(_14749_),
    .Y(_14750_),
    .A1(_14747_),
    .A2(_14748_));
 sg13g2_nor2b_1 _45578_ (.A(_14750_),
    .B_N(net5246),
    .Y(_14751_));
 sg13g2_o21ai_1 _45579_ (.B1(net6867),
    .Y(_14752_),
    .A1(net5246),
    .A2(_10369_));
 sg13g2_o21ai_1 _45580_ (.B1(_14728_),
    .Y(_00976_),
    .A1(_14751_),
    .A2(_14752_));
 sg13g2_a21oi_1 _45581_ (.A1(_10769_),
    .A2(_14713_),
    .Y(_14753_),
    .B1(_10320_));
 sg13g2_xor2_1 _45582_ (.B(_14753_),
    .A(_10311_),
    .X(_14754_));
 sg13g2_nand2_1 _45583_ (.Y(_14755_),
    .A(net5684),
    .B(_10307_));
 sg13g2_o21ai_1 _45584_ (.B1(_14755_),
    .Y(_14756_),
    .A1(net5684),
    .A2(_14754_));
 sg13g2_inv_1 _45585_ (.Y(_14757_),
    .A(_14756_));
 sg13g2_xnor2_1 _45586_ (.Y(_14758_),
    .A(net5372),
    .B(_14756_));
 sg13g2_inv_1 _45587_ (.Y(_14759_),
    .A(_14758_));
 sg13g2_nor2b_1 _45588_ (.A(_14733_),
    .B_N(_14744_),
    .Y(_14760_));
 sg13g2_xnor2_1 _45589_ (.Y(_14761_),
    .A(_14758_),
    .B(_14760_));
 sg13g2_o21ai_1 _45590_ (.B1(net5939),
    .Y(_14762_),
    .A1(net5484),
    .A2(_14756_));
 sg13g2_a21oi_1 _45591_ (.A1(net5478),
    .A2(_14761_),
    .Y(_14763_),
    .B1(_14762_));
 sg13g2_a221oi_1 _45592_ (.B2(net5888),
    .C1(_14763_),
    .B1(_14732_),
    .A1(net5973),
    .Y(_14764_),
    .A2(_10325_));
 sg13g2_o21ai_1 _45593_ (.B1(net6867),
    .Y(_14765_),
    .A1(net5246),
    .A2(_10325_));
 sg13g2_a21oi_1 _45594_ (.A1(net5246),
    .A2(_14764_),
    .Y(_14766_),
    .B1(_14765_));
 sg13g2_a21o_1 _45595_ (.A2(net6395),
    .A1(net3606),
    .B1(_14766_),
    .X(_00977_));
 sg13g2_nand2_1 _45596_ (.Y(_14767_),
    .A(net5692),
    .B(_10315_));
 sg13g2_a21oi_1 _45597_ (.A1(_10310_),
    .A2(_14753_),
    .Y(_14768_),
    .B1(_10308_));
 sg13g2_xnor2_1 _45598_ (.Y(_14769_),
    .A(_10316_),
    .B(_14768_));
 sg13g2_o21ai_1 _45599_ (.B1(_14767_),
    .Y(_14770_),
    .A1(net5684),
    .A2(_14769_));
 sg13g2_nor2_1 _45600_ (.A(net5478),
    .B(_14770_),
    .Y(_14771_));
 sg13g2_and2_1 _45601_ (.A(net5372),
    .B(_14770_),
    .X(_14772_));
 sg13g2_xnor2_1 _45602_ (.Y(_14773_),
    .A(net5432),
    .B(_14770_));
 sg13g2_a21oi_1 _45603_ (.A1(net5372),
    .A2(_14756_),
    .Y(_14774_),
    .B1(_14733_));
 sg13g2_inv_1 _45604_ (.Y(_14775_),
    .A(_14774_));
 sg13g2_a22oi_1 _45605_ (.Y(_14776_),
    .B1(_14774_),
    .B2(_14744_),
    .A2(_14757_),
    .A1(net5433));
 sg13g2_xnor2_1 _45606_ (.Y(_14777_),
    .A(_14773_),
    .B(_14776_));
 sg13g2_a21oi_1 _45607_ (.A1(net5478),
    .A2(_14777_),
    .Y(_14778_),
    .B1(_14771_));
 sg13g2_nand2_1 _45608_ (.Y(_14779_),
    .A(net5221),
    .B(_14778_));
 sg13g2_a22oi_1 _45609_ (.Y(_14780_),
    .B1(_14756_),
    .B2(net5200),
    .A2(_10319_),
    .A1(net5157));
 sg13g2_a21oi_1 _45610_ (.A1(_14779_),
    .A2(_14780_),
    .Y(_14781_),
    .B1(net6838));
 sg13g2_a21o_1 _45611_ (.A2(net6397),
    .A1(net3575),
    .B1(_14781_),
    .X(_00978_));
 sg13g2_nand2_1 _45612_ (.Y(_14782_),
    .A(net5684),
    .B(_10345_));
 sg13g2_a21oi_1 _45613_ (.A1(_10329_),
    .A2(_14712_),
    .Y(_14783_),
    .B1(_10772_));
 sg13g2_xnor2_1 _45614_ (.Y(_14784_),
    .A(_10348_),
    .B(_14783_));
 sg13g2_o21ai_1 _45615_ (.B1(_14782_),
    .Y(_14785_),
    .A1(net5684),
    .A2(_14784_));
 sg13g2_xnor2_1 _45616_ (.Y(_14786_),
    .A(net5433),
    .B(_14785_));
 sg13g2_a21oi_1 _45617_ (.A1(_14773_),
    .A2(_14776_),
    .Y(_14787_),
    .B1(_14772_));
 sg13g2_xor2_1 _45618_ (.B(_14787_),
    .A(_14786_),
    .X(_14788_));
 sg13g2_o21ai_1 _45619_ (.B1(net5939),
    .Y(_14789_),
    .A1(net5478),
    .A2(_14785_));
 sg13g2_a21o_1 _45620_ (.A2(_14788_),
    .A1(net5479),
    .B1(_14789_),
    .X(_14790_));
 sg13g2_a22oi_1 _45621_ (.Y(_14791_),
    .B1(_14770_),
    .B2(net5888),
    .A2(_10307_),
    .A1(net5973));
 sg13g2_nand3_1 _45622_ (.B(_14790_),
    .C(_14791_),
    .A(net5250),
    .Y(_14792_));
 sg13g2_nor2_1 _45623_ (.A(net5250),
    .B(_10307_),
    .Y(_14793_));
 sg13g2_nor2_1 _45624_ (.A(net6838),
    .B(_14793_),
    .Y(_14794_));
 sg13g2_a22oi_1 _45625_ (.Y(_14795_),
    .B1(_14792_),
    .B2(_14794_),
    .A2(net6397),
    .A1(net3601));
 sg13g2_inv_1 _45626_ (.Y(_00979_),
    .A(_14795_));
 sg13g2_o21ai_1 _45627_ (.B1(_10346_),
    .Y(_14796_),
    .A1(_10348_),
    .A2(_14783_));
 sg13g2_xor2_1 _45628_ (.B(_14796_),
    .A(_10352_),
    .X(_14797_));
 sg13g2_nor2_1 _45629_ (.A(net5743),
    .B(_10351_),
    .Y(_14798_));
 sg13g2_a21oi_2 _45630_ (.B1(_14798_),
    .Y(_14799_),
    .A2(_14797_),
    .A1(net5743));
 sg13g2_nor2_1 _45631_ (.A(net5478),
    .B(_14799_),
    .Y(_14800_));
 sg13g2_nand2_1 _45632_ (.Y(_14801_),
    .A(net5371),
    .B(_14799_));
 sg13g2_xnor2_1 _45633_ (.Y(_14802_),
    .A(net5371),
    .B(_14799_));
 sg13g2_inv_1 _45634_ (.Y(_14803_),
    .A(_14802_));
 sg13g2_and2_1 _45635_ (.A(_14773_),
    .B(_14786_),
    .X(_14804_));
 sg13g2_a22oi_1 _45636_ (.Y(_14805_),
    .B1(_14804_),
    .B2(_14775_),
    .A2(_14785_),
    .A1(net5372));
 sg13g2_nand2b_1 _45637_ (.Y(_14806_),
    .B(_14805_),
    .A_N(_14772_));
 sg13g2_and3_1 _45638_ (.X(_14807_),
    .A(_14734_),
    .B(_14759_),
    .C(_14804_));
 sg13g2_inv_1 _45639_ (.Y(_14808_),
    .A(_14807_));
 sg13g2_a21oi_1 _45640_ (.A1(_14740_),
    .A2(_14743_),
    .Y(_14809_),
    .B1(_14808_));
 sg13g2_nor2_1 _45641_ (.A(_14806_),
    .B(_14809_),
    .Y(_14810_));
 sg13g2_o21ai_1 _45642_ (.B1(_14803_),
    .Y(_14811_),
    .A1(_14806_),
    .A2(_14809_));
 sg13g2_xnor2_1 _45643_ (.Y(_14812_),
    .A(_14802_),
    .B(_14810_));
 sg13g2_a21oi_1 _45644_ (.A1(net5478),
    .A2(_14812_),
    .Y(_14813_),
    .B1(_14800_));
 sg13g2_a22oi_1 _45645_ (.Y(_14814_),
    .B1(_14813_),
    .B2(net5221),
    .A2(_14785_),
    .A1(net5200));
 sg13g2_a22oi_1 _45646_ (.Y(_14815_),
    .B1(net5096),
    .B2(_10315_),
    .A2(net6395),
    .A1(net2310));
 sg13g2_o21ai_1 _45647_ (.B1(_14815_),
    .Y(_00980_),
    .A1(net6838),
    .A2(_14814_));
 sg13g2_nor2_1 _45648_ (.A(net5743),
    .B(_10339_),
    .Y(_14816_));
 sg13g2_o21ai_1 _45649_ (.B1(_10773_),
    .Y(_14817_),
    .A1(_10348_),
    .A2(_14783_));
 sg13g2_o21ai_1 _45650_ (.B1(_14817_),
    .Y(_14818_),
    .A1(net5611),
    .A2(_10351_));
 sg13g2_xnor2_1 _45651_ (.Y(_14819_),
    .A(_10341_),
    .B(_14818_));
 sg13g2_a21oi_2 _45652_ (.B1(_14816_),
    .Y(_14820_),
    .A2(_14819_),
    .A1(net5743));
 sg13g2_inv_1 _45653_ (.Y(_14821_),
    .A(_14820_));
 sg13g2_xnor2_1 _45654_ (.Y(_14822_),
    .A(net5371),
    .B(_14820_));
 sg13g2_nand2_1 _45655_ (.Y(_14823_),
    .A(_14801_),
    .B(_14811_));
 sg13g2_xor2_1 _45656_ (.B(_14823_),
    .A(_14822_),
    .X(_14824_));
 sg13g2_o21ai_1 _45657_ (.B1(net5939),
    .Y(_14825_),
    .A1(net5478),
    .A2(_14820_));
 sg13g2_a21oi_1 _45658_ (.A1(net5478),
    .A2(_14824_),
    .Y(_14826_),
    .B1(_14825_));
 sg13g2_a22oi_1 _45659_ (.Y(_14827_),
    .B1(_14799_),
    .B2(net5888),
    .A2(_10345_),
    .A1(net5973));
 sg13g2_nand2_1 _45660_ (.Y(_14828_),
    .A(net5244),
    .B(_14827_));
 sg13g2_nor2_1 _45661_ (.A(net5244),
    .B(_10345_),
    .Y(_14829_));
 sg13g2_o21ai_1 _45662_ (.B1(net6870),
    .Y(_14830_),
    .A1(_14826_),
    .A2(_14828_));
 sg13g2_nand2_1 _45663_ (.Y(_14831_),
    .A(net2633),
    .B(net6397));
 sg13g2_o21ai_1 _45664_ (.B1(_14831_),
    .Y(_00981_),
    .A1(_14829_),
    .A2(_14830_));
 sg13g2_nand2_1 _45665_ (.Y(_14832_),
    .A(net1191),
    .B(net6397));
 sg13g2_nand2_1 _45666_ (.Y(_14833_),
    .A(net5684),
    .B(_10332_));
 sg13g2_o21ai_1 _45667_ (.B1(_10340_),
    .Y(_14834_),
    .A1(_10341_),
    .A2(_14818_));
 sg13g2_xor2_1 _45668_ (.B(_14834_),
    .A(_10334_),
    .X(_14835_));
 sg13g2_o21ai_1 _45669_ (.B1(_14833_),
    .Y(_14836_),
    .A1(net5684),
    .A2(_14835_));
 sg13g2_xnor2_1 _45670_ (.Y(_14837_),
    .A(net5371),
    .B(_14836_));
 sg13g2_o21ai_1 _45671_ (.B1(net5371),
    .Y(_14838_),
    .A1(_14799_),
    .A2(_14820_));
 sg13g2_a22oi_1 _45672_ (.Y(_14839_),
    .B1(_14838_),
    .B2(_14811_),
    .A2(_14821_),
    .A1(net5433));
 sg13g2_a221oi_1 _45673_ (.B2(_14811_),
    .C1(_14837_),
    .B1(_14838_),
    .A1(net5433),
    .Y(_14840_),
    .A2(_14821_));
 sg13g2_xor2_1 _45674_ (.B(_14839_),
    .A(_14837_),
    .X(_14841_));
 sg13g2_o21ai_1 _45675_ (.B1(net5940),
    .Y(_14842_),
    .A1(net5479),
    .A2(_14836_));
 sg13g2_a21oi_1 _45676_ (.A1(net5479),
    .A2(_14841_),
    .Y(_14843_),
    .B1(_14842_));
 sg13g2_a22oi_1 _45677_ (.Y(_14844_),
    .B1(_14820_),
    .B2(net5888),
    .A2(_10351_),
    .A1(net5973));
 sg13g2_nand2_1 _45678_ (.Y(_14845_),
    .A(net5244),
    .B(_14844_));
 sg13g2_nor2_1 _45679_ (.A(_14843_),
    .B(_14845_),
    .Y(_14846_));
 sg13g2_o21ai_1 _45680_ (.B1(net6870),
    .Y(_14847_),
    .A1(net5244),
    .A2(_10351_));
 sg13g2_o21ai_1 _45681_ (.B1(_14832_),
    .Y(_00982_),
    .A1(_14846_),
    .A2(_14847_));
 sg13g2_nand2_1 _45682_ (.Y(_14848_),
    .A(net2450),
    .B(net6397));
 sg13g2_nand2_1 _45683_ (.Y(_14849_),
    .A(net5682),
    .B(_10259_));
 sg13g2_nand2b_1 _45684_ (.Y(_14850_),
    .B(_14712_),
    .A_N(_10354_));
 sg13g2_and2_1 _45685_ (.A(_10776_),
    .B(_14850_),
    .X(_14851_));
 sg13g2_xnor2_1 _45686_ (.Y(_14852_),
    .A(_10261_),
    .B(_14851_));
 sg13g2_o21ai_1 _45687_ (.B1(_14849_),
    .Y(_14853_),
    .A1(net5683),
    .A2(_14852_));
 sg13g2_xnor2_1 _45688_ (.Y(_14854_),
    .A(net5432),
    .B(_14853_));
 sg13g2_a21oi_1 _45689_ (.A1(net5371),
    .A2(_14836_),
    .Y(_14855_),
    .B1(_14840_));
 sg13g2_xor2_1 _45690_ (.B(_14855_),
    .A(_14854_),
    .X(_14856_));
 sg13g2_o21ai_1 _45691_ (.B1(net5941),
    .Y(_14857_),
    .A1(net5477),
    .A2(_14853_));
 sg13g2_a21oi_1 _45692_ (.A1(net5479),
    .A2(_14856_),
    .Y(_14858_),
    .B1(_14857_));
 sg13g2_a22oi_1 _45693_ (.Y(_14859_),
    .B1(_14836_),
    .B2(net5888),
    .A2(_10339_),
    .A1(net5973));
 sg13g2_nand2_1 _45694_ (.Y(_14860_),
    .A(net5245),
    .B(_14859_));
 sg13g2_nor2_1 _45695_ (.A(_14858_),
    .B(_14860_),
    .Y(_14861_));
 sg13g2_o21ai_1 _45696_ (.B1(net6870),
    .Y(_14862_),
    .A1(net5244),
    .A2(_10339_));
 sg13g2_o21ai_1 _45697_ (.B1(_14848_),
    .Y(_00983_),
    .A1(_14861_),
    .A2(_14862_));
 sg13g2_nand2_1 _45698_ (.Y(_14863_),
    .A(net5682),
    .B(_10253_));
 sg13g2_o21ai_1 _45699_ (.B1(_10260_),
    .Y(_14864_),
    .A1(_10261_),
    .A2(_14851_));
 sg13g2_o21ai_1 _45700_ (.B1(_14864_),
    .Y(_14865_),
    .A1(net5609),
    .A2(_10253_));
 sg13g2_xor2_1 _45701_ (.B(_14864_),
    .A(_10255_),
    .X(_14866_));
 sg13g2_o21ai_1 _45702_ (.B1(_14863_),
    .Y(_14867_),
    .A1(net5682),
    .A2(_14866_));
 sg13g2_nor2_1 _45703_ (.A(net5477),
    .B(_14867_),
    .Y(_14868_));
 sg13g2_nand2_1 _45704_ (.Y(_14869_),
    .A(net5370),
    .B(_14867_));
 sg13g2_xnor2_1 _45705_ (.Y(_14870_),
    .A(net5373),
    .B(_14867_));
 sg13g2_inv_1 _45706_ (.Y(_14871_),
    .A(_14870_));
 sg13g2_nand2b_1 _45707_ (.Y(_14872_),
    .B(_14854_),
    .A_N(_14837_));
 sg13g2_nor3_1 _45708_ (.A(_14802_),
    .B(_14822_),
    .C(_14872_),
    .Y(_14873_));
 sg13g2_and2_1 _45709_ (.A(_14807_),
    .B(_14873_),
    .X(_14874_));
 sg13g2_inv_1 _45710_ (.Y(_14875_),
    .A(_14874_));
 sg13g2_a21oi_1 _45711_ (.A1(_14740_),
    .A2(_14743_),
    .Y(_14876_),
    .B1(_14875_));
 sg13g2_o21ai_1 _45712_ (.B1(net5371),
    .Y(_14877_),
    .A1(_14836_),
    .A2(_14853_));
 sg13g2_o21ai_1 _45713_ (.B1(_14877_),
    .Y(_14878_),
    .A1(_14838_),
    .A2(_14872_));
 sg13g2_a21o_1 _45714_ (.A2(_14873_),
    .A1(_14806_),
    .B1(_14878_),
    .X(_14879_));
 sg13g2_o21ai_1 _45715_ (.B1(_14871_),
    .Y(_14880_),
    .A1(_14876_),
    .A2(_14879_));
 sg13g2_or3_1 _45716_ (.A(_14871_),
    .B(_14876_),
    .C(_14879_),
    .X(_14881_));
 sg13g2_nand2_1 _45717_ (.Y(_14882_),
    .A(_14880_),
    .B(_14881_));
 sg13g2_a21oi_1 _45718_ (.A1(net5480),
    .A2(_14882_),
    .Y(_14883_),
    .B1(_14868_));
 sg13g2_a22oi_1 _45719_ (.Y(_14884_),
    .B1(_14883_),
    .B2(net5222),
    .A2(_14853_),
    .A1(net5201));
 sg13g2_a22oi_1 _45720_ (.Y(_14885_),
    .B1(net5096),
    .B2(_10332_),
    .A2(net6397),
    .A1(net3017));
 sg13g2_o21ai_1 _45721_ (.B1(_14885_),
    .Y(_00984_),
    .A1(net6838),
    .A2(_14884_));
 sg13g2_nand2_1 _45722_ (.Y(_14886_),
    .A(_14869_),
    .B(_14880_));
 sg13g2_nand2_1 _45723_ (.Y(_14887_),
    .A(_10254_),
    .B(_14865_));
 sg13g2_xnor2_1 _45724_ (.Y(_14888_),
    .A(_10242_),
    .B(_14887_));
 sg13g2_nor2_1 _45725_ (.A(net5682),
    .B(_14888_),
    .Y(_14889_));
 sg13g2_a21oi_2 _45726_ (.B1(_14889_),
    .Y(_14890_),
    .A2(_10238_),
    .A1(net5682));
 sg13g2_nor2_1 _45727_ (.A(net5370),
    .B(_14890_),
    .Y(_14891_));
 sg13g2_xnor2_1 _45728_ (.Y(_14892_),
    .A(net5370),
    .B(_14890_));
 sg13g2_xor2_1 _45729_ (.B(_14892_),
    .A(_14886_),
    .X(_14893_));
 sg13g2_o21ai_1 _45730_ (.B1(net5222),
    .Y(_14894_),
    .A1(net5477),
    .A2(_14890_));
 sg13g2_a21oi_1 _45731_ (.A1(net5477),
    .A2(_14893_),
    .Y(_14895_),
    .B1(_14894_));
 sg13g2_a21oi_1 _45732_ (.A1(net5202),
    .A2(_14867_),
    .Y(_14896_),
    .B1(_14895_));
 sg13g2_a22oi_1 _45733_ (.Y(_14897_),
    .B1(net5095),
    .B2(_10259_),
    .A2(net6393),
    .A1(net3543));
 sg13g2_o21ai_1 _45734_ (.B1(_14897_),
    .Y(_00985_),
    .A1(net6837),
    .A2(_14896_));
 sg13g2_nand2_1 _45735_ (.Y(_14898_),
    .A(net5682),
    .B(_10247_));
 sg13g2_a21oi_1 _45736_ (.A1(_10241_),
    .A2(_14887_),
    .Y(_14899_),
    .B1(_10239_));
 sg13g2_xnor2_1 _45737_ (.Y(_14900_),
    .A(_10249_),
    .B(_14899_));
 sg13g2_o21ai_1 _45738_ (.B1(_14898_),
    .Y(_14901_),
    .A1(net5682),
    .A2(_14900_));
 sg13g2_and2_1 _45739_ (.A(net5370),
    .B(_14901_),
    .X(_14902_));
 sg13g2_xnor2_1 _45740_ (.Y(_14903_),
    .A(net5432),
    .B(_14901_));
 sg13g2_o21ai_1 _45741_ (.B1(net5370),
    .Y(_14904_),
    .A1(_14867_),
    .A2(_14890_));
 sg13g2_a21oi_1 _45742_ (.A1(_14880_),
    .A2(_14904_),
    .Y(_14905_),
    .B1(_14891_));
 sg13g2_xnor2_1 _45743_ (.Y(_14906_),
    .A(_14903_),
    .B(_14905_));
 sg13g2_a21oi_1 _45744_ (.A1(net5477),
    .A2(_14906_),
    .Y(_14907_),
    .B1(net5151));
 sg13g2_o21ai_1 _45745_ (.B1(_14907_),
    .Y(_14908_),
    .A1(net5477),
    .A2(_14901_));
 sg13g2_a22oi_1 _45746_ (.Y(_14909_),
    .B1(_14890_),
    .B2(net5202),
    .A2(_10253_),
    .A1(net5157));
 sg13g2_a21oi_1 _45747_ (.A1(_14908_),
    .A2(_14909_),
    .Y(_14910_),
    .B1(net6837));
 sg13g2_a21o_1 _45748_ (.A2(net6390),
    .A1(net3504),
    .B1(_14910_),
    .X(_00986_));
 sg13g2_nand2b_1 _45749_ (.Y(_14911_),
    .B(_10262_),
    .A_N(_14851_));
 sg13g2_a21oi_1 _45750_ (.A1(_10780_),
    .A2(_14911_),
    .Y(_14912_),
    .B1(_10287_));
 sg13g2_and3_1 _45751_ (.X(_14913_),
    .A(_10287_),
    .B(_10780_),
    .C(_14911_));
 sg13g2_nor3_1 _45752_ (.A(net5683),
    .B(_14912_),
    .C(_14913_),
    .Y(_14914_));
 sg13g2_a21oi_2 _45753_ (.B1(_14914_),
    .Y(_14915_),
    .A2(_10284_),
    .A1(net5682));
 sg13g2_inv_1 _45754_ (.Y(_14916_),
    .A(_14915_));
 sg13g2_nor2_1 _45755_ (.A(net5432),
    .B(_14915_),
    .Y(_14917_));
 sg13g2_xnor2_1 _45756_ (.Y(_14918_),
    .A(net5373),
    .B(_14915_));
 sg13g2_a21oi_1 _45757_ (.A1(_14903_),
    .A2(_14905_),
    .Y(_14919_),
    .B1(_14902_));
 sg13g2_xnor2_1 _45758_ (.Y(_14920_),
    .A(_14918_),
    .B(_14919_));
 sg13g2_a21oi_1 _45759_ (.A1(net5552),
    .A2(_14915_),
    .Y(_14921_),
    .B1(net5920));
 sg13g2_o21ai_1 _45760_ (.B1(_14921_),
    .Y(_14922_),
    .A1(net5552),
    .A2(_14920_));
 sg13g2_nor2_1 _45761_ (.A(net6003),
    .B(_10238_),
    .Y(_14923_));
 sg13g2_a21oi_1 _45762_ (.A1(net5886),
    .A2(_14901_),
    .Y(_14924_),
    .B1(_14923_));
 sg13g2_and3_1 _45763_ (.X(_14925_),
    .A(net5257),
    .B(_14922_),
    .C(_14924_));
 sg13g2_nand3_1 _45764_ (.B(net5315),
    .C(_10238_),
    .A(net5319),
    .Y(_14926_));
 sg13g2_nand2_1 _45765_ (.Y(_14927_),
    .A(net6870),
    .B(_14926_));
 sg13g2_nand2_1 _45766_ (.Y(_14928_),
    .A(net2880),
    .B(net6393));
 sg13g2_o21ai_1 _45767_ (.B1(_14928_),
    .Y(_00987_),
    .A1(_14925_),
    .A2(_14927_));
 sg13g2_nand2_1 _45768_ (.Y(_14929_),
    .A(net2809),
    .B(net6390));
 sg13g2_nor2_1 _45769_ (.A(net5743),
    .B(_10292_),
    .Y(_14930_));
 sg13g2_a21oi_1 _45770_ (.A1(net5608),
    .A2(_10284_),
    .Y(_14931_),
    .B1(_14912_));
 sg13g2_xnor2_1 _45771_ (.Y(_14932_),
    .A(_10295_),
    .B(_14931_));
 sg13g2_a21oi_2 _45772_ (.B1(_14930_),
    .Y(_14933_),
    .A2(_14932_),
    .A1(net5743));
 sg13g2_nor2_1 _45773_ (.A(net5432),
    .B(_14933_),
    .Y(_14934_));
 sg13g2_nand2_1 _45774_ (.Y(_14935_),
    .A(net5432),
    .B(_14933_));
 sg13g2_nand2b_1 _45775_ (.Y(_14936_),
    .B(_14935_),
    .A_N(_14934_));
 sg13g2_nand2_1 _45776_ (.Y(_14937_),
    .A(_14903_),
    .B(_14918_));
 sg13g2_or2_1 _45777_ (.X(_14938_),
    .B(_14937_),
    .A(_14892_));
 sg13g2_nor2_1 _45778_ (.A(_14904_),
    .B(_14937_),
    .Y(_14939_));
 sg13g2_nor3_1 _45779_ (.A(_14902_),
    .B(_14917_),
    .C(_14939_),
    .Y(_14940_));
 sg13g2_o21ai_1 _45780_ (.B1(_14940_),
    .Y(_14941_),
    .A1(_14880_),
    .A2(_14938_));
 sg13g2_xnor2_1 _45781_ (.Y(_14942_),
    .A(_14936_),
    .B(_14941_));
 sg13g2_a21oi_1 _45782_ (.A1(net5552),
    .A2(_14933_),
    .Y(_14943_),
    .B1(net5920));
 sg13g2_o21ai_1 _45783_ (.B1(_14943_),
    .Y(_14944_),
    .A1(net5552),
    .A2(_14942_));
 sg13g2_a22oi_1 _45784_ (.Y(_14945_),
    .B1(_14916_),
    .B2(net5886),
    .A2(_10247_),
    .A1(net5970));
 sg13g2_nand3_1 _45785_ (.B(_14944_),
    .C(_14945_),
    .A(net5244),
    .Y(_14946_));
 sg13g2_o21ai_1 _45786_ (.B1(_14946_),
    .Y(_14947_),
    .A1(net5244),
    .A2(_10247_));
 sg13g2_o21ai_1 _45787_ (.B1(_14929_),
    .Y(_00988_),
    .A1(net6837),
    .A2(_14947_));
 sg13g2_a21oi_1 _45788_ (.A1(_14935_),
    .A2(_14941_),
    .Y(_14948_),
    .B1(_14934_));
 sg13g2_nand2_1 _45789_ (.Y(_14949_),
    .A(net5683),
    .B(_10274_));
 sg13g2_o21ai_1 _45790_ (.B1(_10293_),
    .Y(_14950_),
    .A1(_10782_),
    .A2(_14912_));
 sg13g2_nor2_1 _45791_ (.A(_10277_),
    .B(_14950_),
    .Y(_14951_));
 sg13g2_xor2_1 _45792_ (.B(_14950_),
    .A(_10277_),
    .X(_14952_));
 sg13g2_o21ai_1 _45793_ (.B1(_14949_),
    .Y(_14953_),
    .A1(net5683),
    .A2(_14952_));
 sg13g2_inv_1 _45794_ (.Y(_14954_),
    .A(_14953_));
 sg13g2_nor2_1 _45795_ (.A(net5370),
    .B(_14954_),
    .Y(_14955_));
 sg13g2_nand2_1 _45796_ (.Y(_14956_),
    .A(net5370),
    .B(_14954_));
 sg13g2_nor2b_1 _45797_ (.A(_14955_),
    .B_N(_14956_),
    .Y(_14957_));
 sg13g2_a21oi_1 _45798_ (.A1(_14948_),
    .A2(_14957_),
    .Y(_14958_),
    .B1(net5552));
 sg13g2_o21ai_1 _45799_ (.B1(_14958_),
    .Y(_14959_),
    .A1(_14948_),
    .A2(_14957_));
 sg13g2_a21oi_1 _45800_ (.A1(net5552),
    .A2(_14953_),
    .Y(_14960_),
    .B1(net5920));
 sg13g2_nand2_1 _45801_ (.Y(_14961_),
    .A(net5970),
    .B(_10284_));
 sg13g2_o21ai_1 _45802_ (.B1(_14961_),
    .Y(_14962_),
    .A1(net5880),
    .A2(_14933_));
 sg13g2_a221oi_1 _45803_ (.B2(_14960_),
    .C1(_14962_),
    .B1(_14959_),
    .A1(net5319),
    .Y(_14963_),
    .A2(net5315));
 sg13g2_o21ai_1 _45804_ (.B1(net6870),
    .Y(_14964_),
    .A1(net5244),
    .A2(_10284_));
 sg13g2_nand2_1 _45805_ (.Y(_14965_),
    .A(net3347),
    .B(net6393));
 sg13g2_o21ai_1 _45806_ (.B1(_14965_),
    .Y(_00989_),
    .A1(_14963_),
    .A2(_14964_));
 sg13g2_o21ai_1 _45807_ (.B1(_14956_),
    .Y(_14966_),
    .A1(_14948_),
    .A2(_14955_));
 sg13g2_nor2_1 _45808_ (.A(_10275_),
    .B(_14951_),
    .Y(_14967_));
 sg13g2_xnor2_1 _45809_ (.Y(_14968_),
    .A(_10267_),
    .B(_14967_));
 sg13g2_nor2_1 _45810_ (.A(net5683),
    .B(_14968_),
    .Y(_14969_));
 sg13g2_a21oi_2 _45811_ (.B1(_14969_),
    .Y(_14970_),
    .A2(_10266_),
    .A1(net5683));
 sg13g2_xnor2_1 _45812_ (.Y(_14971_),
    .A(net5370),
    .B(_14970_));
 sg13g2_or3_1 _45813_ (.A(net5552),
    .B(_14966_),
    .C(_14971_),
    .X(_14972_));
 sg13g2_and2_1 _45814_ (.A(net5477),
    .B(_14971_),
    .X(_14973_));
 sg13g2_a221oi_1 _45815_ (.B2(_14966_),
    .C1(net5151),
    .B1(_14973_),
    .A1(net5552),
    .Y(_14974_),
    .A2(_14970_));
 sg13g2_nor2_1 _45816_ (.A(net5241),
    .B(_10292_),
    .Y(_14975_));
 sg13g2_a221oi_1 _45817_ (.B2(_14974_),
    .C1(_14975_),
    .B1(_14972_),
    .A1(net5202),
    .Y(_14976_),
    .A2(_14954_));
 sg13g2_nand2_1 _45818_ (.Y(_14977_),
    .A(net3493),
    .B(net6390));
 sg13g2_o21ai_1 _45819_ (.B1(_14977_),
    .Y(_00990_),
    .A1(net6837),
    .A2(_14976_));
 sg13g2_a21oi_1 _45820_ (.A1(net5477),
    .A2(_14970_),
    .Y(_14978_),
    .B1(net5432));
 sg13g2_a21o_1 _45821_ (.A2(_14973_),
    .A1(_14966_),
    .B1(_14978_),
    .X(_14979_));
 sg13g2_nand3_1 _45822_ (.B(_10268_),
    .C(_10273_),
    .A(net5970),
    .Y(_14980_));
 sg13g2_o21ai_1 _45823_ (.B1(_14980_),
    .Y(_14981_),
    .A1(net5880),
    .A2(_14970_));
 sg13g2_a221oi_1 _45824_ (.B2(_14979_),
    .C1(_14981_),
    .B1(net5941),
    .A1(net5319),
    .Y(_14982_),
    .A2(net5315));
 sg13g2_nand3_1 _45825_ (.B(net5315),
    .C(_10274_),
    .A(net5319),
    .Y(_14983_));
 sg13g2_nand2_1 _45826_ (.Y(_14984_),
    .A(net6870),
    .B(_14983_));
 sg13g2_nand2_1 _45827_ (.Y(_14985_),
    .A(net2888),
    .B(net6390));
 sg13g2_o21ai_1 _45828_ (.B1(_14985_),
    .Y(_00991_),
    .A1(_14982_),
    .A2(_14984_));
 sg13g2_nor2_1 _45829_ (.A(net5257),
    .B(_10266_),
    .Y(_14986_));
 sg13g2_xnor2_1 _45830_ (.Y(_14987_),
    .A(net5480),
    .B(net5439));
 sg13g2_a22oi_1 _45831_ (.Y(_14988_),
    .B1(_14987_),
    .B2(net5941),
    .A2(net5382),
    .A1(net5886));
 sg13g2_nand2_1 _45832_ (.Y(_14989_),
    .A(net5970),
    .B(_10266_));
 sg13g2_nand3_1 _45833_ (.B(_14988_),
    .C(_14989_),
    .A(net5257),
    .Y(_14990_));
 sg13g2_nor2_1 _45834_ (.A(net6837),
    .B(_14986_),
    .Y(_14991_));
 sg13g2_a22oi_1 _45835_ (.Y(_14992_),
    .B1(_14990_),
    .B2(_14991_),
    .A2(net6401),
    .A1(net3405));
 sg13g2_inv_1 _45836_ (.Y(_00992_),
    .A(_14992_));
 sg13g2_nand2_1 _45837_ (.Y(_14993_),
    .A(net2988),
    .B(net6401));
 sg13g2_nand2_1 _45838_ (.Y(_14994_),
    .A(net5970),
    .B(net5613));
 sg13g2_and3_1 _45839_ (.X(_14995_),
    .A(net5257),
    .B(_14988_),
    .C(_14994_));
 sg13g2_o21ai_1 _45840_ (.B1(net6870),
    .Y(_14996_),
    .A1(net5257),
    .A2(net5613));
 sg13g2_o21ai_1 _45841_ (.B1(_14993_),
    .Y(_00993_),
    .A1(_14995_),
    .A2(_14996_));
 sg13g2_a21oi_1 _45842_ (.A1(inv_done),
    .A2(_18625_),
    .Y(_14997_),
    .B1(_18623_));
 sg13g2_nand2_2 _45843_ (.Y(_14998_),
    .A(_18622_),
    .B(_18626_));
 sg13g2_nor2_1 _45844_ (.A(net3591),
    .B(net6698),
    .Y(_14999_));
 sg13g2_nand2_2 _45845_ (.Y(_15000_),
    .A(_18445_),
    .B(_18446_));
 sg13g2_nor3_2 _45846_ (.A(\u_inv.d_reg[171] ),
    .B(\u_inv.d_reg[170] ),
    .C(_15000_),
    .Y(_15001_));
 sg13g2_nor3_1 _45847_ (.A(\u_inv.d_reg[174] ),
    .B(\u_inv.d_reg[173] ),
    .C(\u_inv.d_reg[172] ),
    .Y(_15002_));
 sg13g2_nand2_1 _45848_ (.Y(_15003_),
    .A(_15001_),
    .B(_15002_));
 sg13g2_nand4_1 _45849_ (.B(_18460_),
    .C(_18461_),
    .A(_18459_),
    .Y(_15004_),
    .D(_18462_));
 sg13g2_nor4_1 _45850_ (.A(\u_inv.d_reg[157] ),
    .B(\u_inv.d_reg[156] ),
    .C(\u_inv.d_reg[151] ),
    .D(_15004_),
    .Y(_15005_));
 sg13g2_nand4_1 _45851_ (.B(_18465_),
    .C(_18466_),
    .A(_18464_),
    .Y(_15006_),
    .D(_15005_));
 sg13g2_nand2_1 _45852_ (.Y(_15007_),
    .A(_18469_),
    .B(_18470_));
 sg13g2_nand3_1 _45853_ (.B(_18469_),
    .C(_18470_),
    .A(_18468_),
    .Y(_15008_));
 sg13g2_nor3_1 _45854_ (.A(\u_inv.d_reg[0] ),
    .B(\u_inv.d_reg[2] ),
    .C(net7293),
    .Y(_15009_));
 sg13g2_nand3_1 _45855_ (.B(_18612_),
    .C(_18613_),
    .A(_18357_),
    .Y(_15010_));
 sg13g2_or4_1 _45856_ (.A(net7293),
    .B(\u_inv.d_reg[3] ),
    .C(\u_inv.d_reg[2] ),
    .D(net7294),
    .X(_15011_));
 sg13g2_nand2b_1 _45857_ (.Y(_15012_),
    .B(_18610_),
    .A_N(_15011_));
 sg13g2_or4_1 _45858_ (.A(_15011_),
    .B(\u_inv.d_reg[5] ),
    .C(\u_inv.d_reg[4] ),
    .D(\u_inv.d_reg[6] ),
    .X(_15013_));
 sg13g2_nor3_1 _45859_ (.A(\u_inv.d_reg[8] ),
    .B(\u_inv.d_reg[7] ),
    .C(_15013_),
    .Y(_15014_));
 sg13g2_or4_1 _45860_ (.A(\u_inv.d_reg[9] ),
    .B(_15013_),
    .C(\u_inv.d_reg[7] ),
    .D(\u_inv.d_reg[8] ),
    .X(_15015_));
 sg13g2_nor3_1 _45861_ (.A(\u_inv.d_reg[11] ),
    .B(\u_inv.d_reg[10] ),
    .C(_15015_),
    .Y(_15016_));
 sg13g2_or4_1 _45862_ (.A(\u_inv.d_reg[12] ),
    .B(\u_inv.d_reg[11] ),
    .C(_15015_),
    .D(net7292),
    .X(_15017_));
 sg13g2_nor3_1 _45863_ (.A(\u_inv.d_reg[14] ),
    .B(\u_inv.d_reg[13] ),
    .C(_15017_),
    .Y(_15018_));
 sg13g2_nor4_2 _45864_ (.A(\u_inv.d_reg[15] ),
    .B(_15017_),
    .C(\u_inv.d_reg[13] ),
    .Y(_15019_),
    .D(\u_inv.d_reg[14] ));
 sg13g2_and2_1 _45865_ (.A(_18598_),
    .B(_15019_),
    .X(_15020_));
 sg13g2_nand4_1 _45866_ (.B(_18597_),
    .C(_18598_),
    .A(_15019_),
    .Y(_15021_),
    .D(_18596_));
 sg13g2_nor3_1 _45867_ (.A(\u_inv.d_reg[20] ),
    .B(\u_inv.d_reg[19] ),
    .C(net1096),
    .Y(_15022_));
 sg13g2_or4_1 _45868_ (.A(\u_inv.d_reg[21] ),
    .B(\u_inv.d_reg[20] ),
    .C(net1096),
    .D(\u_inv.d_reg[19] ),
    .X(_15023_));
 sg13g2_nor3_1 _45869_ (.A(\u_inv.d_reg[23] ),
    .B(net7291),
    .C(_15023_),
    .Y(_15024_));
 sg13g2_or4_1 _45870_ (.A(\u_inv.d_reg[24] ),
    .B(\u_inv.d_reg[23] ),
    .C(_15023_),
    .D(\u_inv.d_reg[22] ),
    .X(_15025_));
 sg13g2_nor3_1 _45871_ (.A(\u_inv.d_reg[26] ),
    .B(\u_inv.d_reg[25] ),
    .C(_15025_),
    .Y(_15026_));
 sg13g2_or4_1 _45872_ (.A(\u_inv.d_reg[27] ),
    .B(\u_inv.d_reg[26] ),
    .C(_15025_),
    .D(\u_inv.d_reg[25] ),
    .X(_15027_));
 sg13g2_nor3_1 _45873_ (.A(\u_inv.d_reg[29] ),
    .B(\u_inv.d_reg[28] ),
    .C(_15027_),
    .Y(_15028_));
 sg13g2_nor4_2 _45874_ (.A(\u_inv.d_reg[30] ),
    .B(_15027_),
    .C(\u_inv.d_reg[28] ),
    .Y(_15029_),
    .D(\u_inv.d_reg[29] ));
 sg13g2_nand2_1 _45875_ (.Y(_15030_),
    .A(_18583_),
    .B(_15029_));
 sg13g2_and4_1 _45876_ (.A(_15029_),
    .B(_18582_),
    .C(_18583_),
    .D(_18581_),
    .X(_15031_));
 sg13g2_nand2_1 _45877_ (.Y(_15032_),
    .A(_18580_),
    .B(_15031_));
 sg13g2_nand4_1 _45878_ (.B(_18579_),
    .C(_18580_),
    .A(_15031_),
    .Y(_15033_),
    .D(_18578_));
 sg13g2_nand2b_1 _45879_ (.Y(_15034_),
    .B(_18577_),
    .A_N(net1137));
 sg13g2_nor4_2 _45880_ (.A(\u_inv.d_reg[39] ),
    .B(\u_inv.d_reg[38] ),
    .C(net1107),
    .Y(_15035_),
    .D(\u_inv.d_reg[37] ));
 sg13g2_nor2_1 _45881_ (.A(\u_inv.d_reg[41] ),
    .B(\u_inv.d_reg[40] ),
    .Y(_15036_));
 sg13g2_nand2_1 _45882_ (.Y(_15037_),
    .A(_15035_),
    .B(_15036_));
 sg13g2_and4_2 _45883_ (.A(_15035_),
    .B(_18572_),
    .C(_18571_),
    .D(_15036_),
    .X(_15038_));
 sg13g2_nor4_1 _45884_ (.A(\u_inv.d_reg[47] ),
    .B(\u_inv.d_reg[46] ),
    .C(\u_inv.d_reg[45] ),
    .D(\u_inv.d_reg[44] ),
    .Y(_15039_));
 sg13g2_nand2_1 _45885_ (.Y(_15040_),
    .A(_15038_),
    .B(_15039_));
 sg13g2_nor2_1 _45886_ (.A(\u_inv.d_reg[49] ),
    .B(\u_inv.d_reg[48] ),
    .Y(_15041_));
 sg13g2_nand3_1 _45887_ (.B(_15039_),
    .C(_15041_),
    .A(_15038_),
    .Y(_15042_));
 sg13g2_nand4_1 _45888_ (.B(_18564_),
    .C(_15039_),
    .A(_15038_),
    .Y(_15043_),
    .D(_15041_));
 sg13g2_nor3_1 _45889_ (.A(\u_inv.d_reg[52] ),
    .B(\u_inv.d_reg[51] ),
    .C(net1091),
    .Y(_15044_));
 sg13g2_nor4_2 _45890_ (.A(net1091),
    .B(\u_inv.d_reg[52] ),
    .C(\u_inv.d_reg[51] ),
    .Y(_15045_),
    .D(\u_inv.d_reg[53] ));
 sg13g2_nor2_2 _45891_ (.A(\u_inv.d_reg[55] ),
    .B(\u_inv.d_reg[54] ),
    .Y(_15046_));
 sg13g2_nand2_1 _45892_ (.Y(_15047_),
    .A(_15045_),
    .B(_15046_));
 sg13g2_nor2_1 _45893_ (.A(\u_inv.d_reg[57] ),
    .B(\u_inv.d_reg[56] ),
    .Y(_15048_));
 sg13g2_nand3_1 _45894_ (.B(_15046_),
    .C(_15048_),
    .A(net1090),
    .Y(_15049_));
 sg13g2_nand4_1 _45895_ (.B(_18556_),
    .C(_15046_),
    .A(_15045_),
    .Y(_15050_),
    .D(_15048_));
 sg13g2_nor3_1 _45896_ (.A(\u_inv.d_reg[60] ),
    .B(\u_inv.d_reg[59] ),
    .C(net1084),
    .Y(_15051_));
 sg13g2_nor4_2 _45897_ (.A(\u_inv.d_reg[61] ),
    .B(\u_inv.d_reg[60] ),
    .C(net1084),
    .Y(_15052_),
    .D(\u_inv.d_reg[59] ));
 sg13g2_nor2_2 _45898_ (.A(\u_inv.d_reg[63] ),
    .B(\u_inv.d_reg[62] ),
    .Y(_15053_));
 sg13g2_nand2_1 _45899_ (.Y(_15054_),
    .A(net1072),
    .B(_15053_));
 sg13g2_nor3_1 _45900_ (.A(\u_inv.d_reg[65] ),
    .B(\u_inv.d_reg[64] ),
    .C(_15054_),
    .Y(_15055_));
 sg13g2_and2_1 _45901_ (.A(_18548_),
    .B(_15055_),
    .X(_15056_));
 sg13g2_nor4_1 _45902_ (.A(\u_inv.d_reg[67] ),
    .B(\u_inv.d_reg[66] ),
    .C(\u_inv.d_reg[65] ),
    .D(\u_inv.d_reg[64] ),
    .Y(_15057_));
 sg13g2_nand2_1 _45903_ (.Y(_15058_),
    .A(_18547_),
    .B(_15056_));
 sg13g2_nor2_1 _45904_ (.A(\u_inv.d_reg[69] ),
    .B(\u_inv.d_reg[68] ),
    .Y(_15059_));
 sg13g2_nand4_1 _45905_ (.B(_15053_),
    .C(_15057_),
    .A(net1072),
    .Y(_15060_),
    .D(_15059_));
 sg13g2_nand2_1 _45906_ (.Y(_15061_),
    .A(_18543_),
    .B(_18544_));
 sg13g2_or2_1 _45907_ (.X(_15062_),
    .B(_15061_),
    .A(net1100));
 sg13g2_nand2_1 _45908_ (.Y(_15063_),
    .A(_18541_),
    .B(_18542_));
 sg13g2_or4_1 _45909_ (.A(\u_inv.d_reg[74] ),
    .B(_15063_),
    .C(_15061_),
    .D(net1100),
    .X(_15064_));
 sg13g2_nand2b_1 _45910_ (.Y(_15065_),
    .B(_18539_),
    .A_N(_15064_));
 sg13g2_nor2_1 _45911_ (.A(\u_inv.d_reg[76] ),
    .B(_15065_),
    .Y(_15066_));
 sg13g2_nor2_1 _45912_ (.A(\u_inv.d_reg[78] ),
    .B(\u_inv.d_reg[77] ),
    .Y(_15067_));
 sg13g2_nand3_1 _45913_ (.B(_18538_),
    .C(_15067_),
    .A(_18535_),
    .Y(_15068_));
 sg13g2_nor2_1 _45914_ (.A(_15065_),
    .B(_15068_),
    .Y(_15069_));
 sg13g2_nor4_2 _45915_ (.A(\u_inv.d_reg[80] ),
    .B(\u_inv.d_reg[75] ),
    .C(_15068_),
    .Y(_15070_),
    .D(_15064_));
 sg13g2_nor3_1 _45916_ (.A(\u_inv.d_reg[83] ),
    .B(\u_inv.d_reg[82] ),
    .C(net7290),
    .Y(_15071_));
 sg13g2_nand2_1 _45917_ (.Y(_15072_),
    .A(net1095),
    .B(_15071_));
 sg13g2_nor2_1 _45918_ (.A(\u_inv.d_reg[85] ),
    .B(\u_inv.d_reg[84] ),
    .Y(_15073_));
 sg13g2_nand3_1 _45919_ (.B(_15071_),
    .C(_15073_),
    .A(net1095),
    .Y(_15074_));
 sg13g2_nor2_1 _45920_ (.A(\u_inv.d_reg[87] ),
    .B(\u_inv.d_reg[86] ),
    .Y(_15075_));
 sg13g2_nand4_1 _45921_ (.B(_15071_),
    .C(_15073_),
    .A(_15075_),
    .Y(_15076_),
    .D(net1095));
 sg13g2_nand2_1 _45922_ (.Y(_15077_),
    .A(_18525_),
    .B(_18526_));
 sg13g2_or2_1 _45923_ (.X(_15078_),
    .B(_15077_),
    .A(net1082));
 sg13g2_nor4_2 _45924_ (.A(\u_inv.d_reg[91] ),
    .B(\u_inv.d_reg[90] ),
    .C(_15077_),
    .Y(_15079_),
    .D(net1082));
 sg13g2_nor4_1 _45925_ (.A(\u_inv.d_reg[95] ),
    .B(\u_inv.d_reg[94] ),
    .C(\u_inv.d_reg[93] ),
    .D(\u_inv.d_reg[92] ),
    .Y(_15080_));
 sg13g2_nand2_1 _45926_ (.Y(_15081_),
    .A(_18517_),
    .B(_18518_));
 sg13g2_nor3_1 _45927_ (.A(\u_inv.d_reg[99] ),
    .B(\u_inv.d_reg[98] ),
    .C(_15081_),
    .Y(_15082_));
 sg13g2_nand3_1 _45928_ (.B(_15080_),
    .C(_15082_),
    .A(_15079_),
    .Y(_15083_));
 sg13g2_nor2_1 _45929_ (.A(\u_inv.d_reg[101] ),
    .B(\u_inv.d_reg[100] ),
    .Y(_15084_));
 sg13g2_nand4_1 _45930_ (.B(_15080_),
    .C(_15082_),
    .A(_15084_),
    .Y(_15085_),
    .D(_15079_));
 sg13g2_nand2_1 _45931_ (.Y(_15086_),
    .A(_18511_),
    .B(_18512_));
 sg13g2_or2_1 _45932_ (.X(_15087_),
    .B(_15086_),
    .A(net1075));
 sg13g2_nand2_2 _45933_ (.Y(_15088_),
    .A(_18509_),
    .B(_18510_));
 sg13g2_nor4_2 _45934_ (.A(\u_inv.d_reg[106] ),
    .B(_15088_),
    .C(_15086_),
    .Y(_15089_),
    .D(net1075));
 sg13g2_nor4_2 _45935_ (.A(\u_inv.d_reg[111] ),
    .B(\u_inv.d_reg[110] ),
    .C(\u_inv.d_reg[109] ),
    .Y(_15090_),
    .D(\u_inv.d_reg[108] ));
 sg13g2_nand3_1 _45936_ (.B(net1092),
    .C(_15090_),
    .A(_18507_),
    .Y(_15091_));
 sg13g2_nor4_1 _45937_ (.A(\u_inv.d_reg[115] ),
    .B(\u_inv.d_reg[114] ),
    .C(\u_inv.d_reg[113] ),
    .D(\u_inv.d_reg[112] ),
    .Y(_15092_));
 sg13g2_nand4_1 _45938_ (.B(_18507_),
    .C(_15090_),
    .A(net1092),
    .Y(_15093_),
    .D(_15092_));
 sg13g2_nand3b_1 _45939_ (.B(_18498_),
    .C(_18497_),
    .Y(_15094_),
    .A_N(net1087));
 sg13g2_nor3_2 _45940_ (.A(_15094_),
    .B(\u_inv.d_reg[118] ),
    .C(\u_inv.d_reg[119] ),
    .Y(_15095_));
 sg13g2_nor3_1 _45941_ (.A(\u_inv.d_reg[122] ),
    .B(\u_inv.d_reg[121] ),
    .C(\u_inv.d_reg[120] ),
    .Y(_15096_));
 sg13g2_nand2_1 _45942_ (.Y(_15097_),
    .A(_18491_),
    .B(_15096_));
 sg13g2_nor2_1 _45943_ (.A(\u_inv.d_reg[124] ),
    .B(_15097_),
    .Y(_15098_));
 sg13g2_nand2_1 _45944_ (.Y(_15099_),
    .A(_18488_),
    .B(_18489_));
 sg13g2_nor2_1 _45945_ (.A(\u_inv.d_reg[127] ),
    .B(_15099_),
    .Y(_15100_));
 sg13g2_nand3_1 _45946_ (.B(_15098_),
    .C(_15095_),
    .A(_15100_),
    .Y(_15101_));
 sg13g2_nand2_1 _45947_ (.Y(_15102_),
    .A(_18477_),
    .B(_18478_));
 sg13g2_nand4_1 _45948_ (.B(_18476_),
    .C(_18477_),
    .A(_18475_),
    .Y(_15103_),
    .D(_18478_));
 sg13g2_nand2b_1 _45949_ (.Y(_15104_),
    .B(_18474_),
    .A_N(_15103_));
 sg13g2_nor4_1 _45950_ (.A(\u_inv.d_reg[135] ),
    .B(\u_inv.d_reg[134] ),
    .C(\u_inv.d_reg[133] ),
    .D(\u_inv.d_reg[132] ),
    .Y(_15105_));
 sg13g2_nor3_1 _45951_ (.A(\u_inv.d_reg[143] ),
    .B(\u_inv.d_reg[142] ),
    .C(\u_inv.d_reg[131] ),
    .Y(_15106_));
 sg13g2_nand2_1 _45952_ (.Y(_15107_),
    .A(_18485_),
    .B(_18486_));
 sg13g2_nor2_1 _45953_ (.A(net7289),
    .B(_15107_),
    .Y(_15108_));
 sg13g2_nand3_1 _45954_ (.B(_15106_),
    .C(_15108_),
    .A(_15105_),
    .Y(_15109_));
 sg13g2_or4_1 _45955_ (.A(\u_inv.d_reg[141] ),
    .B(_15109_),
    .C(_15104_),
    .D(net1073),
    .X(_15110_));
 sg13g2_or3_2 _45956_ (.A(\u_inv.d_reg[147] ),
    .B(_15110_),
    .C(_15008_),
    .X(_15111_));
 sg13g2_or4_1 _45957_ (.A(\u_inv.d_reg[159] ),
    .B(_15111_),
    .C(_15006_),
    .D(\u_inv.d_reg[158] ),
    .X(_15112_));
 sg13g2_nand2_1 _45958_ (.Y(_15113_),
    .A(_18453_),
    .B(_18454_));
 sg13g2_nor2_1 _45959_ (.A(\u_inv.d_reg[162] ),
    .B(_15113_),
    .Y(_15114_));
 sg13g2_inv_1 _45960_ (.Y(_15115_),
    .A(_15114_));
 sg13g2_nor2_1 _45961_ (.A(\u_inv.d_reg[165] ),
    .B(\u_inv.d_reg[164] ),
    .Y(_15116_));
 sg13g2_nor3_1 _45962_ (.A(\u_inv.d_reg[167] ),
    .B(\u_inv.d_reg[166] ),
    .C(\u_inv.d_reg[163] ),
    .Y(_15117_));
 sg13g2_nand3_1 _45963_ (.B(_15116_),
    .C(_15117_),
    .A(_15114_),
    .Y(_15118_));
 sg13g2_or2_2 _45964_ (.X(_15119_),
    .B(_15112_),
    .A(_15118_));
 sg13g2_inv_4 _45965_ (.A(_15119_),
    .Y(_15120_));
 sg13g2_nand4_1 _45966_ (.B(_15001_),
    .C(_15002_),
    .A(_15120_),
    .Y(_15121_),
    .D(_18439_));
 sg13g2_nor4_1 _45967_ (.A(\u_inv.d_reg[179] ),
    .B(\u_inv.d_reg[178] ),
    .C(\u_inv.d_reg[177] ),
    .D(\u_inv.d_reg[176] ),
    .Y(_15122_));
 sg13g2_nand3_1 _45968_ (.B(_18434_),
    .C(_15122_),
    .A(_18433_),
    .Y(_15123_));
 sg13g2_or4_1 _45969_ (.A(\u_inv.d_reg[183] ),
    .B(\u_inv.d_reg[182] ),
    .C(_15123_),
    .D(net1085),
    .X(_15124_));
 sg13g2_nand2_1 _45970_ (.Y(_15125_),
    .A(_18429_),
    .B(_18430_));
 sg13g2_nand2b_1 _45971_ (.Y(_15126_),
    .B(_18428_),
    .A_N(_15125_));
 sg13g2_nand2b_1 _45972_ (.Y(_15127_),
    .B(_18427_),
    .A_N(_15126_));
 sg13g2_nand3b_1 _45973_ (.B(_18426_),
    .C(_18425_),
    .Y(_15128_),
    .A_N(_15127_));
 sg13g2_nor4_2 _45974_ (.A(\u_inv.d_reg[191] ),
    .B(\u_inv.d_reg[190] ),
    .C(_15128_),
    .Y(_15129_),
    .D(_15124_));
 sg13g2_nand3_1 _45975_ (.B(_18421_),
    .C(_18422_),
    .A(_18420_),
    .Y(_15130_));
 sg13g2_nor4_1 _45976_ (.A(\u_inv.d_reg[197] ),
    .B(\u_inv.d_reg[196] ),
    .C(\u_inv.d_reg[195] ),
    .D(_15130_),
    .Y(_15131_));
 sg13g2_nand2_1 _45977_ (.Y(_15132_),
    .A(_15129_),
    .B(_15131_));
 sg13g2_nand4_1 _45978_ (.B(_18416_),
    .C(_18415_),
    .A(_15129_),
    .Y(_15133_),
    .D(_15131_));
 sg13g2_nand4_1 _45979_ (.B(_18412_),
    .C(_18413_),
    .A(_18411_),
    .Y(_15134_),
    .D(_18414_));
 sg13g2_nand3b_1 _45980_ (.B(_18410_),
    .C(_18409_),
    .Y(_15135_),
    .A_N(_15134_));
 sg13g2_or4_1 _45981_ (.A(\u_inv.d_reg[207] ),
    .B(\u_inv.d_reg[206] ),
    .C(_15135_),
    .D(net1079),
    .X(_15136_));
 sg13g2_nand2_1 _45982_ (.Y(_15137_),
    .A(_18405_),
    .B(_18406_));
 sg13g2_nand4_1 _45983_ (.B(_18404_),
    .C(_18405_),
    .A(_18403_),
    .Y(_15138_),
    .D(_18406_));
 sg13g2_nand3b_1 _45984_ (.B(_18402_),
    .C(_18401_),
    .Y(_15139_),
    .A_N(_15138_));
 sg13g2_nor4_2 _45985_ (.A(\u_inv.d_reg[215] ),
    .B(\u_inv.d_reg[214] ),
    .C(_15139_),
    .Y(_15140_),
    .D(_15136_));
 sg13g2_nor3_1 _45986_ (.A(\u_inv.d_reg[218] ),
    .B(\u_inv.d_reg[217] ),
    .C(\u_inv.d_reg[216] ),
    .Y(_15141_));
 sg13g2_nand2_1 _45987_ (.Y(_15142_),
    .A(_18395_),
    .B(_15141_));
 sg13g2_nand3_1 _45988_ (.B(_18395_),
    .C(_15141_),
    .A(_18394_),
    .Y(_15143_));
 sg13g2_nor2_1 _45989_ (.A(\u_inv.d_reg[221] ),
    .B(_15143_),
    .Y(_15144_));
 sg13g2_nand4_1 _45990_ (.B(_18392_),
    .C(_18391_),
    .A(_15140_),
    .Y(_15145_),
    .D(_15144_));
 sg13g2_nand4_1 _45991_ (.B(_18388_),
    .C(_18389_),
    .A(_18387_),
    .Y(_15146_),
    .D(_18390_));
 sg13g2_nand2b_1 _45992_ (.Y(_15147_),
    .B(_18386_),
    .A_N(_15146_));
 sg13g2_nand2b_1 _45993_ (.Y(_15148_),
    .B(_18385_),
    .A_N(_15147_));
 sg13g2_nor3_1 _45994_ (.A(\u_inv.d_reg[231] ),
    .B(\u_inv.d_reg[230] ),
    .C(_15148_),
    .Y(_15149_));
 sg13g2_nand2b_1 _45995_ (.Y(_15150_),
    .B(_15149_),
    .A_N(net1069));
 sg13g2_nor4_1 _45996_ (.A(\u_inv.d_reg[235] ),
    .B(\u_inv.d_reg[234] ),
    .C(\u_inv.d_reg[233] ),
    .D(\u_inv.d_reg[232] ),
    .Y(_15151_));
 sg13g2_nand3b_1 _45997_ (.B(_15149_),
    .C(_15151_),
    .Y(_15152_),
    .A_N(net1068));
 sg13g2_nor4_1 _45998_ (.A(\u_inv.d_reg[239] ),
    .B(\u_inv.d_reg[238] ),
    .C(\u_inv.d_reg[237] ),
    .D(\u_inv.d_reg[236] ),
    .Y(_15153_));
 sg13g2_nand2b_2 _45999_ (.Y(_15154_),
    .B(_15153_),
    .A_N(net1141));
 sg13g2_nor4_1 _46000_ (.A(\u_inv.d_reg[243] ),
    .B(\u_inv.d_reg[242] ),
    .C(net7287),
    .D(net7288),
    .Y(_15155_));
 sg13g2_nand2b_1 _46001_ (.Y(_15156_),
    .B(_15155_),
    .A_N(_15154_));
 sg13g2_nand3b_1 _46002_ (.B(_18370_),
    .C(_18369_),
    .Y(_15157_),
    .A_N(_15156_));
 sg13g2_nand3b_1 _46003_ (.B(_18368_),
    .C(_18367_),
    .Y(_15158_),
    .A_N(_15157_));
 sg13g2_nand4_1 _46004_ (.B(_18364_),
    .C(_18365_),
    .A(_18363_),
    .Y(_15159_),
    .D(_18366_));
 sg13g2_nor3_2 _46005_ (.A(\u_inv.d_reg[252] ),
    .B(_15159_),
    .C(_15158_),
    .Y(_15160_));
 sg13g2_nand2_1 _46006_ (.Y(_15161_),
    .A(net7255),
    .B(_15158_));
 sg13g2_nand2_1 _46007_ (.Y(_15162_),
    .A(net7255),
    .B(_15159_));
 sg13g2_nor2_2 _46008_ (.A(_15160_),
    .B(net7163),
    .Y(_15163_));
 sg13g2_o21ai_1 _46009_ (.B1(net7258),
    .Y(_15164_),
    .A1(\u_inv.d_reg[254] ),
    .A2(\u_inv.d_reg[253] ));
 sg13g2_nor2b_2 _46010_ (.A(_15163_),
    .B_N(_15164_),
    .Y(_15165_));
 sg13g2_nand2_1 _46011_ (.Y(_15166_),
    .A(net7258),
    .B(\u_inv.d_reg[255] ));
 sg13g2_and2_2 _46012_ (.A(_15166_),
    .B(_15165_),
    .X(_15167_));
 sg13g2_xnor2_1 _46013_ (.Y(_15168_),
    .A(_15167_),
    .B(\u_inv.d_reg[256] ));
 sg13g2_xnor2_1 _46014_ (.Y(_15169_),
    .A(_18358_),
    .B(net1124));
 sg13g2_o21ai_1 _46015_ (.B1(net7255),
    .Y(_15170_),
    .A1(\u_inv.d_reg[253] ),
    .A2(net1136));
 sg13g2_xnor2_1 _46016_ (.Y(_15171_),
    .A(_18360_),
    .B(_15170_));
 sg13g2_nor3_1 _46017_ (.A(\u_inv.d_reg[249] ),
    .B(\u_inv.d_reg[248] ),
    .C(net1102),
    .Y(_15172_));
 sg13g2_nor2_1 _46018_ (.A(net7163),
    .B(_15172_),
    .Y(_15173_));
 sg13g2_xnor2_1 _46019_ (.Y(_15174_),
    .A(\u_inv.d_reg[250] ),
    .B(_15173_));
 sg13g2_xnor2_1 _46020_ (.Y(_15175_),
    .A(_18359_),
    .B(net1145));
 sg13g2_nor2_1 _46021_ (.A(_15174_),
    .B(_15175_),
    .Y(_15176_));
 sg13g2_xnor2_1 _46022_ (.Y(_15177_),
    .A(_18361_),
    .B(net1135));
 sg13g2_nand2_1 _46023_ (.Y(_15178_),
    .A(_15161_),
    .B(_15162_));
 sg13g2_xnor2_1 _46024_ (.Y(_15179_),
    .A(_18362_),
    .B(_15178_));
 sg13g2_xnor2_1 _46025_ (.Y(_15180_),
    .A(_18366_),
    .B(_15161_));
 sg13g2_nand2_1 _46026_ (.Y(_15181_),
    .A(net7253),
    .B(net1119));
 sg13g2_o21ai_1 _46027_ (.B1(net7253),
    .Y(_15182_),
    .A1(\u_inv.d_reg[246] ),
    .A2(net1120));
 sg13g2_xnor2_1 _46028_ (.Y(_15183_),
    .A(_18367_),
    .B(_15182_));
 sg13g2_and2_1 _46029_ (.A(net7253),
    .B(_15156_),
    .X(_15184_));
 sg13g2_o21ai_1 _46030_ (.B1(net7253),
    .Y(_15185_),
    .A1(\u_inv.d_reg[244] ),
    .A2(_15156_));
 sg13g2_xnor2_1 _46031_ (.Y(_15186_),
    .A(\u_inv.d_reg[245] ),
    .B(_15185_));
 sg13g2_xnor2_1 _46032_ (.Y(_15187_),
    .A(_18370_),
    .B(_15184_));
 sg13g2_nand2_1 _46033_ (.Y(_15188_),
    .A(_15186_),
    .B(_15187_));
 sg13g2_nor3_1 _46034_ (.A(net7287),
    .B(net7288),
    .C(net1118),
    .Y(_15189_));
 sg13g2_a21o_1 _46035_ (.A2(_15189_),
    .A1(_18372_),
    .B1(_18371_),
    .X(_15190_));
 sg13g2_a22oi_1 _46036_ (.Y(_15191_),
    .B1(_15184_),
    .B2(_15190_),
    .A2(\u_inv.d_reg[243] ),
    .A1(net7163));
 sg13g2_nor4_1 _46037_ (.A(_15180_),
    .B(_15183_),
    .C(_15188_),
    .D(_15191_),
    .Y(_15192_));
 sg13g2_nand4_1 _46038_ (.B(_15177_),
    .C(_15179_),
    .A(_15176_),
    .Y(_15193_),
    .D(_15192_));
 sg13g2_and2_1 _46039_ (.A(_18364_),
    .B(_15172_),
    .X(_15194_));
 sg13g2_o21ai_1 _46040_ (.B1(_15178_),
    .Y(_15195_),
    .A1(_18363_),
    .A2(_15194_));
 sg13g2_o21ai_1 _46041_ (.B1(_15195_),
    .Y(_15196_),
    .A1(net7255),
    .A2(_18363_));
 sg13g2_o21ai_1 _46042_ (.B1(net7255),
    .Y(_15197_),
    .A1(\u_inv.d_reg[248] ),
    .A2(net1105));
 sg13g2_xnor2_1 _46043_ (.Y(_15198_),
    .A(_18365_),
    .B(_15197_));
 sg13g2_inv_1 _46044_ (.Y(_15199_),
    .A(_15198_));
 sg13g2_xnor2_1 _46045_ (.Y(_15200_),
    .A(_18368_),
    .B(_15181_));
 sg13g2_nor2_1 _46046_ (.A(net7163),
    .B(_15189_),
    .Y(_15201_));
 sg13g2_xnor2_1 _46047_ (.Y(_15202_),
    .A(\u_inv.d_reg[242] ),
    .B(_15201_));
 sg13g2_nand2_1 _46048_ (.Y(_15203_),
    .A(net7253),
    .B(_15154_));
 sg13g2_nor3_1 _46049_ (.A(\u_inv.d_reg[237] ),
    .B(\u_inv.d_reg[236] ),
    .C(net1112),
    .Y(_15204_));
 sg13g2_a21oi_1 _46050_ (.A1(_18376_),
    .A2(_15204_),
    .Y(_15205_),
    .B1(_18375_));
 sg13g2_nor2_1 _46051_ (.A(_15203_),
    .B(_15205_),
    .Y(_15206_));
 sg13g2_a21oi_2 _46052_ (.B1(_15206_),
    .Y(_15207_),
    .A2(net3025),
    .A1(net7163));
 sg13g2_nand2_1 _46053_ (.Y(_15208_),
    .A(net7253),
    .B(_15152_));
 sg13g2_nor3_1 _46054_ (.A(\u_inv.d_reg[233] ),
    .B(\u_inv.d_reg[232] ),
    .C(_15150_),
    .Y(_15209_));
 sg13g2_a21oi_1 _46055_ (.A1(_18380_),
    .A2(_15209_),
    .Y(_15210_),
    .B1(_18379_));
 sg13g2_nor2_1 _46056_ (.A(_15208_),
    .B(_15210_),
    .Y(_15211_));
 sg13g2_a21oi_2 _46057_ (.B1(_15211_),
    .Y(_15212_),
    .A2(\u_inv.d_reg[235] ),
    .A1(net7163));
 sg13g2_o21ai_1 _46058_ (.B1(net7252),
    .Y(_15213_),
    .A1(\u_inv.d_reg[224] ),
    .A2(net1069));
 sg13g2_xnor2_1 _46059_ (.Y(_15214_),
    .A(_18389_),
    .B(_15213_));
 sg13g2_and2_1 _46060_ (.A(net7252),
    .B(net1069),
    .X(_15215_));
 sg13g2_xnor2_1 _46061_ (.Y(_15216_),
    .A(\u_inv.d_reg[224] ),
    .B(_15215_));
 sg13g2_nor2_1 _46062_ (.A(_15214_),
    .B(_15216_),
    .Y(_15217_));
 sg13g2_inv_1 _46063_ (.Y(_15218_),
    .A(_15217_));
 sg13g2_nor3_1 _46064_ (.A(\u_inv.d_reg[225] ),
    .B(\u_inv.d_reg[224] ),
    .C(net1069),
    .Y(_15219_));
 sg13g2_nor2_1 _46065_ (.A(net7164),
    .B(_15219_),
    .Y(_15220_));
 sg13g2_xnor2_1 _46066_ (.Y(_15221_),
    .A(\u_inv.d_reg[226] ),
    .B(_15220_));
 sg13g2_o21ai_1 _46067_ (.B1(net7252),
    .Y(_15222_),
    .A1(\u_inv.d_reg[232] ),
    .A2(_15150_));
 sg13g2_xnor2_1 _46068_ (.Y(_15223_),
    .A(_18381_),
    .B(_15222_));
 sg13g2_o21ai_1 _46069_ (.B1(net7252),
    .Y(_15224_),
    .A1(net1069),
    .A2(_15148_));
 sg13g2_inv_1 _46070_ (.Y(_15225_),
    .A(_15224_));
 sg13g2_a21oi_1 _46071_ (.A1(net7252),
    .A2(\u_inv.d_reg[230] ),
    .Y(_15226_),
    .B1(_15225_));
 sg13g2_xnor2_1 _46072_ (.Y(_15227_),
    .A(\u_inv.d_reg[231] ),
    .B(_15226_));
 sg13g2_nand2b_1 _46073_ (.Y(_15228_),
    .B(_15227_),
    .A_N(_15223_));
 sg13g2_nor4_1 _46074_ (.A(_15212_),
    .B(_15218_),
    .C(_15221_),
    .D(_15228_),
    .Y(_15229_));
 sg13g2_o21ai_1 _46075_ (.B1(net7253),
    .Y(_15230_),
    .A1(net7288),
    .A2(net1117));
 sg13g2_xnor2_1 _46076_ (.Y(_15231_),
    .A(net7287),
    .B(_15230_));
 sg13g2_nor2_1 _46077_ (.A(net7163),
    .B(_15204_),
    .Y(_15232_));
 sg13g2_xnor2_1 _46078_ (.Y(_15233_),
    .A(\u_inv.d_reg[238] ),
    .B(_15232_));
 sg13g2_inv_2 _46079_ (.Y(_15234_),
    .A(_15233_));
 sg13g2_xnor2_1 _46080_ (.Y(_15235_),
    .A(_18374_),
    .B(_15203_));
 sg13g2_nor2_1 _46081_ (.A(net7164),
    .B(_15209_),
    .Y(_15236_));
 sg13g2_xnor2_1 _46082_ (.Y(_15237_),
    .A(\u_inv.d_reg[234] ),
    .B(_15236_));
 sg13g2_o21ai_1 _46083_ (.B1(net7253),
    .Y(_15238_),
    .A1(\u_inv.d_reg[236] ),
    .A2(net1141));
 sg13g2_xnor2_1 _46084_ (.Y(_15239_),
    .A(\u_inv.d_reg[237] ),
    .B(_15238_));
 sg13g2_and2_1 _46085_ (.A(_18388_),
    .B(_15219_),
    .X(_15240_));
 sg13g2_a21o_1 _46086_ (.A2(_15146_),
    .A1(net7254),
    .B1(_15215_),
    .X(_15241_));
 sg13g2_o21ai_1 _46087_ (.B1(_15241_),
    .Y(_15242_),
    .A1(_18387_),
    .A2(_15240_));
 sg13g2_o21ai_1 _46088_ (.B1(_15242_),
    .Y(_15243_),
    .A1(net7252),
    .A2(_18387_));
 sg13g2_nand2_1 _46089_ (.Y(_15244_),
    .A(_15239_),
    .B(_15243_));
 sg13g2_nand2_1 _46090_ (.Y(_15245_),
    .A(net7260),
    .B(_15132_));
 sg13g2_o21ai_1 _46091_ (.B1(net7260),
    .Y(_15246_),
    .A1(\u_inv.d_reg[198] ),
    .A2(_15132_));
 sg13g2_xnor2_1 _46092_ (.Y(_15247_),
    .A(\u_inv.d_reg[199] ),
    .B(_15246_));
 sg13g2_o21ai_1 _46093_ (.B1(net7265),
    .Y(_15248_),
    .A1(\u_inv.d_reg[176] ),
    .A2(net1085));
 sg13g2_xnor2_1 _46094_ (.Y(_15249_),
    .A(_18437_),
    .B(_15248_));
 sg13g2_nand2_1 _46095_ (.Y(_15250_),
    .A(net7262),
    .B(net1085));
 sg13g2_xnor2_1 _46096_ (.Y(_15251_),
    .A(_18438_),
    .B(_15250_));
 sg13g2_or2_1 _46097_ (.X(_15252_),
    .B(_15251_),
    .A(_15249_));
 sg13g2_and2_1 _46098_ (.A(net7261),
    .B(_15124_),
    .X(_15253_));
 sg13g2_a21o_1 _46099_ (.A2(_15128_),
    .A1(net7261),
    .B1(_15253_),
    .X(_15254_));
 sg13g2_xnor2_1 _46100_ (.Y(_15255_),
    .A(\u_inv.d_reg[190] ),
    .B(_15254_));
 sg13g2_nor2_2 _46101_ (.A(net7165),
    .B(_15129_),
    .Y(_15256_));
 sg13g2_xnor2_1 _46102_ (.Y(_15257_),
    .A(_18422_),
    .B(_15256_));
 sg13g2_xnor2_1 _46103_ (.Y(_15258_),
    .A(\u_inv.d_reg[192] ),
    .B(_15256_));
 sg13g2_nor3_1 _46104_ (.A(\u_inv.d_reg[177] ),
    .B(\u_inv.d_reg[176] ),
    .C(net1085),
    .Y(_15259_));
 sg13g2_nor2_1 _46105_ (.A(net7165),
    .B(_15259_),
    .Y(_15260_));
 sg13g2_xnor2_1 _46106_ (.Y(_15261_),
    .A(\u_inv.d_reg[178] ),
    .B(_15260_));
 sg13g2_nor4_1 _46107_ (.A(_15252_),
    .B(_15255_),
    .C(_15258_),
    .D(_15261_),
    .Y(_15262_));
 sg13g2_a21oi_1 _46108_ (.A1(net7260),
    .A2(_15130_),
    .Y(_15263_),
    .B1(_15256_));
 sg13g2_a21o_1 _46109_ (.A2(_15263_),
    .A1(_18419_),
    .B1(net7165),
    .X(_15264_));
 sg13g2_o21ai_1 _46110_ (.B1(_15264_),
    .Y(_15265_),
    .A1(net7165),
    .A2(_18418_));
 sg13g2_xnor2_1 _46111_ (.Y(_15266_),
    .A(_18417_),
    .B(_15265_));
 sg13g2_or4_1 _46112_ (.A(\u_inv.d_reg[150] ),
    .B(\u_inv.d_reg[149] ),
    .C(\u_inv.d_reg[148] ),
    .D(_15111_),
    .X(_15267_));
 sg13g2_nand2_1 _46113_ (.Y(_15268_),
    .A(net7271),
    .B(_15267_));
 sg13g2_o21ai_1 _46114_ (.B1(net7271),
    .Y(_15269_),
    .A1(\u_inv.d_reg[151] ),
    .A2(_15267_));
 sg13g2_o21ai_1 _46115_ (.B1(net7271),
    .Y(_15270_),
    .A1(\u_inv.d_reg[153] ),
    .A2(\u_inv.d_reg[152] ));
 sg13g2_and2_1 _46116_ (.A(_15269_),
    .B(_15270_),
    .X(_15271_));
 sg13g2_o21ai_1 _46117_ (.B1(net7271),
    .Y(_15272_),
    .A1(\u_inv.d_reg[155] ),
    .A2(\u_inv.d_reg[154] ));
 sg13g2_nand2_1 _46118_ (.Y(_15273_),
    .A(_15271_),
    .B(_15272_));
 sg13g2_o21ai_1 _46119_ (.B1(net7271),
    .Y(_15274_),
    .A1(\u_inv.d_reg[156] ),
    .A2(_15273_));
 sg13g2_xnor2_1 _46120_ (.Y(_15275_),
    .A(net3762),
    .B(_15274_));
 sg13g2_xnor2_1 _46121_ (.Y(_15276_),
    .A(_18457_),
    .B(_15274_));
 sg13g2_and2_1 _46122_ (.A(net7271),
    .B(_15111_),
    .X(_15277_));
 sg13g2_o21ai_1 _46123_ (.B1(net7267),
    .Y(_15278_),
    .A1(_15006_),
    .A2(_15111_));
 sg13g2_xnor2_1 _46124_ (.Y(_15279_),
    .A(_18456_),
    .B(_15278_));
 sg13g2_xnor2_1 _46125_ (.Y(_15280_),
    .A(\u_inv.d_reg[156] ),
    .B(_15273_));
 sg13g2_nor3_2 _46126_ (.A(_15276_),
    .B(_15279_),
    .C(_15280_),
    .Y(_15281_));
 sg13g2_nand4_1 _46127_ (.B(_15262_),
    .C(_15266_),
    .A(_15247_),
    .Y(_15282_),
    .D(_15281_));
 sg13g2_a21o_1 _46128_ (.A2(_15127_),
    .A1(net7261),
    .B1(_15253_),
    .X(_15283_));
 sg13g2_a21o_1 _46129_ (.A2(\u_inv.d_reg[188] ),
    .A1(net7261),
    .B1(_15283_),
    .X(_15284_));
 sg13g2_xnor2_1 _46130_ (.Y(_15285_),
    .A(_18425_),
    .B(_15284_));
 sg13g2_xnor2_1 _46131_ (.Y(_15286_),
    .A(net2932),
    .B(_15283_));
 sg13g2_nand2b_2 _46132_ (.Y(_15287_),
    .B(_15285_),
    .A_N(_15286_));
 sg13g2_nand2_1 _46133_ (.Y(_15288_),
    .A(net7266),
    .B(_15112_));
 sg13g2_o21ai_1 _46134_ (.B1(net7266),
    .Y(_15289_),
    .A1(_15112_),
    .A2(_15115_));
 sg13g2_nand3b_1 _46135_ (.B(_15114_),
    .C(_18451_),
    .Y(_15290_),
    .A_N(_15112_));
 sg13g2_nand2_1 _46136_ (.Y(_15291_),
    .A(net7266),
    .B(_15290_));
 sg13g2_xnor2_1 _46137_ (.Y(_15292_),
    .A(\u_inv.d_reg[164] ),
    .B(_15291_));
 sg13g2_o21ai_1 _46138_ (.B1(net7266),
    .Y(_15293_),
    .A1(\u_inv.d_reg[164] ),
    .A2(_15290_));
 sg13g2_xnor2_1 _46139_ (.Y(_15294_),
    .A(\u_inv.d_reg[165] ),
    .B(_15293_));
 sg13g2_nand2_2 _46140_ (.Y(_15295_),
    .A(_15292_),
    .B(_15294_));
 sg13g2_xnor2_1 _46141_ (.Y(_15296_),
    .A(net3768),
    .B(_15263_));
 sg13g2_inv_2 _46142_ (.Y(_15297_),
    .A(_15296_));
 sg13g2_a21oi_1 _46143_ (.A1(net7261),
    .A2(\u_inv.d_reg[190] ),
    .Y(_15298_),
    .B1(_15254_));
 sg13g2_xnor2_1 _46144_ (.Y(_15299_),
    .A(_18423_),
    .B(_15298_));
 sg13g2_nor4_2 _46145_ (.A(_15287_),
    .B(_15295_),
    .C(_15297_),
    .Y(_15300_),
    .D(_15299_));
 sg13g2_o21ai_1 _46146_ (.B1(net7267),
    .Y(_15301_),
    .A1(_15000_),
    .A2(net1126));
 sg13g2_xnor2_1 _46147_ (.Y(_15302_),
    .A(\u_inv.d_reg[170] ),
    .B(_15301_));
 sg13g2_nand2b_1 _46148_ (.Y(_15303_),
    .B(_15108_),
    .A_N(net1073));
 sg13g2_nor2_2 _46149_ (.A(\u_inv.d_reg[131] ),
    .B(_15303_),
    .Y(_15304_));
 sg13g2_nand2_2 _46150_ (.Y(_15305_),
    .A(_15105_),
    .B(_15304_));
 sg13g2_nor3_1 _46151_ (.A(\u_inv.d_reg[141] ),
    .B(_15104_),
    .C(_15305_),
    .Y(_15306_));
 sg13g2_nand2b_1 _46152_ (.Y(_15307_),
    .B(net7269),
    .A_N(_15306_));
 sg13g2_a21oi_1 _46153_ (.A1(_18472_),
    .A2(_15306_),
    .Y(_15308_),
    .B1(net7171));
 sg13g2_xnor2_1 _46154_ (.Y(_15309_),
    .A(\u_inv.d_reg[143] ),
    .B(_15308_));
 sg13g2_inv_4 _46155_ (.A(_15309_),
    .Y(_15310_));
 sg13g2_nand2_1 _46156_ (.Y(_15311_),
    .A(net7266),
    .B(_15119_));
 sg13g2_o21ai_1 _46157_ (.B1(net7267),
    .Y(_15312_),
    .A1(_15003_),
    .A2(net1127));
 sg13g2_xnor2_1 _46158_ (.Y(_15313_),
    .A(\u_inv.d_reg[175] ),
    .B(_15312_));
 sg13g2_a21oi_2 _46159_ (.B1(net7167),
    .Y(_15314_),
    .A2(_15120_),
    .A1(_15001_));
 sg13g2_xnor2_1 _46160_ (.Y(_15315_),
    .A(_18442_),
    .B(_15314_));
 sg13g2_nand4_1 _46161_ (.B(_15310_),
    .C(_15313_),
    .A(_15302_),
    .Y(_15316_),
    .D(_15315_));
 sg13g2_nand2_1 _46162_ (.Y(_15317_),
    .A(net7269),
    .B(_15110_));
 sg13g2_o21ai_1 _46163_ (.B1(net7269),
    .Y(_15318_),
    .A1(\u_inv.d_reg[144] ),
    .A2(_15110_));
 sg13g2_xnor2_1 _46164_ (.Y(_15319_),
    .A(_18469_),
    .B(_15318_));
 sg13g2_inv_1 _46165_ (.Y(_15320_),
    .A(_15319_));
 sg13g2_xnor2_1 _46166_ (.Y(_15321_),
    .A(\u_inv.d_reg[148] ),
    .B(_15277_));
 sg13g2_o21ai_1 _46167_ (.B1(net7269),
    .Y(_15322_),
    .A1(_15008_),
    .A2(net1129));
 sg13g2_xnor2_1 _46168_ (.Y(_15323_),
    .A(\u_inv.d_reg[147] ),
    .B(_15322_));
 sg13g2_inv_1 _46169_ (.Y(_15324_),
    .A(_15323_));
 sg13g2_nor2_1 _46170_ (.A(net7170),
    .B(_15304_),
    .Y(_15325_));
 sg13g2_xnor2_1 _46171_ (.Y(_15326_),
    .A(\u_inv.d_reg[132] ),
    .B(_15325_));
 sg13g2_nor2_2 _46172_ (.A(net7174),
    .B(net1110),
    .Y(_15327_));
 sg13g2_o21ai_1 _46173_ (.B1(net7278),
    .Y(_15328_),
    .A1(\u_inv.d_reg[121] ),
    .A2(\u_inv.d_reg[120] ));
 sg13g2_nor2b_1 _46174_ (.A(_15327_),
    .B_N(_15328_),
    .Y(_15329_));
 sg13g2_xnor2_1 _46175_ (.Y(_15330_),
    .A(_18492_),
    .B(_15329_));
 sg13g2_and2_1 _46176_ (.A(net7278),
    .B(net1073),
    .X(_15331_));
 sg13g2_xnor2_1 _46177_ (.Y(_15332_),
    .A(\u_inv.d_reg[128] ),
    .B(_15331_));
 sg13g2_a21oi_1 _46178_ (.A1(_15095_),
    .A2(_15096_),
    .Y(_15333_),
    .B1(net7174));
 sg13g2_xnor2_1 _46179_ (.Y(_15334_),
    .A(net3764),
    .B(_15333_));
 sg13g2_a21oi_1 _46180_ (.A1(net7278),
    .A2(_15097_),
    .Y(_15335_),
    .B1(_15327_));
 sg13g2_xnor2_1 _46181_ (.Y(_15336_),
    .A(\u_inv.d_reg[124] ),
    .B(_15335_));
 sg13g2_nand2b_2 _46182_ (.Y(_15337_),
    .B(_15336_),
    .A_N(_15334_));
 sg13g2_nor4_1 _46183_ (.A(_15326_),
    .B(_15330_),
    .C(_15332_),
    .D(_15337_),
    .Y(_15338_));
 sg13g2_nand2_1 _46184_ (.Y(_15339_),
    .A(net7275),
    .B(_15303_));
 sg13g2_xnor2_1 _46185_ (.Y(_15340_),
    .A(_18483_),
    .B(_15339_));
 sg13g2_xnor2_1 _46186_ (.Y(_15341_),
    .A(\u_inv.d_reg[131] ),
    .B(_15339_));
 sg13g2_o21ai_1 _46187_ (.B1(net7275),
    .Y(_15342_),
    .A1(net1073),
    .A2(_15107_));
 sg13g2_xnor2_1 _46188_ (.Y(_15343_),
    .A(net7289),
    .B(_15342_));
 sg13g2_inv_1 _46189_ (.Y(_15344_),
    .A(_15343_));
 sg13g2_o21ai_1 _46190_ (.B1(net7269),
    .Y(_15345_),
    .A1(_15007_),
    .A2(net1128));
 sg13g2_xnor2_1 _46191_ (.Y(_15346_),
    .A(\u_inv.d_reg[146] ),
    .B(_15345_));
 sg13g2_nand4_1 _46192_ (.B(_15341_),
    .C(_15343_),
    .A(_15338_),
    .Y(_15347_),
    .D(_15346_));
 sg13g2_nor4_2 _46193_ (.A(_15319_),
    .B(_15321_),
    .C(_15324_),
    .Y(_15348_),
    .D(_15347_));
 sg13g2_xnor2_1 _46194_ (.Y(_15349_),
    .A(\u_inv.d_reg[163] ),
    .B(_15289_));
 sg13g2_o21ai_1 _46195_ (.B1(net7269),
    .Y(_15350_),
    .A1(_15104_),
    .A2(_15305_));
 sg13g2_xnor2_1 _46196_ (.Y(_15351_),
    .A(\u_inv.d_reg[141] ),
    .B(_15350_));
 sg13g2_nand3_1 _46197_ (.B(_15349_),
    .C(_15351_),
    .A(_15348_),
    .Y(_15352_));
 sg13g2_a21oi_1 _46198_ (.A1(_18482_),
    .A2(_15304_),
    .Y(_15353_),
    .B1(net7170));
 sg13g2_xnor2_1 _46199_ (.Y(_15354_),
    .A(_18481_),
    .B(_15353_));
 sg13g2_xnor2_1 _46200_ (.Y(_15355_),
    .A(\u_inv.d_reg[133] ),
    .B(_15353_));
 sg13g2_xnor2_1 _46201_ (.Y(_15356_),
    .A(_18463_),
    .B(_15268_));
 sg13g2_o21ai_1 _46202_ (.B1(net7275),
    .Y(_15357_),
    .A1(\u_inv.d_reg[133] ),
    .A2(\u_inv.d_reg[132] ));
 sg13g2_nor2b_1 _46203_ (.A(_15325_),
    .B_N(_15357_),
    .Y(_15358_));
 sg13g2_inv_1 _46204_ (.Y(_15359_),
    .A(_15358_));
 sg13g2_a21oi_1 _46205_ (.A1(net7275),
    .A2(\u_inv.d_reg[134] ),
    .Y(_15360_),
    .B1(_15359_));
 sg13g2_xnor2_1 _46206_ (.Y(_15361_),
    .A(\u_inv.d_reg[135] ),
    .B(_15360_));
 sg13g2_o21ai_1 _46207_ (.B1(net7271),
    .Y(_15362_),
    .A1(\u_inv.d_reg[148] ),
    .A2(_15111_));
 sg13g2_inv_1 _46208_ (.Y(_15363_),
    .A(_15362_));
 sg13g2_xnor2_1 _46209_ (.Y(_15364_),
    .A(\u_inv.d_reg[149] ),
    .B(_15362_));
 sg13g2_nand2_1 _46210_ (.Y(_15365_),
    .A(_15361_),
    .B(_15364_));
 sg13g2_nor3_1 _46211_ (.A(_15355_),
    .B(_15356_),
    .C(_15365_),
    .Y(_15366_));
 sg13g2_o21ai_1 _46212_ (.B1(net7278),
    .Y(_15367_),
    .A1(\u_inv.d_reg[128] ),
    .A2(net1073));
 sg13g2_xnor2_1 _46213_ (.Y(_15368_),
    .A(_18485_),
    .B(_15367_));
 sg13g2_a21oi_1 _46214_ (.A1(_15095_),
    .A2(_15098_),
    .Y(_15369_),
    .B1(net7174));
 sg13g2_a21oi_1 _46215_ (.A1(net7278),
    .A2(\u_inv.d_reg[125] ),
    .Y(_15370_),
    .B1(_15369_));
 sg13g2_xnor2_1 _46216_ (.Y(_15371_),
    .A(\u_inv.d_reg[126] ),
    .B(_15370_));
 sg13g2_a21oi_1 _46217_ (.A1(net7278),
    .A2(_15099_),
    .Y(_15372_),
    .B1(_15369_));
 sg13g2_xnor2_1 _46218_ (.Y(_15373_),
    .A(\u_inv.d_reg[127] ),
    .B(_15372_));
 sg13g2_nand2_1 _46219_ (.Y(_15374_),
    .A(_15371_),
    .B(_15373_));
 sg13g2_nand2_1 _46220_ (.Y(_15375_),
    .A(net7276),
    .B(net1122));
 sg13g2_o21ai_1 _46221_ (.B1(net7277),
    .Y(_15376_),
    .A1(\u_inv.d_reg[118] ),
    .A2(net1122));
 sg13g2_xnor2_1 _46222_ (.Y(_15377_),
    .A(_18495_),
    .B(_15376_));
 sg13g2_nand2_1 _46223_ (.Y(_15378_),
    .A(net7276),
    .B(net1087));
 sg13g2_o21ai_1 _46224_ (.B1(net7276),
    .Y(_15379_),
    .A1(\u_inv.d_reg[116] ),
    .A2(net1133));
 sg13g2_xnor2_1 _46225_ (.Y(_15380_),
    .A(_18497_),
    .B(_15379_));
 sg13g2_xnor2_1 _46226_ (.Y(_15381_),
    .A(_18498_),
    .B(_15378_));
 sg13g2_a21o_2 _46227_ (.A2(net1092),
    .A1(_18507_),
    .B1(net7173),
    .X(_15382_));
 sg13g2_nand2_1 _46228_ (.Y(_15383_),
    .A(net7284),
    .B(\u_inv.d_reg[108] ));
 sg13g2_nand2_1 _46229_ (.Y(_15384_),
    .A(_15382_),
    .B(_15383_));
 sg13g2_xnor2_1 _46230_ (.Y(_15385_),
    .A(_18505_),
    .B(_15384_));
 sg13g2_xnor2_1 _46231_ (.Y(_15386_),
    .A(_18506_),
    .B(_15382_));
 sg13g2_nor2_1 _46232_ (.A(net7173),
    .B(net1092),
    .Y(_15387_));
 sg13g2_xnor2_1 _46233_ (.Y(_15388_),
    .A(_18507_),
    .B(_15387_));
 sg13g2_nand2_1 _46234_ (.Y(_15389_),
    .A(net7284),
    .B(net1075));
 sg13g2_o21ai_1 _46235_ (.B1(net7284),
    .Y(_15390_),
    .A1(\u_inv.d_reg[102] ),
    .A2(net1075));
 sg13g2_xnor2_1 _46236_ (.Y(_15391_),
    .A(\u_inv.d_reg[103] ),
    .B(_15390_));
 sg13g2_nand2_1 _46237_ (.Y(_15392_),
    .A(net7276),
    .B(_15083_));
 sg13g2_xnor2_1 _46238_ (.Y(_15393_),
    .A(\u_inv.d_reg[100] ),
    .B(_15392_));
 sg13g2_o21ai_1 _46239_ (.B1(net7276),
    .Y(_15394_),
    .A1(\u_inv.d_reg[100] ),
    .A2(_15083_));
 sg13g2_xnor2_1 _46240_ (.Y(_15395_),
    .A(\u_inv.d_reg[101] ),
    .B(_15394_));
 sg13g2_nand2_2 _46241_ (.Y(_15396_),
    .A(net7283),
    .B(_15087_));
 sg13g2_xnor2_1 _46242_ (.Y(_15397_),
    .A(\u_inv.d_reg[104] ),
    .B(_15396_));
 sg13g2_xnor2_1 _46243_ (.Y(_15398_),
    .A(_18510_),
    .B(_15396_));
 sg13g2_nor2_1 _46244_ (.A(net7174),
    .B(net1103),
    .Y(_15399_));
 sg13g2_a21oi_1 _46245_ (.A1(net7276),
    .A2(\u_inv.d_reg[92] ),
    .Y(_15400_),
    .B1(_15399_));
 sg13g2_o21ai_1 _46246_ (.B1(net7276),
    .Y(_15401_),
    .A1(\u_inv.d_reg[94] ),
    .A2(\u_inv.d_reg[93] ));
 sg13g2_nand2_1 _46247_ (.Y(_15402_),
    .A(_15400_),
    .B(_15401_));
 sg13g2_xnor2_1 _46248_ (.Y(_15403_),
    .A(_18519_),
    .B(_15402_));
 sg13g2_a21oi_1 _46249_ (.A1(_15079_),
    .A2(_15080_),
    .Y(_15404_),
    .B1(net7173));
 sg13g2_a21oi_1 _46250_ (.A1(net7283),
    .A2(_15081_),
    .Y(_15405_),
    .B1(_15404_));
 sg13g2_inv_1 _46251_ (.Y(_15406_),
    .A(_15405_));
 sg13g2_xnor2_1 _46252_ (.Y(_15407_),
    .A(\u_inv.d_reg[98] ),
    .B(_15405_));
 sg13g2_a21oi_1 _46253_ (.A1(net7283),
    .A2(\u_inv.d_reg[96] ),
    .Y(_15408_),
    .B1(_15404_));
 sg13g2_xnor2_1 _46254_ (.Y(_15409_),
    .A(\u_inv.d_reg[97] ),
    .B(_15408_));
 sg13g2_xnor2_1 _46255_ (.Y(_15410_),
    .A(_18517_),
    .B(_15408_));
 sg13g2_nand4_1 _46256_ (.B(_15403_),
    .C(_15407_),
    .A(_15397_),
    .Y(_15411_),
    .D(_15409_));
 sg13g2_nor2b_1 _46257_ (.A(_15411_),
    .B_N(_15388_),
    .Y(_15412_));
 sg13g2_nand4_1 _46258_ (.B(_15393_),
    .C(_15395_),
    .A(_15391_),
    .Y(_15413_),
    .D(_15412_));
 sg13g2_o21ai_1 _46259_ (.B1(net7283),
    .Y(_15414_),
    .A1(_15087_),
    .A2(_15088_));
 sg13g2_xnor2_1 _46260_ (.Y(_15415_),
    .A(_18508_),
    .B(_15414_));
 sg13g2_inv_2 _46261_ (.Y(_15416_),
    .A(_15415_));
 sg13g2_o21ai_1 _46262_ (.B1(_15396_),
    .Y(_15417_),
    .A1(net7173),
    .A2(_18510_));
 sg13g2_xnor2_1 _46263_ (.Y(_15418_),
    .A(\u_inv.d_reg[105] ),
    .B(_15417_));
 sg13g2_inv_1 _46264_ (.Y(_15419_),
    .A(_15418_));
 sg13g2_a21o_1 _46265_ (.A2(_15400_),
    .A1(_18521_),
    .B1(net7174),
    .X(_15420_));
 sg13g2_xnor2_1 _46266_ (.Y(_15421_),
    .A(_18520_),
    .B(_15420_));
 sg13g2_xnor2_1 _46267_ (.Y(_15422_),
    .A(_18522_),
    .B(_15399_));
 sg13g2_o21ai_1 _46268_ (.B1(net7277),
    .Y(_15423_),
    .A1(\u_inv.d_reg[90] ),
    .A2(_15078_));
 sg13g2_xnor2_1 _46269_ (.Y(_15424_),
    .A(_18523_),
    .B(_15423_));
 sg13g2_nand2_1 _46270_ (.Y(_15425_),
    .A(net7282),
    .B(net1082));
 sg13g2_xnor2_1 _46271_ (.Y(_15426_),
    .A(\u_inv.d_reg[88] ),
    .B(_15425_));
 sg13g2_inv_1 _46272_ (.Y(_15427_),
    .A(_15426_));
 sg13g2_o21ai_1 _46273_ (.B1(net7282),
    .Y(_15428_),
    .A1(\u_inv.d_reg[86] ),
    .A2(_15074_));
 sg13g2_xnor2_1 _46274_ (.Y(_15429_),
    .A(net3766),
    .B(_15428_));
 sg13g2_nand2_1 _46275_ (.Y(_15430_),
    .A(net7282),
    .B(_15074_));
 sg13g2_xnor2_1 _46276_ (.Y(_15431_),
    .A(_18528_),
    .B(_15430_));
 sg13g2_o21ai_1 _46277_ (.B1(net7282),
    .Y(_15432_),
    .A1(\u_inv.d_reg[84] ),
    .A2(_15072_));
 sg13g2_xnor2_1 _46278_ (.Y(_15433_),
    .A(_18529_),
    .B(_15432_));
 sg13g2_nand2_1 _46279_ (.Y(_15434_),
    .A(net7282),
    .B(_15072_));
 sg13g2_xnor2_1 _46280_ (.Y(_15435_),
    .A(_18530_),
    .B(_15434_));
 sg13g2_nor2_1 _46281_ (.A(_15433_),
    .B(_15435_),
    .Y(_15436_));
 sg13g2_inv_1 _46282_ (.Y(_15437_),
    .A(_15436_));
 sg13g2_nor2_1 _46283_ (.A(net7172),
    .B(net1095),
    .Y(_15438_));
 sg13g2_o21ai_1 _46284_ (.B1(net7282),
    .Y(_15439_),
    .A1(\u_inv.d_reg[82] ),
    .A2(net7290));
 sg13g2_nor2b_1 _46285_ (.A(_15438_),
    .B_N(_15439_),
    .Y(_15440_));
 sg13g2_xnor2_1 _46286_ (.Y(_15441_),
    .A(\u_inv.d_reg[83] ),
    .B(_15440_));
 sg13g2_a21oi_1 _46287_ (.A1(net7281),
    .A2(net7290),
    .Y(_15442_),
    .B1(_15438_));
 sg13g2_xnor2_1 _46288_ (.Y(_15443_),
    .A(_18532_),
    .B(_15442_));
 sg13g2_inv_1 _46289_ (.Y(_15444_),
    .A(_15443_));
 sg13g2_nand2_1 _46290_ (.Y(_15445_),
    .A(_15441_),
    .B(_15444_));
 sg13g2_nor2_1 _46291_ (.A(net7172),
    .B(_15069_),
    .Y(_15446_));
 sg13g2_xnor2_1 _46292_ (.Y(_15447_),
    .A(_18534_),
    .B(_15446_));
 sg13g2_inv_1 _46293_ (.Y(_15448_),
    .A(_15447_));
 sg13g2_nor2_1 _46294_ (.A(net7172),
    .B(_15066_),
    .Y(_15449_));
 sg13g2_a21oi_1 _46295_ (.A1(_18537_),
    .A2(_15066_),
    .Y(_15450_),
    .B1(net7172));
 sg13g2_xnor2_1 _46296_ (.Y(_15451_),
    .A(\u_inv.d_reg[78] ),
    .B(_15450_));
 sg13g2_a21oi_1 _46297_ (.A1(_15066_),
    .A2(_15067_),
    .Y(_15452_),
    .B1(net7172));
 sg13g2_xnor2_1 _46298_ (.Y(_15453_),
    .A(\u_inv.d_reg[79] ),
    .B(_15452_));
 sg13g2_nor3_1 _46299_ (.A(_15448_),
    .B(_15451_),
    .C(_15453_),
    .Y(_15454_));
 sg13g2_xnor2_1 _46300_ (.Y(_15455_),
    .A(_18533_),
    .B(_15438_));
 sg13g2_xnor2_1 _46301_ (.Y(_15456_),
    .A(_18537_),
    .B(_15449_));
 sg13g2_nand2_1 _46302_ (.Y(_15457_),
    .A(net7280),
    .B(_15065_));
 sg13g2_xnor2_1 _46303_ (.Y(_15458_),
    .A(_18538_),
    .B(_15457_));
 sg13g2_inv_1 _46304_ (.Y(_15459_),
    .A(_15458_));
 sg13g2_nand2_1 _46305_ (.Y(_15460_),
    .A(net7280),
    .B(_15064_));
 sg13g2_xnor2_1 _46306_ (.Y(_15461_),
    .A(_18539_),
    .B(_15460_));
 sg13g2_inv_1 _46307_ (.Y(_15462_),
    .A(_15461_));
 sg13g2_o21ai_1 _46308_ (.B1(net7280),
    .Y(_15463_),
    .A1(_15062_),
    .A2(_15063_));
 sg13g2_xnor2_1 _46309_ (.Y(_15464_),
    .A(_18540_),
    .B(_15463_));
 sg13g2_o21ai_1 _46310_ (.B1(net7280),
    .Y(_15465_),
    .A1(\u_inv.d_reg[72] ),
    .A2(_15062_));
 sg13g2_xnor2_1 _46311_ (.Y(_15466_),
    .A(_18541_),
    .B(_15465_));
 sg13g2_nand2_1 _46312_ (.Y(_15467_),
    .A(net7280),
    .B(_15062_));
 sg13g2_xnor2_1 _46313_ (.Y(_15468_),
    .A(_18542_),
    .B(_15467_));
 sg13g2_o21ai_1 _46314_ (.B1(net7281),
    .Y(_15469_),
    .A1(\u_inv.d_reg[70] ),
    .A2(net1100));
 sg13g2_xnor2_1 _46315_ (.Y(_15470_),
    .A(_18543_),
    .B(_15469_));
 sg13g2_nand2_1 _46316_ (.Y(_15471_),
    .A(net7280),
    .B(net1100));
 sg13g2_xnor2_1 _46317_ (.Y(_15472_),
    .A(_18544_),
    .B(_15471_));
 sg13g2_inv_2 _46318_ (.Y(_15473_),
    .A(_15472_));
 sg13g2_o21ai_1 _46319_ (.B1(net7280),
    .Y(_15474_),
    .A1(\u_inv.d_reg[68] ),
    .A2(_15058_));
 sg13g2_xnor2_1 _46320_ (.Y(_15475_),
    .A(\u_inv.d_reg[69] ),
    .B(_15474_));
 sg13g2_nand2_1 _46321_ (.Y(_15476_),
    .A(net7280),
    .B(_15058_));
 sg13g2_xnor2_1 _46322_ (.Y(_15477_),
    .A(_18546_),
    .B(_15476_));
 sg13g2_inv_1 _46323_ (.Y(_15478_),
    .A(_15477_));
 sg13g2_nor2_1 _46324_ (.A(net7172),
    .B(_15056_),
    .Y(_15479_));
 sg13g2_xnor2_1 _46325_ (.Y(_15480_),
    .A(\u_inv.d_reg[67] ),
    .B(_15479_));
 sg13g2_a21oi_1 _46326_ (.A1(net1072),
    .A2(_15053_),
    .Y(_15481_),
    .B1(net7172));
 sg13g2_xnor2_1 _46327_ (.Y(_15482_),
    .A(\u_inv.d_reg[64] ),
    .B(_15481_));
 sg13g2_a21oi_1 _46328_ (.A1(_18552_),
    .A2(net1072),
    .Y(_15483_),
    .B1(net7174));
 sg13g2_xnor2_1 _46329_ (.Y(_15484_),
    .A(\u_inv.d_reg[63] ),
    .B(_15483_));
 sg13g2_nor2_1 _46330_ (.A(net7174),
    .B(net1072),
    .Y(_15485_));
 sg13g2_xnor2_1 _46331_ (.Y(_15486_),
    .A(\u_inv.d_reg[62] ),
    .B(_15485_));
 sg13g2_nor2_1 _46332_ (.A(net7174),
    .B(_15051_),
    .Y(_15487_));
 sg13g2_xnor2_1 _46333_ (.Y(_15488_),
    .A(\u_inv.d_reg[61] ),
    .B(_15487_));
 sg13g2_o21ai_1 _46334_ (.B1(net7279),
    .Y(_15489_),
    .A1(\u_inv.d_reg[59] ),
    .A2(net1084));
 sg13g2_xnor2_1 _46335_ (.Y(_15490_),
    .A(_18554_),
    .B(_15489_));
 sg13g2_nand2_1 _46336_ (.Y(_15491_),
    .A(net7279),
    .B(net1084));
 sg13g2_xnor2_1 _46337_ (.Y(_15492_),
    .A(_18555_),
    .B(_15491_));
 sg13g2_nand2_1 _46338_ (.Y(_15493_),
    .A(net7279),
    .B(_15049_));
 sg13g2_xnor2_1 _46339_ (.Y(_15494_),
    .A(_18556_),
    .B(_15493_));
 sg13g2_inv_1 _46340_ (.Y(_15495_),
    .A(_15494_));
 sg13g2_o21ai_1 _46341_ (.B1(net7279),
    .Y(_15496_),
    .A1(\u_inv.d_reg[56] ),
    .A2(_15047_));
 sg13g2_xnor2_1 _46342_ (.Y(_15497_),
    .A(\u_inv.d_reg[57] ),
    .B(_15496_));
 sg13g2_a21oi_1 _46343_ (.A1(net1089),
    .A2(_15046_),
    .Y(_15498_),
    .B1(net7169));
 sg13g2_xnor2_1 _46344_ (.Y(_15499_),
    .A(_18558_),
    .B(_15498_));
 sg13g2_xnor2_1 _46345_ (.Y(_15500_),
    .A(\u_inv.d_reg[56] ),
    .B(_15498_));
 sg13g2_a21oi_1 _46346_ (.A1(_18560_),
    .A2(net1088),
    .Y(_15501_),
    .B1(net7169));
 sg13g2_xnor2_1 _46347_ (.Y(_15502_),
    .A(net2775),
    .B(_15501_));
 sg13g2_nor2_1 _46348_ (.A(net7169),
    .B(_15045_),
    .Y(_15503_));
 sg13g2_xnor2_1 _46349_ (.Y(_15504_),
    .A(\u_inv.d_reg[54] ),
    .B(_15503_));
 sg13g2_nor2_1 _46350_ (.A(net7170),
    .B(_15044_),
    .Y(_15505_));
 sg13g2_xnor2_1 _46351_ (.Y(_15506_),
    .A(\u_inv.d_reg[53] ),
    .B(_15505_));
 sg13g2_o21ai_1 _46352_ (.B1(net7274),
    .Y(_15507_),
    .A1(\u_inv.d_reg[51] ),
    .A2(net1091));
 sg13g2_xnor2_1 _46353_ (.Y(_15508_),
    .A(_18562_),
    .B(_15507_));
 sg13g2_nand2_1 _46354_ (.Y(_15509_),
    .A(net7274),
    .B(net1091));
 sg13g2_xnor2_1 _46355_ (.Y(_15510_),
    .A(_18563_),
    .B(_15509_));
 sg13g2_nand2_1 _46356_ (.Y(_15511_),
    .A(net7274),
    .B(_15042_));
 sg13g2_xnor2_1 _46357_ (.Y(_15512_),
    .A(_18564_),
    .B(_15511_));
 sg13g2_a21o_1 _46358_ (.A2(_15038_),
    .A1(_18570_),
    .B1(net7169),
    .X(_15513_));
 sg13g2_o21ai_1 _46359_ (.B1(net7274),
    .Y(_15514_),
    .A1(\u_inv.d_reg[46] ),
    .A2(\u_inv.d_reg[45] ));
 sg13g2_nand2_1 _46360_ (.Y(_15515_),
    .A(_15513_),
    .B(_15514_));
 sg13g2_xnor2_1 _46361_ (.Y(_15516_),
    .A(\u_inv.d_reg[47] ),
    .B(_15515_));
 sg13g2_o21ai_1 _46362_ (.B1(_15513_),
    .Y(_15517_),
    .A1(net7169),
    .A2(_18569_));
 sg13g2_xnor2_1 _46363_ (.Y(_15518_),
    .A(\u_inv.d_reg[46] ),
    .B(_15517_));
 sg13g2_nand2_1 _46364_ (.Y(_15519_),
    .A(net7274),
    .B(_15040_));
 sg13g2_xnor2_1 _46365_ (.Y(_15520_),
    .A(_18566_),
    .B(_15519_));
 sg13g2_nor3_1 _46366_ (.A(_15516_),
    .B(_15518_),
    .C(_15520_),
    .Y(_15521_));
 sg13g2_o21ai_1 _46367_ (.B1(net7274),
    .Y(_15522_),
    .A1(\u_inv.d_reg[48] ),
    .A2(_15040_));
 sg13g2_xnor2_1 _46368_ (.Y(_15523_),
    .A(_18565_),
    .B(_15522_));
 sg13g2_xnor2_1 _46369_ (.Y(_15524_),
    .A(_18569_),
    .B(_15513_));
 sg13g2_nor2_1 _46370_ (.A(net7169),
    .B(_15038_),
    .Y(_15525_));
 sg13g2_xnor2_1 _46371_ (.Y(_15526_),
    .A(\u_inv.d_reg[44] ),
    .B(_15525_));
 sg13g2_o21ai_1 _46372_ (.B1(net7273),
    .Y(_15527_),
    .A1(\u_inv.d_reg[42] ),
    .A2(_15037_));
 sg13g2_xnor2_1 _46373_ (.Y(_15528_),
    .A(net3765),
    .B(_15527_));
 sg13g2_xnor2_1 _46374_ (.Y(_15529_),
    .A(_18571_),
    .B(_15527_));
 sg13g2_nand2_1 _46375_ (.Y(_15530_),
    .A(net7273),
    .B(_15037_));
 sg13g2_xnor2_1 _46376_ (.Y(_15531_),
    .A(_18572_),
    .B(_15530_));
 sg13g2_a21oi_1 _46377_ (.A1(_18574_),
    .A2(net1106),
    .Y(_15532_),
    .B1(net7169));
 sg13g2_xnor2_1 _46378_ (.Y(_15533_),
    .A(\u_inv.d_reg[41] ),
    .B(_15532_));
 sg13g2_nor2_1 _46379_ (.A(net7169),
    .B(_15035_),
    .Y(_15534_));
 sg13g2_xnor2_1 _46380_ (.Y(_15535_),
    .A(\u_inv.d_reg[40] ),
    .B(_15534_));
 sg13g2_o21ai_1 _46381_ (.B1(net7273),
    .Y(_15536_),
    .A1(\u_inv.d_reg[38] ),
    .A2(_15034_));
 sg13g2_xnor2_1 _46382_ (.Y(_15537_),
    .A(_18575_),
    .B(_15536_));
 sg13g2_nand2_1 _46383_ (.Y(_15538_),
    .A(net7273),
    .B(_15034_));
 sg13g2_xnor2_1 _46384_ (.Y(_15539_),
    .A(_18576_),
    .B(_15538_));
 sg13g2_nand2_1 _46385_ (.Y(_15540_),
    .A(net7273),
    .B(net1137));
 sg13g2_xnor2_1 _46386_ (.Y(_15541_),
    .A(_18577_),
    .B(_15540_));
 sg13g2_o21ai_1 _46387_ (.B1(net7273),
    .Y(_15542_),
    .A1(\u_inv.d_reg[35] ),
    .A2(_15032_));
 sg13g2_xnor2_1 _46388_ (.Y(_15543_),
    .A(_18578_),
    .B(_15542_));
 sg13g2_nand2_1 _46389_ (.Y(_15544_),
    .A(net7273),
    .B(_15032_));
 sg13g2_xnor2_1 _46390_ (.Y(_15545_),
    .A(_18579_),
    .B(_15544_));
 sg13g2_nand2b_2 _46391_ (.Y(_15546_),
    .B(net7273),
    .A_N(_15031_));
 sg13g2_xnor2_1 _46392_ (.Y(_15547_),
    .A(\u_inv.d_reg[34] ),
    .B(_15546_));
 sg13g2_xnor2_1 _46393_ (.Y(_15548_),
    .A(_18580_),
    .B(_15546_));
 sg13g2_nand2_1 _46394_ (.Y(_15549_),
    .A(net7272),
    .B(_15030_));
 sg13g2_xnor2_1 _46395_ (.Y(_15550_),
    .A(\u_inv.d_reg[32] ),
    .B(_15549_));
 sg13g2_nor2_1 _46396_ (.A(net7171),
    .B(_15029_),
    .Y(_15551_));
 sg13g2_xnor2_1 _46397_ (.Y(_15552_),
    .A(\u_inv.d_reg[31] ),
    .B(_15551_));
 sg13g2_nor2_1 _46398_ (.A(net7171),
    .B(_15028_),
    .Y(_15553_));
 sg13g2_xnor2_1 _46399_ (.Y(_15554_),
    .A(\u_inv.d_reg[30] ),
    .B(_15553_));
 sg13g2_o21ai_1 _46400_ (.B1(net7272),
    .Y(_15555_),
    .A1(\u_inv.d_reg[28] ),
    .A2(_15027_));
 sg13g2_xnor2_1 _46401_ (.Y(_15556_),
    .A(_18585_),
    .B(_15555_));
 sg13g2_nand2_1 _46402_ (.Y(_15557_),
    .A(net7272),
    .B(_15027_));
 sg13g2_xnor2_1 _46403_ (.Y(_15558_),
    .A(\u_inv.d_reg[28] ),
    .B(_15557_));
 sg13g2_xnor2_1 _46404_ (.Y(_15559_),
    .A(_18586_),
    .B(_15557_));
 sg13g2_nor2_1 _46405_ (.A(net7166),
    .B(_15026_),
    .Y(_15560_));
 sg13g2_xnor2_1 _46406_ (.Y(_15561_),
    .A(_18587_),
    .B(_15560_));
 sg13g2_o21ai_1 _46407_ (.B1(net7272),
    .Y(_15562_),
    .A1(\u_inv.d_reg[25] ),
    .A2(_15025_));
 sg13g2_xnor2_1 _46408_ (.Y(_15563_),
    .A(_18588_),
    .B(_15562_));
 sg13g2_inv_2 _46409_ (.Y(_15564_),
    .A(_15563_));
 sg13g2_nand2_1 _46410_ (.Y(_15565_),
    .A(_15561_),
    .B(_15564_));
 sg13g2_nand2_1 _46411_ (.Y(_15566_),
    .A(net7265),
    .B(_15025_));
 sg13g2_xnor2_1 _46412_ (.Y(_15567_),
    .A(_18589_),
    .B(_15566_));
 sg13g2_inv_1 _46413_ (.Y(_15568_),
    .A(_15567_));
 sg13g2_o21ai_1 _46414_ (.B1(net7265),
    .Y(_15569_),
    .A1(net7291),
    .A2(net1132));
 sg13g2_xnor2_1 _46415_ (.Y(_15570_),
    .A(_18591_),
    .B(_15569_));
 sg13g2_nand2b_1 _46416_ (.Y(_15571_),
    .B(net7265),
    .A_N(_15022_));
 sg13g2_xnor2_1 _46417_ (.Y(_15572_),
    .A(\u_inv.d_reg[21] ),
    .B(_15571_));
 sg13g2_xnor2_1 _46418_ (.Y(_15573_),
    .A(_18593_),
    .B(_15571_));
 sg13g2_o21ai_1 _46419_ (.B1(net7265),
    .Y(_15574_),
    .A1(\u_inv.d_reg[19] ),
    .A2(net1096));
 sg13g2_xnor2_1 _46420_ (.Y(_15575_),
    .A(\u_inv.d_reg[20] ),
    .B(_15574_));
 sg13g2_xnor2_1 _46421_ (.Y(_15576_),
    .A(_18594_),
    .B(_15574_));
 sg13g2_nand2_1 _46422_ (.Y(_15577_),
    .A(net7265),
    .B(net1096));
 sg13g2_xnor2_1 _46423_ (.Y(_15578_),
    .A(_18595_),
    .B(_15577_));
 sg13g2_a21oi_1 _46424_ (.A1(_18597_),
    .A2(_15020_),
    .Y(_15579_),
    .B1(net7166));
 sg13g2_xnor2_1 _46425_ (.Y(_15580_),
    .A(\u_inv.d_reg[18] ),
    .B(_15579_));
 sg13g2_or2_1 _46426_ (.X(_15581_),
    .B(_15580_),
    .A(_15578_));
 sg13g2_nand2_1 _46427_ (.Y(_15582_),
    .A(net7268),
    .B(_15023_));
 sg13g2_xnor2_1 _46428_ (.Y(_15583_),
    .A(net7291),
    .B(_15582_));
 sg13g2_xnor2_1 _46429_ (.Y(_15584_),
    .A(_18592_),
    .B(_15582_));
 sg13g2_a21oi_1 _46430_ (.A1(_18598_),
    .A2(net1114),
    .Y(_15585_),
    .B1(net7166));
 sg13g2_xnor2_1 _46431_ (.Y(_15586_),
    .A(\u_inv.d_reg[17] ),
    .B(_15585_));
 sg13g2_nor2_1 _46432_ (.A(net7166),
    .B(net1113),
    .Y(_15587_));
 sg13g2_xnor2_1 _46433_ (.Y(_15588_),
    .A(\u_inv.d_reg[16] ),
    .B(_15587_));
 sg13g2_or2_1 _46434_ (.X(_15589_),
    .B(_15588_),
    .A(_15586_));
 sg13g2_or4_1 _46435_ (.A(_15573_),
    .B(_15576_),
    .C(_15581_),
    .D(_15589_),
    .X(_15590_));
 sg13g2_nor3_1 _46436_ (.A(_15570_),
    .B(_15584_),
    .C(_15590_),
    .Y(_15591_));
 sg13g2_nor2_1 _46437_ (.A(net7166),
    .B(_15018_),
    .Y(_15592_));
 sg13g2_xnor2_1 _46438_ (.Y(_15593_),
    .A(\u_inv.d_reg[15] ),
    .B(_15592_));
 sg13g2_o21ai_1 _46439_ (.B1(net7265),
    .Y(_15594_),
    .A1(\u_inv.d_reg[13] ),
    .A2(_15017_));
 sg13g2_xnor2_1 _46440_ (.Y(_15595_),
    .A(_18600_),
    .B(_15594_));
 sg13g2_nand2_1 _46441_ (.Y(_15596_),
    .A(net7265),
    .B(_15017_));
 sg13g2_xnor2_1 _46442_ (.Y(_15597_),
    .A(_18601_),
    .B(_15596_));
 sg13g2_nor2_1 _46443_ (.A(net7165),
    .B(_15016_),
    .Y(_15598_));
 sg13g2_xnor2_1 _46444_ (.Y(_15599_),
    .A(\u_inv.d_reg[12] ),
    .B(_15598_));
 sg13g2_nor2_1 _46445_ (.A(_15597_),
    .B(_15599_),
    .Y(_15600_));
 sg13g2_o21ai_1 _46446_ (.B1(net7263),
    .Y(_15601_),
    .A1(net7292),
    .A2(_15015_));
 sg13g2_xnor2_1 _46447_ (.Y(_15602_),
    .A(\u_inv.d_reg[11] ),
    .B(_15601_));
 sg13g2_xnor2_1 _46448_ (.Y(_15603_),
    .A(_18603_),
    .B(_15601_));
 sg13g2_nor2_1 _46449_ (.A(net7165),
    .B(_15014_),
    .Y(_15604_));
 sg13g2_xnor2_1 _46450_ (.Y(_15605_),
    .A(_18605_),
    .B(_15604_));
 sg13g2_o21ai_1 _46451_ (.B1(net7263),
    .Y(_15606_),
    .A1(\u_inv.d_reg[7] ),
    .A2(net1125));
 sg13g2_xnor2_1 _46452_ (.Y(_15607_),
    .A(_18606_),
    .B(_15606_));
 sg13g2_and2_1 _46453_ (.A(net7263),
    .B(_15013_),
    .X(_15608_));
 sg13g2_xnor2_1 _46454_ (.Y(_15609_),
    .A(\u_inv.d_reg[7] ),
    .B(_15608_));
 sg13g2_xnor2_1 _46455_ (.Y(_15610_),
    .A(_18607_),
    .B(_15608_));
 sg13g2_nor2_1 _46456_ (.A(net7165),
    .B(_15009_),
    .Y(_15611_));
 sg13g2_xnor2_1 _46457_ (.Y(_15612_),
    .A(\u_inv.d_reg[3] ),
    .B(_15611_));
 sg13g2_nand2_1 _46458_ (.Y(_15613_),
    .A(net7260),
    .B(net7294));
 sg13g2_xnor2_1 _46459_ (.Y(_15614_),
    .A(net7293),
    .B(_15613_));
 sg13g2_and2_1 _46460_ (.A(net7294),
    .B(_15614_),
    .X(_15615_));
 sg13g2_o21ai_1 _46461_ (.B1(net7260),
    .Y(_15616_),
    .A1(\u_inv.d_reg[0] ),
    .A2(\u_inv.d_reg[1] ));
 sg13g2_xnor2_1 _46462_ (.Y(_15617_),
    .A(\u_inv.d_reg[2] ),
    .B(_15616_));
 sg13g2_nand2_1 _46463_ (.Y(_15618_),
    .A(_15615_),
    .B(_15617_));
 sg13g2_or2_1 _46464_ (.X(_15619_),
    .B(_15618_),
    .A(_15612_));
 sg13g2_nand2_1 _46465_ (.Y(_15620_),
    .A(net7263),
    .B(net1116));
 sg13g2_xnor2_1 _46466_ (.Y(_15621_),
    .A(\u_inv.d_reg[4] ),
    .B(_15620_));
 sg13g2_xnor2_1 _46467_ (.Y(_15622_),
    .A(_18610_),
    .B(_15620_));
 sg13g2_nand2_1 _46468_ (.Y(_15623_),
    .A(_15619_),
    .B(_15622_));
 sg13g2_o21ai_1 _46469_ (.B1(net7263),
    .Y(_15624_),
    .A1(\u_inv.d_reg[4] ),
    .A2(_15011_));
 sg13g2_xnor2_1 _46470_ (.Y(_15625_),
    .A(\u_inv.d_reg[5] ),
    .B(_15624_));
 sg13g2_xnor2_1 _46471_ (.Y(_15626_),
    .A(_18609_),
    .B(_15624_));
 sg13g2_a21oi_1 _46472_ (.A1(_15619_),
    .A2(_15622_),
    .Y(_15627_),
    .B1(_15626_));
 sg13g2_o21ai_1 _46473_ (.B1(net7263),
    .Y(_15628_),
    .A1(\u_inv.d_reg[5] ),
    .A2(_15012_));
 sg13g2_xnor2_1 _46474_ (.Y(_15629_),
    .A(_18608_),
    .B(_15628_));
 sg13g2_nand3_1 _46475_ (.B(_15609_),
    .C(_15629_),
    .A(_15607_),
    .Y(_15630_));
 sg13g2_or3_1 _46476_ (.A(_15605_),
    .B(_15627_),
    .C(_15630_),
    .X(_15631_));
 sg13g2_nand2_1 _46477_ (.Y(_15632_),
    .A(net7263),
    .B(_15015_));
 sg13g2_xnor2_1 _46478_ (.Y(_15633_),
    .A(net7292),
    .B(_15632_));
 sg13g2_nand4_1 _46479_ (.B(_15602_),
    .C(_15631_),
    .A(_15600_),
    .Y(_15634_),
    .D(_15633_));
 sg13g2_nor3_2 _46480_ (.A(_15593_),
    .B(_15595_),
    .C(_15634_),
    .Y(_15635_));
 sg13g2_nor2_1 _46481_ (.A(net7166),
    .B(_15024_),
    .Y(_15636_));
 sg13g2_xnor2_1 _46482_ (.Y(_15637_),
    .A(\u_inv.d_reg[24] ),
    .B(_15636_));
 sg13g2_inv_1 _46483_ (.Y(_15638_),
    .A(_15637_));
 sg13g2_nand4_1 _46484_ (.B(_15591_),
    .C(_15635_),
    .A(_15568_),
    .Y(_15639_),
    .D(_15638_));
 sg13g2_or4_1 _46485_ (.A(_15556_),
    .B(_15559_),
    .C(_15565_),
    .D(_15639_),
    .X(_15640_));
 sg13g2_or3_1 _46486_ (.A(_15552_),
    .B(_15554_),
    .C(_15640_),
    .X(_15641_));
 sg13g2_nand2b_1 _46487_ (.Y(_15642_),
    .B(_15641_),
    .A_N(_15550_));
 sg13g2_o21ai_1 _46488_ (.B1(net7272),
    .Y(_15643_),
    .A1(\u_inv.d_reg[32] ),
    .A2(_15030_));
 sg13g2_or2_1 _46489_ (.X(_15644_),
    .B(_15643_),
    .A(_18581_));
 sg13g2_nand2_1 _46490_ (.Y(_15645_),
    .A(_18581_),
    .B(_15643_));
 sg13g2_and2_1 _46491_ (.A(_15644_),
    .B(_15645_),
    .X(_15646_));
 sg13g2_nand3_1 _46492_ (.B(_15642_),
    .C(_15646_),
    .A(_15547_),
    .Y(_15647_));
 sg13g2_or4_1 _46493_ (.A(_15541_),
    .B(_15543_),
    .C(_15545_),
    .D(_15647_),
    .X(_15648_));
 sg13g2_or3_1 _46494_ (.A(_15537_),
    .B(_15539_),
    .C(_15648_),
    .X(_15649_));
 sg13g2_nor4_1 _46495_ (.A(_15531_),
    .B(_15533_),
    .C(_15535_),
    .D(_15649_),
    .Y(_15650_));
 sg13g2_nand2_1 _46496_ (.Y(_15651_),
    .A(_15528_),
    .B(_15650_));
 sg13g2_nor4_1 _46497_ (.A(_15523_),
    .B(_15524_),
    .C(_15526_),
    .D(_15651_),
    .Y(_15652_));
 sg13g2_nand2_1 _46498_ (.Y(_15653_),
    .A(_15521_),
    .B(_15652_));
 sg13g2_or4_1 _46499_ (.A(_15508_),
    .B(_15510_),
    .C(_15512_),
    .D(_15653_),
    .X(_15654_));
 sg13g2_nor4_1 _46500_ (.A(_15502_),
    .B(_15504_),
    .C(_15506_),
    .D(_15654_),
    .Y(_15655_));
 sg13g2_nand4_1 _46501_ (.B(_15497_),
    .C(_15499_),
    .A(_15495_),
    .Y(_15656_),
    .D(_15655_));
 sg13g2_or3_1 _46502_ (.A(_15490_),
    .B(_15492_),
    .C(_15656_),
    .X(_15657_));
 sg13g2_or4_1 _46503_ (.A(_15484_),
    .B(_15486_),
    .C(_15488_),
    .D(_15657_),
    .X(_15658_));
 sg13g2_o21ai_1 _46504_ (.B1(net7281),
    .Y(_15659_),
    .A1(\u_inv.d_reg[64] ),
    .A2(_15054_));
 sg13g2_xnor2_1 _46505_ (.Y(_15660_),
    .A(_18549_),
    .B(_15659_));
 sg13g2_nor2_1 _46506_ (.A(net7172),
    .B(_15055_),
    .Y(_15661_));
 sg13g2_xnor2_1 _46507_ (.Y(_15662_),
    .A(\u_inv.d_reg[66] ),
    .B(_15661_));
 sg13g2_or2_1 _46508_ (.X(_15663_),
    .B(_15662_),
    .A(_15660_));
 sg13g2_nor4_1 _46509_ (.A(_15480_),
    .B(_15482_),
    .C(_15658_),
    .D(_15663_),
    .Y(_15664_));
 sg13g2_nand4_1 _46510_ (.B(_15475_),
    .C(_15478_),
    .A(_15473_),
    .Y(_15665_),
    .D(_15664_));
 sg13g2_or4_1 _46511_ (.A(_15466_),
    .B(_15468_),
    .C(_15470_),
    .D(_15665_),
    .X(_15666_));
 sg13g2_nor4_1 _46512_ (.A(_15458_),
    .B(_15461_),
    .C(_15464_),
    .D(_15666_),
    .Y(_15667_));
 sg13g2_nand4_1 _46513_ (.B(_15455_),
    .C(_15456_),
    .A(_15454_),
    .Y(_15668_),
    .D(_15667_));
 sg13g2_nor4_1 _46514_ (.A(_15431_),
    .B(_15437_),
    .C(_15445_),
    .D(_15668_),
    .Y(_15669_));
 sg13g2_nand3_1 _46515_ (.B(_15429_),
    .C(_15669_),
    .A(_15426_),
    .Y(_15670_));
 sg13g2_o21ai_1 _46516_ (.B1(net7283),
    .Y(_15671_),
    .A1(\u_inv.d_reg[88] ),
    .A2(net1082));
 sg13g2_xnor2_1 _46517_ (.Y(_15672_),
    .A(_18525_),
    .B(_15671_));
 sg13g2_inv_1 _46518_ (.Y(_15673_),
    .A(_15672_));
 sg13g2_nand2_1 _46519_ (.Y(_15674_),
    .A(net7277),
    .B(_15078_));
 sg13g2_xnor2_1 _46520_ (.Y(_15675_),
    .A(_18524_),
    .B(_15674_));
 sg13g2_nor4_1 _46521_ (.A(_15424_),
    .B(_15670_),
    .C(_15672_),
    .D(_15675_),
    .Y(_15676_));
 sg13g2_xnor2_1 _46522_ (.Y(_15677_),
    .A(\u_inv.d_reg[96] ),
    .B(_15404_));
 sg13g2_inv_1 _46523_ (.Y(_15678_),
    .A(_15677_));
 sg13g2_xnor2_1 _46524_ (.Y(_15679_),
    .A(\u_inv.d_reg[93] ),
    .B(_15400_));
 sg13g2_nand4_1 _46525_ (.B(_15676_),
    .C(_15678_),
    .A(_15422_),
    .Y(_15680_),
    .D(_15679_));
 sg13g2_a21oi_1 _46526_ (.A1(net7276),
    .A2(\u_inv.d_reg[98] ),
    .Y(_15681_),
    .B1(_15406_));
 sg13g2_xnor2_1 _46527_ (.Y(_15682_),
    .A(\u_inv.d_reg[99] ),
    .B(_15681_));
 sg13g2_xnor2_1 _46528_ (.Y(_15683_),
    .A(_18512_),
    .B(_15389_));
 sg13g2_nand2b_1 _46529_ (.Y(_15684_),
    .B(_15682_),
    .A_N(_15683_));
 sg13g2_or4_1 _46530_ (.A(_15418_),
    .B(_15421_),
    .C(_15680_),
    .D(_15684_),
    .X(_15685_));
 sg13g2_nor4_1 _46531_ (.A(_15386_),
    .B(_15413_),
    .C(_15415_),
    .D(_15685_),
    .Y(_15686_));
 sg13g2_o21ai_1 _46532_ (.B1(net7284),
    .Y(_15687_),
    .A1(\u_inv.d_reg[110] ),
    .A2(\u_inv.d_reg[109] ));
 sg13g2_nand3_1 _46533_ (.B(_15383_),
    .C(_15687_),
    .A(_15382_),
    .Y(_15688_));
 sg13g2_xnor2_1 _46534_ (.Y(_15689_),
    .A(_18503_),
    .B(_15688_));
 sg13g2_a21oi_1 _46535_ (.A1(net7284),
    .A2(\u_inv.d_reg[109] ),
    .Y(_15690_),
    .B1(_15384_));
 sg13g2_xnor2_1 _46536_ (.Y(_15691_),
    .A(\u_inv.d_reg[110] ),
    .B(_15690_));
 sg13g2_nand4_1 _46537_ (.B(_15686_),
    .C(_15689_),
    .A(_15385_),
    .Y(_15692_),
    .D(_15691_));
 sg13g2_nor4_1 _46538_ (.A(_15377_),
    .B(_15380_),
    .C(_15381_),
    .D(_15692_),
    .Y(_15693_));
 sg13g2_xnor2_1 _46539_ (.Y(_15694_),
    .A(_18489_),
    .B(_15369_));
 sg13g2_nand2_1 _46540_ (.Y(_15695_),
    .A(net7283),
    .B(_15091_));
 sg13g2_o21ai_1 _46541_ (.B1(_15695_),
    .Y(_15696_),
    .A1(net7173),
    .A2(_18502_));
 sg13g2_xnor2_1 _46542_ (.Y(_15697_),
    .A(_18501_),
    .B(_15696_));
 sg13g2_xnor2_1 _46543_ (.Y(_15698_),
    .A(\u_inv.d_reg[112] ),
    .B(_15695_));
 sg13g2_a21oi_1 _46544_ (.A1(net7283),
    .A2(\u_inv.d_reg[113] ),
    .Y(_15699_),
    .B1(_15696_));
 sg13g2_xnor2_1 _46545_ (.Y(_15700_),
    .A(\u_inv.d_reg[114] ),
    .B(_15699_));
 sg13g2_o21ai_1 _46546_ (.B1(net7283),
    .Y(_15701_),
    .A1(\u_inv.d_reg[114] ),
    .A2(\u_inv.d_reg[113] ));
 sg13g2_nor2b_1 _46547_ (.A(_15696_),
    .B_N(_15701_),
    .Y(_15702_));
 sg13g2_xnor2_1 _46548_ (.Y(_15703_),
    .A(\u_inv.d_reg[115] ),
    .B(_15702_));
 sg13g2_xnor2_1 _46549_ (.Y(_15704_),
    .A(_18496_),
    .B(_15375_));
 sg13g2_nor2b_1 _46550_ (.A(_15704_),
    .B_N(_15703_),
    .Y(_15705_));
 sg13g2_nand4_1 _46551_ (.B(_15698_),
    .C(_15700_),
    .A(_15697_),
    .Y(_15706_),
    .D(_15705_));
 sg13g2_nor2b_1 _46552_ (.A(_15706_),
    .B_N(_15694_),
    .Y(_15707_));
 sg13g2_a21oi_1 _46553_ (.A1(net7278),
    .A2(\u_inv.d_reg[120] ),
    .Y(_15708_),
    .B1(_15327_));
 sg13g2_xnor2_1 _46554_ (.Y(_15709_),
    .A(_18493_),
    .B(_15708_));
 sg13g2_xnor2_1 _46555_ (.Y(_15710_),
    .A(\u_inv.d_reg[120] ),
    .B(_15327_));
 sg13g2_nor2_1 _46556_ (.A(_15709_),
    .B(_15710_),
    .Y(_15711_));
 sg13g2_xnor2_1 _46557_ (.Y(_15712_),
    .A(_18470_),
    .B(_15317_));
 sg13g2_inv_4 _46558_ (.A(_15712_),
    .Y(_15713_));
 sg13g2_nand4_1 _46559_ (.B(_15707_),
    .C(_15711_),
    .A(_15693_),
    .Y(_15714_),
    .D(_15713_));
 sg13g2_nor3_2 _46560_ (.A(_15368_),
    .B(_15374_),
    .C(_15714_),
    .Y(_15715_));
 sg13g2_xnor2_1 _46561_ (.Y(_15716_),
    .A(\u_inv.d_reg[160] ),
    .B(_15288_));
 sg13g2_xnor2_1 _46562_ (.Y(_15717_),
    .A(\u_inv.d_reg[134] ),
    .B(_15358_));
 sg13g2_nand4_1 _46563_ (.B(_15715_),
    .C(_15716_),
    .A(_15366_),
    .Y(_15718_),
    .D(_15717_));
 sg13g2_o21ai_1 _46564_ (.B1(net7262),
    .Y(_15719_),
    .A1(net1085),
    .A2(_15123_));
 sg13g2_inv_1 _46565_ (.Y(_15720_),
    .A(_15719_));
 sg13g2_a21oi_1 _46566_ (.A1(net7268),
    .A2(\u_inv.d_reg[182] ),
    .Y(_15721_),
    .B1(_15720_));
 sg13g2_xnor2_1 _46567_ (.Y(_15722_),
    .A(\u_inv.d_reg[183] ),
    .B(_15721_));
 sg13g2_nand2_1 _46568_ (.Y(_15723_),
    .A(net7270),
    .B(_15305_));
 sg13g2_o21ai_1 _46569_ (.B1(net7270),
    .Y(_15724_),
    .A1(\u_inv.d_reg[136] ),
    .A2(_15305_));
 sg13g2_xnor2_1 _46570_ (.Y(_15725_),
    .A(net3761),
    .B(_15724_));
 sg13g2_xnor2_1 _46571_ (.Y(_15726_),
    .A(_18477_),
    .B(_15724_));
 sg13g2_xnor2_1 _46572_ (.Y(_15727_),
    .A(_18478_),
    .B(_15723_));
 sg13g2_o21ai_1 _46573_ (.B1(net7270),
    .Y(_15728_),
    .A1(_15102_),
    .A2(_15305_));
 sg13g2_xnor2_1 _46574_ (.Y(_15729_),
    .A(net3770),
    .B(_15728_));
 sg13g2_nor3_1 _46575_ (.A(\u_inv.d_reg[138] ),
    .B(_15102_),
    .C(_15305_),
    .Y(_15730_));
 sg13g2_nand2b_1 _46576_ (.Y(_15731_),
    .B(net7270),
    .A_N(_15730_));
 sg13g2_xnor2_1 _46577_ (.Y(_15732_),
    .A(\u_inv.d_reg[139] ),
    .B(_15731_));
 sg13g2_nand2_1 _46578_ (.Y(_15733_),
    .A(_15729_),
    .B(_15732_));
 sg13g2_nor3_2 _46579_ (.A(_15726_),
    .B(_15727_),
    .C(_15733_),
    .Y(_15734_));
 sg13g2_o21ai_1 _46580_ (.B1(net7267),
    .Y(_15735_),
    .A1(\u_inv.d_reg[168] ),
    .A2(_15119_));
 sg13g2_xnor2_1 _46581_ (.Y(_15736_),
    .A(\u_inv.d_reg[169] ),
    .B(_15735_));
 sg13g2_xnor2_1 _46582_ (.Y(_15737_),
    .A(\u_inv.d_reg[154] ),
    .B(_15271_));
 sg13g2_nand4_1 _46583_ (.B(_15734_),
    .C(_15736_),
    .A(_15722_),
    .Y(_15738_),
    .D(_15737_));
 sg13g2_nor4_1 _46584_ (.A(_15316_),
    .B(_15352_),
    .C(_15718_),
    .D(_15738_),
    .Y(_15739_));
 sg13g2_nor2_1 _46585_ (.A(net7167),
    .B(_15116_),
    .Y(_15740_));
 sg13g2_a21oi_1 _46586_ (.A1(net7266),
    .A2(_15290_),
    .Y(_15741_),
    .B1(_15740_));
 sg13g2_xnor2_1 _46587_ (.Y(_15742_),
    .A(\u_inv.d_reg[166] ),
    .B(_15741_));
 sg13g2_o21ai_1 _46588_ (.B1(net7267),
    .Y(_15743_),
    .A1(\u_inv.d_reg[173] ),
    .A2(\u_inv.d_reg[172] ));
 sg13g2_nor2b_1 _46589_ (.A(_15314_),
    .B_N(_15743_),
    .Y(_15744_));
 sg13g2_xnor2_1 _46590_ (.Y(_15745_),
    .A(\u_inv.d_reg[174] ),
    .B(_15744_));
 sg13g2_nand2_1 _46591_ (.Y(_15746_),
    .A(_15742_),
    .B(_15745_));
 sg13g2_nor3_1 _46592_ (.A(\u_inv.d_reg[170] ),
    .B(_15000_),
    .C(_15119_),
    .Y(_15747_));
 sg13g2_nand2b_1 _46593_ (.Y(_15748_),
    .B(\u_inv.d_reg[171] ),
    .A_N(_15747_));
 sg13g2_a22oi_1 _46594_ (.Y(_15749_),
    .B1(_15314_),
    .B2(_15748_),
    .A2(\u_inv.d_reg[171] ),
    .A1(net7166));
 sg13g2_o21ai_1 _46595_ (.B1(_15271_),
    .Y(_15750_),
    .A1(net7167),
    .A2(_18460_));
 sg13g2_xnor2_1 _46596_ (.Y(_15751_),
    .A(\u_inv.d_reg[155] ),
    .B(_15750_));
 sg13g2_xnor2_1 _46597_ (.Y(_15752_),
    .A(_18459_),
    .B(_15750_));
 sg13g2_nor3_1 _46598_ (.A(_15746_),
    .B(_15749_),
    .C(_15751_),
    .Y(_15753_));
 sg13g2_a21oi_1 _46599_ (.A1(net7271),
    .A2(\u_inv.d_reg[149] ),
    .Y(_15754_),
    .B1(_15363_));
 sg13g2_xnor2_1 _46600_ (.Y(_15755_),
    .A(\u_inv.d_reg[150] ),
    .B(_15754_));
 sg13g2_xnor2_1 _46601_ (.Y(_15756_),
    .A(\u_inv.d_reg[168] ),
    .B(_15311_));
 sg13g2_o21ai_1 _46602_ (.B1(_15278_),
    .Y(_15757_),
    .A1(net7167),
    .A2(_18456_));
 sg13g2_xnor2_1 _46603_ (.Y(_15758_),
    .A(_18455_),
    .B(_15757_));
 sg13g2_nand3_1 _46604_ (.B(_15756_),
    .C(_15758_),
    .A(_15755_),
    .Y(_15759_));
 sg13g2_o21ai_1 _46605_ (.B1(net7266),
    .Y(_15760_),
    .A1(_15112_),
    .A2(_15113_));
 sg13g2_xnor2_1 _46606_ (.Y(_15761_),
    .A(\u_inv.d_reg[162] ),
    .B(_15760_));
 sg13g2_o21ai_1 _46607_ (.B1(net7266),
    .Y(_15762_),
    .A1(\u_inv.d_reg[160] ),
    .A2(_15112_));
 sg13g2_xnor2_1 _46608_ (.Y(_15763_),
    .A(\u_inv.d_reg[161] ),
    .B(_15762_));
 sg13g2_xnor2_1 _46609_ (.Y(_15764_),
    .A(_18472_),
    .B(_15307_));
 sg13g2_inv_1 _46610_ (.Y(_15765_),
    .A(_15764_));
 sg13g2_o21ai_1 _46611_ (.B1(net7269),
    .Y(_15766_),
    .A1(_15103_),
    .A2(_15305_));
 sg13g2_xnor2_1 _46612_ (.Y(_15767_),
    .A(\u_inv.d_reg[140] ),
    .B(_15766_));
 sg13g2_nand4_1 _46613_ (.B(_15763_),
    .C(_15765_),
    .A(_15761_),
    .Y(_15768_),
    .D(_15767_));
 sg13g2_a21oi_1 _46614_ (.A1(net7267),
    .A2(\u_inv.d_reg[172] ),
    .Y(_15769_),
    .B1(_15314_));
 sg13g2_xnor2_1 _46615_ (.Y(_15770_),
    .A(\u_inv.d_reg[173] ),
    .B(_15769_));
 sg13g2_inv_1 _46616_ (.Y(_15771_),
    .A(_15770_));
 sg13g2_o21ai_1 _46617_ (.B1(_15269_),
    .Y(_15772_),
    .A1(net7167),
    .A2(_18462_));
 sg13g2_xnor2_1 _46618_ (.Y(_15773_),
    .A(\u_inv.d_reg[153] ),
    .B(_15772_));
 sg13g2_xnor2_1 _46619_ (.Y(_15774_),
    .A(_18462_),
    .B(_15269_));
 sg13g2_or2_1 _46620_ (.X(_15775_),
    .B(_15774_),
    .A(_15773_));
 sg13g2_nor4_1 _46621_ (.A(_15759_),
    .B(_15768_),
    .C(_15771_),
    .D(_15775_),
    .Y(_15776_));
 sg13g2_nand4_1 _46622_ (.B(_15739_),
    .C(_15753_),
    .A(_15300_),
    .Y(_15777_),
    .D(_15776_));
 sg13g2_and2_1 _46623_ (.A(net7257),
    .B(net1079),
    .X(_15778_));
 sg13g2_o21ai_1 _46624_ (.B1(net7260),
    .Y(_15779_),
    .A1(\u_inv.d_reg[200] ),
    .A2(net1130));
 sg13g2_xnor2_1 _46625_ (.Y(_15780_),
    .A(net3763),
    .B(_15779_));
 sg13g2_xnor2_1 _46626_ (.Y(_15781_),
    .A(_18414_),
    .B(_15778_));
 sg13g2_nand2_1 _46627_ (.Y(_15782_),
    .A(_15780_),
    .B(_15781_));
 sg13g2_nor3_1 _46628_ (.A(\u_inv.d_reg[210] ),
    .B(_15136_),
    .C(_15137_),
    .Y(_15783_));
 sg13g2_nor2_1 _46629_ (.A(net7164),
    .B(_15783_),
    .Y(_15784_));
 sg13g2_and2_1 _46630_ (.A(net7256),
    .B(_15136_),
    .X(_15785_));
 sg13g2_o21ai_1 _46631_ (.B1(net7256),
    .Y(_15786_),
    .A1(_15136_),
    .A2(_15138_));
 sg13g2_xnor2_1 _46632_ (.Y(_15787_),
    .A(_18403_),
    .B(_15784_));
 sg13g2_inv_1 _46633_ (.Y(_15788_),
    .A(_15787_));
 sg13g2_nor4_1 _46634_ (.A(_15282_),
    .B(_15777_),
    .C(_15782_),
    .D(_15788_),
    .Y(_15789_));
 sg13g2_xnor2_1 _46635_ (.Y(_15790_),
    .A(_18418_),
    .B(_15264_));
 sg13g2_a21oi_1 _46636_ (.A1(net7260),
    .A2(\u_inv.d_reg[192] ),
    .Y(_15791_),
    .B1(_15256_));
 sg13g2_a21o_1 _46637_ (.A2(_15791_),
    .A1(_18421_),
    .B1(net7165),
    .X(_15792_));
 sg13g2_xnor2_1 _46638_ (.Y(_15793_),
    .A(net3772),
    .B(_15792_));
 sg13g2_inv_2 _46639_ (.Y(_15794_),
    .A(_15793_));
 sg13g2_o21ai_1 _46640_ (.B1(net7260),
    .Y(_15795_),
    .A1(net1079),
    .A2(_15134_));
 sg13g2_inv_1 _46641_ (.Y(_15796_),
    .A(_15795_));
 sg13g2_o21ai_1 _46642_ (.B1(net7257),
    .Y(_15797_),
    .A1(net1079),
    .A2(_15135_));
 sg13g2_xnor2_1 _46643_ (.Y(_15798_),
    .A(_18408_),
    .B(_15797_));
 sg13g2_a21o_1 _46644_ (.A2(_15741_),
    .A1(_18448_),
    .B1(net7166),
    .X(_15799_));
 sg13g2_xnor2_1 _46645_ (.Y(_15800_),
    .A(_18447_),
    .B(_15799_));
 sg13g2_nor2_1 _46646_ (.A(net7168),
    .B(_15122_),
    .Y(_15801_));
 sg13g2_a21oi_1 _46647_ (.A1(net7262),
    .A2(net1085),
    .Y(_15802_),
    .B1(_15801_));
 sg13g2_inv_1 _46648_ (.Y(_15803_),
    .A(_15802_));
 sg13g2_a21oi_1 _46649_ (.A1(net7262),
    .A2(\u_inv.d_reg[180] ),
    .Y(_15804_),
    .B1(_15803_));
 sg13g2_xnor2_1 _46650_ (.Y(_15805_),
    .A(\u_inv.d_reg[181] ),
    .B(_15804_));
 sg13g2_xnor2_1 _46651_ (.Y(_15806_),
    .A(\u_inv.d_reg[182] ),
    .B(_15719_));
 sg13g2_xnor2_1 _46652_ (.Y(_15807_),
    .A(\u_inv.d_reg[180] ),
    .B(_15802_));
 sg13g2_nand3_1 _46653_ (.B(_15806_),
    .C(_15807_),
    .A(_15805_),
    .Y(_15808_));
 sg13g2_o21ai_1 _46654_ (.B1(net7261),
    .Y(_15809_),
    .A1(_15124_),
    .A2(_15126_));
 sg13g2_xnor2_1 _46655_ (.Y(_15810_),
    .A(\u_inv.d_reg[187] ),
    .B(_15809_));
 sg13g2_o21ai_1 _46656_ (.B1(net7261),
    .Y(_15811_),
    .A1(_15124_),
    .A2(_15125_));
 sg13g2_xnor2_1 _46657_ (.Y(_15812_),
    .A(\u_inv.d_reg[186] ),
    .B(_15811_));
 sg13g2_nand2_1 _46658_ (.Y(_15813_),
    .A(_15810_),
    .B(_15812_));
 sg13g2_nor3_1 _46659_ (.A(_15800_),
    .B(_15808_),
    .C(_15813_),
    .Y(_15814_));
 sg13g2_xnor2_1 _46660_ (.Y(_15815_),
    .A(_18416_),
    .B(_15245_));
 sg13g2_xnor2_1 _46661_ (.Y(_15816_),
    .A(\u_inv.d_reg[193] ),
    .B(_15791_));
 sg13g2_inv_1 _46662_ (.Y(_15817_),
    .A(_15816_));
 sg13g2_o21ai_1 _46663_ (.B1(net7261),
    .Y(_15818_),
    .A1(\u_inv.d_reg[184] ),
    .A2(net1115));
 sg13g2_xnor2_1 _46664_ (.Y(_15819_),
    .A(\u_inv.d_reg[185] ),
    .B(_15818_));
 sg13g2_xnor2_1 _46665_ (.Y(_15820_),
    .A(net2940),
    .B(_15253_));
 sg13g2_inv_1 _46666_ (.Y(_15821_),
    .A(_15820_));
 sg13g2_nand2_1 _46667_ (.Y(_15822_),
    .A(_15819_),
    .B(_15821_));
 sg13g2_a21o_1 _46668_ (.A2(_15259_),
    .A1(_18436_),
    .B1(_18435_),
    .X(_15823_));
 sg13g2_a22oi_1 _46669_ (.Y(_15824_),
    .B1(_15803_),
    .B2(_15823_),
    .A2(\u_inv.d_reg[179] ),
    .A1(net7168));
 sg13g2_nor4_1 _46670_ (.A(_15815_),
    .B(_15817_),
    .C(_15822_),
    .D(_15824_),
    .Y(_15825_));
 sg13g2_nand3b_1 _46671_ (.B(_18414_),
    .C(_18413_),
    .Y(_15826_),
    .A_N(net1079));
 sg13g2_nand2_1 _46672_ (.Y(_15827_),
    .A(net7264),
    .B(_15826_));
 sg13g2_xnor2_1 _46673_ (.Y(_15828_),
    .A(\u_inv.d_reg[202] ),
    .B(_15827_));
 sg13g2_xnor2_1 _46674_ (.Y(_15829_),
    .A(_18406_),
    .B(_15785_));
 sg13g2_nand4_1 _46675_ (.B(_15825_),
    .C(_15828_),
    .A(_15814_),
    .Y(_15830_),
    .D(_15829_));
 sg13g2_nor4_1 _46676_ (.A(_15790_),
    .B(_15794_),
    .C(_15798_),
    .D(_15830_),
    .Y(_15831_));
 sg13g2_o21ai_1 _46677_ (.B1(net7257),
    .Y(_15832_),
    .A1(_15136_),
    .A2(_15137_));
 sg13g2_xnor2_1 _46678_ (.Y(_15833_),
    .A(\u_inv.d_reg[210] ),
    .B(_15832_));
 sg13g2_o21ai_1 _46679_ (.B1(_15797_),
    .Y(_15834_),
    .A1(net7164),
    .A2(_18408_));
 sg13g2_xnor2_1 _46680_ (.Y(_15835_),
    .A(net3767),
    .B(_15834_));
 sg13g2_inv_1 _46681_ (.Y(_15836_),
    .A(_15835_));
 sg13g2_nor2_2 _46682_ (.A(net7164),
    .B(_15140_),
    .Y(_15837_));
 sg13g2_xnor2_1 _46683_ (.Y(_15838_),
    .A(_18398_),
    .B(_15837_));
 sg13g2_nand3_1 _46684_ (.B(_15836_),
    .C(_15838_),
    .A(_15833_),
    .Y(_15839_));
 sg13g2_o21ai_1 _46685_ (.B1(\u_inv.d_reg[203] ),
    .Y(_15840_),
    .A1(\u_inv.d_reg[202] ),
    .A2(_15826_));
 sg13g2_a22oi_1 _46686_ (.Y(_15841_),
    .B1(_15796_),
    .B2(_15840_),
    .A2(\u_inv.d_reg[203] ),
    .A1(net7164));
 sg13g2_o21ai_1 _46687_ (.B1(net7256),
    .Y(_15842_),
    .A1(_15136_),
    .A2(_15139_));
 sg13g2_inv_1 _46688_ (.Y(_15843_),
    .A(_15842_));
 sg13g2_xnor2_1 _46689_ (.Y(_15844_),
    .A(net3771),
    .B(_15842_));
 sg13g2_inv_1 _46690_ (.Y(_15845_),
    .A(_15844_));
 sg13g2_o21ai_1 _46691_ (.B1(_15795_),
    .Y(_15846_),
    .A1(net7164),
    .A2(_18410_));
 sg13g2_xnor2_1 _46692_ (.Y(_15847_),
    .A(_18409_),
    .B(_15846_));
 sg13g2_xnor2_1 _46693_ (.Y(_15848_),
    .A(net2833),
    .B(_15795_));
 sg13g2_nand2_1 _46694_ (.Y(_15849_),
    .A(_15847_),
    .B(_15848_));
 sg13g2_o21ai_1 _46695_ (.B1(net7257),
    .Y(_15850_),
    .A1(\u_inv.d_reg[208] ),
    .A2(_15136_));
 sg13g2_xnor2_1 _46696_ (.Y(_15851_),
    .A(\u_inv.d_reg[209] ),
    .B(_15850_));
 sg13g2_nand2b_1 _46697_ (.Y(_15852_),
    .B(_15851_),
    .A_N(_15849_));
 sg13g2_nor4_1 _46698_ (.A(_15839_),
    .B(_15841_),
    .C(_15845_),
    .D(_15852_),
    .Y(_15853_));
 sg13g2_xnor2_1 _46699_ (.Y(_15854_),
    .A(_15208_),
    .B(_18378_));
 sg13g2_nand2_1 _46700_ (.Y(_15855_),
    .A(_15140_),
    .B(_15144_));
 sg13g2_nand2_1 _46701_ (.Y(_15856_),
    .A(net7259),
    .B(_15855_));
 sg13g2_xnor2_1 _46702_ (.Y(_15857_),
    .A(_18392_),
    .B(_15856_));
 sg13g2_a21oi_1 _46703_ (.A1(net7256),
    .A2(\u_inv.d_reg[216] ),
    .Y(_15858_),
    .B1(_15837_));
 sg13g2_xnor2_1 _46704_ (.Y(_15859_),
    .A(\u_inv.d_reg[217] ),
    .B(_15858_));
 sg13g2_nand2b_1 _46705_ (.Y(_15860_),
    .B(_15859_),
    .A_N(_15857_));
 sg13g2_a21oi_1 _46706_ (.A1(net7256),
    .A2(\u_inv.d_reg[214] ),
    .Y(_15861_),
    .B1(_15843_));
 sg13g2_xnor2_1 _46707_ (.Y(_15862_),
    .A(_18399_),
    .B(_15861_));
 sg13g2_xnor2_1 _46708_ (.Y(_15863_),
    .A(_18402_),
    .B(_15786_));
 sg13g2_nand2_1 _46709_ (.Y(_15864_),
    .A(net7257),
    .B(\u_inv.d_reg[212] ));
 sg13g2_and2_1 _46710_ (.A(_15786_),
    .B(_15864_),
    .X(_15865_));
 sg13g2_xnor2_1 _46711_ (.Y(_15866_),
    .A(_18401_),
    .B(_15865_));
 sg13g2_inv_1 _46712_ (.Y(_15867_),
    .A(_15866_));
 sg13g2_or2_1 _46713_ (.X(_15868_),
    .B(_15866_),
    .A(_15863_));
 sg13g2_nor4_1 _46714_ (.A(net1123),
    .B(_15860_),
    .C(_15862_),
    .D(_15868_),
    .Y(_15869_));
 sg13g2_and4_2 _46715_ (.A(_15789_),
    .B(_15831_),
    .C(_15869_),
    .D(_15853_),
    .X(_15870_));
 sg13g2_o21ai_1 _46716_ (.B1(net7259),
    .Y(_15871_),
    .A1(\u_inv.d_reg[222] ),
    .A2(_15855_));
 sg13g2_xnor2_1 _46717_ (.Y(_15872_),
    .A(_18391_),
    .B(_15871_));
 sg13g2_nand2_1 _46718_ (.Y(_15873_),
    .A(net7252),
    .B(_15150_));
 sg13g2_xnor2_1 _46719_ (.Y(_15874_),
    .A(_18382_),
    .B(_15873_));
 sg13g2_a21o_1 _46720_ (.A2(_15141_),
    .A1(net1099),
    .B1(net7176),
    .X(_15875_));
 sg13g2_xnor2_1 _46721_ (.Y(_15876_),
    .A(\u_inv.d_reg[219] ),
    .B(_15875_));
 sg13g2_o21ai_1 _46722_ (.B1(net7256),
    .Y(_15877_),
    .A1(\u_inv.d_reg[217] ),
    .A2(\u_inv.d_reg[216] ));
 sg13g2_nor2b_1 _46723_ (.A(_15837_),
    .B_N(_15877_),
    .Y(_15878_));
 sg13g2_xnor2_1 _46724_ (.Y(_15879_),
    .A(\u_inv.d_reg[218] ),
    .B(_15878_));
 sg13g2_nand2_1 _46725_ (.Y(_15880_),
    .A(_15876_),
    .B(_15879_));
 sg13g2_nor3_1 _46726_ (.A(_15872_),
    .B(_15874_),
    .C(_15880_),
    .Y(_15881_));
 sg13g2_o21ai_1 _46727_ (.B1(net7252),
    .Y(_15882_),
    .A1(net1069),
    .A2(_15147_));
 sg13g2_xnor2_1 _46728_ (.Y(_15883_),
    .A(\u_inv.d_reg[229] ),
    .B(_15882_));
 sg13g2_xnor2_1 _46729_ (.Y(_15884_),
    .A(_18386_),
    .B(_15241_));
 sg13g2_and2_1 _46730_ (.A(_15883_),
    .B(_15884_),
    .X(_15885_));
 sg13g2_a21oi_1 _46731_ (.A1(net7256),
    .A2(_15143_),
    .Y(_15886_),
    .B1(_15837_));
 sg13g2_xnor2_1 _46732_ (.Y(_15887_),
    .A(\u_inv.d_reg[221] ),
    .B(_15886_));
 sg13g2_a21oi_1 _46733_ (.A1(net7256),
    .A2(_15142_),
    .Y(_15888_),
    .B1(_15837_));
 sg13g2_xnor2_1 _46734_ (.Y(_15889_),
    .A(\u_inv.d_reg[220] ),
    .B(_15888_));
 sg13g2_nand2_1 _46735_ (.Y(_15890_),
    .A(_15887_),
    .B(_15889_));
 sg13g2_inv_1 _46736_ (.Y(_15891_),
    .A(_15890_));
 sg13g2_xnor2_1 _46737_ (.Y(_15892_),
    .A(\u_inv.d_reg[230] ),
    .B(_15224_));
 sg13g2_nor2b_1 _46738_ (.A(_15890_),
    .B_N(_15892_),
    .Y(_15893_));
 sg13g2_nand4_1 _46739_ (.B(_15881_),
    .C(_15885_),
    .A(_15870_),
    .Y(_15894_),
    .D(_15893_));
 sg13g2_nor4_1 _46740_ (.A(_15235_),
    .B(_15237_),
    .C(_15244_),
    .D(_15894_),
    .Y(_15895_));
 sg13g2_nand4_1 _46741_ (.B(_15231_),
    .C(_15895_),
    .A(_15229_),
    .Y(_15896_),
    .D(_15234_));
 sg13g2_nor4_2 _46742_ (.A(_15200_),
    .B(_15202_),
    .C(_15207_),
    .Y(_15897_),
    .D(_15896_));
 sg13g2_nand3_1 _46743_ (.B(_15199_),
    .C(_15897_),
    .A(_15196_),
    .Y(_15898_));
 sg13g2_nor4_2 _46744_ (.A(_15898_),
    .B(_15171_),
    .C(_15193_),
    .Y(_15899_),
    .D(net5347));
 sg13g2_inv_8 _46745_ (.Y(_15900_),
    .A(net5308));
 sg13g2_nor2_2 _46746_ (.A(net5358),
    .B(net5312),
    .Y(_15901_));
 sg13g2_or2_1 _46747_ (.X(_15902_),
    .B(net5308),
    .A(net5356));
 sg13g2_xnor2_1 _46748_ (.Y(_15903_),
    .A(_18357_),
    .B(net5179));
 sg13g2_a21oi_1 _46749_ (.A1(net6698),
    .A2(_15903_),
    .Y(_00994_),
    .B1(_14999_));
 sg13g2_a21oi_1 _46750_ (.A1(_18357_),
    .A2(_18613_),
    .Y(_15904_),
    .B1(_15615_));
 sg13g2_nor2_1 _46751_ (.A(net5353),
    .B(_15904_),
    .Y(_15905_));
 sg13g2_a21oi_1 _46752_ (.A1(net5191),
    .A2(_15904_),
    .Y(_15906_),
    .B1(_15905_));
 sg13g2_nand2_1 _46753_ (.Y(_15907_),
    .A(_15614_),
    .B(net5180));
 sg13g2_nor2_1 _46754_ (.A(net6617),
    .B(_15906_),
    .Y(_15908_));
 sg13g2_a22oi_1 _46755_ (.Y(_00995_),
    .B1(_15907_),
    .B2(_15908_),
    .A2(net6617),
    .A1(_18267_));
 sg13g2_a21oi_1 _46756_ (.A1(_15615_),
    .A2(net5307),
    .Y(_15909_),
    .B1(_15617_));
 sg13g2_nor2_1 _46757_ (.A(_15618_),
    .B(net5192),
    .Y(_15910_));
 sg13g2_nor3_1 _46758_ (.A(net5353),
    .B(_15909_),
    .C(_15910_),
    .Y(_15911_));
 sg13g2_o21ai_1 _46759_ (.B1(_15617_),
    .Y(_15912_),
    .A1(net7294),
    .A2(net7293));
 sg13g2_a21oi_1 _46760_ (.A1(_15010_),
    .A2(_15912_),
    .Y(_15913_),
    .B1(net5327));
 sg13g2_nor3_1 _46761_ (.A(net6617),
    .B(_15911_),
    .C(_15913_),
    .Y(_15914_));
 sg13g2_a21oi_1 _46762_ (.A1(_18269_),
    .A2(net6617),
    .Y(_00996_),
    .B1(_15914_));
 sg13g2_o21ai_1 _46763_ (.B1(_15612_),
    .Y(_15915_),
    .A1(_15618_),
    .A2(net5192));
 sg13g2_o21ai_1 _46764_ (.B1(net5327),
    .Y(_15916_),
    .A1(_15619_),
    .A2(net5192));
 sg13g2_nand2b_1 _46765_ (.Y(_15917_),
    .B(_15915_),
    .A_N(_15916_));
 sg13g2_o21ai_1 _46766_ (.B1(_15011_),
    .Y(_15918_),
    .A1(_15009_),
    .A2(_15612_));
 sg13g2_a21oi_1 _46767_ (.A1(net5353),
    .A2(_15918_),
    .Y(_15919_),
    .B1(net6617));
 sg13g2_a22oi_1 _46768_ (.Y(_00997_),
    .B1(_15917_),
    .B2(_15919_),
    .A2(net6617),
    .A1(_18268_));
 sg13g2_nand2_1 _46769_ (.Y(_15920_),
    .A(_15619_),
    .B(net5307));
 sg13g2_a21oi_1 _46770_ (.A1(_15622_),
    .A2(_15920_),
    .Y(_15921_),
    .B1(net5353));
 sg13g2_o21ai_1 _46771_ (.B1(_15921_),
    .Y(_15922_),
    .A1(_15622_),
    .A2(_15920_));
 sg13g2_a21oi_1 _46772_ (.A1(_15011_),
    .A2(_15621_),
    .Y(_15923_),
    .B1(net5327));
 sg13g2_a21oi_1 _46773_ (.A1(_15012_),
    .A2(_15923_),
    .Y(_15924_),
    .B1(net6617));
 sg13g2_a22oi_1 _46774_ (.Y(_00998_),
    .B1(_15922_),
    .B2(_15924_),
    .A2(net6617),
    .A1(_18270_));
 sg13g2_nor2_1 _46775_ (.A(net2111),
    .B(net6697),
    .Y(_15925_));
 sg13g2_a21oi_1 _46776_ (.A1(_15623_),
    .A2(net5307),
    .Y(_15926_),
    .B1(_15923_));
 sg13g2_xnor2_1 _46777_ (.Y(_15927_),
    .A(_15626_),
    .B(_15926_));
 sg13g2_a21oi_1 _46778_ (.A1(net6697),
    .A2(_15927_),
    .Y(_00999_),
    .B1(_15925_));
 sg13g2_nor2_1 _46779_ (.A(net2551),
    .B(net6697),
    .Y(_15928_));
 sg13g2_a21oi_1 _46780_ (.A1(_15011_),
    .A2(_15621_),
    .Y(_15929_),
    .B1(_15625_));
 sg13g2_nor2_1 _46781_ (.A(net5327),
    .B(_15929_),
    .Y(_15930_));
 sg13g2_nor2b_1 _46782_ (.A(_15627_),
    .B_N(net5307),
    .Y(_15931_));
 sg13g2_or2_1 _46783_ (.X(_15932_),
    .B(_15931_),
    .A(_15930_));
 sg13g2_xor2_1 _46784_ (.B(_15932_),
    .A(_15629_),
    .X(_15933_));
 sg13g2_a21oi_1 _46785_ (.A1(net6697),
    .A2(_15933_),
    .Y(_01000_),
    .B1(_15928_));
 sg13g2_nor2_1 _46786_ (.A(net1383),
    .B(net6697),
    .Y(_15934_));
 sg13g2_nor3_1 _46787_ (.A(net5327),
    .B(_15629_),
    .C(_15929_),
    .Y(_15935_));
 sg13g2_nand2_1 _46788_ (.Y(_15936_),
    .A(_15629_),
    .B(_15931_));
 sg13g2_nand2b_1 _46789_ (.Y(_15937_),
    .B(_15936_),
    .A_N(_15935_));
 sg13g2_xnor2_1 _46790_ (.Y(_15938_),
    .A(_15610_),
    .B(_15937_));
 sg13g2_a21oi_1 _46791_ (.A1(net6697),
    .A2(_15938_),
    .Y(_01001_),
    .B1(_15934_));
 sg13g2_nor2_1 _46792_ (.A(net2099),
    .B(net6699),
    .Y(_15939_));
 sg13g2_nor2_1 _46793_ (.A(_15610_),
    .B(_15936_),
    .Y(_15940_));
 sg13g2_a21oi_1 _46794_ (.A1(_15610_),
    .A2(_15935_),
    .Y(_15941_),
    .B1(_15940_));
 sg13g2_xnor2_1 _46795_ (.Y(_15942_),
    .A(_15607_),
    .B(_15941_));
 sg13g2_a21oi_1 _46796_ (.A1(net6699),
    .A2(_15942_),
    .Y(_01002_),
    .B1(_15939_));
 sg13g2_nor2_1 _46797_ (.A(net2236),
    .B(net6699),
    .Y(_15943_));
 sg13g2_nand2b_1 _46798_ (.Y(_15944_),
    .B(net5327),
    .A_N(_15607_));
 sg13g2_nor4_1 _46799_ (.A(_15607_),
    .B(_15609_),
    .C(_15629_),
    .D(_15929_),
    .Y(_15945_));
 sg13g2_o21ai_1 _46800_ (.B1(_15944_),
    .Y(_15946_),
    .A1(_15940_),
    .A2(_15945_));
 sg13g2_xor2_1 _46801_ (.B(_15946_),
    .A(_15605_),
    .X(_15947_));
 sg13g2_a21oi_1 _46802_ (.A1(net6699),
    .A2(_15947_),
    .Y(_01003_),
    .B1(_15943_));
 sg13g2_a21oi_1 _46803_ (.A1(_15605_),
    .A2(_15945_),
    .Y(_15948_),
    .B1(net5328));
 sg13g2_a21oi_1 _46804_ (.A1(_15631_),
    .A2(net5307),
    .Y(_15949_),
    .B1(_15948_));
 sg13g2_xnor2_1 _46805_ (.Y(_15950_),
    .A(_15633_),
    .B(_15949_));
 sg13g2_mux2_1 _46806_ (.A0(net3328),
    .A1(_15950_),
    .S(net6699),
    .X(_01004_));
 sg13g2_nor2_1 _46807_ (.A(net1793),
    .B(net6700),
    .Y(_15951_));
 sg13g2_a21oi_1 _46808_ (.A1(_15605_),
    .A2(_15945_),
    .Y(_15952_),
    .B1(_15633_));
 sg13g2_and3_1 _46809_ (.X(_15953_),
    .A(_15631_),
    .B(_15633_),
    .C(net5307));
 sg13g2_a21oi_1 _46810_ (.A1(net5354),
    .A2(_15952_),
    .Y(_15954_),
    .B1(_15953_));
 sg13g2_xnor2_1 _46811_ (.Y(_15955_),
    .A(_15603_),
    .B(_15954_));
 sg13g2_a21oi_1 _46812_ (.A1(net6699),
    .A2(_15955_),
    .Y(_01005_),
    .B1(_15951_));
 sg13g2_nor2_1 _46813_ (.A(net1848),
    .B(net6699),
    .Y(_15956_));
 sg13g2_nand3_1 _46814_ (.B(_15603_),
    .C(_15952_),
    .A(net5354),
    .Y(_15957_));
 sg13g2_and2_1 _46815_ (.A(_15602_),
    .B(_15953_),
    .X(_15958_));
 sg13g2_inv_1 _46816_ (.Y(_15959_),
    .A(_15958_));
 sg13g2_nand2_1 _46817_ (.Y(_15960_),
    .A(_15957_),
    .B(_15959_));
 sg13g2_xor2_1 _46818_ (.B(_15960_),
    .A(_15599_),
    .X(_15961_));
 sg13g2_a21oi_1 _46819_ (.A1(net6699),
    .A2(_15961_),
    .Y(_01006_),
    .B1(_15956_));
 sg13g2_nor2_1 _46820_ (.A(net2136),
    .B(net6700),
    .Y(_15962_));
 sg13g2_nand3_1 _46821_ (.B(_15603_),
    .C(_15952_),
    .A(_15599_),
    .Y(_15963_));
 sg13g2_a22oi_1 _46822_ (.Y(_15964_),
    .B1(_15959_),
    .B2(_15963_),
    .A2(_15599_),
    .A1(net5328));
 sg13g2_xor2_1 _46823_ (.B(_15964_),
    .A(_15597_),
    .X(_15965_));
 sg13g2_a21oi_1 _46824_ (.A1(net6700),
    .A2(_15965_),
    .Y(_01007_),
    .B1(_15962_));
 sg13g2_nor2_1 _46825_ (.A(net1910),
    .B(net6700),
    .Y(_15966_));
 sg13g2_and4_1 _46826_ (.A(_15597_),
    .B(_15599_),
    .C(_15603_),
    .D(_15952_),
    .X(_15967_));
 sg13g2_and2_1 _46827_ (.A(_15600_),
    .B(_15958_),
    .X(_15968_));
 sg13g2_a21oi_1 _46828_ (.A1(net5354),
    .A2(_15967_),
    .Y(_15969_),
    .B1(_15968_));
 sg13g2_xnor2_1 _46829_ (.Y(_15970_),
    .A(_15595_),
    .B(_15969_));
 sg13g2_a21oi_1 _46830_ (.A1(net6700),
    .A2(_15970_),
    .Y(_01008_),
    .B1(_15966_));
 sg13g2_nor2_1 _46831_ (.A(net1485),
    .B(net6700),
    .Y(_15971_));
 sg13g2_and2_1 _46832_ (.A(_15595_),
    .B(_15967_),
    .X(_15972_));
 sg13g2_nand2_1 _46833_ (.Y(_15973_),
    .A(net5328),
    .B(_15595_));
 sg13g2_o21ai_1 _46834_ (.B1(_15973_),
    .Y(_15974_),
    .A1(_15968_),
    .A2(_15972_));
 sg13g2_xnor2_1 _46835_ (.Y(_15975_),
    .A(_15593_),
    .B(_15974_));
 sg13g2_a21oi_1 _46836_ (.A1(net6700),
    .A2(_15975_),
    .Y(_01009_),
    .B1(_15971_));
 sg13g2_nor2_1 _46837_ (.A(net1513),
    .B(net6704),
    .Y(_15976_));
 sg13g2_and3_1 _46838_ (.X(_15977_),
    .A(net5355),
    .B(_15593_),
    .C(_15972_));
 sg13g2_and2_1 _46839_ (.A(_15635_),
    .B(net5308),
    .X(_15978_));
 sg13g2_nor2_1 _46840_ (.A(_15977_),
    .B(_15978_),
    .Y(_15979_));
 sg13g2_xnor2_1 _46841_ (.Y(_15980_),
    .A(_15588_),
    .B(_15979_));
 sg13g2_a21oi_1 _46842_ (.A1(net6704),
    .A2(_15980_),
    .Y(_01010_),
    .B1(_15976_));
 sg13g2_nor2_1 _46843_ (.A(net2412),
    .B(net6704),
    .Y(_15981_));
 sg13g2_and4_1 _46844_ (.A(_15588_),
    .B(_15593_),
    .C(_15595_),
    .D(_15967_),
    .X(_15982_));
 sg13g2_nand2_1 _46845_ (.Y(_15983_),
    .A(net5330),
    .B(_15588_));
 sg13g2_o21ai_1 _46846_ (.B1(_15983_),
    .Y(_15984_),
    .A1(_15978_),
    .A2(_15982_));
 sg13g2_xnor2_1 _46847_ (.Y(_15985_),
    .A(_15586_),
    .B(_15984_));
 sg13g2_a21oi_1 _46848_ (.A1(net6704),
    .A2(_15985_),
    .Y(_01011_),
    .B1(_15981_));
 sg13g2_nand2_1 _46849_ (.Y(_15986_),
    .A(_15586_),
    .B(_15982_));
 sg13g2_nand2b_2 _46850_ (.Y(_15987_),
    .B(_15978_),
    .A_N(_15589_));
 sg13g2_o21ai_1 _46851_ (.B1(_15987_),
    .Y(_15988_),
    .A1(net5330),
    .A2(_15986_));
 sg13g2_xor2_1 _46852_ (.B(_15988_),
    .A(_15580_),
    .X(_15989_));
 sg13g2_nand2_1 _46853_ (.Y(_15990_),
    .A(net1201),
    .B(net6622));
 sg13g2_o21ai_1 _46854_ (.B1(_15990_),
    .Y(_01012_),
    .A1(net6621),
    .A2(_15989_));
 sg13g2_nor2_1 _46855_ (.A(net2297),
    .B(net6706),
    .Y(_15991_));
 sg13g2_nand3_1 _46856_ (.B(_15586_),
    .C(_15982_),
    .A(_15580_),
    .Y(_15992_));
 sg13g2_a22oi_1 _46857_ (.Y(_15993_),
    .B1(_15987_),
    .B2(_15992_),
    .A2(_15580_),
    .A1(net5331));
 sg13g2_xor2_1 _46858_ (.B(_15993_),
    .A(_15578_),
    .X(_15994_));
 sg13g2_a21oi_1 _46859_ (.A1(net6706),
    .A2(_15994_),
    .Y(_01013_),
    .B1(_15991_));
 sg13g2_nor2_1 _46860_ (.A(net2155),
    .B(net6705),
    .Y(_15995_));
 sg13g2_nand4_1 _46861_ (.B(_15580_),
    .C(_15586_),
    .A(_15578_),
    .Y(_15996_),
    .D(_15982_));
 sg13g2_nor2_1 _46862_ (.A(net5330),
    .B(_15996_),
    .Y(_15997_));
 sg13g2_nor2_1 _46863_ (.A(_15581_),
    .B(_15987_),
    .Y(_15998_));
 sg13g2_or2_1 _46864_ (.X(_15999_),
    .B(_15998_),
    .A(_15997_));
 sg13g2_xnor2_1 _46865_ (.Y(_16000_),
    .A(_15575_),
    .B(_15999_));
 sg13g2_a21oi_1 _46866_ (.A1(net6704),
    .A2(_16000_),
    .Y(_01014_),
    .B1(_15995_));
 sg13g2_nor2_1 _46867_ (.A(net1968),
    .B(net6710),
    .Y(_16001_));
 sg13g2_nand2_1 _46868_ (.Y(_16002_),
    .A(net5330),
    .B(_15576_));
 sg13g2_nor2_1 _46869_ (.A(_15575_),
    .B(_15996_),
    .Y(_16003_));
 sg13g2_o21ai_1 _46870_ (.B1(_16002_),
    .Y(_16004_),
    .A1(_15998_),
    .A2(_16003_));
 sg13g2_xnor2_1 _46871_ (.Y(_16005_),
    .A(_15573_),
    .B(_16004_));
 sg13g2_a21oi_1 _46872_ (.A1(net6706),
    .A2(_16005_),
    .Y(_01015_),
    .B1(_16001_));
 sg13g2_nor2_1 _46873_ (.A(net1998),
    .B(net6705),
    .Y(_16006_));
 sg13g2_nor4_1 _46874_ (.A(net5330),
    .B(_15572_),
    .C(_15575_),
    .D(_15996_),
    .Y(_16007_));
 sg13g2_nor4_1 _46875_ (.A(_15573_),
    .B(_15576_),
    .C(_15581_),
    .D(_15987_),
    .Y(_16008_));
 sg13g2_nor2_1 _46876_ (.A(_16007_),
    .B(_16008_),
    .Y(_16009_));
 sg13g2_xnor2_1 _46877_ (.Y(_16010_),
    .A(_15584_),
    .B(_16009_));
 sg13g2_a21oi_1 _46878_ (.A1(net6705),
    .A2(_16010_),
    .Y(_01016_),
    .B1(_16006_));
 sg13g2_nor2_1 _46879_ (.A(net2005),
    .B(net6705),
    .Y(_16011_));
 sg13g2_nand2_1 _46880_ (.Y(_16012_),
    .A(net5330),
    .B(_15584_));
 sg13g2_nor4_2 _46881_ (.A(_15572_),
    .B(_15575_),
    .C(_15583_),
    .Y(_16013_),
    .D(_15996_));
 sg13g2_o21ai_1 _46882_ (.B1(_16012_),
    .Y(_16014_),
    .A1(_16008_),
    .A2(_16013_));
 sg13g2_xnor2_1 _46883_ (.Y(_16015_),
    .A(_15570_),
    .B(_16014_));
 sg13g2_a21oi_1 _46884_ (.A1(net6704),
    .A2(_16015_),
    .Y(_01017_),
    .B1(_16011_));
 sg13g2_nand2_1 _46885_ (.Y(_16016_),
    .A(_15570_),
    .B(_16013_));
 sg13g2_nand2_1 _46886_ (.Y(_16017_),
    .A(_15591_),
    .B(_15978_));
 sg13g2_o21ai_1 _46887_ (.B1(_16017_),
    .Y(_16018_),
    .A1(net5330),
    .A2(_16016_));
 sg13g2_xnor2_1 _46888_ (.Y(_16019_),
    .A(_15638_),
    .B(_16018_));
 sg13g2_nand2_1 _46889_ (.Y(_16020_),
    .A(net1190),
    .B(net6621));
 sg13g2_o21ai_1 _46890_ (.B1(_16020_),
    .Y(_01018_),
    .A1(net6621),
    .A2(_16019_));
 sg13g2_nor2_1 _46891_ (.A(net2128),
    .B(net6704),
    .Y(_16021_));
 sg13g2_nand3_1 _46892_ (.B(_15637_),
    .C(_16013_),
    .A(_15570_),
    .Y(_16022_));
 sg13g2_a22oi_1 _46893_ (.Y(_16023_),
    .B1(_16017_),
    .B2(_16022_),
    .A2(_15637_),
    .A1(net5330));
 sg13g2_xnor2_1 _46894_ (.Y(_16024_),
    .A(_15568_),
    .B(_16023_));
 sg13g2_a21oi_1 _46895_ (.A1(net6704),
    .A2(_16024_),
    .Y(_01019_),
    .B1(_16021_));
 sg13g2_nor2_1 _46896_ (.A(net1732),
    .B(net6706),
    .Y(_16025_));
 sg13g2_nand4_1 _46897_ (.B(_15570_),
    .C(_15637_),
    .A(_16013_),
    .Y(_16026_),
    .D(_15567_));
 sg13g2_nand2b_1 _46898_ (.Y(_16027_),
    .B(net5312),
    .A_N(_15639_));
 sg13g2_inv_1 _46899_ (.Y(_16028_),
    .A(_16027_));
 sg13g2_o21ai_1 _46900_ (.B1(_16027_),
    .Y(_16029_),
    .A1(net5331),
    .A2(net1108));
 sg13g2_xnor2_1 _46901_ (.Y(_16030_),
    .A(_15564_),
    .B(_16029_));
 sg13g2_a21oi_1 _46902_ (.A1(net6706),
    .A2(_16030_),
    .Y(_01020_),
    .B1(_16025_));
 sg13g2_nand2_1 _46903_ (.Y(_16031_),
    .A(net5331),
    .B(_15563_));
 sg13g2_nor2_1 _46904_ (.A(_15564_),
    .B(net1108),
    .Y(_16032_));
 sg13g2_o21ai_1 _46905_ (.B1(_16031_),
    .Y(_16033_),
    .A1(_16028_),
    .A2(_16032_));
 sg13g2_xnor2_1 _46906_ (.Y(_16034_),
    .A(_15561_),
    .B(_16033_));
 sg13g2_mux2_1 _46907_ (.A0(net3173),
    .A1(_16034_),
    .S(net6706),
    .X(_01021_));
 sg13g2_nor2_1 _46908_ (.A(net2058),
    .B(net6711),
    .Y(_16035_));
 sg13g2_nor4_1 _46909_ (.A(net5333),
    .B(_15561_),
    .C(_15564_),
    .D(net1108),
    .Y(_16036_));
 sg13g2_nor2_1 _46910_ (.A(_15565_),
    .B(_16027_),
    .Y(_16037_));
 sg13g2_nor2_1 _46911_ (.A(_16036_),
    .B(_16037_),
    .Y(_16038_));
 sg13g2_xnor2_1 _46912_ (.Y(_16039_),
    .A(_15559_),
    .B(_16038_));
 sg13g2_a21oi_1 _46913_ (.A1(net6711),
    .A2(_16039_),
    .Y(_01022_),
    .B1(_16035_));
 sg13g2_nor2_1 _46914_ (.A(net2106),
    .B(net6711),
    .Y(_16040_));
 sg13g2_nand2_1 _46915_ (.Y(_16041_),
    .A(net5333),
    .B(_15559_));
 sg13g2_nor4_2 _46916_ (.A(_15558_),
    .B(_15561_),
    .C(_15564_),
    .Y(_16042_),
    .D(net1108));
 sg13g2_o21ai_1 _46917_ (.B1(_16041_),
    .Y(_16043_),
    .A1(_16037_),
    .A2(_16042_));
 sg13g2_xnor2_1 _46918_ (.Y(_16044_),
    .A(_15556_),
    .B(_16043_));
 sg13g2_a21oi_1 _46919_ (.A1(net6711),
    .A2(_16044_),
    .Y(_01023_),
    .B1(_16040_));
 sg13g2_nor2_1 _46920_ (.A(net2037),
    .B(net6711),
    .Y(_16045_));
 sg13g2_nand3_1 _46921_ (.B(_15556_),
    .C(_16042_),
    .A(net5361),
    .Y(_16046_));
 sg13g2_nand3b_1 _46922_ (.B(_15558_),
    .C(_16037_),
    .Y(_16047_),
    .A_N(_15556_));
 sg13g2_nand2_1 _46923_ (.Y(_16048_),
    .A(_16046_),
    .B(_16047_));
 sg13g2_xor2_1 _46924_ (.B(_16048_),
    .A(_15554_),
    .X(_16049_));
 sg13g2_a21oi_1 _46925_ (.A1(net6711),
    .A2(_16049_),
    .Y(_01024_),
    .B1(_16045_));
 sg13g2_nor2_1 _46926_ (.A(net1896),
    .B(net6711),
    .Y(_16050_));
 sg13g2_and3_1 _46927_ (.X(_16051_),
    .A(_15554_),
    .B(_15556_),
    .C(_16042_));
 sg13g2_inv_1 _46928_ (.Y(_16052_),
    .A(_16051_));
 sg13g2_a22oi_1 _46929_ (.Y(_16053_),
    .B1(_16047_),
    .B2(_16052_),
    .A2(_15554_),
    .A1(net5333));
 sg13g2_xor2_1 _46930_ (.B(_16053_),
    .A(_15552_),
    .X(_16054_));
 sg13g2_a21oi_1 _46931_ (.A1(net6711),
    .A2(_16054_),
    .Y(_01025_),
    .B1(_16050_));
 sg13g2_nand4_1 _46932_ (.B(_15554_),
    .C(_15556_),
    .A(_15552_),
    .Y(_16055_),
    .D(_16042_));
 sg13g2_a22oi_1 _46933_ (.Y(_16056_),
    .B1(_16055_),
    .B2(net5361),
    .A2(net5312),
    .A1(_15641_));
 sg13g2_xnor2_1 _46934_ (.Y(_16057_),
    .A(_15550_),
    .B(_16056_));
 sg13g2_mux2_1 _46935_ (.A0(net2648),
    .A1(_16057_),
    .S(net6715),
    .X(_01026_));
 sg13g2_nand2_1 _46936_ (.Y(_16058_),
    .A(_15550_),
    .B(_16055_));
 sg13g2_a21oi_1 _46937_ (.A1(net5361),
    .A2(_16058_),
    .Y(_16059_),
    .B1(net5312));
 sg13g2_nand2_1 _46938_ (.Y(_16060_),
    .A(_15646_),
    .B(_16059_));
 sg13g2_nor2_1 _46939_ (.A(_15646_),
    .B(_16059_),
    .Y(_16061_));
 sg13g2_nor2_1 _46940_ (.A(net6626),
    .B(_16061_),
    .Y(_16062_));
 sg13g2_a22oi_1 _46941_ (.Y(_01027_),
    .B1(_16060_),
    .B2(_16062_),
    .A2(net6626),
    .A1(_18271_));
 sg13g2_nor2_1 _46942_ (.A(net5309),
    .B(_16061_),
    .Y(_16063_));
 sg13g2_xnor2_1 _46943_ (.Y(_16064_),
    .A(_15548_),
    .B(_16063_));
 sg13g2_nand2_1 _46944_ (.Y(_16065_),
    .A(net1196),
    .B(net6626));
 sg13g2_o21ai_1 _46945_ (.B1(_16065_),
    .Y(_01028_),
    .A1(net6626),
    .A2(_16064_));
 sg13g2_nor2_1 _46946_ (.A(net1525),
    .B(net6719),
    .Y(_16066_));
 sg13g2_nand2_1 _46947_ (.Y(_16067_),
    .A(net5334),
    .B(_15548_));
 sg13g2_a221oi_1 _46948_ (.B2(_16055_),
    .C1(_15547_),
    .B1(_15550_),
    .A1(_15644_),
    .Y(_16068_),
    .A2(_15645_));
 sg13g2_o21ai_1 _46949_ (.B1(_16067_),
    .Y(_16069_),
    .A1(net5309),
    .A2(net1142));
 sg13g2_xnor2_1 _46950_ (.Y(_16070_),
    .A(_15545_),
    .B(_16069_));
 sg13g2_a21oi_1 _46951_ (.A1(net6719),
    .A2(_16070_),
    .Y(_01029_),
    .B1(_16066_));
 sg13g2_nor2_1 _46952_ (.A(net1563),
    .B(net6717),
    .Y(_16071_));
 sg13g2_and2_1 _46953_ (.A(_15545_),
    .B(net1142),
    .X(_16072_));
 sg13g2_a21oi_1 _46954_ (.A1(net5362),
    .A2(_16072_),
    .Y(_16073_),
    .B1(net5309));
 sg13g2_xnor2_1 _46955_ (.Y(_16074_),
    .A(_15543_),
    .B(_16073_));
 sg13g2_a21oi_1 _46956_ (.A1(net6717),
    .A2(_16074_),
    .Y(_01030_),
    .B1(_16071_));
 sg13g2_nor2_1 _46957_ (.A(net2313),
    .B(net6720),
    .Y(_16075_));
 sg13g2_nand2_1 _46958_ (.Y(_16076_),
    .A(_15543_),
    .B(_16072_));
 sg13g2_a22oi_1 _46959_ (.Y(_16077_),
    .B1(net5194),
    .B2(_16076_),
    .A2(_15543_),
    .A1(net5334));
 sg13g2_xor2_1 _46960_ (.B(_16077_),
    .A(_15541_),
    .X(_16078_));
 sg13g2_a21oi_1 _46961_ (.A1(net6720),
    .A2(_16078_),
    .Y(_01031_),
    .B1(_16075_));
 sg13g2_nor2_1 _46962_ (.A(net1596),
    .B(net6719),
    .Y(_16079_));
 sg13g2_and4_1 _46963_ (.A(_15541_),
    .B(_15543_),
    .C(_15545_),
    .D(net1142),
    .X(_16080_));
 sg13g2_a21oi_1 _46964_ (.A1(net5362),
    .A2(_16080_),
    .Y(_16081_),
    .B1(net5309));
 sg13g2_xnor2_1 _46965_ (.Y(_16082_),
    .A(_15539_),
    .B(_16081_));
 sg13g2_a21oi_1 _46966_ (.A1(net6719),
    .A2(_16082_),
    .Y(_01032_),
    .B1(_16079_));
 sg13g2_nor2_1 _46967_ (.A(net1986),
    .B(net6719),
    .Y(_16083_));
 sg13g2_nand2_1 _46968_ (.Y(_16084_),
    .A(net5334),
    .B(_15539_));
 sg13g2_and2_1 _46969_ (.A(_15539_),
    .B(_16080_),
    .X(_16085_));
 sg13g2_o21ai_1 _46970_ (.B1(_16084_),
    .Y(_16086_),
    .A1(net5309),
    .A2(_16085_));
 sg13g2_xnor2_1 _46971_ (.Y(_16087_),
    .A(_15537_),
    .B(_16086_));
 sg13g2_a21oi_1 _46972_ (.A1(net6719),
    .A2(_16087_),
    .Y(_01033_),
    .B1(_16083_));
 sg13g2_nor2_1 _46973_ (.A(net2040),
    .B(net6717),
    .Y(_16088_));
 sg13g2_nand3_1 _46974_ (.B(_15537_),
    .C(_16085_),
    .A(net5362),
    .Y(_16089_));
 sg13g2_nor2b_1 _46975_ (.A(net5309),
    .B_N(_16089_),
    .Y(_16090_));
 sg13g2_xnor2_1 _46976_ (.Y(_16091_),
    .A(_15535_),
    .B(_16090_));
 sg13g2_a21oi_1 _46977_ (.A1(net6717),
    .A2(_16091_),
    .Y(_01034_),
    .B1(_16088_));
 sg13g2_nor2_1 _46978_ (.A(net2219),
    .B(net6716),
    .Y(_16092_));
 sg13g2_nand2_1 _46979_ (.Y(_16093_),
    .A(net5334),
    .B(_15535_));
 sg13g2_and4_1 _46980_ (.A(_15535_),
    .B(_15537_),
    .C(_15539_),
    .D(_16080_),
    .X(_16094_));
 sg13g2_o21ai_1 _46981_ (.B1(_16093_),
    .Y(_16095_),
    .A1(net5309),
    .A2(_16094_));
 sg13g2_xnor2_1 _46982_ (.Y(_16096_),
    .A(_15533_),
    .B(_16095_));
 sg13g2_a21oi_1 _46983_ (.A1(net6716),
    .A2(_16096_),
    .Y(_01035_),
    .B1(_16092_));
 sg13g2_nor2_1 _46984_ (.A(net1994),
    .B(net6716),
    .Y(_16097_));
 sg13g2_nand2_1 _46985_ (.Y(_16098_),
    .A(_15533_),
    .B(_16094_));
 sg13g2_o21ai_1 _46986_ (.B1(net5194),
    .Y(_16099_),
    .A1(net5334),
    .A2(_16098_));
 sg13g2_xor2_1 _46987_ (.B(_16099_),
    .A(_15531_),
    .X(_16100_));
 sg13g2_a21oi_1 _46988_ (.A1(net6716),
    .A2(_16100_),
    .Y(_01036_),
    .B1(_16097_));
 sg13g2_nor2_1 _46989_ (.A(net1407),
    .B(net6716),
    .Y(_16101_));
 sg13g2_nand3_1 _46990_ (.B(_15533_),
    .C(_16094_),
    .A(_15531_),
    .Y(_16102_));
 sg13g2_a22oi_1 _46991_ (.Y(_16103_),
    .B1(net5194),
    .B2(_16102_),
    .A2(_15531_),
    .A1(net5334));
 sg13g2_xnor2_1 _46992_ (.Y(_16104_),
    .A(_15528_),
    .B(_16103_));
 sg13g2_a21oi_1 _46993_ (.A1(net6716),
    .A2(_16104_),
    .Y(_01037_),
    .B1(_16101_));
 sg13g2_nor2_1 _46994_ (.A(net2066),
    .B(net6717),
    .Y(_16105_));
 sg13g2_and4_1 _46995_ (.A(_15529_),
    .B(_15531_),
    .C(_15533_),
    .D(_16094_),
    .X(_16106_));
 sg13g2_a21oi_1 _46996_ (.A1(net5362),
    .A2(_16106_),
    .Y(_16107_),
    .B1(net5310));
 sg13g2_xnor2_1 _46997_ (.Y(_16108_),
    .A(_15526_),
    .B(_16107_));
 sg13g2_a21oi_1 _46998_ (.A1(net6718),
    .A2(_16108_),
    .Y(_01038_),
    .B1(_16105_));
 sg13g2_nor2_1 _46999_ (.A(net2210),
    .B(net6716),
    .Y(_16109_));
 sg13g2_nand2_1 _47000_ (.Y(_16110_),
    .A(net5334),
    .B(_15526_));
 sg13g2_and2_1 _47001_ (.A(_15526_),
    .B(_16106_),
    .X(_16111_));
 sg13g2_o21ai_1 _47002_ (.B1(_16110_),
    .Y(_16112_),
    .A1(net5310),
    .A2(_16111_));
 sg13g2_xnor2_1 _47003_ (.Y(_16113_),
    .A(_15524_),
    .B(_16112_));
 sg13g2_a21oi_1 _47004_ (.A1(net6716),
    .A2(_16113_),
    .Y(_01039_),
    .B1(_16109_));
 sg13g2_nor2_1 _47005_ (.A(net2217),
    .B(net6721),
    .Y(_16114_));
 sg13g2_nand3_1 _47006_ (.B(_15524_),
    .C(_16111_),
    .A(net5362),
    .Y(_16115_));
 sg13g2_nor2b_1 _47007_ (.A(net5310),
    .B_N(_16115_),
    .Y(_16116_));
 sg13g2_xnor2_1 _47008_ (.Y(_16117_),
    .A(_15518_),
    .B(_16116_));
 sg13g2_a21oi_1 _47009_ (.A1(net6721),
    .A2(_16117_),
    .Y(_01040_),
    .B1(_16114_));
 sg13g2_nor2_1 _47010_ (.A(net2379),
    .B(net6717),
    .Y(_16118_));
 sg13g2_nand2_1 _47011_ (.Y(_16119_),
    .A(net5334),
    .B(_15518_));
 sg13g2_and4_1 _47012_ (.A(_15518_),
    .B(_15524_),
    .C(_15526_),
    .D(_16106_),
    .X(_16120_));
 sg13g2_o21ai_1 _47013_ (.B1(_16119_),
    .Y(_16121_),
    .A1(net5309),
    .A2(_16120_));
 sg13g2_xnor2_1 _47014_ (.Y(_16122_),
    .A(_15516_),
    .B(_16121_));
 sg13g2_a21oi_1 _47015_ (.A1(net6718),
    .A2(_16122_),
    .Y(_01041_),
    .B1(_16118_));
 sg13g2_nor2_1 _47016_ (.A(net2237),
    .B(net6718),
    .Y(_16123_));
 sg13g2_nand2_1 _47017_ (.Y(_16124_),
    .A(_15516_),
    .B(_16120_));
 sg13g2_o21ai_1 _47018_ (.B1(net5194),
    .Y(_16125_),
    .A1(net5335),
    .A2(_16124_));
 sg13g2_xor2_1 _47019_ (.B(_16125_),
    .A(_15520_),
    .X(_16126_));
 sg13g2_a21oi_1 _47020_ (.A1(net6718),
    .A2(_16126_),
    .Y(_01042_),
    .B1(_16123_));
 sg13g2_nor2_1 _47021_ (.A(net3180),
    .B(net6724),
    .Y(_16127_));
 sg13g2_nand3_1 _47022_ (.B(_15520_),
    .C(_16120_),
    .A(_15516_),
    .Y(_16128_));
 sg13g2_a22oi_1 _47023_ (.Y(_16129_),
    .B1(net5194),
    .B2(_16128_),
    .A2(_15520_),
    .A1(net5335));
 sg13g2_xor2_1 _47024_ (.B(_16129_),
    .A(_15523_),
    .X(_16130_));
 sg13g2_a21oi_1 _47025_ (.A1(net6720),
    .A2(_16130_),
    .Y(_01043_),
    .B1(_16127_));
 sg13g2_nor2_1 _47026_ (.A(net2218),
    .B(net6721),
    .Y(_16131_));
 sg13g2_and4_1 _47027_ (.A(_15516_),
    .B(_15520_),
    .C(_15523_),
    .D(_16120_),
    .X(_16132_));
 sg13g2_a21oi_1 _47028_ (.A1(net5362),
    .A2(_16132_),
    .Y(_16133_),
    .B1(net5311));
 sg13g2_xnor2_1 _47029_ (.Y(_16134_),
    .A(_15512_),
    .B(_16133_));
 sg13g2_a21oi_1 _47030_ (.A1(net6721),
    .A2(_16134_),
    .Y(_01044_),
    .B1(_16131_));
 sg13g2_nor2_1 _47031_ (.A(net2511),
    .B(net6721),
    .Y(_16135_));
 sg13g2_nand2_1 _47032_ (.Y(_16136_),
    .A(net5335),
    .B(_15512_));
 sg13g2_and2_1 _47033_ (.A(_15512_),
    .B(_16132_),
    .X(_16137_));
 sg13g2_o21ai_1 _47034_ (.B1(_16136_),
    .Y(_16138_),
    .A1(net5311),
    .A2(_16137_));
 sg13g2_xnor2_1 _47035_ (.Y(_16139_),
    .A(_15510_),
    .B(_16138_));
 sg13g2_a21oi_1 _47036_ (.A1(net6721),
    .A2(_16139_),
    .Y(_01045_),
    .B1(_16135_));
 sg13g2_nor2_1 _47037_ (.A(net1822),
    .B(net6727),
    .Y(_16140_));
 sg13g2_nand3_1 _47038_ (.B(_15510_),
    .C(_16137_),
    .A(net5362),
    .Y(_16141_));
 sg13g2_nor2b_1 _47039_ (.A(net5311),
    .B_N(_16141_),
    .Y(_16142_));
 sg13g2_xnor2_1 _47040_ (.Y(_16143_),
    .A(_15508_),
    .B(_16142_));
 sg13g2_a21oi_1 _47041_ (.A1(net6727),
    .A2(_16143_),
    .Y(_01046_),
    .B1(_16140_));
 sg13g2_nor2_1 _47042_ (.A(net2638),
    .B(net6721),
    .Y(_16144_));
 sg13g2_nand2_1 _47043_ (.Y(_16145_),
    .A(net5335),
    .B(_15508_));
 sg13g2_and4_1 _47044_ (.A(_15508_),
    .B(_15510_),
    .C(_15512_),
    .D(_16132_),
    .X(_16146_));
 sg13g2_o21ai_1 _47045_ (.B1(_16145_),
    .Y(_16147_),
    .A1(net5311),
    .A2(_16146_));
 sg13g2_xnor2_1 _47046_ (.Y(_16148_),
    .A(_15506_),
    .B(_16147_));
 sg13g2_a21oi_1 _47047_ (.A1(net6721),
    .A2(_16148_),
    .Y(_01047_),
    .B1(_16144_));
 sg13g2_nand2_1 _47048_ (.Y(_16149_),
    .A(_15506_),
    .B(_16146_));
 sg13g2_o21ai_1 _47049_ (.B1(net5193),
    .Y(_16150_),
    .A1(net5337),
    .A2(_16149_));
 sg13g2_xor2_1 _47050_ (.B(_16150_),
    .A(_15504_),
    .X(_16151_));
 sg13g2_nand2_1 _47051_ (.Y(_16152_),
    .A(net1698),
    .B(net6635));
 sg13g2_o21ai_1 _47052_ (.B1(_16152_),
    .Y(_01048_),
    .A1(net6635),
    .A2(_16151_));
 sg13g2_nor2_1 _47053_ (.A(net2499),
    .B(net6726),
    .Y(_16153_));
 sg13g2_nand3_1 _47054_ (.B(_15506_),
    .C(_16146_),
    .A(_15504_),
    .Y(_16154_));
 sg13g2_a22oi_1 _47055_ (.Y(_16155_),
    .B1(net5193),
    .B2(_16154_),
    .A2(_15504_),
    .A1(net5337));
 sg13g2_xor2_1 _47056_ (.B(_16155_),
    .A(_15502_),
    .X(_16156_));
 sg13g2_a21oi_1 _47057_ (.A1(net6726),
    .A2(_16156_),
    .Y(_01049_),
    .B1(_16153_));
 sg13g2_nor2_1 _47058_ (.A(net2081),
    .B(net6727),
    .Y(_16157_));
 sg13g2_nand4_1 _47059_ (.B(_15504_),
    .C(_15506_),
    .A(_15502_),
    .Y(_16158_),
    .D(_16146_));
 sg13g2_nor2_1 _47060_ (.A(net5337),
    .B(_16158_),
    .Y(_16159_));
 sg13g2_nor2_1 _47061_ (.A(net5313),
    .B(_16159_),
    .Y(_16160_));
 sg13g2_xnor2_1 _47062_ (.Y(_16161_),
    .A(_15500_),
    .B(_16160_));
 sg13g2_a21oi_1 _47063_ (.A1(net6727),
    .A2(_16161_),
    .Y(_01050_),
    .B1(_16157_));
 sg13g2_nor2_1 _47064_ (.A(net2838),
    .B(net6729),
    .Y(_16162_));
 sg13g2_nand2b_1 _47065_ (.Y(_16163_),
    .B(_15500_),
    .A_N(_16158_));
 sg13g2_a22oi_1 _47066_ (.Y(_16164_),
    .B1(net5193),
    .B2(_16163_),
    .A2(_15500_),
    .A1(net5337));
 sg13g2_xnor2_1 _47067_ (.Y(_16165_),
    .A(_15497_),
    .B(_16164_));
 sg13g2_a21oi_1 _47068_ (.A1(net6729),
    .A2(_16165_),
    .Y(_01051_),
    .B1(_16162_));
 sg13g2_nor2_1 _47069_ (.A(net2873),
    .B(net6726),
    .Y(_16166_));
 sg13g2_nor3_1 _47070_ (.A(net5337),
    .B(_15497_),
    .C(_16163_),
    .Y(_16167_));
 sg13g2_nor2_1 _47071_ (.A(net5313),
    .B(_16167_),
    .Y(_16168_));
 sg13g2_xnor2_1 _47072_ (.Y(_16169_),
    .A(_15494_),
    .B(_16168_));
 sg13g2_a21oi_1 _47073_ (.A1(net6726),
    .A2(_16169_),
    .Y(_01052_),
    .B1(_16166_));
 sg13g2_nor2_1 _47074_ (.A(net2752),
    .B(net6725),
    .Y(_16170_));
 sg13g2_nor4_2 _47075_ (.A(_15495_),
    .B(_15497_),
    .C(_15499_),
    .Y(_16171_),
    .D(_16158_));
 sg13g2_nand2_1 _47076_ (.Y(_16172_),
    .A(net5337),
    .B(_15494_));
 sg13g2_o21ai_1 _47077_ (.B1(_16172_),
    .Y(_16173_),
    .A1(net5313),
    .A2(_16171_));
 sg13g2_xnor2_1 _47078_ (.Y(_16174_),
    .A(_15492_),
    .B(_16173_));
 sg13g2_a21oi_1 _47079_ (.A1(net6725),
    .A2(_16174_),
    .Y(_01053_),
    .B1(_16170_));
 sg13g2_nor2_1 _47080_ (.A(net2068),
    .B(net6725),
    .Y(_16175_));
 sg13g2_nand2_1 _47081_ (.Y(_16176_),
    .A(_15492_),
    .B(_16171_));
 sg13g2_o21ai_1 _47082_ (.B1(net5193),
    .Y(_16177_),
    .A1(net5340),
    .A2(_16176_));
 sg13g2_xor2_1 _47083_ (.B(_16177_),
    .A(_15490_),
    .X(_16178_));
 sg13g2_a21oi_1 _47084_ (.A1(net6725),
    .A2(_16178_),
    .Y(_01054_),
    .B1(_16175_));
 sg13g2_nand3_1 _47085_ (.B(_15492_),
    .C(_16171_),
    .A(_15490_),
    .Y(_16179_));
 sg13g2_a22oi_1 _47086_ (.Y(_16180_),
    .B1(net5193),
    .B2(_16179_),
    .A2(_15490_),
    .A1(net5337));
 sg13g2_xnor2_1 _47087_ (.Y(_16181_),
    .A(_15488_),
    .B(_16180_));
 sg13g2_mux2_1 _47088_ (.A0(net3490),
    .A1(_16181_),
    .S(net6725),
    .X(_01055_));
 sg13g2_nor2_1 _47089_ (.A(net2566),
    .B(net6725),
    .Y(_16182_));
 sg13g2_and4_1 _47090_ (.A(_15488_),
    .B(_15490_),
    .C(_15492_),
    .D(_16171_),
    .X(_16183_));
 sg13g2_a21oi_1 _47091_ (.A1(net5368),
    .A2(_16183_),
    .Y(_16184_),
    .B1(net5313));
 sg13g2_xnor2_1 _47092_ (.Y(_16185_),
    .A(_15486_),
    .B(_16184_));
 sg13g2_a21oi_1 _47093_ (.A1(net6725),
    .A2(_16185_),
    .Y(_01056_),
    .B1(_16182_));
 sg13g2_nor2_1 _47094_ (.A(net2558),
    .B(net6725),
    .Y(_16186_));
 sg13g2_nand2_1 _47095_ (.Y(_16187_),
    .A(net5337),
    .B(_15486_));
 sg13g2_and2_1 _47096_ (.A(_15486_),
    .B(_16183_),
    .X(_16188_));
 sg13g2_o21ai_1 _47097_ (.B1(_16187_),
    .Y(_16189_),
    .A1(net5313),
    .A2(_16188_));
 sg13g2_xnor2_1 _47098_ (.Y(_16190_),
    .A(_15484_),
    .B(_16189_));
 sg13g2_a21oi_1 _47099_ (.A1(net6726),
    .A2(_16190_),
    .Y(_01057_),
    .B1(_16186_));
 sg13g2_nor2_1 _47100_ (.A(net3189),
    .B(net6739),
    .Y(_16191_));
 sg13g2_and3_1 _47101_ (.X(_16192_),
    .A(net5368),
    .B(_15484_),
    .C(_16188_));
 sg13g2_nor2_1 _47102_ (.A(net5313),
    .B(_16192_),
    .Y(_16193_));
 sg13g2_xnor2_1 _47103_ (.Y(_16194_),
    .A(_15482_),
    .B(_16193_));
 sg13g2_a21oi_1 _47104_ (.A1(net6736),
    .A2(_16194_),
    .Y(_01058_),
    .B1(_16191_));
 sg13g2_and4_1 _47105_ (.A(_15482_),
    .B(_15484_),
    .C(_15486_),
    .D(_16183_),
    .X(_16195_));
 sg13g2_and2_1 _47106_ (.A(_15660_),
    .B(_16195_),
    .X(_16196_));
 sg13g2_nor2_1 _47107_ (.A(net5342),
    .B(_16196_),
    .Y(_16197_));
 sg13g2_or2_1 _47108_ (.X(_16198_),
    .B(_16195_),
    .A(_15660_));
 sg13g2_a221oi_1 _47109_ (.B2(_16198_),
    .C1(net6630),
    .B1(_16197_),
    .A1(net5342),
    .Y(_16199_),
    .A2(_15660_));
 sg13g2_a22oi_1 _47110_ (.Y(_16200_),
    .B1(net5193),
    .B2(_16199_),
    .A2(net6632),
    .A1(net2711));
 sg13g2_inv_1 _47111_ (.Y(_01059_),
    .A(_16200_));
 sg13g2_nor2_1 _47112_ (.A(net5187),
    .B(_16197_),
    .Y(_16201_));
 sg13g2_xnor2_1 _47113_ (.Y(_16202_),
    .A(_15662_),
    .B(_16201_));
 sg13g2_mux2_1 _47114_ (.A0(net2859),
    .A1(_16202_),
    .S(net6743),
    .X(_01060_));
 sg13g2_nor2_1 _47115_ (.A(net2250),
    .B(net6743),
    .Y(_16203_));
 sg13g2_nand2_1 _47116_ (.Y(_16204_),
    .A(_15662_),
    .B(_16196_));
 sg13g2_nor2_1 _47117_ (.A(net5342),
    .B(_16204_),
    .Y(_16205_));
 sg13g2_nor2_1 _47118_ (.A(net5313),
    .B(_16205_),
    .Y(_16206_));
 sg13g2_xnor2_1 _47119_ (.Y(_16207_),
    .A(_15480_),
    .B(_16206_));
 sg13g2_a21oi_1 _47120_ (.A1(net6743),
    .A2(_16207_),
    .Y(_01061_),
    .B1(_16203_));
 sg13g2_nor2b_1 _47121_ (.A(_16204_),
    .B_N(_15480_),
    .Y(_16208_));
 sg13g2_nand4_1 _47122_ (.B(_15660_),
    .C(_15662_),
    .A(_15480_),
    .Y(_16209_),
    .D(_16195_));
 sg13g2_o21ai_1 _47123_ (.B1(net5174),
    .Y(_16210_),
    .A1(net5341),
    .A2(_16208_));
 sg13g2_xnor2_1 _47124_ (.Y(_16211_),
    .A(_15477_),
    .B(_16210_));
 sg13g2_nand2_1 _47125_ (.Y(_16212_),
    .A(net1360),
    .B(net6632));
 sg13g2_o21ai_1 _47126_ (.B1(_16212_),
    .Y(_01062_),
    .A1(net6632),
    .A2(_16211_));
 sg13g2_nand2_1 _47127_ (.Y(_16213_),
    .A(_15475_),
    .B(net5193));
 sg13g2_nand2_1 _47128_ (.Y(_16214_),
    .A(_15477_),
    .B(_16208_));
 sg13g2_nor2_1 _47129_ (.A(_15475_),
    .B(_16214_),
    .Y(_16215_));
 sg13g2_nor2_1 _47130_ (.A(net5341),
    .B(_16215_),
    .Y(_16216_));
 sg13g2_nand2_1 _47131_ (.Y(_16217_),
    .A(_15475_),
    .B(_16214_));
 sg13g2_a221oi_1 _47132_ (.B2(_16217_),
    .C1(net6631),
    .B1(_16216_),
    .A1(net5341),
    .Y(_16218_),
    .A2(_16213_));
 sg13g2_a21o_1 _47133_ (.A2(net6630),
    .A1(net3057),
    .B1(_16218_),
    .X(_01063_));
 sg13g2_nor2_1 _47134_ (.A(net1923),
    .B(net6743),
    .Y(_16219_));
 sg13g2_nor2_1 _47135_ (.A(net5188),
    .B(_16216_),
    .Y(_16220_));
 sg13g2_xnor2_1 _47136_ (.Y(_16221_),
    .A(_15473_),
    .B(_16220_));
 sg13g2_a21oi_1 _47137_ (.A1(net6743),
    .A2(_16221_),
    .Y(_01064_),
    .B1(_16219_));
 sg13g2_nor2_1 _47138_ (.A(net2630),
    .B(net6740),
    .Y(_16222_));
 sg13g2_xnor2_1 _47139_ (.Y(_16223_),
    .A(net5366),
    .B(_15473_));
 sg13g2_nor3_1 _47140_ (.A(net5188),
    .B(_16216_),
    .C(_16223_),
    .Y(_16224_));
 sg13g2_xor2_1 _47141_ (.B(_16224_),
    .A(_15470_),
    .X(_16225_));
 sg13g2_a21oi_1 _47142_ (.A1(net6740),
    .A2(_16225_),
    .Y(_01065_),
    .B1(_16222_));
 sg13g2_nor2_1 _47143_ (.A(net1406),
    .B(net6743),
    .Y(_16226_));
 sg13g2_nand2_1 _47144_ (.Y(_16227_),
    .A(_15470_),
    .B(_15472_));
 sg13g2_nor4_2 _47145_ (.A(_15475_),
    .B(_15478_),
    .C(_16209_),
    .Y(_16228_),
    .D(_16227_));
 sg13g2_a21oi_1 _47146_ (.A1(net5366),
    .A2(_16228_),
    .Y(_16229_),
    .B1(net5313));
 sg13g2_xnor2_1 _47147_ (.Y(_16230_),
    .A(_15468_),
    .B(_16229_));
 sg13g2_a21oi_1 _47148_ (.A1(net6743),
    .A2(_16230_),
    .Y(_01066_),
    .B1(_16226_));
 sg13g2_o21ai_1 _47149_ (.B1(net5341),
    .Y(_16231_),
    .A1(_15466_),
    .A2(net1140));
 sg13g2_a21oi_1 _47150_ (.A1(_15468_),
    .A2(_16228_),
    .Y(_16232_),
    .B1(_15466_));
 sg13g2_and3_1 _47151_ (.X(_16233_),
    .A(_15466_),
    .B(_15468_),
    .C(_16228_));
 sg13g2_nand2b_1 _47152_ (.Y(_16234_),
    .B(net5367),
    .A_N(_16233_));
 sg13g2_nor2_1 _47153_ (.A(_16232_),
    .B(_16234_),
    .Y(_16235_));
 sg13g2_nor2_1 _47154_ (.A(net6631),
    .B(_16235_),
    .Y(_16236_));
 sg13g2_a22oi_1 _47155_ (.Y(_16237_),
    .B1(_16231_),
    .B2(_16236_),
    .A2(net6630),
    .A1(net3174));
 sg13g2_inv_1 _47156_ (.Y(_01067_),
    .A(_16237_));
 sg13g2_nor2_1 _47157_ (.A(net2373),
    .B(net6740),
    .Y(_16238_));
 sg13g2_nand2_1 _47158_ (.Y(_16239_),
    .A(net5174),
    .B(_16234_));
 sg13g2_xnor2_1 _47159_ (.Y(_16240_),
    .A(_15464_),
    .B(_16239_));
 sg13g2_a21oi_1 _47160_ (.A1(net6740),
    .A2(_16240_),
    .Y(_01068_),
    .B1(_16238_));
 sg13g2_nor2_1 _47161_ (.A(net2161),
    .B(net6740),
    .Y(_16241_));
 sg13g2_nand4_1 _47162_ (.B(_15466_),
    .C(_15468_),
    .A(_15464_),
    .Y(_16242_),
    .D(_16228_));
 sg13g2_nor2_1 _47163_ (.A(net5341),
    .B(_16242_),
    .Y(_16243_));
 sg13g2_nor2_1 _47164_ (.A(net1140),
    .B(_16243_),
    .Y(_16244_));
 sg13g2_xnor2_1 _47165_ (.Y(_16245_),
    .A(_15461_),
    .B(_16244_));
 sg13g2_a21oi_1 _47166_ (.A1(net6740),
    .A2(_16245_),
    .Y(_01069_),
    .B1(_16241_));
 sg13g2_nor2_1 _47167_ (.A(_15462_),
    .B(_16242_),
    .Y(_16246_));
 sg13g2_o21ai_1 _47168_ (.B1(net5176),
    .Y(_16247_),
    .A1(net5341),
    .A2(_16246_));
 sg13g2_xnor2_1 _47169_ (.Y(_16248_),
    .A(_15458_),
    .B(_16247_));
 sg13g2_nand2_1 _47170_ (.Y(_16249_),
    .A(net1207),
    .B(net6630));
 sg13g2_o21ai_1 _47171_ (.B1(_16249_),
    .Y(_01070_),
    .A1(net6630),
    .A2(_16248_));
 sg13g2_nand2_1 _47172_ (.Y(_16250_),
    .A(_15458_),
    .B(_16246_));
 sg13g2_nor4_2 _47173_ (.A(_15456_),
    .B(_15459_),
    .C(_15462_),
    .Y(_16251_),
    .D(_16242_));
 sg13g2_xnor2_1 _47174_ (.Y(_16252_),
    .A(_15456_),
    .B(_16250_));
 sg13g2_a221oi_1 _47175_ (.B2(net5367),
    .C1(net6630),
    .B1(_16252_),
    .A1(_15456_),
    .Y(_16253_),
    .A2(net5188));
 sg13g2_a21oi_1 _47176_ (.A1(_18272_),
    .A2(net6632),
    .Y(_01071_),
    .B1(_16253_));
 sg13g2_nor2_1 _47177_ (.A(net5341),
    .B(_16251_),
    .Y(_16254_));
 sg13g2_nor2_1 _47178_ (.A(net5188),
    .B(_16254_),
    .Y(_16255_));
 sg13g2_xor2_1 _47179_ (.B(_16255_),
    .A(_15451_),
    .X(_16256_));
 sg13g2_nor2_1 _47180_ (.A(net1627),
    .B(net6740),
    .Y(_16257_));
 sg13g2_a21oi_1 _47181_ (.A1(net6740),
    .A2(_16256_),
    .Y(_01072_),
    .B1(_16257_));
 sg13g2_nor2_1 _47182_ (.A(net1991),
    .B(net6741),
    .Y(_16258_));
 sg13g2_xnor2_1 _47183_ (.Y(_16259_),
    .A(net5367),
    .B(_15451_));
 sg13g2_nand2_1 _47184_ (.Y(_16260_),
    .A(_16255_),
    .B(_16259_));
 sg13g2_xnor2_1 _47185_ (.Y(_16261_),
    .A(_15453_),
    .B(_16260_));
 sg13g2_a21oi_1 _47186_ (.A1(net6741),
    .A2(_16261_),
    .Y(_01073_),
    .B1(_16258_));
 sg13g2_nor2_1 _47187_ (.A(net2135),
    .B(net6741),
    .Y(_16262_));
 sg13g2_and2_1 _47188_ (.A(_15451_),
    .B(_15453_),
    .X(_16263_));
 sg13g2_nand2_1 _47189_ (.Y(_16264_),
    .A(_16251_),
    .B(_16263_));
 sg13g2_a21oi_1 _47190_ (.A1(net5367),
    .A2(_16264_),
    .Y(_16265_),
    .B1(net5188));
 sg13g2_xnor2_1 _47191_ (.Y(_16266_),
    .A(_15447_),
    .B(_16265_));
 sg13g2_a21oi_1 _47192_ (.A1(net6741),
    .A2(_16266_),
    .Y(_01074_),
    .B1(_16262_));
 sg13g2_nand2_1 _47193_ (.Y(_16267_),
    .A(_15455_),
    .B(net5194));
 sg13g2_nor2_1 _47194_ (.A(_15447_),
    .B(_15455_),
    .Y(_16268_));
 sg13g2_nor2b_1 _47195_ (.A(_16264_),
    .B_N(_16268_),
    .Y(_16269_));
 sg13g2_nor2_1 _47196_ (.A(net5341),
    .B(_16269_),
    .Y(_16270_));
 sg13g2_o21ai_1 _47197_ (.B1(_15455_),
    .Y(_16271_),
    .A1(_15447_),
    .A2(_16264_));
 sg13g2_a221oi_1 _47198_ (.B2(_16271_),
    .C1(net6630),
    .B1(_16270_),
    .A1(net5342),
    .Y(_16272_),
    .A2(_16267_));
 sg13g2_a21o_1 _47199_ (.A2(net6630),
    .A1(net2936),
    .B1(_16272_),
    .X(_01075_));
 sg13g2_nor2_1 _47200_ (.A(net2046),
    .B(net6742),
    .Y(_16273_));
 sg13g2_nor2_1 _47201_ (.A(net5187),
    .B(_16270_),
    .Y(_16274_));
 sg13g2_xnor2_1 _47202_ (.Y(_16275_),
    .A(_15444_),
    .B(_16274_));
 sg13g2_a21oi_1 _47203_ (.A1(net6742),
    .A2(_16275_),
    .Y(_01076_),
    .B1(_16273_));
 sg13g2_nand4_1 _47204_ (.B(_15443_),
    .C(_16263_),
    .A(_16251_),
    .Y(_16276_),
    .D(_16268_));
 sg13g2_nor2_1 _47205_ (.A(_15441_),
    .B(net1101),
    .Y(_16277_));
 sg13g2_xnor2_1 _47206_ (.Y(_16278_),
    .A(_15441_),
    .B(net1101));
 sg13g2_a221oi_1 _47207_ (.B2(net5367),
    .C1(net6631),
    .B1(_16278_),
    .A1(_15441_),
    .Y(_16279_),
    .A2(net5188));
 sg13g2_a21oi_1 _47208_ (.A1(_18273_),
    .A2(net6631),
    .Y(_01077_),
    .B1(_16279_));
 sg13g2_nor2_1 _47209_ (.A(net2131),
    .B(net6737),
    .Y(_16280_));
 sg13g2_o21ai_1 _47210_ (.B1(net5174),
    .Y(_16281_),
    .A1(net5343),
    .A2(_16277_));
 sg13g2_xnor2_1 _47211_ (.Y(_16282_),
    .A(_15435_),
    .B(_16281_));
 sg13g2_a21oi_1 _47212_ (.A1(net6737),
    .A2(_16282_),
    .Y(_01078_),
    .B1(_16280_));
 sg13g2_nand2_1 _47213_ (.Y(_16283_),
    .A(_15433_),
    .B(_15435_));
 sg13g2_nor3_2 _47214_ (.A(_15441_),
    .B(net1101),
    .C(_16283_),
    .Y(_16284_));
 sg13g2_nor2_1 _47215_ (.A(_15436_),
    .B(_16284_),
    .Y(_16285_));
 sg13g2_o21ai_1 _47216_ (.B1(_16285_),
    .Y(_16286_),
    .A1(_15433_),
    .A2(_16277_));
 sg13g2_a21oi_1 _47217_ (.A1(net5366),
    .A2(_16286_),
    .Y(_16287_),
    .B1(net6631));
 sg13g2_o21ai_1 _47218_ (.B1(_16287_),
    .Y(_16288_),
    .A1(_15433_),
    .A2(net5174));
 sg13g2_o21ai_1 _47219_ (.B1(_16288_),
    .Y(_16289_),
    .A1(net3316),
    .A2(net6737));
 sg13g2_inv_1 _47220_ (.Y(_01079_),
    .A(_16289_));
 sg13g2_nor2_1 _47221_ (.A(net2449),
    .B(net6737),
    .Y(_16290_));
 sg13g2_o21ai_1 _47222_ (.B1(net5174),
    .Y(_16291_),
    .A1(net5343),
    .A2(_16284_));
 sg13g2_xnor2_1 _47223_ (.Y(_16292_),
    .A(_15431_),
    .B(_16291_));
 sg13g2_a21oi_1 _47224_ (.A1(net6737),
    .A2(_16292_),
    .Y(_01080_),
    .B1(_16290_));
 sg13g2_nor2_1 _47225_ (.A(net2315),
    .B(net6737),
    .Y(_16293_));
 sg13g2_xnor2_1 _47226_ (.Y(_16294_),
    .A(net5343),
    .B(_15431_));
 sg13g2_nor2_1 _47227_ (.A(_16291_),
    .B(_16294_),
    .Y(_16295_));
 sg13g2_xnor2_1 _47228_ (.Y(_16296_),
    .A(_15429_),
    .B(_16295_));
 sg13g2_a21oi_1 _47229_ (.A1(net6737),
    .A2(_16296_),
    .Y(_01081_),
    .B1(_16293_));
 sg13g2_nor2b_1 _47230_ (.A(_15429_),
    .B_N(_15431_),
    .Y(_16297_));
 sg13g2_nand2_1 _47231_ (.Y(_16298_),
    .A(_16284_),
    .B(_16297_));
 sg13g2_a21oi_1 _47232_ (.A1(net5366),
    .A2(_16298_),
    .Y(_16299_),
    .B1(net5187));
 sg13g2_xnor2_1 _47233_ (.Y(_16300_),
    .A(_15426_),
    .B(_16299_));
 sg13g2_nand2_1 _47234_ (.Y(_16301_),
    .A(net1240),
    .B(net6631));
 sg13g2_o21ai_1 _47235_ (.B1(_16301_),
    .Y(_01082_),
    .A1(net6633),
    .A2(_16300_));
 sg13g2_nor2_1 _47236_ (.A(net2644),
    .B(net6742),
    .Y(_16302_));
 sg13g2_nor3_1 _47237_ (.A(_15426_),
    .B(_15673_),
    .C(_16298_),
    .Y(_16303_));
 sg13g2_nand4_1 _47238_ (.B(_15672_),
    .C(_16284_),
    .A(_15427_),
    .Y(_16304_),
    .D(_16297_));
 sg13g2_o21ai_1 _47239_ (.B1(_15673_),
    .Y(_16305_),
    .A1(_15426_),
    .A2(_16298_));
 sg13g2_nand2_1 _47240_ (.Y(_16306_),
    .A(_16304_),
    .B(_16305_));
 sg13g2_a22oi_1 _47241_ (.Y(_16307_),
    .B1(_16306_),
    .B2(net5366),
    .A2(net5187),
    .A1(_15673_));
 sg13g2_a21oi_1 _47242_ (.A1(net6738),
    .A2(_16307_),
    .Y(_01083_),
    .B1(_16302_));
 sg13g2_nor2_1 _47243_ (.A(net1566),
    .B(net6738),
    .Y(_16308_));
 sg13g2_o21ai_1 _47244_ (.B1(net5174),
    .Y(_16309_),
    .A1(net5343),
    .A2(_16303_));
 sg13g2_xnor2_1 _47245_ (.Y(_16310_),
    .A(_15675_),
    .B(_16309_));
 sg13g2_a21oi_1 _47246_ (.A1(net6738),
    .A2(_16310_),
    .Y(_01084_),
    .B1(_16308_));
 sg13g2_nand2_1 _47247_ (.Y(_16311_),
    .A(_15675_),
    .B(_16303_));
 sg13g2_nand3b_1 _47248_ (.B(_15675_),
    .C(_15424_),
    .Y(_16312_),
    .A_N(_16304_));
 sg13g2_xor2_1 _47249_ (.B(_16311_),
    .A(_15424_),
    .X(_16313_));
 sg13g2_a21oi_1 _47250_ (.A1(net5366),
    .A2(_16313_),
    .Y(_16314_),
    .B1(net6633));
 sg13g2_o21ai_1 _47251_ (.B1(_16314_),
    .Y(_16315_),
    .A1(_15424_),
    .A2(net5174));
 sg13g2_o21ai_1 _47252_ (.B1(_16315_),
    .Y(_16316_),
    .A1(net3370),
    .A2(net6739));
 sg13g2_inv_1 _47253_ (.Y(_01085_),
    .A(_16316_));
 sg13g2_a21oi_1 _47254_ (.A1(net5366),
    .A2(_16312_),
    .Y(_16317_),
    .B1(net5187));
 sg13g2_xnor2_1 _47255_ (.Y(_16318_),
    .A(_15422_),
    .B(_16317_));
 sg13g2_nand2_1 _47256_ (.Y(_16319_),
    .A(net1208),
    .B(net6631));
 sg13g2_o21ai_1 _47257_ (.B1(_16319_),
    .Y(_01086_),
    .A1(net6633),
    .A2(_16318_));
 sg13g2_nor3_1 _47258_ (.A(_15422_),
    .B(_15679_),
    .C(_16312_),
    .Y(_16320_));
 sg13g2_o21ai_1 _47259_ (.B1(_15679_),
    .Y(_16321_),
    .A1(_15422_),
    .A2(_16312_));
 sg13g2_nand2b_1 _47260_ (.Y(_16322_),
    .B(_16321_),
    .A_N(_16320_));
 sg13g2_a221oi_1 _47261_ (.B2(net5366),
    .C1(net6633),
    .B1(_16322_),
    .A1(_15679_),
    .Y(_16323_),
    .A2(net5187));
 sg13g2_a21oi_1 _47262_ (.A1(_18274_),
    .A2(net6633),
    .Y(_01087_),
    .B1(_16323_));
 sg13g2_o21ai_1 _47263_ (.B1(net5174),
    .Y(_16324_),
    .A1(net5343),
    .A2(_16320_));
 sg13g2_xnor2_1 _47264_ (.Y(_16325_),
    .A(_15421_),
    .B(_16324_));
 sg13g2_nor2_1 _47265_ (.A(net1645),
    .B(net6738),
    .Y(_16326_));
 sg13g2_a21oi_1 _47266_ (.A1(net6738),
    .A2(_16325_),
    .Y(_01088_),
    .B1(_16326_));
 sg13g2_nor2_1 _47267_ (.A(net2162),
    .B(net6737),
    .Y(_16327_));
 sg13g2_xnor2_1 _47268_ (.Y(_16328_),
    .A(net5343),
    .B(_15421_));
 sg13g2_nor2_1 _47269_ (.A(_16324_),
    .B(_16328_),
    .Y(_16329_));
 sg13g2_xnor2_1 _47270_ (.Y(_16330_),
    .A(_15403_),
    .B(_16329_));
 sg13g2_a21oi_1 _47271_ (.A1(net6739),
    .A2(_16330_),
    .Y(_01089_),
    .B1(_16327_));
 sg13g2_nor2_1 _47272_ (.A(net2061),
    .B(net6730),
    .Y(_16331_));
 sg13g2_nand2b_1 _47273_ (.Y(_16332_),
    .B(_15421_),
    .A_N(_15403_));
 sg13g2_nor4_2 _47274_ (.A(_15422_),
    .B(_15679_),
    .C(_16312_),
    .Y(_16333_),
    .D(_16332_));
 sg13g2_o21ai_1 _47275_ (.B1(net5175),
    .Y(_16334_),
    .A1(net5338),
    .A2(_16333_));
 sg13g2_xnor2_1 _47276_ (.Y(_16335_),
    .A(_15677_),
    .B(_16334_));
 sg13g2_a21oi_1 _47277_ (.A1(net6730),
    .A2(_16335_),
    .Y(_01090_),
    .B1(_16331_));
 sg13g2_nor2_1 _47278_ (.A(net2258),
    .B(net6731),
    .Y(_16336_));
 sg13g2_nand3_1 _47279_ (.B(_15677_),
    .C(_16333_),
    .A(_15410_),
    .Y(_16337_));
 sg13g2_a21o_1 _47280_ (.A2(_16333_),
    .A1(_15677_),
    .B1(_15410_),
    .X(_16338_));
 sg13g2_nand2_1 _47281_ (.Y(_16339_),
    .A(_16337_),
    .B(_16338_));
 sg13g2_a22oi_1 _47282_ (.Y(_16340_),
    .B1(_16339_),
    .B2(net5364),
    .A2(net5187),
    .A1(_15409_));
 sg13g2_a21oi_1 _47283_ (.A1(net6730),
    .A2(_16340_),
    .Y(_01091_),
    .B1(_16336_));
 sg13g2_a21oi_1 _47284_ (.A1(net5364),
    .A2(_16337_),
    .Y(_16341_),
    .B1(net5185));
 sg13g2_xnor2_1 _47285_ (.Y(_16342_),
    .A(_15407_),
    .B(_16341_));
 sg13g2_nand2_1 _47286_ (.Y(_16343_),
    .A(net1202),
    .B(net6628));
 sg13g2_o21ai_1 _47287_ (.B1(_16343_),
    .Y(_01092_),
    .A1(net6628),
    .A2(_16342_));
 sg13g2_nor2_1 _47288_ (.A(net1721),
    .B(net6730),
    .Y(_16344_));
 sg13g2_or3_1 _47289_ (.A(_15407_),
    .B(_15682_),
    .C(_16337_),
    .X(_16345_));
 sg13g2_o21ai_1 _47290_ (.B1(_15682_),
    .Y(_16346_),
    .A1(_15407_),
    .A2(_16337_));
 sg13g2_nand2_1 _47291_ (.Y(_16347_),
    .A(_16345_),
    .B(_16346_));
 sg13g2_a22oi_1 _47292_ (.Y(_16348_),
    .B1(_16347_),
    .B2(net5364),
    .A2(net5185),
    .A1(_15682_));
 sg13g2_a21oi_1 _47293_ (.A1(net6730),
    .A2(_16348_),
    .Y(_01093_),
    .B1(_16344_));
 sg13g2_nor2_1 _47294_ (.A(net2544),
    .B(net6730),
    .Y(_16349_));
 sg13g2_a21oi_1 _47295_ (.A1(net5364),
    .A2(_16345_),
    .Y(_16350_),
    .B1(net5185));
 sg13g2_xnor2_1 _47296_ (.Y(_16351_),
    .A(_15393_),
    .B(_16350_));
 sg13g2_a21oi_1 _47297_ (.A1(net6730),
    .A2(_16351_),
    .Y(_01094_),
    .B1(_16349_));
 sg13g2_nor4_1 _47298_ (.A(_15393_),
    .B(_15407_),
    .C(_15409_),
    .D(_15678_),
    .Y(_16352_));
 sg13g2_nor2_1 _47299_ (.A(_15395_),
    .B(_15682_),
    .Y(_16353_));
 sg13g2_and3_2 _47300_ (.X(_16354_),
    .A(_16333_),
    .B(_16352_),
    .C(_16353_));
 sg13g2_o21ai_1 _47301_ (.B1(_15395_),
    .Y(_16355_),
    .A1(_15393_),
    .A2(_16345_));
 sg13g2_nand2b_1 _47302_ (.Y(_16356_),
    .B(_16355_),
    .A_N(_16354_));
 sg13g2_a221oi_1 _47303_ (.B2(net5364),
    .C1(net6634),
    .B1(_16356_),
    .A1(_15395_),
    .Y(_16357_),
    .A2(net5187));
 sg13g2_a21oi_1 _47304_ (.A1(_18275_),
    .A2(net6634),
    .Y(_01095_),
    .B1(_16357_));
 sg13g2_o21ai_1 _47305_ (.B1(net5175),
    .Y(_16358_),
    .A1(net5338),
    .A2(_16354_));
 sg13g2_xnor2_1 _47306_ (.Y(_16359_),
    .A(_15683_),
    .B(_16358_));
 sg13g2_nand2_1 _47307_ (.Y(_16360_),
    .A(net1244),
    .B(net6634));
 sg13g2_o21ai_1 _47308_ (.B1(_16360_),
    .Y(_01096_),
    .A1(net6634),
    .A2(_16359_));
 sg13g2_nor2_1 _47309_ (.A(net1752),
    .B(net6730),
    .Y(_16361_));
 sg13g2_xnor2_1 _47310_ (.Y(_16362_),
    .A(net5338),
    .B(_15683_));
 sg13g2_nor2_1 _47311_ (.A(_16358_),
    .B(_16362_),
    .Y(_16363_));
 sg13g2_xnor2_1 _47312_ (.Y(_16364_),
    .A(_15391_),
    .B(_16363_));
 sg13g2_a21oi_1 _47313_ (.A1(net6731),
    .A2(_16364_),
    .Y(_01097_),
    .B1(_16361_));
 sg13g2_nand2b_1 _47314_ (.Y(_16365_),
    .B(_15683_),
    .A_N(_15391_));
 sg13g2_inv_1 _47315_ (.Y(_16366_),
    .A(_16365_));
 sg13g2_nand2_1 _47316_ (.Y(_16367_),
    .A(_16354_),
    .B(_16366_));
 sg13g2_a21oi_1 _47317_ (.A1(net5364),
    .A2(_16367_),
    .Y(_16368_),
    .B1(net5186));
 sg13g2_xnor2_1 _47318_ (.Y(_16369_),
    .A(_15397_),
    .B(_16368_));
 sg13g2_nand2_1 _47319_ (.Y(_16370_),
    .A(net1209),
    .B(net6628));
 sg13g2_o21ai_1 _47320_ (.B1(_16370_),
    .Y(_01098_),
    .A1(net6628),
    .A2(_16369_));
 sg13g2_nor2_1 _47321_ (.A(net2390),
    .B(net6731),
    .Y(_16371_));
 sg13g2_nand4_1 _47322_ (.B(_15418_),
    .C(_16354_),
    .A(_15398_),
    .Y(_16372_),
    .D(_16366_));
 sg13g2_o21ai_1 _47323_ (.B1(_15419_),
    .Y(_16373_),
    .A1(_15397_),
    .A2(_16367_));
 sg13g2_nand2_1 _47324_ (.Y(_16374_),
    .A(_16372_),
    .B(_16373_));
 sg13g2_a22oi_1 _47325_ (.Y(_16375_),
    .B1(_16374_),
    .B2(net5364),
    .A2(net5185),
    .A1(_15419_));
 sg13g2_a21oi_1 _47326_ (.A1(net6734),
    .A2(_16375_),
    .Y(_01099_),
    .B1(_16371_));
 sg13g2_nor2_1 _47327_ (.A(net1995),
    .B(net6731),
    .Y(_16376_));
 sg13g2_a21oi_1 _47328_ (.A1(net5363),
    .A2(_16372_),
    .Y(_16377_),
    .B1(net5185));
 sg13g2_xnor2_1 _47329_ (.Y(_16378_),
    .A(_15416_),
    .B(_16377_));
 sg13g2_a21oi_1 _47330_ (.A1(net6731),
    .A2(_16378_),
    .Y(_01100_),
    .B1(_16376_));
 sg13g2_nor3_1 _47331_ (.A(_15388_),
    .B(_15416_),
    .C(_16372_),
    .Y(_16379_));
 sg13g2_o21ai_1 _47332_ (.B1(_15388_),
    .Y(_16380_),
    .A1(_15416_),
    .A2(_16372_));
 sg13g2_nand2b_1 _47333_ (.Y(_16381_),
    .B(_16380_),
    .A_N(_16379_));
 sg13g2_a221oi_1 _47334_ (.B2(net5363),
    .C1(net6627),
    .B1(_16381_),
    .A1(_15388_),
    .Y(_16382_),
    .A2(net5185));
 sg13g2_a21oi_1 _47335_ (.A1(_18276_),
    .A2(net6628),
    .Y(_01101_),
    .B1(_16382_));
 sg13g2_nor2_1 _47336_ (.A(net1607),
    .B(net6733),
    .Y(_16383_));
 sg13g2_o21ai_1 _47337_ (.B1(net5175),
    .Y(_16384_),
    .A1(net5338),
    .A2(_16379_));
 sg13g2_xnor2_1 _47338_ (.Y(_16385_),
    .A(_15386_),
    .B(_16384_));
 sg13g2_a21oi_1 _47339_ (.A1(net6733),
    .A2(_16385_),
    .Y(_01102_),
    .B1(_16383_));
 sg13g2_nand2_1 _47340_ (.Y(_16386_),
    .A(_15386_),
    .B(_16379_));
 sg13g2_or2_1 _47341_ (.X(_16387_),
    .B(_16386_),
    .A(_15385_));
 sg13g2_xnor2_1 _47342_ (.Y(_16388_),
    .A(_15385_),
    .B(_16386_));
 sg13g2_a221oi_1 _47343_ (.B2(net5363),
    .C1(net6628),
    .B1(_16388_),
    .A1(_15385_),
    .Y(_16389_),
    .A2(net5186));
 sg13g2_a21oi_1 _47344_ (.A1(_18277_),
    .A2(net6628),
    .Y(_01103_),
    .B1(_16389_));
 sg13g2_nor2_1 _47345_ (.A(net1837),
    .B(net6734),
    .Y(_16390_));
 sg13g2_a21oi_2 _47346_ (.B1(net5186),
    .Y(_16391_),
    .A2(_16387_),
    .A1(net5365));
 sg13g2_xnor2_1 _47347_ (.Y(_16392_),
    .A(_15691_),
    .B(_16391_));
 sg13g2_a21oi_1 _47348_ (.A1(net6734),
    .A2(_16392_),
    .Y(_01104_),
    .B1(_16390_));
 sg13g2_nor2_1 _47349_ (.A(net1944),
    .B(net6734),
    .Y(_16393_));
 sg13g2_xnor2_1 _47350_ (.Y(_16394_),
    .A(net5339),
    .B(_15691_));
 sg13g2_nand2_1 _47351_ (.Y(_16395_),
    .A(_16391_),
    .B(_16394_));
 sg13g2_xor2_1 _47352_ (.B(_16395_),
    .A(_15689_),
    .X(_16396_));
 sg13g2_a21oi_1 _47353_ (.A1(net6734),
    .A2(_16396_),
    .Y(_01105_),
    .B1(_16393_));
 sg13g2_nor2_1 _47354_ (.A(net2183),
    .B(net6734),
    .Y(_16397_));
 sg13g2_or3_1 _47355_ (.A(_15689_),
    .B(_15691_),
    .C(_16387_),
    .X(_16398_));
 sg13g2_a21oi_1 _47356_ (.A1(net5363),
    .A2(_16398_),
    .Y(_16399_),
    .B1(net5185));
 sg13g2_xnor2_1 _47357_ (.Y(_16400_),
    .A(_15698_),
    .B(_16399_));
 sg13g2_a21oi_1 _47358_ (.A1(net6734),
    .A2(_16400_),
    .Y(_01106_),
    .B1(_16397_));
 sg13g2_nor2_1 _47359_ (.A(net2281),
    .B(net6734),
    .Y(_16401_));
 sg13g2_nor3_2 _47360_ (.A(_15697_),
    .B(_15698_),
    .C(_16398_),
    .Y(_16402_));
 sg13g2_o21ai_1 _47361_ (.B1(_15697_),
    .Y(_16403_),
    .A1(_15698_),
    .A2(_16398_));
 sg13g2_nand2b_1 _47362_ (.Y(_16404_),
    .B(_16403_),
    .A_N(_16402_));
 sg13g2_a22oi_1 _47363_ (.Y(_16405_),
    .B1(_16404_),
    .B2(net5363),
    .A2(net5185),
    .A1(_15697_));
 sg13g2_a21oi_1 _47364_ (.A1(net6735),
    .A2(_16405_),
    .Y(_01107_),
    .B1(_16401_));
 sg13g2_nor2_1 _47365_ (.A(net1862),
    .B(net6733),
    .Y(_16406_));
 sg13g2_o21ai_1 _47366_ (.B1(net5175),
    .Y(_16407_),
    .A1(net5339),
    .A2(_16402_));
 sg13g2_xor2_1 _47367_ (.B(_16407_),
    .A(_15700_),
    .X(_16408_));
 sg13g2_a21oi_1 _47368_ (.A1(net6732),
    .A2(_16408_),
    .Y(_01108_),
    .B1(_16406_));
 sg13g2_nand2_1 _47369_ (.Y(_16409_),
    .A(_15703_),
    .B(net5193));
 sg13g2_nand2b_2 _47370_ (.Y(_16410_),
    .B(_16402_),
    .A_N(_15700_));
 sg13g2_nand2_1 _47371_ (.Y(_16411_),
    .A(_15703_),
    .B(_16410_));
 sg13g2_nor2_1 _47372_ (.A(_15703_),
    .B(_16410_),
    .Y(_16412_));
 sg13g2_nor2_1 _47373_ (.A(net5339),
    .B(_16412_),
    .Y(_16413_));
 sg13g2_a221oi_1 _47374_ (.B2(_16413_),
    .C1(net6627),
    .B1(_16411_),
    .A1(net5338),
    .Y(_16414_),
    .A2(_16409_));
 sg13g2_a21oi_1 _47375_ (.A1(net1603),
    .A2(net6629),
    .Y(_16415_),
    .B1(_16414_));
 sg13g2_inv_1 _47376_ (.Y(_01109_),
    .A(_16415_));
 sg13g2_nor2_1 _47377_ (.A(net5186),
    .B(_16413_),
    .Y(_16416_));
 sg13g2_xor2_1 _47378_ (.B(_16416_),
    .A(_15381_),
    .X(_16417_));
 sg13g2_nand2_1 _47379_ (.Y(_16418_),
    .A(net1214),
    .B(net6627));
 sg13g2_o21ai_1 _47380_ (.B1(_16418_),
    .Y(_01110_),
    .A1(net6627),
    .A2(_16417_));
 sg13g2_nand2_1 _47381_ (.Y(_16419_),
    .A(_15380_),
    .B(_15381_));
 sg13g2_nand3_1 _47382_ (.B(_15381_),
    .C(_16412_),
    .A(_15380_),
    .Y(_16420_));
 sg13g2_o21ai_1 _47383_ (.B1(_16420_),
    .Y(_16421_),
    .A1(_15380_),
    .A2(_15381_));
 sg13g2_a21oi_1 _47384_ (.A1(net5363),
    .A2(_16421_),
    .Y(_16422_),
    .B1(net6627));
 sg13g2_o21ai_1 _47385_ (.B1(_16422_),
    .Y(_16423_),
    .A1(_15380_),
    .A2(_16416_));
 sg13g2_o21ai_1 _47386_ (.B1(_16423_),
    .Y(_16424_),
    .A1(net3454),
    .A2(net6732));
 sg13g2_inv_1 _47387_ (.Y(_01111_),
    .A(_16424_));
 sg13g2_nor2_1 _47388_ (.A(net2190),
    .B(net6733),
    .Y(_16425_));
 sg13g2_a21oi_1 _47389_ (.A1(net5363),
    .A2(_16420_),
    .Y(_16426_),
    .B1(net5186));
 sg13g2_xor2_1 _47390_ (.B(_16426_),
    .A(_15704_),
    .X(_16427_));
 sg13g2_a21oi_1 _47391_ (.A1(net6733),
    .A2(_16427_),
    .Y(_01112_),
    .B1(_16425_));
 sg13g2_nor2_1 _47392_ (.A(net2047),
    .B(net6728),
    .Y(_16428_));
 sg13g2_xnor2_1 _47393_ (.Y(_16429_),
    .A(net5365),
    .B(_15704_));
 sg13g2_nand2_1 _47394_ (.Y(_16430_),
    .A(_16426_),
    .B(_16429_));
 sg13g2_xnor2_1 _47395_ (.Y(_16431_),
    .A(_15377_),
    .B(_16430_));
 sg13g2_a21oi_1 _47396_ (.A1(net6728),
    .A2(_16431_),
    .Y(_01113_),
    .B1(_16428_));
 sg13g2_nor2_1 _47397_ (.A(net2338),
    .B(net6732),
    .Y(_16432_));
 sg13g2_nand2_1 _47398_ (.Y(_16433_),
    .A(_15377_),
    .B(_15704_));
 sg13g2_nor2_1 _47399_ (.A(_16420_),
    .B(_16433_),
    .Y(_16434_));
 sg13g2_o21ai_1 _47400_ (.B1(net5175),
    .Y(_16435_),
    .A1(net5338),
    .A2(_16434_));
 sg13g2_xnor2_1 _47401_ (.Y(_16436_),
    .A(_15710_),
    .B(_16435_));
 sg13g2_a21oi_1 _47402_ (.A1(net6732),
    .A2(_16436_),
    .Y(_01114_),
    .B1(_16432_));
 sg13g2_nand2_1 _47403_ (.Y(_16437_),
    .A(_15709_),
    .B(_15710_));
 sg13g2_nor4_1 _47404_ (.A(_15703_),
    .B(_16419_),
    .C(_16433_),
    .D(_16437_),
    .Y(_16438_));
 sg13g2_nor2b_2 _47405_ (.A(_16410_),
    .B_N(_16438_),
    .Y(_16439_));
 sg13g2_nor2_1 _47406_ (.A(_15711_),
    .B(_16439_),
    .Y(_16440_));
 sg13g2_o21ai_1 _47407_ (.B1(_16440_),
    .Y(_16441_),
    .A1(_15709_),
    .A2(_16434_));
 sg13g2_a21oi_1 _47408_ (.A1(net5365),
    .A2(_16441_),
    .Y(_16442_),
    .B1(net6627));
 sg13g2_o21ai_1 _47409_ (.B1(_16442_),
    .Y(_16443_),
    .A1(_15709_),
    .A2(net5175));
 sg13g2_o21ai_1 _47410_ (.B1(_16443_),
    .Y(_16444_),
    .A1(net3320),
    .A2(net6728));
 sg13g2_inv_1 _47411_ (.Y(_01115_),
    .A(_16444_));
 sg13g2_nor2_1 _47412_ (.A(net2057),
    .B(net6728),
    .Y(_16445_));
 sg13g2_o21ai_1 _47413_ (.B1(net5175),
    .Y(_16446_),
    .A1(net5338),
    .A2(_16439_));
 sg13g2_xnor2_1 _47414_ (.Y(_16447_),
    .A(_15330_),
    .B(_16446_));
 sg13g2_a21oi_1 _47415_ (.A1(net6728),
    .A2(_16447_),
    .Y(_01116_),
    .B1(_16445_));
 sg13g2_nor2_1 _47416_ (.A(net2145),
    .B(net6729),
    .Y(_16448_));
 sg13g2_xnor2_1 _47417_ (.Y(_16449_),
    .A(net5338),
    .B(_15330_));
 sg13g2_nor2_1 _47418_ (.A(_16446_),
    .B(_16449_),
    .Y(_16450_));
 sg13g2_xor2_1 _47419_ (.B(_16450_),
    .A(_15334_),
    .X(_16451_));
 sg13g2_a21oi_1 _47420_ (.A1(net6728),
    .A2(_16451_),
    .Y(_01117_),
    .B1(_16448_));
 sg13g2_nor2_1 _47421_ (.A(net1893),
    .B(net6728),
    .Y(_16452_));
 sg13g2_and2_1 _47422_ (.A(_15330_),
    .B(_15334_),
    .X(_16453_));
 sg13g2_nand2_1 _47423_ (.Y(_16454_),
    .A(_16439_),
    .B(_16453_));
 sg13g2_a21oi_1 _47424_ (.A1(net5365),
    .A2(_16454_),
    .Y(_16455_),
    .B1(net5189));
 sg13g2_xnor2_1 _47425_ (.Y(_16456_),
    .A(_15336_),
    .B(_16455_));
 sg13g2_a21oi_1 _47426_ (.A1(net6728),
    .A2(_16456_),
    .Y(_01118_),
    .B1(_16452_));
 sg13g2_nor2b_1 _47427_ (.A(_15336_),
    .B_N(_16453_),
    .Y(_16457_));
 sg13g2_nand3b_1 _47428_ (.B(_16439_),
    .C(_16457_),
    .Y(_16458_),
    .A_N(_15694_));
 sg13g2_o21ai_1 _47429_ (.B1(_15694_),
    .Y(_16459_),
    .A1(_15336_),
    .A2(_16454_));
 sg13g2_nand2_1 _47430_ (.Y(_16460_),
    .A(_16458_),
    .B(_16459_));
 sg13g2_a221oi_1 _47431_ (.B2(net5365),
    .C1(net6627),
    .B1(_16460_),
    .A1(_15694_),
    .Y(_16461_),
    .A2(net5186));
 sg13g2_a21oi_1 _47432_ (.A1(_18278_),
    .A2(net6627),
    .Y(_01119_),
    .B1(_16461_));
 sg13g2_nor2_1 _47433_ (.A(net1569),
    .B(net6732),
    .Y(_16462_));
 sg13g2_a21oi_2 _47434_ (.B1(net5186),
    .Y(_16463_),
    .A2(_16458_),
    .A1(net5363));
 sg13g2_xnor2_1 _47435_ (.Y(_16464_),
    .A(_15371_),
    .B(_16463_));
 sg13g2_a21oi_1 _47436_ (.A1(net6732),
    .A2(_16464_),
    .Y(_01120_),
    .B1(_16462_));
 sg13g2_nor2_1 _47437_ (.A(net1905),
    .B(net6732),
    .Y(_16465_));
 sg13g2_xnor2_1 _47438_ (.Y(_16466_),
    .A(net5339),
    .B(_15371_));
 sg13g2_nand2_1 _47439_ (.Y(_16467_),
    .A(_16463_),
    .B(_16466_));
 sg13g2_xor2_1 _47440_ (.B(_16467_),
    .A(_15373_),
    .X(_16468_));
 sg13g2_a21oi_1 _47441_ (.A1(net6732),
    .A2(_16468_),
    .Y(_01121_),
    .B1(_16465_));
 sg13g2_nor4_1 _47442_ (.A(_15371_),
    .B(_15373_),
    .C(_15694_),
    .D(_15700_),
    .Y(_16469_));
 sg13g2_nand4_1 _47443_ (.B(_16438_),
    .C(_16402_),
    .A(_16457_),
    .Y(_16470_),
    .D(_16469_));
 sg13g2_a21oi_1 _47444_ (.A1(net5365),
    .A2(net1093),
    .Y(_16471_),
    .B1(net5189));
 sg13g2_xor2_1 _47445_ (.B(_16471_),
    .A(_15332_),
    .X(_16472_));
 sg13g2_nand2_1 _47446_ (.Y(_16473_),
    .A(net1339),
    .B(net6629));
 sg13g2_o21ai_1 _47447_ (.B1(_16473_),
    .Y(_01122_),
    .A1(net6629),
    .A2(_16472_));
 sg13g2_nor2b_1 _47448_ (.A(net1093),
    .B_N(_15332_),
    .Y(_16474_));
 sg13g2_nand2_1 _47449_ (.Y(_16475_),
    .A(_15332_),
    .B(_15368_));
 sg13g2_nor2_1 _47450_ (.A(net1093),
    .B(_16475_),
    .Y(_16476_));
 sg13g2_xnor2_1 _47451_ (.Y(_16477_),
    .A(_15368_),
    .B(_16474_));
 sg13g2_a21oi_1 _47452_ (.A1(net5365),
    .A2(_16477_),
    .Y(_16478_),
    .B1(net6629));
 sg13g2_o21ai_1 _47453_ (.B1(_16478_),
    .Y(_16479_),
    .A1(_15368_),
    .A2(net5175));
 sg13g2_o21ai_1 _47454_ (.B1(_16479_),
    .Y(_16480_),
    .A1(net3283),
    .A2(net6729));
 sg13g2_inv_1 _47455_ (.Y(_01123_),
    .A(_16480_));
 sg13g2_nor2_1 _47456_ (.A(net1673),
    .B(net6723),
    .Y(_16481_));
 sg13g2_o21ai_1 _47457_ (.B1(net5173),
    .Y(_16482_),
    .A1(net5336),
    .A2(_16476_));
 sg13g2_xnor2_1 _47458_ (.Y(_16483_),
    .A(_15344_),
    .B(_16482_));
 sg13g2_a21oi_1 _47459_ (.A1(net6722),
    .A2(_16483_),
    .Y(_01124_),
    .B1(_16481_));
 sg13g2_nor2_1 _47460_ (.A(_15341_),
    .B(_15343_),
    .Y(_16484_));
 sg13g2_o21ai_1 _47461_ (.B1(net5336),
    .Y(_16485_),
    .A1(net5310),
    .A2(_16484_));
 sg13g2_nand2_1 _47462_ (.Y(_16486_),
    .A(_16476_),
    .B(_16484_));
 sg13g2_nand2_1 _47463_ (.Y(_16487_),
    .A(net5369),
    .B(_16486_));
 sg13g2_a21oi_1 _47464_ (.A1(_15344_),
    .A2(_16476_),
    .Y(_16488_),
    .B1(_15340_));
 sg13g2_o21ai_1 _47465_ (.B1(net6722),
    .Y(_16489_),
    .A1(_16487_),
    .A2(_16488_));
 sg13g2_a21oi_1 _47466_ (.A1(_15340_),
    .A2(net5184),
    .Y(_16490_),
    .B1(_16489_));
 sg13g2_a22oi_1 _47467_ (.Y(_16491_),
    .B1(_16485_),
    .B2(_16490_),
    .A2(net6626),
    .A1(net3067));
 sg13g2_inv_1 _47468_ (.Y(_01125_),
    .A(_16491_));
 sg13g2_nor2_1 _47469_ (.A(net1881),
    .B(net6722),
    .Y(_16492_));
 sg13g2_nand2_1 _47470_ (.Y(_16493_),
    .A(net5176),
    .B(_16487_));
 sg13g2_xnor2_1 _47471_ (.Y(_16494_),
    .A(_15326_),
    .B(_16493_));
 sg13g2_a21oi_1 _47472_ (.A1(net6722),
    .A2(_16494_),
    .Y(_01126_),
    .B1(_16492_));
 sg13g2_nor2b_1 _47473_ (.A(_16486_),
    .B_N(_15326_),
    .Y(_16495_));
 sg13g2_xnor2_1 _47474_ (.Y(_16496_),
    .A(_15355_),
    .B(_16495_));
 sg13g2_a221oi_1 _47475_ (.B2(net5362),
    .C1(net6626),
    .B1(_16496_),
    .A1(_15354_),
    .Y(_16497_),
    .A2(net5184));
 sg13g2_a21oi_1 _47476_ (.A1(_18279_),
    .A2(net6626),
    .Y(_01127_),
    .B1(_16497_));
 sg13g2_nor2_1 _47477_ (.A(net2582),
    .B(net6723),
    .Y(_16498_));
 sg13g2_a21oi_1 _47478_ (.A1(_15355_),
    .A2(_16495_),
    .Y(_16499_),
    .B1(net5336));
 sg13g2_nor2_1 _47479_ (.A(net5184),
    .B(_16499_),
    .Y(_16500_));
 sg13g2_xnor2_1 _47480_ (.Y(_16501_),
    .A(_15717_),
    .B(_16500_));
 sg13g2_a21oi_1 _47481_ (.A1(net6722),
    .A2(_16501_),
    .Y(_01128_),
    .B1(_16498_));
 sg13g2_nor2_1 _47482_ (.A(net1799),
    .B(net6723),
    .Y(_16502_));
 sg13g2_xnor2_1 _47483_ (.Y(_16503_),
    .A(net5336),
    .B(_15717_));
 sg13g2_nand2_1 _47484_ (.Y(_16504_),
    .A(_16500_),
    .B(_16503_));
 sg13g2_xor2_1 _47485_ (.B(_16504_),
    .A(_15361_),
    .X(_16505_));
 sg13g2_a21oi_1 _47486_ (.A1(net6722),
    .A2(_16505_),
    .Y(_01129_),
    .B1(_16502_));
 sg13g2_nor2_1 _47487_ (.A(net1847),
    .B(net6714),
    .Y(_16506_));
 sg13g2_nor4_1 _47488_ (.A(_15354_),
    .B(_15361_),
    .C(_15717_),
    .D(_16475_),
    .Y(_16507_));
 sg13g2_nand3_1 _47489_ (.B(_16484_),
    .C(_16507_),
    .A(_15326_),
    .Y(_16508_));
 sg13g2_nor2_1 _47490_ (.A(net1093),
    .B(_16508_),
    .Y(_16509_));
 sg13g2_o21ai_1 _47491_ (.B1(net5173),
    .Y(_16510_),
    .A1(net5333),
    .A2(_16509_));
 sg13g2_xnor2_1 _47492_ (.Y(_16511_),
    .A(_15727_),
    .B(_16510_));
 sg13g2_a21oi_1 _47493_ (.A1(net6714),
    .A2(_16511_),
    .Y(_01130_),
    .B1(_16506_));
 sg13g2_nand2_1 _47494_ (.Y(_16512_),
    .A(_15726_),
    .B(_15727_));
 sg13g2_nand3_1 _47495_ (.B(_15727_),
    .C(_16509_),
    .A(_15726_),
    .Y(_16513_));
 sg13g2_a21oi_1 _47496_ (.A1(_15727_),
    .A2(_16509_),
    .Y(_16514_),
    .B1(_15726_));
 sg13g2_nand2b_1 _47497_ (.Y(_16515_),
    .B(_16513_),
    .A_N(_16514_));
 sg13g2_a221oi_1 _47498_ (.B2(net5360),
    .C1(net6626),
    .B1(_16515_),
    .A1(_15725_),
    .Y(_16516_),
    .A2(net5183));
 sg13g2_a21oi_1 _47499_ (.A1(_18280_),
    .A2(net6636),
    .Y(_01131_),
    .B1(_16516_));
 sg13g2_nor2_1 _47500_ (.A(net1741),
    .B(net6722),
    .Y(_16517_));
 sg13g2_a21oi_1 _47501_ (.A1(net5360),
    .A2(_16513_),
    .Y(_16518_),
    .B1(net5183));
 sg13g2_xnor2_1 _47502_ (.Y(_16519_),
    .A(_15729_),
    .B(_16518_));
 sg13g2_a21oi_1 _47503_ (.A1(net6722),
    .A2(_16519_),
    .Y(_01132_),
    .B1(_16517_));
 sg13g2_or4_1 _47504_ (.A(_15729_),
    .B(_15732_),
    .C(net1093),
    .D(_16512_),
    .X(_16520_));
 sg13g2_or2_1 _47505_ (.X(_16521_),
    .B(_16520_),
    .A(_16508_));
 sg13g2_o21ai_1 _47506_ (.B1(_15732_),
    .Y(_16522_),
    .A1(_15729_),
    .A2(_16513_));
 sg13g2_nand2_1 _47507_ (.Y(_16523_),
    .A(_16521_),
    .B(_16522_));
 sg13g2_a221oi_1 _47508_ (.B2(net5360),
    .C1(net6625),
    .B1(_16523_),
    .A1(_15732_),
    .Y(_16524_),
    .A2(net5183));
 sg13g2_a21oi_1 _47509_ (.A1(_18281_),
    .A2(net6624),
    .Y(_01133_),
    .B1(_16524_));
 sg13g2_nor2_1 _47510_ (.A(net2717),
    .B(net6714),
    .Y(_16525_));
 sg13g2_a21oi_1 _47511_ (.A1(net5360),
    .A2(_16521_),
    .Y(_16526_),
    .B1(net5183));
 sg13g2_xnor2_1 _47512_ (.Y(_16527_),
    .A(_15767_),
    .B(_16526_));
 sg13g2_a21oi_1 _47513_ (.A1(net6714),
    .A2(_16527_),
    .Y(_01134_),
    .B1(_16525_));
 sg13g2_or2_1 _47514_ (.X(_16528_),
    .B(_15767_),
    .A(_15351_));
 sg13g2_nor2_1 _47515_ (.A(_16521_),
    .B(_16528_),
    .Y(_16529_));
 sg13g2_o21ai_1 _47516_ (.B1(_15351_),
    .Y(_16530_),
    .A1(_15767_),
    .A2(_16521_));
 sg13g2_nand2b_1 _47517_ (.Y(_16531_),
    .B(_16530_),
    .A_N(_16529_));
 sg13g2_a221oi_1 _47518_ (.B2(net5360),
    .C1(net6624),
    .B1(_16531_),
    .A1(_15351_),
    .Y(_16532_),
    .A2(net5182));
 sg13g2_a21oi_1 _47519_ (.A1(_18282_),
    .A2(net6624),
    .Y(_01135_),
    .B1(_16532_));
 sg13g2_nor2_1 _47520_ (.A(net1620),
    .B(net6714),
    .Y(_16533_));
 sg13g2_o21ai_1 _47521_ (.B1(net5173),
    .Y(_16534_),
    .A1(net5333),
    .A2(_16529_));
 sg13g2_xnor2_1 _47522_ (.Y(_16535_),
    .A(_15764_),
    .B(_16534_));
 sg13g2_a21oi_1 _47523_ (.A1(net6715),
    .A2(_16535_),
    .Y(_01136_),
    .B1(_16533_));
 sg13g2_nor2_1 _47524_ (.A(net1441),
    .B(net6715),
    .Y(_16536_));
 sg13g2_xnor2_1 _47525_ (.Y(_16537_),
    .A(net5333),
    .B(_15764_));
 sg13g2_nor2_1 _47526_ (.A(_16534_),
    .B(_16537_),
    .Y(_16538_));
 sg13g2_xnor2_1 _47527_ (.Y(_16539_),
    .A(_15310_),
    .B(_16538_));
 sg13g2_a21oi_1 _47528_ (.A1(net6715),
    .A2(_16539_),
    .Y(_01137_),
    .B1(_16536_));
 sg13g2_nand2_2 _47529_ (.Y(_16540_),
    .A(_15309_),
    .B(_15764_));
 sg13g2_nor3_2 _47530_ (.A(_16521_),
    .B(_16528_),
    .C(_16540_),
    .Y(_16541_));
 sg13g2_o21ai_1 _47531_ (.B1(net5173),
    .Y(_16542_),
    .A1(net5333),
    .A2(_16541_));
 sg13g2_xnor2_1 _47532_ (.Y(_16543_),
    .A(_15712_),
    .B(_16542_));
 sg13g2_nand2_1 _47533_ (.Y(_16544_),
    .A(net1178),
    .B(net6624));
 sg13g2_o21ai_1 _47534_ (.B1(_16544_),
    .Y(_01138_),
    .A1(net6624),
    .A2(_16543_));
 sg13g2_nand2_1 _47535_ (.Y(_16545_),
    .A(_15712_),
    .B(_16541_));
 sg13g2_nand3_1 _47536_ (.B(_15712_),
    .C(_16541_),
    .A(_15319_),
    .Y(_16546_));
 sg13g2_xnor2_1 _47537_ (.Y(_16547_),
    .A(_15320_),
    .B(_16545_));
 sg13g2_a21oi_1 _47538_ (.A1(net5358),
    .A2(_16547_),
    .Y(_16548_),
    .B1(net6624));
 sg13g2_o21ai_1 _47539_ (.B1(_16548_),
    .Y(_16549_),
    .A1(_15319_),
    .A2(net5173));
 sg13g2_o21ai_1 _47540_ (.B1(_16549_),
    .Y(_16550_),
    .A1(net3212),
    .A2(net6713));
 sg13g2_inv_1 _47541_ (.Y(_01139_),
    .A(_16550_));
 sg13g2_nor2_1 _47542_ (.A(net1703),
    .B(net6713),
    .Y(_16551_));
 sg13g2_a21oi_1 _47543_ (.A1(net5358),
    .A2(_16546_),
    .Y(_16552_),
    .B1(net5182));
 sg13g2_xnor2_1 _47544_ (.Y(_16553_),
    .A(_15346_),
    .B(_16552_));
 sg13g2_a21oi_1 _47545_ (.A1(net6713),
    .A2(_16553_),
    .Y(_01140_),
    .B1(_16551_));
 sg13g2_or3_1 _47546_ (.A(_15320_),
    .B(_15323_),
    .C(_15346_),
    .X(_16554_));
 sg13g2_nor2_1 _47547_ (.A(_16545_),
    .B(_16554_),
    .Y(_16555_));
 sg13g2_o21ai_1 _47548_ (.B1(_15323_),
    .Y(_16556_),
    .A1(_15346_),
    .A2(_16546_));
 sg13g2_nand2b_1 _47549_ (.Y(_16557_),
    .B(_16556_),
    .A_N(_16555_));
 sg13g2_a221oi_1 _47550_ (.B2(net5359),
    .C1(net6624),
    .B1(_16557_),
    .A1(_15323_),
    .Y(_16558_),
    .A2(net5183));
 sg13g2_a21oi_1 _47551_ (.A1(_18283_),
    .A2(net6624),
    .Y(_01141_),
    .B1(_16558_));
 sg13g2_nor2_1 _47552_ (.A(net1437),
    .B(net6714),
    .Y(_16559_));
 sg13g2_o21ai_1 _47553_ (.B1(net5173),
    .Y(_16560_),
    .A1(net5344),
    .A2(_16555_));
 sg13g2_xnor2_1 _47554_ (.Y(_16561_),
    .A(_15321_),
    .B(_16560_));
 sg13g2_a21oi_1 _47555_ (.A1(net6713),
    .A2(_16561_),
    .Y(_01142_),
    .B1(_16559_));
 sg13g2_nand2_1 _47556_ (.Y(_16562_),
    .A(_15321_),
    .B(_16555_));
 sg13g2_xnor2_1 _47557_ (.Y(_16563_),
    .A(_15364_),
    .B(_16562_));
 sg13g2_a221oi_1 _47558_ (.B2(net5359),
    .C1(net6625),
    .B1(_16563_),
    .A1(_15364_),
    .Y(_16564_),
    .A2(net5182));
 sg13g2_a21oi_1 _47559_ (.A1(_18284_),
    .A2(net6623),
    .Y(_01143_),
    .B1(_16564_));
 sg13g2_o21ai_1 _47560_ (.B1(net5359),
    .Y(_16565_),
    .A1(_15364_),
    .A2(_16562_));
 sg13g2_and2_1 _47561_ (.A(net5173),
    .B(_16565_),
    .X(_16566_));
 sg13g2_xnor2_1 _47562_ (.Y(_16567_),
    .A(_15755_),
    .B(_16566_));
 sg13g2_nor2_1 _47563_ (.A(net1583),
    .B(net6713),
    .Y(_16568_));
 sg13g2_a21oi_1 _47564_ (.A1(net6712),
    .A2(_16567_),
    .Y(_01144_),
    .B1(_16568_));
 sg13g2_nor2_1 _47565_ (.A(net2067),
    .B(net6713),
    .Y(_16569_));
 sg13g2_xnor2_1 _47566_ (.Y(_16570_),
    .A(net5333),
    .B(_15755_));
 sg13g2_nand2_1 _47567_ (.Y(_16571_),
    .A(_16566_),
    .B(_16570_));
 sg13g2_xnor2_1 _47568_ (.Y(_16572_),
    .A(_15356_),
    .B(_16571_));
 sg13g2_a21oi_1 _47569_ (.A1(net6712),
    .A2(_16572_),
    .Y(_01145_),
    .B1(_16569_));
 sg13g2_nor2_1 _47570_ (.A(net2184),
    .B(net6713),
    .Y(_16573_));
 sg13g2_nand3_1 _47571_ (.B(_15356_),
    .C(_15712_),
    .A(_15321_),
    .Y(_16574_));
 sg13g2_nor4_1 _47572_ (.A(_15364_),
    .B(_15755_),
    .C(_16554_),
    .D(_16574_),
    .Y(_16575_));
 sg13g2_nand2_1 _47573_ (.Y(_16576_),
    .A(_16541_),
    .B(_16575_));
 sg13g2_a21oi_1 _47574_ (.A1(net5359),
    .A2(_16576_),
    .Y(_16577_),
    .B1(net5182));
 sg13g2_xor2_1 _47575_ (.B(_16577_),
    .A(_15774_),
    .X(_16578_));
 sg13g2_a21oi_1 _47576_ (.A1(net6714),
    .A2(_16578_),
    .Y(_01146_),
    .B1(_16573_));
 sg13g2_nand2b_1 _47577_ (.Y(_16579_),
    .B(_16576_),
    .A_N(_15773_));
 sg13g2_nand4_1 _47578_ (.B(_15774_),
    .C(_16541_),
    .A(_15773_),
    .Y(_16580_),
    .D(_16575_));
 sg13g2_nand3_1 _47579_ (.B(_16579_),
    .C(_16580_),
    .A(_15775_),
    .Y(_16581_));
 sg13g2_a21oi_1 _47580_ (.A1(net5358),
    .A2(_16581_),
    .Y(_16582_),
    .B1(net6623));
 sg13g2_o21ai_1 _47581_ (.B1(_16582_),
    .Y(_16583_),
    .A1(_15773_),
    .A2(net5172));
 sg13g2_o21ai_1 _47582_ (.B1(_16583_),
    .Y(_16584_),
    .A1(net3486),
    .A2(net6708));
 sg13g2_inv_1 _47583_ (.Y(_01147_),
    .A(_16584_));
 sg13g2_nor2_1 _47584_ (.A(net1759),
    .B(net6712),
    .Y(_16585_));
 sg13g2_a21oi_1 _47585_ (.A1(net5358),
    .A2(_16580_),
    .Y(_16586_),
    .B1(net5182));
 sg13g2_xnor2_1 _47586_ (.Y(_16587_),
    .A(_15737_),
    .B(_16586_));
 sg13g2_a21oi_1 _47587_ (.A1(net6712),
    .A2(_16587_),
    .Y(_01148_),
    .B1(_16585_));
 sg13g2_nor3_1 _47588_ (.A(_15737_),
    .B(_15752_),
    .C(_16580_),
    .Y(_16588_));
 sg13g2_o21ai_1 _47589_ (.B1(_15752_),
    .Y(_16589_),
    .A1(_15737_),
    .A2(_16580_));
 sg13g2_nand2b_1 _47590_ (.Y(_16590_),
    .B(_16589_),
    .A_N(_16588_));
 sg13g2_a221oi_1 _47591_ (.B2(net5358),
    .C1(net6623),
    .B1(_16590_),
    .A1(_15752_),
    .Y(_16591_),
    .A2(net5182));
 sg13g2_a21oi_1 _47592_ (.A1(_18285_),
    .A2(net6623),
    .Y(_01149_),
    .B1(_16591_));
 sg13g2_o21ai_1 _47593_ (.B1(net5173),
    .Y(_16592_),
    .A1(net5332),
    .A2(_16588_));
 sg13g2_xnor2_1 _47594_ (.Y(_16593_),
    .A(_15280_),
    .B(_16592_));
 sg13g2_nand2_1 _47595_ (.Y(_16594_),
    .A(net1210),
    .B(net6623));
 sg13g2_o21ai_1 _47596_ (.B1(_16594_),
    .Y(_01150_),
    .A1(net6623),
    .A2(_16593_));
 sg13g2_nand3_1 _47597_ (.B(_15280_),
    .C(_16588_),
    .A(_15276_),
    .Y(_16595_));
 sg13g2_a21o_1 _47598_ (.A2(_16588_),
    .A1(_15280_),
    .B1(_15276_),
    .X(_16596_));
 sg13g2_nand2_1 _47599_ (.Y(_16597_),
    .A(_16595_),
    .B(_16596_));
 sg13g2_a221oi_1 _47600_ (.B2(net5358),
    .C1(net6623),
    .B1(_16597_),
    .A1(_15275_),
    .Y(_16598_),
    .A2(net5182));
 sg13g2_a21oi_1 _47601_ (.A1(_18286_),
    .A2(net6623),
    .Y(_01151_),
    .B1(_16598_));
 sg13g2_a21oi_1 _47602_ (.A1(net5358),
    .A2(_16595_),
    .Y(_16599_),
    .B1(net5182));
 sg13g2_xor2_1 _47603_ (.B(_16599_),
    .A(_15279_),
    .X(_16600_));
 sg13g2_nor2_1 _47604_ (.A(net1846),
    .B(net6712),
    .Y(_16601_));
 sg13g2_a21oi_1 _47605_ (.A1(net6712),
    .A2(_16600_),
    .Y(_01152_),
    .B1(_16601_));
 sg13g2_nor2_1 _47606_ (.A(net1459),
    .B(net6712),
    .Y(_16602_));
 sg13g2_mux2_1 _47607_ (.A0(_15279_),
    .A1(_15281_),
    .S(net5332),
    .X(_16603_));
 sg13g2_nand2_1 _47608_ (.Y(_16604_),
    .A(_16599_),
    .B(_16603_));
 sg13g2_xor2_1 _47609_ (.B(_16604_),
    .A(_15758_),
    .X(_16605_));
 sg13g2_a21oi_1 _47610_ (.A1(net6712),
    .A2(_16605_),
    .Y(_01153_),
    .B1(_16602_));
 sg13g2_nor2_1 _47611_ (.A(net1856),
    .B(net6708),
    .Y(_16606_));
 sg13g2_nand4_1 _47612_ (.B(_15773_),
    .C(_15774_),
    .A(_15276_),
    .Y(_16607_),
    .D(_16575_));
 sg13g2_or3_1 _47613_ (.A(_16508_),
    .B(_16540_),
    .C(_16607_),
    .X(_16608_));
 sg13g2_nor2_1 _47614_ (.A(_15758_),
    .B(_16528_),
    .Y(_16609_));
 sg13g2_nand4_1 _47615_ (.B(_15280_),
    .C(_15751_),
    .A(_15279_),
    .Y(_16610_),
    .D(_16609_));
 sg13g2_nor4_2 _47616_ (.A(_15737_),
    .B(_16520_),
    .C(_16608_),
    .Y(_16611_),
    .D(_16610_));
 sg13g2_o21ai_1 _47617_ (.B1(net5171),
    .Y(_16612_),
    .A1(net5332),
    .A2(_16611_));
 sg13g2_xor2_1 _47618_ (.B(_16612_),
    .A(_15716_),
    .X(_16613_));
 sg13g2_a21oi_1 _47619_ (.A1(net6707),
    .A2(_16613_),
    .Y(_01154_),
    .B1(_16606_));
 sg13g2_nor2_1 _47620_ (.A(net1959),
    .B(net6708),
    .Y(_16614_));
 sg13g2_nand2b_1 _47621_ (.Y(_16615_),
    .B(_16611_),
    .A_N(_15716_));
 sg13g2_nor2_1 _47622_ (.A(_15763_),
    .B(_16615_),
    .Y(_16616_));
 sg13g2_xnor2_1 _47623_ (.Y(_16617_),
    .A(_15763_),
    .B(_16615_));
 sg13g2_a22oi_1 _47624_ (.Y(_16618_),
    .B1(_16617_),
    .B2(net5356),
    .A2(net5180),
    .A1(_15763_));
 sg13g2_a21oi_1 _47625_ (.A1(net6708),
    .A2(_16618_),
    .Y(_01155_),
    .B1(_16614_));
 sg13g2_nor2_1 _47626_ (.A(net2176),
    .B(net6708),
    .Y(_16619_));
 sg13g2_o21ai_1 _47627_ (.B1(net5171),
    .Y(_16620_),
    .A1(net5332),
    .A2(_16616_));
 sg13g2_xor2_1 _47628_ (.B(_16620_),
    .A(_15761_),
    .X(_16621_));
 sg13g2_a21oi_1 _47629_ (.A1(net6707),
    .A2(_16621_),
    .Y(_01156_),
    .B1(_16619_));
 sg13g2_nor3_1 _47630_ (.A(_15761_),
    .B(_15763_),
    .C(_16615_),
    .Y(_16622_));
 sg13g2_nand2b_1 _47631_ (.Y(_16623_),
    .B(_16622_),
    .A_N(_15349_));
 sg13g2_xnor2_1 _47632_ (.Y(_16624_),
    .A(_15349_),
    .B(_16622_));
 sg13g2_o21ai_1 _47633_ (.B1(net6709),
    .Y(_16625_),
    .A1(net5332),
    .A2(_16624_));
 sg13g2_a21oi_1 _47634_ (.A1(_15349_),
    .A2(net5181),
    .Y(_16626_),
    .B1(_16625_));
 sg13g2_a21oi_1 _47635_ (.A1(_18287_),
    .A2(net6621),
    .Y(_01157_),
    .B1(_16626_));
 sg13g2_nor2_1 _47636_ (.A(net1440),
    .B(net6707),
    .Y(_16627_));
 sg13g2_a21oi_1 _47637_ (.A1(net5356),
    .A2(_16623_),
    .Y(_16628_),
    .B1(net5181));
 sg13g2_xnor2_1 _47638_ (.Y(_16629_),
    .A(_15292_),
    .B(_16628_));
 sg13g2_a21oi_1 _47639_ (.A1(net6707),
    .A2(_16629_),
    .Y(_01158_),
    .B1(_16627_));
 sg13g2_nor2_1 _47640_ (.A(_15292_),
    .B(_15294_),
    .Y(_16630_));
 sg13g2_nand2b_1 _47641_ (.Y(_16631_),
    .B(_16630_),
    .A_N(_16623_));
 sg13g2_o21ai_1 _47642_ (.B1(_15294_),
    .Y(_16632_),
    .A1(_15292_),
    .A2(_16623_));
 sg13g2_nand2_1 _47643_ (.Y(_16633_),
    .A(_16631_),
    .B(_16632_));
 sg13g2_a221oi_1 _47644_ (.B2(net5356),
    .C1(net6621),
    .B1(_16633_),
    .A1(_15294_),
    .Y(_16634_),
    .A2(net5180));
 sg13g2_a21oi_1 _47645_ (.A1(_18288_),
    .A2(net6621),
    .Y(_01159_),
    .B1(_16634_));
 sg13g2_nor2_1 _47646_ (.A(net1819),
    .B(net6707),
    .Y(_16635_));
 sg13g2_a21oi_1 _47647_ (.A1(net1134),
    .A2(_16631_),
    .Y(_16636_),
    .B1(net5181));
 sg13g2_xnor2_1 _47648_ (.Y(_16637_),
    .A(_15742_),
    .B(_16636_));
 sg13g2_a21oi_1 _47649_ (.A1(net6707),
    .A2(_16637_),
    .Y(_01160_),
    .B1(_16635_));
 sg13g2_nor2_1 _47650_ (.A(net2065),
    .B(net6707),
    .Y(_16638_));
 sg13g2_xnor2_1 _47651_ (.Y(_16639_),
    .A(net5332),
    .B(_15742_));
 sg13g2_nand2_1 _47652_ (.Y(_16640_),
    .A(_16636_),
    .B(_16639_));
 sg13g2_xnor2_1 _47653_ (.Y(_16641_),
    .A(_15800_),
    .B(_16640_));
 sg13g2_a21oi_1 _47654_ (.A1(net6707),
    .A2(_16641_),
    .Y(_01161_),
    .B1(_16638_));
 sg13g2_nor2_1 _47655_ (.A(net1922),
    .B(net6709),
    .Y(_16642_));
 sg13g2_nor4_1 _47656_ (.A(_15349_),
    .B(_15716_),
    .C(_15761_),
    .D(_15763_),
    .Y(_16643_));
 sg13g2_nor2b_1 _47657_ (.A(_15742_),
    .B_N(_16643_),
    .Y(_16644_));
 sg13g2_and4_1 _47658_ (.A(_15800_),
    .B(_16611_),
    .C(_16630_),
    .D(_16644_),
    .X(_16645_));
 sg13g2_o21ai_1 _47659_ (.B1(net5172),
    .Y(_16646_),
    .A1(net5332),
    .A2(_16645_));
 sg13g2_xor2_1 _47660_ (.B(_16646_),
    .A(_15756_),
    .X(_16647_));
 sg13g2_a21oi_1 _47661_ (.A1(net6709),
    .A2(_16647_),
    .Y(_01162_),
    .B1(_16642_));
 sg13g2_nor2_1 _47662_ (.A(net1892),
    .B(net6709),
    .Y(_16648_));
 sg13g2_nand2b_1 _47663_ (.Y(_16649_),
    .B(_16645_),
    .A_N(_15756_));
 sg13g2_or2_1 _47664_ (.X(_16650_),
    .B(_16649_),
    .A(_15736_));
 sg13g2_xnor2_1 _47665_ (.Y(_16651_),
    .A(_15736_),
    .B(_16649_));
 sg13g2_a22oi_1 _47666_ (.Y(_16652_),
    .B1(_16651_),
    .B2(net5356),
    .A2(net5181),
    .A1(_15736_));
 sg13g2_a21oi_1 _47667_ (.A1(net6709),
    .A2(_16652_),
    .Y(_01163_),
    .B1(_16648_));
 sg13g2_nor2_1 _47668_ (.A(net2011),
    .B(net6709),
    .Y(_16653_));
 sg13g2_a21oi_1 _47669_ (.A1(net5356),
    .A2(_16650_),
    .Y(_16654_),
    .B1(net5181));
 sg13g2_xnor2_1 _47670_ (.Y(_16655_),
    .A(_15302_),
    .B(_16654_));
 sg13g2_a21oi_1 _47671_ (.A1(net6709),
    .A2(_16655_),
    .Y(_01164_),
    .B1(_16653_));
 sg13g2_nor2_1 _47672_ (.A(_15302_),
    .B(_16650_),
    .Y(_16656_));
 sg13g2_nand2_1 _47673_ (.Y(_16657_),
    .A(_15749_),
    .B(_16656_));
 sg13g2_xnor2_1 _47674_ (.Y(_16658_),
    .A(_15749_),
    .B(_16656_));
 sg13g2_a21oi_1 _47675_ (.A1(net5355),
    .A2(_16658_),
    .Y(_16659_),
    .B1(net6621));
 sg13g2_o21ai_1 _47676_ (.B1(_16659_),
    .Y(_16660_),
    .A1(_15749_),
    .A2(net5171));
 sg13g2_o21ai_1 _47677_ (.B1(_16660_),
    .Y(_16661_),
    .A1(net3362),
    .A2(net6709));
 sg13g2_inv_1 _47678_ (.Y(_01165_),
    .A(_16661_));
 sg13g2_a21oi_1 _47679_ (.A1(net5355),
    .A2(_16657_),
    .Y(_16662_),
    .B1(net5180));
 sg13g2_xnor2_1 _47680_ (.Y(_16663_),
    .A(_15315_),
    .B(_16662_));
 sg13g2_nand2_1 _47681_ (.Y(_16664_),
    .A(net1197),
    .B(net6619));
 sg13g2_o21ai_1 _47682_ (.B1(_16664_),
    .Y(_01166_),
    .A1(net6619),
    .A2(_16663_));
 sg13g2_o21ai_1 _47683_ (.B1(net5355),
    .Y(_16665_),
    .A1(_15315_),
    .A2(_16657_));
 sg13g2_nand2_1 _47684_ (.Y(_16666_),
    .A(net5171),
    .B(_16665_));
 sg13g2_nor3_1 _47685_ (.A(_15315_),
    .B(_15770_),
    .C(_16657_),
    .Y(_16667_));
 sg13g2_inv_1 _47686_ (.Y(_16668_),
    .A(_16667_));
 sg13g2_a221oi_1 _47687_ (.B2(net5355),
    .C1(net6620),
    .B1(_16667_),
    .A1(_15770_),
    .Y(_16669_),
    .A2(_16666_));
 sg13g2_a21oi_1 _47688_ (.A1(_18289_),
    .A2(net6619),
    .Y(_01167_),
    .B1(_16669_));
 sg13g2_nor2_1 _47689_ (.A(net2255),
    .B(net6702),
    .Y(_16670_));
 sg13g2_o21ai_1 _47690_ (.B1(net5171),
    .Y(_16671_),
    .A1(net5329),
    .A2(_16667_));
 sg13g2_xor2_1 _47691_ (.B(_16671_),
    .A(_15745_),
    .X(_16672_));
 sg13g2_a21oi_1 _47692_ (.A1(net6702),
    .A2(_16672_),
    .Y(_01168_),
    .B1(_16670_));
 sg13g2_nor2_1 _47693_ (.A(net1887),
    .B(net6702),
    .Y(_16673_));
 sg13g2_xnor2_1 _47694_ (.Y(_16674_),
    .A(net5355),
    .B(_15745_));
 sg13g2_nor2_1 _47695_ (.A(_16671_),
    .B(_16674_),
    .Y(_16675_));
 sg13g2_xnor2_1 _47696_ (.Y(_16676_),
    .A(_15313_),
    .B(_16675_));
 sg13g2_a21oi_1 _47697_ (.A1(net6702),
    .A2(_16676_),
    .Y(_01169_),
    .B1(_16673_));
 sg13g2_nor3_2 _47698_ (.A(_15313_),
    .B(_15745_),
    .C(_16668_),
    .Y(_16677_));
 sg13g2_o21ai_1 _47699_ (.B1(net5171),
    .Y(_16678_),
    .A1(net5329),
    .A2(_16677_));
 sg13g2_xnor2_1 _47700_ (.Y(_16679_),
    .A(_15251_),
    .B(_16678_));
 sg13g2_nor2_1 _47701_ (.A(net1530),
    .B(net6697),
    .Y(_16680_));
 sg13g2_a21oi_1 _47702_ (.A1(net6702),
    .A2(_16679_),
    .Y(_01170_),
    .B1(_16680_));
 sg13g2_nand2b_1 _47703_ (.Y(_16681_),
    .B(_16678_),
    .A_N(_15249_));
 sg13g2_nand3_1 _47704_ (.B(_15251_),
    .C(_16677_),
    .A(_15249_),
    .Y(_16682_));
 sg13g2_a21oi_1 _47705_ (.A1(_15252_),
    .A2(_16682_),
    .Y(_16683_),
    .B1(net5329));
 sg13g2_nor2_1 _47706_ (.A(net6618),
    .B(_16683_),
    .Y(_16684_));
 sg13g2_a22oi_1 _47707_ (.Y(_01171_),
    .B1(_16681_),
    .B2(_16684_),
    .A2(net6618),
    .A1(_18290_));
 sg13g2_nor2_1 _47708_ (.A(net1662),
    .B(net6694),
    .Y(_16685_));
 sg13g2_a21oi_1 _47709_ (.A1(net5353),
    .A2(_16682_),
    .Y(_16686_),
    .B1(net5180));
 sg13g2_xor2_1 _47710_ (.B(_16686_),
    .A(_15261_),
    .X(_16687_));
 sg13g2_a21oi_1 _47711_ (.A1(net6694),
    .A2(_16687_),
    .Y(_01172_),
    .B1(_16685_));
 sg13g2_nor2b_1 _47712_ (.A(_16682_),
    .B_N(_15261_),
    .Y(_16688_));
 sg13g2_a21oi_1 _47713_ (.A1(net5355),
    .A2(_16688_),
    .Y(_16689_),
    .B1(_15824_));
 sg13g2_nand2_1 _47714_ (.Y(_16690_),
    .A(net5191),
    .B(_16689_));
 sg13g2_nand2_1 _47715_ (.Y(_16691_),
    .A(_15261_),
    .B(_15824_));
 sg13g2_nor2_1 _47716_ (.A(_16682_),
    .B(_16691_),
    .Y(_16692_));
 sg13g2_nand2_1 _47717_ (.Y(_16693_),
    .A(net5354),
    .B(_16692_));
 sg13g2_nand3_1 _47718_ (.B(_16690_),
    .C(_16693_),
    .A(net6702),
    .Y(_16694_));
 sg13g2_o21ai_1 _47719_ (.B1(_16694_),
    .Y(_16695_),
    .A1(net3421),
    .A2(net6701));
 sg13g2_inv_1 _47720_ (.Y(_01173_),
    .A(_16695_));
 sg13g2_a21oi_1 _47721_ (.A1(net5354),
    .A2(_16692_),
    .Y(_16696_),
    .B1(net5307));
 sg13g2_xor2_1 _47722_ (.B(_16696_),
    .A(_15807_),
    .X(_16697_));
 sg13g2_nor2_1 _47723_ (.A(net1882),
    .B(net6701),
    .Y(_16698_));
 sg13g2_a21oi_1 _47724_ (.A1(net6701),
    .A2(_16697_),
    .Y(_01174_),
    .B1(_16698_));
 sg13g2_nand2b_1 _47725_ (.Y(_16699_),
    .B(_16692_),
    .A_N(_15807_));
 sg13g2_o21ai_1 _47726_ (.B1(_15805_),
    .Y(_16700_),
    .A1(net5327),
    .A2(_16699_));
 sg13g2_nand2b_1 _47727_ (.Y(_16701_),
    .B(net5191),
    .A_N(_16700_));
 sg13g2_nor3_1 _47728_ (.A(net5328),
    .B(_15805_),
    .C(_16699_),
    .Y(_16702_));
 sg13g2_nor2_1 _47729_ (.A(net6619),
    .B(_16702_),
    .Y(_16703_));
 sg13g2_a22oi_1 _47730_ (.Y(_01175_),
    .B1(_16701_),
    .B2(_16703_),
    .A2(net6619),
    .A1(_18291_));
 sg13g2_nor2_1 _47731_ (.A(net5307),
    .B(_16702_),
    .Y(_16704_));
 sg13g2_xor2_1 _47732_ (.B(_16704_),
    .A(_15806_),
    .X(_16705_));
 sg13g2_nand2_1 _47733_ (.Y(_16706_),
    .A(net1247),
    .B(net6620));
 sg13g2_o21ai_1 _47734_ (.B1(_16706_),
    .Y(_01176_),
    .A1(net6620),
    .A2(_16705_));
 sg13g2_nor2_1 _47735_ (.A(net1677),
    .B(net6701),
    .Y(_16707_));
 sg13g2_or3_1 _47736_ (.A(_15805_),
    .B(_15806_),
    .C(_15807_),
    .X(_16708_));
 sg13g2_a22oi_1 _47737_ (.Y(_16709_),
    .B1(_16708_),
    .B2(net5356),
    .A2(_16693_),
    .A1(net5191));
 sg13g2_xnor2_1 _47738_ (.Y(_16710_),
    .A(_15722_),
    .B(_16709_));
 sg13g2_a21oi_1 _47739_ (.A1(net6703),
    .A2(_16710_),
    .Y(_01177_),
    .B1(_16707_));
 sg13g2_nor3_1 _47740_ (.A(_15722_),
    .B(_16691_),
    .C(_16708_),
    .Y(_16711_));
 sg13g2_nor2b_1 _47741_ (.A(_16682_),
    .B_N(_16711_),
    .Y(_16712_));
 sg13g2_o21ai_1 _47742_ (.B1(net5171),
    .Y(_16713_),
    .A1(net5329),
    .A2(_16712_));
 sg13g2_xnor2_1 _47743_ (.Y(_16714_),
    .A(_15820_),
    .B(_16713_));
 sg13g2_nor2_1 _47744_ (.A(net1938),
    .B(net6698),
    .Y(_16715_));
 sg13g2_a21oi_1 _47745_ (.A1(net6698),
    .A2(_16714_),
    .Y(_01178_),
    .B1(_16715_));
 sg13g2_nor2_1 _47746_ (.A(_15819_),
    .B(_15821_),
    .Y(_16716_));
 sg13g2_nand2_2 _47747_ (.Y(_16717_),
    .A(_16712_),
    .B(_16716_));
 sg13g2_nand2_1 _47748_ (.Y(_16718_),
    .A(_15822_),
    .B(_16717_));
 sg13g2_a221oi_1 _47749_ (.B2(net5353),
    .C1(net6619),
    .B1(_16718_),
    .A1(_15819_),
    .Y(_16719_),
    .A2(_16713_));
 sg13g2_a21oi_1 _47750_ (.A1(_18292_),
    .A2(net6618),
    .Y(_01179_),
    .B1(_16719_));
 sg13g2_a21oi_1 _47751_ (.A1(net5353),
    .A2(_16717_),
    .Y(_16720_),
    .B1(net5180));
 sg13g2_xnor2_1 _47752_ (.Y(_16721_),
    .A(_15812_),
    .B(_16720_));
 sg13g2_nor2_1 _47753_ (.A(net1853),
    .B(net6698),
    .Y(_16722_));
 sg13g2_a21oi_1 _47754_ (.A1(net6702),
    .A2(_16721_),
    .Y(_01180_),
    .B1(_16722_));
 sg13g2_or2_1 _47755_ (.X(_16723_),
    .B(_15812_),
    .A(_15810_));
 sg13g2_o21ai_1 _47756_ (.B1(_15813_),
    .Y(_16724_),
    .A1(_16717_),
    .A2(_16723_));
 sg13g2_a21oi_1 _47757_ (.A1(_15810_),
    .A2(_16717_),
    .Y(_16725_),
    .B1(_16724_));
 sg13g2_o21ai_1 _47758_ (.B1(net6702),
    .Y(_16726_),
    .A1(net5327),
    .A2(_16725_));
 sg13g2_a21oi_1 _47759_ (.A1(_15810_),
    .A2(net5180),
    .Y(_16727_),
    .B1(_16726_));
 sg13g2_a21oi_1 _47760_ (.A1(_18293_),
    .A2(net6616),
    .Y(_01181_),
    .B1(_16727_));
 sg13g2_o21ai_1 _47761_ (.B1(net5354),
    .Y(_16728_),
    .A1(_16717_),
    .A2(_16723_));
 sg13g2_nand2_1 _47762_ (.Y(_16729_),
    .A(net5171),
    .B(_16728_));
 sg13g2_xnor2_1 _47763_ (.Y(_16730_),
    .A(_15286_),
    .B(_16729_));
 sg13g2_nand2_1 _47764_ (.Y(_16731_),
    .A(net1205),
    .B(net6618));
 sg13g2_o21ai_1 _47765_ (.B1(_16731_),
    .Y(_01182_),
    .A1(net6618),
    .A2(_16730_));
 sg13g2_nand2b_1 _47766_ (.Y(_16732_),
    .B(_15286_),
    .A_N(_15285_));
 sg13g2_or3_1 _47767_ (.A(_16717_),
    .B(_16723_),
    .C(_16732_),
    .X(_16733_));
 sg13g2_nand2_1 _47768_ (.Y(_16734_),
    .A(_15287_),
    .B(_16733_));
 sg13g2_a221oi_1 _47769_ (.B2(net5354),
    .C1(net6618),
    .B1(_16734_),
    .A1(_15285_),
    .Y(_16735_),
    .A2(_16729_));
 sg13g2_a21oi_1 _47770_ (.A1(_18294_),
    .A2(net6616),
    .Y(_01183_),
    .B1(_16735_));
 sg13g2_a21oi_1 _47771_ (.A1(net5353),
    .A2(_16733_),
    .Y(_16736_),
    .B1(net5180));
 sg13g2_xor2_1 _47772_ (.B(_16736_),
    .A(_15255_),
    .X(_16737_));
 sg13g2_nor2_1 _47773_ (.A(net2125),
    .B(net6693),
    .Y(_16738_));
 sg13g2_a21oi_1 _47774_ (.A1(net6693),
    .A2(_16737_),
    .Y(_01184_),
    .B1(_16738_));
 sg13g2_nor2_1 _47775_ (.A(net1985),
    .B(net6698),
    .Y(_16739_));
 sg13g2_nand2b_1 _47776_ (.Y(_16740_),
    .B(_15255_),
    .A_N(_16733_));
 sg13g2_a22oi_1 _47777_ (.Y(_16741_),
    .B1(net5192),
    .B2(_16740_),
    .A2(_15255_),
    .A1(net5329));
 sg13g2_xor2_1 _47778_ (.B(_16741_),
    .A(_15299_),
    .X(_16742_));
 sg13g2_a21oi_1 _47779_ (.A1(net6697),
    .A2(_16742_),
    .Y(_01185_),
    .B1(_16739_));
 sg13g2_nor4_2 _47780_ (.A(_15313_),
    .B(_15315_),
    .C(_15745_),
    .Y(_16743_),
    .D(_15770_));
 sg13g2_and4_1 _47781_ (.A(_15249_),
    .B(_15251_),
    .C(_15299_),
    .D(_16743_),
    .X(_16744_));
 sg13g2_nor3_2 _47782_ (.A(_15302_),
    .B(_15736_),
    .C(_15756_),
    .Y(_16745_));
 sg13g2_nand4_1 _47783_ (.B(_16711_),
    .C(_16716_),
    .A(_15749_),
    .Y(_16746_),
    .D(_16745_));
 sg13g2_nor3_1 _47784_ (.A(_16723_),
    .B(_16732_),
    .C(_16746_),
    .Y(_16747_));
 sg13g2_nand4_1 _47785_ (.B(_16744_),
    .C(_16645_),
    .A(_15255_),
    .Y(_16748_),
    .D(_16747_));
 sg13g2_nand2b_1 _47786_ (.Y(_16749_),
    .B(_15258_),
    .A_N(net1111));
 sg13g2_nand2_1 _47787_ (.Y(_16750_),
    .A(net5351),
    .B(_16749_));
 sg13g2_a21oi_1 _47788_ (.A1(_15257_),
    .A2(net1111),
    .Y(_16751_),
    .B1(_16750_));
 sg13g2_o21ai_1 _47789_ (.B1(net6695),
    .Y(_16752_),
    .A1(net5352),
    .A2(_15257_));
 sg13g2_nor3_1 _47790_ (.A(net5306),
    .B(_16751_),
    .C(_16752_),
    .Y(_16753_));
 sg13g2_a21o_1 _47791_ (.A2(net6615),
    .A1(net2285),
    .B1(_16753_),
    .X(_01186_));
 sg13g2_nand2_1 _47792_ (.Y(_16754_),
    .A(net5170),
    .B(_16750_));
 sg13g2_xnor2_1 _47793_ (.Y(_16755_),
    .A(_15817_),
    .B(_16754_));
 sg13g2_nor2_1 _47794_ (.A(net2213),
    .B(net6693),
    .Y(_16756_));
 sg13g2_a21oi_1 _47795_ (.A1(net6693),
    .A2(_16755_),
    .Y(_01187_),
    .B1(_16756_));
 sg13g2_nor2_1 _47796_ (.A(net2051),
    .B(net6693),
    .Y(_16757_));
 sg13g2_xnor2_1 _47797_ (.Y(_16758_),
    .A(net5351),
    .B(_15816_));
 sg13g2_nor2_1 _47798_ (.A(_16754_),
    .B(_16758_),
    .Y(_16759_));
 sg13g2_xnor2_1 _47799_ (.Y(_16760_),
    .A(_15793_),
    .B(_16759_));
 sg13g2_a21oi_1 _47800_ (.A1(net6693),
    .A2(_16760_),
    .Y(_01188_),
    .B1(_16757_));
 sg13g2_nor2_1 _47801_ (.A(net1674),
    .B(net6693),
    .Y(_16761_));
 sg13g2_a21oi_1 _47802_ (.A1(_15794_),
    .A2(_16759_),
    .Y(_16762_),
    .B1(net5306));
 sg13g2_xnor2_1 _47803_ (.Y(_16763_),
    .A(_15297_),
    .B(_16762_));
 sg13g2_a21oi_1 _47804_ (.A1(net6693),
    .A2(_16763_),
    .Y(_01189_),
    .B1(_16761_));
 sg13g2_nor2_1 _47805_ (.A(net1859),
    .B(net6692),
    .Y(_16764_));
 sg13g2_nand3_1 _47806_ (.B(_15794_),
    .C(_15817_),
    .A(_15297_),
    .Y(_16765_));
 sg13g2_nor2_1 _47807_ (.A(_16749_),
    .B(_16765_),
    .Y(_16766_));
 sg13g2_a21oi_1 _47808_ (.A1(net5351),
    .A2(_16766_),
    .Y(_16767_),
    .B1(net5306));
 sg13g2_xnor2_1 _47809_ (.Y(_16768_),
    .A(_15790_),
    .B(_16767_));
 sg13g2_a21oi_1 _47810_ (.A1(net6692),
    .A2(_16768_),
    .Y(_01190_),
    .B1(_16764_));
 sg13g2_nor2_1 _47811_ (.A(net2001),
    .B(net6691),
    .Y(_16769_));
 sg13g2_nand2_1 _47812_ (.Y(_16770_),
    .A(_15790_),
    .B(_16766_));
 sg13g2_nor2_1 _47813_ (.A(_15266_),
    .B(_16770_),
    .Y(_16771_));
 sg13g2_xnor2_1 _47814_ (.Y(_16772_),
    .A(_15266_),
    .B(_16770_));
 sg13g2_a22oi_1 _47815_ (.Y(_16773_),
    .B1(_16772_),
    .B2(net5351),
    .A2(net5179),
    .A1(_15266_));
 sg13g2_a21oi_1 _47816_ (.A1(net6691),
    .A2(_16773_),
    .Y(_01191_),
    .B1(_16769_));
 sg13g2_o21ai_1 _47817_ (.B1(net5170),
    .Y(_16774_),
    .A1(net5326),
    .A2(_16771_));
 sg13g2_inv_1 _47818_ (.Y(_16775_),
    .A(_16774_));
 sg13g2_xnor2_1 _47819_ (.Y(_16776_),
    .A(_15815_),
    .B(_16774_));
 sg13g2_nand2_1 _47820_ (.Y(_16777_),
    .A(net1198),
    .B(net6614));
 sg13g2_o21ai_1 _47821_ (.B1(_16777_),
    .Y(_01192_),
    .A1(net6614),
    .A2(_16776_));
 sg13g2_nor2_1 _47822_ (.A(net2013),
    .B(net6694),
    .Y(_16778_));
 sg13g2_nand2_1 _47823_ (.Y(_16779_),
    .A(_15815_),
    .B(_16771_));
 sg13g2_a22oi_1 _47824_ (.Y(_16780_),
    .B1(net5191),
    .B2(_16779_),
    .A2(_15815_),
    .A1(net5326));
 sg13g2_xnor2_1 _47825_ (.Y(_16781_),
    .A(_15247_),
    .B(_16780_));
 sg13g2_a21oi_1 _47826_ (.A1(net6694),
    .A2(_16781_),
    .Y(_01193_),
    .B1(_16778_));
 sg13g2_nor2_1 _47827_ (.A(net2187),
    .B(net6694),
    .Y(_16782_));
 sg13g2_nor2b_1 _47828_ (.A(_15247_),
    .B_N(_15815_),
    .Y(_16783_));
 sg13g2_o21ai_1 _47829_ (.B1(_16775_),
    .Y(_16784_),
    .A1(net5326),
    .A2(_16783_));
 sg13g2_xor2_1 _47830_ (.B(_16784_),
    .A(_15781_),
    .X(_16785_));
 sg13g2_a21oi_1 _47831_ (.A1(net6694),
    .A2(_16785_),
    .Y(_01194_),
    .B1(_16782_));
 sg13g2_nand2_1 _47832_ (.Y(_16786_),
    .A(_15790_),
    .B(_16783_));
 sg13g2_nor4_1 _47833_ (.A(_15266_),
    .B(_15780_),
    .C(_15781_),
    .D(_16786_),
    .Y(_16787_));
 sg13g2_nand2_1 _47834_ (.Y(_16788_),
    .A(_16766_),
    .B(_16787_));
 sg13g2_nand2_1 _47835_ (.Y(_16789_),
    .A(_15782_),
    .B(_16788_));
 sg13g2_a221oi_1 _47836_ (.B2(net5351),
    .C1(net6616),
    .B1(_16789_),
    .A1(_15780_),
    .Y(_16790_),
    .A2(_16784_));
 sg13g2_a21oi_1 _47837_ (.A1(_18295_),
    .A2(net6616),
    .Y(_01195_),
    .B1(_16790_));
 sg13g2_nor2_1 _47838_ (.A(net1932),
    .B(net6691),
    .Y(_16791_));
 sg13g2_a21oi_1 _47839_ (.A1(net5350),
    .A2(_16788_),
    .Y(_16792_),
    .B1(net5179));
 sg13g2_xnor2_1 _47840_ (.Y(_16793_),
    .A(_15828_),
    .B(_16792_));
 sg13g2_a21oi_1 _47841_ (.A1(net6690),
    .A2(_16793_),
    .Y(_01196_),
    .B1(_16791_));
 sg13g2_nor2_1 _47842_ (.A(_15828_),
    .B(_16788_),
    .Y(_16794_));
 sg13g2_a21o_1 _47843_ (.A2(_16794_),
    .A1(net5350),
    .B1(_15841_),
    .X(_16795_));
 sg13g2_and2_1 _47844_ (.A(_15841_),
    .B(_16794_),
    .X(_16796_));
 sg13g2_a21oi_1 _47845_ (.A1(net5350),
    .A2(_16796_),
    .Y(_16797_),
    .B1(net6614));
 sg13g2_o21ai_1 _47846_ (.B1(_16797_),
    .Y(_16798_),
    .A1(net5306),
    .A2(_16795_));
 sg13g2_o21ai_1 _47847_ (.B1(_16798_),
    .Y(_16799_),
    .A1(net3222),
    .A2(net6681));
 sg13g2_inv_1 _47848_ (.Y(_01197_),
    .A(_16799_));
 sg13g2_nor2_1 _47849_ (.A(net2096),
    .B(net6690),
    .Y(_16800_));
 sg13g2_o21ai_1 _47850_ (.B1(net5170),
    .Y(_16801_),
    .A1(net5326),
    .A2(_16796_));
 sg13g2_xor2_1 _47851_ (.B(_16801_),
    .A(_15848_),
    .X(_16802_));
 sg13g2_a21oi_1 _47852_ (.A1(net6690),
    .A2(_16802_),
    .Y(_01198_),
    .B1(_16800_));
 sg13g2_nor2_1 _47853_ (.A(_15847_),
    .B(_15848_),
    .Y(_16803_));
 sg13g2_nand2_1 _47854_ (.Y(_16804_),
    .A(_16796_),
    .B(_16803_));
 sg13g2_nand2_1 _47855_ (.Y(_16805_),
    .A(_15849_),
    .B(_16804_));
 sg13g2_a221oi_1 _47856_ (.B2(net5350),
    .C1(net6615),
    .B1(_16805_),
    .A1(_15847_),
    .Y(_16806_),
    .A2(_16801_));
 sg13g2_a21oi_1 _47857_ (.A1(_18296_),
    .A2(net6614),
    .Y(_01199_),
    .B1(_16806_));
 sg13g2_nor2_1 _47858_ (.A(net2757),
    .B(net6690),
    .Y(_16807_));
 sg13g2_a21oi_1 _47859_ (.A1(net5350),
    .A2(_16804_),
    .Y(_16808_),
    .B1(net5179));
 sg13g2_xor2_1 _47860_ (.B(_16808_),
    .A(_15798_),
    .X(_16809_));
 sg13g2_a21oi_1 _47861_ (.A1(net6690),
    .A2(_16809_),
    .Y(_01200_),
    .B1(_16807_));
 sg13g2_nor2_1 _47862_ (.A(net2518),
    .B(net6692),
    .Y(_16810_));
 sg13g2_xnor2_1 _47863_ (.Y(_16811_),
    .A(net5350),
    .B(_15798_));
 sg13g2_nand2_1 _47864_ (.Y(_16812_),
    .A(_16808_),
    .B(_16811_));
 sg13g2_xnor2_1 _47865_ (.Y(_16813_),
    .A(_15835_),
    .B(_16812_));
 sg13g2_a21oi_1 _47866_ (.A1(net6692),
    .A2(_16813_),
    .Y(_01201_),
    .B1(_16810_));
 sg13g2_nor2_1 _47867_ (.A(_15257_),
    .B(_15828_),
    .Y(_16814_));
 sg13g2_nand3_1 _47868_ (.B(_15835_),
    .C(_16803_),
    .A(_15798_),
    .Y(_16815_));
 sg13g2_nor2_1 _47869_ (.A(_16765_),
    .B(_16815_),
    .Y(_16816_));
 sg13g2_nand4_1 _47870_ (.B(_16787_),
    .C(_16814_),
    .A(_15841_),
    .Y(_16817_),
    .D(_16816_));
 sg13g2_nor2_2 _47871_ (.A(net1111),
    .B(_16817_),
    .Y(_16818_));
 sg13g2_a21oi_1 _47872_ (.A1(net5350),
    .A2(_16818_),
    .Y(_16819_),
    .B1(net5308));
 sg13g2_xor2_1 _47873_ (.B(_16819_),
    .A(_15829_),
    .X(_16820_));
 sg13g2_nand2_1 _47874_ (.Y(_16821_),
    .A(net1291),
    .B(net6614));
 sg13g2_o21ai_1 _47875_ (.B1(_16821_),
    .Y(_01202_),
    .A1(net6614),
    .A2(_16820_));
 sg13g2_nor2_1 _47876_ (.A(net1984),
    .B(net6691),
    .Y(_16822_));
 sg13g2_nand2b_1 _47877_ (.Y(_16823_),
    .B(_16818_),
    .A_N(_15829_));
 sg13g2_nor2_1 _47878_ (.A(_15851_),
    .B(_16823_),
    .Y(_16824_));
 sg13g2_xnor2_1 _47879_ (.Y(_16825_),
    .A(_15851_),
    .B(_16823_));
 sg13g2_a22oi_1 _47880_ (.Y(_16826_),
    .B1(_16825_),
    .B2(net5351),
    .A2(net5179),
    .A1(_15851_));
 sg13g2_a21oi_1 _47881_ (.A1(net6690),
    .A2(_16826_),
    .Y(_01203_),
    .B1(_16822_));
 sg13g2_nor2_1 _47882_ (.A(net1794),
    .B(net6681),
    .Y(_16827_));
 sg13g2_a21oi_1 _47883_ (.A1(net5350),
    .A2(_16824_),
    .Y(_16828_),
    .B1(net5306));
 sg13g2_xor2_1 _47884_ (.B(_16828_),
    .A(_15833_),
    .X(_16829_));
 sg13g2_a21oi_1 _47885_ (.A1(net6681),
    .A2(_16829_),
    .Y(_01204_),
    .B1(_16827_));
 sg13g2_nand2b_1 _47886_ (.Y(_16830_),
    .B(_16824_),
    .A_N(_15833_));
 sg13g2_o21ai_1 _47887_ (.B1(_15787_),
    .Y(_16831_),
    .A1(net5326),
    .A2(_16830_));
 sg13g2_or2_1 _47888_ (.X(_16832_),
    .B(_16831_),
    .A(net5308));
 sg13g2_nor4_1 _47889_ (.A(_15787_),
    .B(_15829_),
    .C(_15833_),
    .D(_15851_),
    .Y(_16833_));
 sg13g2_nor2_1 _47890_ (.A(_15787_),
    .B(_16830_),
    .Y(_16834_));
 sg13g2_a21oi_1 _47891_ (.A1(net5352),
    .A2(_16834_),
    .Y(_16835_),
    .B1(net6622));
 sg13g2_a22oi_1 _47892_ (.Y(_01205_),
    .B1(_16832_),
    .B2(_16835_),
    .A2(net6615),
    .A1(_18297_));
 sg13g2_o21ai_1 _47893_ (.B1(net5170),
    .Y(_16836_),
    .A1(net5326),
    .A2(_16834_));
 sg13g2_xnor2_1 _47894_ (.Y(_16837_),
    .A(_15863_),
    .B(_16836_));
 sg13g2_nor2_1 _47895_ (.A(net2078),
    .B(net6691),
    .Y(_16838_));
 sg13g2_a21oi_1 _47896_ (.A1(net6691),
    .A2(_16837_),
    .Y(_01206_),
    .B1(_16838_));
 sg13g2_nand3_1 _47897_ (.B(_15866_),
    .C(_16834_),
    .A(_15863_),
    .Y(_16839_));
 sg13g2_nand2_1 _47898_ (.Y(_16840_),
    .A(_15868_),
    .B(_16839_));
 sg13g2_a221oi_1 _47899_ (.B2(net5351),
    .C1(net6614),
    .B1(_16840_),
    .A1(_15867_),
    .Y(_16841_),
    .A2(_16836_));
 sg13g2_a21oi_1 _47900_ (.A1(_18298_),
    .A2(net6614),
    .Y(_01207_),
    .B1(_16841_));
 sg13g2_nor2_1 _47901_ (.A(net3305),
    .B(net6690),
    .Y(_16842_));
 sg13g2_a21oi_1 _47902_ (.A1(net5352),
    .A2(_16839_),
    .Y(_16843_),
    .B1(net5179));
 sg13g2_xnor2_1 _47903_ (.Y(_16844_),
    .A(_15844_),
    .B(_16843_));
 sg13g2_a21oi_1 _47904_ (.A1(net6690),
    .A2(_16844_),
    .Y(_01208_),
    .B1(_16842_));
 sg13g2_nor2_1 _47905_ (.A(net3172),
    .B(net6695),
    .Y(_16845_));
 sg13g2_xnor2_1 _47906_ (.Y(_16846_),
    .A(net5352),
    .B(_15845_));
 sg13g2_nand2_1 _47907_ (.Y(_16847_),
    .A(_16843_),
    .B(_16846_));
 sg13g2_xnor2_1 _47908_ (.Y(_16848_),
    .A(_15862_),
    .B(_16847_));
 sg13g2_a21oi_1 _47909_ (.A1(net6695),
    .A2(_16848_),
    .Y(_01209_),
    .B1(_16845_));
 sg13g2_and4_1 _47910_ (.A(_15845_),
    .B(_15863_),
    .C(_15866_),
    .D(_16833_),
    .X(_16849_));
 sg13g2_nand3_1 _47911_ (.B(_16849_),
    .C(_16818_),
    .A(_15862_),
    .Y(_16850_));
 sg13g2_o21ai_1 _47912_ (.B1(net5191),
    .Y(_16851_),
    .A1(net5323),
    .A2(net1138));
 sg13g2_xnor2_1 _47913_ (.Y(_16852_),
    .A(_15838_),
    .B(_16851_));
 sg13g2_nand2_1 _47914_ (.Y(_16853_),
    .A(net1246),
    .B(net6613));
 sg13g2_o21ai_1 _47915_ (.B1(_16853_),
    .Y(_01210_),
    .A1(net6613),
    .A2(_16852_));
 sg13g2_nor2_1 _47916_ (.A(net1543),
    .B(net6680),
    .Y(_16854_));
 sg13g2_nor2_1 _47917_ (.A(_15838_),
    .B(_15859_),
    .Y(_16855_));
 sg13g2_nand2b_1 _47918_ (.Y(_16856_),
    .B(_16855_),
    .A_N(net1138));
 sg13g2_o21ai_1 _47919_ (.B1(_15859_),
    .Y(_16857_),
    .A1(_15838_),
    .A2(net1138));
 sg13g2_nand2_1 _47920_ (.Y(_16858_),
    .A(_16856_),
    .B(_16857_));
 sg13g2_a22oi_1 _47921_ (.Y(_16859_),
    .B1(_16858_),
    .B2(net5357),
    .A2(net5178),
    .A1(_15859_));
 sg13g2_a21oi_1 _47922_ (.A1(net6679),
    .A2(_16859_),
    .Y(_01211_),
    .B1(_16854_));
 sg13g2_nor2_1 _47923_ (.A(net1899),
    .B(net6680),
    .Y(_16860_));
 sg13g2_nand2_1 _47924_ (.Y(_16861_),
    .A(net5347),
    .B(_16856_));
 sg13g2_nand2_1 _47925_ (.Y(_16862_),
    .A(net5169),
    .B(_16861_));
 sg13g2_xor2_1 _47926_ (.B(_16862_),
    .A(_15879_),
    .X(_16863_));
 sg13g2_a21oi_1 _47927_ (.A1(net6679),
    .A2(_16863_),
    .Y(_01212_),
    .B1(_16860_));
 sg13g2_nand2_1 _47928_ (.Y(_16864_),
    .A(net1224),
    .B(net6613));
 sg13g2_nor2_1 _47929_ (.A(_15876_),
    .B(_15879_),
    .Y(_16865_));
 sg13g2_o21ai_1 _47930_ (.B1(_16861_),
    .Y(_16866_),
    .A1(net5323),
    .A2(_16865_));
 sg13g2_o21ai_1 _47931_ (.B1(_15876_),
    .Y(_16867_),
    .A1(_15879_),
    .A2(_16856_));
 sg13g2_o21ai_1 _47932_ (.B1(net6685),
    .Y(_16868_),
    .A1(net5347),
    .A2(_15876_));
 sg13g2_a21o_1 _47933_ (.A2(_16867_),
    .A1(_16866_),
    .B1(_16868_),
    .X(_16869_));
 sg13g2_o21ai_1 _47934_ (.B1(_16864_),
    .Y(_01213_),
    .A1(net5306),
    .A2(_16869_));
 sg13g2_nor2_1 _47935_ (.A(net2029),
    .B(net6680),
    .Y(_16870_));
 sg13g2_nor2_1 _47936_ (.A(net5178),
    .B(_16866_),
    .Y(_16871_));
 sg13g2_xnor2_1 _47937_ (.Y(_16872_),
    .A(_15889_),
    .B(_16871_));
 sg13g2_a21oi_1 _47938_ (.A1(net6679),
    .A2(_16872_),
    .Y(_01214_),
    .B1(_16870_));
 sg13g2_o21ai_1 _47939_ (.B1(_15887_),
    .Y(_16873_),
    .A1(net5178),
    .A2(_16866_));
 sg13g2_nand2_1 _47940_ (.Y(_16874_),
    .A(_16855_),
    .B(_16865_));
 sg13g2_nor4_2 _47941_ (.A(_15887_),
    .B(_15889_),
    .C(net1138),
    .Y(_16875_),
    .D(_16874_));
 sg13g2_o21ai_1 _47942_ (.B1(net5347),
    .Y(_16876_),
    .A1(_15891_),
    .A2(_16875_));
 sg13g2_nand3_1 _47943_ (.B(_16873_),
    .C(_16876_),
    .A(net6685),
    .Y(_16877_));
 sg13g2_o21ai_1 _47944_ (.B1(_16877_),
    .Y(_16878_),
    .A1(net3365),
    .A2(net6685));
 sg13g2_inv_1 _47945_ (.Y(_01215_),
    .A(_16878_));
 sg13g2_o21ai_1 _47946_ (.B1(net5169),
    .Y(_16879_),
    .A1(net5323),
    .A2(_16875_));
 sg13g2_xnor2_1 _47947_ (.Y(_16880_),
    .A(_15857_),
    .B(_16879_));
 sg13g2_nor2_1 _47948_ (.A(net1606),
    .B(net6684),
    .Y(_16881_));
 sg13g2_a21oi_1 _47949_ (.A1(net6685),
    .A2(_16880_),
    .Y(_01216_),
    .B1(_16881_));
 sg13g2_nor2_1 _47950_ (.A(net1663),
    .B(net6678),
    .Y(_16882_));
 sg13g2_xnor2_1 _47951_ (.Y(_16883_),
    .A(net5323),
    .B(_15857_));
 sg13g2_nor2_1 _47952_ (.A(_16879_),
    .B(_16883_),
    .Y(_16884_));
 sg13g2_xor2_1 _47953_ (.B(_16884_),
    .A(_15872_),
    .X(_16885_));
 sg13g2_a21oi_1 _47954_ (.A1(net6684),
    .A2(_16885_),
    .Y(_01217_),
    .B1(_16882_));
 sg13g2_nand3_1 _47955_ (.B(_15872_),
    .C(_16875_),
    .A(_15857_),
    .Y(_16886_));
 sg13g2_a21o_1 _47956_ (.A2(_16886_),
    .A1(net5346),
    .B1(net5177),
    .X(_16887_));
 sg13g2_xnor2_1 _47957_ (.Y(_16888_),
    .A(_15216_),
    .B(_16887_));
 sg13g2_nand2_1 _47958_ (.Y(_16889_),
    .A(net1231),
    .B(net6609));
 sg13g2_o21ai_1 _47959_ (.B1(_16889_),
    .Y(_01218_),
    .A1(net6609),
    .A2(_16888_));
 sg13g2_nand2b_1 _47960_ (.Y(_16890_),
    .B(_16887_),
    .A_N(_15214_));
 sg13g2_nand2_1 _47961_ (.Y(_16891_),
    .A(_15214_),
    .B(_15216_));
 sg13g2_nor2_1 _47962_ (.A(_16886_),
    .B(_16891_),
    .Y(_16892_));
 sg13g2_o21ai_1 _47963_ (.B1(net5346),
    .Y(_16893_),
    .A1(_15217_),
    .A2(_16892_));
 sg13g2_nand3_1 _47964_ (.B(_16890_),
    .C(_16893_),
    .A(net6682),
    .Y(_16894_));
 sg13g2_o21ai_1 _47965_ (.B1(_16894_),
    .Y(_16895_),
    .A1(net3497),
    .A2(net6682));
 sg13g2_inv_1 _47966_ (.Y(_01219_),
    .A(_16895_));
 sg13g2_a21oi_1 _47967_ (.A1(net5347),
    .A2(_16892_),
    .Y(_16896_),
    .B1(net5305));
 sg13g2_nand2_1 _47968_ (.Y(_16897_),
    .A(_15221_),
    .B(_16892_));
 sg13g2_xnor2_1 _47969_ (.Y(_16898_),
    .A(_15221_),
    .B(_16896_));
 sg13g2_nand2_1 _47970_ (.Y(_16899_),
    .A(net1226),
    .B(net6613));
 sg13g2_o21ai_1 _47971_ (.B1(_16899_),
    .Y(_01220_),
    .A1(net6609),
    .A2(_16898_));
 sg13g2_o21ai_1 _47972_ (.B1(_15243_),
    .Y(_16900_),
    .A1(net5323),
    .A2(_16897_));
 sg13g2_or2_1 _47973_ (.X(_16901_),
    .B(_16900_),
    .A(net5305));
 sg13g2_nor3_1 _47974_ (.A(net5323),
    .B(_15243_),
    .C(_16897_),
    .Y(_16902_));
 sg13g2_nor2_1 _47975_ (.A(net6610),
    .B(_16902_),
    .Y(_16903_));
 sg13g2_nor2_1 _47976_ (.A(_15243_),
    .B(_16897_),
    .Y(_16904_));
 sg13g2_a22oi_1 _47977_ (.Y(_01221_),
    .B1(_16901_),
    .B2(_16903_),
    .A2(net6609),
    .A1(_18309_));
 sg13g2_o21ai_1 _47978_ (.B1(net5169),
    .Y(_16905_),
    .A1(net5323),
    .A2(_16904_));
 sg13g2_xor2_1 _47979_ (.B(_16905_),
    .A(_15884_),
    .X(_16906_));
 sg13g2_nand2_1 _47980_ (.Y(_16907_),
    .A(net1182),
    .B(net6611));
 sg13g2_o21ai_1 _47981_ (.B1(_16907_),
    .Y(_01222_),
    .A1(net6609),
    .A2(_16906_));
 sg13g2_nor2_1 _47982_ (.A(net1505),
    .B(net6684),
    .Y(_16908_));
 sg13g2_nor2_1 _47983_ (.A(_15883_),
    .B(_15884_),
    .Y(_16909_));
 sg13g2_nand2_1 _47984_ (.Y(_16910_),
    .A(_16902_),
    .B(_16909_));
 sg13g2_nand3_1 _47985_ (.B(_16904_),
    .C(_16909_),
    .A(net5347),
    .Y(_16911_));
 sg13g2_inv_1 _47986_ (.Y(_16912_),
    .A(_16911_));
 sg13g2_a221oi_1 _47987_ (.B2(_15883_),
    .C1(_16912_),
    .B1(_16905_),
    .A1(net5347),
    .Y(_16913_),
    .A2(_15885_));
 sg13g2_a21oi_1 _47988_ (.A1(net6684),
    .A2(_16913_),
    .Y(_01223_),
    .B1(_16908_));
 sg13g2_and3_1 _47989_ (.X(_16914_),
    .A(_15892_),
    .B(net5191),
    .C(_16910_));
 sg13g2_nor2_1 _47990_ (.A(_15892_),
    .B(_16910_),
    .Y(_16915_));
 sg13g2_nor3_1 _47991_ (.A(net6609),
    .B(_16914_),
    .C(_16915_),
    .Y(_16916_));
 sg13g2_a21oi_1 _47992_ (.A1(_18312_),
    .A2(net6610),
    .Y(_01224_),
    .B1(_16916_));
 sg13g2_nor2_1 _47993_ (.A(net1422),
    .B(net6684),
    .Y(_16917_));
 sg13g2_nor2_1 _47994_ (.A(net5305),
    .B(_16915_),
    .Y(_16918_));
 sg13g2_xor2_1 _47995_ (.B(_16918_),
    .A(_15227_),
    .X(_16919_));
 sg13g2_a21oi_1 _47996_ (.A1(net6684),
    .A2(_16919_),
    .Y(_01225_),
    .B1(_16917_));
 sg13g2_nor3_1 _47997_ (.A(_15227_),
    .B(_15892_),
    .C(_16891_),
    .Y(_16920_));
 sg13g2_nand2_1 _47998_ (.Y(_16921_),
    .A(_16909_),
    .B(_16920_));
 sg13g2_nand2b_1 _47999_ (.Y(_16922_),
    .B(_15221_),
    .A_N(_15243_));
 sg13g2_or3_1 _48000_ (.A(_16886_),
    .B(_16921_),
    .C(_16922_),
    .X(_16923_));
 sg13g2_o21ai_1 _48001_ (.B1(net5191),
    .Y(_16924_),
    .A1(net5324),
    .A2(_16923_));
 sg13g2_nor2b_1 _48002_ (.A(_16923_),
    .B_N(_15874_),
    .Y(_16925_));
 sg13g2_xor2_1 _48003_ (.B(_16924_),
    .A(_15874_),
    .X(_16926_));
 sg13g2_nand2_1 _48004_ (.Y(_16927_),
    .A(net1301),
    .B(net6611));
 sg13g2_o21ai_1 _48005_ (.B1(_16927_),
    .Y(_01226_),
    .A1(net6611),
    .A2(_16926_));
 sg13g2_and2_1 _48006_ (.A(_15223_),
    .B(_16925_),
    .X(_16928_));
 sg13g2_a21oi_1 _48007_ (.A1(net5346),
    .A2(_16925_),
    .Y(_16929_),
    .B1(_15223_));
 sg13g2_a21oi_1 _48008_ (.A1(net5346),
    .A2(_16928_),
    .Y(_16930_),
    .B1(_16929_));
 sg13g2_nor3_1 _48009_ (.A(net6609),
    .B(net5305),
    .C(_16930_),
    .Y(_16931_));
 sg13g2_a21o_1 _48010_ (.A2(net6609),
    .A1(net2112),
    .B1(_16931_),
    .X(_01227_));
 sg13g2_nor2_1 _48011_ (.A(net1384),
    .B(net6682),
    .Y(_16932_));
 sg13g2_a21oi_1 _48012_ (.A1(net5346),
    .A2(_16928_),
    .Y(_16933_),
    .B1(net5305));
 sg13g2_xnor2_1 _48013_ (.Y(_16934_),
    .A(_15237_),
    .B(_16933_));
 sg13g2_a21oi_1 _48014_ (.A1(net6682),
    .A2(_16934_),
    .Y(_01228_),
    .B1(_16932_));
 sg13g2_nand4_1 _48015_ (.B(_15223_),
    .C(_15237_),
    .A(_15212_),
    .Y(_16935_),
    .D(_15874_));
 sg13g2_nor2_2 _48016_ (.A(_16923_),
    .B(_16935_),
    .Y(_16936_));
 sg13g2_a21oi_1 _48017_ (.A1(_15237_),
    .A2(_16928_),
    .Y(_16937_),
    .B1(_15212_));
 sg13g2_o21ai_1 _48018_ (.B1(net5346),
    .Y(_16938_),
    .A1(_16936_),
    .A2(_16937_));
 sg13g2_and2_1 _48019_ (.A(net6682),
    .B(_16938_),
    .X(_16939_));
 sg13g2_o21ai_1 _48020_ (.B1(_16939_),
    .Y(_16940_),
    .A1(_15212_),
    .A2(net5169));
 sg13g2_o21ai_1 _48021_ (.B1(_16940_),
    .Y(_16941_),
    .A1(net3635),
    .A2(net6682));
 sg13g2_inv_1 _48022_ (.Y(_01229_),
    .A(_16941_));
 sg13g2_nor2_1 _48023_ (.A(net2148),
    .B(net6685),
    .Y(_16942_));
 sg13g2_o21ai_1 _48024_ (.B1(net5169),
    .Y(_16943_),
    .A1(net5324),
    .A2(_16936_));
 sg13g2_xnor2_1 _48025_ (.Y(_16944_),
    .A(net1123),
    .B(_16943_));
 sg13g2_a21oi_1 _48026_ (.A1(net6685),
    .A2(_16944_),
    .Y(_01230_),
    .B1(_16942_));
 sg13g2_nand2_1 _48027_ (.Y(_16945_),
    .A(net1123),
    .B(_16936_));
 sg13g2_nor2b_1 _48028_ (.A(_15239_),
    .B_N(net1123),
    .Y(_16946_));
 sg13g2_xnor2_1 _48029_ (.Y(_16947_),
    .A(_15239_),
    .B(_16945_));
 sg13g2_a221oi_1 _48030_ (.B2(net5346),
    .C1(net6610),
    .B1(_16947_),
    .A1(_15239_),
    .Y(_16948_),
    .A2(net5177));
 sg13g2_a21oi_1 _48031_ (.A1(_18315_),
    .A2(net6610),
    .Y(_01231_),
    .B1(_16948_));
 sg13g2_nor2_1 _48032_ (.A(net2276),
    .B(net6682),
    .Y(_16949_));
 sg13g2_a21oi_1 _48033_ (.A1(_16936_),
    .A2(_16946_),
    .Y(_16950_),
    .B1(net5324));
 sg13g2_nor2_1 _48034_ (.A(net5177),
    .B(_16950_),
    .Y(_16951_));
 sg13g2_xnor2_1 _48035_ (.Y(_16952_),
    .A(_15234_),
    .B(_16951_));
 sg13g2_a21oi_1 _48036_ (.A1(net6683),
    .A2(_16952_),
    .Y(_01232_),
    .B1(_16949_));
 sg13g2_nor2_1 _48037_ (.A(net1681),
    .B(net6683),
    .Y(_16953_));
 sg13g2_xnor2_1 _48038_ (.Y(_16954_),
    .A(net5346),
    .B(_15234_));
 sg13g2_nor3_1 _48039_ (.A(net5177),
    .B(_16950_),
    .C(_16954_),
    .Y(_16955_));
 sg13g2_nand3_1 _48040_ (.B(_15233_),
    .C(_16946_),
    .A(_15207_),
    .Y(_16956_));
 sg13g2_nor3_1 _48041_ (.A(_16923_),
    .B(_16935_),
    .C(_16956_),
    .Y(_16957_));
 sg13g2_xor2_1 _48042_ (.B(_16955_),
    .A(_15207_),
    .X(_16958_));
 sg13g2_a21oi_1 _48043_ (.A1(net6683),
    .A2(_16958_),
    .Y(_01233_),
    .B1(_16953_));
 sg13g2_nor2_1 _48044_ (.A(net1933),
    .B(net6686),
    .Y(_16959_));
 sg13g2_nor4_1 _48045_ (.A(net5323),
    .B(_16923_),
    .C(_16935_),
    .D(_16956_),
    .Y(_16960_));
 sg13g2_nor2_1 _48046_ (.A(net5305),
    .B(_16960_),
    .Y(_16961_));
 sg13g2_xnor2_1 _48047_ (.Y(_16962_),
    .A(_15235_),
    .B(_16961_));
 sg13g2_a21oi_1 _48048_ (.A1(net6682),
    .A2(_16962_),
    .Y(_01234_),
    .B1(_16959_));
 sg13g2_nand2_1 _48049_ (.Y(_16963_),
    .A(_15235_),
    .B(_16957_));
 sg13g2_nor2_1 _48050_ (.A(net1904),
    .B(net6686),
    .Y(_16964_));
 sg13g2_nor2b_1 _48051_ (.A(_15231_),
    .B_N(_15235_),
    .Y(_16965_));
 sg13g2_nor2_1 _48052_ (.A(_15231_),
    .B(_16963_),
    .Y(_16966_));
 sg13g2_xnor2_1 _48053_ (.Y(_16967_),
    .A(_15231_),
    .B(_16963_));
 sg13g2_a22oi_1 _48054_ (.Y(_16968_),
    .B1(_16967_),
    .B2(net5357),
    .A2(net5177),
    .A1(_15231_));
 sg13g2_a21oi_1 _48055_ (.A1(net6686),
    .A2(_16968_),
    .Y(_01235_),
    .B1(_16964_));
 sg13g2_nor2_1 _48056_ (.A(net1880),
    .B(net6687),
    .Y(_16969_));
 sg13g2_o21ai_1 _48057_ (.B1(net5169),
    .Y(_16970_),
    .A1(net5325),
    .A2(_16966_));
 sg13g2_xnor2_1 _48058_ (.Y(_16971_),
    .A(_15202_),
    .B(_16970_));
 sg13g2_a21oi_1 _48059_ (.A1(net6686),
    .A2(_16971_),
    .Y(_01236_),
    .B1(_16969_));
 sg13g2_nand4_1 _48060_ (.B(_15202_),
    .C(_16957_),
    .A(_15191_),
    .Y(_16972_),
    .D(_16965_));
 sg13g2_and2_1 _48061_ (.A(_15202_),
    .B(_16966_),
    .X(_16973_));
 sg13g2_o21ai_1 _48062_ (.B1(_16972_),
    .Y(_16974_),
    .A1(_15191_),
    .A2(_16973_));
 sg13g2_o21ai_1 _48063_ (.B1(net6689),
    .Y(_16975_),
    .A1(_15191_),
    .A2(net5169));
 sg13g2_a21oi_1 _48064_ (.A1(net5348),
    .A2(_16974_),
    .Y(_16976_),
    .B1(_16975_));
 sg13g2_a21oi_1 _48065_ (.A1(_18319_),
    .A2(net6612),
    .Y(_01237_),
    .B1(_16976_));
 sg13g2_nor2_1 _48066_ (.A(net2259),
    .B(net6689),
    .Y(_16977_));
 sg13g2_a21o_1 _48067_ (.A2(_16972_),
    .A1(net5348),
    .B1(net5177),
    .X(_16978_));
 sg13g2_xor2_1 _48068_ (.B(_16978_),
    .A(_15187_),
    .X(_16979_));
 sg13g2_a21oi_1 _48069_ (.A1(net6689),
    .A2(_16979_),
    .Y(_01238_),
    .B1(_16977_));
 sg13g2_or3_1 _48070_ (.A(_15186_),
    .B(_15187_),
    .C(_16972_),
    .X(_16980_));
 sg13g2_nand2_1 _48071_ (.Y(_16981_),
    .A(_15188_),
    .B(_16980_));
 sg13g2_a221oi_1 _48072_ (.B2(net5348),
    .C1(net6611),
    .B1(_16981_),
    .A1(_15186_),
    .Y(_16982_),
    .A2(_16978_));
 sg13g2_a21oi_1 _48073_ (.A1(_18321_),
    .A2(net6612),
    .Y(_01239_),
    .B1(_16982_));
 sg13g2_nor2_1 _48074_ (.A(net2098),
    .B(net6687),
    .Y(_16983_));
 sg13g2_a21o_1 _48075_ (.A2(_16980_),
    .A1(net5347),
    .B1(net5177),
    .X(_16984_));
 sg13g2_xnor2_1 _48076_ (.Y(_16985_),
    .A(_15200_),
    .B(_16984_));
 sg13g2_a21oi_1 _48077_ (.A1(net6683),
    .A2(_16985_),
    .Y(_01240_),
    .B1(_16983_));
 sg13g2_nor2_1 _48078_ (.A(net2868),
    .B(net6686),
    .Y(_16986_));
 sg13g2_nor2_1 _48079_ (.A(net5324),
    .B(_15200_),
    .Y(_16987_));
 sg13g2_nor2_2 _48080_ (.A(_16987_),
    .B(_16984_),
    .Y(_16988_));
 sg13g2_xor2_1 _48081_ (.B(_16988_),
    .A(_15183_),
    .X(_16989_));
 sg13g2_a21oi_2 _48082_ (.B1(_16986_),
    .Y(_01241_),
    .A2(net6686),
    .A1(_16989_));
 sg13g2_nand2_1 _48083_ (.Y(_16990_),
    .A(_15183_),
    .B(_15200_));
 sg13g2_nor2_1 _48084_ (.A(_16980_),
    .B(_16990_),
    .Y(_16991_));
 sg13g2_or2_1 _48085_ (.X(_16992_),
    .B(_16990_),
    .A(_16980_));
 sg13g2_nand2_1 _48086_ (.Y(_16993_),
    .A(net5348),
    .B(_16991_));
 sg13g2_nor2_1 _48087_ (.A(_15180_),
    .B(net5305),
    .Y(_16994_));
 sg13g2_and2_1 _48088_ (.A(_15180_),
    .B(_16991_),
    .X(_16995_));
 sg13g2_a221oi_1 _48089_ (.B2(net5348),
    .C1(net6612),
    .B1(_16995_),
    .A1(_16993_),
    .Y(_16996_),
    .A2(_16994_));
 sg13g2_a21oi_1 _48090_ (.A1(_18326_),
    .A2(net6613),
    .Y(_01242_),
    .B1(_16996_));
 sg13g2_nor2_1 _48091_ (.A(net2002),
    .B(net6687),
    .Y(_16997_));
 sg13g2_and2_1 _48092_ (.A(_15198_),
    .B(_16995_),
    .X(_16998_));
 sg13g2_xnor2_1 _48093_ (.Y(_16999_),
    .A(_15198_),
    .B(_16995_));
 sg13g2_a22oi_1 _48094_ (.Y(_17000_),
    .B1(_16999_),
    .B2(net5357),
    .A2(net5177),
    .A1(_15199_));
 sg13g2_a21oi_1 _48095_ (.A1(net6686),
    .A2(_17000_),
    .Y(_01243_),
    .B1(_16997_));
 sg13g2_nor2_1 _48096_ (.A(net1644),
    .B(net6687),
    .Y(_17001_));
 sg13g2_o21ai_1 _48097_ (.B1(net5169),
    .Y(_17002_),
    .A1(net5325),
    .A2(_16998_));
 sg13g2_xnor2_1 _48098_ (.Y(_17003_),
    .A(_15174_),
    .B(_17002_));
 sg13g2_a21oi_1 _48099_ (.A1(net6687),
    .A2(_17003_),
    .Y(_01244_),
    .B1(_17001_));
 sg13g2_nor2_1 _48100_ (.A(_15174_),
    .B(net5306),
    .Y(_17004_));
 sg13g2_nand3_1 _48101_ (.B(_15180_),
    .C(_15198_),
    .A(_15174_),
    .Y(_17005_));
 sg13g2_o21ai_1 _48102_ (.B1(_15196_),
    .Y(_17006_),
    .A1(_17002_),
    .A2(_17004_));
 sg13g2_or2_1 _48103_ (.X(_17007_),
    .B(_17005_),
    .A(_15196_));
 sg13g2_nor2_1 _48104_ (.A(_16993_),
    .B(_17007_),
    .Y(_17008_));
 sg13g2_nor2_1 _48105_ (.A(net6612),
    .B(_17008_),
    .Y(_17009_));
 sg13g2_a22oi_1 _48106_ (.Y(_01245_),
    .B1(_17006_),
    .B2(_17009_),
    .A2(net6612),
    .A1(_18327_));
 sg13g2_nor2_1 _48107_ (.A(net1965),
    .B(net6688),
    .Y(_17010_));
 sg13g2_nor2_1 _48108_ (.A(net5305),
    .B(_17008_),
    .Y(_17011_));
 sg13g2_xor2_1 _48109_ (.B(_17011_),
    .A(_15179_),
    .X(_17012_));
 sg13g2_a21oi_1 _48110_ (.A1(net6686),
    .A2(_17012_),
    .Y(_01246_),
    .B1(_17010_));
 sg13g2_nor4_1 _48111_ (.A(_15177_),
    .B(_15179_),
    .C(_16992_),
    .D(_17007_),
    .Y(_17013_));
 sg13g2_nor3_1 _48112_ (.A(_15179_),
    .B(_16992_),
    .C(_17007_),
    .Y(_17014_));
 sg13g2_nor2b_1 _48113_ (.A(_17014_),
    .B_N(_15177_),
    .Y(_17015_));
 sg13g2_o21ai_1 _48114_ (.B1(net5348),
    .Y(_17016_),
    .A1(_17013_),
    .A2(_17015_));
 sg13g2_a21oi_1 _48115_ (.A1(_15177_),
    .A2(net5178),
    .Y(_17017_),
    .B1(net6612));
 sg13g2_a22oi_1 _48116_ (.Y(_01247_),
    .B1(_17016_),
    .B2(_17017_),
    .A2(net6612),
    .A1(_18329_));
 sg13g2_o21ai_1 _48117_ (.B1(net5170),
    .Y(_17018_),
    .A1(net5325),
    .A2(_17013_));
 sg13g2_xnor2_1 _48118_ (.Y(_17019_),
    .A(_15171_),
    .B(_17018_));
 sg13g2_nor2_1 _48119_ (.A(net2193),
    .B(net6688),
    .Y(_17020_));
 sg13g2_a21oi_1 _48120_ (.A1(net6688),
    .A2(_17019_),
    .Y(_01248_),
    .B1(_17020_));
 sg13g2_nor2_1 _48121_ (.A(net1508),
    .B(net6688),
    .Y(_17021_));
 sg13g2_xnor2_1 _48122_ (.Y(_17022_),
    .A(net5325),
    .B(_15171_));
 sg13g2_nor2_1 _48123_ (.A(_17018_),
    .B(_17022_),
    .Y(_17023_));
 sg13g2_xor2_1 _48124_ (.B(_17023_),
    .A(_15175_),
    .X(_17024_));
 sg13g2_a21oi_1 _48125_ (.A1(net6688),
    .A2(_17024_),
    .Y(_01249_),
    .B1(_17021_));
 sg13g2_a21oi_1 _48126_ (.A1(net7088),
    .A2(net6205),
    .Y(_17025_),
    .B1(net6388));
 sg13g2_nand3_1 _48127_ (.B(net7095),
    .C(net6062),
    .A(net2703),
    .Y(_17026_));
 sg13g2_o21ai_1 _48128_ (.B1(_17026_),
    .Y(_01250_),
    .A1(_18357_),
    .A2(net6062));
 sg13g2_nand3_1 _48129_ (.B(net7095),
    .C(net6062),
    .A(net1680),
    .Y(_17027_));
 sg13g2_o21ai_1 _48130_ (.B1(_17027_),
    .Y(_01251_),
    .A1(_18613_),
    .A2(net6062));
 sg13g2_nand3_1 _48131_ (.B(net7095),
    .C(net6062),
    .A(net2514),
    .Y(_17028_));
 sg13g2_o21ai_1 _48132_ (.B1(_17028_),
    .Y(_01252_),
    .A1(_18612_),
    .A2(net6062));
 sg13g2_nand3_1 _48133_ (.B(net7097),
    .C(net6062),
    .A(net2974),
    .Y(_17029_));
 sg13g2_o21ai_1 _48134_ (.B1(_17029_),
    .Y(_01253_),
    .A1(_18611_),
    .A2(net6062));
 sg13g2_nand3_1 _48135_ (.B(net7097),
    .C(net6063),
    .A(net2819),
    .Y(_17030_));
 sg13g2_o21ai_1 _48136_ (.B1(_17030_),
    .Y(_01254_),
    .A1(_18610_),
    .A2(net6063));
 sg13g2_nand3_1 _48137_ (.B(net7097),
    .C(net6063),
    .A(net2464),
    .Y(_17031_));
 sg13g2_o21ai_1 _48138_ (.B1(_17031_),
    .Y(_01255_),
    .A1(_18609_),
    .A2(net6063));
 sg13g2_nand3_1 _48139_ (.B(net7097),
    .C(net6063),
    .A(net2805),
    .Y(_17032_));
 sg13g2_o21ai_1 _48140_ (.B1(_17032_),
    .Y(_01256_),
    .A1(_18608_),
    .A2(net6063));
 sg13g2_nand3_1 _48141_ (.B(net7096),
    .C(net6063),
    .A(net2736),
    .Y(_17033_));
 sg13g2_o21ai_1 _48142_ (.B1(_17033_),
    .Y(_01257_),
    .A1(_18607_),
    .A2(net6063));
 sg13g2_nand3_1 _48143_ (.B(net7096),
    .C(net6081),
    .A(net1823),
    .Y(_17034_));
 sg13g2_o21ai_1 _48144_ (.B1(_17034_),
    .Y(_01258_),
    .A1(_18606_),
    .A2(net6080));
 sg13g2_nand3_1 _48145_ (.B(net7097),
    .C(net6081),
    .A(net3145),
    .Y(_17035_));
 sg13g2_o21ai_1 _48146_ (.B1(_17035_),
    .Y(_01259_),
    .A1(_18605_),
    .A2(net6081));
 sg13g2_nand3_1 _48147_ (.B(net7096),
    .C(net6077),
    .A(net2977),
    .Y(_17036_));
 sg13g2_o21ai_1 _48148_ (.B1(_17036_),
    .Y(_01260_),
    .A1(_18604_),
    .A2(net6077));
 sg13g2_nand3_1 _48149_ (.B(net7096),
    .C(net6080),
    .A(net1389),
    .Y(_17037_));
 sg13g2_o21ai_1 _48150_ (.B1(_17037_),
    .Y(_01261_),
    .A1(_18603_),
    .A2(net6080));
 sg13g2_nand3_1 _48151_ (.B(net7104),
    .C(net6079),
    .A(net2807),
    .Y(_17038_));
 sg13g2_o21ai_1 _48152_ (.B1(_17038_),
    .Y(_01262_),
    .A1(_18602_),
    .A2(net6079));
 sg13g2_nand3_1 _48153_ (.B(net7104),
    .C(net6079),
    .A(net2482),
    .Y(_17039_));
 sg13g2_o21ai_1 _48154_ (.B1(_17039_),
    .Y(_01263_),
    .A1(_18601_),
    .A2(net6079));
 sg13g2_nand3_1 _48155_ (.B(net7104),
    .C(net6078),
    .A(net2945),
    .Y(_17040_));
 sg13g2_o21ai_1 _48156_ (.B1(_17040_),
    .Y(_01264_),
    .A1(_18600_),
    .A2(net6079));
 sg13g2_nand3_1 _48157_ (.B(net7104),
    .C(net6081),
    .A(net2797),
    .Y(_17041_));
 sg13g2_o21ai_1 _48158_ (.B1(_17041_),
    .Y(_01265_),
    .A1(_18599_),
    .A2(net6079));
 sg13g2_nand3_1 _48159_ (.B(net7107),
    .C(net6084),
    .A(net3078),
    .Y(_17042_));
 sg13g2_o21ai_1 _48160_ (.B1(_17042_),
    .Y(_01266_),
    .A1(_18598_),
    .A2(net6084));
 sg13g2_nand3_1 _48161_ (.B(net7107),
    .C(net6084),
    .A(net2968),
    .Y(_17043_));
 sg13g2_o21ai_1 _48162_ (.B1(_17043_),
    .Y(_01267_),
    .A1(_18597_),
    .A2(net6084));
 sg13g2_nand3_1 _48163_ (.B(net7104),
    .C(net6084),
    .A(net7299),
    .Y(_17044_));
 sg13g2_o21ai_1 _48164_ (.B1(_17044_),
    .Y(_01268_),
    .A1(_18596_),
    .A2(net6084));
 sg13g2_nand3_1 _48165_ (.B(net7104),
    .C(net6084),
    .A(net3383),
    .Y(_17045_));
 sg13g2_o21ai_1 _48166_ (.B1(_17045_),
    .Y(_01269_),
    .A1(_18595_),
    .A2(net6085));
 sg13g2_nand3_1 _48167_ (.B(net7106),
    .C(net6084),
    .A(net3293),
    .Y(_17046_));
 sg13g2_o21ai_1 _48168_ (.B1(_17046_),
    .Y(_01270_),
    .A1(_18594_),
    .A2(net6085));
 sg13g2_nand3_1 _48169_ (.B(net7105),
    .C(net6083),
    .A(net3080),
    .Y(_17047_));
 sg13g2_o21ai_1 _48170_ (.B1(_17047_),
    .Y(_01271_),
    .A1(_18593_),
    .A2(net6083));
 sg13g2_nand3_1 _48171_ (.B(net7105),
    .C(net6082),
    .A(net3210),
    .Y(_17048_));
 sg13g2_o21ai_1 _48172_ (.B1(_17048_),
    .Y(_01272_),
    .A1(_18592_),
    .A2(net6083));
 sg13g2_nand3_1 _48173_ (.B(net7105),
    .C(net6082),
    .A(net3142),
    .Y(_17049_));
 sg13g2_o21ai_1 _48174_ (.B1(_17049_),
    .Y(_01273_),
    .A1(_18591_),
    .A2(net6083));
 sg13g2_nand3_1 _48175_ (.B(net7106),
    .C(net6085),
    .A(net2537),
    .Y(_17050_));
 sg13g2_o21ai_1 _48176_ (.B1(_17050_),
    .Y(_01274_),
    .A1(_18590_),
    .A2(net6086));
 sg13g2_nand3_1 _48177_ (.B(net7106),
    .C(net6085),
    .A(net2948),
    .Y(_17051_));
 sg13g2_o21ai_1 _48178_ (.B1(_17051_),
    .Y(_01275_),
    .A1(_18589_),
    .A2(net6085));
 sg13g2_nand3_1 _48179_ (.B(net7106),
    .C(net6085),
    .A(net3133),
    .Y(_17052_));
 sg13g2_o21ai_1 _48180_ (.B1(_17052_),
    .Y(_01276_),
    .A1(_18588_),
    .A2(net6085));
 sg13g2_nand3_1 _48181_ (.B(net7106),
    .C(net6100),
    .A(net2038),
    .Y(_17053_));
 sg13g2_o21ai_1 _48182_ (.B1(_17053_),
    .Y(_01277_),
    .A1(_18587_),
    .A2(net6100));
 sg13g2_nand3_1 _48183_ (.B(net7106),
    .C(net6100),
    .A(net2268),
    .Y(_17054_));
 sg13g2_o21ai_1 _48184_ (.B1(_17054_),
    .Y(_01278_),
    .A1(_18586_),
    .A2(net6100));
 sg13g2_nand3_1 _48185_ (.B(net7114),
    .C(net6100),
    .A(net1915),
    .Y(_17055_));
 sg13g2_o21ai_1 _48186_ (.B1(_17055_),
    .Y(_01279_),
    .A1(_18585_),
    .A2(net6100));
 sg13g2_nand3_1 _48187_ (.B(net7114),
    .C(net6100),
    .A(net3471),
    .Y(_17056_));
 sg13g2_o21ai_1 _48188_ (.B1(_17056_),
    .Y(_01280_),
    .A1(_18584_),
    .A2(net6100));
 sg13g2_nand3_1 _48189_ (.B(net7115),
    .C(net6101),
    .A(net1742),
    .Y(_17057_));
 sg13g2_o21ai_1 _48190_ (.B1(_17057_),
    .Y(_01281_),
    .A1(_18583_),
    .A2(net6101));
 sg13g2_nand3_1 _48191_ (.B(net7116),
    .C(net6107),
    .A(net2100),
    .Y(_17058_));
 sg13g2_o21ai_1 _48192_ (.B1(_17058_),
    .Y(_01282_),
    .A1(_18582_),
    .A2(net6107));
 sg13g2_nand3_1 _48193_ (.B(net7116),
    .C(net6108),
    .A(net3096),
    .Y(_17059_));
 sg13g2_o21ai_1 _48194_ (.B1(_17059_),
    .Y(_01283_),
    .A1(_18581_),
    .A2(net6108));
 sg13g2_nand3_1 _48195_ (.B(net7116),
    .C(net6108),
    .A(net1955),
    .Y(_17060_));
 sg13g2_o21ai_1 _48196_ (.B1(_17060_),
    .Y(_01284_),
    .A1(_18580_),
    .A2(net6108));
 sg13g2_nand3_1 _48197_ (.B(net7117),
    .C(net6108),
    .A(net2646),
    .Y(_17061_));
 sg13g2_o21ai_1 _48198_ (.B1(_17061_),
    .Y(_01285_),
    .A1(_18579_),
    .A2(net6108));
 sg13g2_nand3_1 _48199_ (.B(net7116),
    .C(net6109),
    .A(net2705),
    .Y(_17062_));
 sg13g2_o21ai_1 _48200_ (.B1(_17062_),
    .Y(_01286_),
    .A1(_18578_),
    .A2(net6109));
 sg13g2_nand3_1 _48201_ (.B(net7116),
    .C(net6108),
    .A(net2764),
    .Y(_17063_));
 sg13g2_o21ai_1 _48202_ (.B1(_17063_),
    .Y(_01287_),
    .A1(_18577_),
    .A2(net6109));
 sg13g2_nand3_1 _48203_ (.B(net7116),
    .C(net6109),
    .A(net2762),
    .Y(_17064_));
 sg13g2_o21ai_1 _48204_ (.B1(_17064_),
    .Y(_01288_),
    .A1(_18576_),
    .A2(net6108));
 sg13g2_nand3_1 _48205_ (.B(net7116),
    .C(net6109),
    .A(net3163),
    .Y(_17065_));
 sg13g2_o21ai_1 _48206_ (.B1(_17065_),
    .Y(_01289_),
    .A1(_18575_),
    .A2(net6109));
 sg13g2_nand3_1 _48207_ (.B(net7116),
    .C(net6121),
    .A(net3323),
    .Y(_17066_));
 sg13g2_o21ai_1 _48208_ (.B1(_17066_),
    .Y(_01290_),
    .A1(_18574_),
    .A2(net6121));
 sg13g2_nand3_1 _48209_ (.B(net7121),
    .C(net6121),
    .A(net3416),
    .Y(_17067_));
 sg13g2_o21ai_1 _48210_ (.B1(_17067_),
    .Y(_01291_),
    .A1(_18573_),
    .A2(net6121));
 sg13g2_nand3_1 _48211_ (.B(net7121),
    .C(net6121),
    .A(net1724),
    .Y(_17068_));
 sg13g2_o21ai_1 _48212_ (.B1(_17068_),
    .Y(_01292_),
    .A1(_18572_),
    .A2(net6122));
 sg13g2_nand3_1 _48213_ (.B(net7121),
    .C(net6121),
    .A(net3011),
    .Y(_17069_));
 sg13g2_o21ai_1 _48214_ (.B1(_17069_),
    .Y(_01293_),
    .A1(_18571_),
    .A2(net6122));
 sg13g2_nand3_1 _48215_ (.B(net7121),
    .C(net6121),
    .A(net3124),
    .Y(_17070_));
 sg13g2_o21ai_1 _48216_ (.B1(_17070_),
    .Y(_01294_),
    .A1(_18570_),
    .A2(net6121));
 sg13g2_nand3_1 _48217_ (.B(net7121),
    .C(net6122),
    .A(net3353),
    .Y(_17071_));
 sg13g2_o21ai_1 _48218_ (.B1(_17071_),
    .Y(_01295_),
    .A1(_18569_),
    .A2(net6122));
 sg13g2_nand3_1 _48219_ (.B(net7128),
    .C(net6134),
    .A(net2662),
    .Y(_17072_));
 sg13g2_o21ai_1 _48220_ (.B1(_17072_),
    .Y(_01296_),
    .A1(_18568_),
    .A2(net6134));
 sg13g2_nand3_1 _48221_ (.B(net7128),
    .C(net6134),
    .A(net3045),
    .Y(_17073_));
 sg13g2_o21ai_1 _48222_ (.B1(_17073_),
    .Y(_01297_),
    .A1(_18567_),
    .A2(net6134));
 sg13g2_nand3_1 _48223_ (.B(net7121),
    .C(net6124),
    .A(net2480),
    .Y(_17074_));
 sg13g2_o21ai_1 _48224_ (.B1(_17074_),
    .Y(_01298_),
    .A1(_18566_),
    .A2(net6124));
 sg13g2_nand3_1 _48225_ (.B(net7121),
    .C(net6124),
    .A(net2916),
    .Y(_17075_));
 sg13g2_o21ai_1 _48226_ (.B1(_17075_),
    .Y(_01299_),
    .A1(_18565_),
    .A2(net6124));
 sg13g2_nand3_1 _48227_ (.B(net7121),
    .C(net6124),
    .A(net1238),
    .Y(_17076_));
 sg13g2_o21ai_1 _48228_ (.B1(_17076_),
    .Y(_01300_),
    .A1(_18564_),
    .A2(net6124));
 sg13g2_nand3_1 _48229_ (.B(net7122),
    .C(net6130),
    .A(net3579),
    .Y(_17077_));
 sg13g2_o21ai_1 _48230_ (.B1(_17077_),
    .Y(_01301_),
    .A1(_18563_),
    .A2(net6130));
 sg13g2_nand3_1 _48231_ (.B(net7124),
    .C(net6131),
    .A(net3408),
    .Y(_17078_));
 sg13g2_o21ai_1 _48232_ (.B1(_17078_),
    .Y(_01302_),
    .A1(_18562_),
    .A2(net6131));
 sg13g2_nand3_1 _48233_ (.B(net7124),
    .C(net6130),
    .A(net3236),
    .Y(_17079_));
 sg13g2_o21ai_1 _48234_ (.B1(_17079_),
    .Y(_01303_),
    .A1(_18561_),
    .A2(net6130));
 sg13g2_nand3_1 _48235_ (.B(net7125),
    .C(net6138),
    .A(net2910),
    .Y(_17080_));
 sg13g2_o21ai_1 _48236_ (.B1(_17080_),
    .Y(_01304_),
    .A1(_18560_),
    .A2(net6138));
 sg13g2_nand3_1 _48237_ (.B(net7125),
    .C(net6138),
    .A(net2483),
    .Y(_17081_));
 sg13g2_o21ai_1 _48238_ (.B1(_17081_),
    .Y(_01305_),
    .A1(_18559_),
    .A2(net6138));
 sg13g2_nand3_1 _48239_ (.B(net7125),
    .C(net6136),
    .A(net3583),
    .Y(_17082_));
 sg13g2_o21ai_1 _48240_ (.B1(_17082_),
    .Y(_01306_),
    .A1(_18558_),
    .A2(net6136));
 sg13g2_nand3_1 _48241_ (.B(net7125),
    .C(net6136),
    .A(\u_inv.d_next[57] ),
    .Y(_17083_));
 sg13g2_o21ai_1 _48242_ (.B1(_17083_),
    .Y(_01307_),
    .A1(_18557_),
    .A2(net6136));
 sg13g2_nand3_1 _48243_ (.B(net7125),
    .C(net6136),
    .A(net2614),
    .Y(_17084_));
 sg13g2_o21ai_1 _48244_ (.B1(_17084_),
    .Y(_01308_),
    .A1(_18556_),
    .A2(net6136));
 sg13g2_nand3_1 _48245_ (.B(net7127),
    .C(net6137),
    .A(net2979),
    .Y(_17085_));
 sg13g2_o21ai_1 _48246_ (.B1(_17085_),
    .Y(_01309_),
    .A1(_18555_),
    .A2(net6137));
 sg13g2_nand3_1 _48247_ (.B(net7125),
    .C(net6137),
    .A(net2120),
    .Y(_17086_));
 sg13g2_o21ai_1 _48248_ (.B1(_17086_),
    .Y(_01310_),
    .A1(_18554_),
    .A2(net6156));
 sg13g2_nand3_1 _48249_ (.B(net7125),
    .C(net6136),
    .A(net3074),
    .Y(_17087_));
 sg13g2_o21ai_1 _48250_ (.B1(_17087_),
    .Y(_01311_),
    .A1(_18553_),
    .A2(net6136));
 sg13g2_nand3_1 _48251_ (.B(net7125),
    .C(net6137),
    .A(net2436),
    .Y(_17088_));
 sg13g2_o21ai_1 _48252_ (.B1(_17088_),
    .Y(_01312_),
    .A1(_18552_),
    .A2(net6156));
 sg13g2_nand3_1 _48253_ (.B(net7127),
    .C(net6137),
    .A(net3009),
    .Y(_17089_));
 sg13g2_o21ai_1 _48254_ (.B1(_17089_),
    .Y(_01313_),
    .A1(_18551_),
    .A2(net6137));
 sg13g2_nand3_1 _48255_ (.B(net7142),
    .C(net6183),
    .A(net2253),
    .Y(_17090_));
 sg13g2_o21ai_1 _48256_ (.B1(_17090_),
    .Y(_01314_),
    .A1(_18550_),
    .A2(net6183));
 sg13g2_nand3_1 _48257_ (.B(net7142),
    .C(net6183),
    .A(net2814),
    .Y(_17091_));
 sg13g2_o21ai_1 _48258_ (.B1(_17091_),
    .Y(_01315_),
    .A1(_18549_),
    .A2(net6183));
 sg13g2_nand3_1 _48259_ (.B(net7142),
    .C(net6185),
    .A(net2521),
    .Y(_17092_));
 sg13g2_o21ai_1 _48260_ (.B1(_17092_),
    .Y(_01316_),
    .A1(_18548_),
    .A2(net6183));
 sg13g2_nand3_1 _48261_ (.B(net7142),
    .C(net6183),
    .A(net3199),
    .Y(_17093_));
 sg13g2_o21ai_1 _48262_ (.B1(_17093_),
    .Y(_01317_),
    .A1(_18547_),
    .A2(net6183));
 sg13g2_nand3_1 _48263_ (.B(net7142),
    .C(net6183),
    .A(net3340),
    .Y(_17094_));
 sg13g2_o21ai_1 _48264_ (.B1(_17094_),
    .Y(_01318_),
    .A1(_18546_),
    .A2(net6169));
 sg13g2_nand3_1 _48265_ (.B(net7145),
    .C(net6189),
    .A(net3239),
    .Y(_17095_));
 sg13g2_o21ai_1 _48266_ (.B1(_17095_),
    .Y(_01319_),
    .A1(_18545_),
    .A2(net6189));
 sg13g2_nand3_1 _48267_ (.B(net7138),
    .C(net6189),
    .A(net7297),
    .Y(_17096_));
 sg13g2_o21ai_1 _48268_ (.B1(_17096_),
    .Y(_01320_),
    .A1(_18544_),
    .A2(net6169));
 sg13g2_nand3_1 _48269_ (.B(net7138),
    .C(net6169),
    .A(net2804),
    .Y(_17097_));
 sg13g2_o21ai_1 _48270_ (.B1(_17097_),
    .Y(_01321_),
    .A1(_18543_),
    .A2(net6169));
 sg13g2_nand3_1 _48271_ (.B(net7145),
    .C(net6189),
    .A(net3523),
    .Y(_17098_));
 sg13g2_o21ai_1 _48272_ (.B1(_17098_),
    .Y(_01322_),
    .A1(_18542_),
    .A2(net6180));
 sg13g2_nand3_1 _48273_ (.B(net7145),
    .C(net6189),
    .A(net3260),
    .Y(_17099_));
 sg13g2_o21ai_1 _48274_ (.B1(_17099_),
    .Y(_01323_),
    .A1(_18541_),
    .A2(net6189));
 sg13g2_nand3_1 _48275_ (.B(net7139),
    .C(net6179),
    .A(net3477),
    .Y(_17100_));
 sg13g2_o21ai_1 _48276_ (.B1(_17100_),
    .Y(_01324_),
    .A1(_18540_),
    .A2(net6179));
 sg13g2_nand3_1 _48277_ (.B(net7139),
    .C(net6179),
    .A(net3393),
    .Y(_17101_));
 sg13g2_o21ai_1 _48278_ (.B1(_17101_),
    .Y(_01325_),
    .A1(_18539_),
    .A2(net6179));
 sg13g2_nand3_1 _48279_ (.B(net7138),
    .C(net6181),
    .A(net2585),
    .Y(_17102_));
 sg13g2_o21ai_1 _48280_ (.B1(_17102_),
    .Y(_01326_),
    .A1(_18538_),
    .A2(net6181));
 sg13g2_nand3_1 _48281_ (.B(net7139),
    .C(net6180),
    .A(net1849),
    .Y(_17103_));
 sg13g2_o21ai_1 _48282_ (.B1(_17103_),
    .Y(_01327_),
    .A1(_18537_),
    .A2(net6181));
 sg13g2_nand3_1 _48283_ (.B(net7139),
    .C(net6180),
    .A(net3274),
    .Y(_17104_));
 sg13g2_o21ai_1 _48284_ (.B1(_17104_),
    .Y(_01328_),
    .A1(_18536_),
    .A2(net6180));
 sg13g2_nand3_1 _48285_ (.B(net7138),
    .C(net6181),
    .A(net2325),
    .Y(_17105_));
 sg13g2_o21ai_1 _48286_ (.B1(_17105_),
    .Y(_01329_),
    .A1(_18535_),
    .A2(net6181));
 sg13g2_nand3_1 _48287_ (.B(net7141),
    .C(net6169),
    .A(net2366),
    .Y(_17106_));
 sg13g2_o21ai_1 _48288_ (.B1(_17106_),
    .Y(_01330_),
    .A1(_18534_),
    .A2(net6168));
 sg13g2_nand3_1 _48289_ (.B(net7142),
    .C(net6185),
    .A(\u_inv.d_next[81] ),
    .Y(_17107_));
 sg13g2_o21ai_1 _48290_ (.B1(_17107_),
    .Y(_01331_),
    .A1(_18533_),
    .A2(net6168));
 sg13g2_nand3_1 _48291_ (.B(net7141),
    .C(net6168),
    .A(net2746),
    .Y(_17108_));
 sg13g2_o21ai_1 _48292_ (.B1(_17108_),
    .Y(_01332_),
    .A1(_18532_),
    .A2(net6168));
 sg13g2_nand3_1 _48293_ (.B(net7133),
    .C(net6153),
    .A(net3462),
    .Y(_17109_));
 sg13g2_o21ai_1 _48294_ (.B1(_17109_),
    .Y(_01333_),
    .A1(_18531_),
    .A2(net6159));
 sg13g2_nand3_1 _48295_ (.B(net7134),
    .C(net6158),
    .A(net3334),
    .Y(_17110_));
 sg13g2_o21ai_1 _48296_ (.B1(_17110_),
    .Y(_01334_),
    .A1(_18530_),
    .A2(net6158));
 sg13g2_nand3_1 _48297_ (.B(net7134),
    .C(net6159),
    .A(net2119),
    .Y(_17111_));
 sg13g2_o21ai_1 _48298_ (.B1(_17111_),
    .Y(_01335_),
    .A1(_18529_),
    .A2(net6159));
 sg13g2_nand3_1 _48299_ (.B(net7134),
    .C(net6158),
    .A(net3510),
    .Y(_17112_));
 sg13g2_o21ai_1 _48300_ (.B1(_17112_),
    .Y(_01336_),
    .A1(_18528_),
    .A2(net6158));
 sg13g2_nand3_1 _48301_ (.B(net7134),
    .C(net6158),
    .A(net3494),
    .Y(_17113_));
 sg13g2_o21ai_1 _48302_ (.B1(_17113_),
    .Y(_01337_),
    .A1(_18527_),
    .A2(net6158));
 sg13g2_nand3_1 _48303_ (.B(net7134),
    .C(net6157),
    .A(net2538),
    .Y(_17114_));
 sg13g2_o21ai_1 _48304_ (.B1(_17114_),
    .Y(_01338_),
    .A1(_18526_),
    .A2(net6157));
 sg13g2_nand3_1 _48305_ (.B(net7134),
    .C(net6157),
    .A(net3566),
    .Y(_17115_));
 sg13g2_o21ai_1 _48306_ (.B1(_17115_),
    .Y(_01339_),
    .A1(_18525_),
    .A2(net6157));
 sg13g2_nand3_1 _48307_ (.B(net7134),
    .C(net6157),
    .A(net2316),
    .Y(_17116_));
 sg13g2_o21ai_1 _48308_ (.B1(_17116_),
    .Y(_01340_),
    .A1(_18524_),
    .A2(net6158));
 sg13g2_nand3_1 _48309_ (.B(net7134),
    .C(net6157),
    .A(net1638),
    .Y(_17117_));
 sg13g2_o21ai_1 _48310_ (.B1(_17117_),
    .Y(_01341_),
    .A1(_18523_),
    .A2(net6157));
 sg13g2_nand3_1 _48311_ (.B(net7135),
    .C(net6160),
    .A(net2475),
    .Y(_17118_));
 sg13g2_o21ai_1 _48312_ (.B1(_17118_),
    .Y(_01342_),
    .A1(_18522_),
    .A2(net6160));
 sg13g2_nand3_1 _48313_ (.B(net7135),
    .C(net6160),
    .A(net3175),
    .Y(_17119_));
 sg13g2_o21ai_1 _48314_ (.B1(_17119_),
    .Y(_01343_),
    .A1(_18521_),
    .A2(net6160));
 sg13g2_nand3_1 _48315_ (.B(net7137),
    .C(net6160),
    .A(net2083),
    .Y(_17120_));
 sg13g2_o21ai_1 _48316_ (.B1(_17120_),
    .Y(_01344_),
    .A1(_18520_),
    .A2(net6160));
 sg13g2_nand3_1 _48317_ (.B(net7136),
    .C(net6159),
    .A(\u_inv.d_next[95] ),
    .Y(_17121_));
 sg13g2_o21ai_1 _48318_ (.B1(_17121_),
    .Y(_01345_),
    .A1(_18519_),
    .A2(net6157));
 sg13g2_nand3_1 _48319_ (.B(net7142),
    .C(net6184),
    .A(net2319),
    .Y(_17122_));
 sg13g2_o21ai_1 _48320_ (.B1(_17122_),
    .Y(_01346_),
    .A1(_18518_),
    .A2(net6184));
 sg13g2_nand3_1 _48321_ (.B(net7146),
    .C(net6184),
    .A(net3652),
    .Y(_17123_));
 sg13g2_o21ai_1 _48322_ (.B1(_17123_),
    .Y(_01347_),
    .A1(_18517_),
    .A2(net6162));
 sg13g2_nand3_1 _48323_ (.B(net7146),
    .C(net6184),
    .A(net2972),
    .Y(_17124_));
 sg13g2_o21ai_1 _48324_ (.B1(_17124_),
    .Y(_01348_),
    .A1(_18516_),
    .A2(net6184));
 sg13g2_nand3_1 _48325_ (.B(net7143),
    .C(net6186),
    .A(net3664),
    .Y(_17125_));
 sg13g2_o21ai_1 _48326_ (.B1(_17125_),
    .Y(_01349_),
    .A1(_18515_),
    .A2(net6184));
 sg13g2_nand3_1 _48327_ (.B(net7143),
    .C(net6186),
    .A(net1701),
    .Y(_17126_));
 sg13g2_o21ai_1 _48328_ (.B1(_17126_),
    .Y(_01350_),
    .A1(_18514_),
    .A2(net6189));
 sg13g2_nand3_1 _48329_ (.B(net7143),
    .C(net6186),
    .A(net3119),
    .Y(_17127_));
 sg13g2_o21ai_1 _48330_ (.B1(_17127_),
    .Y(_01351_),
    .A1(_18513_),
    .A2(net6187));
 sg13g2_nand3_1 _48331_ (.B(net7143),
    .C(net6187),
    .A(net2992),
    .Y(_17128_));
 sg13g2_o21ai_1 _48332_ (.B1(_17128_),
    .Y(_01352_),
    .A1(_18512_),
    .A2(net6186));
 sg13g2_nand3_1 _48333_ (.B(net7143),
    .C(net6186),
    .A(net3342),
    .Y(_17129_));
 sg13g2_o21ai_1 _48334_ (.B1(_17129_),
    .Y(_01353_),
    .A1(_18511_),
    .A2(net6186));
 sg13g2_nand3_1 _48335_ (.B(net7143),
    .C(net6186),
    .A(net2862),
    .Y(_17130_));
 sg13g2_o21ai_1 _48336_ (.B1(_17130_),
    .Y(_01354_),
    .A1(_18510_),
    .A2(net6186));
 sg13g2_nand3_1 _48337_ (.B(net7144),
    .C(net6188),
    .A(net2986),
    .Y(_17131_));
 sg13g2_o21ai_1 _48338_ (.B1(_17131_),
    .Y(_01355_),
    .A1(_18509_),
    .A2(net6188));
 sg13g2_nand3_1 _48339_ (.B(net7144),
    .C(net6188),
    .A(net2663),
    .Y(_17132_));
 sg13g2_o21ai_1 _48340_ (.B1(_17132_),
    .Y(_01356_),
    .A1(_18508_),
    .A2(net6188));
 sg13g2_nand3_1 _48341_ (.B(net7144),
    .C(net6188),
    .A(net2869),
    .Y(_17133_));
 sg13g2_o21ai_1 _48342_ (.B1(_17133_),
    .Y(_01357_),
    .A1(_18507_),
    .A2(net6188));
 sg13g2_nand3_1 _48343_ (.B(net7143),
    .C(net6187),
    .A(net3321),
    .Y(_17134_));
 sg13g2_o21ai_1 _48344_ (.B1(_17134_),
    .Y(_01358_),
    .A1(_18506_),
    .A2(net6187));
 sg13g2_nand3_1 _48345_ (.B(net7143),
    .C(net6187),
    .A(net2665),
    .Y(_17135_));
 sg13g2_o21ai_1 _48346_ (.B1(_17135_),
    .Y(_01359_),
    .A1(_18505_),
    .A2(net6187));
 sg13g2_nand3_1 _48347_ (.B(net7144),
    .C(net6187),
    .A(net2134),
    .Y(_17136_));
 sg13g2_o21ai_1 _48348_ (.B1(_17136_),
    .Y(_01360_),
    .A1(_18504_),
    .A2(net6188));
 sg13g2_nand3_1 _48349_ (.B(net7144),
    .C(net6184),
    .A(\u_inv.d_next[111] ),
    .Y(_17137_));
 sg13g2_o21ai_1 _48350_ (.B1(_17137_),
    .Y(_01361_),
    .A1(_18503_),
    .A2(net6185));
 sg13g2_nand3_1 _48351_ (.B(net7142),
    .C(net6184),
    .A(net3327),
    .Y(_17138_));
 sg13g2_o21ai_1 _48352_ (.B1(_17138_),
    .Y(_01362_),
    .A1(_18502_),
    .A2(net6162));
 sg13g2_nand3_1 _48353_ (.B(net7135),
    .C(net6162),
    .A(net3052),
    .Y(_17139_));
 sg13g2_o21ai_1 _48354_ (.B1(_17139_),
    .Y(_01363_),
    .A1(_18501_),
    .A2(net6163));
 sg13g2_dfrbpq_1 _48355_ (.RESET_B(net7565),
    .D(net1798),
    .Q(\u_inv.input_reg[95] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _48356_ (.RESET_B(net7536),
    .D(net1547),
    .Q(\u_inv.input_reg[96] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _48357_ (.RESET_B(net7537),
    .D(net1366),
    .Q(\u_inv.input_reg[97] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _48358_ (.RESET_B(net7531),
    .D(net1659),
    .Q(\u_inv.input_reg[98] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _48359_ (.RESET_B(net7533),
    .D(net1323),
    .Q(\u_inv.input_reg[99] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _48360_ (.RESET_B(net7536),
    .D(net1946),
    .Q(\u_inv.input_reg[100] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _48361_ (.RESET_B(net7534),
    .D(net1801),
    .Q(\u_inv.input_reg[101] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _48362_ (.RESET_B(net7535),
    .D(net1864),
    .Q(\u_inv.input_reg[102] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _48363_ (.RESET_B(net7531),
    .D(net1410),
    .Q(\u_inv.input_reg[103] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _48364_ (.RESET_B(net7534),
    .D(net1683),
    .Q(\u_inv.input_reg[104] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _48365_ (.RESET_B(net7535),
    .D(net1364),
    .Q(\u_inv.input_reg[105] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _48366_ (.RESET_B(net7534),
    .D(net2371),
    .Q(\u_inv.input_reg[106] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _48367_ (.RESET_B(net7548),
    .D(net1277),
    .Q(\u_inv.input_reg[107] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _48368_ (.RESET_B(net7545),
    .D(net1690),
    .Q(\u_inv.input_reg[108] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _48369_ (.RESET_B(net7530),
    .D(net1763),
    .Q(\u_inv.input_reg[109] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _48370_ (.RESET_B(net7530),
    .D(net1593),
    .Q(\u_inv.input_reg[110] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _48371_ (.RESET_B(net7530),
    .D(net1734),
    .Q(\u_inv.input_reg[111] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _48372_ (.RESET_B(net7540),
    .D(net1398),
    .Q(\u_inv.input_reg[112] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _48373_ (.RESET_B(net7540),
    .D(net1536),
    .Q(\u_inv.input_reg[113] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _48374_ (.RESET_B(net7530),
    .D(net1749),
    .Q(\u_inv.input_reg[114] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _48375_ (.RESET_B(net7540),
    .D(net2016),
    .Q(\u_inv.input_reg[115] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _48376_ (.RESET_B(net7542),
    .D(net2513),
    .Q(\u_inv.input_reg[116] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_1 _48377_ (.RESET_B(net7524),
    .D(net1430),
    .Q(\u_inv.input_reg[117] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_1 _48378_ (.RESET_B(net7540),
    .D(net1729),
    .Q(\u_inv.input_reg[118] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _48379_ (.RESET_B(net7530),
    .D(_00026_),
    .Q(\u_inv.input_reg[119] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _48380_ (.RESET_B(net7542),
    .D(net1317),
    .Q(\u_inv.input_reg[120] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _48381_ (.RESET_B(net7542),
    .D(_00028_),
    .Q(\u_inv.input_reg[121] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _48382_ (.RESET_B(net7529),
    .D(net1657),
    .Q(\u_inv.input_reg[122] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _48383_ (.RESET_B(net7524),
    .D(net1259),
    .Q(\u_inv.input_reg[123] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _48384_ (.RESET_B(net7523),
    .D(net3171),
    .Q(\u_inv.input_reg[124] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _48385_ (.RESET_B(net7523),
    .D(net3166),
    .Q(\u_inv.input_reg[125] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_1 _48386_ (.RESET_B(net7530),
    .D(net2999),
    .Q(\u_inv.input_reg[126] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _48387_ (.RESET_B(net7520),
    .D(net1907),
    .Q(\u_inv.input_reg[127] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _48388_ (.RESET_B(net7520),
    .D(net2318),
    .Q(\u_inv.input_reg[128] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _48389_ (.RESET_B(net7520),
    .D(net1641),
    .Q(\u_inv.input_reg[129] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _48390_ (.RESET_B(net7520),
    .D(net2400),
    .Q(\u_inv.input_reg[130] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _48391_ (.RESET_B(net7525),
    .D(net1382),
    .Q(\u_inv.input_reg[131] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _48392_ (.RESET_B(net7516),
    .D(net1272),
    .Q(\u_inv.input_reg[132] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_1 _48393_ (.RESET_B(net7516),
    .D(net1532),
    .Q(\u_inv.input_reg[133] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_1 _48394_ (.RESET_B(net7499),
    .D(net1686),
    .Q(\u_inv.input_reg[134] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_1 _48395_ (.RESET_B(net7499),
    .D(net2553),
    .Q(\u_inv.input_reg[135] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _48396_ (.RESET_B(net7511),
    .D(net2601),
    .Q(\u_inv.input_reg[136] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _48397_ (.RESET_B(net7509),
    .D(net2970),
    .Q(\u_inv.input_reg[137] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_1 _48398_ (.RESET_B(net7500),
    .D(net2230),
    .Q(\u_inv.input_reg[138] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _48399_ (.RESET_B(net7500),
    .D(net2474),
    .Q(\u_inv.input_reg[139] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_1 _48400_ (.RESET_B(net7500),
    .D(net1912),
    .Q(\u_inv.input_reg[140] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_1 _48401_ (.RESET_B(net7500),
    .D(net2263),
    .Q(\u_inv.input_reg[141] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_1 _48402_ (.RESET_B(net7500),
    .D(net1961),
    .Q(\u_inv.input_reg[142] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _48403_ (.RESET_B(net7500),
    .D(net1338),
    .Q(\u_inv.input_reg[143] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_1 _48404_ (.RESET_B(net7498),
    .D(net2363),
    .Q(\u_inv.input_reg[144] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_1 _48405_ (.RESET_B(net7499),
    .D(net2358),
    .Q(\u_inv.input_reg[145] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_1 _48406_ (.RESET_B(net7498),
    .D(net2792),
    .Q(\u_inv.input_reg[146] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_1 _48407_ (.RESET_B(net7498),
    .D(net2496),
    .Q(\u_inv.input_reg[147] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_1 _48408_ (.RESET_B(net7498),
    .D(net1886),
    .Q(\u_inv.input_reg[148] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_1 _48409_ (.RESET_B(net7498),
    .D(net2893),
    .Q(\u_inv.input_reg[149] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_1 _48410_ (.RESET_B(net7498),
    .D(net1805),
    .Q(\u_inv.input_reg[150] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_1 _48411_ (.RESET_B(net7501),
    .D(net2239),
    .Q(\u_inv.input_reg[151] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_1 _48412_ (.RESET_B(net7498),
    .D(net1499),
    .Q(\u_inv.input_reg[152] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_1 _48413_ (.RESET_B(net7496),
    .D(net1556),
    .Q(\u_inv.input_reg[153] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_1 _48414_ (.RESET_B(net7497),
    .D(net2042),
    .Q(\u_inv.input_reg[154] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_1 _48415_ (.RESET_B(net7495),
    .D(net2090),
    .Q(\u_inv.input_reg[155] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_1 _48416_ (.RESET_B(net7497),
    .D(net1414),
    .Q(\u_inv.input_reg[156] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_1 _48417_ (.RESET_B(net7497),
    .D(net2022),
    .Q(\u_inv.input_reg[157] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_1 _48418_ (.RESET_B(net7495),
    .D(net1503),
    .Q(\u_inv.input_reg[158] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_1 _48419_ (.RESET_B(net7495),
    .D(net2049),
    .Q(\u_inv.input_reg[159] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_1 _48420_ (.RESET_B(net7497),
    .D(net2478),
    .Q(\u_inv.input_reg[160] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_1 _48421_ (.RESET_B(net7489),
    .D(net1562),
    .Q(\u_inv.input_reg[161] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_1 _48422_ (.RESET_B(net7485),
    .D(net1455),
    .Q(\u_inv.input_reg[162] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _48423_ (.RESET_B(net7487),
    .D(_00070_),
    .Q(\u_inv.input_reg[163] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_1 _48424_ (.RESET_B(net7485),
    .D(net1981),
    .Q(\u_inv.input_reg[164] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _48425_ (.RESET_B(net7483),
    .D(net1884),
    .Q(\u_inv.input_reg[165] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_1 _48426_ (.RESET_B(net7479),
    .D(net1357),
    .Q(\u_inv.input_reg[166] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_1 _48427_ (.RESET_B(net7484),
    .D(net1517),
    .Q(\u_inv.input_reg[167] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _48428_ (.RESET_B(net7471),
    .D(net2354),
    .Q(\u_inv.input_reg[168] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_1 _48429_ (.RESET_B(net7471),
    .D(_00076_),
    .Q(\u_inv.input_reg[169] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _48430_ (.RESET_B(net7475),
    .D(net1931),
    .Q(\u_inv.input_reg[170] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _48431_ (.RESET_B(net7475),
    .D(net1520),
    .Q(\u_inv.input_reg[171] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _48432_ (.RESET_B(net7474),
    .D(net1330),
    .Q(\u_inv.input_reg[172] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _48433_ (.RESET_B(net7474),
    .D(net1288),
    .Q(\u_inv.input_reg[173] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _48434_ (.RESET_B(net7473),
    .D(net1631),
    .Q(\u_inv.input_reg[174] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _48435_ (.RESET_B(net7473),
    .D(net1979),
    .Q(\u_inv.input_reg[175] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _48436_ (.RESET_B(net7471),
    .D(net1552),
    .Q(\u_inv.input_reg[176] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _48437_ (.RESET_B(net7471),
    .D(net1571),
    .Q(\u_inv.input_reg[177] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _48438_ (.RESET_B(net7471),
    .D(net1405),
    .Q(\u_inv.input_reg[178] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _48439_ (.RESET_B(net7465),
    .D(net1582),
    .Q(\u_inv.input_reg[179] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _48440_ (.RESET_B(net7465),
    .D(net1545),
    .Q(\u_inv.input_reg[180] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_1 _48441_ (.RESET_B(net7465),
    .D(net1394),
    .Q(\u_inv.input_reg[181] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _48442_ (.RESET_B(net7469),
    .D(net1836),
    .Q(\u_inv.input_reg[182] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _48443_ (.RESET_B(net7471),
    .D(net2290),
    .Q(\u_inv.input_reg[183] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _48444_ (.RESET_B(net7464),
    .D(net1813),
    .Q(\u_inv.input_reg[184] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _48445_ (.RESET_B(net7464),
    .D(net1818),
    .Q(\u_inv.input_reg[185] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _48446_ (.RESET_B(net7464),
    .D(net2060),
    .Q(\u_inv.input_reg[186] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _48447_ (.RESET_B(net7464),
    .D(_00094_),
    .Q(\u_inv.input_reg[187] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_1 _48448_ (.RESET_B(net7458),
    .D(net1873),
    .Q(\u_inv.input_reg[188] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _48449_ (.RESET_B(net7464),
    .D(_00096_),
    .Q(\u_inv.input_reg[189] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _48450_ (.RESET_B(net7458),
    .D(net2000),
    .Q(\u_inv.input_reg[190] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _48451_ (.RESET_B(net7458),
    .D(net1463),
    .Q(\u_inv.input_reg[191] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _48452_ (.RESET_B(net7456),
    .D(net1283),
    .Q(\u_inv.input_reg[192] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _48453_ (.RESET_B(net7419),
    .D(net1807),
    .Q(\u_inv.input_reg[193] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _48454_ (.RESET_B(net7420),
    .D(net1714),
    .Q(\u_inv.input_reg[194] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _48455_ (.RESET_B(net7418),
    .D(net1784),
    .Q(\u_inv.input_reg[195] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _48456_ (.RESET_B(net7419),
    .D(net1705),
    .Q(\u_inv.input_reg[196] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _48457_ (.RESET_B(net7419),
    .D(net1834),
    .Q(\u_inv.input_reg[197] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _48458_ (.RESET_B(net7418),
    .D(net1457),
    .Q(\u_inv.input_reg[198] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _48459_ (.RESET_B(net7420),
    .D(net1426),
    .Q(\u_inv.input_reg[199] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _48460_ (.RESET_B(net7417),
    .D(net1341),
    .Q(\u_inv.input_reg[200] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _48461_ (.RESET_B(net7456),
    .D(_00108_),
    .Q(\u_inv.input_reg[201] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _48462_ (.RESET_B(net7417),
    .D(net1661),
    .Q(\u_inv.input_reg[202] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _48463_ (.RESET_B(net7457),
    .D(_00110_),
    .Q(\u_inv.input_reg[203] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _48464_ (.RESET_B(net7420),
    .D(net2485),
    .Q(\u_inv.input_reg[204] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _48465_ (.RESET_B(net7418),
    .D(net2261),
    .Q(\u_inv.input_reg[205] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _48466_ (.RESET_B(net7416),
    .D(net1929),
    .Q(\u_inv.input_reg[206] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _48467_ (.RESET_B(net7419),
    .D(net2719),
    .Q(\u_inv.input_reg[207] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _48468_ (.RESET_B(net7417),
    .D(net1482),
    .Q(\u_inv.input_reg[208] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _48469_ (.RESET_B(net7418),
    .D(net2302),
    .Q(\u_inv.input_reg[209] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _48470_ (.RESET_B(net7417),
    .D(net1529),
    .Q(\u_inv.input_reg[210] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _48471_ (.RESET_B(net7417),
    .D(net1218),
    .Q(\u_inv.input_reg[211] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _48472_ (.RESET_B(net7417),
    .D(net1700),
    .Q(\u_inv.input_reg[212] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _48473_ (.RESET_B(net7418),
    .D(net2458),
    .Q(\u_inv.input_reg[213] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _48474_ (.RESET_B(net7417),
    .D(net2273),
    .Q(\u_inv.input_reg[214] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _48475_ (.RESET_B(net7415),
    .D(net1629),
    .Q(\u_inv.input_reg[215] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _48476_ (.RESET_B(net7421),
    .D(net1626),
    .Q(\u_inv.input_reg[216] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _48477_ (.RESET_B(net7421),
    .D(net1311),
    .Q(\u_inv.input_reg[217] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _48478_ (.RESET_B(net7424),
    .D(net1470),
    .Q(\u_inv.input_reg[218] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _48479_ (.RESET_B(net7421),
    .D(net2524),
    .Q(\u_inv.input_reg[219] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _48480_ (.RESET_B(net7415),
    .D(net1313),
    .Q(\u_inv.input_reg[220] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _48481_ (.RESET_B(net7415),
    .D(net1869),
    .Q(\u_inv.input_reg[221] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _48482_ (.RESET_B(net7421),
    .D(net1796),
    .Q(\u_inv.input_reg[222] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _48483_ (.RESET_B(net7415),
    .D(_00130_),
    .Q(\u_inv.input_reg[223] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _48484_ (.RESET_B(net7415),
    .D(net1400),
    .Q(\u_inv.input_reg[224] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _48485_ (.RESET_B(net7415),
    .D(net1839),
    .Q(\u_inv.input_reg[225] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _48486_ (.RESET_B(net7414),
    .D(net1396),
    .Q(\u_inv.input_reg[226] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _48487_ (.RESET_B(net7416),
    .D(net1653),
    .Q(\u_inv.input_reg[227] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _48488_ (.RESET_B(net7414),
    .D(net1560),
    .Q(\u_inv.input_reg[228] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _48489_ (.RESET_B(net7414),
    .D(net1611),
    .Q(\u_inv.input_reg[229] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _48490_ (.RESET_B(net7416),
    .D(net1402),
    .Q(\u_inv.input_reg[230] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _48491_ (.RESET_B(net7414),
    .D(net2094),
    .Q(\u_inv.input_reg[231] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _48492_ (.RESET_B(net7430),
    .D(net1386),
    .Q(\u_inv.input_reg[232] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _48493_ (.RESET_B(net7415),
    .D(net1378),
    .Q(\u_inv.input_reg[233] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _48494_ (.RESET_B(net7430),
    .D(net1515),
    .Q(\u_inv.input_reg[234] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _48495_ (.RESET_B(net7430),
    .D(net1943),
    .Q(\u_inv.input_reg[235] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _48496_ (.RESET_B(net7430),
    .D(net1439),
    .Q(\u_inv.input_reg[236] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _48497_ (.RESET_B(net7430),
    .D(net1290),
    .Q(\u_inv.input_reg[237] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _48498_ (.RESET_B(net7430),
    .D(net1605),
    .Q(\u_inv.input_reg[238] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _48499_ (.RESET_B(net7430),
    .D(net1334),
    .Q(\u_inv.input_reg[239] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _48500_ (.RESET_B(net7434),
    .D(net1328),
    .Q(\u_inv.input_reg[240] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _48501_ (.RESET_B(net7434),
    .D(net1321),
    .Q(\u_inv.input_reg[241] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _48502_ (.RESET_B(net7432),
    .D(net1476),
    .Q(\u_inv.input_reg[242] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _48503_ (.RESET_B(net7434),
    .D(net1428),
    .Q(\u_inv.input_reg[243] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _48504_ (.RESET_B(net7432),
    .D(net1707),
    .Q(\u_inv.input_reg[244] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _48505_ (.RESET_B(net7448),
    .D(net1565),
    .Q(\u_inv.input_reg[245] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _48506_ (.RESET_B(net7432),
    .D(net1368),
    .Q(\u_inv.input_reg[246] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _48507_ (.RESET_B(net7448),
    .D(net1309),
    .Q(\u_inv.input_reg[247] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _48508_ (.RESET_B(net7437),
    .D(net1716),
    .Q(\u_inv.input_reg[248] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _48509_ (.RESET_B(net7437),
    .D(net1990),
    .Q(\u_inv.input_reg[249] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _48510_ (.RESET_B(net7437),
    .D(net2324),
    .Q(\u_inv.input_reg[250] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _48511_ (.RESET_B(net7435),
    .D(net1964),
    .Q(\u_inv.input_reg[251] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _48512_ (.RESET_B(net7439),
    .D(net2506),
    .Q(\u_inv.input_reg[252] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _48513_ (.RESET_B(net7439),
    .D(net1315),
    .Q(\u_inv.input_reg[253] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _48514_ (.RESET_B(net7439),
    .D(net1776),
    .Q(\u_inv.input_reg[254] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _48515_ (.RESET_B(net7439),
    .D(net1803),
    .Q(\u_inv.input_reg[255] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _48516_ (.RESET_B(net7453),
    .D(net1160),
    .Q(parity_error),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _48517_ (.RESET_B(net7435),
    .D(_00164_),
    .Q(\u_trng.bit_cnt[0] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _48518_ (.RESET_B(net7435),
    .D(_00165_),
    .Q(\u_trng.bit_cnt[1] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _48519_ (.RESET_B(net7435),
    .D(net1152),
    .Q(\u_trng.bit_cnt[2] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _48520_ (.RESET_B(net7450),
    .D(net3748),
    .Q(\state[0] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _48521_ (.RESET_B(net7450),
    .D(_00168_),
    .Q(\state[1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _48522_ (.RESET_B(net7451),
    .D(_00169_),
    .Q(\byte_cnt[0] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _48523_ (.RESET_B(net7451),
    .D(net1168),
    .Q(\byte_cnt[1] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _48524_ (.RESET_B(net7451),
    .D(_00171_),
    .Q(\byte_cnt[2] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _48525_ (.RESET_B(net7451),
    .D(net1154),
    .Q(\byte_cnt[3] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _48526_ (.RESET_B(net7451),
    .D(_00173_),
    .Q(\byte_cnt[4] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _48527_ (.RESET_B(net7450),
    .D(net2487),
    .Q(\byte_cnt[5] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _48528_ (.RESET_B(net7451),
    .D(net2612),
    .Q(inv_go),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _48529_ (.RESET_B(net7453),
    .D(net1731),
    .Q(\shift_reg[0] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _48530_ (.RESET_B(net7470),
    .D(net1970),
    .Q(\shift_reg[1] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _48531_ (.RESET_B(net7453),
    .D(net1522),
    .Q(\shift_reg[2] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _48532_ (.RESET_B(net7453),
    .D(net1575),
    .Q(\shift_reg[3] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _48533_ (.RESET_B(net7454),
    .D(net3403),
    .Q(\shift_reg[4] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _48534_ (.RESET_B(net7454),
    .D(net3672),
    .Q(\shift_reg[5] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _48535_ (.RESET_B(net7453),
    .D(net3451),
    .Q(\shift_reg[6] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _48536_ (.RESET_B(net7494),
    .D(_00182_),
    .Q(\shift_reg[7] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _48537_ (.RESET_B(net7459),
    .D(net1495),
    .Q(\shift_reg[8] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _48538_ (.RESET_B(net7468),
    .D(net1325),
    .Q(\shift_reg[9] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _48539_ (.RESET_B(net7458),
    .D(_00185_),
    .Q(\shift_reg[10] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _48540_ (.RESET_B(net7462),
    .D(_00186_),
    .Q(\shift_reg[11] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _48541_ (.RESET_B(net7457),
    .D(net2467),
    .Q(\shift_reg[12] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _48542_ (.RESET_B(net7469),
    .D(net1200),
    .Q(\shift_reg[13] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _48543_ (.RESET_B(net7459),
    .D(net2829),
    .Q(\shift_reg[14] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _48544_ (.RESET_B(net7481),
    .D(_00190_),
    .Q(\shift_reg[15] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _48545_ (.RESET_B(net7456),
    .D(_00191_),
    .Q(\shift_reg[16] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _48546_ (.RESET_B(net7463),
    .D(_00192_),
    .Q(\shift_reg[17] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _48547_ (.RESET_B(net7471),
    .D(_00193_),
    .Q(\shift_reg[18] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _48548_ (.RESET_B(net7463),
    .D(_00194_),
    .Q(\shift_reg[19] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _48549_ (.RESET_B(net7463),
    .D(_00195_),
    .Q(\shift_reg[20] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _48550_ (.RESET_B(net7463),
    .D(_00196_),
    .Q(\shift_reg[21] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _48551_ (.RESET_B(net7463),
    .D(_00197_),
    .Q(\shift_reg[22] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _48552_ (.RESET_B(net7479),
    .D(net2779),
    .Q(\shift_reg[23] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _48553_ (.RESET_B(net7482),
    .D(net3527),
    .Q(\shift_reg[24] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _48554_ (.RESET_B(net7478),
    .D(_00200_),
    .Q(\shift_reg[25] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _48555_ (.RESET_B(net7484),
    .D(net3337),
    .Q(\shift_reg[26] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_2 _48556_ (.RESET_B(net7485),
    .D(net3400),
    .Q(\shift_reg[27] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_2 _48557_ (.RESET_B(net7478),
    .D(_00203_),
    .Q(\shift_reg[28] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _48558_ (.RESET_B(net7483),
    .D(net3247),
    .Q(\shift_reg[29] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _48559_ (.RESET_B(net7482),
    .D(net3207),
    .Q(\shift_reg[30] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _48560_ (.RESET_B(net7483),
    .D(_00206_),
    .Q(\shift_reg[31] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_2 _48561_ (.RESET_B(net7488),
    .D(net2597),
    .Q(\shift_reg[32] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _48562_ (.RESET_B(net7489),
    .D(net2803),
    .Q(\shift_reg[33] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _48563_ (.RESET_B(net7485),
    .D(net3192),
    .Q(\shift_reg[34] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_2 _48564_ (.RESET_B(net7485),
    .D(net3279),
    .Q(\shift_reg[35] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_2 _48565_ (.RESET_B(net7490),
    .D(net2931),
    .Q(\shift_reg[36] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _48566_ (.RESET_B(net7490),
    .D(net3016),
    .Q(\shift_reg[37] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _48567_ (.RESET_B(net7488),
    .D(_00213_),
    .Q(\shift_reg[38] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _48568_ (.RESET_B(net7496),
    .D(net2252),
    .Q(\shift_reg[39] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _48569_ (.RESET_B(net7488),
    .D(_00215_),
    .Q(\shift_reg[40] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _48570_ (.RESET_B(net7490),
    .D(_00216_),
    .Q(\shift_reg[41] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _48571_ (.RESET_B(net7495),
    .D(_00217_),
    .Q(\shift_reg[42] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _48572_ (.RESET_B(net7496),
    .D(_00218_),
    .Q(\shift_reg[43] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _48573_ (.RESET_B(net7513),
    .D(net2782),
    .Q(\shift_reg[44] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _48574_ (.RESET_B(net7514),
    .D(net1765),
    .Q(\shift_reg[45] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _48575_ (.RESET_B(net7498),
    .D(_00221_),
    .Q(\shift_reg[46] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _48576_ (.RESET_B(net7512),
    .D(_00222_),
    .Q(\shift_reg[47] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _48577_ (.RESET_B(net7512),
    .D(net2823),
    .Q(\shift_reg[48] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_2 _48578_ (.RESET_B(net7512),
    .D(net3101),
    .Q(\shift_reg[49] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _48579_ (.RESET_B(net7513),
    .D(net2734),
    .Q(\shift_reg[50] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _48580_ (.RESET_B(net7513),
    .D(net2954),
    .Q(\shift_reg[51] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_2 _48581_ (.RESET_B(net7513),
    .D(_00227_),
    .Q(\shift_reg[52] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_2 _48582_ (.RESET_B(net7519),
    .D(_00228_),
    .Q(\shift_reg[53] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_2 _48583_ (.RESET_B(net7513),
    .D(net3468),
    .Q(\shift_reg[54] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _48584_ (.RESET_B(net7513),
    .D(net3041),
    .Q(\shift_reg[55] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _48585_ (.RESET_B(net7517),
    .D(_00231_),
    .Q(\shift_reg[56] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_2 _48586_ (.RESET_B(net7517),
    .D(net2771),
    .Q(\shift_reg[57] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _48587_ (.RESET_B(net7517),
    .D(_00233_),
    .Q(\shift_reg[58] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_2 _48588_ (.RESET_B(net7517),
    .D(_00234_),
    .Q(\shift_reg[59] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _48589_ (.RESET_B(net7518),
    .D(_00235_),
    .Q(\shift_reg[60] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_2 _48590_ (.RESET_B(net7518),
    .D(_00236_),
    .Q(\shift_reg[61] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_2 _48591_ (.RESET_B(net7518),
    .D(net3453),
    .Q(\shift_reg[62] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_2 _48592_ (.RESET_B(net7519),
    .D(_00238_),
    .Q(\shift_reg[63] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_2 _48593_ (.RESET_B(net7519),
    .D(_00239_),
    .Q(\shift_reg[64] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_2 _48594_ (.RESET_B(net7528),
    .D(net2901),
    .Q(\shift_reg[65] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _48595_ (.RESET_B(net7526),
    .D(_00241_),
    .Q(\shift_reg[66] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _48596_ (.RESET_B(net7526),
    .D(net3140),
    .Q(\shift_reg[67] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_2 _48597_ (.RESET_B(net7526),
    .D(net3269),
    .Q(\shift_reg[68] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _48598_ (.RESET_B(net7528),
    .D(net2622),
    .Q(\shift_reg[69] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _48599_ (.RESET_B(net7528),
    .D(net3431),
    .Q(\shift_reg[70] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _48600_ (.RESET_B(net7527),
    .D(net3219),
    .Q(\shift_reg[71] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _48601_ (.RESET_B(net7531),
    .D(_00247_),
    .Q(\shift_reg[72] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_2 _48602_ (.RESET_B(net7531),
    .D(_00248_),
    .Q(\shift_reg[73] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _48603_ (.RESET_B(net7527),
    .D(_00249_),
    .Q(\shift_reg[74] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_2 _48604_ (.RESET_B(net7531),
    .D(_00250_),
    .Q(\shift_reg[75] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _48605_ (.RESET_B(net7527),
    .D(_00251_),
    .Q(\shift_reg[76] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _48606_ (.RESET_B(net7527),
    .D(net3444),
    .Q(\shift_reg[77] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _48607_ (.RESET_B(net7527),
    .D(net3428),
    .Q(\shift_reg[78] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _48608_ (.RESET_B(net7531),
    .D(_00254_),
    .Q(\shift_reg[79] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _48609_ (.RESET_B(net7550),
    .D(net2702),
    .Q(\shift_reg[80] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_2 _48610_ (.RESET_B(net7550),
    .D(net2995),
    .Q(\shift_reg[81] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_2 _48611_ (.RESET_B(net7550),
    .D(net2817),
    .Q(\shift_reg[82] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_2 _48612_ (.RESET_B(net7551),
    .D(net2435),
    .Q(\shift_reg[83] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_2 _48613_ (.RESET_B(net7550),
    .D(net2913),
    .Q(\shift_reg[84] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_2 _48614_ (.RESET_B(net7533),
    .D(net3127),
    .Q(\shift_reg[85] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_2 _48615_ (.RESET_B(net7551),
    .D(net3089),
    .Q(\shift_reg[86] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_2 _48616_ (.RESET_B(net7551),
    .D(net3169),
    .Q(\shift_reg[87] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_2 _48617_ (.RESET_B(net7559),
    .D(net2411),
    .Q(\shift_reg[88] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_2 _48618_ (.RESET_B(net7559),
    .D(_00264_),
    .Q(\shift_reg[89] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_2 _48619_ (.RESET_B(net7558),
    .D(_00265_),
    .Q(\shift_reg[90] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_2 _48620_ (.RESET_B(net7558),
    .D(_00266_),
    .Q(\shift_reg[91] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_2 _48621_ (.RESET_B(net7558),
    .D(_00267_),
    .Q(\shift_reg[92] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_2 _48622_ (.RESET_B(net7551),
    .D(net3087),
    .Q(\shift_reg[93] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_2 _48623_ (.RESET_B(net7564),
    .D(_00269_),
    .Q(\shift_reg[94] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_2 _48624_ (.RESET_B(net7558),
    .D(net3049),
    .Q(\shift_reg[95] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_2 _48625_ (.RESET_B(net7558),
    .D(_00271_),
    .Q(\shift_reg[96] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_2 _48626_ (.RESET_B(net7558),
    .D(_00272_),
    .Q(\shift_reg[97] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_2 _48627_ (.RESET_B(net7555),
    .D(net3123),
    .Q(\shift_reg[98] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_2 _48628_ (.RESET_B(net7556),
    .D(net2572),
    .Q(\shift_reg[99] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_2 _48629_ (.RESET_B(net7563),
    .D(net2854),
    .Q(\shift_reg[100] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_2 _48630_ (.RESET_B(net7555),
    .D(net2935),
    .Q(\shift_reg[101] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_2 _48631_ (.RESET_B(net7553),
    .D(net3194),
    .Q(\shift_reg[102] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_2 _48632_ (.RESET_B(net7563),
    .D(_00278_),
    .Q(\shift_reg[103] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_2 _48633_ (.RESET_B(net7555),
    .D(_00279_),
    .Q(\shift_reg[104] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_2 _48634_ (.RESET_B(net7555),
    .D(_00280_),
    .Q(\shift_reg[105] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_2 _48635_ (.RESET_B(net7554),
    .D(_00281_),
    .Q(\shift_reg[106] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_2 _48636_ (.RESET_B(net7565),
    .D(_00282_),
    .Q(\shift_reg[107] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_2 _48637_ (.RESET_B(net7554),
    .D(_00283_),
    .Q(\shift_reg[108] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_2 _48638_ (.RESET_B(net7556),
    .D(_00284_),
    .Q(\shift_reg[109] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_2 _48639_ (.RESET_B(net7553),
    .D(_00285_),
    .Q(\shift_reg[110] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_2 _48640_ (.RESET_B(net7556),
    .D(_00286_),
    .Q(\shift_reg[111] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_2 _48641_ (.RESET_B(net7534),
    .D(net2555),
    .Q(\shift_reg[112] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _48642_ (.RESET_B(net7534),
    .D(net2652),
    .Q(\shift_reg[113] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_2 _48643_ (.RESET_B(net7535),
    .D(net2915),
    .Q(\shift_reg[114] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_2 _48644_ (.RESET_B(net7536),
    .D(net3148),
    .Q(\shift_reg[115] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_2 _48645_ (.RESET_B(net7536),
    .D(net3184),
    .Q(\shift_reg[116] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_2 _48646_ (.RESET_B(net7534),
    .D(net2116),
    .Q(\shift_reg[117] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_2 _48647_ (.RESET_B(net7536),
    .D(net2924),
    .Q(\shift_reg[118] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_2 _48648_ (.RESET_B(net7548),
    .D(_00294_),
    .Q(\shift_reg[119] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_2 _48649_ (.RESET_B(net7546),
    .D(net2335),
    .Q(\shift_reg[120] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _48650_ (.RESET_B(net7546),
    .D(net2424),
    .Q(\shift_reg[121] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _48651_ (.RESET_B(net7545),
    .D(net2452),
    .Q(\shift_reg[122] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _48652_ (.RESET_B(net7545),
    .D(net1977),
    .Q(\shift_reg[123] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_2 _48653_ (.RESET_B(net7545),
    .D(net2348),
    .Q(\shift_reg[124] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _48654_ (.RESET_B(net7540),
    .D(_00300_),
    .Q(\shift_reg[125] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_2 _48655_ (.RESET_B(net7540),
    .D(_00301_),
    .Q(\shift_reg[126] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_2 _48656_ (.RESET_B(net7540),
    .D(net1937),
    .Q(\shift_reg[127] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_2 _48657_ (.RESET_B(net7538),
    .D(net2020),
    .Q(\shift_reg[128] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _48658_ (.RESET_B(net7539),
    .D(_00304_),
    .Q(\shift_reg[129] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _48659_ (.RESET_B(net7539),
    .D(_00305_),
    .Q(\shift_reg[130] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _48660_ (.RESET_B(net7539),
    .D(_00306_),
    .Q(\shift_reg[131] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _48661_ (.RESET_B(net7539),
    .D(_00307_),
    .Q(\shift_reg[132] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _48662_ (.RESET_B(net7523),
    .D(net2577),
    .Q(\shift_reg[133] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _48663_ (.RESET_B(net7538),
    .D(net2429),
    .Q(\shift_reg[134] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_2 _48664_ (.RESET_B(net7538),
    .D(_00310_),
    .Q(\shift_reg[135] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_2 _48665_ (.RESET_B(net7542),
    .D(net1975),
    .Q(\shift_reg[136] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _48666_ (.RESET_B(net7542),
    .D(net2292),
    .Q(\shift_reg[137] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_2 _48667_ (.RESET_B(net7541),
    .D(_00313_),
    .Q(\shift_reg[138] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_2 _48668_ (.RESET_B(net7541),
    .D(_00314_),
    .Q(\shift_reg[139] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _48669_ (.RESET_B(net7542),
    .D(_00315_),
    .Q(\shift_reg[140] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _48670_ (.RESET_B(net7523),
    .D(_00316_),
    .Q(\shift_reg[141] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _48671_ (.RESET_B(net7541),
    .D(_00317_),
    .Q(\shift_reg[142] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_2 _48672_ (.RESET_B(net7541),
    .D(_00318_),
    .Q(\shift_reg[143] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_2 _48673_ (.RESET_B(net7523),
    .D(_00319_),
    .Q(\shift_reg[144] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _48674_ (.RESET_B(net7523),
    .D(_00320_),
    .Q(\shift_reg[145] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _48675_ (.RESET_B(net7522),
    .D(_00321_),
    .Q(\shift_reg[146] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _48676_ (.RESET_B(net7524),
    .D(_00322_),
    .Q(\shift_reg[147] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _48677_ (.RESET_B(net7522),
    .D(_00323_),
    .Q(\shift_reg[148] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _48678_ (.RESET_B(net7521),
    .D(_00324_),
    .Q(\shift_reg[149] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _48679_ (.RESET_B(net7510),
    .D(_00325_),
    .Q(\shift_reg[150] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _48680_ (.RESET_B(net7521),
    .D(_00326_),
    .Q(\shift_reg[151] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _48681_ (.RESET_B(net7521),
    .D(net3257),
    .Q(\shift_reg[152] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _48682_ (.RESET_B(net7508),
    .D(net3099),
    .Q(\shift_reg[153] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _48683_ (.RESET_B(net7510),
    .D(net3333),
    .Q(\shift_reg[154] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _48684_ (.RESET_B(net7508),
    .D(net2751),
    .Q(\shift_reg[155] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _48685_ (.RESET_B(net7507),
    .D(net3382),
    .Q(\shift_reg[156] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _48686_ (.RESET_B(net7510),
    .D(net2899),
    .Q(\shift_reg[157] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _48687_ (.RESET_B(net7507),
    .D(net3302),
    .Q(\shift_reg[158] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _48688_ (.RESET_B(net7507),
    .D(net3330),
    .Q(\shift_reg[159] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _48689_ (.RESET_B(net7508),
    .D(_00335_),
    .Q(\shift_reg[160] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _48690_ (.RESET_B(net7509),
    .D(_00336_),
    .Q(\shift_reg[161] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_2 _48691_ (.RESET_B(net7509),
    .D(net3249),
    .Q(\shift_reg[162] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _48692_ (.RESET_B(net7509),
    .D(_00338_),
    .Q(\shift_reg[163] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_2 _48693_ (.RESET_B(net7507),
    .D(net3108),
    .Q(\shift_reg[164] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_2 _48694_ (.RESET_B(net7507),
    .D(_00340_),
    .Q(\shift_reg[165] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_2 _48695_ (.RESET_B(net7505),
    .D(_00341_),
    .Q(\shift_reg[166] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _48696_ (.RESET_B(net7505),
    .D(net3243),
    .Q(\shift_reg[167] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _48697_ (.RESET_B(net7507),
    .D(_00343_),
    .Q(\shift_reg[168] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _48698_ (.RESET_B(net7507),
    .D(_00344_),
    .Q(\shift_reg[169] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_2 _48699_ (.RESET_B(net7504),
    .D(_00345_),
    .Q(\shift_reg[170] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _48700_ (.RESET_B(net7505),
    .D(net3352),
    .Q(\shift_reg[171] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_2 _48701_ (.RESET_B(net7505),
    .D(_00347_),
    .Q(\shift_reg[172] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_2 _48702_ (.RESET_B(net7503),
    .D(_00348_),
    .Q(\shift_reg[173] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _48703_ (.RESET_B(net7502),
    .D(_00349_),
    .Q(\shift_reg[174] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _48704_ (.RESET_B(net7502),
    .D(_00350_),
    .Q(\shift_reg[175] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _48705_ (.RESET_B(net7503),
    .D(net3522),
    .Q(\shift_reg[176] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _48706_ (.RESET_B(net7502),
    .D(net3282),
    .Q(\shift_reg[177] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_2 _48707_ (.RESET_B(net7493),
    .D(_00353_),
    .Q(\shift_reg[178] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _48708_ (.RESET_B(net7493),
    .D(net2794),
    .Q(\shift_reg[179] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _48709_ (.RESET_B(net7493),
    .D(net3311),
    .Q(\shift_reg[180] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _48710_ (.RESET_B(net7502),
    .D(net3499),
    .Q(\shift_reg[181] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _48711_ (.RESET_B(net7494),
    .D(net3224),
    .Q(\shift_reg[182] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _48712_ (.RESET_B(net7491),
    .D(net3178),
    .Q(\shift_reg[183] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _48713_ (.RESET_B(net7474),
    .D(_00359_),
    .Q(\shift_reg[184] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _48714_ (.RESET_B(net7474),
    .D(_00360_),
    .Q(\shift_reg[185] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _48715_ (.RESET_B(net7475),
    .D(net2679),
    .Q(\shift_reg[186] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _48716_ (.RESET_B(net7475),
    .D(net2294),
    .Q(\shift_reg[187] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_2 _48717_ (.RESET_B(net7486),
    .D(_00363_),
    .Q(\shift_reg[188] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _48718_ (.RESET_B(net7486),
    .D(_00364_),
    .Q(\shift_reg[189] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _48719_ (.RESET_B(net7474),
    .D(net2234),
    .Q(\shift_reg[190] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _48720_ (.RESET_B(net7481),
    .D(_00366_),
    .Q(\shift_reg[191] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _48721_ (.RESET_B(net7474),
    .D(_00367_),
    .Q(\shift_reg[192] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _48722_ (.RESET_B(net7473),
    .D(net2212),
    .Q(\shift_reg[193] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _48723_ (.RESET_B(net7473),
    .D(net2322),
    .Q(\shift_reg[194] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _48724_ (.RESET_B(net7473),
    .D(net2352),
    .Q(\shift_reg[195] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _48725_ (.RESET_B(net7473),
    .D(net2605),
    .Q(\shift_reg[196] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _48726_ (.RESET_B(net7473),
    .D(net2536),
    .Q(\shift_reg[197] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _48727_ (.RESET_B(net7472),
    .D(_00373_),
    .Q(\shift_reg[198] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _48728_ (.RESET_B(net7472),
    .D(net2557),
    .Q(\shift_reg[199] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _48729_ (.RESET_B(net7472),
    .D(_00375_),
    .Q(\shift_reg[200] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _48730_ (.RESET_B(net7472),
    .D(_00376_),
    .Q(\shift_reg[201] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _48731_ (.RESET_B(net7472),
    .D(_00377_),
    .Q(\shift_reg[202] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _48732_ (.RESET_B(net7466),
    .D(net2278),
    .Q(\shift_reg[203] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _48733_ (.RESET_B(net7466),
    .D(_00379_),
    .Q(\shift_reg[204] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _48734_ (.RESET_B(net7466),
    .D(net2249),
    .Q(\shift_reg[205] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _48735_ (.RESET_B(net7465),
    .D(net2508),
    .Q(\shift_reg[206] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _48736_ (.RESET_B(net7465),
    .D(_00382_),
    .Q(\shift_reg[207] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _48737_ (.RESET_B(net7464),
    .D(_00383_),
    .Q(\shift_reg[208] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _48738_ (.RESET_B(net7458),
    .D(net2547),
    .Q(\shift_reg[209] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _48739_ (.RESET_B(net7464),
    .D(_00385_),
    .Q(\shift_reg[210] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _48740_ (.RESET_B(net7461),
    .D(_00386_),
    .Q(\shift_reg[211] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _48741_ (.RESET_B(net7461),
    .D(net3003),
    .Q(\shift_reg[212] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _48742_ (.RESET_B(net7468),
    .D(_00388_),
    .Q(\shift_reg[213] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _48743_ (.RESET_B(net7456),
    .D(_00389_),
    .Q(\shift_reg[214] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _48744_ (.RESET_B(net7461),
    .D(_00390_),
    .Q(\shift_reg[215] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _48745_ (.RESET_B(net7461),
    .D(_00391_),
    .Q(\shift_reg[216] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _48746_ (.RESET_B(net7456),
    .D(net2172),
    .Q(\shift_reg[217] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _48747_ (.RESET_B(net7458),
    .D(_00393_),
    .Q(\shift_reg[218] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _48748_ (.RESET_B(net7456),
    .D(net2729),
    .Q(\shift_reg[219] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _48749_ (.RESET_B(net7461),
    .D(net2962),
    .Q(\shift_reg[220] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _48750_ (.RESET_B(net7461),
    .D(net3235),
    .Q(\shift_reg[221] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _48751_ (.RESET_B(net7456),
    .D(_00397_),
    .Q(\shift_reg[222] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _48752_ (.RESET_B(net7461),
    .D(_00398_),
    .Q(\shift_reg[223] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _48753_ (.RESET_B(net7460),
    .D(net3433),
    .Q(\shift_reg[224] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _48754_ (.RESET_B(net7457),
    .D(_00400_),
    .Q(\shift_reg[225] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _48755_ (.RESET_B(net7459),
    .D(net3229),
    .Q(\shift_reg[226] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _48756_ (.RESET_B(net7459),
    .D(_00402_),
    .Q(\shift_reg[227] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _48757_ (.RESET_B(net7459),
    .D(_00403_),
    .Q(\shift_reg[228] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _48758_ (.RESET_B(net7460),
    .D(_00404_),
    .Q(\shift_reg[229] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _48759_ (.RESET_B(net7417),
    .D(net2632),
    .Q(\shift_reg[230] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _48760_ (.RESET_B(net7426),
    .D(net3319),
    .Q(\shift_reg[231] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _48761_ (.RESET_B(net7421),
    .D(net2520),
    .Q(\shift_reg[232] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _48762_ (.RESET_B(net7421),
    .D(net2175),
    .Q(\shift_reg[233] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _48763_ (.RESET_B(net7426),
    .D(net2743),
    .Q(\shift_reg[234] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _48764_ (.RESET_B(net7426),
    .D(net2801),
    .Q(\shift_reg[235] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _48765_ (.RESET_B(net7421),
    .D(net2247),
    .Q(\shift_reg[236] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _48766_ (.RESET_B(net7427),
    .D(net3263),
    .Q(\shift_reg[237] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _48767_ (.RESET_B(net7421),
    .D(net2331),
    .Q(\shift_reg[238] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _48768_ (.RESET_B(net7422),
    .D(net1852),
    .Q(\shift_reg[239] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _48769_ (.RESET_B(net7414),
    .D(_00415_),
    .Q(\shift_reg[240] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _48770_ (.RESET_B(net7422),
    .D(net2550),
    .Q(\shift_reg[241] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _48771_ (.RESET_B(net7422),
    .D(net3063),
    .Q(\shift_reg[242] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _48772_ (.RESET_B(net7422),
    .D(net2404),
    .Q(\shift_reg[243] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _48773_ (.RESET_B(net7414),
    .D(net2139),
    .Q(\shift_reg[244] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _48774_ (.RESET_B(net7422),
    .D(net2609),
    .Q(\shift_reg[245] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _48775_ (.RESET_B(net7414),
    .D(net2392),
    .Q(\shift_reg[246] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _48776_ (.RESET_B(net7414),
    .D(net2271),
    .Q(\shift_reg[247] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _48777_ (.RESET_B(net7431),
    .D(_00423_),
    .Q(\shift_reg[248] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _48778_ (.RESET_B(net7441),
    .D(_00424_),
    .Q(\shift_reg[249] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _48779_ (.RESET_B(net7431),
    .D(net2565),
    .Q(\shift_reg[250] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _48780_ (.RESET_B(net7441),
    .D(net3021),
    .Q(\shift_reg[251] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _48781_ (.RESET_B(net7430),
    .D(net2510),
    .Q(\shift_reg[252] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _48782_ (.RESET_B(net7441),
    .D(_00428_),
    .Q(\shift_reg[253] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _48783_ (.RESET_B(net7431),
    .D(_00429_),
    .Q(\shift_reg[254] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _48784_ (.RESET_B(net7431),
    .D(_00430_),
    .Q(\shift_reg[255] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _48785_ (.RESET_B(net7432),
    .D(net2650),
    .Q(\shift_reg[256] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _48786_ (.RESET_B(net7432),
    .D(net2209),
    .Q(\shift_reg[257] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _48787_ (.RESET_B(net7432),
    .D(net2157),
    .Q(\shift_reg[258] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _48788_ (.RESET_B(net7432),
    .D(net2159),
    .Q(\shift_reg[259] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _48789_ (.RESET_B(net7433),
    .D(_00435_),
    .Q(\shift_reg[260] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _48790_ (.RESET_B(net7444),
    .D(net2983),
    .Q(\shift_reg[261] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _48791_ (.RESET_B(net7433),
    .D(net2110),
    .Q(\shift_reg[262] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _48792_ (.RESET_B(net7433),
    .D(net2288),
    .Q(\shift_reg[263] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _48793_ (.RESET_B(net7448),
    .D(net2627),
    .Q(\shift_reg[264] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _48794_ (.RESET_B(net7438),
    .D(_00440_),
    .Q(\shift_reg[265] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _48795_ (.RESET_B(net7437),
    .D(_00441_),
    .Q(\shift_reg[266] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _48796_ (.RESET_B(net7450),
    .D(net2861),
    .Q(\shift_reg[267] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _48797_ (.RESET_B(net7439),
    .D(net2575),
    .Q(\shift_reg[268] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _48798_ (.RESET_B(net7450),
    .D(net2929),
    .Q(\shift_reg[269] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _48799_ (.RESET_B(net7439),
    .D(_00445_),
    .Q(\shift_reg[270] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _48800_ (.RESET_B(net7439),
    .D(net2431),
    .Q(\shift_reg[271] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _48801_ (.RESET_B(net7450),
    .D(net1181),
    .Q(next_loaded),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _48802_ (.RESET_B(net7438),
    .D(_00448_),
    .Q(pipe_pending),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _48803_ (.RESET_B(net7450),
    .D(net10),
    .Q(wr_prev),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _48804_ (.RESET_B(net7438),
    .D(net11),
    .Q(rd_prev),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _48805_ (.RESET_B(net7438),
    .D(net2852),
    .Q(\trng_data[0] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _48806_ (.RESET_B(net7435),
    .D(net2280),
    .Q(\trng_data[1] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _48807_ (.RESET_B(net7436),
    .D(net2265),
    .Q(\trng_data[2] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _48808_ (.RESET_B(net7436),
    .D(net2063),
    .Q(\trng_data[3] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _48809_ (.RESET_B(net7436),
    .D(_00453_),
    .Q(\trng_data[4] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _48810_ (.RESET_B(net7437),
    .D(_00454_),
    .Q(\trng_data[5] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _48811_ (.RESET_B(net7437),
    .D(net1918),
    .Q(\trng_data[6] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _48812_ (.RESET_B(net7437),
    .D(net1362),
    .Q(\trng_data[7] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _48813_ (.RESET_B(net7436),
    .D(\u_trng.entropy_raw ),
    .Q(\u_trng.entropy_ff1 ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _48814_ (.RESET_B(net7435),
    .D(net1177),
    .Q(\u_trng.have_prev ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _48815_ (.RESET_B(net7437),
    .D(net2543),
    .Q(\u_trng.prev_sample ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _48816_ (.RESET_B(net7435),
    .D(net1223),
    .Q(trng_ready),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _48817_ (.RESET_B(net7450),
    .D(net1148),
    .Q(\u_inv.input_valid ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _48818_ (.RESET_B(net7435),
    .D(net1146),
    .Q(\u_trng.entropy_bit ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _48819_ (.RESET_B(net136),
    .D(_00460_),
    .Q(\u_inv.f_next[0] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _48820_ (.RESET_B(net135),
    .D(_00461_),
    .Q(\u_inv.f_next[1] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_2 _48821_ (.RESET_B(net134),
    .D(_00462_),
    .Q(\u_inv.f_next[2] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _48822_ (.RESET_B(net133),
    .D(_00463_),
    .Q(\u_inv.f_next[3] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _48823_ (.RESET_B(net132),
    .D(_00464_),
    .Q(\u_inv.f_next[4] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _48824_ (.RESET_B(net131),
    .D(_00465_),
    .Q(\u_inv.f_next[5] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _48825_ (.RESET_B(net130),
    .D(_00466_),
    .Q(\u_inv.f_next[6] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _48826_ (.RESET_B(net129),
    .D(_00467_),
    .Q(\u_inv.f_next[7] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _48827_ (.RESET_B(net128),
    .D(_00468_),
    .Q(\u_inv.f_next[8] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _48828_ (.RESET_B(net127),
    .D(_00469_),
    .Q(\u_inv.f_next[9] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _48829_ (.RESET_B(net126),
    .D(_00470_),
    .Q(\u_inv.f_next[10] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _48830_ (.RESET_B(net125),
    .D(_00471_),
    .Q(\u_inv.f_next[11] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _48831_ (.RESET_B(net124),
    .D(_00472_),
    .Q(\u_inv.f_next[12] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _48832_ (.RESET_B(net123),
    .D(_00473_),
    .Q(\u_inv.f_next[13] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _48833_ (.RESET_B(net122),
    .D(_00474_),
    .Q(\u_inv.f_next[14] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _48834_ (.RESET_B(net121),
    .D(_00475_),
    .Q(\u_inv.f_next[15] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _48835_ (.RESET_B(net120),
    .D(_00476_),
    .Q(\u_inv.f_next[16] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _48836_ (.RESET_B(net119),
    .D(_00477_),
    .Q(\u_inv.f_next[17] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _48837_ (.RESET_B(net118),
    .D(_00478_),
    .Q(\u_inv.f_next[18] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _48838_ (.RESET_B(net117),
    .D(_00479_),
    .Q(\u_inv.f_next[19] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _48839_ (.RESET_B(net116),
    .D(_00480_),
    .Q(\u_inv.f_next[20] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _48840_ (.RESET_B(net115),
    .D(_00481_),
    .Q(\u_inv.f_next[21] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _48841_ (.RESET_B(net114),
    .D(_00482_),
    .Q(\u_inv.f_next[22] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _48842_ (.RESET_B(net113),
    .D(_00483_),
    .Q(\u_inv.f_next[23] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _48843_ (.RESET_B(net112),
    .D(_00484_),
    .Q(\u_inv.f_next[24] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _48844_ (.RESET_B(net111),
    .D(_00485_),
    .Q(\u_inv.f_next[25] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _48845_ (.RESET_B(net110),
    .D(_00486_),
    .Q(\u_inv.f_next[26] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _48846_ (.RESET_B(net109),
    .D(_00487_),
    .Q(\u_inv.f_next[27] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _48847_ (.RESET_B(net108),
    .D(_00488_),
    .Q(\u_inv.f_next[28] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _48848_ (.RESET_B(net107),
    .D(_00489_),
    .Q(\u_inv.f_next[29] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _48849_ (.RESET_B(net106),
    .D(_00490_),
    .Q(\u_inv.f_next[30] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _48850_ (.RESET_B(net105),
    .D(_00491_),
    .Q(\u_inv.f_next[31] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _48851_ (.RESET_B(net104),
    .D(_00492_),
    .Q(\u_inv.f_next[32] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_2 _48852_ (.RESET_B(net103),
    .D(_00493_),
    .Q(\u_inv.f_next[33] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _48853_ (.RESET_B(net102),
    .D(_00494_),
    .Q(\u_inv.f_next[34] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_2 _48854_ (.RESET_B(net101),
    .D(_00495_),
    .Q(\u_inv.f_next[35] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _48855_ (.RESET_B(net100),
    .D(_00496_),
    .Q(\u_inv.f_next[36] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _48856_ (.RESET_B(net99),
    .D(net1447),
    .Q(\u_inv.f_next[37] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _48857_ (.RESET_B(net98),
    .D(_00498_),
    .Q(\u_inv.f_next[38] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_2 _48858_ (.RESET_B(net97),
    .D(_00499_),
    .Q(\u_inv.f_next[39] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_2 _48859_ (.RESET_B(net96),
    .D(_00500_),
    .Q(\u_inv.f_next[40] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_2 _48860_ (.RESET_B(net95),
    .D(_00501_),
    .Q(\u_inv.f_next[41] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_2 _48861_ (.RESET_B(net94),
    .D(_00502_),
    .Q(\u_inv.f_next[42] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_2 _48862_ (.RESET_B(net93),
    .D(_00503_),
    .Q(\u_inv.f_next[43] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_2 _48863_ (.RESET_B(net92),
    .D(_00504_),
    .Q(\u_inv.f_next[44] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_2 _48864_ (.RESET_B(net91),
    .D(net1285),
    .Q(\u_inv.f_next[45] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_2 _48865_ (.RESET_B(net90),
    .D(_00506_),
    .Q(\u_inv.f_next[46] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_2 _48866_ (.RESET_B(net89),
    .D(_00507_),
    .Q(\u_inv.f_next[47] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_2 _48867_ (.RESET_B(net88),
    .D(_00508_),
    .Q(\u_inv.f_next[48] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_2 _48868_ (.RESET_B(net87),
    .D(_00509_),
    .Q(\u_inv.f_next[49] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_2 _48869_ (.RESET_B(net86),
    .D(_00510_),
    .Q(\u_inv.f_next[50] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_2 _48870_ (.RESET_B(net85),
    .D(_00511_),
    .Q(\u_inv.f_next[51] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_2 _48871_ (.RESET_B(net84),
    .D(_00512_),
    .Q(\u_inv.f_next[52] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_2 _48872_ (.RESET_B(net83),
    .D(_00513_),
    .Q(\u_inv.f_next[53] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_2 _48873_ (.RESET_B(net82),
    .D(_00514_),
    .Q(\u_inv.f_next[54] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_2 _48874_ (.RESET_B(net81),
    .D(_00515_),
    .Q(\u_inv.f_next[55] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_2 _48875_ (.RESET_B(net80),
    .D(_00516_),
    .Q(\u_inv.f_next[56] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_2 _48876_ (.RESET_B(net79),
    .D(_00517_),
    .Q(\u_inv.f_next[57] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_2 _48877_ (.RESET_B(net78),
    .D(_00518_),
    .Q(\u_inv.f_next[58] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_2 _48878_ (.RESET_B(net77),
    .D(_00519_),
    .Q(\u_inv.f_next[59] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _48879_ (.RESET_B(net76),
    .D(_00520_),
    .Q(\u_inv.f_next[60] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_2 _48880_ (.RESET_B(net75),
    .D(_00521_),
    .Q(\u_inv.f_next[61] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _48881_ (.RESET_B(net74),
    .D(_00522_),
    .Q(\u_inv.f_next[62] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_2 _48882_ (.RESET_B(net73),
    .D(_00523_),
    .Q(\u_inv.f_next[63] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_2 _48883_ (.RESET_B(net72),
    .D(_00524_),
    .Q(\u_inv.f_next[64] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_2 _48884_ (.RESET_B(net71),
    .D(_00525_),
    .Q(\u_inv.f_next[65] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_2 _48885_ (.RESET_B(net70),
    .D(_00526_),
    .Q(\u_inv.f_next[66] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_2 _48886_ (.RESET_B(net69),
    .D(_00527_),
    .Q(\u_inv.f_next[67] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_2 _48887_ (.RESET_B(net68),
    .D(_00528_),
    .Q(\u_inv.f_next[68] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_2 _48888_ (.RESET_B(net67),
    .D(_00529_),
    .Q(\u_inv.f_next[69] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_2 _48889_ (.RESET_B(net66),
    .D(_00530_),
    .Q(\u_inv.f_next[70] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_2 _48890_ (.RESET_B(net65),
    .D(_00531_),
    .Q(\u_inv.f_next[71] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_2 _48891_ (.RESET_B(net64),
    .D(_00532_),
    .Q(\u_inv.f_next[72] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_2 _48892_ (.RESET_B(net63),
    .D(_00533_),
    .Q(\u_inv.f_next[73] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_2 _48893_ (.RESET_B(net62),
    .D(_00534_),
    .Q(\u_inv.f_next[74] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_2 _48894_ (.RESET_B(net61),
    .D(_00535_),
    .Q(\u_inv.f_next[75] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_2 _48895_ (.RESET_B(net60),
    .D(_00536_),
    .Q(\u_inv.f_next[76] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_2 _48896_ (.RESET_B(net59),
    .D(_00537_),
    .Q(\u_inv.f_next[77] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_2 _48897_ (.RESET_B(net58),
    .D(_00538_),
    .Q(\u_inv.f_next[78] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_2 _48898_ (.RESET_B(net57),
    .D(_00539_),
    .Q(\u_inv.f_next[79] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_2 _48899_ (.RESET_B(net56),
    .D(_00540_),
    .Q(\u_inv.f_next[80] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_2 _48900_ (.RESET_B(net55),
    .D(_00541_),
    .Q(\u_inv.f_next[81] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_2 _48901_ (.RESET_B(net54),
    .D(_00542_),
    .Q(\u_inv.f_next[82] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_2 _48902_ (.RESET_B(net53),
    .D(_00543_),
    .Q(\u_inv.f_next[83] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_2 _48903_ (.RESET_B(net52),
    .D(_00544_),
    .Q(\u_inv.f_next[84] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_2 _48904_ (.RESET_B(net51),
    .D(_00545_),
    .Q(\u_inv.f_next[85] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _48905_ (.RESET_B(net50),
    .D(_00546_),
    .Q(\u_inv.f_next[86] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _48906_ (.RESET_B(net49),
    .D(_00547_),
    .Q(\u_inv.f_next[87] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_2 _48907_ (.RESET_B(net48),
    .D(_00548_),
    .Q(\u_inv.f_next[88] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_2 _48908_ (.RESET_B(net47),
    .D(_00549_),
    .Q(\u_inv.f_next[89] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_2 _48909_ (.RESET_B(net46),
    .D(_00550_),
    .Q(\u_inv.f_next[90] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_2 _48910_ (.RESET_B(net45),
    .D(_00551_),
    .Q(\u_inv.f_next[91] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_2 _48911_ (.RESET_B(net44),
    .D(_00552_),
    .Q(\u_inv.f_next[92] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_2 _48912_ (.RESET_B(net43),
    .D(_00553_),
    .Q(\u_inv.f_next[93] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _48913_ (.RESET_B(net42),
    .D(_00554_),
    .Q(\u_inv.f_next[94] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_2 _48914_ (.RESET_B(net41),
    .D(_00555_),
    .Q(\u_inv.f_next[95] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_2 _48915_ (.RESET_B(net40),
    .D(_00556_),
    .Q(\u_inv.f_next[96] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_2 _48916_ (.RESET_B(net39),
    .D(_00557_),
    .Q(\u_inv.f_next[97] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_2 _48917_ (.RESET_B(net38),
    .D(_00558_),
    .Q(\u_inv.f_next[98] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_2 _48918_ (.RESET_B(net37),
    .D(_00559_),
    .Q(\u_inv.f_next[99] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _48919_ (.RESET_B(net36),
    .D(_00560_),
    .Q(\u_inv.f_next[100] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _48920_ (.RESET_B(net35),
    .D(_00561_),
    .Q(\u_inv.f_next[101] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_2 _48921_ (.RESET_B(net34),
    .D(_00562_),
    .Q(\u_inv.f_next[102] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_2 _48922_ (.RESET_B(net33),
    .D(_00563_),
    .Q(\u_inv.f_next[103] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _48923_ (.RESET_B(net32),
    .D(_00564_),
    .Q(\u_inv.f_next[104] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _48924_ (.RESET_B(net31),
    .D(_00565_),
    .Q(\u_inv.f_next[105] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _48925_ (.RESET_B(net30),
    .D(_00566_),
    .Q(\u_inv.f_next[106] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_2 _48926_ (.RESET_B(net29),
    .D(_00567_),
    .Q(\u_inv.f_next[107] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_2 _48927_ (.RESET_B(net28),
    .D(_00568_),
    .Q(\u_inv.f_next[108] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _48928_ (.RESET_B(net27),
    .D(_00569_),
    .Q(\u_inv.f_next[109] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _48929_ (.RESET_B(net26),
    .D(_00570_),
    .Q(\u_inv.f_next[110] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _48930_ (.RESET_B(net25),
    .D(_00571_),
    .Q(\u_inv.f_next[111] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _48931_ (.RESET_B(net24),
    .D(_00572_),
    .Q(\u_inv.f_next[112] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_2 _48932_ (.RESET_B(net23),
    .D(_00573_),
    .Q(\u_inv.f_next[113] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _48933_ (.RESET_B(net22),
    .D(_00574_),
    .Q(\u_inv.f_next[114] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _48934_ (.RESET_B(net21),
    .D(_00575_),
    .Q(\u_inv.f_next[115] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _48935_ (.RESET_B(net1058),
    .D(net2144),
    .Q(\u_inv.f_next[116] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _48936_ (.RESET_B(net1057),
    .D(_00577_),
    .Q(\u_inv.f_next[117] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_2 _48937_ (.RESET_B(net1056),
    .D(_00578_),
    .Q(\u_inv.f_next[118] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _48938_ (.RESET_B(net1055),
    .D(_00579_),
    .Q(\u_inv.f_next[119] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_2 _48939_ (.RESET_B(net1054),
    .D(_00580_),
    .Q(\u_inv.f_next[120] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_2 _48940_ (.RESET_B(net1053),
    .D(_00581_),
    .Q(\u_inv.f_next[121] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_2 _48941_ (.RESET_B(net1052),
    .D(_00582_),
    .Q(\u_inv.f_next[122] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_2 _48942_ (.RESET_B(net1051),
    .D(_00583_),
    .Q(\u_inv.f_next[123] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_2 _48943_ (.RESET_B(net1050),
    .D(_00584_),
    .Q(\u_inv.f_next[124] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _48944_ (.RESET_B(net1049),
    .D(_00585_),
    .Q(\u_inv.f_next[125] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _48945_ (.RESET_B(net1048),
    .D(_00586_),
    .Q(\u_inv.f_next[126] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_2 _48946_ (.RESET_B(net1047),
    .D(_00587_),
    .Q(\u_inv.f_next[127] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_2 _48947_ (.RESET_B(net1046),
    .D(_00588_),
    .Q(\u_inv.f_next[128] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_2 _48948_ (.RESET_B(net1045),
    .D(_00589_),
    .Q(\u_inv.f_next[129] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_2 _48949_ (.RESET_B(net1044),
    .D(_00590_),
    .Q(\u_inv.f_next[130] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _48950_ (.RESET_B(net1043),
    .D(_00591_),
    .Q(\u_inv.f_next[131] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _48951_ (.RESET_B(net1042),
    .D(_00592_),
    .Q(\u_inv.f_next[132] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _48952_ (.RESET_B(net1041),
    .D(_00593_),
    .Q(\u_inv.f_next[133] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _48953_ (.RESET_B(net1040),
    .D(_00594_),
    .Q(\u_inv.f_next[134] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _48954_ (.RESET_B(net1039),
    .D(_00595_),
    .Q(\u_inv.f_next[135] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _48955_ (.RESET_B(net1038),
    .D(_00596_),
    .Q(\u_inv.f_next[136] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _48956_ (.RESET_B(net1037),
    .D(_00597_),
    .Q(\u_inv.f_next[137] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _48957_ (.RESET_B(net1036),
    .D(_00598_),
    .Q(\u_inv.f_next[138] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _48958_ (.RESET_B(net1035),
    .D(_00599_),
    .Q(\u_inv.f_next[139] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _48959_ (.RESET_B(net1034),
    .D(_00600_),
    .Q(\u_inv.f_next[140] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _48960_ (.RESET_B(net1033),
    .D(_00601_),
    .Q(\u_inv.f_next[141] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _48961_ (.RESET_B(net1032),
    .D(_00602_),
    .Q(\u_inv.f_next[142] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _48962_ (.RESET_B(net1031),
    .D(_00603_),
    .Q(\u_inv.f_next[143] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _48963_ (.RESET_B(net1030),
    .D(_00604_),
    .Q(\u_inv.f_next[144] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _48964_ (.RESET_B(net1029),
    .D(net1474),
    .Q(\u_inv.f_next[145] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _48965_ (.RESET_B(net1028),
    .D(_00606_),
    .Q(\u_inv.f_next[146] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _48966_ (.RESET_B(net1027),
    .D(_00607_),
    .Q(\u_inv.f_next[147] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _48967_ (.RESET_B(net1026),
    .D(_00608_),
    .Q(\u_inv.f_next[148] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _48968_ (.RESET_B(net1025),
    .D(_00609_),
    .Q(\u_inv.f_next[149] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _48969_ (.RESET_B(net1024),
    .D(_00610_),
    .Q(\u_inv.f_next[150] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _48970_ (.RESET_B(net1023),
    .D(_00611_),
    .Q(\u_inv.f_next[151] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _48971_ (.RESET_B(net1022),
    .D(_00612_),
    .Q(\u_inv.f_next[152] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _48972_ (.RESET_B(net1021),
    .D(_00613_),
    .Q(\u_inv.f_next[153] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _48973_ (.RESET_B(net1020),
    .D(_00614_),
    .Q(\u_inv.f_next[154] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _48974_ (.RESET_B(net1019),
    .D(_00615_),
    .Q(\u_inv.f_next[155] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _48975_ (.RESET_B(net1018),
    .D(_00616_),
    .Q(\u_inv.f_next[156] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _48976_ (.RESET_B(net1017),
    .D(_00617_),
    .Q(\u_inv.f_next[157] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _48977_ (.RESET_B(net1016),
    .D(_00618_),
    .Q(\u_inv.f_next[158] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _48978_ (.RESET_B(net1015),
    .D(_00619_),
    .Q(\u_inv.f_next[159] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _48979_ (.RESET_B(net1014),
    .D(_00620_),
    .Q(\u_inv.f_next[160] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _48980_ (.RESET_B(net1013),
    .D(_00621_),
    .Q(\u_inv.f_next[161] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _48981_ (.RESET_B(net1012),
    .D(_00622_),
    .Q(\u_inv.f_next[162] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _48982_ (.RESET_B(net1011),
    .D(net3007),
    .Q(\u_inv.f_next[163] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _48983_ (.RESET_B(net1010),
    .D(_00624_),
    .Q(\u_inv.f_next[164] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _48984_ (.RESET_B(net1009),
    .D(net1512),
    .Q(\u_inv.f_next[165] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _48985_ (.RESET_B(net1008),
    .D(_00626_),
    .Q(\u_inv.f_next[166] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _48986_ (.RESET_B(net1007),
    .D(_00627_),
    .Q(\u_inv.f_next[167] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _48987_ (.RESET_B(net1006),
    .D(_00628_),
    .Q(\u_inv.f_next[168] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _48988_ (.RESET_B(net1005),
    .D(_00629_),
    .Q(\u_inv.f_next[169] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _48989_ (.RESET_B(net1004),
    .D(_00630_),
    .Q(\u_inv.f_next[170] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _48990_ (.RESET_B(net1003),
    .D(_00631_),
    .Q(\u_inv.f_next[171] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _48991_ (.RESET_B(net1002),
    .D(_00632_),
    .Q(\u_inv.f_next[172] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _48992_ (.RESET_B(net1001),
    .D(_00633_),
    .Q(\u_inv.f_next[173] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _48993_ (.RESET_B(net1000),
    .D(_00634_),
    .Q(\u_inv.f_next[174] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _48994_ (.RESET_B(net999),
    .D(_00635_),
    .Q(\u_inv.f_next[175] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _48995_ (.RESET_B(net998),
    .D(_00636_),
    .Q(\u_inv.f_next[176] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _48996_ (.RESET_B(net997),
    .D(_00637_),
    .Q(\u_inv.f_next[177] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _48997_ (.RESET_B(net996),
    .D(_00638_),
    .Q(\u_inv.f_next[178] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _48998_ (.RESET_B(net995),
    .D(_00639_),
    .Q(\u_inv.f_next[179] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _48999_ (.RESET_B(net994),
    .D(_00640_),
    .Q(\u_inv.f_next[180] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _49000_ (.RESET_B(net993),
    .D(_00641_),
    .Q(\u_inv.f_next[181] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _49001_ (.RESET_B(net992),
    .D(_00642_),
    .Q(\u_inv.f_next[182] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_2 _49002_ (.RESET_B(net991),
    .D(_00643_),
    .Q(\u_inv.f_next[183] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _49003_ (.RESET_B(net990),
    .D(_00644_),
    .Q(\u_inv.f_next[184] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _49004_ (.RESET_B(net989),
    .D(_00645_),
    .Q(\u_inv.f_next[185] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_2 _49005_ (.RESET_B(net988),
    .D(_00646_),
    .Q(\u_inv.f_next[186] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_2 _49006_ (.RESET_B(net987),
    .D(_00647_),
    .Q(\u_inv.f_next[187] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_2 _49007_ (.RESET_B(net986),
    .D(_00648_),
    .Q(\u_inv.f_next[188] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_2 _49008_ (.RESET_B(net985),
    .D(_00649_),
    .Q(\u_inv.f_next[189] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_2 _49009_ (.RESET_B(net984),
    .D(_00650_),
    .Q(\u_inv.f_next[190] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_2 _49010_ (.RESET_B(net983),
    .D(_00651_),
    .Q(\u_inv.f_next[191] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_2 _49011_ (.RESET_B(net982),
    .D(_00652_),
    .Q(\u_inv.f_next[192] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_2 _49012_ (.RESET_B(net981),
    .D(_00653_),
    .Q(\u_inv.f_next[193] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_2 _49013_ (.RESET_B(net980),
    .D(_00654_),
    .Q(\u_inv.f_next[194] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_2 _49014_ (.RESET_B(net979),
    .D(_00655_),
    .Q(\u_inv.f_next[195] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_2 _49015_ (.RESET_B(net978),
    .D(_00656_),
    .Q(\u_inv.f_next[196] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_2 _49016_ (.RESET_B(net977),
    .D(_00657_),
    .Q(\u_inv.f_next[197] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_2 _49017_ (.RESET_B(net976),
    .D(_00658_),
    .Q(\u_inv.f_next[198] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_2 _49018_ (.RESET_B(net975),
    .D(_00659_),
    .Q(\u_inv.f_next[199] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _49019_ (.RESET_B(net974),
    .D(_00660_),
    .Q(\u_inv.f_next[200] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _49020_ (.RESET_B(net973),
    .D(_00661_),
    .Q(\u_inv.f_next[201] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_2 _49021_ (.RESET_B(net972),
    .D(_00662_),
    .Q(\u_inv.f_next[202] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_2 _49022_ (.RESET_B(net971),
    .D(_00663_),
    .Q(\u_inv.f_next[203] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_2 _49023_ (.RESET_B(net970),
    .D(_00664_),
    .Q(\u_inv.f_next[204] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_2 _49024_ (.RESET_B(net969),
    .D(net1927),
    .Q(\u_inv.f_next[205] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _49025_ (.RESET_B(net968),
    .D(_00666_),
    .Q(\u_inv.f_next[206] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _49026_ (.RESET_B(net967),
    .D(_00667_),
    .Q(\u_inv.f_next[207] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _49027_ (.RESET_B(net966),
    .D(_00668_),
    .Q(\u_inv.f_next[208] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_2 _49028_ (.RESET_B(net965),
    .D(_00669_),
    .Q(\u_inv.f_next[209] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _49029_ (.RESET_B(net964),
    .D(_00670_),
    .Q(\u_inv.f_next[210] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _49030_ (.RESET_B(net963),
    .D(_00671_),
    .Q(\u_inv.f_next[211] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_2 _49031_ (.RESET_B(net962),
    .D(_00672_),
    .Q(\u_inv.f_next[212] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _49032_ (.RESET_B(net961),
    .D(_00673_),
    .Q(\u_inv.f_next[213] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _49033_ (.RESET_B(net960),
    .D(_00674_),
    .Q(\u_inv.f_next[214] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _49034_ (.RESET_B(net959),
    .D(_00675_),
    .Q(\u_inv.f_next[215] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_2 _49035_ (.RESET_B(net958),
    .D(_00676_),
    .Q(\u_inv.f_next[216] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _49036_ (.RESET_B(net957),
    .D(_00677_),
    .Q(\u_inv.f_next[217] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _49037_ (.RESET_B(net956),
    .D(_00678_),
    .Q(\u_inv.f_next[218] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _49038_ (.RESET_B(net955),
    .D(net1727),
    .Q(\u_inv.f_next[219] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _49039_ (.RESET_B(net954),
    .D(_00680_),
    .Q(\u_inv.f_next[220] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _49040_ (.RESET_B(net953),
    .D(_00681_),
    .Q(\u_inv.f_next[221] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _49041_ (.RESET_B(net952),
    .D(_00682_),
    .Q(\u_inv.f_next[222] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _49042_ (.RESET_B(net951),
    .D(_00683_),
    .Q(\u_inv.f_next[223] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _49043_ (.RESET_B(net950),
    .D(_00684_),
    .Q(\u_inv.f_next[224] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _49044_ (.RESET_B(net949),
    .D(_00685_),
    .Q(\u_inv.f_next[225] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _49045_ (.RESET_B(net948),
    .D(_00686_),
    .Q(\u_inv.f_next[226] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _49046_ (.RESET_B(net947),
    .D(_00687_),
    .Q(\u_inv.f_next[227] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _49047_ (.RESET_B(net946),
    .D(_00688_),
    .Q(\u_inv.f_next[228] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _49048_ (.RESET_B(net945),
    .D(_00689_),
    .Q(\u_inv.f_next[229] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _49049_ (.RESET_B(net944),
    .D(_00690_),
    .Q(\u_inv.f_next[230] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _49050_ (.RESET_B(net943),
    .D(_00691_),
    .Q(\u_inv.f_next[231] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _49051_ (.RESET_B(net942),
    .D(_00692_),
    .Q(\u_inv.f_next[232] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _49052_ (.RESET_B(net941),
    .D(_00693_),
    .Q(\u_inv.f_next[233] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _49053_ (.RESET_B(net940),
    .D(_00694_),
    .Q(\u_inv.f_next[234] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _49054_ (.RESET_B(net939),
    .D(_00695_),
    .Q(\u_inv.f_next[235] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _49055_ (.RESET_B(net938),
    .D(_00696_),
    .Q(\u_inv.f_next[236] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _49056_ (.RESET_B(net937),
    .D(_00697_),
    .Q(\u_inv.f_next[237] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _49057_ (.RESET_B(net936),
    .D(_00698_),
    .Q(\u_inv.f_next[238] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _49058_ (.RESET_B(net935),
    .D(_00699_),
    .Q(\u_inv.f_next[239] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _49059_ (.RESET_B(net934),
    .D(_00700_),
    .Q(\u_inv.f_next[240] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _49060_ (.RESET_B(net933),
    .D(_00701_),
    .Q(\u_inv.f_next[241] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _49061_ (.RESET_B(net932),
    .D(_00702_),
    .Q(\u_inv.f_next[242] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _49062_ (.RESET_B(net931),
    .D(_00703_),
    .Q(\u_inv.f_next[243] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _49063_ (.RESET_B(net930),
    .D(_00704_),
    .Q(\u_inv.f_next[244] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _49064_ (.RESET_B(net929),
    .D(_00705_),
    .Q(\u_inv.f_next[245] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _49065_ (.RESET_B(net928),
    .D(_00706_),
    .Q(\u_inv.f_next[246] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _49066_ (.RESET_B(net927),
    .D(_00707_),
    .Q(\u_inv.f_next[247] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _49067_ (.RESET_B(net926),
    .D(_00708_),
    .Q(\u_inv.f_next[248] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _49068_ (.RESET_B(net925),
    .D(_00709_),
    .Q(\u_inv.f_next[249] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _49069_ (.RESET_B(net924),
    .D(_00710_),
    .Q(\u_inv.f_next[250] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _49070_ (.RESET_B(net923),
    .D(_00711_),
    .Q(\u_inv.f_next[251] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _49071_ (.RESET_B(net922),
    .D(_00712_),
    .Q(\u_inv.f_next[252] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _49072_ (.RESET_B(net921),
    .D(_00713_),
    .Q(\u_inv.f_next[253] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _49073_ (.RESET_B(net920),
    .D(_00714_),
    .Q(\u_inv.f_next[254] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _49074_ (.RESET_B(net919),
    .D(_00715_),
    .Q(\u_inv.f_next[255] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _49075_ (.RESET_B(net918),
    .D(_00716_),
    .Q(\u_inv.f_next[256] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _49076_ (.RESET_B(net7441),
    .D(_00717_),
    .Q(\perf_double[0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _49077_ (.RESET_B(net7441),
    .D(_00718_),
    .Q(\perf_double[1] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _49078_ (.RESET_B(net7441),
    .D(_00719_),
    .Q(\perf_double[2] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _49079_ (.RESET_B(net7442),
    .D(_00720_),
    .Q(\perf_double[3] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _49080_ (.RESET_B(net7441),
    .D(_00721_),
    .Q(\perf_double[4] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _49081_ (.RESET_B(net7442),
    .D(_00722_),
    .Q(\perf_double[5] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _49082_ (.RESET_B(net7432),
    .D(_00723_),
    .Q(\perf_double[6] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _49083_ (.RESET_B(net7443),
    .D(_00724_),
    .Q(\perf_double[7] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _49084_ (.RESET_B(net7443),
    .D(_00725_),
    .Q(\perf_double[8] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _49085_ (.RESET_B(net7443),
    .D(_00726_),
    .Q(\perf_double[9] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _49086_ (.RESET_B(net7449),
    .D(net1770),
    .Q(inv_done),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _49087_ (.RESET_B(net7443),
    .D(_00727_),
    .Q(\perf_total[0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _49088_ (.RESET_B(net7443),
    .D(_00728_),
    .Q(\perf_total[1] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _49089_ (.RESET_B(net7443),
    .D(net1267),
    .Q(\perf_total[2] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _49090_ (.RESET_B(net7448),
    .D(net1162),
    .Q(\perf_total[3] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _49091_ (.RESET_B(net7448),
    .D(net1195),
    .Q(\perf_total[4] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _49092_ (.RESET_B(net7448),
    .D(net1156),
    .Q(\perf_total[5] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _49093_ (.RESET_B(net7448),
    .D(_00733_),
    .Q(\perf_total[6] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _49094_ (.RESET_B(net7448),
    .D(_00734_),
    .Q(\perf_total[7] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _49095_ (.RESET_B(net7449),
    .D(_00735_),
    .Q(\perf_total[8] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _49096_ (.RESET_B(net7449),
    .D(net1281),
    .Q(\perf_total[9] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _49097_ (.RESET_B(net916),
    .D(_00737_),
    .Q(\u_inv.d_next[0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _49098_ (.RESET_B(net915),
    .D(_00738_),
    .Q(\u_inv.d_next[1] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _49099_ (.RESET_B(net913),
    .D(_00739_),
    .Q(\u_inv.d_next[2] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _49100_ (.RESET_B(net911),
    .D(_00740_),
    .Q(\u_inv.d_next[3] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _49101_ (.RESET_B(net909),
    .D(_00741_),
    .Q(\u_inv.d_next[4] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _49102_ (.RESET_B(net908),
    .D(_00742_),
    .Q(\u_inv.d_next[5] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _49103_ (.RESET_B(net906),
    .D(_00743_),
    .Q(\u_inv.d_next[6] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _49104_ (.RESET_B(net904),
    .D(_00744_),
    .Q(\u_inv.d_next[7] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _49105_ (.RESET_B(net902),
    .D(_00745_),
    .Q(\u_inv.d_next[8] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _49106_ (.RESET_B(net901),
    .D(_00746_),
    .Q(\u_inv.d_next[9] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _49107_ (.RESET_B(net899),
    .D(_00747_),
    .Q(\u_inv.d_next[10] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _49108_ (.RESET_B(net897),
    .D(_00748_),
    .Q(\u_inv.d_next[11] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _49109_ (.RESET_B(net895),
    .D(_00749_),
    .Q(\u_inv.d_next[12] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _49110_ (.RESET_B(net894),
    .D(_00750_),
    .Q(\u_inv.d_next[13] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _49111_ (.RESET_B(net892),
    .D(_00751_),
    .Q(\u_inv.d_next[14] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _49112_ (.RESET_B(net890),
    .D(_00752_),
    .Q(\u_inv.d_next[15] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _49113_ (.RESET_B(net888),
    .D(_00753_),
    .Q(\u_inv.d_next[16] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _49114_ (.RESET_B(net887),
    .D(_00754_),
    .Q(\u_inv.d_next[17] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_1 _49115_ (.RESET_B(net885),
    .D(_00755_),
    .Q(\u_inv.d_next[18] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _49116_ (.RESET_B(net883),
    .D(_00756_),
    .Q(\u_inv.d_next[19] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _49117_ (.RESET_B(net881),
    .D(_00757_),
    .Q(\u_inv.d_next[20] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _49118_ (.RESET_B(net880),
    .D(_00758_),
    .Q(\u_inv.d_next[21] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_2 _49119_ (.RESET_B(net878),
    .D(_00759_),
    .Q(\u_inv.d_next[22] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _49120_ (.RESET_B(net876),
    .D(_00760_),
    .Q(\u_inv.d_next[23] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_2 _49121_ (.RESET_B(net874),
    .D(_00761_),
    .Q(\u_inv.d_next[24] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_2 _49122_ (.RESET_B(net873),
    .D(_00762_),
    .Q(\u_inv.d_next[25] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _49123_ (.RESET_B(net871),
    .D(_00763_),
    .Q(\u_inv.d_next[26] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_2 _49124_ (.RESET_B(net869),
    .D(_00764_),
    .Q(\u_inv.d_next[27] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_2 _49125_ (.RESET_B(net867),
    .D(_00765_),
    .Q(\u_inv.d_next[28] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_2 _49126_ (.RESET_B(net866),
    .D(_00766_),
    .Q(\u_inv.d_next[29] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_2 _49127_ (.RESET_B(net864),
    .D(_00767_),
    .Q(\u_inv.d_next[30] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _49128_ (.RESET_B(net862),
    .D(_00768_),
    .Q(\u_inv.d_next[31] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _49129_ (.RESET_B(net860),
    .D(_00769_),
    .Q(\u_inv.d_next[32] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _49130_ (.RESET_B(net859),
    .D(_00770_),
    .Q(\u_inv.d_next[33] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _49131_ (.RESET_B(net857),
    .D(_00771_),
    .Q(\u_inv.d_next[34] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _49132_ (.RESET_B(net855),
    .D(_00772_),
    .Q(\u_inv.d_next[35] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _49133_ (.RESET_B(net853),
    .D(_00773_),
    .Q(\u_inv.d_next[36] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _49134_ (.RESET_B(net852),
    .D(_00774_),
    .Q(\u_inv.d_next[37] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _49135_ (.RESET_B(net850),
    .D(_00775_),
    .Q(\u_inv.d_next[38] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _49136_ (.RESET_B(net848),
    .D(_00776_),
    .Q(\u_inv.d_next[39] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _49137_ (.RESET_B(net846),
    .D(_00777_),
    .Q(\u_inv.d_next[40] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _49138_ (.RESET_B(net845),
    .D(_00778_),
    .Q(\u_inv.d_next[41] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _49139_ (.RESET_B(net843),
    .D(_00779_),
    .Q(\u_inv.d_next[42] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _49140_ (.RESET_B(net841),
    .D(_00780_),
    .Q(\u_inv.d_next[43] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _49141_ (.RESET_B(net839),
    .D(_00781_),
    .Q(\u_inv.d_next[44] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _49142_ (.RESET_B(net838),
    .D(_00782_),
    .Q(\u_inv.d_next[45] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _49143_ (.RESET_B(net836),
    .D(_00783_),
    .Q(\u_inv.d_next[46] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _49144_ (.RESET_B(net834),
    .D(_00784_),
    .Q(\u_inv.d_next[47] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _49145_ (.RESET_B(net832),
    .D(_00785_),
    .Q(\u_inv.d_next[48] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _49146_ (.RESET_B(net831),
    .D(_00786_),
    .Q(\u_inv.d_next[49] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _49147_ (.RESET_B(net829),
    .D(_00787_),
    .Q(\u_inv.d_next[50] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _49148_ (.RESET_B(net827),
    .D(_00788_),
    .Q(\u_inv.d_next[51] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _49149_ (.RESET_B(net825),
    .D(_00789_),
    .Q(\u_inv.d_next[52] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _49150_ (.RESET_B(net824),
    .D(_00790_),
    .Q(\u_inv.d_next[53] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _49151_ (.RESET_B(net822),
    .D(_00791_),
    .Q(\u_inv.d_next[54] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _49152_ (.RESET_B(net820),
    .D(_00792_),
    .Q(\u_inv.d_next[55] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _49153_ (.RESET_B(net818),
    .D(_00793_),
    .Q(\u_inv.d_next[56] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _49154_ (.RESET_B(net817),
    .D(_00794_),
    .Q(\u_inv.d_next[57] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _49155_ (.RESET_B(net815),
    .D(_00795_),
    .Q(\u_inv.d_next[58] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _49156_ (.RESET_B(net813),
    .D(_00796_),
    .Q(\u_inv.d_next[59] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _49157_ (.RESET_B(net811),
    .D(_00797_),
    .Q(\u_inv.d_next[60] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _49158_ (.RESET_B(net810),
    .D(_00798_),
    .Q(\u_inv.d_next[61] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _49159_ (.RESET_B(net808),
    .D(_00799_),
    .Q(\u_inv.d_next[62] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _49160_ (.RESET_B(net806),
    .D(_00800_),
    .Q(\u_inv.d_next[63] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _49161_ (.RESET_B(net804),
    .D(_00801_),
    .Q(\u_inv.d_next[64] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _49162_ (.RESET_B(net803),
    .D(_00802_),
    .Q(\u_inv.d_next[65] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _49163_ (.RESET_B(net801),
    .D(_00803_),
    .Q(\u_inv.d_next[66] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _49164_ (.RESET_B(net799),
    .D(_00804_),
    .Q(\u_inv.d_next[67] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _49165_ (.RESET_B(net797),
    .D(_00805_),
    .Q(\u_inv.d_next[68] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _49166_ (.RESET_B(net796),
    .D(_00806_),
    .Q(\u_inv.d_next[69] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_1 _49167_ (.RESET_B(net794),
    .D(_00807_),
    .Q(\u_inv.d_next[70] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _49168_ (.RESET_B(net792),
    .D(_00808_),
    .Q(\u_inv.d_next[71] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _49169_ (.RESET_B(net790),
    .D(_00809_),
    .Q(\u_inv.d_next[72] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _49170_ (.RESET_B(net789),
    .D(_00810_),
    .Q(\u_inv.d_next[73] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _49171_ (.RESET_B(net787),
    .D(_00811_),
    .Q(\u_inv.d_next[74] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _49172_ (.RESET_B(net785),
    .D(_00812_),
    .Q(\u_inv.d_next[75] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _49173_ (.RESET_B(net783),
    .D(_00813_),
    .Q(\u_inv.d_next[76] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_2 _49174_ (.RESET_B(net782),
    .D(_00814_),
    .Q(\u_inv.d_next[77] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_2 _49175_ (.RESET_B(net780),
    .D(_00815_),
    .Q(\u_inv.d_next[78] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _49176_ (.RESET_B(net778),
    .D(_00816_),
    .Q(\u_inv.d_next[79] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _49177_ (.RESET_B(net776),
    .D(_00817_),
    .Q(\u_inv.d_next[80] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _49178_ (.RESET_B(net775),
    .D(_00818_),
    .Q(\u_inv.d_next[81] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _49179_ (.RESET_B(net773),
    .D(_00819_),
    .Q(\u_inv.d_next[82] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _49180_ (.RESET_B(net771),
    .D(_00820_),
    .Q(\u_inv.d_next[83] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _49181_ (.RESET_B(net769),
    .D(_00821_),
    .Q(\u_inv.d_next[84] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _49182_ (.RESET_B(net768),
    .D(_00822_),
    .Q(\u_inv.d_next[85] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _49183_ (.RESET_B(net766),
    .D(_00823_),
    .Q(\u_inv.d_next[86] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _49184_ (.RESET_B(net764),
    .D(_00824_),
    .Q(\u_inv.d_next[87] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _49185_ (.RESET_B(net762),
    .D(_00825_),
    .Q(\u_inv.d_next[88] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _49186_ (.RESET_B(net761),
    .D(_00826_),
    .Q(\u_inv.d_next[89] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _49187_ (.RESET_B(net759),
    .D(_00827_),
    .Q(\u_inv.d_next[90] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _49188_ (.RESET_B(net757),
    .D(_00828_),
    .Q(\u_inv.d_next[91] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _49189_ (.RESET_B(net755),
    .D(_00829_),
    .Q(\u_inv.d_next[92] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _49190_ (.RESET_B(net754),
    .D(_00830_),
    .Q(\u_inv.d_next[93] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _49191_ (.RESET_B(net752),
    .D(_00831_),
    .Q(\u_inv.d_next[94] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _49192_ (.RESET_B(net750),
    .D(_00832_),
    .Q(\u_inv.d_next[95] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _49193_ (.RESET_B(net748),
    .D(_00833_),
    .Q(\u_inv.d_next[96] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _49194_ (.RESET_B(net747),
    .D(_00834_),
    .Q(\u_inv.d_next[97] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _49195_ (.RESET_B(net745),
    .D(_00835_),
    .Q(\u_inv.d_next[98] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _49196_ (.RESET_B(net743),
    .D(_00836_),
    .Q(\u_inv.d_next[99] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _49197_ (.RESET_B(net741),
    .D(_00837_),
    .Q(\u_inv.d_next[100] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _49198_ (.RESET_B(net740),
    .D(_00838_),
    .Q(\u_inv.d_next[101] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _49199_ (.RESET_B(net738),
    .D(_00839_),
    .Q(\u_inv.d_next[102] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _49200_ (.RESET_B(net736),
    .D(_00840_),
    .Q(\u_inv.d_next[103] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _49201_ (.RESET_B(net734),
    .D(_00841_),
    .Q(\u_inv.d_next[104] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _49202_ (.RESET_B(net733),
    .D(_00842_),
    .Q(\u_inv.d_next[105] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _49203_ (.RESET_B(net731),
    .D(_00843_),
    .Q(\u_inv.d_next[106] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _49204_ (.RESET_B(net729),
    .D(_00844_),
    .Q(\u_inv.d_next[107] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _49205_ (.RESET_B(net727),
    .D(_00845_),
    .Q(\u_inv.d_next[108] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _49206_ (.RESET_B(net726),
    .D(_00846_),
    .Q(\u_inv.d_next[109] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _49207_ (.RESET_B(net724),
    .D(_00847_),
    .Q(\u_inv.d_next[110] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _49208_ (.RESET_B(net722),
    .D(_00848_),
    .Q(\u_inv.d_next[111] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _49209_ (.RESET_B(net720),
    .D(_00849_),
    .Q(\u_inv.d_next[112] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _49210_ (.RESET_B(net719),
    .D(_00850_),
    .Q(\u_inv.d_next[113] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _49211_ (.RESET_B(net717),
    .D(_00851_),
    .Q(\u_inv.d_next[114] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _49212_ (.RESET_B(net715),
    .D(_00852_),
    .Q(\u_inv.d_next[115] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _49213_ (.RESET_B(net713),
    .D(_00853_),
    .Q(\u_inv.d_next[116] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _49214_ (.RESET_B(net712),
    .D(_00854_),
    .Q(\u_inv.d_next[117] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _49215_ (.RESET_B(net710),
    .D(_00855_),
    .Q(\u_inv.d_next[118] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _49216_ (.RESET_B(net708),
    .D(_00856_),
    .Q(\u_inv.d_next[119] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _49217_ (.RESET_B(net706),
    .D(_00857_),
    .Q(\u_inv.d_next[120] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _49218_ (.RESET_B(net705),
    .D(_00858_),
    .Q(\u_inv.d_next[121] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _49219_ (.RESET_B(net703),
    .D(_00859_),
    .Q(\u_inv.d_next[122] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _49220_ (.RESET_B(net701),
    .D(_00860_),
    .Q(\u_inv.d_next[123] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _49221_ (.RESET_B(net699),
    .D(_00861_),
    .Q(\u_inv.d_next[124] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _49222_ (.RESET_B(net698),
    .D(_00862_),
    .Q(\u_inv.d_next[125] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _49223_ (.RESET_B(net696),
    .D(_00863_),
    .Q(\u_inv.d_next[126] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _49224_ (.RESET_B(net694),
    .D(_00864_),
    .Q(\u_inv.d_next[127] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _49225_ (.RESET_B(net692),
    .D(_00865_),
    .Q(\u_inv.d_next[128] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _49226_ (.RESET_B(net691),
    .D(_00866_),
    .Q(\u_inv.d_next[129] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _49227_ (.RESET_B(net689),
    .D(_00867_),
    .Q(\u_inv.d_next[130] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _49228_ (.RESET_B(net687),
    .D(_00868_),
    .Q(\u_inv.d_next[131] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _49229_ (.RESET_B(net685),
    .D(_00869_),
    .Q(\u_inv.d_next[132] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _49230_ (.RESET_B(net684),
    .D(_00870_),
    .Q(\u_inv.d_next[133] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _49231_ (.RESET_B(net682),
    .D(_00871_),
    .Q(\u_inv.d_next[134] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _49232_ (.RESET_B(net680),
    .D(_00872_),
    .Q(\u_inv.d_next[135] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _49233_ (.RESET_B(net678),
    .D(_00873_),
    .Q(\u_inv.d_next[136] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _49234_ (.RESET_B(net677),
    .D(_00874_),
    .Q(\u_inv.d_next[137] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _49235_ (.RESET_B(net675),
    .D(_00875_),
    .Q(\u_inv.d_next[138] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _49236_ (.RESET_B(net673),
    .D(_00876_),
    .Q(\u_inv.d_next[139] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _49237_ (.RESET_B(net671),
    .D(_00877_),
    .Q(\u_inv.d_next[140] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _49238_ (.RESET_B(net670),
    .D(_00878_),
    .Q(\u_inv.d_next[141] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _49239_ (.RESET_B(net668),
    .D(_00879_),
    .Q(\u_inv.d_next[142] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _49240_ (.RESET_B(net666),
    .D(_00880_),
    .Q(\u_inv.d_next[143] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _49241_ (.RESET_B(net664),
    .D(_00881_),
    .Q(\u_inv.d_next[144] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _49242_ (.RESET_B(net663),
    .D(_00882_),
    .Q(\u_inv.d_next[145] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _49243_ (.RESET_B(net661),
    .D(_00883_),
    .Q(\u_inv.d_next[146] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _49244_ (.RESET_B(net659),
    .D(_00884_),
    .Q(\u_inv.d_next[147] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _49245_ (.RESET_B(net657),
    .D(_00885_),
    .Q(\u_inv.d_next[148] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _49246_ (.RESET_B(net656),
    .D(_00886_),
    .Q(\u_inv.d_next[149] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _49247_ (.RESET_B(net654),
    .D(_00887_),
    .Q(\u_inv.d_next[150] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _49248_ (.RESET_B(net652),
    .D(_00888_),
    .Q(\u_inv.d_next[151] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _49249_ (.RESET_B(net650),
    .D(_00889_),
    .Q(\u_inv.d_next[152] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _49250_ (.RESET_B(net649),
    .D(_00890_),
    .Q(\u_inv.d_next[153] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _49251_ (.RESET_B(net647),
    .D(_00891_),
    .Q(\u_inv.d_next[154] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _49252_ (.RESET_B(net645),
    .D(_00892_),
    .Q(\u_inv.d_next[155] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _49253_ (.RESET_B(net643),
    .D(_00893_),
    .Q(\u_inv.d_next[156] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _49254_ (.RESET_B(net642),
    .D(_00894_),
    .Q(\u_inv.d_next[157] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _49255_ (.RESET_B(net640),
    .D(_00895_),
    .Q(\u_inv.d_next[158] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _49256_ (.RESET_B(net638),
    .D(_00896_),
    .Q(\u_inv.d_next[159] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _49257_ (.RESET_B(net636),
    .D(_00897_),
    .Q(\u_inv.d_next[160] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _49258_ (.RESET_B(net635),
    .D(_00898_),
    .Q(\u_inv.d_next[161] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _49259_ (.RESET_B(net633),
    .D(_00899_),
    .Q(\u_inv.d_next[162] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _49260_ (.RESET_B(net631),
    .D(_00900_),
    .Q(\u_inv.d_next[163] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _49261_ (.RESET_B(net629),
    .D(_00901_),
    .Q(\u_inv.d_next[164] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _49262_ (.RESET_B(net628),
    .D(_00902_),
    .Q(\u_inv.d_next[165] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _49263_ (.RESET_B(net626),
    .D(_00903_),
    .Q(\u_inv.d_next[166] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _49264_ (.RESET_B(net624),
    .D(_00904_),
    .Q(\u_inv.d_next[167] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _49265_ (.RESET_B(net622),
    .D(_00905_),
    .Q(\u_inv.d_next[168] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _49266_ (.RESET_B(net621),
    .D(_00906_),
    .Q(\u_inv.d_next[169] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _49267_ (.RESET_B(net619),
    .D(_00907_),
    .Q(\u_inv.d_next[170] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _49268_ (.RESET_B(net617),
    .D(_00908_),
    .Q(\u_inv.d_next[171] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _49269_ (.RESET_B(net615),
    .D(_00909_),
    .Q(\u_inv.d_next[172] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _49270_ (.RESET_B(net614),
    .D(_00910_),
    .Q(\u_inv.d_next[173] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _49271_ (.RESET_B(net612),
    .D(_00911_),
    .Q(\u_inv.d_next[174] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _49272_ (.RESET_B(net610),
    .D(_00912_),
    .Q(\u_inv.d_next[175] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _49273_ (.RESET_B(net608),
    .D(_00913_),
    .Q(\u_inv.d_next[176] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _49274_ (.RESET_B(net607),
    .D(_00914_),
    .Q(\u_inv.d_next[177] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _49275_ (.RESET_B(net605),
    .D(_00915_),
    .Q(\u_inv.d_next[178] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _49276_ (.RESET_B(net603),
    .D(_00916_),
    .Q(\u_inv.d_next[179] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _49277_ (.RESET_B(net601),
    .D(_00917_),
    .Q(\u_inv.d_next[180] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _49278_ (.RESET_B(net600),
    .D(_00918_),
    .Q(\u_inv.d_next[181] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _49279_ (.RESET_B(net598),
    .D(_00919_),
    .Q(\u_inv.d_next[182] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _49280_ (.RESET_B(net596),
    .D(_00920_),
    .Q(\u_inv.d_next[183] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _49281_ (.RESET_B(net594),
    .D(_00921_),
    .Q(\u_inv.d_next[184] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _49282_ (.RESET_B(net593),
    .D(_00922_),
    .Q(\u_inv.d_next[185] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _49283_ (.RESET_B(net591),
    .D(_00923_),
    .Q(\u_inv.d_next[186] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _49284_ (.RESET_B(net589),
    .D(_00924_),
    .Q(\u_inv.d_next[187] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _49285_ (.RESET_B(net587),
    .D(_00925_),
    .Q(\u_inv.d_next[188] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _49286_ (.RESET_B(net586),
    .D(_00926_),
    .Q(\u_inv.d_next[189] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_2 _49287_ (.RESET_B(net584),
    .D(_00927_),
    .Q(\u_inv.d_next[190] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _49288_ (.RESET_B(net582),
    .D(_00928_),
    .Q(\u_inv.d_next[191] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _49289_ (.RESET_B(net580),
    .D(_00929_),
    .Q(\u_inv.d_next[192] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _49290_ (.RESET_B(net579),
    .D(_00930_),
    .Q(\u_inv.d_next[193] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _49291_ (.RESET_B(net577),
    .D(_00931_),
    .Q(\u_inv.d_next[194] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _49292_ (.RESET_B(net575),
    .D(_00932_),
    .Q(\u_inv.d_next[195] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _49293_ (.RESET_B(net573),
    .D(_00933_),
    .Q(\u_inv.d_next[196] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _49294_ (.RESET_B(net572),
    .D(_00934_),
    .Q(\u_inv.d_next[197] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _49295_ (.RESET_B(net570),
    .D(_00935_),
    .Q(\u_inv.d_next[198] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _49296_ (.RESET_B(net568),
    .D(_00936_),
    .Q(\u_inv.d_next[199] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _49297_ (.RESET_B(net566),
    .D(_00937_),
    .Q(\u_inv.d_next[200] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _49298_ (.RESET_B(net565),
    .D(_00938_),
    .Q(\u_inv.d_next[201] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _49299_ (.RESET_B(net563),
    .D(_00939_),
    .Q(\u_inv.d_next[202] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _49300_ (.RESET_B(net561),
    .D(_00940_),
    .Q(\u_inv.d_next[203] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_2 _49301_ (.RESET_B(net559),
    .D(_00941_),
    .Q(\u_inv.d_next[204] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _49302_ (.RESET_B(net558),
    .D(_00942_),
    .Q(\u_inv.d_next[205] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_2 _49303_ (.RESET_B(net556),
    .D(_00943_),
    .Q(\u_inv.d_next[206] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _49304_ (.RESET_B(net554),
    .D(_00944_),
    .Q(\u_inv.d_next[207] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _49305_ (.RESET_B(net552),
    .D(_00945_),
    .Q(\u_inv.d_next[208] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _49306_ (.RESET_B(net551),
    .D(_00946_),
    .Q(\u_inv.d_next[209] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_2 _49307_ (.RESET_B(net549),
    .D(_00947_),
    .Q(\u_inv.d_next[210] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _49308_ (.RESET_B(net547),
    .D(_00948_),
    .Q(\u_inv.d_next[211] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _49309_ (.RESET_B(net545),
    .D(_00949_),
    .Q(\u_inv.d_next[212] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _49310_ (.RESET_B(net544),
    .D(_00950_),
    .Q(\u_inv.d_next[213] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _49311_ (.RESET_B(net542),
    .D(_00951_),
    .Q(\u_inv.d_next[214] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _49312_ (.RESET_B(net540),
    .D(_00952_),
    .Q(\u_inv.d_next[215] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_2 _49313_ (.RESET_B(net538),
    .D(_00953_),
    .Q(\u_inv.d_next[216] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _49314_ (.RESET_B(net537),
    .D(_00954_),
    .Q(\u_inv.d_next[217] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _49315_ (.RESET_B(net535),
    .D(_00955_),
    .Q(\u_inv.d_next[218] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _49316_ (.RESET_B(net533),
    .D(_00956_),
    .Q(\u_inv.d_next[219] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _49317_ (.RESET_B(net531),
    .D(_00957_),
    .Q(\u_inv.d_next[220] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _49318_ (.RESET_B(net530),
    .D(_00958_),
    .Q(\u_inv.d_next[221] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_2 _49319_ (.RESET_B(net528),
    .D(_00959_),
    .Q(\u_inv.d_next[222] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _49320_ (.RESET_B(net526),
    .D(_00960_),
    .Q(\u_inv.d_next[223] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _49321_ (.RESET_B(net524),
    .D(_00961_),
    .Q(\u_inv.d_next[224] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _49322_ (.RESET_B(net523),
    .D(_00962_),
    .Q(\u_inv.d_next[225] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _49323_ (.RESET_B(net521),
    .D(_00963_),
    .Q(\u_inv.d_next[226] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _49324_ (.RESET_B(net519),
    .D(_00964_),
    .Q(\u_inv.d_next[227] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _49325_ (.RESET_B(net517),
    .D(_00965_),
    .Q(\u_inv.d_next[228] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _49326_ (.RESET_B(net516),
    .D(_00966_),
    .Q(\u_inv.d_next[229] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _49327_ (.RESET_B(net514),
    .D(_00967_),
    .Q(\u_inv.d_next[230] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _49328_ (.RESET_B(net512),
    .D(_00968_),
    .Q(\u_inv.d_next[231] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _49329_ (.RESET_B(net510),
    .D(_00969_),
    .Q(\u_inv.d_next[232] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _49330_ (.RESET_B(net509),
    .D(_00970_),
    .Q(\u_inv.d_next[233] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _49331_ (.RESET_B(net507),
    .D(_00971_),
    .Q(\u_inv.d_next[234] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _49332_ (.RESET_B(net505),
    .D(_00972_),
    .Q(\u_inv.d_next[235] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _49333_ (.RESET_B(net503),
    .D(_00973_),
    .Q(\u_inv.d_next[236] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _49334_ (.RESET_B(net502),
    .D(_00974_),
    .Q(\u_inv.d_next[237] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _49335_ (.RESET_B(net500),
    .D(_00975_),
    .Q(\u_inv.d_next[238] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _49336_ (.RESET_B(net498),
    .D(_00976_),
    .Q(\u_inv.d_next[239] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _49337_ (.RESET_B(net496),
    .D(_00977_),
    .Q(\u_inv.d_next[240] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _49338_ (.RESET_B(net495),
    .D(_00978_),
    .Q(\u_inv.d_next[241] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _49339_ (.RESET_B(net493),
    .D(_00979_),
    .Q(\u_inv.d_next[242] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _49340_ (.RESET_B(net491),
    .D(_00980_),
    .Q(\u_inv.d_next[243] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _49341_ (.RESET_B(net489),
    .D(_00981_),
    .Q(\u_inv.d_next[244] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _49342_ (.RESET_B(net488),
    .D(_00982_),
    .Q(\u_inv.d_next[245] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _49343_ (.RESET_B(net486),
    .D(_00983_),
    .Q(\u_inv.d_next[246] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _49344_ (.RESET_B(net484),
    .D(_00984_),
    .Q(\u_inv.d_next[247] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _49345_ (.RESET_B(net482),
    .D(_00985_),
    .Q(\u_inv.d_next[248] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _49346_ (.RESET_B(net481),
    .D(_00986_),
    .Q(\u_inv.d_next[249] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _49347_ (.RESET_B(net479),
    .D(_00987_),
    .Q(\u_inv.d_next[250] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _49348_ (.RESET_B(net477),
    .D(_00988_),
    .Q(\u_inv.d_next[251] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _49349_ (.RESET_B(net475),
    .D(_00989_),
    .Q(\u_inv.d_next[252] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _49350_ (.RESET_B(net474),
    .D(_00990_),
    .Q(\u_inv.d_next[253] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _49351_ (.RESET_B(net472),
    .D(_00991_),
    .Q(\u_inv.d_next[254] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _49352_ (.RESET_B(net470),
    .D(_00992_),
    .Q(\u_inv.d_next[255] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _49353_ (.RESET_B(net468),
    .D(_00993_),
    .Q(\u_inv.d_next[256] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _49354_ (.RESET_B(net7475),
    .D(net3592),
    .Q(\inv_result[0] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _49355_ (.RESET_B(net7480),
    .D(net2180),
    .Q(\inv_result[1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _49356_ (.RESET_B(net7478),
    .D(net1489),
    .Q(\inv_result[2] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _49357_ (.RESET_B(net7478),
    .D(net2337),
    .Q(\inv_result[3] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _49358_ (.RESET_B(net7479),
    .D(net2470),
    .Q(\inv_result[4] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _49359_ (.RESET_B(net7478),
    .D(_00999_),
    .Q(\inv_result[5] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _49360_ (.RESET_B(net7479),
    .D(_01000_),
    .Q(\inv_result[6] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_2 _49361_ (.RESET_B(net7479),
    .D(_01001_),
    .Q(\inv_result[7] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _49362_ (.RESET_B(net7479),
    .D(_01002_),
    .Q(\inv_result[8] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _49363_ (.RESET_B(net7479),
    .D(_01003_),
    .Q(\inv_result[9] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_1 _49364_ (.RESET_B(net7483),
    .D(_01004_),
    .Q(\inv_result[10] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _49365_ (.RESET_B(net7483),
    .D(_01005_),
    .Q(\inv_result[11] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _49366_ (.RESET_B(net7483),
    .D(_01006_),
    .Q(\inv_result[12] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_1 _49367_ (.RESET_B(net7483),
    .D(_01007_),
    .Q(\inv_result[13] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_1 _49368_ (.RESET_B(net7483),
    .D(_01008_),
    .Q(\inv_result[14] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _49369_ (.RESET_B(net7484),
    .D(_01009_),
    .Q(\inv_result[15] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_1 _49370_ (.RESET_B(net7488),
    .D(_01010_),
    .Q(\inv_result[16] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_1 _49371_ (.RESET_B(net7489),
    .D(_01011_),
    .Q(\inv_result[17] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_2 _49372_ (.RESET_B(net7489),
    .D(_01012_),
    .Q(\inv_result[18] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _49373_ (.RESET_B(net7490),
    .D(_01013_),
    .Q(\inv_result[19] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _49374_ (.RESET_B(net7488),
    .D(_01014_),
    .Q(\inv_result[20] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _49375_ (.RESET_B(net7490),
    .D(_01015_),
    .Q(\inv_result[21] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _49376_ (.RESET_B(net7489),
    .D(_01016_),
    .Q(\inv_result[22] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _49377_ (.RESET_B(net7488),
    .D(_01017_),
    .Q(\inv_result[23] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _49378_ (.RESET_B(net7489),
    .D(_01018_),
    .Q(\inv_result[24] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _49379_ (.RESET_B(net7488),
    .D(_01019_),
    .Q(\inv_result[25] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _49380_ (.RESET_B(net7495),
    .D(_01020_),
    .Q(\inv_result[26] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_1 _49381_ (.RESET_B(net7495),
    .D(_01021_),
    .Q(\inv_result[27] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_1 _49382_ (.RESET_B(net7496),
    .D(_01022_),
    .Q(\inv_result[28] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_1 _49383_ (.RESET_B(net7496),
    .D(_01023_),
    .Q(\inv_result[29] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_1 _49384_ (.RESET_B(net7496),
    .D(_01024_),
    .Q(\inv_result[30] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_1 _49385_ (.RESET_B(net7496),
    .D(_01025_),
    .Q(\inv_result[31] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _49386_ (.RESET_B(net7499),
    .D(_01026_),
    .Q(\inv_result[32] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _49387_ (.RESET_B(net7515),
    .D(_01027_),
    .Q(\inv_result[33] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _49388_ (.RESET_B(net7515),
    .D(_01028_),
    .Q(\inv_result[34] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _49389_ (.RESET_B(net7512),
    .D(_01029_),
    .Q(\inv_result[35] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _49390_ (.RESET_B(net7515),
    .D(_01030_),
    .Q(\inv_result[36] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _49391_ (.RESET_B(net7516),
    .D(_01031_),
    .Q(\inv_result[37] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _49392_ (.RESET_B(net7512),
    .D(_01032_),
    .Q(\inv_result[38] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _49393_ (.RESET_B(net7512),
    .D(_01033_),
    .Q(\inv_result[39] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_1 _49394_ (.RESET_B(net7513),
    .D(_01034_),
    .Q(\inv_result[40] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_1 _49395_ (.RESET_B(net7512),
    .D(_01035_),
    .Q(\inv_result[41] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_1 _49396_ (.RESET_B(net7514),
    .D(_01036_),
    .Q(\inv_result[42] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _49397_ (.RESET_B(net7513),
    .D(_01037_),
    .Q(\inv_result[43] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _49398_ (.RESET_B(net7514),
    .D(_01038_),
    .Q(\inv_result[44] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_1 _49399_ (.RESET_B(net7514),
    .D(_01039_),
    .Q(\inv_result[45] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_1 _49400_ (.RESET_B(net7518),
    .D(_01040_),
    .Q(\inv_result[46] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_1 _49401_ (.RESET_B(net7514),
    .D(_01041_),
    .Q(\inv_result[47] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _49402_ (.RESET_B(net7514),
    .D(_01042_),
    .Q(\inv_result[48] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _49403_ (.RESET_B(net7516),
    .D(_01043_),
    .Q(\inv_result[49] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _49404_ (.RESET_B(net7519),
    .D(_01044_),
    .Q(\inv_result[50] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _49405_ (.RESET_B(net7518),
    .D(_01045_),
    .Q(\inv_result[51] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _49406_ (.RESET_B(net7519),
    .D(_01046_),
    .Q(\inv_result[52] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_2 _49407_ (.RESET_B(net7519),
    .D(_01047_),
    .Q(\inv_result[53] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_2 _49408_ (.RESET_B(net7529),
    .D(_01048_),
    .Q(\inv_result[54] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_2 _49409_ (.RESET_B(net7529),
    .D(_01049_),
    .Q(\inv_result[55] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_2 _49410_ (.RESET_B(net7526),
    .D(_01050_),
    .Q(\inv_result[56] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _49411_ (.RESET_B(net7529),
    .D(_01051_),
    .Q(\inv_result[57] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_2 _49412_ (.RESET_B(net7520),
    .D(_01052_),
    .Q(\inv_result[58] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_2 _49413_ (.RESET_B(net7529),
    .D(_01053_),
    .Q(\inv_result[59] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_2 _49414_ (.RESET_B(net7529),
    .D(_01054_),
    .Q(\inv_result[60] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_2 _49415_ (.RESET_B(net7529),
    .D(_01055_),
    .Q(\inv_result[61] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _49416_ (.RESET_B(net7529),
    .D(_01056_),
    .Q(\inv_result[62] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _49417_ (.RESET_B(net7530),
    .D(_01057_),
    .Q(\inv_result[63] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _49418_ (.RESET_B(net7536),
    .D(_01058_),
    .Q(\inv_result[64] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_2 _49419_ (.RESET_B(net7550),
    .D(_01059_),
    .Q(\inv_result[65] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_2 _49420_ (.RESET_B(net7551),
    .D(_01060_),
    .Q(\inv_result[66] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_2 _49421_ (.RESET_B(net7551),
    .D(_01061_),
    .Q(\inv_result[67] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_2 _49422_ (.RESET_B(net7556),
    .D(_01062_),
    .Q(\inv_result[68] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_2 _49423_ (.RESET_B(net7555),
    .D(_01063_),
    .Q(\inv_result[69] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_2 _49424_ (.RESET_B(net7551),
    .D(_01064_),
    .Q(\inv_result[70] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_2 _49425_ (.RESET_B(net7563),
    .D(_01065_),
    .Q(\inv_result[71] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_2 _49426_ (.RESET_B(net7558),
    .D(_01066_),
    .Q(\inv_result[72] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_2 _49427_ (.RESET_B(net7556),
    .D(_01067_),
    .Q(\inv_result[73] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_2 _49428_ (.RESET_B(net7563),
    .D(_01068_),
    .Q(\inv_result[74] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_2 _49429_ (.RESET_B(net7563),
    .D(_01069_),
    .Q(\inv_result[75] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_2 _49430_ (.RESET_B(net7563),
    .D(_01070_),
    .Q(\inv_result[76] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_2 _49431_ (.RESET_B(net7551),
    .D(_01071_),
    .Q(\inv_result[77] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_2 _49432_ (.RESET_B(net7564),
    .D(_01072_),
    .Q(\inv_result[78] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_2 _49433_ (.RESET_B(net7563),
    .D(_01073_),
    .Q(\inv_result[79] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_2 _49434_ (.RESET_B(net7563),
    .D(_01074_),
    .Q(\inv_result[80] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_2 _49435_ (.RESET_B(net7555),
    .D(_01075_),
    .Q(\inv_result[81] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _49436_ (.RESET_B(net7555),
    .D(_01076_),
    .Q(\inv_result[82] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_2 _49437_ (.RESET_B(net7555),
    .D(_01077_),
    .Q(\inv_result[83] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_2 _49438_ (.RESET_B(net7553),
    .D(_01078_),
    .Q(\inv_result[84] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_2 _49439_ (.RESET_B(net7553),
    .D(_01079_),
    .Q(\inv_result[85] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _49440_ (.RESET_B(net7553),
    .D(_01080_),
    .Q(\inv_result[86] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_2 _49441_ (.RESET_B(net7554),
    .D(_01081_),
    .Q(\inv_result[87] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_2 _49442_ (.RESET_B(net7553),
    .D(_01082_),
    .Q(\inv_result[88] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_2 _49443_ (.RESET_B(net7554),
    .D(_01083_),
    .Q(\inv_result[89] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_2 _49444_ (.RESET_B(net7554),
    .D(_01084_),
    .Q(\inv_result[90] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _49445_ (.RESET_B(net7536),
    .D(_01085_),
    .Q(\inv_result[91] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_2 _49446_ (.RESET_B(net7554),
    .D(_01086_),
    .Q(\inv_result[92] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _49447_ (.RESET_B(net7536),
    .D(_01087_),
    .Q(\inv_result[93] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_2 _49448_ (.RESET_B(net7553),
    .D(_01088_),
    .Q(\inv_result[94] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _49449_ (.RESET_B(net7553),
    .D(_01089_),
    .Q(\inv_result[95] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _49450_ (.RESET_B(net7534),
    .D(_01090_),
    .Q(\inv_result[96] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _49451_ (.RESET_B(net7545),
    .D(_01091_),
    .Q(\inv_result[97] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _49452_ (.RESET_B(net7545),
    .D(_01092_),
    .Q(\inv_result[98] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _49453_ (.RESET_B(net7534),
    .D(_01093_),
    .Q(\inv_result[99] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _49454_ (.RESET_B(net7546),
    .D(_01094_),
    .Q(\inv_result[100] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _49455_ (.RESET_B(net7546),
    .D(_01095_),
    .Q(\inv_result[101] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _49456_ (.RESET_B(net7548),
    .D(_01096_),
    .Q(\inv_result[102] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _49457_ (.RESET_B(net7546),
    .D(_01097_),
    .Q(\inv_result[103] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _49458_ (.RESET_B(net7547),
    .D(_01098_),
    .Q(\inv_result[104] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_1 _49459_ (.RESET_B(net7546),
    .D(_01099_),
    .Q(\inv_result[105] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _49460_ (.RESET_B(net7540),
    .D(_01100_),
    .Q(\inv_result[106] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_2 _49461_ (.RESET_B(net7545),
    .D(_01101_),
    .Q(\inv_result[107] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _49462_ (.RESET_B(net7547),
    .D(_01102_),
    .Q(\inv_result[108] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _49463_ (.RESET_B(net7545),
    .D(_01103_),
    .Q(\inv_result[109] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _49464_ (.RESET_B(net7547),
    .D(_01104_),
    .Q(\inv_result[110] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_2 _49465_ (.RESET_B(net7547),
    .D(_01105_),
    .Q(\inv_result[111] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _49466_ (.RESET_B(net7549),
    .D(_01106_),
    .Q(\inv_result[112] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _49467_ (.RESET_B(net7547),
    .D(_01107_),
    .Q(\inv_result[113] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _49468_ (.RESET_B(net7547),
    .D(_01108_),
    .Q(\inv_result[114] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _49469_ (.RESET_B(net7541),
    .D(_01109_),
    .Q(\inv_result[115] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _49470_ (.RESET_B(net7542),
    .D(_01110_),
    .Q(\inv_result[116] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _49471_ (.RESET_B(net7543),
    .D(_01111_),
    .Q(\inv_result[117] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _49472_ (.RESET_B(net7538),
    .D(_01112_),
    .Q(\inv_result[118] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _49473_ (.RESET_B(net7538),
    .D(_01113_),
    .Q(\inv_result[119] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_1 _49474_ (.RESET_B(net7543),
    .D(_01114_),
    .Q(\inv_result[120] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _49475_ (.RESET_B(net7538),
    .D(_01115_),
    .Q(\inv_result[121] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _49476_ (.RESET_B(net7541),
    .D(_01116_),
    .Q(\inv_result[122] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _49477_ (.RESET_B(net7538),
    .D(_01117_),
    .Q(\inv_result[123] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_1 _49478_ (.RESET_B(net7542),
    .D(_01118_),
    .Q(\inv_result[124] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _49479_ (.RESET_B(net7543),
    .D(_01119_),
    .Q(\inv_result[125] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _49480_ (.RESET_B(net7543),
    .D(_01120_),
    .Q(\inv_result[126] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _49481_ (.RESET_B(net7538),
    .D(_01121_),
    .Q(\inv_result[127] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _49482_ (.RESET_B(net7523),
    .D(_01122_),
    .Q(\inv_result[128] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _49483_ (.RESET_B(net7523),
    .D(_01123_),
    .Q(\inv_result[129] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _49484_ (.RESET_B(net7521),
    .D(_01124_),
    .Q(\inv_result[130] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _49485_ (.RESET_B(net7524),
    .D(_01125_),
    .Q(\inv_result[131] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _49486_ (.RESET_B(net7522),
    .D(_01126_),
    .Q(\inv_result[132] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _49487_ (.RESET_B(net7522),
    .D(_01127_),
    .Q(\inv_result[133] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_1 _49488_ (.RESET_B(net7524),
    .D(_01128_),
    .Q(\inv_result[134] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _49489_ (.RESET_B(net7521),
    .D(_01129_),
    .Q(\inv_result[135] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _49490_ (.RESET_B(net7521),
    .D(_01130_),
    .Q(\inv_result[136] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _49491_ (.RESET_B(net7521),
    .D(_01131_),
    .Q(\inv_result[137] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_1 _49492_ (.RESET_B(net7521),
    .D(_01132_),
    .Q(\inv_result[138] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _49493_ (.RESET_B(net7510),
    .D(_01133_),
    .Q(\inv_result[139] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _49494_ (.RESET_B(net7510),
    .D(_01134_),
    .Q(\inv_result[140] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _49495_ (.RESET_B(net7510),
    .D(_01135_),
    .Q(\inv_result[141] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _49496_ (.RESET_B(net7510),
    .D(_01136_),
    .Q(\inv_result[142] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _49497_ (.RESET_B(net7508),
    .D(_01137_),
    .Q(\inv_result[143] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _49498_ (.RESET_B(net7508),
    .D(_01138_),
    .Q(\inv_result[144] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _49499_ (.RESET_B(net7508),
    .D(_01139_),
    .Q(\inv_result[145] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _49500_ (.RESET_B(net7508),
    .D(_01140_),
    .Q(\inv_result[146] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _49501_ (.RESET_B(net7508),
    .D(_01141_),
    .Q(\inv_result[147] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _49502_ (.RESET_B(net7506),
    .D(_01142_),
    .Q(\inv_result[148] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _49503_ (.RESET_B(net7506),
    .D(_01143_),
    .Q(\inv_result[149] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _49504_ (.RESET_B(net7507),
    .D(_01144_),
    .Q(\inv_result[150] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _49505_ (.RESET_B(net7504),
    .D(_01145_),
    .Q(\inv_result[151] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _49506_ (.RESET_B(net7504),
    .D(_01146_),
    .Q(\inv_result[152] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _49507_ (.RESET_B(net7502),
    .D(_01147_),
    .Q(\inv_result[153] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _49508_ (.RESET_B(net7505),
    .D(_01148_),
    .Q(\inv_result[154] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _49509_ (.RESET_B(net7504),
    .D(_01149_),
    .Q(\inv_result[155] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _49510_ (.RESET_B(net7504),
    .D(_01150_),
    .Q(\inv_result[156] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _49511_ (.RESET_B(net7504),
    .D(_01151_),
    .Q(\inv_result[157] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _49512_ (.RESET_B(net7504),
    .D(_01152_),
    .Q(\inv_result[158] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _49513_ (.RESET_B(net7504),
    .D(_01153_),
    .Q(\inv_result[159] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _49514_ (.RESET_B(net7503),
    .D(_01154_),
    .Q(\inv_result[160] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _49515_ (.RESET_B(net7502),
    .D(_01155_),
    .Q(\inv_result[161] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _49516_ (.RESET_B(net7502),
    .D(_01156_),
    .Q(\inv_result[162] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _49517_ (.RESET_B(net7502),
    .D(_01157_),
    .Q(\inv_result[163] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _49518_ (.RESET_B(net7493),
    .D(_01158_),
    .Q(\inv_result[164] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _49519_ (.RESET_B(net7493),
    .D(_01159_),
    .Q(\inv_result[165] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _49520_ (.RESET_B(net7493),
    .D(_01160_),
    .Q(\inv_result[166] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _49521_ (.RESET_B(net7493),
    .D(_01161_),
    .Q(\inv_result[167] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _49522_ (.RESET_B(net7491),
    .D(_01162_),
    .Q(\inv_result[168] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _49523_ (.RESET_B(net7487),
    .D(_01163_),
    .Q(\inv_result[169] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _49524_ (.RESET_B(net7487),
    .D(_01164_),
    .Q(\inv_result[170] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _49525_ (.RESET_B(net7487),
    .D(_01165_),
    .Q(\inv_result[171] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _49526_ (.RESET_B(net7486),
    .D(_01166_),
    .Q(\inv_result[172] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _49527_ (.RESET_B(net7487),
    .D(_01167_),
    .Q(\inv_result[173] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _49528_ (.RESET_B(net7486),
    .D(_01168_),
    .Q(\inv_result[174] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _49529_ (.RESET_B(net7486),
    .D(_01169_),
    .Q(\inv_result[175] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _49530_ (.RESET_B(net7480),
    .D(_01170_),
    .Q(\inv_result[176] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _49531_ (.RESET_B(net7480),
    .D(_01171_),
    .Q(\inv_result[177] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _49532_ (.RESET_B(net7476),
    .D(_01172_),
    .Q(\inv_result[178] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _49533_ (.RESET_B(net7486),
    .D(_01173_),
    .Q(\inv_result[179] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _49534_ (.RESET_B(net7480),
    .D(_01174_),
    .Q(\inv_result[180] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _49535_ (.RESET_B(net7486),
    .D(_01175_),
    .Q(\inv_result[181] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _49536_ (.RESET_B(net7481),
    .D(_01176_),
    .Q(\inv_result[182] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _49537_ (.RESET_B(net7486),
    .D(_01177_),
    .Q(\inv_result[183] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _49538_ (.RESET_B(net7481),
    .D(_01178_),
    .Q(\inv_result[184] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _49539_ (.RESET_B(net7480),
    .D(_01179_),
    .Q(\inv_result[185] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _49540_ (.RESET_B(net7480),
    .D(_01180_),
    .Q(\inv_result[186] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _49541_ (.RESET_B(net7474),
    .D(net1229),
    .Q(\inv_result[187] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _49542_ (.RESET_B(net7480),
    .D(_01182_),
    .Q(\inv_result[188] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _49543_ (.RESET_B(net7476),
    .D(_01183_),
    .Q(\inv_result[189] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _49544_ (.RESET_B(net7476),
    .D(_01184_),
    .Q(\inv_result[190] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _49545_ (.RESET_B(net7480),
    .D(_01185_),
    .Q(\inv_result[191] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _49546_ (.RESET_B(net7468),
    .D(_01186_),
    .Q(\inv_result[192] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _49547_ (.RESET_B(net7474),
    .D(_01187_),
    .Q(\inv_result[193] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _49548_ (.RESET_B(net7476),
    .D(_01188_),
    .Q(\inv_result[194] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _49549_ (.RESET_B(net7476),
    .D(_01189_),
    .Q(\inv_result[195] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _49550_ (.RESET_B(net7468),
    .D(_01190_),
    .Q(\inv_result[196] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _49551_ (.RESET_B(net7465),
    .D(_01191_),
    .Q(\inv_result[197] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _49552_ (.RESET_B(net7467),
    .D(_01192_),
    .Q(\inv_result[198] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _49553_ (.RESET_B(net7472),
    .D(net2014),
    .Q(\inv_result[199] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _49554_ (.RESET_B(net7472),
    .D(_01194_),
    .Q(\inv_result[200] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _49555_ (.RESET_B(net7472),
    .D(_01195_),
    .Q(\inv_result[201] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _49556_ (.RESET_B(net7467),
    .D(_01196_),
    .Q(\inv_result[202] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _49557_ (.RESET_B(net7468),
    .D(_01197_),
    .Q(\inv_result[203] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _49558_ (.RESET_B(net7467),
    .D(_01198_),
    .Q(\inv_result[204] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _49559_ (.RESET_B(net7466),
    .D(_01199_),
    .Q(\inv_result[205] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _49560_ (.RESET_B(net7466),
    .D(_01200_),
    .Q(\inv_result[206] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _49561_ (.RESET_B(net7466),
    .D(_01201_),
    .Q(\inv_result[207] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _49562_ (.RESET_B(net7466),
    .D(_01202_),
    .Q(\inv_result[208] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _49563_ (.RESET_B(net7465),
    .D(_01203_),
    .Q(\inv_result[209] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _49564_ (.RESET_B(net7461),
    .D(_01204_),
    .Q(\inv_result[210] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _49565_ (.RESET_B(net7467),
    .D(_01205_),
    .Q(\inv_result[211] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _49566_ (.RESET_B(net7467),
    .D(_01206_),
    .Q(\inv_result[212] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _49567_ (.RESET_B(net7465),
    .D(_01207_),
    .Q(\inv_result[213] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _49568_ (.RESET_B(net7467),
    .D(_01208_),
    .Q(\inv_result[214] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _49569_ (.RESET_B(net7467),
    .D(_01209_),
    .Q(\inv_result[215] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _49570_ (.RESET_B(net7460),
    .D(_01210_),
    .Q(\inv_result[216] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _49571_ (.RESET_B(net7459),
    .D(_01211_),
    .Q(\inv_result[217] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _49572_ (.RESET_B(net7460),
    .D(_01212_),
    .Q(\inv_result[218] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _49573_ (.RESET_B(net7460),
    .D(_01213_),
    .Q(\inv_result[219] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _49574_ (.RESET_B(net7460),
    .D(_01214_),
    .Q(\inv_result[220] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _49575_ (.RESET_B(net7427),
    .D(_01215_),
    .Q(\inv_result[221] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _49576_ (.RESET_B(net7427),
    .D(_01216_),
    .Q(\inv_result[222] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _49577_ (.RESET_B(net7428),
    .D(_01217_),
    .Q(\inv_result[223] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _49578_ (.RESET_B(net7446),
    .D(_01218_),
    .Q(\inv_result[224] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _49579_ (.RESET_B(net7446),
    .D(_01219_),
    .Q(\inv_result[225] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _49580_ (.RESET_B(net7427),
    .D(_01220_),
    .Q(\inv_result[226] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _49581_ (.RESET_B(net7427),
    .D(_01221_),
    .Q(\inv_result[227] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _49582_ (.RESET_B(net7427),
    .D(_01222_),
    .Q(\inv_result[228] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _49583_ (.RESET_B(net7427),
    .D(_01223_),
    .Q(\inv_result[229] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _49584_ (.RESET_B(net7428),
    .D(_01224_),
    .Q(\inv_result[230] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _49585_ (.RESET_B(net7446),
    .D(_01225_),
    .Q(\inv_result[231] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _49586_ (.RESET_B(net7470),
    .D(_01226_),
    .Q(\inv_result[232] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _49587_ (.RESET_B(net7442),
    .D(_01227_),
    .Q(\inv_result[233] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _49588_ (.RESET_B(net7446),
    .D(_01228_),
    .Q(\inv_result[234] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _49589_ (.RESET_B(net7442),
    .D(_01229_),
    .Q(\inv_result[235] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _49590_ (.RESET_B(net7446),
    .D(_01230_),
    .Q(\inv_result[236] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _49591_ (.RESET_B(net7442),
    .D(_01231_),
    .Q(\inv_result[237] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _49592_ (.RESET_B(net7446),
    .D(_01232_),
    .Q(\inv_result[238] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _49593_ (.RESET_B(net7446),
    .D(_01233_),
    .Q(\inv_result[239] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _49594_ (.RESET_B(net7445),
    .D(_01234_),
    .Q(\inv_result[240] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _49595_ (.RESET_B(net7443),
    .D(_01235_),
    .Q(\inv_result[241] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _49596_ (.RESET_B(net7447),
    .D(_01236_),
    .Q(\inv_result[242] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _49597_ (.RESET_B(net7470),
    .D(_01237_),
    .Q(\inv_result[243] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _49598_ (.RESET_B(net7470),
    .D(_01238_),
    .Q(\inv_result[244] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _49599_ (.RESET_B(net7443),
    .D(_01239_),
    .Q(\inv_result[245] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _49600_ (.RESET_B(net7445),
    .D(_01240_),
    .Q(\inv_result[246] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _49601_ (.RESET_B(net7445),
    .D(_01241_),
    .Q(\inv_result[247] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _49602_ (.RESET_B(net7444),
    .D(_01242_),
    .Q(\inv_result[248] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _49603_ (.RESET_B(net7445),
    .D(_01243_),
    .Q(\inv_result[249] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _49604_ (.RESET_B(net7445),
    .D(_01244_),
    .Q(\inv_result[250] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _49605_ (.RESET_B(net7445),
    .D(_01245_),
    .Q(\inv_result[251] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _49606_ (.RESET_B(net7445),
    .D(_01246_),
    .Q(\inv_result[252] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _49607_ (.RESET_B(net7445),
    .D(_01247_),
    .Q(\inv_result[253] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _49608_ (.RESET_B(net7453),
    .D(_01248_),
    .Q(\inv_result[254] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _49609_ (.RESET_B(net7453),
    .D(_01249_),
    .Q(\inv_result[255] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _49610_ (.RESET_B(net467),
    .D(net2704),
    .Q(\u_inv.d_reg[0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _49611_ (.RESET_B(net465),
    .D(_01251_),
    .Q(\u_inv.d_reg[1] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _49612_ (.RESET_B(net463),
    .D(net2515),
    .Q(\u_inv.d_reg[2] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _49613_ (.RESET_B(net461),
    .D(net2975),
    .Q(\u_inv.d_reg[3] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _49614_ (.RESET_B(net460),
    .D(net2820),
    .Q(\u_inv.d_reg[4] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _49615_ (.RESET_B(net458),
    .D(net2465),
    .Q(\u_inv.d_reg[5] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _49616_ (.RESET_B(net456),
    .D(net2806),
    .Q(\u_inv.d_reg[6] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _49617_ (.RESET_B(net454),
    .D(net2737),
    .Q(\u_inv.d_reg[7] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _49618_ (.RESET_B(net453),
    .D(net1824),
    .Q(\u_inv.d_reg[8] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _49619_ (.RESET_B(net451),
    .D(net3146),
    .Q(\u_inv.d_reg[9] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_1 _49620_ (.RESET_B(net449),
    .D(net2978),
    .Q(\u_inv.d_reg[10] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _49621_ (.RESET_B(net447),
    .D(net1390),
    .Q(\u_inv.d_reg[11] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _49622_ (.RESET_B(net446),
    .D(net2808),
    .Q(\u_inv.d_reg[12] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _49623_ (.RESET_B(net444),
    .D(_01263_),
    .Q(\u_inv.d_reg[13] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _49624_ (.RESET_B(net442),
    .D(net2946),
    .Q(\u_inv.d_reg[14] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _49625_ (.RESET_B(net440),
    .D(net2798),
    .Q(\u_inv.d_reg[15] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _49626_ (.RESET_B(net439),
    .D(net3079),
    .Q(\u_inv.d_reg[16] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _49627_ (.RESET_B(net437),
    .D(_01267_),
    .Q(\u_inv.d_reg[17] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _49628_ (.RESET_B(net435),
    .D(_01268_),
    .Q(\u_inv.d_reg[18] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _49629_ (.RESET_B(net433),
    .D(net3384),
    .Q(\u_inv.d_reg[19] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _49630_ (.RESET_B(net432),
    .D(net3294),
    .Q(\u_inv.d_reg[20] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _49631_ (.RESET_B(net430),
    .D(net3081),
    .Q(\u_inv.d_reg[21] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _49632_ (.RESET_B(net428),
    .D(net3211),
    .Q(\u_inv.d_reg[22] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _49633_ (.RESET_B(net426),
    .D(net3143),
    .Q(\u_inv.d_reg[23] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _49634_ (.RESET_B(net425),
    .D(_01274_),
    .Q(\u_inv.d_reg[24] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _49635_ (.RESET_B(net423),
    .D(net2949),
    .Q(\u_inv.d_reg[25] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _49636_ (.RESET_B(net421),
    .D(net3134),
    .Q(\u_inv.d_reg[26] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _49637_ (.RESET_B(net419),
    .D(net2039),
    .Q(\u_inv.d_reg[27] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _49638_ (.RESET_B(net418),
    .D(net2269),
    .Q(\u_inv.d_reg[28] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _49639_ (.RESET_B(net416),
    .D(net1916),
    .Q(\u_inv.d_reg[29] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _49640_ (.RESET_B(net414),
    .D(net3472),
    .Q(\u_inv.d_reg[30] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _49641_ (.RESET_B(net412),
    .D(net1743),
    .Q(\u_inv.d_reg[31] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _49642_ (.RESET_B(net411),
    .D(net2101),
    .Q(\u_inv.d_reg[32] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _49643_ (.RESET_B(net409),
    .D(net3097),
    .Q(\u_inv.d_reg[33] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _49644_ (.RESET_B(net407),
    .D(net1956),
    .Q(\u_inv.d_reg[34] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _49645_ (.RESET_B(net405),
    .D(net2647),
    .Q(\u_inv.d_reg[35] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _49646_ (.RESET_B(net404),
    .D(net2706),
    .Q(\u_inv.d_reg[36] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _49647_ (.RESET_B(net402),
    .D(net2765),
    .Q(\u_inv.d_reg[37] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _49648_ (.RESET_B(net400),
    .D(net2763),
    .Q(\u_inv.d_reg[38] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _49649_ (.RESET_B(net398),
    .D(net3164),
    .Q(\u_inv.d_reg[39] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _49650_ (.RESET_B(net397),
    .D(net3324),
    .Q(\u_inv.d_reg[40] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_2 _49651_ (.RESET_B(net395),
    .D(net3417),
    .Q(\u_inv.d_reg[41] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _49652_ (.RESET_B(net393),
    .D(net1725),
    .Q(\u_inv.d_reg[42] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_2 _49653_ (.RESET_B(net391),
    .D(net3012),
    .Q(\u_inv.d_reg[43] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_2 _49654_ (.RESET_B(net390),
    .D(net3125),
    .Q(\u_inv.d_reg[44] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _49655_ (.RESET_B(net388),
    .D(net3354),
    .Q(\u_inv.d_reg[45] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _49656_ (.RESET_B(net386),
    .D(_01296_),
    .Q(\u_inv.d_reg[46] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _49657_ (.RESET_B(net384),
    .D(net3046),
    .Q(\u_inv.d_reg[47] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _49658_ (.RESET_B(net383),
    .D(net2481),
    .Q(\u_inv.d_reg[48] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _49659_ (.RESET_B(net381),
    .D(_01299_),
    .Q(\u_inv.d_reg[49] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _49660_ (.RESET_B(net379),
    .D(net1239),
    .Q(\u_inv.d_reg[50] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _49661_ (.RESET_B(net377),
    .D(net3580),
    .Q(\u_inv.d_reg[51] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _49662_ (.RESET_B(net376),
    .D(_01302_),
    .Q(\u_inv.d_reg[52] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_2 _49663_ (.RESET_B(net374),
    .D(net3237),
    .Q(\u_inv.d_reg[53] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_2 _49664_ (.RESET_B(net372),
    .D(net2911),
    .Q(\u_inv.d_reg[54] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_2 _49665_ (.RESET_B(net370),
    .D(_01305_),
    .Q(\u_inv.d_reg[55] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_2 _49666_ (.RESET_B(net369),
    .D(net3584),
    .Q(\u_inv.d_reg[56] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_2 _49667_ (.RESET_B(net367),
    .D(net2444),
    .Q(\u_inv.d_reg[57] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_2 _49668_ (.RESET_B(net365),
    .D(net2615),
    .Q(\u_inv.d_reg[58] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _49669_ (.RESET_B(net363),
    .D(_01309_),
    .Q(\u_inv.d_reg[59] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _49670_ (.RESET_B(net362),
    .D(net2121),
    .Q(\u_inv.d_reg[60] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _49671_ (.RESET_B(net360),
    .D(net3075),
    .Q(\u_inv.d_reg[61] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _49672_ (.RESET_B(net358),
    .D(_01312_),
    .Q(\u_inv.d_reg[62] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _49673_ (.RESET_B(net356),
    .D(net3010),
    .Q(\u_inv.d_reg[63] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _49674_ (.RESET_B(net355),
    .D(net2254),
    .Q(\u_inv.d_reg[64] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _49675_ (.RESET_B(net353),
    .D(net2815),
    .Q(\u_inv.d_reg[65] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _49676_ (.RESET_B(net351),
    .D(net2522),
    .Q(\u_inv.d_reg[66] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _49677_ (.RESET_B(net349),
    .D(net3200),
    .Q(\u_inv.d_reg[67] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _49678_ (.RESET_B(net348),
    .D(net3341),
    .Q(\u_inv.d_reg[68] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _49679_ (.RESET_B(net346),
    .D(net3240),
    .Q(\u_inv.d_reg[69] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _49680_ (.RESET_B(net344),
    .D(_01320_),
    .Q(\u_inv.d_reg[70] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _49681_ (.RESET_B(net342),
    .D(_01321_),
    .Q(\u_inv.d_reg[71] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_2 _49682_ (.RESET_B(net341),
    .D(net3524),
    .Q(\u_inv.d_reg[72] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_2 _49683_ (.RESET_B(net339),
    .D(_01323_),
    .Q(\u_inv.d_reg[73] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _49684_ (.RESET_B(net337),
    .D(net3478),
    .Q(\u_inv.d_reg[74] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _49685_ (.RESET_B(net335),
    .D(net3394),
    .Q(\u_inv.d_reg[75] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _49686_ (.RESET_B(net334),
    .D(net2586),
    .Q(\u_inv.d_reg[76] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _49687_ (.RESET_B(net332),
    .D(net1850),
    .Q(\u_inv.d_reg[77] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _49688_ (.RESET_B(net330),
    .D(net3275),
    .Q(\u_inv.d_reg[78] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _49689_ (.RESET_B(net328),
    .D(net2326),
    .Q(\u_inv.d_reg[79] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _49690_ (.RESET_B(net327),
    .D(net2367),
    .Q(\u_inv.d_reg[80] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _49691_ (.RESET_B(net325),
    .D(net2732),
    .Q(\u_inv.d_reg[81] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _49692_ (.RESET_B(net323),
    .D(net2747),
    .Q(\u_inv.d_reg[82] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _49693_ (.RESET_B(net321),
    .D(net3463),
    .Q(\u_inv.d_reg[83] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _49694_ (.RESET_B(net320),
    .D(net3335),
    .Q(\u_inv.d_reg[84] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _49695_ (.RESET_B(net318),
    .D(_01335_),
    .Q(\u_inv.d_reg[85] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _49696_ (.RESET_B(net316),
    .D(net3511),
    .Q(\u_inv.d_reg[86] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _49697_ (.RESET_B(net314),
    .D(net3495),
    .Q(\u_inv.d_reg[87] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _49698_ (.RESET_B(net313),
    .D(net2539),
    .Q(\u_inv.d_reg[88] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _49699_ (.RESET_B(net311),
    .D(net3567),
    .Q(\u_inv.d_reg[89] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _49700_ (.RESET_B(net309),
    .D(_01340_),
    .Q(\u_inv.d_reg[90] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _49701_ (.RESET_B(net307),
    .D(net1639),
    .Q(\u_inv.d_reg[91] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _49702_ (.RESET_B(net306),
    .D(net2476),
    .Q(\u_inv.d_reg[92] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _49703_ (.RESET_B(net304),
    .D(net3176),
    .Q(\u_inv.d_reg[93] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _49704_ (.RESET_B(net302),
    .D(net2084),
    .Q(\u_inv.d_reg[94] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _49705_ (.RESET_B(net300),
    .D(net3641),
    .Q(\u_inv.d_reg[95] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _49706_ (.RESET_B(net299),
    .D(net2320),
    .Q(\u_inv.d_reg[96] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _49707_ (.RESET_B(net297),
    .D(net3653),
    .Q(\u_inv.d_reg[97] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _49708_ (.RESET_B(net296),
    .D(net2973),
    .Q(\u_inv.d_reg[98] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _49709_ (.RESET_B(net294),
    .D(net3665),
    .Q(\u_inv.d_reg[99] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _49710_ (.RESET_B(net293),
    .D(net1702),
    .Q(\u_inv.d_reg[100] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _49711_ (.RESET_B(net291),
    .D(net3120),
    .Q(\u_inv.d_reg[101] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _49712_ (.RESET_B(net290),
    .D(_01352_),
    .Q(\u_inv.d_reg[102] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _49713_ (.RESET_B(net288),
    .D(net3343),
    .Q(\u_inv.d_reg[103] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _49714_ (.RESET_B(net287),
    .D(net2863),
    .Q(\u_inv.d_reg[104] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _49715_ (.RESET_B(net285),
    .D(net2987),
    .Q(\u_inv.d_reg[105] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _49716_ (.RESET_B(net284),
    .D(net2664),
    .Q(\u_inv.d_reg[106] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _49717_ (.RESET_B(net282),
    .D(net2870),
    .Q(\u_inv.d_reg[107] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _49718_ (.RESET_B(net281),
    .D(net3322),
    .Q(\u_inv.d_reg[108] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _49719_ (.RESET_B(net279),
    .D(net2666),
    .Q(\u_inv.d_reg[109] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _49720_ (.RESET_B(net278),
    .D(_01360_),
    .Q(\u_inv.d_reg[110] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _49721_ (.RESET_B(net276),
    .D(net3605),
    .Q(\u_inv.d_reg[111] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _49722_ (.RESET_B(net275),
    .D(_01362_),
    .Q(\u_inv.d_reg[112] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _49723_ (.RESET_B(net273),
    .D(net3053),
    .Q(\u_inv.d_reg[113] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _49724_ (.RESET_B(net272),
    .D(_01364_),
    .Q(\u_inv.d_reg[114] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _49725_ (.RESET_B(net270),
    .D(net2329),
    .Q(\u_inv.d_reg[115] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _49726_ (.RESET_B(net269),
    .D(net2981),
    .Q(\u_inv.d_reg[116] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _49727_ (.RESET_B(net267),
    .D(net2878),
    .Q(\u_inv.d_reg[117] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _49728_ (.RESET_B(net266),
    .D(_01368_),
    .Q(\u_inv.d_reg[118] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _49729_ (.RESET_B(net264),
    .D(net2891),
    .Q(\u_inv.d_reg[119] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _49730_ (.RESET_B(net263),
    .D(net2226),
    .Q(\u_inv.d_reg[120] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _49731_ (.RESET_B(net261),
    .D(net3129),
    .Q(\u_inv.d_reg[121] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _49732_ (.RESET_B(net260),
    .D(net3158),
    .Q(\u_inv.d_reg[122] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _49733_ (.RESET_B(net258),
    .D(net2398),
    .Q(\u_inv.d_reg[123] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _49734_ (.RESET_B(net257),
    .D(net2438),
    .Q(\u_inv.d_reg[124] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _49735_ (.RESET_B(net255),
    .D(net3361),
    .Q(\u_inv.d_reg[125] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _49736_ (.RESET_B(net253),
    .D(net2402),
    .Q(\u_inv.d_reg[126] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _49737_ (.RESET_B(net251),
    .D(_01377_),
    .Q(\u_inv.d_reg[127] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _49738_ (.RESET_B(net250),
    .D(net2588),
    .Q(\u_inv.d_reg[128] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _49739_ (.RESET_B(net248),
    .D(net3300),
    .Q(\u_inv.d_reg[129] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _49740_ (.RESET_B(net246),
    .D(net1243),
    .Q(\u_inv.d_reg[130] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _49741_ (.RESET_B(net244),
    .D(net3364),
    .Q(\u_inv.d_reg[131] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _49742_ (.RESET_B(net243),
    .D(net3414),
    .Q(\u_inv.d_reg[132] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _49743_ (.RESET_B(net241),
    .D(_01383_),
    .Q(\u_inv.d_reg[133] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _49744_ (.RESET_B(net239),
    .D(_01384_),
    .Q(\u_inv.d_reg[134] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _49745_ (.RESET_B(net237),
    .D(net3476),
    .Q(\u_inv.d_reg[135] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _49746_ (.RESET_B(net236),
    .D(net2827),
    .Q(\u_inv.d_reg[136] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _49747_ (.RESET_B(net234),
    .D(net3308),
    .Q(\u_inv.d_reg[137] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _49748_ (.RESET_B(net232),
    .D(_01388_),
    .Q(\u_inv.d_reg[138] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _49749_ (.RESET_B(net230),
    .D(net3569),
    .Q(\u_inv.d_reg[139] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _49750_ (.RESET_B(net229),
    .D(net2607),
    .Q(\u_inv.d_reg[140] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _49751_ (.RESET_B(net227),
    .D(net3254),
    .Q(\u_inv.d_reg[141] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _49752_ (.RESET_B(net225),
    .D(_01392_),
    .Q(\u_inv.d_reg[142] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _49753_ (.RESET_B(net223),
    .D(net3397),
    .Q(\u_inv.d_reg[143] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _49754_ (.RESET_B(net222),
    .D(net2727),
    .Q(\u_inv.d_reg[144] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _49755_ (.RESET_B(net220),
    .D(net2836),
    .Q(\u_inv.d_reg[145] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _49756_ (.RESET_B(net218),
    .D(_01396_),
    .Q(\u_inv.d_reg[146] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _49757_ (.RESET_B(net216),
    .D(net3626),
    .Q(\u_inv.d_reg[147] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _49758_ (.RESET_B(net215),
    .D(net3367),
    .Q(\u_inv.d_reg[148] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _49759_ (.RESET_B(net213),
    .D(net1903),
    .Q(\u_inv.d_reg[149] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _49760_ (.RESET_B(net211),
    .D(_01400_),
    .Q(\u_inv.d_reg[150] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _49761_ (.RESET_B(net209),
    .D(_01401_),
    .Q(\u_inv.d_reg[151] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _49762_ (.RESET_B(net208),
    .D(net2590),
    .Q(\u_inv.d_reg[152] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _49763_ (.RESET_B(net206),
    .D(_01403_),
    .Q(\u_inv.d_reg[153] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _49764_ (.RESET_B(net204),
    .D(net2887),
    .Q(\u_inv.d_reg[154] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _49765_ (.RESET_B(net202),
    .D(net2951),
    .Q(\u_inv.d_reg[155] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _49766_ (.RESET_B(net201),
    .D(net2670),
    .Q(\u_inv.d_reg[156] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _49767_ (.RESET_B(net199),
    .D(net3221),
    .Q(\u_inv.d_reg[157] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _49768_ (.RESET_B(net197),
    .D(net2472),
    .Q(\u_inv.d_reg[158] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _49769_ (.RESET_B(net195),
    .D(net3315),
    .Q(\u_inv.d_reg[159] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _49770_ (.RESET_B(net194),
    .D(net3106),
    .Q(\u_inv.d_reg[160] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _49771_ (.RESET_B(net192),
    .D(net2267),
    .Q(\u_inv.d_reg[161] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _49772_ (.RESET_B(net190),
    .D(_01412_),
    .Q(\u_inv.d_reg[162] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _49773_ (.RESET_B(net188),
    .D(net1497),
    .Q(\u_inv.d_reg[163] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _49774_ (.RESET_B(net186),
    .D(net2713),
    .Q(\u_inv.d_reg[164] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _49775_ (.RESET_B(net184),
    .D(net1540),
    .Q(\u_inv.d_reg[165] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _49776_ (.RESET_B(net183),
    .D(_01416_),
    .Q(\u_inv.d_reg[166] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _49777_ (.RESET_B(net181),
    .D(net3182),
    .Q(\u_inv.d_reg[167] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _49778_ (.RESET_B(net180),
    .D(net3059),
    .Q(\u_inv.d_reg[168] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _49779_ (.RESET_B(net178),
    .D(net3562),
    .Q(\u_inv.d_reg[169] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _49780_ (.RESET_B(net177),
    .D(_01420_),
    .Q(\u_inv.d_reg[170] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _49781_ (.RESET_B(net175),
    .D(net2197),
    .Q(\u_inv.d_reg[171] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _49782_ (.RESET_B(net174),
    .D(net3066),
    .Q(\u_inv.d_reg[172] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _49783_ (.RESET_B(net172),
    .D(net2192),
    .Q(\u_inv.d_reg[173] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _49784_ (.RESET_B(net171),
    .D(_01424_),
    .Q(\u_inv.d_reg[174] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _49785_ (.RESET_B(net169),
    .D(net2579),
    .Q(\u_inv.d_reg[175] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _49786_ (.RESET_B(net168),
    .D(net3112),
    .Q(\u_inv.d_reg[176] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _49787_ (.RESET_B(net166),
    .D(net2708),
    .Q(\u_inv.d_reg[177] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _49788_ (.RESET_B(net165),
    .D(net2075),
    .Q(\u_inv.d_reg[178] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _49789_ (.RESET_B(net163),
    .D(_01429_),
    .Q(\u_inv.d_reg[179] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_2 _49790_ (.RESET_B(net162),
    .D(net2032),
    .Q(\u_inv.d_reg[180] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _49791_ (.RESET_B(net160),
    .D(net1983),
    .Q(\u_inv.d_reg[181] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _49792_ (.RESET_B(net159),
    .D(_01432_),
    .Q(\u_inv.d_reg[182] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _49793_ (.RESET_B(net157),
    .D(net2655),
    .Q(\u_inv.d_reg[183] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _49794_ (.RESET_B(net156),
    .D(_01434_),
    .Q(\u_inv.d_reg[184] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _49795_ (.RESET_B(net154),
    .D(net3375),
    .Q(\u_inv.d_reg[185] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _49796_ (.RESET_B(net153),
    .D(net2441),
    .Q(\u_inv.d_reg[186] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _49797_ (.RESET_B(net151),
    .D(net1484),
    .Q(\u_inv.d_reg[187] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _49798_ (.RESET_B(net150),
    .D(_01438_),
    .Q(\u_inv.d_reg[188] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _49799_ (.RESET_B(net148),
    .D(net3466),
    .Q(\u_inv.d_reg[189] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _49800_ (.RESET_B(net147),
    .D(_01440_),
    .Q(\u_inv.d_reg[190] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _49801_ (.RESET_B(net145),
    .D(net3540),
    .Q(\u_inv.d_reg[191] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _49802_ (.RESET_B(net144),
    .D(net2926),
    .Q(\u_inv.d_reg[192] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _49803_ (.RESET_B(net142),
    .D(_01443_),
    .Q(\u_inv.d_reg[193] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _49804_ (.RESET_B(net141),
    .D(net2448),
    .Q(\u_inv.d_reg[194] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _49805_ (.RESET_B(net139),
    .D(net3390),
    .Q(\u_inv.d_reg[195] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _49806_ (.RESET_B(net138),
    .D(net3550),
    .Q(\u_inv.d_reg[196] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _49807_ (.RESET_B(net917),
    .D(_01447_),
    .Q(\u_inv.d_reg[197] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _49808_ (.RESET_B(net914),
    .D(_01448_),
    .Q(\u_inv.d_reg[198] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _49809_ (.RESET_B(net910),
    .D(net3028),
    .Q(\u_inv.d_reg[199] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _49810_ (.RESET_B(net907),
    .D(net2692),
    .Q(\u_inv.d_reg[200] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _49811_ (.RESET_B(net903),
    .D(net2773),
    .Q(\u_inv.d_reg[201] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _49812_ (.RESET_B(net900),
    .D(_01452_),
    .Q(\u_inv.d_reg[202] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _49813_ (.RESET_B(net896),
    .D(net3456),
    .Q(\u_inv.d_reg[203] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _49814_ (.RESET_B(net893),
    .D(_01454_),
    .Q(\u_inv.d_reg[204] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _49815_ (.RESET_B(net889),
    .D(net2825),
    .Q(\u_inv.d_reg[205] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _49816_ (.RESET_B(net886),
    .D(_01456_),
    .Q(\u_inv.d_reg[206] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _49817_ (.RESET_B(net882),
    .D(net2722),
    .Q(\u_inv.d_reg[207] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _49818_ (.RESET_B(net879),
    .D(net3426),
    .Q(\u_inv.d_reg[208] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _49819_ (.RESET_B(net875),
    .D(net3272),
    .Q(\u_inv.d_reg[209] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _49820_ (.RESET_B(net872),
    .D(net2872),
    .Q(\u_inv.d_reg[210] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _49821_ (.RESET_B(net868),
    .D(net2788),
    .Q(\u_inv.d_reg[211] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _49822_ (.RESET_B(net865),
    .D(net2284),
    .Q(\u_inv.d_reg[212] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _49823_ (.RESET_B(net861),
    .D(net3621),
    .Q(\u_inv.d_reg[213] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _49824_ (.RESET_B(net858),
    .D(net2921),
    .Q(\u_inv.d_reg[214] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _49825_ (.RESET_B(net854),
    .D(net3582),
    .Q(\u_inv.d_reg[215] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _49826_ (.RESET_B(net851),
    .D(net2299),
    .Q(\u_inv.d_reg[216] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _49827_ (.RESET_B(net847),
    .D(net3507),
    .Q(\u_inv.d_reg[217] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _49828_ (.RESET_B(net844),
    .D(net2369),
    .Q(\u_inv.d_reg[218] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _49829_ (.RESET_B(net840),
    .D(net2123),
    .Q(\u_inv.d_reg[219] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _49830_ (.RESET_B(net837),
    .D(net1988),
    .Q(\u_inv.d_reg[220] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _49831_ (.RESET_B(net833),
    .D(net2418),
    .Q(\u_inv.d_reg[221] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _49832_ (.RESET_B(net830),
    .D(net2034),
    .Q(\u_inv.d_reg[222] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _49833_ (.RESET_B(net826),
    .D(net3071),
    .Q(\u_inv.d_reg[223] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _49834_ (.RESET_B(net823),
    .D(net2990),
    .Q(\u_inv.d_reg[224] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _49835_ (.RESET_B(net819),
    .D(_01475_),
    .Q(\u_inv.d_reg[225] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _49836_ (.RESET_B(net816),
    .D(_01476_),
    .Q(\u_inv.d_reg[226] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _49837_ (.RESET_B(net812),
    .D(net3377),
    .Q(\u_inv.d_reg[227] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _49838_ (.RESET_B(net809),
    .D(_01478_),
    .Q(\u_inv.d_reg[228] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _49839_ (.RESET_B(net805),
    .D(net3446),
    .Q(\u_inv.d_reg[229] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _49840_ (.RESET_B(net802),
    .D(_01480_),
    .Q(\u_inv.d_reg[230] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _49841_ (.RESET_B(net798),
    .D(net3150),
    .Q(\u_inv.d_reg[231] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _49842_ (.RESET_B(net795),
    .D(_01482_),
    .Q(\u_inv.d_reg[232] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _49843_ (.RESET_B(net791),
    .D(net3162),
    .Q(\u_inv.d_reg[233] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _49844_ (.RESET_B(net788),
    .D(_01484_),
    .Q(\u_inv.d_reg[234] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _49845_ (.RESET_B(net784),
    .D(net3594),
    .Q(\u_inv.d_reg[235] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _49846_ (.RESET_B(net781),
    .D(_01486_),
    .Q(\u_inv.d_reg[236] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _49847_ (.RESET_B(net777),
    .D(net2127),
    .Q(\u_inv.d_reg[237] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _49848_ (.RESET_B(net774),
    .D(_01488_),
    .Q(\u_inv.d_reg[238] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _49849_ (.RESET_B(net770),
    .D(_01489_),
    .Q(\u_inv.d_reg[239] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _49850_ (.RESET_B(net767),
    .D(net3607),
    .Q(\u_inv.d_reg[240] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _49851_ (.RESET_B(net763),
    .D(net3576),
    .Q(\u_inv.d_reg[241] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _49852_ (.RESET_B(net760),
    .D(_01492_),
    .Q(\u_inv.d_reg[242] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _49853_ (.RESET_B(net756),
    .D(net2311),
    .Q(\u_inv.d_reg[243] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _49854_ (.RESET_B(net753),
    .D(_01494_),
    .Q(\u_inv.d_reg[244] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _49855_ (.RESET_B(net749),
    .D(_01495_),
    .Q(\u_inv.d_reg[245] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _49856_ (.RESET_B(net746),
    .D(_01496_),
    .Q(\u_inv.d_reg[246] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _49857_ (.RESET_B(net742),
    .D(net3018),
    .Q(\u_inv.d_reg[247] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _49858_ (.RESET_B(net739),
    .D(net3544),
    .Q(\u_inv.d_reg[248] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _49859_ (.RESET_B(net735),
    .D(net3505),
    .Q(\u_inv.d_reg[249] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _49860_ (.RESET_B(net732),
    .D(_01500_),
    .Q(\u_inv.d_reg[250] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _49861_ (.RESET_B(net728),
    .D(_01501_),
    .Q(\u_inv.d_reg[251] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _49862_ (.RESET_B(net725),
    .D(_01502_),
    .Q(\u_inv.d_reg[252] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _49863_ (.RESET_B(net721),
    .D(_01503_),
    .Q(\u_inv.d_reg[253] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _49864_ (.RESET_B(net718),
    .D(net2889),
    .Q(\u_inv.d_reg[254] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _49865_ (.RESET_B(net714),
    .D(net3406),
    .Q(\u_inv.d_reg[255] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _49866_ (.RESET_B(net711),
    .D(_01506_),
    .Q(\u_inv.d_reg[256] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _49867_ (.RESET_B(net707),
    .D(_01507_),
    .Q(\u_inv.f_reg[0] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_2 _49868_ (.RESET_B(net704),
    .D(net2182),
    .Q(\u_inv.f_reg[1] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_2 _49869_ (.RESET_B(net700),
    .D(net1348),
    .Q(\u_inv.f_reg[2] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_2 _49870_ (.RESET_B(net697),
    .D(net1723),
    .Q(\u_inv.f_reg[3] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_1 _49871_ (.RESET_B(net693),
    .D(net1754),
    .Q(\u_inv.f_reg[4] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _49872_ (.RESET_B(net690),
    .D(net1443),
    .Q(\u_inv.f_reg[5] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _49873_ (.RESET_B(net686),
    .D(net1637),
    .Q(\u_inv.f_reg[6] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_1 _49874_ (.RESET_B(net683),
    .D(net2133),
    .Q(\u_inv.f_reg[7] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _49875_ (.RESET_B(net679),
    .D(net1550),
    .Q(\u_inv.f_reg[8] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _49876_ (.RESET_B(net676),
    .D(net2629),
    .Q(\u_inv.f_reg[9] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _49877_ (.RESET_B(net672),
    .D(net2026),
    .Q(\u_inv.f_reg[10] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_1 _49878_ (.RESET_B(net669),
    .D(_01518_),
    .Q(\u_inv.f_reg[11] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _49879_ (.RESET_B(net665),
    .D(net1697),
    .Q(\u_inv.f_reg[12] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _49880_ (.RESET_B(net662),
    .D(net2840),
    .Q(\u_inv.f_reg[13] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _49881_ (.RESET_B(net658),
    .D(net1832),
    .Q(\u_inv.f_reg[14] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _49882_ (.RESET_B(net655),
    .D(_01522_),
    .Q(\u_inv.f_reg[15] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _49883_ (.RESET_B(net651),
    .D(net1647),
    .Q(\u_inv.f_reg[16] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _49884_ (.RESET_B(net648),
    .D(net1718),
    .Q(\u_inv.f_reg[17] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _49885_ (.RESET_B(net644),
    .D(net2657),
    .Q(\u_inv.f_reg[18] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _49886_ (.RESET_B(net641),
    .D(net3198),
    .Q(\u_inv.f_reg[19] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _49887_ (.RESET_B(net637),
    .D(net1751),
    .Q(\u_inv.f_reg[20] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _49888_ (.RESET_B(net634),
    .D(net2170),
    .Q(\u_inv.f_reg[21] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _49889_ (.RESET_B(net630),
    .D(net2008),
    .Q(\u_inv.f_reg[22] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _49890_ (.RESET_B(net627),
    .D(net2897),
    .Q(\u_inv.f_reg[23] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _49891_ (.RESET_B(net623),
    .D(net2077),
    .Q(\u_inv.f_reg[24] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _49892_ (.RESET_B(net620),
    .D(net3290),
    .Q(\u_inv.f_reg[25] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _49893_ (.RESET_B(net616),
    .D(net1589),
    .Q(\u_inv.f_reg[26] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_1 _49894_ (.RESET_B(net613),
    .D(net1921),
    .Q(\u_inv.f_reg[27] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _49895_ (.RESET_B(net609),
    .D(net2245),
    .Q(\u_inv.f_reg[28] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _49896_ (.RESET_B(net606),
    .D(net3043),
    .Q(\u_inv.f_reg[29] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _49897_ (.RESET_B(net602),
    .D(net1709),
    .Q(\u_inv.f_reg[30] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _49898_ (.RESET_B(net599),
    .D(net2394),
    .Q(\u_inv.f_reg[31] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _49899_ (.RESET_B(net595),
    .D(net2761),
    .Q(\u_inv.f_reg[32] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_2 _49900_ (.RESET_B(net592),
    .D(net2056),
    .Q(\u_inv.f_reg[33] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_2 _49901_ (.RESET_B(net588),
    .D(net1487),
    .Q(\u_inv.f_reg[34] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_2 _49902_ (.RESET_B(net585),
    .D(net2071),
    .Q(\u_inv.f_reg[35] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_2 _49903_ (.RESET_B(net581),
    .D(net1580),
    .Q(\u_inv.f_reg[36] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_2 _49904_ (.RESET_B(net578),
    .D(net1354),
    .Q(\u_inv.f_reg[37] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_2 _49905_ (.RESET_B(net574),
    .D(net1655),
    .Q(\u_inv.f_reg[38] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_2 _49906_ (.RESET_B(net571),
    .D(net2036),
    .Q(\u_inv.f_reg[39] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_2 _49907_ (.RESET_B(net567),
    .D(net2118),
    .Q(\u_inv.f_reg[40] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_2 _49908_ (.RESET_B(net564),
    .D(_01548_),
    .Q(\u_inv.f_reg[41] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_2 _49909_ (.RESET_B(net560),
    .D(net2686),
    .Q(\u_inv.f_reg[42] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_2 _49910_ (.RESET_B(net557),
    .D(net2942),
    .Q(\u_inv.f_reg[43] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_2 _49911_ (.RESET_B(net553),
    .D(net1445),
    .Q(\u_inv.f_reg[44] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _49912_ (.RESET_B(net550),
    .D(_01552_),
    .Q(\u_inv.f_reg[45] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_2 _49913_ (.RESET_B(net546),
    .D(net2080),
    .Q(\u_inv.f_reg[46] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_2 _49914_ (.RESET_B(net543),
    .D(net2599),
    .Q(\u_inv.f_reg[47] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_2 _49915_ (.RESET_B(net539),
    .D(net1507),
    .Q(\u_inv.f_reg[48] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _49916_ (.RESET_B(net536),
    .D(_01556_),
    .Q(\u_inv.f_reg[49] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_2 _49917_ (.RESET_B(net532),
    .D(net1895),
    .Q(\u_inv.f_reg[50] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_2 _49918_ (.RESET_B(net529),
    .D(net2345),
    .Q(\u_inv.f_reg[51] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_2 _49919_ (.RESET_B(net525),
    .D(net2454),
    .Q(\u_inv.f_reg[52] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_2 _49920_ (.RESET_B(net522),
    .D(net2842),
    .Q(\u_inv.f_reg[53] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_2 _49921_ (.RESET_B(net518),
    .D(net2876),
    .Q(\u_inv.f_reg[54] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_2 _49922_ (.RESET_B(net515),
    .D(net1786),
    .Q(\u_inv.f_reg[55] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_2 _49923_ (.RESET_B(net511),
    .D(net2426),
    .Q(\u_inv.f_reg[56] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_2 _49924_ (.RESET_B(net508),
    .D(net3110),
    .Q(\u_inv.f_reg[57] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_2 _49925_ (.RESET_B(net504),
    .D(net2389),
    .Q(\u_inv.f_reg[58] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_2 _49926_ (.RESET_B(net501),
    .D(net1866),
    .Q(\u_inv.f_reg[59] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _49927_ (.RESET_B(net497),
    .D(net1688),
    .Q(\u_inv.f_reg[60] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _49928_ (.RESET_B(net494),
    .D(net2199),
    .Q(\u_inv.f_reg[61] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _49929_ (.RESET_B(net490),
    .D(net1950),
    .Q(\u_inv.f_reg[62] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _49930_ (.RESET_B(net487),
    .D(net2811),
    .Q(\u_inv.f_reg[63] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _49931_ (.RESET_B(net483),
    .D(net1858),
    .Q(\u_inv.f_reg[64] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _49932_ (.RESET_B(net480),
    .D(net2296),
    .Q(\u_inv.f_reg[65] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_2 _49933_ (.RESET_B(net476),
    .D(net2342),
    .Q(\u_inv.f_reg[66] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_2 _49934_ (.RESET_B(net473),
    .D(net2114),
    .Q(\u_inv.f_reg[67] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_2 _49935_ (.RESET_B(net469),
    .D(net2502),
    .Q(\u_inv.f_reg[68] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_2 _49936_ (.RESET_B(net466),
    .D(net3345),
    .Q(\u_inv.f_reg[69] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_2 _49937_ (.RESET_B(net462),
    .D(net1901),
    .Q(\u_inv.f_reg[70] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_2 _49938_ (.RESET_B(net459),
    .D(net2777),
    .Q(\u_inv.f_reg[71] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_2 _49939_ (.RESET_B(net455),
    .D(net1587),
    .Q(\u_inv.f_reg[72] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_2 _49940_ (.RESET_B(net452),
    .D(net1948),
    .Q(\u_inv.f_reg[73] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_2 _49941_ (.RESET_B(net448),
    .D(net2739),
    .Q(\u_inv.f_reg[74] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_2 _49942_ (.RESET_B(net445),
    .D(net3005),
    .Q(\u_inv.f_reg[75] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_2 _49943_ (.RESET_B(net441),
    .D(net2416),
    .Q(\u_inv.f_reg[76] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_2 _49944_ (.RESET_B(net438),
    .D(net1666),
    .Q(\u_inv.f_reg[77] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_2 _49945_ (.RESET_B(net434),
    .D(net2195),
    .Q(\u_inv.f_reg[78] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_2 _49946_ (.RESET_B(net431),
    .D(net2365),
    .Q(\u_inv.f_reg[79] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_2 _49947_ (.RESET_B(net427),
    .D(net2130),
    .Q(\u_inv.f_reg[80] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_2 _49948_ (.RESET_B(net424),
    .D(net2461),
    .Q(\u_inv.f_reg[81] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_2 _49949_ (.RESET_B(net420),
    .D(net2108),
    .Q(\u_inv.f_reg[82] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _49950_ (.RESET_B(net417),
    .D(net1712),
    .Q(\u_inv.f_reg[83] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _49951_ (.RESET_B(net413),
    .D(net3094),
    .Q(\u_inv.f_reg[84] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_2 _49952_ (.RESET_B(net410),
    .D(net2396),
    .Q(\u_inv.f_reg[85] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _49953_ (.RESET_B(net406),
    .D(net2741),
    .Q(\u_inv.f_reg[86] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _49954_ (.RESET_B(net403),
    .D(_01594_),
    .Q(\u_inv.f_reg[87] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_2 _49955_ (.RESET_B(net399),
    .D(net2092),
    .Q(\u_inv.f_reg[88] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_2 _49956_ (.RESET_B(net396),
    .D(net3069),
    .Q(\u_inv.f_reg[89] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_2 _49957_ (.RESET_B(net392),
    .D(net2024),
    .Q(\u_inv.f_reg[90] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_2 _49958_ (.RESET_B(net389),
    .D(net2360),
    .Q(\u_inv.f_reg[91] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_2 _49959_ (.RESET_B(net385),
    .D(net1633),
    .Q(\u_inv.f_reg[92] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _49960_ (.RESET_B(net382),
    .D(net2028),
    .Q(\u_inv.f_reg[93] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _49961_ (.RESET_B(net378),
    .D(net2221),
    .Q(\u_inv.f_reg[94] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_2 _49962_ (.RESET_B(net375),
    .D(net2215),
    .Q(\u_inv.f_reg[95] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_2 _49963_ (.RESET_B(net371),
    .D(net2492),
    .Q(\u_inv.f_reg[96] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _49964_ (.RESET_B(net368),
    .D(net2073),
    .Q(\u_inv.f_reg[97] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_2 _49965_ (.RESET_B(net364),
    .D(net2684),
    .Q(\u_inv.f_reg[98] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_2 _49966_ (.RESET_B(net361),
    .D(net2223),
    .Q(\u_inv.f_reg[99] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _49967_ (.RESET_B(net357),
    .D(net2201),
    .Q(\u_inv.f_reg[100] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_2 _49968_ (.RESET_B(net354),
    .D(net2242),
    .Q(\u_inv.f_reg[101] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_2 _49969_ (.RESET_B(net350),
    .D(net2406),
    .Q(\u_inv.f_reg[102] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_2 _49970_ (.RESET_B(net347),
    .D(net2813),
    .Q(\u_inv.f_reg[103] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_2 _49971_ (.RESET_B(net343),
    .D(net1643),
    .Q(\u_inv.f_reg[104] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _49972_ (.RESET_B(net340),
    .D(_01612_),
    .Q(\u_inv.f_reg[105] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_2 _49973_ (.RESET_B(net336),
    .D(net2918),
    .Q(\u_inv.f_reg[106] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _49974_ (.RESET_B(net333),
    .D(net1855),
    .Q(\u_inv.f_reg[107] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_2 _49975_ (.RESET_B(net329),
    .D(net2710),
    .Q(\u_inv.f_reg[108] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _49976_ (.RESET_B(net326),
    .D(net1432),
    .Q(\u_inv.f_reg[109] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _49977_ (.RESET_B(net322),
    .D(net1875),
    .Q(\u_inv.f_reg[110] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_2 _49978_ (.RESET_B(net319),
    .D(net3209),
    .Q(\u_inv.f_reg[111] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_2 _49979_ (.RESET_B(net315),
    .D(net2340),
    .Q(\u_inv.f_reg[112] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_2 _49980_ (.RESET_B(net312),
    .D(net2010),
    .Q(\u_inv.f_reg[113] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_2 _49981_ (.RESET_B(net308),
    .D(net2414),
    .Q(\u_inv.f_reg[114] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_2 _49982_ (.RESET_B(net305),
    .D(net3051),
    .Q(\u_inv.f_reg[115] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _49983_ (.RESET_B(net301),
    .D(_01623_),
    .Q(\u_inv.f_reg[116] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _49984_ (.RESET_B(net298),
    .D(net2307),
    .Q(\u_inv.f_reg[117] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _49985_ (.RESET_B(net295),
    .D(net1434),
    .Q(\u_inv.f_reg[118] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _49986_ (.RESET_B(net292),
    .D(net1909),
    .Q(\u_inv.f_reg[119] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _49987_ (.RESET_B(net289),
    .D(net1993),
    .Q(\u_inv.f_reg[120] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_2 _49988_ (.RESET_B(net286),
    .D(net1740),
    .Q(\u_inv.f_reg[121] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_2 _49989_ (.RESET_B(net283),
    .D(net2956),
    .Q(\u_inv.f_reg[122] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_2 _49990_ (.RESET_B(net280),
    .D(net1898),
    .Q(\u_inv.f_reg[123] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_2 _49991_ (.RESET_B(net277),
    .D(net3154),
    .Q(\u_inv.f_reg[124] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _49992_ (.RESET_B(net274),
    .D(net2228),
    .Q(\u_inv.f_reg[125] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _49993_ (.RESET_B(net271),
    .D(net3233),
    .Q(\u_inv.f_reg[126] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_2 _49994_ (.RESET_B(net268),
    .D(net2668),
    .Q(\u_inv.f_reg[127] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_2 _49995_ (.RESET_B(net265),
    .D(net2767),
    .Q(\u_inv.f_reg[128] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _49996_ (.RESET_B(net262),
    .D(net2504),
    .Q(\u_inv.f_reg[129] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_2 _49997_ (.RESET_B(net259),
    .D(net1624),
    .Q(\u_inv.f_reg[130] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _49998_ (.RESET_B(net256),
    .D(net2150),
    .Q(\u_inv.f_reg[131] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _49999_ (.RESET_B(net252),
    .D(net2044),
    .Q(\u_inv.f_reg[132] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _50000_ (.RESET_B(net249),
    .D(net3085),
    .Q(\u_inv.f_reg[133] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _50001_ (.RESET_B(net245),
    .D(net2715),
    .Q(\u_inv.f_reg[134] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _50002_ (.RESET_B(net242),
    .D(net3104),
    .Q(\u_inv.f_reg[135] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _50003_ (.RESET_B(net238),
    .D(net2103),
    .Q(\u_inv.f_reg[136] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _50004_ (.RESET_B(net235),
    .D(net1973),
    .Q(\u_inv.f_reg[137] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _50005_ (.RESET_B(net231),
    .D(net1622),
    .Q(\u_inv.f_reg[138] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _50006_ (.RESET_B(net228),
    .D(net3160),
    .Q(\u_inv.f_reg[139] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _50007_ (.RESET_B(net224),
    .D(net2375),
    .Q(\u_inv.f_reg[140] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _50008_ (.RESET_B(net221),
    .D(net2489),
    .Q(\u_inv.f_reg[141] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _50009_ (.RESET_B(net217),
    .D(net2275),
    .Q(\u_inv.f_reg[142] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _50010_ (.RESET_B(net214),
    .D(net3014),
    .Q(\u_inv.f_reg[143] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _50011_ (.RESET_B(net210),
    .D(net1861),
    .Q(\u_inv.f_reg[144] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _50012_ (.RESET_B(net207),
    .D(_01652_),
    .Q(\u_inv.f_reg[145] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _50013_ (.RESET_B(net203),
    .D(net1668),
    .Q(\u_inv.f_reg[146] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _50014_ (.RESET_B(net200),
    .D(net3114),
    .Q(\u_inv.f_reg[147] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _50015_ (.RESET_B(net196),
    .D(net2769),
    .Q(\u_inv.f_reg[148] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _50016_ (.RESET_B(net193),
    .D(net2905),
    .Q(\u_inv.f_reg[149] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _50017_ (.RESET_B(net189),
    .D(net1821),
    .Q(\u_inv.f_reg[150] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _50018_ (.RESET_B(net185),
    .D(_01658_),
    .Q(\u_inv.f_reg[151] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _50019_ (.RESET_B(net182),
    .D(net2749),
    .Q(\u_inv.f_reg[152] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _50020_ (.RESET_B(net179),
    .D(net2882),
    .Q(\u_inv.f_reg[153] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _50021_ (.RESET_B(net176),
    .D(net1788),
    .Q(\u_inv.f_reg[154] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _50022_ (.RESET_B(net173),
    .D(net2178),
    .Q(\u_inv.f_reg[155] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _50023_ (.RESET_B(net170),
    .D(net1635),
    .Q(\u_inv.f_reg[156] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _50024_ (.RESET_B(net167),
    .D(net2997),
    .Q(\u_inv.f_reg[157] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _50025_ (.RESET_B(net164),
    .D(net2541),
    .Q(\u_inv.f_reg[158] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _50026_ (.RESET_B(net161),
    .D(net2356),
    .Q(\u_inv.f_reg[159] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _50027_ (.RESET_B(net158),
    .D(net2641),
    .Q(\u_inv.f_reg[160] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _50028_ (.RESET_B(net155),
    .D(net2907),
    .Q(\u_inv.f_reg[161] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _50029_ (.RESET_B(net152),
    .D(net1845),
    .Q(\u_inv.f_reg[162] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_1 _50030_ (.RESET_B(net149),
    .D(net1253),
    .Q(\u_inv.f_reg[163] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _50031_ (.RESET_B(net146),
    .D(net2603),
    .Q(\u_inv.f_reg[164] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _50032_ (.RESET_B(net143),
    .D(_01672_),
    .Q(\u_inv.f_reg[165] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _50033_ (.RESET_B(net140),
    .D(net2378),
    .Q(\u_inv.f_reg[166] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _50034_ (.RESET_B(net137),
    .D(net2186),
    .Q(\u_inv.f_reg[167] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _50035_ (.RESET_B(net912),
    .D(net2865),
    .Q(\u_inv.f_reg[168] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _50036_ (.RESET_B(net905),
    .D(net2433),
    .Q(\u_inv.f_reg[169] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _50037_ (.RESET_B(net898),
    .D(net2018),
    .Q(\u_inv.f_reg[170] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _50038_ (.RESET_B(net891),
    .D(_01678_),
    .Q(\u_inv.f_reg[171] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _50039_ (.RESET_B(net884),
    .D(net2617),
    .Q(\u_inv.f_reg[172] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _50040_ (.RESET_B(net877),
    .D(net1790),
    .Q(\u_inv.f_reg[173] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _50041_ (.RESET_B(net870),
    .D(net1778),
    .Q(\u_inv.f_reg[174] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _50042_ (.RESET_B(net863),
    .D(_01682_),
    .Q(\u_inv.f_reg[175] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _50043_ (.RESET_B(net856),
    .D(net3033),
    .Q(\u_inv.f_reg[176] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _50044_ (.RESET_B(net849),
    .D(_01684_),
    .Q(\u_inv.f_reg[177] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _50045_ (.RESET_B(net842),
    .D(net2790),
    .Q(\u_inv.f_reg[178] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_2 _50046_ (.RESET_B(net835),
    .D(_01686_),
    .Q(\u_inv.f_reg[179] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _50047_ (.RESET_B(net828),
    .D(_01687_),
    .Q(\u_inv.f_reg[180] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _50048_ (.RESET_B(net821),
    .D(net2105),
    .Q(\u_inv.f_reg[181] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _50049_ (.RESET_B(net814),
    .D(net2796),
    .Q(\u_inv.f_reg[182] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_1 _50050_ (.RESET_B(net807),
    .D(net1186),
    .Q(\u_inv.f_reg[183] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_2 _50051_ (.RESET_B(net800),
    .D(net1651),
    .Q(\u_inv.f_reg[184] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _50052_ (.RESET_B(net793),
    .D(net3137),
    .Q(\u_inv.f_reg[185] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _50053_ (.RESET_B(net786),
    .D(net2560),
    .Q(\u_inv.f_reg[186] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _50054_ (.RESET_B(net779),
    .D(net2594),
    .Q(\u_inv.f_reg[187] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _50055_ (.RESET_B(net772),
    .D(net1958),
    .Q(\u_inv.f_reg[188] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_1 _50056_ (.RESET_B(net765),
    .D(net1997),
    .Q(\u_inv.f_reg[189] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_2 _50057_ (.RESET_B(net758),
    .D(net2205),
    .Q(\u_inv.f_reg[190] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_2 _50058_ (.RESET_B(net751),
    .D(net2677),
    .Q(\u_inv.f_reg[191] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_2 _50059_ (.RESET_B(net744),
    .D(net3091),
    .Q(\u_inv.f_reg[192] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_2 _50060_ (.RESET_B(net737),
    .D(net2420),
    .Q(\u_inv.f_reg[193] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_2 _50061_ (.RESET_B(net730),
    .D(net2386),
    .Q(\u_inv.f_reg[194] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_2 _50062_ (.RESET_B(net723),
    .D(net2568),
    .Q(\u_inv.f_reg[195] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_2 _50063_ (.RESET_B(net716),
    .D(net3156),
    .Q(\u_inv.f_reg[196] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_2 _50064_ (.RESET_B(net709),
    .D(net2867),
    .Q(\u_inv.f_reg[197] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_2 _50065_ (.RESET_B(net702),
    .D(net1954),
    .Q(\u_inv.f_reg[198] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_2 _50066_ (.RESET_B(net695),
    .D(_01706_),
    .Q(\u_inv.f_reg[199] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_2 _50067_ (.RESET_B(net688),
    .D(net2959),
    .Q(\u_inv.f_reg[200] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _50068_ (.RESET_B(net681),
    .D(net2409),
    .Q(\u_inv.f_reg[201] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_2 _50069_ (.RESET_B(net674),
    .D(net1811),
    .Q(\u_inv.f_reg[202] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_2 _50070_ (.RESET_B(net667),
    .D(net2985),
    .Q(\u_inv.f_reg[203] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_2 _50071_ (.RESET_B(net660),
    .D(net2350),
    .Q(\u_inv.f_reg[204] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_2 _50072_ (.RESET_B(net653),
    .D(net1774),
    .Q(\u_inv.f_reg[205] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_2 _50073_ (.RESET_B(net646),
    .D(net2532),
    .Q(\u_inv.f_reg[206] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_2 _50074_ (.RESET_B(net639),
    .D(net2164),
    .Q(\u_inv.f_reg[207] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_2 _50075_ (.RESET_B(net632),
    .D(net3245),
    .Q(\u_inv.f_reg[208] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_2 _50076_ (.RESET_B(net625),
    .D(net2309),
    .Q(\u_inv.f_reg[209] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_2 _50077_ (.RESET_B(net618),
    .D(net3132),
    .Q(\u_inv.f_reg[210] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_2 _50078_ (.RESET_B(net611),
    .D(net2463),
    .Q(\u_inv.f_reg[211] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_2 _50079_ (.RESET_B(net604),
    .D(net2944),
    .Q(\u_inv.f_reg[212] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_2 _50080_ (.RESET_B(net597),
    .D(net2754),
    .Q(\u_inv.f_reg[213] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_2 _50081_ (.RESET_B(net590),
    .D(net2517),
    .Q(\u_inv.f_reg[214] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_2 _50082_ (.RESET_B(net583),
    .D(net2446),
    .Q(\u_inv.f_reg[215] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_1 _50083_ (.RESET_B(net576),
    .D(_01723_),
    .Q(\u_inv.f_reg[216] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _50084_ (.RESET_B(net569),
    .D(_01724_),
    .Q(\u_inv.f_reg[217] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _50085_ (.RESET_B(net562),
    .D(net2700),
    .Q(\u_inv.f_reg[218] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _50086_ (.RESET_B(net555),
    .D(_01726_),
    .Q(\u_inv.f_reg[219] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _50087_ (.RESET_B(net548),
    .D(net2967),
    .Q(\u_inv.f_reg[220] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _50088_ (.RESET_B(net541),
    .D(net3035),
    .Q(\u_inv.f_reg[221] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_2 _50089_ (.RESET_B(net534),
    .D(net2696),
    .Q(\u_inv.f_reg[222] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_2 _50090_ (.RESET_B(net527),
    .D(net2207),
    .Q(\u_inv.f_reg[223] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_2 _50091_ (.RESET_B(net520),
    .D(net1578),
    .Q(\u_inv.f_reg[224] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_2 _50092_ (.RESET_B(net513),
    .D(net3204),
    .Q(\u_inv.f_reg[225] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_2 _50093_ (.RESET_B(net506),
    .D(net1747),
    .Q(\u_inv.f_reg[226] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _50094_ (.RESET_B(net499),
    .D(net2168),
    .Q(\u_inv.f_reg[227] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _50095_ (.RESET_B(net492),
    .D(net2903),
    .Q(\u_inv.f_reg[228] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _50096_ (.RESET_B(net485),
    .D(net1843),
    .Q(\u_inv.f_reg[229] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _50097_ (.RESET_B(net478),
    .D(net2856),
    .Q(\u_inv.f_reg[230] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _50098_ (.RESET_B(net471),
    .D(_01738_),
    .Q(\u_inv.f_reg[231] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _50099_ (.RESET_B(net464),
    .D(net2885),
    .Q(\u_inv.f_reg[232] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _50100_ (.RESET_B(net457),
    .D(_01740_),
    .Q(\u_inv.f_reg[233] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _50101_ (.RESET_B(net450),
    .D(net3277),
    .Q(\u_inv.f_reg[234] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _50102_ (.RESET_B(net443),
    .D(net2147),
    .Q(\u_inv.f_reg[235] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _50103_ (.RESET_B(net436),
    .D(net3030),
    .Q(\u_inv.f_reg[236] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _50104_ (.RESET_B(net429),
    .D(net2141),
    .Q(\u_inv.f_reg[237] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _50105_ (.RESET_B(net422),
    .D(net1941),
    .Q(\u_inv.f_reg[238] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _50106_ (.RESET_B(net415),
    .D(net2909),
    .Q(\u_inv.f_reg[239] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _50107_ (.RESET_B(net408),
    .D(net2643),
    .Q(\u_inv.f_reg[240] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _50108_ (.RESET_B(net401),
    .D(net2333),
    .Q(\u_inv.f_reg[241] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _50109_ (.RESET_B(net394),
    .D(net2725),
    .Q(\u_inv.f_reg[242] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _50110_ (.RESET_B(net387),
    .D(_01750_),
    .Q(\u_inv.f_reg[243] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _50111_ (.RESET_B(net380),
    .D(net2681),
    .Q(\u_inv.f_reg[244] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _50112_ (.RESET_B(net373),
    .D(net2232),
    .Q(\u_inv.f_reg[245] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _50113_ (.RESET_B(net366),
    .D(net1914),
    .Q(\u_inv.f_reg[246] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _50114_ (.RESET_B(net359),
    .D(net3056),
    .Q(\u_inv.f_reg[247] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _50115_ (.RESET_B(net352),
    .D(net2689),
    .Q(\u_inv.f_reg[248] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _50116_ (.RESET_B(net345),
    .D(net2858),
    .Q(\u_inv.f_reg[249] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _50117_ (.RESET_B(net338),
    .D(net2166),
    .Q(\u_inv.f_reg[250] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _50118_ (.RESET_B(net331),
    .D(net2624),
    .Q(\u_inv.f_reg[251] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _50119_ (.RESET_B(net324),
    .D(net2527),
    .Q(\u_inv.f_reg[252] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _50120_ (.RESET_B(net317),
    .D(net3073),
    .Q(\u_inv.f_reg[253] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _50121_ (.RESET_B(net310),
    .D(net2661),
    .Q(\u_inv.f_reg[254] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _50122_ (.RESET_B(net303),
    .D(net3215),
    .Q(\u_inv.f_reg[255] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _50123_ (.RESET_B(net187),
    .D(_01763_),
    .Q(\u_inv.f_reg[256] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _50124_ (.RESET_B(net7449),
    .D(_24689_[0]),
    .Q(\u_inv.load_input ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _50125_ (.RESET_B(net7453),
    .D(_01764_),
    .Q(\u_inv.state[0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _50126_ (.RESET_B(net7449),
    .D(_01765_),
    .Q(\u_inv.state[1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _50127_ (.RESET_B(net7423),
    .D(_01766_),
    .Q(\perf_triple[0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _50128_ (.RESET_B(net7422),
    .D(_01767_),
    .Q(\perf_triple[1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _50129_ (.RESET_B(net7427),
    .D(_01768_),
    .Q(\perf_triple[2] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _50130_ (.RESET_B(net7423),
    .D(_01769_),
    .Q(\perf_triple[3] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _50131_ (.RESET_B(net7422),
    .D(_01770_),
    .Q(\perf_triple[4] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _50132_ (.RESET_B(net7423),
    .D(_01771_),
    .Q(\perf_triple[5] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _50133_ (.RESET_B(net7423),
    .D(_01772_),
    .Q(\perf_triple[6] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _50134_ (.RESET_B(net7422),
    .D(_01773_),
    .Q(\perf_triple[7] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _50135_ (.RESET_B(net7441),
    .D(_01774_),
    .Q(\perf_triple[8] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _50136_ (.RESET_B(net7442),
    .D(_01775_),
    .Q(\perf_triple[9] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _50137_ (.RESET_B(net254),
    .D(_01776_),
    .Q(\u_inv.delta_double[0] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _50138_ (.RESET_B(net247),
    .D(_01777_),
    .Q(\u_inv.delta_reg[1] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _50139_ (.RESET_B(net240),
    .D(_01778_),
    .Q(\u_inv.delta_reg[2] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _50140_ (.RESET_B(net233),
    .D(_01779_),
    .Q(\u_inv.delta_reg[3] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _50141_ (.RESET_B(net226),
    .D(_01780_),
    .Q(\u_inv.delta_reg[4] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _50142_ (.RESET_B(net219),
    .D(_01781_),
    .Q(\u_inv.delta_reg[5] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _50143_ (.RESET_B(net212),
    .D(net1172),
    .Q(\u_inv.delta_reg[6] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _50144_ (.RESET_B(net205),
    .D(_01783_),
    .Q(\u_inv.delta_reg[7] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _50145_ (.RESET_B(net198),
    .D(_01784_),
    .Q(\u_inv.delta_reg[8] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _50146_ (.RESET_B(net191),
    .D(net1250),
    .Q(\u_inv.delta_reg[9] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _50147_ (.RESET_B(net7426),
    .D(net3744),
    .Q(\u_inv.counter[0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _50148_ (.RESET_B(net7459),
    .D(net1234),
    .Q(\inv_cycles[0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _50149_ (.RESET_B(net7459),
    .D(net2203),
    .Q(\inv_cycles[1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _50150_ (.RESET_B(net7425),
    .D(net2305),
    .Q(\inv_cycles[2] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _50151_ (.RESET_B(net7426),
    .D(net1213),
    .Q(\inv_cycles[3] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _50152_ (.RESET_B(net7426),
    .D(net1204),
    .Q(\inv_cycles[4] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _50153_ (.RESET_B(net7425),
    .D(net1189),
    .Q(\inv_cycles[5] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _50154_ (.RESET_B(net7425),
    .D(net1879),
    .Q(\inv_cycles[6] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _50155_ (.RESET_B(net7424),
    .D(net1767),
    .Q(\inv_cycles[7] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _50156_ (.RESET_B(net7424),
    .D(net1736),
    .Q(\inv_cycles[8] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _50157_ (.RESET_B(net7425),
    .D(net1416),
    .Q(\inv_cycles[9] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _50158_ (.RESET_B(net7419),
    .D(_01797_),
    .Q(\u_inv.counter[1] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _50159_ (.RESET_B(net7419),
    .D(_01798_),
    .Q(\u_inv.counter[2] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _50160_ (.RESET_B(net7419),
    .D(net1619),
    .Q(\u_inv.counter[3] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _50161_ (.RESET_B(net7419),
    .D(_01800_),
    .Q(\u_inv.counter[4] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _50162_ (.RESET_B(net7425),
    .D(_01801_),
    .Q(\u_inv.counter[5] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _50163_ (.RESET_B(net7425),
    .D(_01802_),
    .Q(\u_inv.counter[6] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _50164_ (.RESET_B(net7425),
    .D(_01803_),
    .Q(\u_inv.counter[7] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _50165_ (.RESET_B(net7425),
    .D(net3759),
    .Q(\u_inv.counter[8] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _50166_ (.RESET_B(net7426),
    .D(_01805_),
    .Q(\u_inv.counter[9] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _50167_ (.RESET_B(net7456),
    .D(net1307),
    .Q(\u_inv.input_reg[0] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _50168_ (.RESET_B(net7462),
    .D(net1925),
    .Q(\u_inv.input_reg[1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _50169_ (.RESET_B(net7458),
    .D(net1538),
    .Q(\u_inv.input_reg[2] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _50170_ (.RESET_B(net7463),
    .D(net1649),
    .Q(\u_inv.input_reg[3] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_1 _50171_ (.RESET_B(net7464),
    .D(net1296),
    .Q(\u_inv.input_reg[4] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _50172_ (.RESET_B(net7463),
    .D(net1889),
    .Q(\u_inv.input_reg[5] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_1 _50173_ (.RESET_B(net7463),
    .D(net1568),
    .Q(\u_inv.input_reg[6] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _50174_ (.RESET_B(net7471),
    .D(net1761),
    .Q(\u_inv.input_reg[7] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _50175_ (.RESET_B(net7477),
    .D(net1294),
    .Q(\u_inv.input_reg[8] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_1 _50176_ (.RESET_B(net7477),
    .D(net1392),
    .Q(\u_inv.input_reg[9] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_1 _50177_ (.RESET_B(net7478),
    .D(net1332),
    .Q(\u_inv.input_reg[10] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_1 _50178_ (.RESET_B(net7477),
    .D(net1449),
    .Q(\u_inv.input_reg[11] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_1 _50179_ (.RESET_B(net7478),
    .D(net1275),
    .Q(\u_inv.input_reg[12] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_1 _50180_ (.RESET_B(net7482),
    .D(net1695),
    .Q(\u_inv.input_reg[13] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _50181_ (.RESET_B(net7478),
    .D(net1303),
    .Q(\u_inv.input_reg[14] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _50182_ (.RESET_B(net7484),
    .D(net1613),
    .Q(\u_inv.input_reg[15] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _50183_ (.RESET_B(net7485),
    .D(net1871),
    .Q(\u_inv.input_reg[16] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_1 _50184_ (.RESET_B(net7488),
    .D(net1453),
    .Q(\u_inv.input_reg[17] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_1 _50185_ (.RESET_B(net7485),
    .D(net1370),
    .Q(\u_inv.input_reg[18] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _50186_ (.RESET_B(net7490),
    .D(net2054),
    .Q(\u_inv.input_reg[19] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _50187_ (.RESET_B(net7490),
    .D(net1376),
    .Q(\u_inv.input_reg[20] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _50188_ (.RESET_B(net7491),
    .D(net1693),
    .Q(\u_inv.input_reg[21] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _50189_ (.RESET_B(net7495),
    .D(net1510),
    .Q(\u_inv.input_reg[22] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_1 _50190_ (.RESET_B(net7495),
    .D(net1336),
    .Q(\u_inv.input_reg[23] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_1 _50191_ (.RESET_B(net7490),
    .D(net1451),
    .Q(\u_inv.input_reg[24] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_1 _50192_ (.RESET_B(net7496),
    .D(net1558),
    .Q(\u_inv.input_reg[25] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_1 _50193_ (.RESET_B(net7499),
    .D(net1344),
    .Q(\u_inv.input_reg[26] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_1 _50194_ (.RESET_B(net7512),
    .D(net1319),
    .Q(\u_inv.input_reg[27] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_1 _50195_ (.RESET_B(net7514),
    .D(net1380),
    .Q(\u_inv.input_reg[28] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_1 _50196_ (.RESET_B(net7517),
    .D(net1300),
    .Q(\u_inv.input_reg[29] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_1 _50197_ (.RESET_B(net7518),
    .D(net1745),
    .Q(\u_inv.input_reg[30] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_1 _50198_ (.RESET_B(net7518),
    .D(net1501),
    .Q(\u_inv.input_reg[31] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_1 _50199_ (.RESET_B(net7517),
    .D(net1269),
    .Q(\u_inv.input_reg[32] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_1 _50200_ (.RESET_B(net7517),
    .D(net1421),
    .Q(\u_inv.input_reg[33] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_1 _50201_ (.RESET_B(net7517),
    .D(net1346),
    .Q(\u_inv.input_reg[34] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_1 _50202_ (.RESET_B(net7520),
    .D(net1257),
    .Q(\u_inv.input_reg[35] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _50203_ (.RESET_B(net7526),
    .D(net1265),
    .Q(\u_inv.input_reg[36] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _50204_ (.RESET_B(net7520),
    .D(net1809),
    .Q(\u_inv.input_reg[37] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _50205_ (.RESET_B(net7526),
    .D(net1352),
    .Q(\u_inv.input_reg[38] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _50206_ (.RESET_B(net7526),
    .D(net1305),
    .Q(\u_inv.input_reg[39] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _50207_ (.RESET_B(net7526),
    .D(net1591),
    .Q(\u_inv.input_reg[40] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _50208_ (.RESET_B(net7519),
    .D(net2152),
    .Q(\u_inv.input_reg[41] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _50209_ (.RESET_B(net7527),
    .D(net1756),
    .Q(\u_inv.input_reg[42] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _50210_ (.RESET_B(net7527),
    .D(net1600),
    .Q(\u_inv.input_reg[43] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _50211_ (.RESET_B(net7528),
    .D(net1412),
    .Q(\u_inv.input_reg[44] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _50212_ (.RESET_B(net7527),
    .D(net1877),
    .Q(\u_inv.input_reg[45] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _50213_ (.RESET_B(net7532),
    .D(net1350),
    .Q(\u_inv.input_reg[46] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _50214_ (.RESET_B(net7532),
    .D(net1524),
    .Q(\u_inv.input_reg[47] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _50215_ (.RESET_B(net7531),
    .D(net1263),
    .Q(\u_inv.input_reg[48] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _50216_ (.RESET_B(net7532),
    .D(net1478),
    .Q(\u_inv.input_reg[49] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _50217_ (.RESET_B(net7533),
    .D(net1493),
    .Q(\u_inv.input_reg[50] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _50218_ (.RESET_B(net7537),
    .D(net1491),
    .Q(\u_inv.input_reg[51] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _50219_ (.RESET_B(net7533),
    .D(net1542),
    .Q(\u_inv.input_reg[52] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _50220_ (.RESET_B(net7531),
    .D(net1891),
    .Q(\u_inv.input_reg[53] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _50221_ (.RESET_B(net7533),
    .D(net1468),
    .Q(\u_inv.input_reg[54] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _50222_ (.RESET_B(net7550),
    .D(net1967),
    .Q(\u_inv.input_reg[55] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _50223_ (.RESET_B(net7550),
    .D(net1374),
    .Q(\u_inv.input_reg[56] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _50224_ (.RESET_B(net7557),
    .D(net1598),
    .Q(\u_inv.input_reg[57] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _50225_ (.RESET_B(net7533),
    .D(net1573),
    .Q(\u_inv.input_reg[58] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _50226_ (.RESET_B(net7550),
    .D(net1466),
    .Q(\u_inv.input_reg[59] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _50227_ (.RESET_B(net7533),
    .D(net1671),
    .Q(\u_inv.input_reg[60] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _50228_ (.RESET_B(net7552),
    .D(net1595),
    .Q(\u_inv.input_reg[61] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _50229_ (.RESET_B(net7552),
    .D(net1826),
    .Q(\u_inv.input_reg[62] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _50230_ (.RESET_B(net7552),
    .D(net1418),
    .Q(\u_inv.input_reg[63] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _50231_ (.RESET_B(net7560),
    .D(net1617),
    .Q(\u_inv.input_reg[64] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _50232_ (.RESET_B(net7558),
    .D(net1738),
    .Q(\u_inv.input_reg[65] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _50233_ (.RESET_B(net7560),
    .D(net1602),
    .Q(\u_inv.input_reg[66] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _50234_ (.RESET_B(net7560),
    .D(net1758),
    .Q(\u_inv.input_reg[67] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _50235_ (.RESET_B(net7560),
    .D(net1952),
    .Q(\u_inv.input_reg[68] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _50236_ (.RESET_B(net7561),
    .D(net1781),
    .Q(\u_inv.input_reg[69] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _50237_ (.RESET_B(net7561),
    .D(net1830),
    .Q(\u_inv.input_reg[70] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _50238_ (.RESET_B(net7559),
    .D(net1585),
    .Q(\u_inv.input_reg[71] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _50239_ (.RESET_B(net7561),
    .D(net2086),
    .Q(\u_inv.input_reg[72] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _50240_ (.RESET_B(net7561),
    .D(net1472),
    .Q(\u_inv.input_reg[73] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _50241_ (.RESET_B(net7562),
    .D(net2154),
    .Q(\u_inv.input_reg[74] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _50242_ (.RESET_B(net7561),
    .D(net1676),
    .Q(\u_inv.input_reg[75] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _50243_ (.RESET_B(net7559),
    .D(net2189),
    .Q(\u_inv.input_reg[76] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _50244_ (.RESET_B(net7562),
    .D(net1828),
    .Q(\u_inv.input_reg[77] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _50245_ (.RESET_B(net7562),
    .D(net2004),
    .Q(\u_inv.input_reg[78] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _50246_ (.RESET_B(net7559),
    .D(net1554),
    .Q(\u_inv.input_reg[79] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _50247_ (.RESET_B(net7561),
    .D(net1792),
    .Q(\u_inv.input_reg[80] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _50248_ (.RESET_B(net7561),
    .D(net1816),
    .Q(\u_inv.input_reg[81] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _50249_ (.RESET_B(net7561),
    .D(net1772),
    .Q(\u_inv.input_reg[82] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _50250_ (.RESET_B(net7564),
    .D(net1424),
    .Q(\u_inv.input_reg[83] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _50251_ (.RESET_B(net7564),
    .D(net1359),
    .Q(\u_inv.input_reg[84] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _50252_ (.RESET_B(net7566),
    .D(net1935),
    .Q(\u_inv.input_reg[85] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _50253_ (.RESET_B(net7566),
    .D(net1615),
    .Q(\u_inv.input_reg[86] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _50254_ (.RESET_B(net7566),
    .D(net1372),
    .Q(\u_inv.input_reg[87] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _50255_ (.RESET_B(net7566),
    .D(net1461),
    .Q(\u_inv.input_reg[88] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _50256_ (.RESET_B(net7566),
    .D(net1436),
    .Q(\u_inv.input_reg[89] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _50257_ (.RESET_B(net7566),
    .D(net1720),
    .Q(\u_inv.input_reg[90] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _50258_ (.RESET_B(net7566),
    .D(net1527),
    .Q(\u_inv.input_reg[91] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _50259_ (.RESET_B(net7564),
    .D(net1534),
    .Q(\u_inv.input_reg[92] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _50260_ (.RESET_B(net7567),
    .D(net2088),
    .Q(\u_inv.input_reg[93] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _50261_ (.RESET_B(net7565),
    .D(net1609),
    .Q(\u_inv.input_reg[94] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_tiehi _48933__22 (.L_HI(net22));
 sg13g2_tiehi _48932__23 (.L_HI(net23));
 sg13g2_tiehi _48931__24 (.L_HI(net24));
 sg13g2_tiehi _48930__25 (.L_HI(net25));
 sg13g2_tiehi _48929__26 (.L_HI(net26));
 sg13g2_tiehi _48928__27 (.L_HI(net27));
 sg13g2_tiehi _48927__28 (.L_HI(net28));
 sg13g2_tiehi _48926__29 (.L_HI(net29));
 sg13g2_tiehi _48925__30 (.L_HI(net30));
 sg13g2_tiehi _48924__31 (.L_HI(net31));
 sg13g2_tiehi _48923__32 (.L_HI(net32));
 sg13g2_tiehi _48922__33 (.L_HI(net33));
 sg13g2_tiehi _48921__34 (.L_HI(net34));
 sg13g2_tiehi _48920__35 (.L_HI(net35));
 sg13g2_tiehi _48919__36 (.L_HI(net36));
 sg13g2_tiehi _48918__37 (.L_HI(net37));
 sg13g2_tiehi _48917__38 (.L_HI(net38));
 sg13g2_tiehi _48916__39 (.L_HI(net39));
 sg13g2_tiehi _48915__40 (.L_HI(net40));
 sg13g2_tiehi _48914__41 (.L_HI(net41));
 sg13g2_tiehi _48913__42 (.L_HI(net42));
 sg13g2_tiehi _48912__43 (.L_HI(net43));
 sg13g2_tiehi _48911__44 (.L_HI(net44));
 sg13g2_tiehi _48910__45 (.L_HI(net45));
 sg13g2_tiehi _48909__46 (.L_HI(net46));
 sg13g2_tiehi _48908__47 (.L_HI(net47));
 sg13g2_tiehi _48907__48 (.L_HI(net48));
 sg13g2_tiehi _48906__49 (.L_HI(net49));
 sg13g2_tiehi _48905__50 (.L_HI(net50));
 sg13g2_tiehi _48904__51 (.L_HI(net51));
 sg13g2_tiehi _48903__52 (.L_HI(net52));
 sg13g2_tiehi _48902__53 (.L_HI(net53));
 sg13g2_tiehi _48901__54 (.L_HI(net54));
 sg13g2_tiehi _48900__55 (.L_HI(net55));
 sg13g2_tiehi _48899__56 (.L_HI(net56));
 sg13g2_tiehi _48898__57 (.L_HI(net57));
 sg13g2_tiehi _48897__58 (.L_HI(net58));
 sg13g2_tiehi _48896__59 (.L_HI(net59));
 sg13g2_tiehi _48895__60 (.L_HI(net60));
 sg13g2_tiehi _48894__61 (.L_HI(net61));
 sg13g2_tiehi _48893__62 (.L_HI(net62));
 sg13g2_tiehi _48892__63 (.L_HI(net63));
 sg13g2_tiehi _48891__64 (.L_HI(net64));
 sg13g2_tiehi _48890__65 (.L_HI(net65));
 sg13g2_tiehi _48889__66 (.L_HI(net66));
 sg13g2_tiehi _48888__67 (.L_HI(net67));
 sg13g2_tiehi _48887__68 (.L_HI(net68));
 sg13g2_tiehi _48886__69 (.L_HI(net69));
 sg13g2_tiehi _48885__70 (.L_HI(net70));
 sg13g2_tiehi _48884__71 (.L_HI(net71));
 sg13g2_tiehi _48883__72 (.L_HI(net72));
 sg13g2_tiehi _48882__73 (.L_HI(net73));
 sg13g2_tiehi _48881__74 (.L_HI(net74));
 sg13g2_tiehi _48880__75 (.L_HI(net75));
 sg13g2_tiehi _48879__76 (.L_HI(net76));
 sg13g2_tiehi _48878__77 (.L_HI(net77));
 sg13g2_tiehi _48877__78 (.L_HI(net78));
 sg13g2_tiehi _48876__79 (.L_HI(net79));
 sg13g2_tiehi _48875__80 (.L_HI(net80));
 sg13g2_tiehi _48874__81 (.L_HI(net81));
 sg13g2_tiehi _48873__82 (.L_HI(net82));
 sg13g2_tiehi _48872__83 (.L_HI(net83));
 sg13g2_tiehi _48871__84 (.L_HI(net84));
 sg13g2_tiehi _48870__85 (.L_HI(net85));
 sg13g2_tiehi _48869__86 (.L_HI(net86));
 sg13g2_tiehi _48868__87 (.L_HI(net87));
 sg13g2_tiehi _48867__88 (.L_HI(net88));
 sg13g2_tiehi _48866__89 (.L_HI(net89));
 sg13g2_tiehi _48865__90 (.L_HI(net90));
 sg13g2_tiehi _48864__91 (.L_HI(net91));
 sg13g2_tiehi _48863__92 (.L_HI(net92));
 sg13g2_tiehi _48862__93 (.L_HI(net93));
 sg13g2_tiehi _48861__94 (.L_HI(net94));
 sg13g2_tiehi _48860__95 (.L_HI(net95));
 sg13g2_tiehi _48859__96 (.L_HI(net96));
 sg13g2_tiehi _48858__97 (.L_HI(net97));
 sg13g2_tiehi _48857__98 (.L_HI(net98));
 sg13g2_tiehi _48856__99 (.L_HI(net99));
 sg13g2_tiehi _48855__100 (.L_HI(net100));
 sg13g2_tiehi _48854__101 (.L_HI(net101));
 sg13g2_tiehi _48853__102 (.L_HI(net102));
 sg13g2_tiehi _48852__103 (.L_HI(net103));
 sg13g2_tiehi _48851__104 (.L_HI(net104));
 sg13g2_tiehi _48850__105 (.L_HI(net105));
 sg13g2_tiehi _48849__106 (.L_HI(net106));
 sg13g2_tiehi _48848__107 (.L_HI(net107));
 sg13g2_tiehi _48847__108 (.L_HI(net108));
 sg13g2_tiehi _48846__109 (.L_HI(net109));
 sg13g2_tiehi _48845__110 (.L_HI(net110));
 sg13g2_tiehi _48844__111 (.L_HI(net111));
 sg13g2_tiehi _48843__112 (.L_HI(net112));
 sg13g2_tiehi _48842__113 (.L_HI(net113));
 sg13g2_tiehi _48841__114 (.L_HI(net114));
 sg13g2_tiehi _48840__115 (.L_HI(net115));
 sg13g2_tiehi _48839__116 (.L_HI(net116));
 sg13g2_tiehi _48838__117 (.L_HI(net117));
 sg13g2_tiehi _48837__118 (.L_HI(net118));
 sg13g2_tiehi _48836__119 (.L_HI(net119));
 sg13g2_tiehi _48835__120 (.L_HI(net120));
 sg13g2_tiehi _48834__121 (.L_HI(net121));
 sg13g2_tiehi _48833__122 (.L_HI(net122));
 sg13g2_tiehi _48832__123 (.L_HI(net123));
 sg13g2_tiehi _48831__124 (.L_HI(net124));
 sg13g2_tiehi _48830__125 (.L_HI(net125));
 sg13g2_tiehi _48829__126 (.L_HI(net126));
 sg13g2_tiehi _48828__127 (.L_HI(net127));
 sg13g2_tiehi _48827__128 (.L_HI(net128));
 sg13g2_tiehi _48826__129 (.L_HI(net129));
 sg13g2_tiehi _48825__130 (.L_HI(net130));
 sg13g2_tiehi _48824__131 (.L_HI(net131));
 sg13g2_tiehi _48823__132 (.L_HI(net132));
 sg13g2_tiehi _48822__133 (.L_HI(net133));
 sg13g2_tiehi _48821__134 (.L_HI(net134));
 sg13g2_tiehi _48820__135 (.L_HI(net135));
 sg13g2_tiehi _48819__136 (.L_HI(net136));
 sg13g2_tiehi _50034__137 (.L_HI(net137));
 sg13g2_tiehi _49806__138 (.L_HI(net138));
 sg13g2_tiehi _49805__139 (.L_HI(net139));
 sg13g2_tiehi _50033__140 (.L_HI(net140));
 sg13g2_tiehi _49804__141 (.L_HI(net141));
 sg13g2_tiehi _49803__142 (.L_HI(net142));
 sg13g2_tiehi _50032__143 (.L_HI(net143));
 sg13g2_tiehi _49802__144 (.L_HI(net144));
 sg13g2_tiehi _49801__145 (.L_HI(net145));
 sg13g2_tiehi _50031__146 (.L_HI(net146));
 sg13g2_tiehi _49800__147 (.L_HI(net147));
 sg13g2_tiehi _49799__148 (.L_HI(net148));
 sg13g2_tiehi _50030__149 (.L_HI(net149));
 sg13g2_tiehi _49798__150 (.L_HI(net150));
 sg13g2_tiehi _49797__151 (.L_HI(net151));
 sg13g2_tiehi _50029__152 (.L_HI(net152));
 sg13g2_tiehi _49796__153 (.L_HI(net153));
 sg13g2_tiehi _49795__154 (.L_HI(net154));
 sg13g2_tiehi _50028__155 (.L_HI(net155));
 sg13g2_tiehi _49794__156 (.L_HI(net156));
 sg13g2_tiehi _49793__157 (.L_HI(net157));
 sg13g2_tiehi _50027__158 (.L_HI(net158));
 sg13g2_tiehi _49792__159 (.L_HI(net159));
 sg13g2_tiehi _49791__160 (.L_HI(net160));
 sg13g2_tiehi _50026__161 (.L_HI(net161));
 sg13g2_tiehi _49790__162 (.L_HI(net162));
 sg13g2_tiehi _49789__163 (.L_HI(net163));
 sg13g2_tiehi _50025__164 (.L_HI(net164));
 sg13g2_tiehi _49788__165 (.L_HI(net165));
 sg13g2_tiehi _49787__166 (.L_HI(net166));
 sg13g2_tiehi _50024__167 (.L_HI(net167));
 sg13g2_tiehi _49786__168 (.L_HI(net168));
 sg13g2_tiehi _49785__169 (.L_HI(net169));
 sg13g2_tiehi _50023__170 (.L_HI(net170));
 sg13g2_tiehi _49784__171 (.L_HI(net171));
 sg13g2_tiehi _49783__172 (.L_HI(net172));
 sg13g2_tiehi _50022__173 (.L_HI(net173));
 sg13g2_tiehi _49782__174 (.L_HI(net174));
 sg13g2_tiehi _49781__175 (.L_HI(net175));
 sg13g2_tiehi _50021__176 (.L_HI(net176));
 sg13g2_tiehi _49780__177 (.L_HI(net177));
 sg13g2_tiehi _49779__178 (.L_HI(net178));
 sg13g2_tiehi _50020__179 (.L_HI(net179));
 sg13g2_tiehi _49778__180 (.L_HI(net180));
 sg13g2_tiehi _49777__181 (.L_HI(net181));
 sg13g2_tiehi _50019__182 (.L_HI(net182));
 sg13g2_tiehi _49776__183 (.L_HI(net183));
 sg13g2_tiehi _49775__184 (.L_HI(net184));
 sg13g2_tiehi _50018__185 (.L_HI(net185));
 sg13g2_tiehi _49774__186 (.L_HI(net186));
 sg13g2_tiehi _50123__187 (.L_HI(net187));
 sg13g2_tiehi _49773__188 (.L_HI(net188));
 sg13g2_tiehi _50017__189 (.L_HI(net189));
 sg13g2_tiehi _49772__190 (.L_HI(net190));
 sg13g2_tiehi _50146__191 (.L_HI(net191));
 sg13g2_tiehi _49771__192 (.L_HI(net192));
 sg13g2_tiehi _50016__193 (.L_HI(net193));
 sg13g2_tiehi _49770__194 (.L_HI(net194));
 sg13g2_tiehi _49769__195 (.L_HI(net195));
 sg13g2_tiehi _50015__196 (.L_HI(net196));
 sg13g2_tiehi _49768__197 (.L_HI(net197));
 sg13g2_tiehi _50145__198 (.L_HI(net198));
 sg13g2_tiehi _49767__199 (.L_HI(net199));
 sg13g2_tiehi _50014__200 (.L_HI(net200));
 sg13g2_tiehi _49766__201 (.L_HI(net201));
 sg13g2_tiehi _49765__202 (.L_HI(net202));
 sg13g2_tiehi _50013__203 (.L_HI(net203));
 sg13g2_tiehi _49764__204 (.L_HI(net204));
 sg13g2_tiehi _50144__205 (.L_HI(net205));
 sg13g2_tiehi _49763__206 (.L_HI(net206));
 sg13g2_tiehi _50012__207 (.L_HI(net207));
 sg13g2_tiehi _49762__208 (.L_HI(net208));
 sg13g2_tiehi _49761__209 (.L_HI(net209));
 sg13g2_tiehi _50011__210 (.L_HI(net210));
 sg13g2_tiehi _49760__211 (.L_HI(net211));
 sg13g2_tiehi _50143__212 (.L_HI(net212));
 sg13g2_tiehi _49759__213 (.L_HI(net213));
 sg13g2_tiehi _50010__214 (.L_HI(net214));
 sg13g2_tiehi _49758__215 (.L_HI(net215));
 sg13g2_tiehi _49757__216 (.L_HI(net216));
 sg13g2_tiehi _50009__217 (.L_HI(net217));
 sg13g2_tiehi _49756__218 (.L_HI(net218));
 sg13g2_tiehi _50142__219 (.L_HI(net219));
 sg13g2_tiehi _49755__220 (.L_HI(net220));
 sg13g2_tiehi _50008__221 (.L_HI(net221));
 sg13g2_tiehi _49754__222 (.L_HI(net222));
 sg13g2_tiehi _49753__223 (.L_HI(net223));
 sg13g2_tiehi _50007__224 (.L_HI(net224));
 sg13g2_tiehi _49752__225 (.L_HI(net225));
 sg13g2_tiehi _50141__226 (.L_HI(net226));
 sg13g2_tiehi _49751__227 (.L_HI(net227));
 sg13g2_tiehi _50006__228 (.L_HI(net228));
 sg13g2_tiehi _49750__229 (.L_HI(net229));
 sg13g2_tiehi _49749__230 (.L_HI(net230));
 sg13g2_tiehi _50005__231 (.L_HI(net231));
 sg13g2_tiehi _49748__232 (.L_HI(net232));
 sg13g2_tiehi _50140__233 (.L_HI(net233));
 sg13g2_tiehi _49747__234 (.L_HI(net234));
 sg13g2_tiehi _50004__235 (.L_HI(net235));
 sg13g2_tiehi _49746__236 (.L_HI(net236));
 sg13g2_tiehi _49745__237 (.L_HI(net237));
 sg13g2_tiehi _50003__238 (.L_HI(net238));
 sg13g2_tiehi _49744__239 (.L_HI(net239));
 sg13g2_tiehi _50139__240 (.L_HI(net240));
 sg13g2_tiehi _49743__241 (.L_HI(net241));
 sg13g2_tiehi _50002__242 (.L_HI(net242));
 sg13g2_tiehi _49742__243 (.L_HI(net243));
 sg13g2_tiehi _49741__244 (.L_HI(net244));
 sg13g2_tiehi _50001__245 (.L_HI(net245));
 sg13g2_tiehi _49740__246 (.L_HI(net246));
 sg13g2_tiehi _50138__247 (.L_HI(net247));
 sg13g2_tiehi _49739__248 (.L_HI(net248));
 sg13g2_tiehi _50000__249 (.L_HI(net249));
 sg13g2_tiehi _49738__250 (.L_HI(net250));
 sg13g2_tiehi _49737__251 (.L_HI(net251));
 sg13g2_tiehi _49999__252 (.L_HI(net252));
 sg13g2_tiehi _49736__253 (.L_HI(net253));
 sg13g2_tiehi _50137__254 (.L_HI(net254));
 sg13g2_tiehi _49735__255 (.L_HI(net255));
 sg13g2_tiehi _49998__256 (.L_HI(net256));
 sg13g2_tiehi _49734__257 (.L_HI(net257));
 sg13g2_tiehi _49733__258 (.L_HI(net258));
 sg13g2_tiehi _49997__259 (.L_HI(net259));
 sg13g2_tiehi _49732__260 (.L_HI(net260));
 sg13g2_tiehi _49731__261 (.L_HI(net261));
 sg13g2_tiehi _49996__262 (.L_HI(net262));
 sg13g2_tiehi _49730__263 (.L_HI(net263));
 sg13g2_tiehi _49729__264 (.L_HI(net264));
 sg13g2_tiehi _49995__265 (.L_HI(net265));
 sg13g2_tiehi _49728__266 (.L_HI(net266));
 sg13g2_tiehi _49727__267 (.L_HI(net267));
 sg13g2_tiehi _49994__268 (.L_HI(net268));
 sg13g2_tiehi _49726__269 (.L_HI(net269));
 sg13g2_tiehi _49725__270 (.L_HI(net270));
 sg13g2_tiehi _49993__271 (.L_HI(net271));
 sg13g2_tiehi _49724__272 (.L_HI(net272));
 sg13g2_tiehi _49723__273 (.L_HI(net273));
 sg13g2_tiehi _49992__274 (.L_HI(net274));
 sg13g2_tiehi _49722__275 (.L_HI(net275));
 sg13g2_tiehi _49721__276 (.L_HI(net276));
 sg13g2_tiehi _49991__277 (.L_HI(net277));
 sg13g2_tiehi _49720__278 (.L_HI(net278));
 sg13g2_tiehi _49719__279 (.L_HI(net279));
 sg13g2_tiehi _49990__280 (.L_HI(net280));
 sg13g2_tiehi _49718__281 (.L_HI(net281));
 sg13g2_tiehi _49717__282 (.L_HI(net282));
 sg13g2_tiehi _49989__283 (.L_HI(net283));
 sg13g2_tiehi _49716__284 (.L_HI(net284));
 sg13g2_tiehi _49715__285 (.L_HI(net285));
 sg13g2_tiehi _49988__286 (.L_HI(net286));
 sg13g2_tiehi _49714__287 (.L_HI(net287));
 sg13g2_tiehi _49713__288 (.L_HI(net288));
 sg13g2_tiehi _49987__289 (.L_HI(net289));
 sg13g2_tiehi _49712__290 (.L_HI(net290));
 sg13g2_tiehi _49711__291 (.L_HI(net291));
 sg13g2_tiehi _49986__292 (.L_HI(net292));
 sg13g2_tiehi _49710__293 (.L_HI(net293));
 sg13g2_tiehi _49709__294 (.L_HI(net294));
 sg13g2_tiehi _49985__295 (.L_HI(net295));
 sg13g2_tiehi _49708__296 (.L_HI(net296));
 sg13g2_tiehi _49707__297 (.L_HI(net297));
 sg13g2_tiehi _49984__298 (.L_HI(net298));
 sg13g2_tiehi _49706__299 (.L_HI(net299));
 sg13g2_tiehi _49705__300 (.L_HI(net300));
 sg13g2_tiehi _49983__301 (.L_HI(net301));
 sg13g2_tiehi _49704__302 (.L_HI(net302));
 sg13g2_tiehi _50122__303 (.L_HI(net303));
 sg13g2_tiehi _49703__304 (.L_HI(net304));
 sg13g2_tiehi _49982__305 (.L_HI(net305));
 sg13g2_tiehi _49702__306 (.L_HI(net306));
 sg13g2_tiehi _49701__307 (.L_HI(net307));
 sg13g2_tiehi _49981__308 (.L_HI(net308));
 sg13g2_tiehi _49700__309 (.L_HI(net309));
 sg13g2_tiehi _50121__310 (.L_HI(net310));
 sg13g2_tiehi _49699__311 (.L_HI(net311));
 sg13g2_tiehi _49980__312 (.L_HI(net312));
 sg13g2_tiehi _49698__313 (.L_HI(net313));
 sg13g2_tiehi _49697__314 (.L_HI(net314));
 sg13g2_tiehi _49979__315 (.L_HI(net315));
 sg13g2_tiehi _49696__316 (.L_HI(net316));
 sg13g2_tiehi _50120__317 (.L_HI(net317));
 sg13g2_tiehi _49695__318 (.L_HI(net318));
 sg13g2_tiehi _49978__319 (.L_HI(net319));
 sg13g2_tiehi _49694__320 (.L_HI(net320));
 sg13g2_tiehi _49693__321 (.L_HI(net321));
 sg13g2_tiehi _49977__322 (.L_HI(net322));
 sg13g2_tiehi _49692__323 (.L_HI(net323));
 sg13g2_tiehi _50119__324 (.L_HI(net324));
 sg13g2_tiehi _49691__325 (.L_HI(net325));
 sg13g2_tiehi _49976__326 (.L_HI(net326));
 sg13g2_tiehi _49690__327 (.L_HI(net327));
 sg13g2_tiehi _49689__328 (.L_HI(net328));
 sg13g2_tiehi _49975__329 (.L_HI(net329));
 sg13g2_tiehi _49688__330 (.L_HI(net330));
 sg13g2_tiehi _50118__331 (.L_HI(net331));
 sg13g2_tiehi _49687__332 (.L_HI(net332));
 sg13g2_tiehi _49974__333 (.L_HI(net333));
 sg13g2_tiehi _49686__334 (.L_HI(net334));
 sg13g2_tiehi _49685__335 (.L_HI(net335));
 sg13g2_tiehi _49973__336 (.L_HI(net336));
 sg13g2_tiehi _49684__337 (.L_HI(net337));
 sg13g2_tiehi _50117__338 (.L_HI(net338));
 sg13g2_tiehi _49683__339 (.L_HI(net339));
 sg13g2_tiehi _49972__340 (.L_HI(net340));
 sg13g2_tiehi _49682__341 (.L_HI(net341));
 sg13g2_tiehi _49681__342 (.L_HI(net342));
 sg13g2_tiehi _49971__343 (.L_HI(net343));
 sg13g2_tiehi _49680__344 (.L_HI(net344));
 sg13g2_tiehi _50116__345 (.L_HI(net345));
 sg13g2_tiehi _49679__346 (.L_HI(net346));
 sg13g2_tiehi _49970__347 (.L_HI(net347));
 sg13g2_tiehi _49678__348 (.L_HI(net348));
 sg13g2_tiehi _49677__349 (.L_HI(net349));
 sg13g2_tiehi _49969__350 (.L_HI(net350));
 sg13g2_tiehi _49676__351 (.L_HI(net351));
 sg13g2_tiehi _50115__352 (.L_HI(net352));
 sg13g2_tiehi _49675__353 (.L_HI(net353));
 sg13g2_tiehi _49968__354 (.L_HI(net354));
 sg13g2_tiehi _49674__355 (.L_HI(net355));
 sg13g2_tiehi _49673__356 (.L_HI(net356));
 sg13g2_tiehi _49967__357 (.L_HI(net357));
 sg13g2_tiehi _49672__358 (.L_HI(net358));
 sg13g2_tiehi _50114__359 (.L_HI(net359));
 sg13g2_tiehi _49671__360 (.L_HI(net360));
 sg13g2_tiehi _49966__361 (.L_HI(net361));
 sg13g2_tiehi _49670__362 (.L_HI(net362));
 sg13g2_tiehi _49669__363 (.L_HI(net363));
 sg13g2_tiehi _49965__364 (.L_HI(net364));
 sg13g2_tiehi _49668__365 (.L_HI(net365));
 sg13g2_tiehi _50113__366 (.L_HI(net366));
 sg13g2_tiehi _49667__367 (.L_HI(net367));
 sg13g2_tiehi _49964__368 (.L_HI(net368));
 sg13g2_tiehi _49666__369 (.L_HI(net369));
 sg13g2_tiehi _49665__370 (.L_HI(net370));
 sg13g2_tiehi _49963__371 (.L_HI(net371));
 sg13g2_tiehi _49664__372 (.L_HI(net372));
 sg13g2_tiehi _50112__373 (.L_HI(net373));
 sg13g2_tiehi _49663__374 (.L_HI(net374));
 sg13g2_tiehi _49962__375 (.L_HI(net375));
 sg13g2_tiehi _49662__376 (.L_HI(net376));
 sg13g2_tiehi _49661__377 (.L_HI(net377));
 sg13g2_tiehi _49961__378 (.L_HI(net378));
 sg13g2_tiehi _49660__379 (.L_HI(net379));
 sg13g2_tiehi _50111__380 (.L_HI(net380));
 sg13g2_tiehi _49659__381 (.L_HI(net381));
 sg13g2_tiehi _49960__382 (.L_HI(net382));
 sg13g2_tiehi _49658__383 (.L_HI(net383));
 sg13g2_tiehi _49657__384 (.L_HI(net384));
 sg13g2_tiehi _49959__385 (.L_HI(net385));
 sg13g2_tiehi _49656__386 (.L_HI(net386));
 sg13g2_tiehi _50110__387 (.L_HI(net387));
 sg13g2_tiehi _49655__388 (.L_HI(net388));
 sg13g2_tiehi _49958__389 (.L_HI(net389));
 sg13g2_tiehi _49654__390 (.L_HI(net390));
 sg13g2_tiehi _49653__391 (.L_HI(net391));
 sg13g2_tiehi _49957__392 (.L_HI(net392));
 sg13g2_tiehi _49652__393 (.L_HI(net393));
 sg13g2_tiehi _50109__394 (.L_HI(net394));
 sg13g2_tiehi _49651__395 (.L_HI(net395));
 sg13g2_tiehi _49956__396 (.L_HI(net396));
 sg13g2_tiehi _49650__397 (.L_HI(net397));
 sg13g2_tiehi _49649__398 (.L_HI(net398));
 sg13g2_tiehi _49955__399 (.L_HI(net399));
 sg13g2_tiehi _49648__400 (.L_HI(net400));
 sg13g2_tiehi _50108__401 (.L_HI(net401));
 sg13g2_tiehi _49647__402 (.L_HI(net402));
 sg13g2_tiehi _49954__403 (.L_HI(net403));
 sg13g2_tiehi _49646__404 (.L_HI(net404));
 sg13g2_tiehi _49645__405 (.L_HI(net405));
 sg13g2_tiehi _49953__406 (.L_HI(net406));
 sg13g2_tiehi _49644__407 (.L_HI(net407));
 sg13g2_tiehi _50107__408 (.L_HI(net408));
 sg13g2_tiehi _49643__409 (.L_HI(net409));
 sg13g2_tiehi _49952__410 (.L_HI(net410));
 sg13g2_tiehi _49642__411 (.L_HI(net411));
 sg13g2_tiehi _49641__412 (.L_HI(net412));
 sg13g2_tiehi _49951__413 (.L_HI(net413));
 sg13g2_tiehi _49640__414 (.L_HI(net414));
 sg13g2_tiehi _50106__415 (.L_HI(net415));
 sg13g2_tiehi _49639__416 (.L_HI(net416));
 sg13g2_tiehi _49950__417 (.L_HI(net417));
 sg13g2_tiehi _49638__418 (.L_HI(net418));
 sg13g2_tiehi _49637__419 (.L_HI(net419));
 sg13g2_tiehi _49949__420 (.L_HI(net420));
 sg13g2_tiehi _49636__421 (.L_HI(net421));
 sg13g2_tiehi _50105__422 (.L_HI(net422));
 sg13g2_tiehi _49635__423 (.L_HI(net423));
 sg13g2_tiehi _49948__424 (.L_HI(net424));
 sg13g2_tiehi _49634__425 (.L_HI(net425));
 sg13g2_tiehi _49633__426 (.L_HI(net426));
 sg13g2_tiehi _49947__427 (.L_HI(net427));
 sg13g2_tiehi _49632__428 (.L_HI(net428));
 sg13g2_tiehi _50104__429 (.L_HI(net429));
 sg13g2_tiehi _49631__430 (.L_HI(net430));
 sg13g2_tiehi _49946__431 (.L_HI(net431));
 sg13g2_tiehi _49630__432 (.L_HI(net432));
 sg13g2_tiehi _49629__433 (.L_HI(net433));
 sg13g2_tiehi _49945__434 (.L_HI(net434));
 sg13g2_tiehi _49628__435 (.L_HI(net435));
 sg13g2_tiehi _50103__436 (.L_HI(net436));
 sg13g2_tiehi _49627__437 (.L_HI(net437));
 sg13g2_tiehi _49944__438 (.L_HI(net438));
 sg13g2_tiehi _49626__439 (.L_HI(net439));
 sg13g2_tiehi _49625__440 (.L_HI(net440));
 sg13g2_tiehi _49943__441 (.L_HI(net441));
 sg13g2_tiehi _49624__442 (.L_HI(net442));
 sg13g2_tiehi _50102__443 (.L_HI(net443));
 sg13g2_tiehi _49623__444 (.L_HI(net444));
 sg13g2_tiehi _49942__445 (.L_HI(net445));
 sg13g2_tiehi _49622__446 (.L_HI(net446));
 sg13g2_tiehi _49621__447 (.L_HI(net447));
 sg13g2_tiehi _49941__448 (.L_HI(net448));
 sg13g2_tiehi _49620__449 (.L_HI(net449));
 sg13g2_tiehi _50101__450 (.L_HI(net450));
 sg13g2_tiehi _49619__451 (.L_HI(net451));
 sg13g2_tiehi _49940__452 (.L_HI(net452));
 sg13g2_tiehi _49618__453 (.L_HI(net453));
 sg13g2_tiehi _49617__454 (.L_HI(net454));
 sg13g2_tiehi _49939__455 (.L_HI(net455));
 sg13g2_tiehi _49616__456 (.L_HI(net456));
 sg13g2_tiehi _50100__457 (.L_HI(net457));
 sg13g2_tiehi _49615__458 (.L_HI(net458));
 sg13g2_tiehi _49938__459 (.L_HI(net459));
 sg13g2_tiehi _49614__460 (.L_HI(net460));
 sg13g2_tiehi _49613__461 (.L_HI(net461));
 sg13g2_tiehi _49937__462 (.L_HI(net462));
 sg13g2_tiehi _49612__463 (.L_HI(net463));
 sg13g2_tiehi _50099__464 (.L_HI(net464));
 sg13g2_tiehi _49611__465 (.L_HI(net465));
 sg13g2_tiehi _49936__466 (.L_HI(net466));
 sg13g2_tiehi _49610__467 (.L_HI(net467));
 sg13g2_tiehi _49353__468 (.L_HI(net468));
 sg13g2_tiehi _49935__469 (.L_HI(net469));
 sg13g2_tiehi _49352__470 (.L_HI(net470));
 sg13g2_tiehi _50098__471 (.L_HI(net471));
 sg13g2_tiehi _49351__472 (.L_HI(net472));
 sg13g2_tiehi _49934__473 (.L_HI(net473));
 sg13g2_tiehi _49350__474 (.L_HI(net474));
 sg13g2_tiehi _49349__475 (.L_HI(net475));
 sg13g2_tiehi _49933__476 (.L_HI(net476));
 sg13g2_tiehi _49348__477 (.L_HI(net477));
 sg13g2_tiehi _50097__478 (.L_HI(net478));
 sg13g2_tiehi _49347__479 (.L_HI(net479));
 sg13g2_tiehi _49932__480 (.L_HI(net480));
 sg13g2_tiehi _49346__481 (.L_HI(net481));
 sg13g2_tiehi _49345__482 (.L_HI(net482));
 sg13g2_tiehi _49931__483 (.L_HI(net483));
 sg13g2_tiehi _49344__484 (.L_HI(net484));
 sg13g2_tiehi _50096__485 (.L_HI(net485));
 sg13g2_tiehi _49343__486 (.L_HI(net486));
 sg13g2_tiehi _49930__487 (.L_HI(net487));
 sg13g2_tiehi _49342__488 (.L_HI(net488));
 sg13g2_tiehi _49341__489 (.L_HI(net489));
 sg13g2_tiehi _49929__490 (.L_HI(net490));
 sg13g2_tiehi _49340__491 (.L_HI(net491));
 sg13g2_tiehi _50095__492 (.L_HI(net492));
 sg13g2_tiehi _49339__493 (.L_HI(net493));
 sg13g2_tiehi _49928__494 (.L_HI(net494));
 sg13g2_tiehi _49338__495 (.L_HI(net495));
 sg13g2_tiehi _49337__496 (.L_HI(net496));
 sg13g2_tiehi _49927__497 (.L_HI(net497));
 sg13g2_tiehi _49336__498 (.L_HI(net498));
 sg13g2_tiehi _50094__499 (.L_HI(net499));
 sg13g2_tiehi _49335__500 (.L_HI(net500));
 sg13g2_tiehi _49926__501 (.L_HI(net501));
 sg13g2_tiehi _49334__502 (.L_HI(net502));
 sg13g2_tiehi _49333__503 (.L_HI(net503));
 sg13g2_tiehi _49925__504 (.L_HI(net504));
 sg13g2_tiehi _49332__505 (.L_HI(net505));
 sg13g2_tiehi _50093__506 (.L_HI(net506));
 sg13g2_tiehi _49331__507 (.L_HI(net507));
 sg13g2_tiehi _49924__508 (.L_HI(net508));
 sg13g2_tiehi _49330__509 (.L_HI(net509));
 sg13g2_tiehi _49329__510 (.L_HI(net510));
 sg13g2_tiehi _49923__511 (.L_HI(net511));
 sg13g2_tiehi _49328__512 (.L_HI(net512));
 sg13g2_tiehi _50092__513 (.L_HI(net513));
 sg13g2_tiehi _49327__514 (.L_HI(net514));
 sg13g2_tiehi _49922__515 (.L_HI(net515));
 sg13g2_tiehi _49326__516 (.L_HI(net516));
 sg13g2_tiehi _49325__517 (.L_HI(net517));
 sg13g2_tiehi _49921__518 (.L_HI(net518));
 sg13g2_tiehi _49324__519 (.L_HI(net519));
 sg13g2_tiehi _50091__520 (.L_HI(net520));
 sg13g2_tiehi _49323__521 (.L_HI(net521));
 sg13g2_tiehi _49920__522 (.L_HI(net522));
 sg13g2_tiehi _49322__523 (.L_HI(net523));
 sg13g2_tiehi _49321__524 (.L_HI(net524));
 sg13g2_tiehi _49919__525 (.L_HI(net525));
 sg13g2_tiehi _49320__526 (.L_HI(net526));
 sg13g2_tiehi _50090__527 (.L_HI(net527));
 sg13g2_tiehi _49319__528 (.L_HI(net528));
 sg13g2_tiehi _49918__529 (.L_HI(net529));
 sg13g2_tiehi _49318__530 (.L_HI(net530));
 sg13g2_tiehi _49317__531 (.L_HI(net531));
 sg13g2_tiehi _49917__532 (.L_HI(net532));
 sg13g2_tiehi _49316__533 (.L_HI(net533));
 sg13g2_tiehi _50089__534 (.L_HI(net534));
 sg13g2_tiehi _49315__535 (.L_HI(net535));
 sg13g2_tiehi _49916__536 (.L_HI(net536));
 sg13g2_tiehi _49314__537 (.L_HI(net537));
 sg13g2_tiehi _49313__538 (.L_HI(net538));
 sg13g2_tiehi _49915__539 (.L_HI(net539));
 sg13g2_tiehi _49312__540 (.L_HI(net540));
 sg13g2_tiehi _50088__541 (.L_HI(net541));
 sg13g2_tiehi _49311__542 (.L_HI(net542));
 sg13g2_tiehi _49914__543 (.L_HI(net543));
 sg13g2_tiehi _49310__544 (.L_HI(net544));
 sg13g2_tiehi _49309__545 (.L_HI(net545));
 sg13g2_tiehi _49913__546 (.L_HI(net546));
 sg13g2_tiehi _49308__547 (.L_HI(net547));
 sg13g2_tiehi _50087__548 (.L_HI(net548));
 sg13g2_tiehi _49307__549 (.L_HI(net549));
 sg13g2_tiehi _49912__550 (.L_HI(net550));
 sg13g2_tiehi _49306__551 (.L_HI(net551));
 sg13g2_tiehi _49305__552 (.L_HI(net552));
 sg13g2_tiehi _49911__553 (.L_HI(net553));
 sg13g2_tiehi _49304__554 (.L_HI(net554));
 sg13g2_tiehi _50086__555 (.L_HI(net555));
 sg13g2_tiehi _49303__556 (.L_HI(net556));
 sg13g2_tiehi _49910__557 (.L_HI(net557));
 sg13g2_tiehi _49302__558 (.L_HI(net558));
 sg13g2_tiehi _49301__559 (.L_HI(net559));
 sg13g2_tiehi _49909__560 (.L_HI(net560));
 sg13g2_tiehi _49300__561 (.L_HI(net561));
 sg13g2_tiehi _50085__562 (.L_HI(net562));
 sg13g2_tiehi _49299__563 (.L_HI(net563));
 sg13g2_tiehi _49908__564 (.L_HI(net564));
 sg13g2_tiehi _49298__565 (.L_HI(net565));
 sg13g2_tiehi _49297__566 (.L_HI(net566));
 sg13g2_tiehi _49907__567 (.L_HI(net567));
 sg13g2_tiehi _49296__568 (.L_HI(net568));
 sg13g2_tiehi _50084__569 (.L_HI(net569));
 sg13g2_tiehi _49295__570 (.L_HI(net570));
 sg13g2_tiehi _49906__571 (.L_HI(net571));
 sg13g2_tiehi _49294__572 (.L_HI(net572));
 sg13g2_tiehi _49293__573 (.L_HI(net573));
 sg13g2_tiehi _49905__574 (.L_HI(net574));
 sg13g2_tiehi _49292__575 (.L_HI(net575));
 sg13g2_tiehi _50083__576 (.L_HI(net576));
 sg13g2_tiehi _49291__577 (.L_HI(net577));
 sg13g2_tiehi _49904__578 (.L_HI(net578));
 sg13g2_tiehi _49290__579 (.L_HI(net579));
 sg13g2_tiehi _49289__580 (.L_HI(net580));
 sg13g2_tiehi _49903__581 (.L_HI(net581));
 sg13g2_tiehi _49288__582 (.L_HI(net582));
 sg13g2_tiehi _50082__583 (.L_HI(net583));
 sg13g2_tiehi _49287__584 (.L_HI(net584));
 sg13g2_tiehi _49902__585 (.L_HI(net585));
 sg13g2_tiehi _49286__586 (.L_HI(net586));
 sg13g2_tiehi _49285__587 (.L_HI(net587));
 sg13g2_tiehi _49901__588 (.L_HI(net588));
 sg13g2_tiehi _49284__589 (.L_HI(net589));
 sg13g2_tiehi _50081__590 (.L_HI(net590));
 sg13g2_tiehi _49283__591 (.L_HI(net591));
 sg13g2_tiehi _49900__592 (.L_HI(net592));
 sg13g2_tiehi _49282__593 (.L_HI(net593));
 sg13g2_tiehi _49281__594 (.L_HI(net594));
 sg13g2_tiehi _49899__595 (.L_HI(net595));
 sg13g2_tiehi _49280__596 (.L_HI(net596));
 sg13g2_tiehi _50080__597 (.L_HI(net597));
 sg13g2_tiehi _49279__598 (.L_HI(net598));
 sg13g2_tiehi _49898__599 (.L_HI(net599));
 sg13g2_tiehi _49278__600 (.L_HI(net600));
 sg13g2_tiehi _49277__601 (.L_HI(net601));
 sg13g2_tiehi _49897__602 (.L_HI(net602));
 sg13g2_tiehi _49276__603 (.L_HI(net603));
 sg13g2_tiehi _50079__604 (.L_HI(net604));
 sg13g2_tiehi _49275__605 (.L_HI(net605));
 sg13g2_tiehi _49896__606 (.L_HI(net606));
 sg13g2_tiehi _49274__607 (.L_HI(net607));
 sg13g2_tiehi _49273__608 (.L_HI(net608));
 sg13g2_tiehi _49895__609 (.L_HI(net609));
 sg13g2_tiehi _49272__610 (.L_HI(net610));
 sg13g2_tiehi _50078__611 (.L_HI(net611));
 sg13g2_tiehi _49271__612 (.L_HI(net612));
 sg13g2_tiehi _49894__613 (.L_HI(net613));
 sg13g2_tiehi _49270__614 (.L_HI(net614));
 sg13g2_tiehi _49269__615 (.L_HI(net615));
 sg13g2_tiehi _49893__616 (.L_HI(net616));
 sg13g2_tiehi _49268__617 (.L_HI(net617));
 sg13g2_tiehi _50077__618 (.L_HI(net618));
 sg13g2_tiehi _49267__619 (.L_HI(net619));
 sg13g2_tiehi _49892__620 (.L_HI(net620));
 sg13g2_tiehi _49266__621 (.L_HI(net621));
 sg13g2_tiehi _49265__622 (.L_HI(net622));
 sg13g2_tiehi _49891__623 (.L_HI(net623));
 sg13g2_tiehi _49264__624 (.L_HI(net624));
 sg13g2_tiehi _50076__625 (.L_HI(net625));
 sg13g2_tiehi _49263__626 (.L_HI(net626));
 sg13g2_tiehi _49890__627 (.L_HI(net627));
 sg13g2_tiehi _49262__628 (.L_HI(net628));
 sg13g2_tiehi _49261__629 (.L_HI(net629));
 sg13g2_tiehi _49889__630 (.L_HI(net630));
 sg13g2_tiehi _49260__631 (.L_HI(net631));
 sg13g2_tiehi _50075__632 (.L_HI(net632));
 sg13g2_tiehi _49259__633 (.L_HI(net633));
 sg13g2_tiehi _49888__634 (.L_HI(net634));
 sg13g2_tiehi _49258__635 (.L_HI(net635));
 sg13g2_tiehi _49257__636 (.L_HI(net636));
 sg13g2_tiehi _49887__637 (.L_HI(net637));
 sg13g2_tiehi _49256__638 (.L_HI(net638));
 sg13g2_tiehi _50074__639 (.L_HI(net639));
 sg13g2_tiehi _49255__640 (.L_HI(net640));
 sg13g2_tiehi _49886__641 (.L_HI(net641));
 sg13g2_tiehi _49254__642 (.L_HI(net642));
 sg13g2_tiehi _49253__643 (.L_HI(net643));
 sg13g2_tiehi _49885__644 (.L_HI(net644));
 sg13g2_tiehi _49252__645 (.L_HI(net645));
 sg13g2_tiehi _50073__646 (.L_HI(net646));
 sg13g2_tiehi _49251__647 (.L_HI(net647));
 sg13g2_tiehi _49884__648 (.L_HI(net648));
 sg13g2_tiehi _49250__649 (.L_HI(net649));
 sg13g2_tiehi _49249__650 (.L_HI(net650));
 sg13g2_tiehi _49883__651 (.L_HI(net651));
 sg13g2_tiehi _49248__652 (.L_HI(net652));
 sg13g2_tiehi _50072__653 (.L_HI(net653));
 sg13g2_tiehi _49247__654 (.L_HI(net654));
 sg13g2_tiehi _49882__655 (.L_HI(net655));
 sg13g2_tiehi _49246__656 (.L_HI(net656));
 sg13g2_tiehi _49245__657 (.L_HI(net657));
 sg13g2_tiehi _49881__658 (.L_HI(net658));
 sg13g2_tiehi _49244__659 (.L_HI(net659));
 sg13g2_tiehi _50071__660 (.L_HI(net660));
 sg13g2_tiehi _49243__661 (.L_HI(net661));
 sg13g2_tiehi _49880__662 (.L_HI(net662));
 sg13g2_tiehi _49242__663 (.L_HI(net663));
 sg13g2_tiehi _49241__664 (.L_HI(net664));
 sg13g2_tiehi _49879__665 (.L_HI(net665));
 sg13g2_tiehi _49240__666 (.L_HI(net666));
 sg13g2_tiehi _50070__667 (.L_HI(net667));
 sg13g2_tiehi _49239__668 (.L_HI(net668));
 sg13g2_tiehi _49878__669 (.L_HI(net669));
 sg13g2_tiehi _49238__670 (.L_HI(net670));
 sg13g2_tiehi _49237__671 (.L_HI(net671));
 sg13g2_tiehi _49877__672 (.L_HI(net672));
 sg13g2_tiehi _49236__673 (.L_HI(net673));
 sg13g2_tiehi _50069__674 (.L_HI(net674));
 sg13g2_tiehi _49235__675 (.L_HI(net675));
 sg13g2_tiehi _49876__676 (.L_HI(net676));
 sg13g2_tiehi _49234__677 (.L_HI(net677));
 sg13g2_tiehi _49233__678 (.L_HI(net678));
 sg13g2_tiehi _49875__679 (.L_HI(net679));
 sg13g2_tiehi _49232__680 (.L_HI(net680));
 sg13g2_tiehi _50068__681 (.L_HI(net681));
 sg13g2_tiehi _49231__682 (.L_HI(net682));
 sg13g2_tiehi _49874__683 (.L_HI(net683));
 sg13g2_tiehi _49230__684 (.L_HI(net684));
 sg13g2_tiehi _49229__685 (.L_HI(net685));
 sg13g2_tiehi _49873__686 (.L_HI(net686));
 sg13g2_tiehi _49228__687 (.L_HI(net687));
 sg13g2_tiehi _50067__688 (.L_HI(net688));
 sg13g2_tiehi _49227__689 (.L_HI(net689));
 sg13g2_tiehi _49872__690 (.L_HI(net690));
 sg13g2_tiehi _49226__691 (.L_HI(net691));
 sg13g2_tiehi _49225__692 (.L_HI(net692));
 sg13g2_tiehi _49871__693 (.L_HI(net693));
 sg13g2_tiehi _49224__694 (.L_HI(net694));
 sg13g2_tiehi _50066__695 (.L_HI(net695));
 sg13g2_tiehi _49223__696 (.L_HI(net696));
 sg13g2_tiehi _49870__697 (.L_HI(net697));
 sg13g2_tiehi _49222__698 (.L_HI(net698));
 sg13g2_tiehi _49221__699 (.L_HI(net699));
 sg13g2_tiehi _49869__700 (.L_HI(net700));
 sg13g2_tiehi _49220__701 (.L_HI(net701));
 sg13g2_tiehi _50065__702 (.L_HI(net702));
 sg13g2_tiehi _49219__703 (.L_HI(net703));
 sg13g2_tiehi _49868__704 (.L_HI(net704));
 sg13g2_tiehi _49218__705 (.L_HI(net705));
 sg13g2_tiehi _49217__706 (.L_HI(net706));
 sg13g2_tiehi _49867__707 (.L_HI(net707));
 sg13g2_tiehi _49216__708 (.L_HI(net708));
 sg13g2_tiehi _50064__709 (.L_HI(net709));
 sg13g2_tiehi _49215__710 (.L_HI(net710));
 sg13g2_tiehi _49866__711 (.L_HI(net711));
 sg13g2_tiehi _49214__712 (.L_HI(net712));
 sg13g2_tiehi _49213__713 (.L_HI(net713));
 sg13g2_tiehi _49865__714 (.L_HI(net714));
 sg13g2_tiehi _49212__715 (.L_HI(net715));
 sg13g2_tiehi _50063__716 (.L_HI(net716));
 sg13g2_tiehi _49211__717 (.L_HI(net717));
 sg13g2_tiehi _49864__718 (.L_HI(net718));
 sg13g2_tiehi _49210__719 (.L_HI(net719));
 sg13g2_tiehi _49209__720 (.L_HI(net720));
 sg13g2_tiehi _49863__721 (.L_HI(net721));
 sg13g2_tiehi _49208__722 (.L_HI(net722));
 sg13g2_tiehi _50062__723 (.L_HI(net723));
 sg13g2_tiehi _49207__724 (.L_HI(net724));
 sg13g2_tiehi _49862__725 (.L_HI(net725));
 sg13g2_tiehi _49206__726 (.L_HI(net726));
 sg13g2_tiehi _49205__727 (.L_HI(net727));
 sg13g2_tiehi _49861__728 (.L_HI(net728));
 sg13g2_tiehi _49204__729 (.L_HI(net729));
 sg13g2_tiehi _50061__730 (.L_HI(net730));
 sg13g2_tiehi _49203__731 (.L_HI(net731));
 sg13g2_tiehi _49860__732 (.L_HI(net732));
 sg13g2_tiehi _49202__733 (.L_HI(net733));
 sg13g2_tiehi _49201__734 (.L_HI(net734));
 sg13g2_tiehi _49859__735 (.L_HI(net735));
 sg13g2_tiehi _49200__736 (.L_HI(net736));
 sg13g2_tiehi _50060__737 (.L_HI(net737));
 sg13g2_tiehi _49199__738 (.L_HI(net738));
 sg13g2_tiehi _49858__739 (.L_HI(net739));
 sg13g2_tiehi _49198__740 (.L_HI(net740));
 sg13g2_tiehi _49197__741 (.L_HI(net741));
 sg13g2_tiehi _49857__742 (.L_HI(net742));
 sg13g2_tiehi _49196__743 (.L_HI(net743));
 sg13g2_tiehi _50059__744 (.L_HI(net744));
 sg13g2_tiehi _49195__745 (.L_HI(net745));
 sg13g2_tiehi _49856__746 (.L_HI(net746));
 sg13g2_tiehi _49194__747 (.L_HI(net747));
 sg13g2_tiehi _49193__748 (.L_HI(net748));
 sg13g2_tiehi _49855__749 (.L_HI(net749));
 sg13g2_tiehi _49192__750 (.L_HI(net750));
 sg13g2_tiehi _50058__751 (.L_HI(net751));
 sg13g2_tiehi _49191__752 (.L_HI(net752));
 sg13g2_tiehi _49854__753 (.L_HI(net753));
 sg13g2_tiehi _49190__754 (.L_HI(net754));
 sg13g2_tiehi _49189__755 (.L_HI(net755));
 sg13g2_tiehi _49853__756 (.L_HI(net756));
 sg13g2_tiehi _49188__757 (.L_HI(net757));
 sg13g2_tiehi _50057__758 (.L_HI(net758));
 sg13g2_tiehi _49187__759 (.L_HI(net759));
 sg13g2_tiehi _49852__760 (.L_HI(net760));
 sg13g2_tiehi _49186__761 (.L_HI(net761));
 sg13g2_tiehi _49185__762 (.L_HI(net762));
 sg13g2_tiehi _49851__763 (.L_HI(net763));
 sg13g2_tiehi _49184__764 (.L_HI(net764));
 sg13g2_tiehi _50056__765 (.L_HI(net765));
 sg13g2_tiehi _49183__766 (.L_HI(net766));
 sg13g2_tiehi _49850__767 (.L_HI(net767));
 sg13g2_tiehi _49182__768 (.L_HI(net768));
 sg13g2_tiehi _49181__769 (.L_HI(net769));
 sg13g2_tiehi _49849__770 (.L_HI(net770));
 sg13g2_tiehi _49180__771 (.L_HI(net771));
 sg13g2_tiehi _50055__772 (.L_HI(net772));
 sg13g2_tiehi _49179__773 (.L_HI(net773));
 sg13g2_tiehi _49848__774 (.L_HI(net774));
 sg13g2_tiehi _49178__775 (.L_HI(net775));
 sg13g2_tiehi _49177__776 (.L_HI(net776));
 sg13g2_tiehi _49847__777 (.L_HI(net777));
 sg13g2_tiehi _49176__778 (.L_HI(net778));
 sg13g2_tiehi _50054__779 (.L_HI(net779));
 sg13g2_tiehi _49175__780 (.L_HI(net780));
 sg13g2_tiehi _49846__781 (.L_HI(net781));
 sg13g2_tiehi _49174__782 (.L_HI(net782));
 sg13g2_tiehi _49173__783 (.L_HI(net783));
 sg13g2_tiehi _49845__784 (.L_HI(net784));
 sg13g2_tiehi _49172__785 (.L_HI(net785));
 sg13g2_tiehi _50053__786 (.L_HI(net786));
 sg13g2_tiehi _49171__787 (.L_HI(net787));
 sg13g2_tiehi _49844__788 (.L_HI(net788));
 sg13g2_tiehi _49170__789 (.L_HI(net789));
 sg13g2_tiehi _49169__790 (.L_HI(net790));
 sg13g2_tiehi _49843__791 (.L_HI(net791));
 sg13g2_tiehi _49168__792 (.L_HI(net792));
 sg13g2_tiehi _50052__793 (.L_HI(net793));
 sg13g2_tiehi _49167__794 (.L_HI(net794));
 sg13g2_tiehi _49842__795 (.L_HI(net795));
 sg13g2_tiehi _49166__796 (.L_HI(net796));
 sg13g2_tiehi _49165__797 (.L_HI(net797));
 sg13g2_tiehi _49841__798 (.L_HI(net798));
 sg13g2_tiehi _49164__799 (.L_HI(net799));
 sg13g2_tiehi _50051__800 (.L_HI(net800));
 sg13g2_tiehi _49163__801 (.L_HI(net801));
 sg13g2_tiehi _49840__802 (.L_HI(net802));
 sg13g2_tiehi _49162__803 (.L_HI(net803));
 sg13g2_tiehi _49161__804 (.L_HI(net804));
 sg13g2_tiehi _49839__805 (.L_HI(net805));
 sg13g2_tiehi _49160__806 (.L_HI(net806));
 sg13g2_tiehi _50050__807 (.L_HI(net807));
 sg13g2_tiehi _49159__808 (.L_HI(net808));
 sg13g2_tiehi _49838__809 (.L_HI(net809));
 sg13g2_tiehi _49158__810 (.L_HI(net810));
 sg13g2_tiehi _49157__811 (.L_HI(net811));
 sg13g2_tiehi _49837__812 (.L_HI(net812));
 sg13g2_tiehi _49156__813 (.L_HI(net813));
 sg13g2_tiehi _50049__814 (.L_HI(net814));
 sg13g2_tiehi _49155__815 (.L_HI(net815));
 sg13g2_tiehi _49836__816 (.L_HI(net816));
 sg13g2_tiehi _49154__817 (.L_HI(net817));
 sg13g2_tiehi _49153__818 (.L_HI(net818));
 sg13g2_tiehi _49835__819 (.L_HI(net819));
 sg13g2_tiehi _49152__820 (.L_HI(net820));
 sg13g2_tiehi _50048__821 (.L_HI(net821));
 sg13g2_tiehi _49151__822 (.L_HI(net822));
 sg13g2_tiehi _49834__823 (.L_HI(net823));
 sg13g2_tiehi _49150__824 (.L_HI(net824));
 sg13g2_tiehi _49149__825 (.L_HI(net825));
 sg13g2_tiehi _49833__826 (.L_HI(net826));
 sg13g2_tiehi _49148__827 (.L_HI(net827));
 sg13g2_tiehi _50047__828 (.L_HI(net828));
 sg13g2_tiehi _49147__829 (.L_HI(net829));
 sg13g2_tiehi _49832__830 (.L_HI(net830));
 sg13g2_tiehi _49146__831 (.L_HI(net831));
 sg13g2_tiehi _49145__832 (.L_HI(net832));
 sg13g2_tiehi _49831__833 (.L_HI(net833));
 sg13g2_tiehi _49144__834 (.L_HI(net834));
 sg13g2_tiehi _50046__835 (.L_HI(net835));
 sg13g2_tiehi _49143__836 (.L_HI(net836));
 sg13g2_tiehi _49830__837 (.L_HI(net837));
 sg13g2_tiehi _49142__838 (.L_HI(net838));
 sg13g2_tiehi _49141__839 (.L_HI(net839));
 sg13g2_tiehi _49829__840 (.L_HI(net840));
 sg13g2_tiehi _49140__841 (.L_HI(net841));
 sg13g2_tiehi _50045__842 (.L_HI(net842));
 sg13g2_tiehi _49139__843 (.L_HI(net843));
 sg13g2_tiehi _49828__844 (.L_HI(net844));
 sg13g2_tiehi _49138__845 (.L_HI(net845));
 sg13g2_tiehi _49137__846 (.L_HI(net846));
 sg13g2_tiehi _49827__847 (.L_HI(net847));
 sg13g2_tiehi _49136__848 (.L_HI(net848));
 sg13g2_tiehi _50044__849 (.L_HI(net849));
 sg13g2_tiehi _49135__850 (.L_HI(net850));
 sg13g2_tiehi _49826__851 (.L_HI(net851));
 sg13g2_tiehi _49134__852 (.L_HI(net852));
 sg13g2_tiehi _49133__853 (.L_HI(net853));
 sg13g2_tiehi _49825__854 (.L_HI(net854));
 sg13g2_tiehi _49132__855 (.L_HI(net855));
 sg13g2_tiehi _50043__856 (.L_HI(net856));
 sg13g2_tiehi _49131__857 (.L_HI(net857));
 sg13g2_tiehi _49824__858 (.L_HI(net858));
 sg13g2_tiehi _49130__859 (.L_HI(net859));
 sg13g2_tiehi _49129__860 (.L_HI(net860));
 sg13g2_tiehi _49823__861 (.L_HI(net861));
 sg13g2_tiehi _49128__862 (.L_HI(net862));
 sg13g2_tiehi _50042__863 (.L_HI(net863));
 sg13g2_tiehi _49127__864 (.L_HI(net864));
 sg13g2_tiehi _49822__865 (.L_HI(net865));
 sg13g2_tiehi _49126__866 (.L_HI(net866));
 sg13g2_tiehi _49125__867 (.L_HI(net867));
 sg13g2_tiehi _49821__868 (.L_HI(net868));
 sg13g2_tiehi _49124__869 (.L_HI(net869));
 sg13g2_tiehi _50041__870 (.L_HI(net870));
 sg13g2_tiehi _49123__871 (.L_HI(net871));
 sg13g2_tiehi _49820__872 (.L_HI(net872));
 sg13g2_tiehi _49122__873 (.L_HI(net873));
 sg13g2_tiehi _49121__874 (.L_HI(net874));
 sg13g2_tiehi _49819__875 (.L_HI(net875));
 sg13g2_tiehi _49120__876 (.L_HI(net876));
 sg13g2_tiehi _50040__877 (.L_HI(net877));
 sg13g2_tiehi _49119__878 (.L_HI(net878));
 sg13g2_tiehi _49818__879 (.L_HI(net879));
 sg13g2_tiehi _49118__880 (.L_HI(net880));
 sg13g2_tiehi _49117__881 (.L_HI(net881));
 sg13g2_tiehi _49817__882 (.L_HI(net882));
 sg13g2_tiehi _49116__883 (.L_HI(net883));
 sg13g2_tiehi _50039__884 (.L_HI(net884));
 sg13g2_tiehi _49115__885 (.L_HI(net885));
 sg13g2_tiehi _49816__886 (.L_HI(net886));
 sg13g2_tiehi _49114__887 (.L_HI(net887));
 sg13g2_tiehi _49113__888 (.L_HI(net888));
 sg13g2_tiehi _49815__889 (.L_HI(net889));
 sg13g2_tiehi _49112__890 (.L_HI(net890));
 sg13g2_tiehi _50038__891 (.L_HI(net891));
 sg13g2_tiehi _49111__892 (.L_HI(net892));
 sg13g2_tiehi _49814__893 (.L_HI(net893));
 sg13g2_tiehi _49110__894 (.L_HI(net894));
 sg13g2_tiehi _49109__895 (.L_HI(net895));
 sg13g2_tiehi _49813__896 (.L_HI(net896));
 sg13g2_tiehi _49108__897 (.L_HI(net897));
 sg13g2_tiehi _50037__898 (.L_HI(net898));
 sg13g2_tiehi _49107__899 (.L_HI(net899));
 sg13g2_tiehi _49812__900 (.L_HI(net900));
 sg13g2_tiehi _49106__901 (.L_HI(net901));
 sg13g2_tiehi _49105__902 (.L_HI(net902));
 sg13g2_tiehi _49811__903 (.L_HI(net903));
 sg13g2_tiehi _49104__904 (.L_HI(net904));
 sg13g2_tiehi _50036__905 (.L_HI(net905));
 sg13g2_tiehi _49103__906 (.L_HI(net906));
 sg13g2_tiehi _49810__907 (.L_HI(net907));
 sg13g2_tiehi _49102__908 (.L_HI(net908));
 sg13g2_tiehi _49101__909 (.L_HI(net909));
 sg13g2_tiehi _49809__910 (.L_HI(net910));
 sg13g2_tiehi _49100__911 (.L_HI(net911));
 sg13g2_tiehi _50035__912 (.L_HI(net912));
 sg13g2_tiehi _49099__913 (.L_HI(net913));
 sg13g2_tiehi _49808__914 (.L_HI(net914));
 sg13g2_tiehi _49098__915 (.L_HI(net915));
 sg13g2_tiehi _49097__916 (.L_HI(net916));
 sg13g2_tiehi _49807__917 (.L_HI(net917));
 sg13g2_tiehi _49075__918 (.L_HI(net918));
 sg13g2_tiehi _49074__919 (.L_HI(net919));
 sg13g2_tiehi _49073__920 (.L_HI(net920));
 sg13g2_tiehi _49072__921 (.L_HI(net921));
 sg13g2_tiehi _49071__922 (.L_HI(net922));
 sg13g2_tiehi _49070__923 (.L_HI(net923));
 sg13g2_tiehi _49069__924 (.L_HI(net924));
 sg13g2_tiehi _49068__925 (.L_HI(net925));
 sg13g2_tiehi _49067__926 (.L_HI(net926));
 sg13g2_tiehi _49066__927 (.L_HI(net927));
 sg13g2_tiehi _49065__928 (.L_HI(net928));
 sg13g2_tiehi _49064__929 (.L_HI(net929));
 sg13g2_tiehi _49063__930 (.L_HI(net930));
 sg13g2_tiehi _49062__931 (.L_HI(net931));
 sg13g2_tiehi _49061__932 (.L_HI(net932));
 sg13g2_tiehi _49060__933 (.L_HI(net933));
 sg13g2_tiehi _49059__934 (.L_HI(net934));
 sg13g2_tiehi _49058__935 (.L_HI(net935));
 sg13g2_tiehi _49057__936 (.L_HI(net936));
 sg13g2_tiehi _49056__937 (.L_HI(net937));
 sg13g2_tiehi _49055__938 (.L_HI(net938));
 sg13g2_tiehi _49054__939 (.L_HI(net939));
 sg13g2_tiehi _49053__940 (.L_HI(net940));
 sg13g2_tiehi _49052__941 (.L_HI(net941));
 sg13g2_tiehi _49051__942 (.L_HI(net942));
 sg13g2_tiehi _49050__943 (.L_HI(net943));
 sg13g2_tiehi _49049__944 (.L_HI(net944));
 sg13g2_tiehi _49048__945 (.L_HI(net945));
 sg13g2_tiehi _49047__946 (.L_HI(net946));
 sg13g2_tiehi _49046__947 (.L_HI(net947));
 sg13g2_tiehi _49045__948 (.L_HI(net948));
 sg13g2_tiehi _49044__949 (.L_HI(net949));
 sg13g2_tiehi _49043__950 (.L_HI(net950));
 sg13g2_tiehi _49042__951 (.L_HI(net951));
 sg13g2_tiehi _49041__952 (.L_HI(net952));
 sg13g2_tiehi _49040__953 (.L_HI(net953));
 sg13g2_tiehi _49039__954 (.L_HI(net954));
 sg13g2_tiehi _49038__955 (.L_HI(net955));
 sg13g2_tiehi _49037__956 (.L_HI(net956));
 sg13g2_tiehi _49036__957 (.L_HI(net957));
 sg13g2_tiehi _49035__958 (.L_HI(net958));
 sg13g2_tiehi _49034__959 (.L_HI(net959));
 sg13g2_tiehi _49033__960 (.L_HI(net960));
 sg13g2_tiehi _49032__961 (.L_HI(net961));
 sg13g2_tiehi _49031__962 (.L_HI(net962));
 sg13g2_tiehi _49030__963 (.L_HI(net963));
 sg13g2_tiehi _49029__964 (.L_HI(net964));
 sg13g2_tiehi _49028__965 (.L_HI(net965));
 sg13g2_tiehi _49027__966 (.L_HI(net966));
 sg13g2_tiehi _49026__967 (.L_HI(net967));
 sg13g2_tiehi _49025__968 (.L_HI(net968));
 sg13g2_tiehi _49024__969 (.L_HI(net969));
 sg13g2_tiehi _49023__970 (.L_HI(net970));
 sg13g2_tiehi _49022__971 (.L_HI(net971));
 sg13g2_tiehi _49021__972 (.L_HI(net972));
 sg13g2_tiehi _49020__973 (.L_HI(net973));
 sg13g2_tiehi _49019__974 (.L_HI(net974));
 sg13g2_tiehi _49018__975 (.L_HI(net975));
 sg13g2_tiehi _49017__976 (.L_HI(net976));
 sg13g2_tiehi _49016__977 (.L_HI(net977));
 sg13g2_tiehi _49015__978 (.L_HI(net978));
 sg13g2_tiehi _49014__979 (.L_HI(net979));
 sg13g2_tiehi _49013__980 (.L_HI(net980));
 sg13g2_tiehi _49012__981 (.L_HI(net981));
 sg13g2_tiehi _49011__982 (.L_HI(net982));
 sg13g2_tiehi _49010__983 (.L_HI(net983));
 sg13g2_tiehi _49009__984 (.L_HI(net984));
 sg13g2_tiehi _49008__985 (.L_HI(net985));
 sg13g2_tiehi _49007__986 (.L_HI(net986));
 sg13g2_tiehi _49006__987 (.L_HI(net987));
 sg13g2_tiehi _49005__988 (.L_HI(net988));
 sg13g2_tiehi _49004__989 (.L_HI(net989));
 sg13g2_tiehi _49003__990 (.L_HI(net990));
 sg13g2_tiehi _49002__991 (.L_HI(net991));
 sg13g2_tiehi _49001__992 (.L_HI(net992));
 sg13g2_tiehi _49000__993 (.L_HI(net993));
 sg13g2_tiehi _48999__994 (.L_HI(net994));
 sg13g2_tiehi _48998__995 (.L_HI(net995));
 sg13g2_tiehi _48997__996 (.L_HI(net996));
 sg13g2_tiehi _48996__997 (.L_HI(net997));
 sg13g2_tiehi _48995__998 (.L_HI(net998));
 sg13g2_tiehi _48994__999 (.L_HI(net999));
 sg13g2_tiehi _48993__1000 (.L_HI(net1000));
 sg13g2_tiehi _48992__1001 (.L_HI(net1001));
 sg13g2_tiehi _48991__1002 (.L_HI(net1002));
 sg13g2_tiehi _48990__1003 (.L_HI(net1003));
 sg13g2_tiehi _48989__1004 (.L_HI(net1004));
 sg13g2_tiehi _48988__1005 (.L_HI(net1005));
 sg13g2_tiehi _48987__1006 (.L_HI(net1006));
 sg13g2_tiehi _48986__1007 (.L_HI(net1007));
 sg13g2_tiehi _48985__1008 (.L_HI(net1008));
 sg13g2_tiehi _48984__1009 (.L_HI(net1009));
 sg13g2_tiehi _48983__1010 (.L_HI(net1010));
 sg13g2_tiehi _48982__1011 (.L_HI(net1011));
 sg13g2_tiehi _48981__1012 (.L_HI(net1012));
 sg13g2_tiehi _48980__1013 (.L_HI(net1013));
 sg13g2_tiehi _48979__1014 (.L_HI(net1014));
 sg13g2_tiehi _48978__1015 (.L_HI(net1015));
 sg13g2_tiehi _48977__1016 (.L_HI(net1016));
 sg13g2_tiehi _48976__1017 (.L_HI(net1017));
 sg13g2_tiehi _48975__1018 (.L_HI(net1018));
 sg13g2_tiehi _48974__1019 (.L_HI(net1019));
 sg13g2_tiehi _48973__1020 (.L_HI(net1020));
 sg13g2_tiehi _48972__1021 (.L_HI(net1021));
 sg13g2_tiehi _48971__1022 (.L_HI(net1022));
 sg13g2_tiehi _48970__1023 (.L_HI(net1023));
 sg13g2_tiehi _48969__1024 (.L_HI(net1024));
 sg13g2_tiehi _48968__1025 (.L_HI(net1025));
 sg13g2_tiehi _48967__1026 (.L_HI(net1026));
 sg13g2_tiehi _48966__1027 (.L_HI(net1027));
 sg13g2_tiehi _48965__1028 (.L_HI(net1028));
 sg13g2_tiehi _48964__1029 (.L_HI(net1029));
 sg13g2_tiehi _48963__1030 (.L_HI(net1030));
 sg13g2_tiehi _48962__1031 (.L_HI(net1031));
 sg13g2_tiehi _48961__1032 (.L_HI(net1032));
 sg13g2_tiehi _48960__1033 (.L_HI(net1033));
 sg13g2_tiehi _48959__1034 (.L_HI(net1034));
 sg13g2_tiehi _48958__1035 (.L_HI(net1035));
 sg13g2_tiehi _48957__1036 (.L_HI(net1036));
 sg13g2_tiehi _48956__1037 (.L_HI(net1037));
 sg13g2_tiehi _48955__1038 (.L_HI(net1038));
 sg13g2_tiehi _48954__1039 (.L_HI(net1039));
 sg13g2_tiehi _48953__1040 (.L_HI(net1040));
 sg13g2_tiehi _48952__1041 (.L_HI(net1041));
 sg13g2_tiehi _48951__1042 (.L_HI(net1042));
 sg13g2_tiehi _48950__1043 (.L_HI(net1043));
 sg13g2_tiehi _48949__1044 (.L_HI(net1044));
 sg13g2_tiehi _48948__1045 (.L_HI(net1045));
 sg13g2_tiehi _48947__1046 (.L_HI(net1046));
 sg13g2_tiehi _48946__1047 (.L_HI(net1047));
 sg13g2_tiehi _48945__1048 (.L_HI(net1048));
 sg13g2_tiehi _48944__1049 (.L_HI(net1049));
 sg13g2_tiehi _48943__1050 (.L_HI(net1050));
 sg13g2_tiehi _48942__1051 (.L_HI(net1051));
 sg13g2_tiehi _48941__1052 (.L_HI(net1052));
 sg13g2_tiehi _48940__1053 (.L_HI(net1053));
 sg13g2_tiehi _48939__1054 (.L_HI(net1054));
 sg13g2_tiehi _48938__1055 (.L_HI(net1055));
 sg13g2_tiehi _48937__1056 (.L_HI(net1056));
 sg13g2_tiehi _48936__1057 (.L_HI(net1057));
 sg13g2_tiehi _48935__1058 (.L_HI(net1058));
 sg13g2_tiehi tt_um_corey_1059 (.L_HI(net1059));
 sg13g2_tiehi tt_um_corey_1060 (.L_HI(net1060));
 sg13g2_tiehi tt_um_corey_1061 (.L_HI(net1061));
 sg13g2_tiehi tt_um_corey_1062 (.L_HI(net1062));
 sg13g2_tiehi tt_um_corey_1063 (.L_HI(net1063));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_corey_15 (.L_LO(net15));
 sg13g2_tielo tt_um_corey_16 (.L_LO(net16));
 sg13g2_tielo tt_um_corey_17 (.L_LO(net17));
 sg13g2_tielo tt_um_corey_18 (.L_LO(net18));
 sg13g2_tielo tt_um_corey_19 (.L_LO(net19));
 sg13g2_tielo tt_um_corey_20 (.L_LO(net20));
 sg13g2_tiehi _48934__21 (.L_HI(net21));
 sg13g2_buf_1 _51312_ (.A(accepting),
    .X(uio_out[0]));
 sg13g2_buf_8 _51313_ (.A(parity_error),
    .X(uio_out[4]));
 sg13g2_buf_1 _51314_ (.A(trng_ready),
    .X(uio_out[6]));
 sg13g2_and2_1 \u_trng.u_ro5.u_and  (.A(net1),
    .B(\u_trng.u_ro5.c[4] ),
    .X(\u_trng.u_ro5.and_out ));
 sg13g2_inv_1 \u_trng.u_ro5.u_i0  (.Y(\u_trng.u_ro5.c[0] ),
    .A(\u_trng.u_ro5.and_out ));
 sg13g2_inv_1 \u_trng.u_ro5.u_i1  (.Y(\u_trng.u_ro5.c[1] ),
    .A(\u_trng.u_ro5.c[0] ));
 sg13g2_inv_1 \u_trng.u_ro5.u_i2  (.Y(\u_trng.u_ro5.c[2] ),
    .A(\u_trng.u_ro5.c[1] ));
 sg13g2_inv_1 \u_trng.u_ro5.u_i3  (.Y(\u_trng.u_ro5.c[3] ),
    .A(\u_trng.u_ro5.c[2] ));
 sg13g2_inv_1 \u_trng.u_ro5.u_i4  (.Y(\u_trng.u_ro5.c[4] ),
    .A(\u_trng.u_ro5.c[3] ));
 sg13g2_and2_1 \u_trng.u_ro7.u_and  (.A(net1),
    .B(\u_trng.u_ro7.c[6] ),
    .X(\u_trng.u_ro7.and_out ));
 sg13g2_inv_1 \u_trng.u_ro7.u_i0  (.Y(\u_trng.u_ro7.c[0] ),
    .A(\u_trng.u_ro7.and_out ));
 sg13g2_inv_1 \u_trng.u_ro7.u_i1  (.Y(\u_trng.u_ro7.c[1] ),
    .A(\u_trng.u_ro7.c[0] ));
 sg13g2_inv_1 \u_trng.u_ro7.u_i2  (.Y(\u_trng.u_ro7.c[2] ),
    .A(\u_trng.u_ro7.c[1] ));
 sg13g2_inv_1 \u_trng.u_ro7.u_i3  (.Y(\u_trng.u_ro7.c[3] ),
    .A(\u_trng.u_ro7.c[2] ));
 sg13g2_inv_1 \u_trng.u_ro7.u_i4  (.Y(\u_trng.u_ro7.c[4] ),
    .A(\u_trng.u_ro7.c[3] ));
 sg13g2_inv_1 \u_trng.u_ro7.u_i5  (.Y(\u_trng.u_ro7.c[5] ),
    .A(\u_trng.u_ro7.c[4] ));
 sg13g2_inv_1 \u_trng.u_ro7.u_i6  (.Y(\u_trng.u_ro7.c[6] ),
    .A(\u_trng.u_ro7.c[5] ));
 sg13g2_and2_1 \u_trng.u_ro9.u_and  (.A(net1),
    .B(\u_trng.u_ro9.c[8] ),
    .X(\u_trng.u_ro9.and_out ));
 sg13g2_inv_1 \u_trng.u_ro9.u_i0  (.Y(\u_trng.u_ro9.c[0] ),
    .A(\u_trng.u_ro9.and_out ));
 sg13g2_inv_1 \u_trng.u_ro9.u_i1  (.Y(\u_trng.u_ro9.c[1] ),
    .A(\u_trng.u_ro9.c[0] ));
 sg13g2_inv_1 \u_trng.u_ro9.u_i2  (.Y(\u_trng.u_ro9.c[2] ),
    .A(\u_trng.u_ro9.c[1] ));
 sg13g2_inv_1 \u_trng.u_ro9.u_i3  (.Y(\u_trng.u_ro9.c[3] ),
    .A(\u_trng.u_ro9.c[2] ));
 sg13g2_inv_1 \u_trng.u_ro9.u_i4  (.Y(\u_trng.u_ro9.c[4] ),
    .A(\u_trng.u_ro9.c[3] ));
 sg13g2_inv_1 \u_trng.u_ro9.u_i5  (.Y(\u_trng.u_ro9.c[5] ),
    .A(\u_trng.u_ro9.c[4] ));
 sg13g2_inv_1 \u_trng.u_ro9.u_i6  (.Y(\u_trng.u_ro9.c[6] ),
    .A(\u_trng.u_ro9.c[5] ));
 sg13g2_inv_1 \u_trng.u_ro9.u_i7  (.Y(\u_trng.u_ro9.c[7] ),
    .A(\u_trng.u_ro9.c[6] ));
 sg13g2_inv_1 \u_trng.u_ro9.u_i8  (.Y(\u_trng.u_ro9.c[8] ),
    .A(\u_trng.u_ro9.c[7] ));
 sg13g2_buf_8 fanout5065 (.A(_02375_),
    .X(net5065));
 sg13g2_buf_8 fanout5066 (.A(_02375_),
    .X(net5066));
 sg13g2_buf_8 fanout5067 (.A(net5069),
    .X(net5067));
 sg13g2_buf_8 fanout5068 (.A(net5069),
    .X(net5068));
 sg13g2_buf_8 fanout5069 (.A(net5070),
    .X(net5069));
 sg13g2_buf_8 fanout5070 (.A(_02377_),
    .X(net5070));
 sg13g2_buf_8 fanout5071 (.A(net5074),
    .X(net5071));
 sg13g2_buf_8 fanout5072 (.A(net5074),
    .X(net5072));
 sg13g2_buf_8 fanout5073 (.A(net5074),
    .X(net5073));
 sg13g2_buf_8 fanout5074 (.A(_02377_),
    .X(net5074));
 sg13g2_buf_8 fanout5075 (.A(net5077),
    .X(net5075));
 sg13g2_buf_1 fanout5076 (.A(net5077),
    .X(net5076));
 sg13g2_buf_8 fanout5077 (.A(net5078),
    .X(net5077));
 sg13g2_buf_8 fanout5078 (.A(net5080),
    .X(net5078));
 sg13g2_buf_8 fanout5079 (.A(net5080),
    .X(net5079));
 sg13g2_buf_8 fanout5080 (.A(net5091),
    .X(net5080));
 sg13g2_buf_8 fanout5081 (.A(net5084),
    .X(net5081));
 sg13g2_buf_8 fanout5082 (.A(net5083),
    .X(net5082));
 sg13g2_buf_2 fanout5083 (.A(net5084),
    .X(net5083));
 sg13g2_buf_8 fanout5084 (.A(net5091),
    .X(net5084));
 sg13g2_buf_8 fanout5085 (.A(net5090),
    .X(net5085));
 sg13g2_buf_2 fanout5086 (.A(net5090),
    .X(net5086));
 sg13g2_buf_8 fanout5087 (.A(net5088),
    .X(net5087));
 sg13g2_buf_8 fanout5088 (.A(net5089),
    .X(net5088));
 sg13g2_buf_8 fanout5089 (.A(net5090),
    .X(net5089));
 sg13g2_buf_8 fanout5090 (.A(net5091),
    .X(net5090));
 sg13g2_buf_8 fanout5091 (.A(_02376_),
    .X(net5091));
 sg13g2_buf_8 fanout5092 (.A(net5093),
    .X(net5092));
 sg13g2_buf_8 fanout5093 (.A(net5094),
    .X(net5093));
 sg13g2_buf_8 fanout5094 (.A(net5100),
    .X(net5094));
 sg13g2_buf_8 fanout5095 (.A(net5100),
    .X(net5095));
 sg13g2_buf_8 fanout5096 (.A(net5100),
    .X(net5096));
 sg13g2_buf_8 fanout5097 (.A(net5099),
    .X(net5097));
 sg13g2_buf_8 fanout5098 (.A(net5099),
    .X(net5098));
 sg13g2_buf_8 fanout5099 (.A(net5100),
    .X(net5099));
 sg13g2_buf_8 fanout5100 (.A(_02374_),
    .X(net5100));
 sg13g2_buf_8 fanout5101 (.A(net5105),
    .X(net5101));
 sg13g2_buf_8 fanout5102 (.A(net5105),
    .X(net5102));
 sg13g2_buf_8 fanout5103 (.A(net5105),
    .X(net5103));
 sg13g2_buf_8 fanout5104 (.A(net5105),
    .X(net5104));
 sg13g2_buf_8 fanout5105 (.A(net5109),
    .X(net5105));
 sg13g2_buf_8 fanout5106 (.A(net5107),
    .X(net5106));
 sg13g2_buf_8 fanout5107 (.A(net5108),
    .X(net5107));
 sg13g2_buf_8 fanout5108 (.A(net5109),
    .X(net5108));
 sg13g2_buf_8 fanout5109 (.A(_02374_),
    .X(net5109));
 sg13g2_buf_8 fanout5110 (.A(net5112),
    .X(net5110));
 sg13g2_buf_8 fanout5111 (.A(net5112),
    .X(net5111));
 sg13g2_buf_8 fanout5112 (.A(net5119),
    .X(net5112));
 sg13g2_buf_8 fanout5113 (.A(net5119),
    .X(net5113));
 sg13g2_buf_1 fanout5114 (.A(net5119),
    .X(net5114));
 sg13g2_buf_8 fanout5115 (.A(net5118),
    .X(net5115));
 sg13g2_buf_2 fanout5116 (.A(net5118),
    .X(net5116));
 sg13g2_buf_8 fanout5117 (.A(net5118),
    .X(net5117));
 sg13g2_buf_8 fanout5118 (.A(net5119),
    .X(net5118));
 sg13g2_buf_8 fanout5119 (.A(_02369_),
    .X(net5119));
 sg13g2_buf_8 fanout5120 (.A(net5121),
    .X(net5120));
 sg13g2_buf_8 fanout5121 (.A(_02364_),
    .X(net5121));
 sg13g2_buf_8 fanout5122 (.A(_02364_),
    .X(net5122));
 sg13g2_buf_8 fanout5123 (.A(net5124),
    .X(net5123));
 sg13g2_buf_8 fanout5124 (.A(net5125),
    .X(net5124));
 sg13g2_buf_8 fanout5125 (.A(net5128),
    .X(net5125));
 sg13g2_buf_8 fanout5126 (.A(net5127),
    .X(net5126));
 sg13g2_buf_8 fanout5127 (.A(net5128),
    .X(net5127));
 sg13g2_buf_8 fanout5128 (.A(_02359_),
    .X(net5128));
 sg13g2_buf_8 fanout5129 (.A(net5136),
    .X(net5129));
 sg13g2_buf_2 fanout5130 (.A(net5136),
    .X(net5130));
 sg13g2_buf_8 fanout5131 (.A(net5132),
    .X(net5131));
 sg13g2_buf_8 fanout5132 (.A(net5133),
    .X(net5132));
 sg13g2_buf_2 fanout5133 (.A(net5136),
    .X(net5133));
 sg13g2_buf_8 fanout5134 (.A(net5135),
    .X(net5134));
 sg13g2_buf_8 fanout5135 (.A(net5136),
    .X(net5135));
 sg13g2_buf_8 fanout5136 (.A(_02358_),
    .X(net5136));
 sg13g2_buf_8 fanout5137 (.A(net5139),
    .X(net5137));
 sg13g2_buf_1 fanout5138 (.A(net5139),
    .X(net5138));
 sg13g2_buf_8 fanout5139 (.A(_02358_),
    .X(net5139));
 sg13g2_buf_8 fanout5140 (.A(net5141),
    .X(net5140));
 sg13g2_buf_8 fanout5141 (.A(net5143),
    .X(net5141));
 sg13g2_buf_8 fanout5142 (.A(net5143),
    .X(net5142));
 sg13g2_buf_8 fanout5143 (.A(net5150),
    .X(net5143));
 sg13g2_buf_8 fanout5144 (.A(net5145),
    .X(net5144));
 sg13g2_buf_8 fanout5145 (.A(net5146),
    .X(net5145));
 sg13g2_buf_8 fanout5146 (.A(net5150),
    .X(net5146));
 sg13g2_buf_8 fanout5147 (.A(net5148),
    .X(net5147));
 sg13g2_buf_8 fanout5148 (.A(net5149),
    .X(net5148));
 sg13g2_buf_8 fanout5149 (.A(net5150),
    .X(net5149));
 sg13g2_buf_8 fanout5150 (.A(_02358_),
    .X(net5150));
 sg13g2_buf_8 fanout5151 (.A(net5153),
    .X(net5151));
 sg13g2_buf_8 fanout5152 (.A(net5153),
    .X(net5152));
 sg13g2_buf_8 fanout5153 (.A(_02357_),
    .X(net5153));
 sg13g2_buf_8 fanout5154 (.A(net5155),
    .X(net5154));
 sg13g2_buf_8 fanout5155 (.A(net5156),
    .X(net5155));
 sg13g2_buf_8 fanout5156 (.A(net5157),
    .X(net5156));
 sg13g2_buf_8 fanout5157 (.A(net5160),
    .X(net5157));
 sg13g2_buf_8 fanout5158 (.A(net5160),
    .X(net5158));
 sg13g2_buf_8 fanout5159 (.A(net5160),
    .X(net5159));
 sg13g2_buf_8 fanout5160 (.A(_02344_),
    .X(net5160));
 sg13g2_buf_8 fanout5161 (.A(net5168),
    .X(net5161));
 sg13g2_buf_2 fanout5162 (.A(net5168),
    .X(net5162));
 sg13g2_buf_8 fanout5163 (.A(net5168),
    .X(net5163));
 sg13g2_buf_8 fanout5164 (.A(net5165),
    .X(net5164));
 sg13g2_buf_8 fanout5165 (.A(net5167),
    .X(net5165));
 sg13g2_buf_8 fanout5166 (.A(net5167),
    .X(net5166));
 sg13g2_buf_8 fanout5167 (.A(net5168),
    .X(net5167));
 sg13g2_buf_8 fanout5168 (.A(_02344_),
    .X(net5168));
 sg13g2_buf_8 fanout5169 (.A(net5170),
    .X(net5169));
 sg13g2_buf_8 fanout5170 (.A(net5172),
    .X(net5170));
 sg13g2_buf_8 fanout5171 (.A(net5172),
    .X(net5171));
 sg13g2_buf_8 fanout5172 (.A(_15902_),
    .X(net5172));
 sg13g2_buf_8 fanout5173 (.A(net5176),
    .X(net5173));
 sg13g2_buf_8 fanout5174 (.A(net5176),
    .X(net5174));
 sg13g2_buf_8 fanout5175 (.A(net5176),
    .X(net5175));
 sg13g2_buf_8 fanout5176 (.A(_15902_),
    .X(net5176));
 sg13g2_buf_8 fanout5177 (.A(net5178),
    .X(net5177));
 sg13g2_buf_8 fanout5178 (.A(net5179),
    .X(net5178));
 sg13g2_buf_16 fanout5179 (.X(net5179),
    .A(net5190));
 sg13g2_buf_8 fanout5180 (.A(net5190),
    .X(net5180));
 sg13g2_buf_1 fanout5181 (.A(net5190),
    .X(net5181));
 sg13g2_buf_8 fanout5182 (.A(net5184),
    .X(net5182));
 sg13g2_buf_1 fanout5183 (.A(net5184),
    .X(net5183));
 sg13g2_buf_8 fanout5184 (.A(net1139),
    .X(net5184));
 sg13g2_buf_8 fanout5185 (.A(net5186),
    .X(net5185));
 sg13g2_buf_8 fanout5186 (.A(net5189),
    .X(net5186));
 sg13g2_buf_8 fanout5187 (.A(net5189),
    .X(net5187));
 sg13g2_buf_8 fanout5188 (.A(net5189),
    .X(net5188));
 sg13g2_buf_8 fanout5189 (.A(net1139),
    .X(net5189));
 sg13g2_buf_8 fanout5190 (.A(_15901_),
    .X(net5190));
 sg13g2_buf_8 fanout5191 (.A(_15900_),
    .X(net5191));
 sg13g2_buf_1 fanout5192 (.A(_15900_),
    .X(net5192));
 sg13g2_buf_8 fanout5193 (.A(net5194),
    .X(net5193));
 sg13g2_buf_8 fanout5194 (.A(_15900_),
    .X(net5194));
 sg13g2_buf_8 fanout5195 (.A(net5197),
    .X(net5195));
 sg13g2_buf_8 fanout5196 (.A(net5197),
    .X(net5196));
 sg13g2_buf_8 fanout5197 (.A(net5208),
    .X(net5197));
 sg13g2_buf_8 fanout5198 (.A(net5199),
    .X(net5198));
 sg13g2_buf_2 fanout5199 (.A(net5208),
    .X(net5199));
 sg13g2_buf_8 fanout5200 (.A(net5202),
    .X(net5200));
 sg13g2_buf_8 fanout5201 (.A(net5202),
    .X(net5201));
 sg13g2_buf_8 fanout5202 (.A(net5208),
    .X(net5202));
 sg13g2_buf_8 fanout5203 (.A(net5208),
    .X(net5203));
 sg13g2_buf_8 fanout5204 (.A(net5208),
    .X(net5204));
 sg13g2_buf_8 fanout5205 (.A(net5207),
    .X(net5205));
 sg13g2_buf_8 fanout5206 (.A(net5207),
    .X(net5206));
 sg13g2_buf_8 fanout5207 (.A(net5208),
    .X(net5207));
 sg13g2_buf_8 fanout5208 (.A(_02363_),
    .X(net5208));
 sg13g2_buf_8 fanout5209 (.A(net5211),
    .X(net5209));
 sg13g2_buf_8 fanout5210 (.A(net5211),
    .X(net5210));
 sg13g2_buf_8 fanout5211 (.A(net5214),
    .X(net5211));
 sg13g2_buf_8 fanout5212 (.A(net5214),
    .X(net5212));
 sg13g2_buf_8 fanout5213 (.A(net5214),
    .X(net5213));
 sg13g2_buf_8 fanout5214 (.A(_02363_),
    .X(net5214));
 sg13g2_buf_8 fanout5215 (.A(net5217),
    .X(net5215));
 sg13g2_buf_2 fanout5216 (.A(net5217),
    .X(net5216));
 sg13g2_buf_8 fanout5217 (.A(net5220),
    .X(net5217));
 sg13g2_buf_8 fanout5218 (.A(net5219),
    .X(net5218));
 sg13g2_buf_8 fanout5219 (.A(net5220),
    .X(net5219));
 sg13g2_buf_8 fanout5220 (.A(_02363_),
    .X(net5220));
 sg13g2_buf_8 fanout5221 (.A(net5222),
    .X(net5221));
 sg13g2_buf_8 fanout5222 (.A(net5234),
    .X(net5222));
 sg13g2_buf_8 fanout5223 (.A(net5234),
    .X(net5223));
 sg13g2_buf_8 fanout5224 (.A(net5225),
    .X(net5224));
 sg13g2_buf_8 fanout5225 (.A(net5227),
    .X(net5225));
 sg13g2_buf_8 fanout5226 (.A(net5227),
    .X(net5226));
 sg13g2_buf_8 fanout5227 (.A(net5234),
    .X(net5227));
 sg13g2_buf_8 fanout5228 (.A(net5229),
    .X(net5228));
 sg13g2_buf_8 fanout5229 (.A(net5233),
    .X(net5229));
 sg13g2_buf_8 fanout5230 (.A(net5231),
    .X(net5230));
 sg13g2_buf_8 fanout5231 (.A(net5232),
    .X(net5231));
 sg13g2_buf_8 fanout5232 (.A(net5233),
    .X(net5232));
 sg13g2_buf_8 fanout5233 (.A(net5234),
    .X(net5233));
 sg13g2_buf_8 fanout5234 (.A(_02356_),
    .X(net5234));
 sg13g2_buf_8 fanout5235 (.A(net5236),
    .X(net5235));
 sg13g2_buf_8 fanout5236 (.A(net5237),
    .X(net5236));
 sg13g2_buf_8 fanout5237 (.A(_02345_),
    .X(net5237));
 sg13g2_buf_8 fanout5238 (.A(_02345_),
    .X(net5238));
 sg13g2_buf_8 fanout5239 (.A(net5240),
    .X(net5239));
 sg13g2_buf_8 fanout5240 (.A(net5241),
    .X(net5240));
 sg13g2_buf_8 fanout5241 (.A(_02343_),
    .X(net5241));
 sg13g2_buf_8 fanout5242 (.A(_02343_),
    .X(net5242));
 sg13g2_buf_8 fanout5243 (.A(_02343_),
    .X(net5243));
 sg13g2_buf_8 fanout5244 (.A(net5245),
    .X(net5244));
 sg13g2_buf_8 fanout5245 (.A(net5276),
    .X(net5245));
 sg13g2_buf_8 fanout5246 (.A(net5250),
    .X(net5246));
 sg13g2_buf_8 fanout5247 (.A(net5249),
    .X(net5247));
 sg13g2_buf_1 fanout5248 (.A(net5249),
    .X(net5248));
 sg13g2_buf_8 fanout5249 (.A(net5250),
    .X(net5249));
 sg13g2_buf_8 fanout5250 (.A(net5276),
    .X(net5250));
 sg13g2_buf_8 fanout5251 (.A(net5256),
    .X(net5251));
 sg13g2_buf_2 fanout5252 (.A(net5256),
    .X(net5252));
 sg13g2_buf_8 fanout5253 (.A(net5254),
    .X(net5253));
 sg13g2_buf_8 fanout5254 (.A(net5255),
    .X(net5254));
 sg13g2_buf_8 fanout5255 (.A(net5256),
    .X(net5255));
 sg13g2_buf_8 fanout5256 (.A(net5257),
    .X(net5256));
 sg13g2_buf_8 fanout5257 (.A(net5276),
    .X(net5257));
 sg13g2_buf_8 fanout5258 (.A(net5260),
    .X(net5258));
 sg13g2_buf_1 fanout5259 (.A(net5266),
    .X(net5259));
 sg13g2_buf_8 fanout5260 (.A(net5266),
    .X(net5260));
 sg13g2_buf_8 fanout5261 (.A(net5262),
    .X(net5261));
 sg13g2_buf_8 fanout5262 (.A(net5266),
    .X(net5262));
 sg13g2_buf_8 fanout5263 (.A(net5264),
    .X(net5263));
 sg13g2_buf_1 fanout5264 (.A(net5265),
    .X(net5264));
 sg13g2_buf_8 fanout5265 (.A(net5266),
    .X(net5265));
 sg13g2_buf_8 fanout5266 (.A(net5276),
    .X(net5266));
 sg13g2_buf_8 fanout5267 (.A(net5270),
    .X(net5267));
 sg13g2_buf_8 fanout5268 (.A(net5270),
    .X(net5268));
 sg13g2_buf_1 fanout5269 (.A(net5270),
    .X(net5269));
 sg13g2_buf_8 fanout5270 (.A(net5275),
    .X(net5270));
 sg13g2_buf_8 fanout5271 (.A(net5272),
    .X(net5271));
 sg13g2_buf_2 fanout5272 (.A(net5273),
    .X(net5272));
 sg13g2_buf_1 fanout5273 (.A(net5275),
    .X(net5273));
 sg13g2_buf_8 fanout5274 (.A(net5275),
    .X(net5274));
 sg13g2_buf_8 fanout5275 (.A(net5276),
    .X(net5275));
 sg13g2_buf_8 fanout5276 (.A(net5304),
    .X(net5276));
 sg13g2_buf_8 fanout5277 (.A(net5278),
    .X(net5277));
 sg13g2_buf_8 fanout5278 (.A(net5284),
    .X(net5278));
 sg13g2_buf_8 fanout5279 (.A(net5284),
    .X(net5279));
 sg13g2_buf_8 fanout5280 (.A(net5283),
    .X(net5280));
 sg13g2_buf_8 fanout5281 (.A(net5283),
    .X(net5281));
 sg13g2_buf_1 fanout5282 (.A(net5283),
    .X(net5282));
 sg13g2_buf_8 fanout5283 (.A(net5284),
    .X(net5283));
 sg13g2_buf_8 fanout5284 (.A(net5304),
    .X(net5284));
 sg13g2_buf_8 fanout5285 (.A(net5286),
    .X(net5285));
 sg13g2_buf_8 fanout5286 (.A(net5287),
    .X(net5286));
 sg13g2_buf_8 fanout5287 (.A(net5288),
    .X(net5287));
 sg13g2_buf_8 fanout5288 (.A(net5304),
    .X(net5288));
 sg13g2_buf_8 fanout5289 (.A(net5292),
    .X(net5289));
 sg13g2_buf_8 fanout5290 (.A(net5292),
    .X(net5290));
 sg13g2_buf_2 fanout5291 (.A(net5292),
    .X(net5291));
 sg13g2_buf_8 fanout5292 (.A(net5303),
    .X(net5292));
 sg13g2_buf_8 fanout5293 (.A(net5294),
    .X(net5293));
 sg13g2_buf_8 fanout5294 (.A(net5303),
    .X(net5294));
 sg13g2_buf_8 fanout5295 (.A(net5302),
    .X(net5295));
 sg13g2_buf_8 fanout5296 (.A(net5302),
    .X(net5296));
 sg13g2_buf_8 fanout5297 (.A(net5298),
    .X(net5297));
 sg13g2_buf_8 fanout5298 (.A(net5302),
    .X(net5298));
 sg13g2_buf_8 fanout5299 (.A(net5301),
    .X(net5299));
 sg13g2_buf_1 fanout5300 (.A(net5301),
    .X(net5300));
 sg13g2_buf_1 fanout5301 (.A(net5302),
    .X(net5301));
 sg13g2_buf_8 fanout5302 (.A(net5303),
    .X(net5302));
 sg13g2_buf_8 fanout5303 (.A(net5304),
    .X(net5303));
 sg13g2_buf_8 fanout5304 (.A(_02334_),
    .X(net5304));
 sg13g2_buf_8 fanout5305 (.A(net5306),
    .X(net5305));
 sg13g2_buf_8 fanout5306 (.A(net5308),
    .X(net5306));
 sg13g2_buf_8 fanout5307 (.A(net5308),
    .X(net5307));
 sg13g2_buf_8 fanout5308 (.A(net1065),
    .X(net5308));
 sg13g2_buf_8 fanout5309 (.A(net5310),
    .X(net5309));
 sg13g2_buf_8 fanout5310 (.A(net5311),
    .X(net5310));
 sg13g2_buf_8 fanout5311 (.A(net5312),
    .X(net5311));
 sg13g2_buf_8 fanout5312 (.A(net5314),
    .X(net5312));
 sg13g2_buf_8 fanout5313 (.A(net1140),
    .X(net5313));
 sg13g2_buf_16 fanout5314 (.X(net5314),
    .A(net1065));
 sg13g2_buf_8 fanout5315 (.A(net5318),
    .X(net5315));
 sg13g2_buf_8 fanout5316 (.A(net5318),
    .X(net5316));
 sg13g2_buf_8 fanout5317 (.A(net5318),
    .X(net5317));
 sg13g2_buf_8 fanout5318 (.A(_02333_),
    .X(net5318));
 sg13g2_buf_8 fanout5319 (.A(net5322),
    .X(net5319));
 sg13g2_buf_8 fanout5320 (.A(net5322),
    .X(net5320));
 sg13g2_buf_8 fanout5321 (.A(net5322),
    .X(net5321));
 sg13g2_buf_8 fanout5322 (.A(_02328_),
    .X(net5322));
 sg13g2_buf_8 fanout5323 (.A(net5325),
    .X(net5323));
 sg13g2_buf_1 fanout5324 (.A(net5325),
    .X(net5324));
 sg13g2_buf_8 fanout5325 (.A(net5326),
    .X(net5325));
 sg13g2_buf_8 fanout5326 (.A(net5345),
    .X(net5326));
 sg13g2_buf_8 fanout5327 (.A(net5329),
    .X(net5327));
 sg13g2_buf_8 fanout5328 (.A(net5329),
    .X(net5328));
 sg13g2_buf_8 fanout5329 (.A(net5345),
    .X(net5329));
 sg13g2_buf_8 fanout5330 (.A(net5331),
    .X(net5330));
 sg13g2_buf_8 fanout5331 (.A(net5332),
    .X(net5331));
 sg13g2_buf_8 fanout5332 (.A(net5345),
    .X(net5332));
 sg13g2_buf_8 fanout5333 (.A(net5344),
    .X(net5333));
 sg13g2_buf_8 fanout5334 (.A(net5335),
    .X(net5334));
 sg13g2_buf_2 fanout5335 (.A(net5336),
    .X(net5335));
 sg13g2_buf_8 fanout5336 (.A(net5344),
    .X(net5336));
 sg13g2_buf_8 fanout5337 (.A(net5340),
    .X(net5337));
 sg13g2_buf_8 fanout5338 (.A(net5340),
    .X(net5338));
 sg13g2_buf_2 fanout5339 (.A(net5340),
    .X(net5339));
 sg13g2_buf_8 fanout5340 (.A(net5344),
    .X(net5340));
 sg13g2_buf_8 fanout5341 (.A(net5342),
    .X(net5341));
 sg13g2_buf_1 fanout5342 (.A(net5343),
    .X(net5342));
 sg13g2_buf_8 fanout5343 (.A(net5344),
    .X(net5343));
 sg13g2_buf_8 fanout5344 (.A(net5345),
    .X(net5344));
 sg13g2_buf_8 fanout5345 (.A(_15169_),
    .X(net5345));
 sg13g2_buf_8 fanout5346 (.A(net5348),
    .X(net5346));
 sg13g2_buf_8 fanout5347 (.A(net5348),
    .X(net5347));
 sg13g2_buf_8 fanout5348 (.A(net5357),
    .X(net5348));
 sg13g2_buf_2 rebuffer78 (.A(_15152_),
    .X(net1141));
 sg13g2_buf_8 fanout5350 (.A(net5351),
    .X(net5350));
 sg13g2_buf_8 fanout5351 (.A(net5352),
    .X(net5351));
 sg13g2_buf_8 fanout5352 (.A(net5357),
    .X(net5352));
 sg13g2_buf_8 fanout5353 (.A(net5354),
    .X(net5353));
 sg13g2_buf_8 fanout5354 (.A(net5355),
    .X(net5354));
 sg13g2_buf_8 fanout5355 (.A(net5356),
    .X(net5355));
 sg13g2_buf_8 fanout5356 (.A(net1134),
    .X(net5356));
 sg13g2_buf_8 fanout5357 (.A(_15168_),
    .X(net5357));
 sg13g2_buf_8 fanout5358 (.A(net5360),
    .X(net5358));
 sg13g2_buf_1 fanout5359 (.A(net5360),
    .X(net5359));
 sg13g2_buf_8 fanout5360 (.A(net5361),
    .X(net5360));
 sg13g2_buf_8 fanout5361 (.A(net5369),
    .X(net5361));
 sg13g2_buf_8 fanout5362 (.A(net5369),
    .X(net5362));
 sg13g2_buf_8 fanout5363 (.A(net5364),
    .X(net5363));
 sg13g2_buf_8 fanout5364 (.A(net5365),
    .X(net5364));
 sg13g2_buf_8 fanout5365 (.A(net5368),
    .X(net5365));
 sg13g2_buf_8 fanout5366 (.A(net5368),
    .X(net5366));
 sg13g2_buf_8 fanout5367 (.A(net5368),
    .X(net5367));
 sg13g2_buf_8 fanout5368 (.A(net5369),
    .X(net5368));
 sg13g2_buf_8 fanout5369 (.A(net1076),
    .X(net5369));
 sg13g2_buf_8 fanout5370 (.A(net5373),
    .X(net5370));
 sg13g2_buf_8 fanout5371 (.A(net5373),
    .X(net5371));
 sg13g2_buf_1 fanout5372 (.A(net5373),
    .X(net5372));
 sg13g2_buf_8 fanout5373 (.A(net5382),
    .X(net5373));
 sg13g2_buf_8 fanout5374 (.A(net5378),
    .X(net5374));
 sg13g2_buf_8 fanout5375 (.A(net5376),
    .X(net5375));
 sg13g2_buf_8 fanout5376 (.A(net5377),
    .X(net5376));
 sg13g2_buf_8 fanout5377 (.A(net5378),
    .X(net5377));
 sg13g2_buf_8 fanout5378 (.A(net5382),
    .X(net5378));
 sg13g2_buf_8 fanout5379 (.A(net5381),
    .X(net5379));
 sg13g2_buf_1 fanout5380 (.A(net5381),
    .X(net5380));
 sg13g2_buf_8 fanout5381 (.A(net5382),
    .X(net5381));
 sg13g2_buf_8 fanout5382 (.A(net5408),
    .X(net5382));
 sg13g2_buf_8 fanout5383 (.A(net5390),
    .X(net5383));
 sg13g2_buf_8 fanout5384 (.A(net5387),
    .X(net5384));
 sg13g2_buf_8 fanout5385 (.A(net5386),
    .X(net5385));
 sg13g2_buf_8 fanout5386 (.A(net5387),
    .X(net5386));
 sg13g2_buf_8 fanout5387 (.A(net5390),
    .X(net5387));
 sg13g2_buf_8 fanout5388 (.A(net5389),
    .X(net5388));
 sg13g2_buf_8 fanout5389 (.A(net5390),
    .X(net5389));
 sg13g2_buf_8 fanout5390 (.A(net5408),
    .X(net5390));
 sg13g2_buf_8 fanout5391 (.A(net5393),
    .X(net5391));
 sg13g2_buf_8 fanout5392 (.A(net5400),
    .X(net5392));
 sg13g2_buf_2 fanout5393 (.A(net5400),
    .X(net5393));
 sg13g2_buf_8 fanout5394 (.A(net5396),
    .X(net5394));
 sg13g2_buf_1 fanout5395 (.A(net5396),
    .X(net5395));
 sg13g2_buf_8 fanout5396 (.A(net5400),
    .X(net5396));
 sg13g2_buf_8 fanout5397 (.A(net5398),
    .X(net5397));
 sg13g2_buf_1 fanout5398 (.A(net5399),
    .X(net5398));
 sg13g2_buf_2 fanout5399 (.A(net5400),
    .X(net5399));
 sg13g2_buf_8 fanout5400 (.A(net5408),
    .X(net5400));
 sg13g2_buf_8 fanout5401 (.A(net5404),
    .X(net5401));
 sg13g2_buf_8 fanout5402 (.A(net5403),
    .X(net5402));
 sg13g2_buf_2 fanout5403 (.A(net5404),
    .X(net5403));
 sg13g2_buf_8 fanout5404 (.A(net5408),
    .X(net5404));
 sg13g2_buf_8 fanout5405 (.A(net5407),
    .X(net5405));
 sg13g2_buf_1 fanout5406 (.A(net5407),
    .X(net5406));
 sg13g2_buf_8 fanout5407 (.A(net5408),
    .X(net5407));
 sg13g2_buf_8 fanout5408 (.A(_10789_),
    .X(net5408));
 sg13g2_buf_8 fanout5409 (.A(net5411),
    .X(net5409));
 sg13g2_buf_8 fanout5410 (.A(net5411),
    .X(net5410));
 sg13g2_buf_8 fanout5411 (.A(net5416),
    .X(net5411));
 sg13g2_buf_8 fanout5412 (.A(net5416),
    .X(net5412));
 sg13g2_buf_8 fanout5413 (.A(net5416),
    .X(net5413));
 sg13g2_buf_8 fanout5414 (.A(net5415),
    .X(net5414));
 sg13g2_buf_8 fanout5415 (.A(net5416),
    .X(net5415));
 sg13g2_buf_8 fanout5416 (.A(_10789_),
    .X(net5416));
 sg13g2_buf_8 fanout5417 (.A(net5420),
    .X(net5417));
 sg13g2_buf_8 fanout5418 (.A(net5419),
    .X(net5418));
 sg13g2_buf_8 fanout5419 (.A(net5420),
    .X(net5419));
 sg13g2_buf_8 fanout5420 (.A(net5431),
    .X(net5420));
 sg13g2_buf_8 fanout5421 (.A(net5431),
    .X(net5421));
 sg13g2_buf_8 fanout5422 (.A(net5424),
    .X(net5422));
 sg13g2_buf_1 fanout5423 (.A(net5424),
    .X(net5423));
 sg13g2_buf_8 fanout5424 (.A(net5431),
    .X(net5424));
 sg13g2_buf_8 fanout5425 (.A(net5429),
    .X(net5425));
 sg13g2_buf_8 fanout5426 (.A(net5429),
    .X(net5426));
 sg13g2_buf_8 fanout5427 (.A(net5429),
    .X(net5427));
 sg13g2_buf_1 fanout5428 (.A(net5429),
    .X(net5428));
 sg13g2_buf_8 fanout5429 (.A(net5430),
    .X(net5429));
 sg13g2_buf_8 fanout5430 (.A(net5431),
    .X(net5430));
 sg13g2_buf_8 fanout5431 (.A(_10789_),
    .X(net5431));
 sg13g2_buf_8 fanout5432 (.A(net5439),
    .X(net5432));
 sg13g2_buf_1 fanout5433 (.A(net5439),
    .X(net5433));
 sg13g2_buf_8 fanout5434 (.A(net5436),
    .X(net5434));
 sg13g2_buf_2 fanout5435 (.A(net5436),
    .X(net5435));
 sg13g2_buf_8 fanout5436 (.A(net5437),
    .X(net5436));
 sg13g2_buf_8 fanout5437 (.A(net5438),
    .X(net5437));
 sg13g2_buf_8 fanout5438 (.A(net5439),
    .X(net5438));
 sg13g2_buf_8 fanout5439 (.A(net5474),
    .X(net5439));
 sg13g2_buf_8 fanout5440 (.A(net5444),
    .X(net5440));
 sg13g2_buf_8 fanout5441 (.A(net5444),
    .X(net5441));
 sg13g2_buf_8 fanout5442 (.A(net5443),
    .X(net5442));
 sg13g2_buf_8 fanout5443 (.A(net5444),
    .X(net5443));
 sg13g2_buf_8 fanout5444 (.A(net5445),
    .X(net5444));
 sg13g2_buf_8 fanout5445 (.A(net5474),
    .X(net5445));
 sg13g2_buf_8 fanout5446 (.A(net5447),
    .X(net5446));
 sg13g2_buf_8 fanout5447 (.A(net5452),
    .X(net5447));
 sg13g2_buf_8 fanout5448 (.A(net5451),
    .X(net5448));
 sg13g2_buf_8 fanout5449 (.A(net5451),
    .X(net5449));
 sg13g2_buf_8 fanout5450 (.A(net5451),
    .X(net5450));
 sg13g2_buf_8 fanout5451 (.A(net5452),
    .X(net5451));
 sg13g2_buf_8 fanout5452 (.A(net5456),
    .X(net5452));
 sg13g2_buf_8 fanout5453 (.A(net5455),
    .X(net5453));
 sg13g2_buf_8 fanout5454 (.A(net5455),
    .X(net5454));
 sg13g2_buf_8 fanout5455 (.A(net5456),
    .X(net5455));
 sg13g2_buf_8 fanout5456 (.A(net5474),
    .X(net5456));
 sg13g2_buf_8 fanout5457 (.A(net5464),
    .X(net5457));
 sg13g2_buf_8 fanout5458 (.A(net5461),
    .X(net5458));
 sg13g2_buf_8 fanout5459 (.A(net5460),
    .X(net5459));
 sg13g2_buf_8 fanout5460 (.A(net5461),
    .X(net5460));
 sg13g2_buf_8 fanout5461 (.A(net5464),
    .X(net5461));
 sg13g2_buf_8 fanout5462 (.A(net5463),
    .X(net5462));
 sg13g2_buf_8 fanout5463 (.A(net5464),
    .X(net5463));
 sg13g2_buf_8 fanout5464 (.A(net5474),
    .X(net5464));
 sg13g2_buf_8 fanout5465 (.A(net5468),
    .X(net5465));
 sg13g2_buf_1 fanout5466 (.A(net5468),
    .X(net5466));
 sg13g2_buf_8 fanout5467 (.A(net5468),
    .X(net5467));
 sg13g2_buf_8 fanout5468 (.A(net5474),
    .X(net5468));
 sg13g2_buf_8 fanout5469 (.A(net5473),
    .X(net5469));
 sg13g2_buf_8 fanout5470 (.A(net5472),
    .X(net5470));
 sg13g2_buf_8 fanout5471 (.A(net5472),
    .X(net5471));
 sg13g2_buf_8 fanout5472 (.A(net5473),
    .X(net5472));
 sg13g2_buf_8 fanout5473 (.A(net5474),
    .X(net5473));
 sg13g2_buf_8 fanout5474 (.A(_10788_),
    .X(net5474));
 sg13g2_buf_8 fanout5475 (.A(_10224_),
    .X(net5475));
 sg13g2_buf_8 fanout5476 (.A(_08849_),
    .X(net5476));
 sg13g2_buf_8 fanout5477 (.A(net5480),
    .X(net5477));
 sg13g2_buf_8 fanout5478 (.A(net5479),
    .X(net5478));
 sg13g2_buf_2 fanout5479 (.A(net5480),
    .X(net5479));
 sg13g2_buf_8 fanout5480 (.A(net5496),
    .X(net5480));
 sg13g2_buf_8 fanout5481 (.A(net5482),
    .X(net5481));
 sg13g2_buf_1 fanout5482 (.A(net5488),
    .X(net5482));
 sg13g2_buf_8 fanout5483 (.A(net5488),
    .X(net5483));
 sg13g2_buf_8 fanout5484 (.A(net5488),
    .X(net5484));
 sg13g2_buf_8 fanout5485 (.A(net5486),
    .X(net5485));
 sg13g2_buf_1 fanout5486 (.A(net5488),
    .X(net5486));
 sg13g2_buf_8 fanout5487 (.A(net5488),
    .X(net5487));
 sg13g2_buf_8 fanout5488 (.A(net5496),
    .X(net5488));
 sg13g2_buf_8 fanout5489 (.A(net5490),
    .X(net5489));
 sg13g2_buf_2 fanout5490 (.A(net5492),
    .X(net5490));
 sg13g2_buf_8 fanout5491 (.A(net5492),
    .X(net5491));
 sg13g2_buf_1 fanout5492 (.A(net5496),
    .X(net5492));
 sg13g2_buf_8 fanout5493 (.A(net5496),
    .X(net5493));
 sg13g2_buf_1 fanout5494 (.A(net5495),
    .X(net5494));
 sg13g2_buf_8 fanout5495 (.A(net5496),
    .X(net5495));
 sg13g2_buf_8 fanout5496 (.A(net5547),
    .X(net5496));
 sg13g2_buf_8 fanout5497 (.A(net5499),
    .X(net5497));
 sg13g2_buf_1 fanout5498 (.A(net5499),
    .X(net5498));
 sg13g2_buf_2 fanout5499 (.A(net5510),
    .X(net5499));
 sg13g2_buf_8 fanout5500 (.A(net5501),
    .X(net5500));
 sg13g2_buf_8 fanout5501 (.A(net5510),
    .X(net5501));
 sg13g2_buf_8 fanout5502 (.A(net5504),
    .X(net5502));
 sg13g2_buf_1 fanout5503 (.A(net5504),
    .X(net5503));
 sg13g2_buf_1 fanout5504 (.A(net5505),
    .X(net5504));
 sg13g2_buf_1 fanout5505 (.A(net5510),
    .X(net5505));
 sg13g2_buf_8 fanout5506 (.A(net5508),
    .X(net5506));
 sg13g2_buf_1 fanout5507 (.A(net5508),
    .X(net5507));
 sg13g2_buf_1 fanout5508 (.A(net5509),
    .X(net5508));
 sg13g2_buf_1 fanout5509 (.A(net5510),
    .X(net5509));
 sg13g2_buf_8 fanout5510 (.A(net5547),
    .X(net5510));
 sg13g2_buf_8 fanout5511 (.A(net5515),
    .X(net5511));
 sg13g2_buf_1 fanout5512 (.A(net5515),
    .X(net5512));
 sg13g2_buf_8 fanout5513 (.A(net5515),
    .X(net5513));
 sg13g2_buf_1 fanout5514 (.A(net5515),
    .X(net5514));
 sg13g2_buf_8 fanout5515 (.A(net5519),
    .X(net5515));
 sg13g2_buf_8 fanout5516 (.A(net5519),
    .X(net5516));
 sg13g2_buf_8 fanout5517 (.A(net5518),
    .X(net5517));
 sg13g2_buf_2 fanout5518 (.A(net5519),
    .X(net5518));
 sg13g2_buf_8 fanout5519 (.A(net5547),
    .X(net5519));
 sg13g2_buf_8 fanout5520 (.A(net5522),
    .X(net5520));
 sg13g2_buf_1 fanout5521 (.A(net5522),
    .X(net5521));
 sg13g2_buf_8 fanout5522 (.A(net5527),
    .X(net5522));
 sg13g2_buf_8 fanout5523 (.A(net5527),
    .X(net5523));
 sg13g2_buf_1 fanout5524 (.A(net5527),
    .X(net5524));
 sg13g2_buf_8 fanout5525 (.A(net5526),
    .X(net5525));
 sg13g2_buf_8 fanout5526 (.A(net5527),
    .X(net5526));
 sg13g2_buf_8 fanout5527 (.A(net5547),
    .X(net5527));
 sg13g2_buf_8 fanout5528 (.A(net5530),
    .X(net5528));
 sg13g2_buf_1 fanout5529 (.A(net5530),
    .X(net5529));
 sg13g2_buf_8 fanout5530 (.A(net5531),
    .X(net5530));
 sg13g2_buf_2 fanout5531 (.A(net5547),
    .X(net5531));
 sg13g2_buf_8 fanout5532 (.A(net5546),
    .X(net5532));
 sg13g2_buf_1 fanout5533 (.A(net5546),
    .X(net5533));
 sg13g2_buf_8 fanout5534 (.A(net5535),
    .X(net5534));
 sg13g2_buf_8 fanout5535 (.A(net5536),
    .X(net5535));
 sg13g2_buf_8 fanout5536 (.A(net5546),
    .X(net5536));
 sg13g2_buf_8 fanout5537 (.A(net5546),
    .X(net5537));
 sg13g2_buf_1 fanout5538 (.A(net5546),
    .X(net5538));
 sg13g2_buf_8 fanout5539 (.A(net5540),
    .X(net5539));
 sg13g2_buf_8 fanout5540 (.A(net5545),
    .X(net5540));
 sg13g2_buf_8 fanout5541 (.A(net5544),
    .X(net5541));
 sg13g2_buf_8 fanout5542 (.A(net5543),
    .X(net5542));
 sg13g2_buf_8 fanout5543 (.A(net5544),
    .X(net5543));
 sg13g2_buf_8 fanout5544 (.A(net5545),
    .X(net5544));
 sg13g2_buf_8 fanout5545 (.A(net5546),
    .X(net5545));
 sg13g2_buf_8 fanout5546 (.A(net5547),
    .X(net5546));
 sg13g2_buf_8 fanout5547 (.A(_08583_),
    .X(net5547));
 sg13g2_buf_8 fanout5548 (.A(net5549),
    .X(net5548));
 sg13g2_buf_8 fanout5549 (.A(net5550),
    .X(net5549));
 sg13g2_buf_8 fanout5550 (.A(net5551),
    .X(net5550));
 sg13g2_buf_1 fanout5551 (.A(net5557),
    .X(net5551));
 sg13g2_buf_8 fanout5552 (.A(net5557),
    .X(net5552));
 sg13g2_buf_8 fanout5553 (.A(net5557),
    .X(net5553));
 sg13g2_buf_1 fanout5554 (.A(net5557),
    .X(net5554));
 sg13g2_buf_8 fanout5555 (.A(net5556),
    .X(net5555));
 sg13g2_buf_8 fanout5556 (.A(net5557),
    .X(net5556));
 sg13g2_buf_8 fanout5557 (.A(net5560),
    .X(net5557));
 sg13g2_buf_8 fanout5558 (.A(net5559),
    .X(net5558));
 sg13g2_buf_8 fanout5559 (.A(net5560),
    .X(net5559));
 sg13g2_buf_8 fanout5560 (.A(net5570),
    .X(net5560));
 sg13g2_buf_8 fanout5561 (.A(net5562),
    .X(net5561));
 sg13g2_buf_8 fanout5562 (.A(net5564),
    .X(net5562));
 sg13g2_buf_8 fanout5563 (.A(net5564),
    .X(net5563));
 sg13g2_buf_8 fanout5564 (.A(net5570),
    .X(net5564));
 sg13g2_buf_8 fanout5565 (.A(net5566),
    .X(net5565));
 sg13g2_buf_8 fanout5566 (.A(net5570),
    .X(net5566));
 sg13g2_buf_8 fanout5567 (.A(net5568),
    .X(net5567));
 sg13g2_buf_8 fanout5568 (.A(net5569),
    .X(net5568));
 sg13g2_buf_8 fanout5569 (.A(net5570),
    .X(net5569));
 sg13g2_buf_8 fanout5570 (.A(_08582_),
    .X(net5570));
 sg13g2_buf_8 fanout5571 (.A(net5572),
    .X(net5571));
 sg13g2_buf_8 fanout5572 (.A(net5573),
    .X(net5572));
 sg13g2_buf_8 fanout5573 (.A(net5576),
    .X(net5573));
 sg13g2_buf_8 fanout5574 (.A(net5575),
    .X(net5574));
 sg13g2_buf_1 fanout5575 (.A(net5576),
    .X(net5575));
 sg13g2_buf_8 fanout5576 (.A(net5590),
    .X(net5576));
 sg13g2_buf_8 fanout5577 (.A(net5590),
    .X(net5577));
 sg13g2_buf_8 fanout5578 (.A(net5579),
    .X(net5578));
 sg13g2_buf_2 fanout5579 (.A(net5580),
    .X(net5579));
 sg13g2_buf_8 fanout5580 (.A(net5590),
    .X(net5580));
 sg13g2_buf_8 fanout5581 (.A(net5584),
    .X(net5581));
 sg13g2_buf_8 fanout5582 (.A(net5584),
    .X(net5582));
 sg13g2_buf_1 fanout5583 (.A(net5584),
    .X(net5583));
 sg13g2_buf_8 fanout5584 (.A(net5585),
    .X(net5584));
 sg13g2_buf_8 fanout5585 (.A(net5590),
    .X(net5585));
 sg13g2_buf_8 fanout5586 (.A(net5589),
    .X(net5586));
 sg13g2_buf_8 fanout5587 (.A(net5589),
    .X(net5587));
 sg13g2_buf_1 fanout5588 (.A(net5589),
    .X(net5588));
 sg13g2_buf_8 fanout5589 (.A(net5590),
    .X(net5589));
 sg13g2_buf_8 fanout5590 (.A(_08578_),
    .X(net5590));
 sg13g2_buf_8 fanout5591 (.A(net5594),
    .X(net5591));
 sg13g2_buf_8 fanout5592 (.A(net5593),
    .X(net5592));
 sg13g2_buf_8 fanout5593 (.A(net5594),
    .X(net5593));
 sg13g2_buf_8 fanout5594 (.A(net5595),
    .X(net5594));
 sg13g2_buf_8 fanout5595 (.A(net5607),
    .X(net5595));
 sg13g2_buf_8 fanout5596 (.A(net5597),
    .X(net5596));
 sg13g2_buf_8 fanout5597 (.A(net5598),
    .X(net5597));
 sg13g2_buf_8 fanout5598 (.A(net5607),
    .X(net5598));
 sg13g2_buf_8 fanout5599 (.A(net5606),
    .X(net5599));
 sg13g2_buf_1 fanout5600 (.A(net5606),
    .X(net5600));
 sg13g2_buf_8 fanout5601 (.A(net5603),
    .X(net5601));
 sg13g2_buf_1 fanout5602 (.A(net5603),
    .X(net5602));
 sg13g2_buf_8 fanout5603 (.A(net5606),
    .X(net5603));
 sg13g2_buf_8 fanout5604 (.A(net5606),
    .X(net5604));
 sg13g2_buf_1 fanout5605 (.A(net5606),
    .X(net5605));
 sg13g2_buf_8 fanout5606 (.A(net5607),
    .X(net5606));
 sg13g2_buf_8 fanout5607 (.A(_08578_),
    .X(net5607));
 sg13g2_buf_8 fanout5608 (.A(net5610),
    .X(net5608));
 sg13g2_buf_8 fanout5609 (.A(net5610),
    .X(net5609));
 sg13g2_buf_2 fanout5610 (.A(net5613),
    .X(net5610));
 sg13g2_buf_8 fanout5611 (.A(net5613),
    .X(net5611));
 sg13g2_buf_1 fanout5612 (.A(net5613),
    .X(net5612));
 sg13g2_buf_8 fanout5613 (.A(net5621),
    .X(net5613));
 sg13g2_buf_8 fanout5614 (.A(net5615),
    .X(net5614));
 sg13g2_buf_8 fanout5615 (.A(net5616),
    .X(net5615));
 sg13g2_buf_8 fanout5616 (.A(net5617),
    .X(net5616));
 sg13g2_buf_8 fanout5617 (.A(net5621),
    .X(net5617));
 sg13g2_buf_8 fanout5618 (.A(net5619),
    .X(net5618));
 sg13g2_buf_8 fanout5619 (.A(net5620),
    .X(net5619));
 sg13g2_buf_8 fanout5620 (.A(net5621),
    .X(net5620));
 sg13g2_buf_8 fanout5621 (.A(net5651),
    .X(net5621));
 sg13g2_buf_8 fanout5622 (.A(net5630),
    .X(net5622));
 sg13g2_buf_8 fanout5623 (.A(net5625),
    .X(net5623));
 sg13g2_buf_1 fanout5624 (.A(net5625),
    .X(net5624));
 sg13g2_buf_8 fanout5625 (.A(net5626),
    .X(net5625));
 sg13g2_buf_8 fanout5626 (.A(net5630),
    .X(net5626));
 sg13g2_buf_8 fanout5627 (.A(net5628),
    .X(net5627));
 sg13g2_buf_8 fanout5628 (.A(net5629),
    .X(net5628));
 sg13g2_buf_8 fanout5629 (.A(net5630),
    .X(net5629));
 sg13g2_buf_8 fanout5630 (.A(net5651),
    .X(net5630));
 sg13g2_buf_8 fanout5631 (.A(net5632),
    .X(net5631));
 sg13g2_buf_8 fanout5632 (.A(net5643),
    .X(net5632));
 sg13g2_buf_8 fanout5633 (.A(net5635),
    .X(net5633));
 sg13g2_buf_8 fanout5634 (.A(net5635),
    .X(net5634));
 sg13g2_buf_2 fanout5635 (.A(net5643),
    .X(net5635));
 sg13g2_buf_8 fanout5636 (.A(net5638),
    .X(net5636));
 sg13g2_buf_1 fanout5637 (.A(net5638),
    .X(net5637));
 sg13g2_buf_8 fanout5638 (.A(net5639),
    .X(net5638));
 sg13g2_buf_8 fanout5639 (.A(net5643),
    .X(net5639));
 sg13g2_buf_8 fanout5640 (.A(net5642),
    .X(net5640));
 sg13g2_buf_8 fanout5641 (.A(net5642),
    .X(net5641));
 sg13g2_buf_2 fanout5642 (.A(net5643),
    .X(net5642));
 sg13g2_buf_8 fanout5643 (.A(net5651),
    .X(net5643));
 sg13g2_buf_8 fanout5644 (.A(net5647),
    .X(net5644));
 sg13g2_buf_1 fanout5645 (.A(net5647),
    .X(net5645));
 sg13g2_buf_8 fanout5646 (.A(net5647),
    .X(net5646));
 sg13g2_buf_8 fanout5647 (.A(net5651),
    .X(net5647));
 sg13g2_buf_8 fanout5648 (.A(net5650),
    .X(net5648));
 sg13g2_buf_1 fanout5649 (.A(net5650),
    .X(net5649));
 sg13g2_buf_8 fanout5650 (.A(net5651),
    .X(net5650));
 sg13g2_buf_8 fanout5651 (.A(_08577_),
    .X(net5651));
 sg13g2_buf_8 fanout5652 (.A(net5653),
    .X(net5652));
 sg13g2_buf_8 fanout5653 (.A(net5663),
    .X(net5653));
 sg13g2_buf_1 fanout5654 (.A(net5663),
    .X(net5654));
 sg13g2_buf_8 fanout5655 (.A(net5657),
    .X(net5655));
 sg13g2_buf_8 fanout5656 (.A(net5657),
    .X(net5656));
 sg13g2_buf_8 fanout5657 (.A(net5663),
    .X(net5657));
 sg13g2_buf_8 fanout5658 (.A(net5662),
    .X(net5658));
 sg13g2_buf_1 fanout5659 (.A(net5662),
    .X(net5659));
 sg13g2_buf_8 fanout5660 (.A(net5662),
    .X(net5660));
 sg13g2_buf_1 fanout5661 (.A(net5662),
    .X(net5661));
 sg13g2_buf_8 fanout5662 (.A(net5663),
    .X(net5662));
 sg13g2_buf_8 fanout5663 (.A(net5681),
    .X(net5663));
 sg13g2_buf_8 fanout5664 (.A(net5665),
    .X(net5664));
 sg13g2_buf_8 fanout5665 (.A(net5666),
    .X(net5665));
 sg13g2_buf_8 fanout5666 (.A(net5681),
    .X(net5666));
 sg13g2_buf_8 fanout5667 (.A(net5668),
    .X(net5667));
 sg13g2_buf_1 fanout5668 (.A(net5669),
    .X(net5668));
 sg13g2_buf_8 fanout5669 (.A(net5681),
    .X(net5669));
 sg13g2_buf_8 fanout5670 (.A(net5671),
    .X(net5670));
 sg13g2_buf_8 fanout5671 (.A(net5681),
    .X(net5671));
 sg13g2_buf_8 fanout5672 (.A(net5680),
    .X(net5672));
 sg13g2_buf_1 fanout5673 (.A(net5680),
    .X(net5673));
 sg13g2_buf_8 fanout5674 (.A(net5680),
    .X(net5674));
 sg13g2_buf_8 fanout5675 (.A(net5680),
    .X(net5675));
 sg13g2_buf_8 fanout5676 (.A(net5680),
    .X(net5676));
 sg13g2_buf_8 fanout5677 (.A(net5678),
    .X(net5677));
 sg13g2_buf_2 fanout5678 (.A(net5679),
    .X(net5678));
 sg13g2_buf_2 fanout5679 (.A(net5680),
    .X(net5679));
 sg13g2_buf_8 fanout5680 (.A(net5681),
    .X(net5680));
 sg13g2_buf_8 fanout5681 (.A(_08577_),
    .X(net5681));
 sg13g2_buf_8 fanout5682 (.A(net5683),
    .X(net5682));
 sg13g2_buf_8 fanout5683 (.A(net5692),
    .X(net5683));
 sg13g2_buf_8 fanout5684 (.A(net5692),
    .X(net5684));
 sg13g2_buf_8 fanout5685 (.A(net5689),
    .X(net5685));
 sg13g2_buf_8 fanout5686 (.A(net5687),
    .X(net5686));
 sg13g2_buf_8 fanout5687 (.A(net5688),
    .X(net5687));
 sg13g2_buf_8 fanout5688 (.A(net5689),
    .X(net5688));
 sg13g2_buf_8 fanout5689 (.A(net5692),
    .X(net5689));
 sg13g2_buf_8 fanout5690 (.A(net5691),
    .X(net5690));
 sg13g2_buf_1 fanout5691 (.A(net5692),
    .X(net5691));
 sg13g2_buf_8 fanout5692 (.A(net5715),
    .X(net5692));
 sg13g2_buf_8 fanout5693 (.A(net5694),
    .X(net5693));
 sg13g2_buf_2 fanout5694 (.A(net5695),
    .X(net5694));
 sg13g2_buf_1 fanout5695 (.A(net5715),
    .X(net5695));
 sg13g2_buf_8 fanout5696 (.A(net5698),
    .X(net5696));
 sg13g2_buf_8 fanout5697 (.A(net5698),
    .X(net5697));
 sg13g2_buf_8 fanout5698 (.A(net5699),
    .X(net5698));
 sg13g2_buf_8 fanout5699 (.A(net5715),
    .X(net5699));
 sg13g2_buf_8 fanout5700 (.A(net5702),
    .X(net5700));
 sg13g2_buf_8 fanout5701 (.A(net5702),
    .X(net5701));
 sg13g2_buf_8 fanout5702 (.A(net5714),
    .X(net5702));
 sg13g2_buf_8 fanout5703 (.A(net5704),
    .X(net5703));
 sg13g2_buf_8 fanout5704 (.A(net5705),
    .X(net5704));
 sg13g2_buf_8 fanout5705 (.A(net5714),
    .X(net5705));
 sg13g2_buf_8 fanout5706 (.A(net5708),
    .X(net5706));
 sg13g2_buf_1 fanout5707 (.A(net5708),
    .X(net5707));
 sg13g2_buf_2 fanout5708 (.A(net5714),
    .X(net5708));
 sg13g2_buf_8 fanout5709 (.A(net5710),
    .X(net5709));
 sg13g2_buf_8 fanout5710 (.A(net5713),
    .X(net5710));
 sg13g2_buf_8 fanout5711 (.A(net5713),
    .X(net5711));
 sg13g2_buf_1 fanout5712 (.A(net5713),
    .X(net5712));
 sg13g2_buf_8 fanout5713 (.A(net5714),
    .X(net5713));
 sg13g2_buf_8 fanout5714 (.A(net5715),
    .X(net5714));
 sg13g2_buf_8 fanout5715 (.A(_05352_),
    .X(net5715));
 sg13g2_buf_8 fanout5716 (.A(net5717),
    .X(net5716));
 sg13g2_buf_1 fanout5717 (.A(net5721),
    .X(net5717));
 sg13g2_buf_8 fanout5718 (.A(net5721),
    .X(net5718));
 sg13g2_buf_8 fanout5719 (.A(net5720),
    .X(net5719));
 sg13g2_buf_8 fanout5720 (.A(net5721),
    .X(net5720));
 sg13g2_buf_8 fanout5721 (.A(net5737),
    .X(net5721));
 sg13g2_buf_8 fanout5722 (.A(net5723),
    .X(net5722));
 sg13g2_buf_8 fanout5723 (.A(net5737),
    .X(net5723));
 sg13g2_buf_8 fanout5724 (.A(net5727),
    .X(net5724));
 sg13g2_buf_8 fanout5725 (.A(net5727),
    .X(net5725));
 sg13g2_buf_8 fanout5726 (.A(net5727),
    .X(net5726));
 sg13g2_buf_8 fanout5727 (.A(net5736),
    .X(net5727));
 sg13g2_buf_8 fanout5728 (.A(net5735),
    .X(net5728));
 sg13g2_buf_8 fanout5729 (.A(net5735),
    .X(net5729));
 sg13g2_buf_8 fanout5730 (.A(net5731),
    .X(net5730));
 sg13g2_buf_8 fanout5731 (.A(net5732),
    .X(net5731));
 sg13g2_buf_8 fanout5732 (.A(net5735),
    .X(net5732));
 sg13g2_buf_8 fanout5733 (.A(net5734),
    .X(net5733));
 sg13g2_buf_8 fanout5734 (.A(net5735),
    .X(net5734));
 sg13g2_buf_8 fanout5735 (.A(net5736),
    .X(net5735));
 sg13g2_buf_8 fanout5736 (.A(net5737),
    .X(net5736));
 sg13g2_buf_8 fanout5737 (.A(_05352_),
    .X(net5737));
 sg13g2_buf_8 fanout5738 (.A(net5740),
    .X(net5738));
 sg13g2_buf_1 fanout5739 (.A(net5740),
    .X(net5739));
 sg13g2_buf_2 fanout5740 (.A(net5743),
    .X(net5740));
 sg13g2_buf_8 fanout5741 (.A(net5742),
    .X(net5741));
 sg13g2_buf_2 fanout5742 (.A(net5743),
    .X(net5742));
 sg13g2_buf_8 fanout5743 (.A(net5749),
    .X(net5743));
 sg13g2_buf_8 fanout5744 (.A(net5745),
    .X(net5744));
 sg13g2_buf_8 fanout5745 (.A(net5749),
    .X(net5745));
 sg13g2_buf_8 fanout5746 (.A(net5747),
    .X(net5746));
 sg13g2_buf_1 fanout5747 (.A(net5749),
    .X(net5747));
 sg13g2_buf_8 fanout5748 (.A(net5749),
    .X(net5748));
 sg13g2_buf_8 fanout5749 (.A(net5773),
    .X(net5749));
 sg13g2_buf_8 fanout5750 (.A(net5753),
    .X(net5750));
 sg13g2_buf_8 fanout5751 (.A(net5753),
    .X(net5751));
 sg13g2_buf_8 fanout5752 (.A(net5753),
    .X(net5752));
 sg13g2_buf_8 fanout5753 (.A(net5773),
    .X(net5753));
 sg13g2_buf_8 fanout5754 (.A(net5757),
    .X(net5754));
 sg13g2_buf_8 fanout5755 (.A(net5757),
    .X(net5755));
 sg13g2_buf_1 fanout5756 (.A(net5757),
    .X(net5756));
 sg13g2_buf_8 fanout5757 (.A(net5773),
    .X(net5757));
 sg13g2_buf_8 fanout5758 (.A(net5759),
    .X(net5758));
 sg13g2_buf_8 fanout5759 (.A(net5762),
    .X(net5759));
 sg13g2_buf_8 fanout5760 (.A(net5761),
    .X(net5760));
 sg13g2_buf_8 fanout5761 (.A(net5762),
    .X(net5761));
 sg13g2_buf_8 fanout5762 (.A(net5772),
    .X(net5762));
 sg13g2_buf_8 fanout5763 (.A(net5764),
    .X(net5763));
 sg13g2_buf_8 fanout5764 (.A(net5772),
    .X(net5764));
 sg13g2_buf_8 fanout5765 (.A(net5766),
    .X(net5765));
 sg13g2_buf_8 fanout5766 (.A(net5767),
    .X(net5766));
 sg13g2_buf_8 fanout5767 (.A(net5772),
    .X(net5767));
 sg13g2_buf_8 fanout5768 (.A(net5770),
    .X(net5768));
 sg13g2_buf_8 fanout5769 (.A(net5770),
    .X(net5769));
 sg13g2_buf_8 fanout5770 (.A(net5771),
    .X(net5770));
 sg13g2_buf_8 fanout5771 (.A(net5772),
    .X(net5771));
 sg13g2_buf_8 fanout5772 (.A(net5773),
    .X(net5772));
 sg13g2_buf_8 fanout5773 (.A(_05351_),
    .X(net5773));
 sg13g2_buf_8 fanout5774 (.A(net5776),
    .X(net5774));
 sg13g2_buf_8 fanout5775 (.A(net5776),
    .X(net5775));
 sg13g2_buf_2 fanout5776 (.A(net5786),
    .X(net5776));
 sg13g2_buf_8 fanout5777 (.A(net5782),
    .X(net5777));
 sg13g2_buf_8 fanout5778 (.A(net5781),
    .X(net5778));
 sg13g2_buf_8 fanout5779 (.A(net5781),
    .X(net5779));
 sg13g2_buf_1 fanout5780 (.A(net5781),
    .X(net5780));
 sg13g2_buf_8 fanout5781 (.A(net5782),
    .X(net5781));
 sg13g2_buf_8 fanout5782 (.A(net5786),
    .X(net5782));
 sg13g2_buf_8 fanout5783 (.A(net5785),
    .X(net5783));
 sg13g2_buf_1 fanout5784 (.A(net5785),
    .X(net5784));
 sg13g2_buf_8 fanout5785 (.A(net5786),
    .X(net5785));
 sg13g2_buf_8 fanout5786 (.A(net5835),
    .X(net5786));
 sg13g2_buf_8 fanout5787 (.A(net5788),
    .X(net5787));
 sg13g2_buf_8 fanout5788 (.A(net5790),
    .X(net5788));
 sg13g2_buf_8 fanout5789 (.A(net5790),
    .X(net5789));
 sg13g2_buf_8 fanout5790 (.A(net5793),
    .X(net5790));
 sg13g2_buf_8 fanout5791 (.A(net5792),
    .X(net5791));
 sg13g2_buf_8 fanout5792 (.A(net5793),
    .X(net5792));
 sg13g2_buf_8 fanout5793 (.A(net5835),
    .X(net5793));
 sg13g2_buf_8 fanout5794 (.A(net5795),
    .X(net5794));
 sg13g2_buf_8 fanout5795 (.A(net5808),
    .X(net5795));
 sg13g2_buf_8 fanout5796 (.A(net5797),
    .X(net5796));
 sg13g2_buf_8 fanout5797 (.A(net5798),
    .X(net5797));
 sg13g2_buf_8 fanout5798 (.A(net5808),
    .X(net5798));
 sg13g2_buf_8 fanout5799 (.A(net5801),
    .X(net5799));
 sg13g2_buf_8 fanout5800 (.A(net5801),
    .X(net5800));
 sg13g2_buf_8 fanout5801 (.A(net5808),
    .X(net5801));
 sg13g2_buf_8 fanout5802 (.A(net5803),
    .X(net5802));
 sg13g2_buf_8 fanout5803 (.A(net5808),
    .X(net5803));
 sg13g2_buf_8 fanout5804 (.A(net5807),
    .X(net5804));
 sg13g2_buf_8 fanout5805 (.A(net5806),
    .X(net5805));
 sg13g2_buf_2 fanout5806 (.A(net5807),
    .X(net5806));
 sg13g2_buf_1 fanout5807 (.A(net5808),
    .X(net5807));
 sg13g2_buf_8 fanout5808 (.A(net5835),
    .X(net5808));
 sg13g2_buf_8 fanout5809 (.A(net5812),
    .X(net5809));
 sg13g2_buf_8 fanout5810 (.A(net5812),
    .X(net5810));
 sg13g2_buf_1 fanout5811 (.A(net5812),
    .X(net5811));
 sg13g2_buf_8 fanout5812 (.A(net5820),
    .X(net5812));
 sg13g2_buf_8 fanout5813 (.A(net5814),
    .X(net5813));
 sg13g2_buf_8 fanout5814 (.A(net5820),
    .X(net5814));
 sg13g2_buf_8 fanout5815 (.A(net5817),
    .X(net5815));
 sg13g2_buf_1 fanout5816 (.A(net5817),
    .X(net5816));
 sg13g2_buf_1 fanout5817 (.A(net5820),
    .X(net5817));
 sg13g2_buf_8 fanout5818 (.A(net5819),
    .X(net5818));
 sg13g2_buf_8 fanout5819 (.A(net5820),
    .X(net5819));
 sg13g2_buf_8 fanout5820 (.A(net5834),
    .X(net5820));
 sg13g2_buf_8 fanout5821 (.A(net5822),
    .X(net5821));
 sg13g2_buf_1 fanout5822 (.A(net5834),
    .X(net5822));
 sg13g2_buf_8 fanout5823 (.A(net5825),
    .X(net5823));
 sg13g2_buf_8 fanout5824 (.A(net5825),
    .X(net5824));
 sg13g2_buf_8 fanout5825 (.A(net5826),
    .X(net5825));
 sg13g2_buf_8 fanout5826 (.A(net5834),
    .X(net5826));
 sg13g2_buf_8 fanout5827 (.A(net5828),
    .X(net5827));
 sg13g2_buf_8 fanout5828 (.A(net5829),
    .X(net5828));
 sg13g2_buf_2 fanout5829 (.A(net5833),
    .X(net5829));
 sg13g2_buf_8 fanout5830 (.A(net5831),
    .X(net5830));
 sg13g2_buf_8 fanout5831 (.A(net5832),
    .X(net5831));
 sg13g2_buf_8 fanout5832 (.A(net5833),
    .X(net5832));
 sg13g2_buf_8 fanout5833 (.A(net5834),
    .X(net5833));
 sg13g2_buf_8 fanout5834 (.A(net5835),
    .X(net5834));
 sg13g2_buf_8 fanout5835 (.A(_05343_),
    .X(net5835));
 sg13g2_buf_8 fanout5836 (.A(net5839),
    .X(net5836));
 sg13g2_buf_8 fanout5837 (.A(net5838),
    .X(net5837));
 sg13g2_buf_8 fanout5838 (.A(net5839),
    .X(net5838));
 sg13g2_buf_8 fanout5839 (.A(net5857),
    .X(net5839));
 sg13g2_buf_8 fanout5840 (.A(net5844),
    .X(net5840));
 sg13g2_buf_2 fanout5841 (.A(net5844),
    .X(net5841));
 sg13g2_buf_8 fanout5842 (.A(net5843),
    .X(net5842));
 sg13g2_buf_8 fanout5843 (.A(net5844),
    .X(net5843));
 sg13g2_buf_8 fanout5844 (.A(net5845),
    .X(net5844));
 sg13g2_buf_8 fanout5845 (.A(net5857),
    .X(net5845));
 sg13g2_buf_8 fanout5846 (.A(net5847),
    .X(net5846));
 sg13g2_buf_1 fanout5847 (.A(net5852),
    .X(net5847));
 sg13g2_buf_8 fanout5848 (.A(net5852),
    .X(net5848));
 sg13g2_buf_8 fanout5849 (.A(net5850),
    .X(net5849));
 sg13g2_buf_8 fanout5850 (.A(net5851),
    .X(net5850));
 sg13g2_buf_8 fanout5851 (.A(net5852),
    .X(net5851));
 sg13g2_buf_8 fanout5852 (.A(net5857),
    .X(net5852));
 sg13g2_buf_8 fanout5853 (.A(net5854),
    .X(net5853));
 sg13g2_buf_8 fanout5854 (.A(net5857),
    .X(net5854));
 sg13g2_buf_8 fanout5855 (.A(net5856),
    .X(net5855));
 sg13g2_buf_8 fanout5856 (.A(net5857),
    .X(net5856));
 sg13g2_buf_8 fanout5857 (.A(net5879),
    .X(net5857));
 sg13g2_buf_8 fanout5858 (.A(net5861),
    .X(net5858));
 sg13g2_buf_2 fanout5859 (.A(net5861),
    .X(net5859));
 sg13g2_buf_8 fanout5860 (.A(net5861),
    .X(net5860));
 sg13g2_buf_8 fanout5861 (.A(net5864),
    .X(net5861));
 sg13g2_buf_8 fanout5862 (.A(net5864),
    .X(net5862));
 sg13g2_buf_8 fanout5863 (.A(net5864),
    .X(net5863));
 sg13g2_buf_8 fanout5864 (.A(net5879),
    .X(net5864));
 sg13g2_buf_8 fanout5865 (.A(net5866),
    .X(net5865));
 sg13g2_buf_8 fanout5866 (.A(net5879),
    .X(net5866));
 sg13g2_buf_8 fanout5867 (.A(net5871),
    .X(net5867));
 sg13g2_buf_8 fanout5868 (.A(net5870),
    .X(net5868));
 sg13g2_buf_1 fanout5869 (.A(net5870),
    .X(net5869));
 sg13g2_buf_8 fanout5870 (.A(net5871),
    .X(net5870));
 sg13g2_buf_8 fanout5871 (.A(net5878),
    .X(net5871));
 sg13g2_buf_8 fanout5872 (.A(net5878),
    .X(net5872));
 sg13g2_buf_8 fanout5873 (.A(net5878),
    .X(net5873));
 sg13g2_buf_8 fanout5874 (.A(net5877),
    .X(net5874));
 sg13g2_buf_8 fanout5875 (.A(net5877),
    .X(net5875));
 sg13g2_buf_8 fanout5876 (.A(net5877),
    .X(net5876));
 sg13g2_buf_8 fanout5877 (.A(net5878),
    .X(net5877));
 sg13g2_buf_8 fanout5878 (.A(net5879),
    .X(net5878));
 sg13g2_buf_8 fanout5879 (.A(_05342_),
    .X(net5879));
 sg13g2_buf_8 fanout5880 (.A(net5883),
    .X(net5880));
 sg13g2_buf_8 fanout5881 (.A(net5882),
    .X(net5881));
 sg13g2_buf_8 fanout5882 (.A(net5883),
    .X(net5882));
 sg13g2_buf_8 fanout5883 (.A(_02362_),
    .X(net5883));
 sg13g2_buf_8 fanout5884 (.A(net5885),
    .X(net5884));
 sg13g2_buf_8 fanout5885 (.A(net5917),
    .X(net5885));
 sg13g2_buf_8 fanout5886 (.A(net5891),
    .X(net5886));
 sg13g2_buf_8 fanout5887 (.A(net5888),
    .X(net5887));
 sg13g2_buf_8 fanout5888 (.A(net5890),
    .X(net5888));
 sg13g2_buf_8 fanout5889 (.A(net5890),
    .X(net5889));
 sg13g2_buf_8 fanout5890 (.A(net5891),
    .X(net5890));
 sg13g2_buf_8 fanout5891 (.A(net5917),
    .X(net5891));
 sg13g2_buf_8 fanout5892 (.A(net5896),
    .X(net5892));
 sg13g2_buf_8 fanout5893 (.A(net5895),
    .X(net5893));
 sg13g2_buf_8 fanout5894 (.A(net5895),
    .X(net5894));
 sg13g2_buf_8 fanout5895 (.A(net5896),
    .X(net5895));
 sg13g2_buf_8 fanout5896 (.A(net5901),
    .X(net5896));
 sg13g2_buf_8 fanout5897 (.A(net5901),
    .X(net5897));
 sg13g2_buf_8 fanout5898 (.A(net5901),
    .X(net5898));
 sg13g2_buf_8 fanout5899 (.A(net5900),
    .X(net5899));
 sg13g2_buf_8 fanout5900 (.A(net5901),
    .X(net5900));
 sg13g2_buf_8 fanout5901 (.A(net5917),
    .X(net5901));
 sg13g2_buf_8 fanout5902 (.A(net5907),
    .X(net5902));
 sg13g2_buf_8 fanout5903 (.A(net5904),
    .X(net5903));
 sg13g2_buf_8 fanout5904 (.A(net5907),
    .X(net5904));
 sg13g2_buf_8 fanout5905 (.A(net5906),
    .X(net5905));
 sg13g2_buf_8 fanout5906 (.A(net5907),
    .X(net5906));
 sg13g2_buf_8 fanout5907 (.A(net5916),
    .X(net5907));
 sg13g2_buf_8 fanout5908 (.A(net5916),
    .X(net5908));
 sg13g2_buf_8 fanout5909 (.A(net5916),
    .X(net5909));
 sg13g2_buf_8 fanout5910 (.A(net5915),
    .X(net5910));
 sg13g2_buf_8 fanout5911 (.A(net5915),
    .X(net5911));
 sg13g2_buf_8 fanout5912 (.A(net5914),
    .X(net5912));
 sg13g2_buf_8 fanout5913 (.A(net5914),
    .X(net5913));
 sg13g2_buf_8 fanout5914 (.A(net5915),
    .X(net5914));
 sg13g2_buf_8 fanout5915 (.A(net5916),
    .X(net5915));
 sg13g2_buf_8 fanout5916 (.A(net5917),
    .X(net5916));
 sg13g2_buf_8 fanout5917 (.A(_02361_),
    .X(net5917));
 sg13g2_buf_8 fanout5918 (.A(net5919),
    .X(net5918));
 sg13g2_buf_8 fanout5919 (.A(net5925),
    .X(net5919));
 sg13g2_buf_8 fanout5920 (.A(net5925),
    .X(net5920));
 sg13g2_buf_1 fanout5921 (.A(net5925),
    .X(net5921));
 sg13g2_buf_8 fanout5922 (.A(net5923),
    .X(net5922));
 sg13g2_buf_8 fanout5923 (.A(net5924),
    .X(net5923));
 sg13g2_buf_8 fanout5924 (.A(net5925),
    .X(net5924));
 sg13g2_buf_8 fanout5925 (.A(_02355_),
    .X(net5925));
 sg13g2_buf_8 fanout5926 (.A(net5929),
    .X(net5926));
 sg13g2_buf_8 fanout5927 (.A(net5928),
    .X(net5927));
 sg13g2_buf_8 fanout5928 (.A(net5929),
    .X(net5928));
 sg13g2_buf_8 fanout5929 (.A(net5934),
    .X(net5929));
 sg13g2_buf_8 fanout5930 (.A(net5934),
    .X(net5930));
 sg13g2_buf_8 fanout5931 (.A(net5934),
    .X(net5931));
 sg13g2_buf_8 fanout5932 (.A(net5933),
    .X(net5932));
 sg13g2_buf_8 fanout5933 (.A(net5934),
    .X(net5933));
 sg13g2_buf_8 fanout5934 (.A(_02355_),
    .X(net5934));
 sg13g2_buf_8 fanout5935 (.A(net5937),
    .X(net5935));
 sg13g2_buf_1 fanout5936 (.A(net5937),
    .X(net5936));
 sg13g2_buf_8 fanout5937 (.A(net5938),
    .X(net5937));
 sg13g2_buf_8 fanout5938 (.A(net5942),
    .X(net5938));
 sg13g2_buf_8 fanout5939 (.A(net5942),
    .X(net5939));
 sg13g2_buf_8 fanout5940 (.A(net5942),
    .X(net5940));
 sg13g2_buf_8 fanout5941 (.A(net5942),
    .X(net5941));
 sg13g2_buf_8 fanout5942 (.A(net5969),
    .X(net5942));
 sg13g2_buf_8 fanout5943 (.A(net5946),
    .X(net5943));
 sg13g2_buf_8 fanout5944 (.A(net5946),
    .X(net5944));
 sg13g2_buf_2 fanout5945 (.A(net5946),
    .X(net5945));
 sg13g2_buf_8 fanout5946 (.A(net5969),
    .X(net5946));
 sg13g2_buf_8 fanout5947 (.A(net5951),
    .X(net5947));
 sg13g2_buf_8 fanout5948 (.A(net5951),
    .X(net5948));
 sg13g2_buf_8 fanout5949 (.A(net5950),
    .X(net5949));
 sg13g2_buf_8 fanout5950 (.A(net5951),
    .X(net5950));
 sg13g2_buf_8 fanout5951 (.A(net5969),
    .X(net5951));
 sg13g2_buf_8 fanout5952 (.A(net5955),
    .X(net5952));
 sg13g2_buf_8 fanout5953 (.A(net5955),
    .X(net5953));
 sg13g2_buf_1 fanout5954 (.A(net5955),
    .X(net5954));
 sg13g2_buf_8 fanout5955 (.A(net5959),
    .X(net5955));
 sg13g2_buf_8 fanout5956 (.A(net5959),
    .X(net5956));
 sg13g2_buf_2 fanout5957 (.A(net5959),
    .X(net5957));
 sg13g2_buf_8 fanout5958 (.A(net5959),
    .X(net5958));
 sg13g2_buf_8 fanout5959 (.A(net5969),
    .X(net5959));
 sg13g2_buf_8 fanout5960 (.A(net5961),
    .X(net5960));
 sg13g2_buf_8 fanout5961 (.A(net5968),
    .X(net5961));
 sg13g2_buf_8 fanout5962 (.A(net5963),
    .X(net5962));
 sg13g2_buf_8 fanout5963 (.A(net5968),
    .X(net5963));
 sg13g2_buf_8 fanout5964 (.A(net5967),
    .X(net5964));
 sg13g2_buf_8 fanout5965 (.A(net5966),
    .X(net5965));
 sg13g2_buf_8 fanout5966 (.A(net5967),
    .X(net5966));
 sg13g2_buf_8 fanout5967 (.A(net5968),
    .X(net5967));
 sg13g2_buf_8 fanout5968 (.A(net5969),
    .X(net5968));
 sg13g2_buf_8 fanout5969 (.A(_02354_),
    .X(net5969));
 sg13g2_buf_8 fanout5970 (.A(net5985),
    .X(net5970));
 sg13g2_buf_1 fanout5971 (.A(net5985),
    .X(net5971));
 sg13g2_buf_8 fanout5972 (.A(net5973),
    .X(net5972));
 sg13g2_buf_8 fanout5973 (.A(net5975),
    .X(net5973));
 sg13g2_buf_8 fanout5974 (.A(net5975),
    .X(net5974));
 sg13g2_buf_8 fanout5975 (.A(net5976),
    .X(net5975));
 sg13g2_buf_8 fanout5976 (.A(net5985),
    .X(net5976));
 sg13g2_buf_8 fanout5977 (.A(net5980),
    .X(net5977));
 sg13g2_buf_8 fanout5978 (.A(net5979),
    .X(net5978));
 sg13g2_buf_8 fanout5979 (.A(net5980),
    .X(net5979));
 sg13g2_buf_8 fanout5980 (.A(net5985),
    .X(net5980));
 sg13g2_buf_8 fanout5981 (.A(net5982),
    .X(net5981));
 sg13g2_buf_8 fanout5982 (.A(net5985),
    .X(net5982));
 sg13g2_buf_8 fanout5983 (.A(net5984),
    .X(net5983));
 sg13g2_buf_8 fanout5984 (.A(net5985),
    .X(net5984));
 sg13g2_buf_8 fanout5985 (.A(_02342_),
    .X(net5985));
 sg13g2_buf_8 fanout5986 (.A(net5988),
    .X(net5986));
 sg13g2_buf_8 fanout5987 (.A(net5988),
    .X(net5987));
 sg13g2_buf_8 fanout5988 (.A(net6002),
    .X(net5988));
 sg13g2_buf_8 fanout5989 (.A(net6002),
    .X(net5989));
 sg13g2_buf_8 fanout5990 (.A(net5991),
    .X(net5990));
 sg13g2_buf_8 fanout5991 (.A(net5992),
    .X(net5991));
 sg13g2_buf_8 fanout5992 (.A(net6002),
    .X(net5992));
 sg13g2_buf_8 fanout5993 (.A(net6002),
    .X(net5993));
 sg13g2_buf_8 fanout5994 (.A(net6002),
    .X(net5994));
 sg13g2_buf_8 fanout5995 (.A(net6000),
    .X(net5995));
 sg13g2_buf_8 fanout5996 (.A(net6000),
    .X(net5996));
 sg13g2_buf_8 fanout5997 (.A(net5998),
    .X(net5997));
 sg13g2_buf_8 fanout5998 (.A(net6000),
    .X(net5998));
 sg13g2_buf_1 fanout5999 (.A(net6000),
    .X(net5999));
 sg13g2_buf_8 fanout6000 (.A(net6001),
    .X(net6000));
 sg13g2_buf_8 fanout6001 (.A(net6002),
    .X(net6001));
 sg13g2_buf_8 fanout6002 (.A(_02342_),
    .X(net6002));
 sg13g2_buf_8 fanout6003 (.A(net6005),
    .X(net6003));
 sg13g2_buf_8 fanout6004 (.A(net6005),
    .X(net6004));
 sg13g2_buf_8 fanout6005 (.A(_02341_),
    .X(net6005));
 sg13g2_buf_8 fanout6006 (.A(_02341_),
    .X(net6006));
 sg13g2_buf_8 fanout6007 (.A(net6008),
    .X(net6007));
 sg13g2_buf_8 fanout6008 (.A(_02341_),
    .X(net6008));
 sg13g2_buf_8 fanout6009 (.A(net6013),
    .X(net6009));
 sg13g2_buf_1 fanout6010 (.A(net6013),
    .X(net6010));
 sg13g2_buf_8 fanout6011 (.A(net6013),
    .X(net6011));
 sg13g2_buf_1 fanout6012 (.A(net6013),
    .X(net6012));
 sg13g2_buf_8 fanout6013 (.A(net6032),
    .X(net6013));
 sg13g2_buf_8 fanout6014 (.A(net6019),
    .X(net6014));
 sg13g2_buf_1 fanout6015 (.A(net6019),
    .X(net6015));
 sg13g2_buf_8 fanout6016 (.A(net6018),
    .X(net6016));
 sg13g2_buf_1 fanout6017 (.A(net6018),
    .X(net6017));
 sg13g2_buf_8 fanout6018 (.A(net6019),
    .X(net6018));
 sg13g2_buf_8 fanout6019 (.A(net6032),
    .X(net6019));
 sg13g2_buf_8 fanout6020 (.A(net6022),
    .X(net6020));
 sg13g2_buf_8 fanout6021 (.A(net6022),
    .X(net6021));
 sg13g2_buf_8 fanout6022 (.A(net6032),
    .X(net6022));
 sg13g2_buf_8 fanout6023 (.A(net6024),
    .X(net6023));
 sg13g2_buf_2 fanout6024 (.A(net6026),
    .X(net6024));
 sg13g2_buf_8 fanout6025 (.A(net6026),
    .X(net6025));
 sg13g2_buf_1 fanout6026 (.A(net6031),
    .X(net6026));
 sg13g2_buf_8 fanout6027 (.A(net6028),
    .X(net6027));
 sg13g2_buf_8 fanout6028 (.A(net6029),
    .X(net6028));
 sg13g2_buf_8 fanout6029 (.A(net6031),
    .X(net6029));
 sg13g2_buf_8 fanout6030 (.A(net6031),
    .X(net6030));
 sg13g2_buf_8 fanout6031 (.A(net6032),
    .X(net6031));
 sg13g2_buf_8 fanout6032 (.A(net6191),
    .X(net6032));
 sg13g2_buf_8 fanout6033 (.A(net6034),
    .X(net6033));
 sg13g2_buf_8 fanout6034 (.A(net6035),
    .X(net6034));
 sg13g2_buf_8 fanout6035 (.A(net6037),
    .X(net6035));
 sg13g2_buf_8 fanout6036 (.A(net6037),
    .X(net6036));
 sg13g2_buf_8 fanout6037 (.A(net6054),
    .X(net6037));
 sg13g2_buf_8 fanout6038 (.A(net6039),
    .X(net6038));
 sg13g2_buf_2 fanout6039 (.A(net6042),
    .X(net6039));
 sg13g2_buf_8 fanout6040 (.A(net6042),
    .X(net6040));
 sg13g2_buf_1 fanout6041 (.A(net6042),
    .X(net6041));
 sg13g2_buf_8 fanout6042 (.A(net6054),
    .X(net6042));
 sg13g2_buf_8 fanout6043 (.A(net6047),
    .X(net6043));
 sg13g2_buf_1 fanout6044 (.A(net6047),
    .X(net6044));
 sg13g2_buf_8 fanout6045 (.A(net6047),
    .X(net6045));
 sg13g2_buf_8 fanout6046 (.A(net6047),
    .X(net6046));
 sg13g2_buf_8 fanout6047 (.A(net6054),
    .X(net6047));
 sg13g2_buf_8 fanout6048 (.A(net6050),
    .X(net6048));
 sg13g2_buf_8 fanout6049 (.A(net6050),
    .X(net6049));
 sg13g2_buf_8 fanout6050 (.A(net6054),
    .X(net6050));
 sg13g2_buf_8 fanout6051 (.A(net6052),
    .X(net6051));
 sg13g2_buf_2 fanout6052 (.A(net6053),
    .X(net6052));
 sg13g2_buf_2 fanout6053 (.A(net6054),
    .X(net6053));
 sg13g2_buf_8 fanout6054 (.A(net6191),
    .X(net6054));
 sg13g2_buf_8 fanout6055 (.A(net6056),
    .X(net6055));
 sg13g2_buf_8 fanout6056 (.A(net6059),
    .X(net6056));
 sg13g2_buf_8 fanout6057 (.A(net6058),
    .X(net6057));
 sg13g2_buf_8 fanout6058 (.A(net6059),
    .X(net6058));
 sg13g2_buf_8 fanout6059 (.A(net6076),
    .X(net6059));
 sg13g2_buf_8 fanout6060 (.A(net6061),
    .X(net6060));
 sg13g2_buf_8 fanout6061 (.A(net6064),
    .X(net6061));
 sg13g2_buf_8 fanout6062 (.A(net6064),
    .X(net6062));
 sg13g2_buf_8 fanout6063 (.A(net6064),
    .X(net6063));
 sg13g2_buf_8 fanout6064 (.A(net6076),
    .X(net6064));
 sg13g2_buf_8 fanout6065 (.A(net6066),
    .X(net6065));
 sg13g2_buf_8 fanout6066 (.A(net6067),
    .X(net6066));
 sg13g2_buf_2 fanout6067 (.A(net6070),
    .X(net6067));
 sg13g2_buf_8 fanout6068 (.A(net6069),
    .X(net6068));
 sg13g2_buf_8 fanout6069 (.A(net6070),
    .X(net6069));
 sg13g2_buf_8 fanout6070 (.A(net6076),
    .X(net6070));
 sg13g2_buf_8 fanout6071 (.A(net6075),
    .X(net6071));
 sg13g2_buf_1 fanout6072 (.A(net6075),
    .X(net6072));
 sg13g2_buf_8 fanout6073 (.A(net6075),
    .X(net6073));
 sg13g2_buf_2 fanout6074 (.A(net6075),
    .X(net6074));
 sg13g2_buf_8 fanout6075 (.A(net6076),
    .X(net6075));
 sg13g2_buf_8 fanout6076 (.A(net6096),
    .X(net6076));
 sg13g2_buf_8 fanout6077 (.A(net6080),
    .X(net6077));
 sg13g2_buf_8 fanout6078 (.A(net6080),
    .X(net6078));
 sg13g2_buf_2 fanout6079 (.A(net6080),
    .X(net6079));
 sg13g2_buf_8 fanout6080 (.A(net6081),
    .X(net6080));
 sg13g2_buf_8 fanout6081 (.A(net6086),
    .X(net6081));
 sg13g2_buf_8 fanout6082 (.A(net6083),
    .X(net6082));
 sg13g2_buf_8 fanout6083 (.A(net6086),
    .X(net6083));
 sg13g2_buf_8 fanout6084 (.A(net6085),
    .X(net6084));
 sg13g2_buf_8 fanout6085 (.A(net6086),
    .X(net6085));
 sg13g2_buf_8 fanout6086 (.A(net6096),
    .X(net6086));
 sg13g2_buf_8 fanout6087 (.A(net6090),
    .X(net6087));
 sg13g2_buf_2 fanout6088 (.A(net6090),
    .X(net6088));
 sg13g2_buf_8 fanout6089 (.A(net6090),
    .X(net6089));
 sg13g2_buf_8 fanout6090 (.A(net6096),
    .X(net6090));
 sg13g2_buf_8 fanout6091 (.A(net6092),
    .X(net6091));
 sg13g2_buf_8 fanout6092 (.A(net6094),
    .X(net6092));
 sg13g2_buf_8 fanout6093 (.A(net6094),
    .X(net6093));
 sg13g2_buf_8 fanout6094 (.A(net6095),
    .X(net6094));
 sg13g2_buf_2 fanout6095 (.A(net6096),
    .X(net6095));
 sg13g2_buf_8 fanout6096 (.A(net6191),
    .X(net6096));
 sg13g2_buf_8 fanout6097 (.A(net6099),
    .X(net6097));
 sg13g2_buf_1 fanout6098 (.A(net6099),
    .X(net6098));
 sg13g2_buf_8 fanout6099 (.A(net6102),
    .X(net6099));
 sg13g2_buf_8 fanout6100 (.A(net6102),
    .X(net6100));
 sg13g2_buf_8 fanout6101 (.A(net6102),
    .X(net6101));
 sg13g2_buf_8 fanout6102 (.A(net6118),
    .X(net6102));
 sg13g2_buf_8 fanout6103 (.A(net6106),
    .X(net6103));
 sg13g2_buf_8 fanout6104 (.A(net6106),
    .X(net6104));
 sg13g2_buf_8 fanout6105 (.A(net6106),
    .X(net6105));
 sg13g2_buf_8 fanout6106 (.A(net6118),
    .X(net6106));
 sg13g2_buf_8 fanout6107 (.A(net6110),
    .X(net6107));
 sg13g2_buf_8 fanout6108 (.A(net6110),
    .X(net6108));
 sg13g2_buf_1 fanout6109 (.A(net6110),
    .X(net6109));
 sg13g2_buf_8 fanout6110 (.A(net6118),
    .X(net6110));
 sg13g2_buf_8 fanout6111 (.A(net6112),
    .X(net6111));
 sg13g2_buf_2 fanout6112 (.A(net6118),
    .X(net6112));
 sg13g2_buf_8 fanout6113 (.A(net6114),
    .X(net6113));
 sg13g2_buf_8 fanout6114 (.A(net6118),
    .X(net6114));
 sg13g2_buf_8 fanout6115 (.A(net6117),
    .X(net6115));
 sg13g2_buf_8 fanout6116 (.A(net6117),
    .X(net6116));
 sg13g2_buf_8 fanout6117 (.A(net6118),
    .X(net6117));
 sg13g2_buf_8 fanout6118 (.A(net6191),
    .X(net6118));
 sg13g2_buf_8 fanout6119 (.A(net6120),
    .X(net6119));
 sg13g2_buf_8 fanout6120 (.A(net6125),
    .X(net6120));
 sg13g2_buf_8 fanout6121 (.A(net6123),
    .X(net6121));
 sg13g2_buf_1 fanout6122 (.A(net6123),
    .X(net6122));
 sg13g2_buf_1 fanout6123 (.A(net6124),
    .X(net6123));
 sg13g2_buf_8 fanout6124 (.A(net6125),
    .X(net6124));
 sg13g2_buf_8 fanout6125 (.A(net6142),
    .X(net6125));
 sg13g2_buf_8 fanout6126 (.A(net6129),
    .X(net6126));
 sg13g2_buf_8 fanout6127 (.A(net6128),
    .X(net6127));
 sg13g2_buf_8 fanout6128 (.A(net6129),
    .X(net6128));
 sg13g2_buf_8 fanout6129 (.A(net6133),
    .X(net6129));
 sg13g2_buf_8 fanout6130 (.A(net6132),
    .X(net6130));
 sg13g2_buf_1 fanout6131 (.A(net6132),
    .X(net6131));
 sg13g2_buf_8 fanout6132 (.A(net6133),
    .X(net6132));
 sg13g2_buf_2 fanout6133 (.A(net6142),
    .X(net6133));
 sg13g2_buf_8 fanout6134 (.A(net6142),
    .X(net6134));
 sg13g2_buf_1 fanout6135 (.A(net6142),
    .X(net6135));
 sg13g2_buf_8 fanout6136 (.A(net6138),
    .X(net6136));
 sg13g2_buf_2 fanout6137 (.A(net6138),
    .X(net6137));
 sg13g2_buf_8 fanout6138 (.A(net6141),
    .X(net6138));
 sg13g2_buf_8 fanout6139 (.A(net6141),
    .X(net6139));
 sg13g2_buf_8 fanout6140 (.A(net6141),
    .X(net6140));
 sg13g2_buf_8 fanout6141 (.A(net6142),
    .X(net6141));
 sg13g2_buf_8 fanout6142 (.A(net6191),
    .X(net6142));
 sg13g2_buf_8 fanout6143 (.A(net6144),
    .X(net6143));
 sg13g2_buf_2 fanout6144 (.A(net6145),
    .X(net6144));
 sg13g2_buf_8 fanout6145 (.A(net6155),
    .X(net6145));
 sg13g2_buf_8 fanout6146 (.A(net6149),
    .X(net6146));
 sg13g2_buf_1 fanout6147 (.A(net6149),
    .X(net6147));
 sg13g2_buf_8 fanout6148 (.A(net6149),
    .X(net6148));
 sg13g2_buf_8 fanout6149 (.A(net6155),
    .X(net6149));
 sg13g2_buf_8 fanout6150 (.A(net6152),
    .X(net6150));
 sg13g2_buf_8 fanout6151 (.A(net6152),
    .X(net6151));
 sg13g2_buf_8 fanout6152 (.A(net6155),
    .X(net6152));
 sg13g2_buf_8 fanout6153 (.A(net6155),
    .X(net6153));
 sg13g2_buf_1 fanout6154 (.A(net6155),
    .X(net6154));
 sg13g2_buf_8 fanout6155 (.A(net6190),
    .X(net6155));
 sg13g2_buf_8 fanout6156 (.A(net6164),
    .X(net6156));
 sg13g2_buf_8 fanout6157 (.A(net6158),
    .X(net6157));
 sg13g2_buf_8 fanout6158 (.A(net6159),
    .X(net6158));
 sg13g2_buf_8 fanout6159 (.A(net6164),
    .X(net6159));
 sg13g2_buf_8 fanout6160 (.A(net6161),
    .X(net6160));
 sg13g2_buf_2 fanout6161 (.A(net6163),
    .X(net6161));
 sg13g2_buf_8 fanout6162 (.A(net6163),
    .X(net6162));
 sg13g2_buf_1 fanout6163 (.A(net6164),
    .X(net6163));
 sg13g2_buf_8 fanout6164 (.A(net6190),
    .X(net6164));
 sg13g2_buf_8 fanout6165 (.A(net6166),
    .X(net6165));
 sg13g2_buf_8 fanout6166 (.A(net6167),
    .X(net6166));
 sg13g2_buf_8 fanout6167 (.A(net6182),
    .X(net6167));
 sg13g2_buf_8 fanout6168 (.A(net6182),
    .X(net6168));
 sg13g2_buf_2 fanout6169 (.A(net6182),
    .X(net6169));
 sg13g2_buf_8 fanout6170 (.A(net6175),
    .X(net6170));
 sg13g2_buf_8 fanout6171 (.A(net6172),
    .X(net6171));
 sg13g2_buf_2 fanout6172 (.A(net6175),
    .X(net6172));
 sg13g2_buf_8 fanout6173 (.A(net6175),
    .X(net6173));
 sg13g2_buf_1 fanout6174 (.A(net6175),
    .X(net6174));
 sg13g2_buf_8 fanout6175 (.A(net6182),
    .X(net6175));
 sg13g2_buf_8 fanout6176 (.A(net6178),
    .X(net6176));
 sg13g2_buf_1 fanout6177 (.A(net6178),
    .X(net6177));
 sg13g2_buf_1 fanout6178 (.A(net6182),
    .X(net6178));
 sg13g2_buf_8 fanout6179 (.A(net6180),
    .X(net6179));
 sg13g2_buf_8 fanout6180 (.A(net6181),
    .X(net6180));
 sg13g2_buf_8 fanout6181 (.A(net6182),
    .X(net6181));
 sg13g2_buf_8 fanout6182 (.A(net6190),
    .X(net6182));
 sg13g2_buf_8 fanout6183 (.A(net6185),
    .X(net6183));
 sg13g2_buf_8 fanout6184 (.A(net6185),
    .X(net6184));
 sg13g2_buf_8 fanout6185 (.A(net6190),
    .X(net6185));
 sg13g2_buf_8 fanout6186 (.A(net6187),
    .X(net6186));
 sg13g2_buf_8 fanout6187 (.A(net6188),
    .X(net6187));
 sg13g2_buf_8 fanout6188 (.A(net6189),
    .X(net6188));
 sg13g2_buf_8 fanout6189 (.A(net6190),
    .X(net6189));
 sg13g2_buf_8 fanout6190 (.A(net6191),
    .X(net6190));
 sg13g2_buf_8 fanout6191 (.A(_17025_),
    .X(net6191));
 sg13g2_buf_8 fanout6192 (.A(net6193),
    .X(net6192));
 sg13g2_buf_8 fanout6193 (.A(net6204),
    .X(net6193));
 sg13g2_buf_8 fanout6194 (.A(net6196),
    .X(net6194));
 sg13g2_buf_8 fanout6195 (.A(net6196),
    .X(net6195));
 sg13g2_buf_8 fanout6196 (.A(net6204),
    .X(net6196));
 sg13g2_buf_8 fanout6197 (.A(net6198),
    .X(net6197));
 sg13g2_buf_8 fanout6198 (.A(net6204),
    .X(net6198));
 sg13g2_buf_8 fanout6199 (.A(net6200),
    .X(net6199));
 sg13g2_buf_1 fanout6200 (.A(net6204),
    .X(net6200));
 sg13g2_buf_8 fanout6201 (.A(net6202),
    .X(net6201));
 sg13g2_buf_8 fanout6202 (.A(net6204),
    .X(net6202));
 sg13g2_buf_1 fanout6203 (.A(net6204),
    .X(net6203));
 sg13g2_buf_8 fanout6204 (.A(net6273),
    .X(net6204));
 sg13g2_buf_8 fanout6205 (.A(net6212),
    .X(net6205));
 sg13g2_buf_8 fanout6206 (.A(net6212),
    .X(net6206));
 sg13g2_buf_8 fanout6207 (.A(net6208),
    .X(net6207));
 sg13g2_buf_8 fanout6208 (.A(net6212),
    .X(net6208));
 sg13g2_buf_8 fanout6209 (.A(net6211),
    .X(net6209));
 sg13g2_buf_2 fanout6210 (.A(net6211),
    .X(net6210));
 sg13g2_buf_8 fanout6211 (.A(net6212),
    .X(net6211));
 sg13g2_buf_8 fanout6212 (.A(net6273),
    .X(net6212));
 sg13g2_buf_8 fanout6213 (.A(net6216),
    .X(net6213));
 sg13g2_buf_1 fanout6214 (.A(net6216),
    .X(net6214));
 sg13g2_buf_8 fanout6215 (.A(net6216),
    .X(net6215));
 sg13g2_buf_8 fanout6216 (.A(net6231),
    .X(net6216));
 sg13g2_buf_8 fanout6217 (.A(net6218),
    .X(net6217));
 sg13g2_buf_8 fanout6218 (.A(net6231),
    .X(net6218));
 sg13g2_buf_8 fanout6219 (.A(net6220),
    .X(net6219));
 sg13g2_buf_8 fanout6220 (.A(net6222),
    .X(net6220));
 sg13g2_buf_8 fanout6221 (.A(net6222),
    .X(net6221));
 sg13g2_buf_8 fanout6222 (.A(net6231),
    .X(net6222));
 sg13g2_buf_8 fanout6223 (.A(net6224),
    .X(net6223));
 sg13g2_buf_8 fanout6224 (.A(net6227),
    .X(net6224));
 sg13g2_buf_8 fanout6225 (.A(net6227),
    .X(net6225));
 sg13g2_buf_8 fanout6226 (.A(net6227),
    .X(net6226));
 sg13g2_buf_8 fanout6227 (.A(net6230),
    .X(net6227));
 sg13g2_buf_8 fanout6228 (.A(net6230),
    .X(net6228));
 sg13g2_buf_8 fanout6229 (.A(net6230),
    .X(net6229));
 sg13g2_buf_8 fanout6230 (.A(net6231),
    .X(net6230));
 sg13g2_buf_8 fanout6231 (.A(net6273),
    .X(net6231));
 sg13g2_buf_8 fanout6232 (.A(net6234),
    .X(net6232));
 sg13g2_buf_8 fanout6233 (.A(net6234),
    .X(net6233));
 sg13g2_buf_8 fanout6234 (.A(net6240),
    .X(net6234));
 sg13g2_buf_8 fanout6235 (.A(net6238),
    .X(net6235));
 sg13g2_buf_2 fanout6236 (.A(net6238),
    .X(net6236));
 sg13g2_buf_8 fanout6237 (.A(net6238),
    .X(net6237));
 sg13g2_buf_8 fanout6238 (.A(net6240),
    .X(net6238));
 sg13g2_buf_8 fanout6239 (.A(net6240),
    .X(net6239));
 sg13g2_buf_8 fanout6240 (.A(net6272),
    .X(net6240));
 sg13g2_buf_8 fanout6241 (.A(net6242),
    .X(net6241));
 sg13g2_buf_8 fanout6242 (.A(net6249),
    .X(net6242));
 sg13g2_buf_1 fanout6243 (.A(net6249),
    .X(net6243));
 sg13g2_buf_8 fanout6244 (.A(net6246),
    .X(net6244));
 sg13g2_buf_8 fanout6245 (.A(net6246),
    .X(net6245));
 sg13g2_buf_8 fanout6246 (.A(net6249),
    .X(net6246));
 sg13g2_buf_8 fanout6247 (.A(net6248),
    .X(net6247));
 sg13g2_buf_8 fanout6248 (.A(net6249),
    .X(net6248));
 sg13g2_buf_8 fanout6249 (.A(net6272),
    .X(net6249));
 sg13g2_buf_8 fanout6250 (.A(net6252),
    .X(net6250));
 sg13g2_buf_8 fanout6251 (.A(net6252),
    .X(net6251));
 sg13g2_buf_8 fanout6252 (.A(net6259),
    .X(net6252));
 sg13g2_buf_8 fanout6253 (.A(net6256),
    .X(net6253));
 sg13g2_buf_2 fanout6254 (.A(net6256),
    .X(net6254));
 sg13g2_buf_8 fanout6255 (.A(net6256),
    .X(net6255));
 sg13g2_buf_8 fanout6256 (.A(net6259),
    .X(net6256));
 sg13g2_buf_8 fanout6257 (.A(net6258),
    .X(net6257));
 sg13g2_buf_8 fanout6258 (.A(net6259),
    .X(net6258));
 sg13g2_buf_8 fanout6259 (.A(net6272),
    .X(net6259));
 sg13g2_buf_8 fanout6260 (.A(net6261),
    .X(net6260));
 sg13g2_buf_1 fanout6261 (.A(net6271),
    .X(net6261));
 sg13g2_buf_8 fanout6262 (.A(net6264),
    .X(net6262));
 sg13g2_buf_1 fanout6263 (.A(net6264),
    .X(net6263));
 sg13g2_buf_8 fanout6264 (.A(net6271),
    .X(net6264));
 sg13g2_buf_8 fanout6265 (.A(net6266),
    .X(net6265));
 sg13g2_buf_2 fanout6266 (.A(net6271),
    .X(net6266));
 sg13g2_buf_8 fanout6267 (.A(net6270),
    .X(net6267));
 sg13g2_buf_8 fanout6268 (.A(net6270),
    .X(net6268));
 sg13g2_buf_1 fanout6269 (.A(net6270),
    .X(net6269));
 sg13g2_buf_8 fanout6270 (.A(net6271),
    .X(net6270));
 sg13g2_buf_8 fanout6271 (.A(net6272),
    .X(net6271));
 sg13g2_buf_8 fanout6272 (.A(net6273),
    .X(net6272));
 sg13g2_buf_8 fanout6273 (.A(_19821_),
    .X(net6273));
 sg13g2_buf_8 fanout6274 (.A(net6278),
    .X(net6274));
 sg13g2_buf_8 fanout6275 (.A(net6278),
    .X(net6275));
 sg13g2_buf_8 fanout6276 (.A(net6277),
    .X(net6276));
 sg13g2_buf_2 fanout6277 (.A(net6278),
    .X(net6277));
 sg13g2_buf_8 fanout6278 (.A(net6282),
    .X(net6278));
 sg13g2_buf_8 fanout6279 (.A(net6280),
    .X(net6279));
 sg13g2_buf_8 fanout6280 (.A(net6281),
    .X(net6280));
 sg13g2_buf_8 fanout6281 (.A(net6282),
    .X(net6281));
 sg13g2_buf_8 fanout6282 (.A(net6371),
    .X(net6282));
 sg13g2_buf_8 fanout6283 (.A(net6284),
    .X(net6283));
 sg13g2_buf_8 fanout6284 (.A(net6285),
    .X(net6284));
 sg13g2_buf_8 fanout6285 (.A(net6296),
    .X(net6285));
 sg13g2_buf_8 fanout6286 (.A(net6296),
    .X(net6286));
 sg13g2_buf_1 fanout6287 (.A(net6296),
    .X(net6287));
 sg13g2_buf_8 fanout6288 (.A(net6289),
    .X(net6288));
 sg13g2_buf_2 fanout6289 (.A(net6293),
    .X(net6289));
 sg13g2_buf_8 fanout6290 (.A(net6291),
    .X(net6290));
 sg13g2_buf_8 fanout6291 (.A(net6292),
    .X(net6291));
 sg13g2_buf_8 fanout6292 (.A(net6293),
    .X(net6292));
 sg13g2_buf_1 fanout6293 (.A(net6296),
    .X(net6293));
 sg13g2_buf_8 fanout6294 (.A(net6295),
    .X(net6294));
 sg13g2_buf_8 fanout6295 (.A(net6296),
    .X(net6295));
 sg13g2_buf_8 fanout6296 (.A(net6371),
    .X(net6296));
 sg13g2_buf_8 fanout6297 (.A(net6300),
    .X(net6297));
 sg13g2_buf_8 fanout6298 (.A(net6300),
    .X(net6298));
 sg13g2_buf_8 fanout6299 (.A(net6300),
    .X(net6299));
 sg13g2_buf_8 fanout6300 (.A(net6317),
    .X(net6300));
 sg13g2_buf_8 fanout6301 (.A(net6306),
    .X(net6301));
 sg13g2_buf_1 fanout6302 (.A(net6306),
    .X(net6302));
 sg13g2_buf_8 fanout6303 (.A(net6306),
    .X(net6303));
 sg13g2_buf_8 fanout6304 (.A(net6305),
    .X(net6304));
 sg13g2_buf_8 fanout6305 (.A(net6306),
    .X(net6305));
 sg13g2_buf_8 fanout6306 (.A(net6317),
    .X(net6306));
 sg13g2_buf_8 fanout6307 (.A(net6310),
    .X(net6307));
 sg13g2_buf_8 fanout6308 (.A(net6309),
    .X(net6308));
 sg13g2_buf_8 fanout6309 (.A(net6310),
    .X(net6309));
 sg13g2_buf_8 fanout6310 (.A(net6317),
    .X(net6310));
 sg13g2_buf_8 fanout6311 (.A(net6313),
    .X(net6311));
 sg13g2_buf_1 fanout6312 (.A(net6313),
    .X(net6312));
 sg13g2_buf_8 fanout6313 (.A(net6314),
    .X(net6313));
 sg13g2_buf_8 fanout6314 (.A(net6317),
    .X(net6314));
 sg13g2_buf_8 fanout6315 (.A(net6316),
    .X(net6315));
 sg13g2_buf_8 fanout6316 (.A(net6317),
    .X(net6316));
 sg13g2_buf_8 fanout6317 (.A(net6371),
    .X(net6317));
 sg13g2_buf_8 fanout6318 (.A(net6324),
    .X(net6318));
 sg13g2_buf_8 fanout6319 (.A(net6324),
    .X(net6319));
 sg13g2_buf_8 fanout6320 (.A(net6321),
    .X(net6320));
 sg13g2_buf_8 fanout6321 (.A(net6324),
    .X(net6321));
 sg13g2_buf_8 fanout6322 (.A(net6323),
    .X(net6322));
 sg13g2_buf_8 fanout6323 (.A(net6324),
    .X(net6323));
 sg13g2_buf_8 fanout6324 (.A(net6330),
    .X(net6324));
 sg13g2_buf_8 fanout6325 (.A(net6327),
    .X(net6325));
 sg13g2_buf_8 fanout6326 (.A(net6327),
    .X(net6326));
 sg13g2_buf_2 fanout6327 (.A(net6330),
    .X(net6327));
 sg13g2_buf_8 fanout6328 (.A(net6330),
    .X(net6328));
 sg13g2_buf_1 fanout6329 (.A(net6330),
    .X(net6329));
 sg13g2_buf_8 fanout6330 (.A(net6370),
    .X(net6330));
 sg13g2_buf_8 fanout6331 (.A(net6334),
    .X(net6331));
 sg13g2_buf_8 fanout6332 (.A(net6333),
    .X(net6332));
 sg13g2_buf_8 fanout6333 (.A(net6334),
    .X(net6333));
 sg13g2_buf_8 fanout6334 (.A(net6370),
    .X(net6334));
 sg13g2_buf_8 fanout6335 (.A(net6337),
    .X(net6335));
 sg13g2_buf_1 fanout6336 (.A(net6337),
    .X(net6336));
 sg13g2_buf_8 fanout6337 (.A(net6342),
    .X(net6337));
 sg13g2_buf_8 fanout6338 (.A(net6339),
    .X(net6338));
 sg13g2_buf_2 fanout6339 (.A(net6340),
    .X(net6339));
 sg13g2_buf_8 fanout6340 (.A(net6341),
    .X(net6340));
 sg13g2_buf_8 fanout6341 (.A(net6342),
    .X(net6341));
 sg13g2_buf_8 fanout6342 (.A(net6370),
    .X(net6342));
 sg13g2_buf_8 fanout6343 (.A(net6346),
    .X(net6343));
 sg13g2_buf_8 fanout6344 (.A(net6346),
    .X(net6344));
 sg13g2_buf_8 fanout6345 (.A(net6346),
    .X(net6345));
 sg13g2_buf_8 fanout6346 (.A(net6356),
    .X(net6346));
 sg13g2_buf_8 fanout6347 (.A(net6348),
    .X(net6347));
 sg13g2_buf_8 fanout6348 (.A(net6356),
    .X(net6348));
 sg13g2_buf_8 fanout6349 (.A(net6355),
    .X(net6349));
 sg13g2_buf_8 fanout6350 (.A(net6351),
    .X(net6350));
 sg13g2_buf_8 fanout6351 (.A(net6352),
    .X(net6351));
 sg13g2_buf_8 fanout6352 (.A(net6355),
    .X(net6352));
 sg13g2_buf_8 fanout6353 (.A(net6354),
    .X(net6353));
 sg13g2_buf_8 fanout6354 (.A(net6355),
    .X(net6354));
 sg13g2_buf_8 fanout6355 (.A(net6356),
    .X(net6355));
 sg13g2_buf_8 fanout6356 (.A(net6370),
    .X(net6356));
 sg13g2_buf_8 fanout6357 (.A(net6358),
    .X(net6357));
 sg13g2_buf_8 fanout6358 (.A(net6369),
    .X(net6358));
 sg13g2_buf_8 fanout6359 (.A(net6360),
    .X(net6359));
 sg13g2_buf_8 fanout6360 (.A(net6361),
    .X(net6360));
 sg13g2_buf_8 fanout6361 (.A(net6369),
    .X(net6361));
 sg13g2_buf_8 fanout6362 (.A(net6369),
    .X(net6362));
 sg13g2_buf_1 fanout6363 (.A(net6369),
    .X(net6363));
 sg13g2_buf_8 fanout6364 (.A(net6368),
    .X(net6364));
 sg13g2_buf_8 fanout6365 (.A(net6368),
    .X(net6365));
 sg13g2_buf_8 fanout6366 (.A(net6368),
    .X(net6366));
 sg13g2_buf_2 fanout6367 (.A(net6368),
    .X(net6367));
 sg13g2_buf_8 fanout6368 (.A(net6369),
    .X(net6368));
 sg13g2_buf_8 fanout6369 (.A(net6370),
    .X(net6369));
 sg13g2_buf_8 fanout6370 (.A(net6371),
    .X(net6370));
 sg13g2_buf_8 fanout6371 (.A(_19820_),
    .X(net6371));
 sg13g2_buf_8 fanout6372 (.A(net6374),
    .X(net6372));
 sg13g2_buf_1 fanout6373 (.A(net6374),
    .X(net6373));
 sg13g2_buf_1 fanout6374 (.A(net6382),
    .X(net6374));
 sg13g2_buf_8 fanout6375 (.A(net6377),
    .X(net6375));
 sg13g2_buf_8 fanout6376 (.A(net6377),
    .X(net6376));
 sg13g2_buf_8 fanout6377 (.A(net6378),
    .X(net6377));
 sg13g2_buf_2 fanout6378 (.A(net6382),
    .X(net6378));
 sg13g2_buf_8 fanout6379 (.A(net6381),
    .X(net6379));
 sg13g2_buf_8 fanout6380 (.A(net6381),
    .X(net6380));
 sg13g2_buf_8 fanout6381 (.A(net6382),
    .X(net6381));
 sg13g2_buf_8 fanout6382 (.A(net6419),
    .X(net6382));
 sg13g2_buf_8 fanout6383 (.A(net6384),
    .X(net6383));
 sg13g2_buf_8 fanout6384 (.A(net6387),
    .X(net6384));
 sg13g2_buf_8 fanout6385 (.A(net6386),
    .X(net6385));
 sg13g2_buf_8 fanout6386 (.A(net6387),
    .X(net6386));
 sg13g2_buf_8 fanout6387 (.A(net6419),
    .X(net6387));
 sg13g2_buf_8 fanout6388 (.A(net6389),
    .X(net6388));
 sg13g2_buf_8 fanout6389 (.A(net6390),
    .X(net6389));
 sg13g2_buf_8 fanout6390 (.A(net6398),
    .X(net6390));
 sg13g2_buf_8 fanout6391 (.A(net6393),
    .X(net6391));
 sg13g2_buf_8 fanout6392 (.A(net6393),
    .X(net6392));
 sg13g2_buf_8 fanout6393 (.A(net6398),
    .X(net6393));
 sg13g2_buf_8 fanout6394 (.A(net6395),
    .X(net6394));
 sg13g2_buf_8 fanout6395 (.A(net6398),
    .X(net6395));
 sg13g2_buf_8 fanout6396 (.A(net6397),
    .X(net6396));
 sg13g2_buf_8 fanout6397 (.A(net6398),
    .X(net6397));
 sg13g2_buf_8 fanout6398 (.A(net6419),
    .X(net6398));
 sg13g2_buf_8 fanout6399 (.A(net6400),
    .X(net6399));
 sg13g2_buf_8 fanout6400 (.A(net6401),
    .X(net6400));
 sg13g2_buf_8 fanout6401 (.A(net6409),
    .X(net6401));
 sg13g2_buf_8 fanout6402 (.A(net6403),
    .X(net6402));
 sg13g2_buf_8 fanout6403 (.A(net6409),
    .X(net6403));
 sg13g2_buf_8 fanout6404 (.A(net6406),
    .X(net6404));
 sg13g2_buf_8 fanout6405 (.A(net6406),
    .X(net6405));
 sg13g2_buf_8 fanout6406 (.A(net6409),
    .X(net6406));
 sg13g2_buf_8 fanout6407 (.A(net6408),
    .X(net6407));
 sg13g2_buf_8 fanout6408 (.A(net6409),
    .X(net6408));
 sg13g2_buf_8 fanout6409 (.A(net6419),
    .X(net6409));
 sg13g2_buf_8 fanout6410 (.A(net6411),
    .X(net6410));
 sg13g2_buf_8 fanout6411 (.A(net6418),
    .X(net6411));
 sg13g2_buf_8 fanout6412 (.A(net6413),
    .X(net6412));
 sg13g2_buf_8 fanout6413 (.A(net6418),
    .X(net6413));
 sg13g2_buf_8 fanout6414 (.A(net6418),
    .X(net6414));
 sg13g2_buf_8 fanout6415 (.A(net6418),
    .X(net6415));
 sg13g2_buf_8 fanout6416 (.A(net6417),
    .X(net6416));
 sg13g2_buf_1 fanout6417 (.A(net6418),
    .X(net6417));
 sg13g2_buf_8 fanout6418 (.A(net6419),
    .X(net6418));
 sg13g2_buf_8 fanout6419 (.A(_19811_),
    .X(net6419));
 sg13g2_buf_8 fanout6420 (.A(net6421),
    .X(net6420));
 sg13g2_buf_8 fanout6421 (.A(net6422),
    .X(net6421));
 sg13g2_buf_8 fanout6422 (.A(net6431),
    .X(net6422));
 sg13g2_buf_1 fanout6423 (.A(net6431),
    .X(net6423));
 sg13g2_buf_8 fanout6424 (.A(net6425),
    .X(net6424));
 sg13g2_buf_8 fanout6425 (.A(net6427),
    .X(net6425));
 sg13g2_buf_8 fanout6426 (.A(net6427),
    .X(net6426));
 sg13g2_buf_8 fanout6427 (.A(net6431),
    .X(net6427));
 sg13g2_buf_8 fanout6428 (.A(net6430),
    .X(net6428));
 sg13g2_buf_8 fanout6429 (.A(net6430),
    .X(net6429));
 sg13g2_buf_8 fanout6430 (.A(net6431),
    .X(net6430));
 sg13g2_buf_8 fanout6431 (.A(net6474),
    .X(net6431));
 sg13g2_buf_8 fanout6432 (.A(net6445),
    .X(net6432));
 sg13g2_buf_2 fanout6433 (.A(net6445),
    .X(net6433));
 sg13g2_buf_8 fanout6434 (.A(net6438),
    .X(net6434));
 sg13g2_buf_1 fanout6435 (.A(net6438),
    .X(net6435));
 sg13g2_buf_8 fanout6436 (.A(net6438),
    .X(net6436));
 sg13g2_buf_2 fanout6437 (.A(net6438),
    .X(net6437));
 sg13g2_buf_8 fanout6438 (.A(net6445),
    .X(net6438));
 sg13g2_buf_8 fanout6439 (.A(net6445),
    .X(net6439));
 sg13g2_buf_2 fanout6440 (.A(net6445),
    .X(net6440));
 sg13g2_buf_8 fanout6441 (.A(net6444),
    .X(net6441));
 sg13g2_buf_8 fanout6442 (.A(net6444),
    .X(net6442));
 sg13g2_buf_1 fanout6443 (.A(net6444),
    .X(net6443));
 sg13g2_buf_8 fanout6444 (.A(net6445),
    .X(net6444));
 sg13g2_buf_8 fanout6445 (.A(net6474),
    .X(net6445));
 sg13g2_buf_8 fanout6446 (.A(net6450),
    .X(net6446));
 sg13g2_buf_8 fanout6447 (.A(net6449),
    .X(net6447));
 sg13g2_buf_8 fanout6448 (.A(net6449),
    .X(net6448));
 sg13g2_buf_8 fanout6449 (.A(net6450),
    .X(net6449));
 sg13g2_buf_8 fanout6450 (.A(net6456),
    .X(net6450));
 sg13g2_buf_8 fanout6451 (.A(net6453),
    .X(net6451));
 sg13g2_buf_2 fanout6452 (.A(net6453),
    .X(net6452));
 sg13g2_buf_8 fanout6453 (.A(net6456),
    .X(net6453));
 sg13g2_buf_8 fanout6454 (.A(net6455),
    .X(net6454));
 sg13g2_buf_1 fanout6455 (.A(net6456),
    .X(net6455));
 sg13g2_buf_8 fanout6456 (.A(net6474),
    .X(net6456));
 sg13g2_buf_8 fanout6457 (.A(net6459),
    .X(net6457));
 sg13g2_buf_8 fanout6458 (.A(net6459),
    .X(net6458));
 sg13g2_buf_8 fanout6459 (.A(net6473),
    .X(net6459));
 sg13g2_buf_8 fanout6460 (.A(net6461),
    .X(net6460));
 sg13g2_buf_8 fanout6461 (.A(net6462),
    .X(net6461));
 sg13g2_buf_8 fanout6462 (.A(net6466),
    .X(net6462));
 sg13g2_buf_8 fanout6463 (.A(net6464),
    .X(net6463));
 sg13g2_buf_8 fanout6464 (.A(net6465),
    .X(net6464));
 sg13g2_buf_1 fanout6465 (.A(net6466),
    .X(net6465));
 sg13g2_buf_8 fanout6466 (.A(net6473),
    .X(net6466));
 sg13g2_buf_8 fanout6467 (.A(net6473),
    .X(net6467));
 sg13g2_buf_8 fanout6468 (.A(net6473),
    .X(net6468));
 sg13g2_buf_8 fanout6469 (.A(net6470),
    .X(net6469));
 sg13g2_buf_8 fanout6470 (.A(net6472),
    .X(net6470));
 sg13g2_buf_8 fanout6471 (.A(net6472),
    .X(net6471));
 sg13g2_buf_8 fanout6472 (.A(net6473),
    .X(net6472));
 sg13g2_buf_8 fanout6473 (.A(net6474),
    .X(net6473));
 sg13g2_buf_8 fanout6474 (.A(_19811_),
    .X(net6474));
 sg13g2_buf_8 fanout6475 (.A(net6478),
    .X(net6475));
 sg13g2_buf_1 fanout6476 (.A(net6478),
    .X(net6476));
 sg13g2_buf_8 fanout6477 (.A(net6478),
    .X(net6477));
 sg13g2_buf_8 fanout6478 (.A(net6484),
    .X(net6478));
 sg13g2_buf_8 fanout6479 (.A(net6480),
    .X(net6479));
 sg13g2_buf_8 fanout6480 (.A(net6484),
    .X(net6480));
 sg13g2_buf_8 fanout6481 (.A(net6483),
    .X(net6481));
 sg13g2_buf_8 fanout6482 (.A(net6483),
    .X(net6482));
 sg13g2_buf_8 fanout6483 (.A(net6484),
    .X(net6483));
 sg13g2_buf_8 fanout6484 (.A(net6510),
    .X(net6484));
 sg13g2_buf_8 fanout6485 (.A(net6487),
    .X(net6485));
 sg13g2_buf_1 fanout6486 (.A(net6487),
    .X(net6486));
 sg13g2_buf_8 fanout6487 (.A(net6490),
    .X(net6487));
 sg13g2_buf_8 fanout6488 (.A(net6489),
    .X(net6488));
 sg13g2_buf_8 fanout6489 (.A(net6490),
    .X(net6489));
 sg13g2_buf_8 fanout6490 (.A(net6510),
    .X(net6490));
 sg13g2_buf_8 fanout6491 (.A(net6494),
    .X(net6491));
 sg13g2_buf_1 fanout6492 (.A(net6494),
    .X(net6492));
 sg13g2_buf_8 fanout6493 (.A(net6494),
    .X(net6493));
 sg13g2_buf_8 fanout6494 (.A(net6499),
    .X(net6494));
 sg13g2_buf_8 fanout6495 (.A(net6497),
    .X(net6495));
 sg13g2_buf_1 fanout6496 (.A(net6497),
    .X(net6496));
 sg13g2_buf_8 fanout6497 (.A(net6499),
    .X(net6497));
 sg13g2_buf_8 fanout6498 (.A(net6499),
    .X(net6498));
 sg13g2_buf_8 fanout6499 (.A(net6510),
    .X(net6499));
 sg13g2_buf_8 fanout6500 (.A(net6503),
    .X(net6500));
 sg13g2_buf_8 fanout6501 (.A(net6502),
    .X(net6501));
 sg13g2_buf_8 fanout6502 (.A(net6503),
    .X(net6502));
 sg13g2_buf_8 fanout6503 (.A(net6504),
    .X(net6503));
 sg13g2_buf_8 fanout6504 (.A(net6509),
    .X(net6504));
 sg13g2_buf_8 fanout6505 (.A(net6507),
    .X(net6505));
 sg13g2_buf_8 fanout6506 (.A(net6507),
    .X(net6506));
 sg13g2_buf_8 fanout6507 (.A(net6509),
    .X(net6507));
 sg13g2_buf_8 fanout6508 (.A(net6509),
    .X(net6508));
 sg13g2_buf_8 fanout6509 (.A(net6510),
    .X(net6509));
 sg13g2_buf_8 fanout6510 (.A(_19810_),
    .X(net6510));
 sg13g2_buf_8 fanout6511 (.A(net6512),
    .X(net6511));
 sg13g2_buf_8 fanout6512 (.A(net6513),
    .X(net6512));
 sg13g2_buf_8 fanout6513 (.A(net6514),
    .X(net6513));
 sg13g2_buf_8 fanout6514 (.A(net6521),
    .X(net6514));
 sg13g2_buf_8 fanout6515 (.A(net6521),
    .X(net6515));
 sg13g2_buf_2 fanout6516 (.A(net6521),
    .X(net6516));
 sg13g2_buf_8 fanout6517 (.A(net6520),
    .X(net6517));
 sg13g2_buf_8 fanout6518 (.A(net6520),
    .X(net6518));
 sg13g2_buf_8 fanout6519 (.A(net6520),
    .X(net6519));
 sg13g2_buf_8 fanout6520 (.A(net6521),
    .X(net6520));
 sg13g2_buf_8 fanout6521 (.A(net6542),
    .X(net6521));
 sg13g2_buf_2 fanout6522 (.A(net6523),
    .X(net6522));
 sg13g2_buf_2 fanout6523 (.A(net6526),
    .X(net6523));
 sg13g2_buf_2 fanout6524 (.A(net6525),
    .X(net6524));
 sg13g2_buf_1 fanout6525 (.A(net6526),
    .X(net6525));
 sg13g2_buf_1 fanout6526 (.A(net6532),
    .X(net6526));
 sg13g2_buf_8 fanout6527 (.A(net6528),
    .X(net6527));
 sg13g2_buf_8 fanout6528 (.A(net6532),
    .X(net6528));
 sg13g2_buf_8 fanout6529 (.A(net6531),
    .X(net6529));
 sg13g2_buf_1 fanout6530 (.A(net6531),
    .X(net6530));
 sg13g2_buf_1 fanout6531 (.A(net6532),
    .X(net6531));
 sg13g2_buf_8 fanout6532 (.A(net6542),
    .X(net6532));
 sg13g2_buf_2 fanout6533 (.A(net6535),
    .X(net6533));
 sg13g2_buf_8 fanout6534 (.A(net6535),
    .X(net6534));
 sg13g2_buf_8 fanout6535 (.A(net6542),
    .X(net6535));
 sg13g2_buf_8 fanout6536 (.A(net6537),
    .X(net6536));
 sg13g2_buf_1 fanout6537 (.A(net6541),
    .X(net6537));
 sg13g2_buf_8 fanout6538 (.A(net6539),
    .X(net6538));
 sg13g2_buf_8 fanout6539 (.A(net6541),
    .X(net6539));
 sg13g2_buf_2 fanout6540 (.A(net6541),
    .X(net6540));
 sg13g2_buf_8 fanout6541 (.A(net6542),
    .X(net6541));
 sg13g2_buf_8 fanout6542 (.A(net6605),
    .X(net6542));
 sg13g2_buf_8 fanout6543 (.A(net6544),
    .X(net6543));
 sg13g2_buf_1 fanout6544 (.A(net6545),
    .X(net6544));
 sg13g2_buf_1 fanout6545 (.A(net6546),
    .X(net6545));
 sg13g2_buf_8 fanout6546 (.A(net6555),
    .X(net6546));
 sg13g2_buf_8 fanout6547 (.A(net6548),
    .X(net6547));
 sg13g2_buf_8 fanout6548 (.A(net6555),
    .X(net6548));
 sg13g2_buf_8 fanout6549 (.A(net6550),
    .X(net6549));
 sg13g2_buf_8 fanout6550 (.A(net6554),
    .X(net6550));
 sg13g2_buf_8 fanout6551 (.A(net6552),
    .X(net6551));
 sg13g2_buf_8 fanout6552 (.A(net6553),
    .X(net6552));
 sg13g2_buf_8 fanout6553 (.A(net6554),
    .X(net6553));
 sg13g2_buf_8 fanout6554 (.A(net6555),
    .X(net6554));
 sg13g2_buf_8 fanout6555 (.A(net6605),
    .X(net6555));
 sg13g2_buf_8 fanout6556 (.A(net6575),
    .X(net6556));
 sg13g2_buf_8 fanout6557 (.A(net6559),
    .X(net6557));
 sg13g2_buf_1 fanout6558 (.A(net6559),
    .X(net6558));
 sg13g2_buf_8 fanout6559 (.A(net6565),
    .X(net6559));
 sg13g2_buf_8 fanout6560 (.A(net6561),
    .X(net6560));
 sg13g2_buf_8 fanout6561 (.A(net6562),
    .X(net6561));
 sg13g2_buf_8 fanout6562 (.A(net6565),
    .X(net6562));
 sg13g2_buf_8 fanout6563 (.A(net6564),
    .X(net6563));
 sg13g2_buf_1 fanout6564 (.A(net6565),
    .X(net6564));
 sg13g2_buf_8 fanout6565 (.A(net6575),
    .X(net6565));
 sg13g2_buf_2 fanout6566 (.A(net6567),
    .X(net6566));
 sg13g2_buf_1 fanout6567 (.A(net6572),
    .X(net6567));
 sg13g2_buf_8 fanout6568 (.A(net6570),
    .X(net6568));
 sg13g2_buf_1 fanout6569 (.A(net6570),
    .X(net6569));
 sg13g2_buf_1 fanout6570 (.A(net6572),
    .X(net6570));
 sg13g2_buf_8 fanout6571 (.A(net6572),
    .X(net6571));
 sg13g2_buf_2 fanout6572 (.A(net6575),
    .X(net6572));
 sg13g2_buf_8 fanout6573 (.A(net6575),
    .X(net6573));
 sg13g2_buf_1 fanout6574 (.A(net6575),
    .X(net6574));
 sg13g2_buf_8 fanout6575 (.A(net6605),
    .X(net6575));
 sg13g2_buf_8 fanout6576 (.A(net6582),
    .X(net6576));
 sg13g2_buf_8 fanout6577 (.A(net6582),
    .X(net6577));
 sg13g2_buf_8 fanout6578 (.A(net6579),
    .X(net6578));
 sg13g2_buf_8 fanout6579 (.A(net6581),
    .X(net6579));
 sg13g2_buf_8 fanout6580 (.A(net6581),
    .X(net6580));
 sg13g2_buf_8 fanout6581 (.A(net6582),
    .X(net6581));
 sg13g2_buf_8 fanout6582 (.A(net6592),
    .X(net6582));
 sg13g2_buf_2 fanout6583 (.A(net6584),
    .X(net6583));
 sg13g2_buf_1 fanout6584 (.A(net6587),
    .X(net6584));
 sg13g2_buf_2 fanout6585 (.A(net6587),
    .X(net6585));
 sg13g2_buf_1 fanout6586 (.A(net6587),
    .X(net6586));
 sg13g2_buf_2 fanout6587 (.A(net6592),
    .X(net6587));
 sg13g2_buf_2 fanout6588 (.A(net6589),
    .X(net6588));
 sg13g2_buf_8 fanout6589 (.A(net6592),
    .X(net6589));
 sg13g2_buf_8 fanout6590 (.A(net6591),
    .X(net6590));
 sg13g2_buf_8 fanout6591 (.A(net6592),
    .X(net6591));
 sg13g2_buf_8 fanout6592 (.A(net6605),
    .X(net6592));
 sg13g2_buf_2 fanout6593 (.A(net6594),
    .X(net6593));
 sg13g2_buf_8 fanout6594 (.A(net6604),
    .X(net6594));
 sg13g2_buf_8 fanout6595 (.A(net6603),
    .X(net6595));
 sg13g2_buf_8 fanout6596 (.A(net6598),
    .X(net6596));
 sg13g2_buf_1 fanout6597 (.A(net6598),
    .X(net6597));
 sg13g2_buf_2 fanout6598 (.A(net6603),
    .X(net6598));
 sg13g2_buf_8 fanout6599 (.A(net6602),
    .X(net6599));
 sg13g2_buf_8 fanout6600 (.A(net6602),
    .X(net6600));
 sg13g2_buf_8 fanout6601 (.A(net6602),
    .X(net6601));
 sg13g2_buf_8 fanout6602 (.A(net6603),
    .X(net6602));
 sg13g2_buf_8 fanout6603 (.A(net6604),
    .X(net6603));
 sg13g2_buf_8 fanout6604 (.A(net6605),
    .X(net6604));
 sg13g2_buf_8 fanout6605 (.A(_18928_),
    .X(net6605));
 sg13g2_buf_8 fanout6606 (.A(net6608),
    .X(net6606));
 sg13g2_buf_8 fanout6607 (.A(net6608),
    .X(net6607));
 sg13g2_buf_8 fanout6608 (.A(_18629_),
    .X(net6608));
 sg13g2_buf_8 fanout6609 (.A(net6610),
    .X(net6609));
 sg13g2_buf_8 fanout6610 (.A(net6611),
    .X(net6610));
 sg13g2_buf_2 fanout6611 (.A(net6612),
    .X(net6611));
 sg13g2_buf_8 fanout6612 (.A(net6613),
    .X(net6612));
 sg13g2_buf_8 fanout6613 (.A(net6622),
    .X(net6613));
 sg13g2_buf_8 fanout6614 (.A(net6615),
    .X(net6614));
 sg13g2_buf_1 fanout6615 (.A(net6616),
    .X(net6615));
 sg13g2_buf_1 fanout6616 (.A(net6622),
    .X(net6616));
 sg13g2_buf_8 fanout6617 (.A(net6619),
    .X(net6617));
 sg13g2_buf_1 fanout6618 (.A(net6619),
    .X(net6618));
 sg13g2_buf_8 fanout6619 (.A(net6620),
    .X(net6619));
 sg13g2_buf_8 fanout6620 (.A(net6621),
    .X(net6620));
 sg13g2_buf_8 fanout6621 (.A(net6622),
    .X(net6621));
 sg13g2_buf_8 fanout6622 (.A(_14998_),
    .X(net6622));
 sg13g2_buf_8 fanout6623 (.A(net6625),
    .X(net6623));
 sg13g2_buf_8 fanout6624 (.A(net6625),
    .X(net6624));
 sg13g2_buf_8 fanout6625 (.A(net6636),
    .X(net6625));
 sg13g2_buf_8 fanout6626 (.A(net6636),
    .X(net6626));
 sg13g2_buf_8 fanout6627 (.A(net6628),
    .X(net6627));
 sg13g2_buf_8 fanout6628 (.A(net6629),
    .X(net6628));
 sg13g2_buf_8 fanout6629 (.A(net6635),
    .X(net6629));
 sg13g2_buf_8 fanout6630 (.A(net6631),
    .X(net6630));
 sg13g2_buf_8 fanout6631 (.A(net6632),
    .X(net6631));
 sg13g2_buf_8 fanout6632 (.A(net6633),
    .X(net6632));
 sg13g2_buf_8 fanout6633 (.A(net6634),
    .X(net6633));
 sg13g2_buf_2 fanout6634 (.A(net6635),
    .X(net6634));
 sg13g2_buf_8 fanout6635 (.A(net6636),
    .X(net6635));
 sg13g2_buf_8 fanout6636 (.A(_14998_),
    .X(net6636));
 sg13g2_buf_8 fanout6637 (.A(net6640),
    .X(net6637));
 sg13g2_buf_8 fanout6638 (.A(net6640),
    .X(net6638));
 sg13g2_buf_1 fanout6639 (.A(net6640),
    .X(net6639));
 sg13g2_buf_8 fanout6640 (.A(net6651),
    .X(net6640));
 sg13g2_buf_8 fanout6641 (.A(net6644),
    .X(net6641));
 sg13g2_buf_8 fanout6642 (.A(net6644),
    .X(net6642));
 sg13g2_buf_1 fanout6643 (.A(net6644),
    .X(net6643));
 sg13g2_buf_8 fanout6644 (.A(net6651),
    .X(net6644));
 sg13g2_buf_8 fanout6645 (.A(net6647),
    .X(net6645));
 sg13g2_buf_1 fanout6646 (.A(net6647),
    .X(net6646));
 sg13g2_buf_8 fanout6647 (.A(net6651),
    .X(net6647));
 sg13g2_buf_8 fanout6648 (.A(net6650),
    .X(net6648));
 sg13g2_buf_8 fanout6649 (.A(net6650),
    .X(net6649));
 sg13g2_buf_8 fanout6650 (.A(net6651),
    .X(net6650));
 sg13g2_buf_8 fanout6651 (.A(net6675),
    .X(net6651));
 sg13g2_buf_8 fanout6652 (.A(net6654),
    .X(net6652));
 sg13g2_buf_1 fanout6653 (.A(net6654),
    .X(net6653));
 sg13g2_buf_8 fanout6654 (.A(net6655),
    .X(net6654));
 sg13g2_buf_2 fanout6655 (.A(net6656),
    .X(net6655));
 sg13g2_buf_8 fanout6656 (.A(net6675),
    .X(net6656));
 sg13g2_buf_8 fanout6657 (.A(net6660),
    .X(net6657));
 sg13g2_buf_8 fanout6658 (.A(net6660),
    .X(net6658));
 sg13g2_buf_8 fanout6659 (.A(net6660),
    .X(net6659));
 sg13g2_buf_8 fanout6660 (.A(net6675),
    .X(net6660));
 sg13g2_buf_8 fanout6661 (.A(net6674),
    .X(net6661));
 sg13g2_buf_1 fanout6662 (.A(net6674),
    .X(net6662));
 sg13g2_buf_8 fanout6663 (.A(net6667),
    .X(net6663));
 sg13g2_buf_8 fanout6664 (.A(net6665),
    .X(net6664));
 sg13g2_buf_2 fanout6665 (.A(net6667),
    .X(net6665));
 sg13g2_buf_8 fanout6666 (.A(net6667),
    .X(net6666));
 sg13g2_buf_8 fanout6667 (.A(net6674),
    .X(net6667));
 sg13g2_buf_8 fanout6668 (.A(net6671),
    .X(net6668));
 sg13g2_buf_8 fanout6669 (.A(net6671),
    .X(net6669));
 sg13g2_buf_8 fanout6670 (.A(net6671),
    .X(net6670));
 sg13g2_buf_8 fanout6671 (.A(net6672),
    .X(net6671));
 sg13g2_buf_8 fanout6672 (.A(net6673),
    .X(net6672));
 sg13g2_buf_1 fanout6673 (.A(net6674),
    .X(net6673));
 sg13g2_buf_8 fanout6674 (.A(net6675),
    .X(net6674));
 sg13g2_buf_8 fanout6675 (.A(_18945_),
    .X(net6675));
 sg13g2_buf_8 fanout6676 (.A(_18908_),
    .X(net6676));
 sg13g2_buf_8 fanout6677 (.A(_18632_),
    .X(net6677));
 sg13g2_buf_8 fanout6678 (.A(net6680),
    .X(net6678));
 sg13g2_buf_8 fanout6679 (.A(net6680),
    .X(net6679));
 sg13g2_buf_8 fanout6680 (.A(net6681),
    .X(net6680));
 sg13g2_buf_8 fanout6681 (.A(net6696),
    .X(net6681));
 sg13g2_buf_8 fanout6682 (.A(net6684),
    .X(net6682));
 sg13g2_buf_1 fanout6683 (.A(net6684),
    .X(net6683));
 sg13g2_buf_8 fanout6684 (.A(net6685),
    .X(net6684));
 sg13g2_buf_8 fanout6685 (.A(net6696),
    .X(net6685));
 sg13g2_buf_8 fanout6686 (.A(net6688),
    .X(net6686));
 sg13g2_buf_1 fanout6687 (.A(net6688),
    .X(net6687));
 sg13g2_buf_8 fanout6688 (.A(net6689),
    .X(net6688));
 sg13g2_buf_1 fanout6689 (.A(net6696),
    .X(net6689));
 sg13g2_buf_8 fanout6690 (.A(net6691),
    .X(net6690));
 sg13g2_buf_8 fanout6691 (.A(net6692),
    .X(net6691));
 sg13g2_buf_1 fanout6692 (.A(net6695),
    .X(net6692));
 sg13g2_buf_8 fanout6693 (.A(net6694),
    .X(net6693));
 sg13g2_buf_8 fanout6694 (.A(net6695),
    .X(net6694));
 sg13g2_buf_8 fanout6695 (.A(net6696),
    .X(net6695));
 sg13g2_buf_8 fanout6696 (.A(net6745),
    .X(net6696));
 sg13g2_buf_8 fanout6697 (.A(net6703),
    .X(net6697));
 sg13g2_buf_1 fanout6698 (.A(net6703),
    .X(net6698));
 sg13g2_buf_8 fanout6699 (.A(net6701),
    .X(net6699));
 sg13g2_buf_2 fanout6700 (.A(net6701),
    .X(net6700));
 sg13g2_buf_8 fanout6701 (.A(net6703),
    .X(net6701));
 sg13g2_buf_8 fanout6702 (.A(net6703),
    .X(net6702));
 sg13g2_buf_8 fanout6703 (.A(net6745),
    .X(net6703));
 sg13g2_buf_8 fanout6704 (.A(net6706),
    .X(net6704));
 sg13g2_buf_1 fanout6705 (.A(net6706),
    .X(net6705));
 sg13g2_buf_8 fanout6706 (.A(net6710),
    .X(net6706));
 sg13g2_buf_8 fanout6707 (.A(net6710),
    .X(net6707));
 sg13g2_buf_1 fanout6708 (.A(net6710),
    .X(net6708));
 sg13g2_buf_8 fanout6709 (.A(net6710),
    .X(net6709));
 sg13g2_buf_8 fanout6710 (.A(net6745),
    .X(net6710));
 sg13g2_buf_8 fanout6711 (.A(net6715),
    .X(net6711));
 sg13g2_buf_8 fanout6712 (.A(net6713),
    .X(net6712));
 sg13g2_buf_8 fanout6713 (.A(net6714),
    .X(net6713));
 sg13g2_buf_8 fanout6714 (.A(net6715),
    .X(net6714));
 sg13g2_buf_8 fanout6715 (.A(net6744),
    .X(net6715));
 sg13g2_buf_8 fanout6716 (.A(net6717),
    .X(net6716));
 sg13g2_buf_8 fanout6717 (.A(net6718),
    .X(net6717));
 sg13g2_buf_2 fanout6718 (.A(net6719),
    .X(net6718));
 sg13g2_buf_2 fanout6719 (.A(net6720),
    .X(net6719));
 sg13g2_buf_1 fanout6720 (.A(net6724),
    .X(net6720));
 sg13g2_buf_8 fanout6721 (.A(net6724),
    .X(net6721));
 sg13g2_buf_8 fanout6722 (.A(net6723),
    .X(net6722));
 sg13g2_buf_2 fanout6723 (.A(net6724),
    .X(net6723));
 sg13g2_buf_8 fanout6724 (.A(net6744),
    .X(net6724));
 sg13g2_buf_8 fanout6725 (.A(net6726),
    .X(net6725));
 sg13g2_buf_2 fanout6726 (.A(net6727),
    .X(net6726));
 sg13g2_buf_8 fanout6727 (.A(net6736),
    .X(net6727));
 sg13g2_buf_8 fanout6728 (.A(net6729),
    .X(net6728));
 sg13g2_buf_8 fanout6729 (.A(net6736),
    .X(net6729));
 sg13g2_buf_2 fanout6730 (.A(net6731),
    .X(net6730));
 sg13g2_buf_1 fanout6731 (.A(net6735),
    .X(net6731));
 sg13g2_buf_8 fanout6732 (.A(net6733),
    .X(net6732));
 sg13g2_buf_2 fanout6733 (.A(net6735),
    .X(net6733));
 sg13g2_buf_8 fanout6734 (.A(net6735),
    .X(net6734));
 sg13g2_buf_1 fanout6735 (.A(net6736),
    .X(net6735));
 sg13g2_buf_8 fanout6736 (.A(net6744),
    .X(net6736));
 sg13g2_buf_8 fanout6737 (.A(net6738),
    .X(net6737));
 sg13g2_buf_2 fanout6738 (.A(net6739),
    .X(net6738));
 sg13g2_buf_1 fanout6739 (.A(net6744),
    .X(net6739));
 sg13g2_buf_8 fanout6740 (.A(net6741),
    .X(net6740));
 sg13g2_buf_2 fanout6741 (.A(net6742),
    .X(net6741));
 sg13g2_buf_1 fanout6742 (.A(net6743),
    .X(net6742));
 sg13g2_buf_8 fanout6743 (.A(net6744),
    .X(net6743));
 sg13g2_buf_8 fanout6744 (.A(net6745),
    .X(net6744));
 sg13g2_buf_8 fanout6745 (.A(_14997_),
    .X(net6745));
 sg13g2_buf_8 fanout6746 (.A(net6758),
    .X(net6746));
 sg13g2_buf_8 fanout6747 (.A(net6748),
    .X(net6747));
 sg13g2_buf_2 fanout6748 (.A(net6749),
    .X(net6748));
 sg13g2_buf_1 fanout6749 (.A(net6752),
    .X(net6749));
 sg13g2_buf_8 fanout6750 (.A(net6752),
    .X(net6750));
 sg13g2_buf_8 fanout6751 (.A(net6752),
    .X(net6751));
 sg13g2_buf_8 fanout6752 (.A(net6758),
    .X(net6752));
 sg13g2_buf_8 fanout6753 (.A(net6754),
    .X(net6753));
 sg13g2_buf_8 fanout6754 (.A(net6756),
    .X(net6754));
 sg13g2_buf_8 fanout6755 (.A(net6756),
    .X(net6755));
 sg13g2_buf_8 fanout6756 (.A(net6757),
    .X(net6756));
 sg13g2_buf_8 fanout6757 (.A(net6758),
    .X(net6757));
 sg13g2_buf_8 fanout6758 (.A(net6787),
    .X(net6758));
 sg13g2_buf_8 fanout6759 (.A(net6760),
    .X(net6759));
 sg13g2_buf_8 fanout6760 (.A(net6764),
    .X(net6760));
 sg13g2_buf_8 fanout6761 (.A(net6764),
    .X(net6761));
 sg13g2_buf_1 fanout6762 (.A(net6764),
    .X(net6762));
 sg13g2_buf_8 fanout6763 (.A(net6764),
    .X(net6763));
 sg13g2_buf_8 fanout6764 (.A(net6787),
    .X(net6764));
 sg13g2_buf_8 fanout6765 (.A(net6767),
    .X(net6765));
 sg13g2_buf_1 fanout6766 (.A(net6767),
    .X(net6766));
 sg13g2_buf_2 fanout6767 (.A(net6769),
    .X(net6767));
 sg13g2_buf_8 fanout6768 (.A(net6769),
    .X(net6768));
 sg13g2_buf_2 fanout6769 (.A(net6787),
    .X(net6769));
 sg13g2_buf_8 fanout6770 (.A(net6773),
    .X(net6770));
 sg13g2_buf_1 fanout6771 (.A(net6773),
    .X(net6771));
 sg13g2_buf_8 fanout6772 (.A(net6773),
    .X(net6772));
 sg13g2_buf_8 fanout6773 (.A(net6777),
    .X(net6773));
 sg13g2_buf_8 fanout6774 (.A(net6777),
    .X(net6774));
 sg13g2_buf_8 fanout6775 (.A(net6777),
    .X(net6775));
 sg13g2_buf_8 fanout6776 (.A(net6777),
    .X(net6776));
 sg13g2_buf_8 fanout6777 (.A(net6787),
    .X(net6777));
 sg13g2_buf_8 fanout6778 (.A(net6781),
    .X(net6778));
 sg13g2_buf_8 fanout6779 (.A(net6781),
    .X(net6779));
 sg13g2_buf_2 fanout6780 (.A(net6781),
    .X(net6780));
 sg13g2_buf_8 fanout6781 (.A(net6786),
    .X(net6781));
 sg13g2_buf_8 fanout6782 (.A(net6783),
    .X(net6782));
 sg13g2_buf_8 fanout6783 (.A(net6784),
    .X(net6783));
 sg13g2_buf_8 fanout6784 (.A(net6786),
    .X(net6784));
 sg13g2_buf_8 fanout6785 (.A(net6786),
    .X(net6785));
 sg13g2_buf_8 fanout6786 (.A(net6787),
    .X(net6786));
 sg13g2_buf_8 fanout6787 (.A(_03354_),
    .X(net6787));
 sg13g2_buf_8 fanout6788 (.A(net6789),
    .X(net6788));
 sg13g2_buf_8 fanout6789 (.A(net6790),
    .X(net6789));
 sg13g2_buf_8 fanout6790 (.A(net6815),
    .X(net6790));
 sg13g2_buf_8 fanout6791 (.A(net6793),
    .X(net6791));
 sg13g2_buf_1 fanout6792 (.A(net6793),
    .X(net6792));
 sg13g2_buf_8 fanout6793 (.A(net6795),
    .X(net6793));
 sg13g2_buf_8 fanout6794 (.A(net6795),
    .X(net6794));
 sg13g2_buf_8 fanout6795 (.A(net6815),
    .X(net6795));
 sg13g2_buf_8 fanout6796 (.A(net6800),
    .X(net6796));
 sg13g2_buf_8 fanout6797 (.A(net6800),
    .X(net6797));
 sg13g2_buf_8 fanout6798 (.A(net6800),
    .X(net6798));
 sg13g2_buf_2 fanout6799 (.A(net6800),
    .X(net6799));
 sg13g2_buf_8 fanout6800 (.A(net6801),
    .X(net6800));
 sg13g2_buf_8 fanout6801 (.A(net6815),
    .X(net6801));
 sg13g2_buf_8 fanout6802 (.A(net6803),
    .X(net6802));
 sg13g2_buf_8 fanout6803 (.A(net6815),
    .X(net6803));
 sg13g2_buf_8 fanout6804 (.A(net6808),
    .X(net6804));
 sg13g2_buf_1 fanout6805 (.A(net6808),
    .X(net6805));
 sg13g2_buf_8 fanout6806 (.A(net6808),
    .X(net6806));
 sg13g2_buf_8 fanout6807 (.A(net6808),
    .X(net6807));
 sg13g2_buf_8 fanout6808 (.A(net6815),
    .X(net6808));
 sg13g2_buf_8 fanout6809 (.A(net6814),
    .X(net6809));
 sg13g2_buf_8 fanout6810 (.A(net6811),
    .X(net6810));
 sg13g2_buf_1 fanout6811 (.A(net6813),
    .X(net6811));
 sg13g2_buf_8 fanout6812 (.A(net6813),
    .X(net6812));
 sg13g2_buf_2 fanout6813 (.A(net6814),
    .X(net6813));
 sg13g2_buf_8 fanout6814 (.A(net6815),
    .X(net6814));
 sg13g2_buf_8 fanout6815 (.A(net6835),
    .X(net6815));
 sg13g2_buf_8 fanout6816 (.A(net6820),
    .X(net6816));
 sg13g2_buf_8 fanout6817 (.A(net6820),
    .X(net6817));
 sg13g2_buf_8 fanout6818 (.A(net6819),
    .X(net6818));
 sg13g2_buf_8 fanout6819 (.A(net6820),
    .X(net6819));
 sg13g2_buf_8 fanout6820 (.A(net6835),
    .X(net6820));
 sg13g2_buf_8 fanout6821 (.A(net6823),
    .X(net6821));
 sg13g2_buf_8 fanout6822 (.A(net6823),
    .X(net6822));
 sg13g2_buf_8 fanout6823 (.A(net6835),
    .X(net6823));
 sg13g2_buf_8 fanout6824 (.A(net6827),
    .X(net6824));
 sg13g2_buf_8 fanout6825 (.A(net6826),
    .X(net6825));
 sg13g2_buf_8 fanout6826 (.A(net6827),
    .X(net6826));
 sg13g2_buf_8 fanout6827 (.A(net6834),
    .X(net6827));
 sg13g2_buf_8 fanout6828 (.A(net6829),
    .X(net6828));
 sg13g2_buf_8 fanout6829 (.A(net6830),
    .X(net6829));
 sg13g2_buf_2 fanout6830 (.A(net6834),
    .X(net6830));
 sg13g2_buf_8 fanout6831 (.A(net6832),
    .X(net6831));
 sg13g2_buf_8 fanout6832 (.A(net6833),
    .X(net6832));
 sg13g2_buf_8 fanout6833 (.A(net6834),
    .X(net6833));
 sg13g2_buf_8 fanout6834 (.A(net6835),
    .X(net6834));
 sg13g2_buf_8 fanout6835 (.A(_03353_),
    .X(net6835));
 sg13g2_buf_8 fanout6836 (.A(net6841),
    .X(net6836));
 sg13g2_buf_8 fanout6837 (.A(net6840),
    .X(net6837));
 sg13g2_buf_8 fanout6838 (.A(net6840),
    .X(net6838));
 sg13g2_buf_8 fanout6839 (.A(net6840),
    .X(net6839));
 sg13g2_buf_8 fanout6840 (.A(net6841),
    .X(net6840));
 sg13g2_buf_8 fanout6841 (.A(net6865),
    .X(net6841));
 sg13g2_buf_8 fanout6842 (.A(net6844),
    .X(net6842));
 sg13g2_buf_8 fanout6843 (.A(net6844),
    .X(net6843));
 sg13g2_buf_8 fanout6844 (.A(net6865),
    .X(net6844));
 sg13g2_buf_8 fanout6845 (.A(net6849),
    .X(net6845));
 sg13g2_buf_8 fanout6846 (.A(net6849),
    .X(net6846));
 sg13g2_buf_8 fanout6847 (.A(net6849),
    .X(net6847));
 sg13g2_buf_1 fanout6848 (.A(net6849),
    .X(net6848));
 sg13g2_buf_8 fanout6849 (.A(net6865),
    .X(net6849));
 sg13g2_buf_8 fanout6850 (.A(net6858),
    .X(net6850));
 sg13g2_buf_8 fanout6851 (.A(net6853),
    .X(net6851));
 sg13g2_buf_1 fanout6852 (.A(net6853),
    .X(net6852));
 sg13g2_buf_8 fanout6853 (.A(net6858),
    .X(net6853));
 sg13g2_buf_8 fanout6854 (.A(net6858),
    .X(net6854));
 sg13g2_buf_8 fanout6855 (.A(net6856),
    .X(net6855));
 sg13g2_buf_8 fanout6856 (.A(net6857),
    .X(net6856));
 sg13g2_buf_8 fanout6857 (.A(net6858),
    .X(net6857));
 sg13g2_buf_8 fanout6858 (.A(net6865),
    .X(net6858));
 sg13g2_buf_8 fanout6859 (.A(net6864),
    .X(net6859));
 sg13g2_buf_8 fanout6860 (.A(net6861),
    .X(net6860));
 sg13g2_buf_8 fanout6861 (.A(net6862),
    .X(net6861));
 sg13g2_buf_8 fanout6862 (.A(net6863),
    .X(net6862));
 sg13g2_buf_8 fanout6863 (.A(net6864),
    .X(net6863));
 sg13g2_buf_8 fanout6864 (.A(net6865),
    .X(net6864));
 sg13g2_buf_8 fanout6865 (.A(_02348_),
    .X(net6865));
 sg13g2_buf_8 fanout6866 (.A(net6871),
    .X(net6866));
 sg13g2_buf_8 fanout6867 (.A(net6868),
    .X(net6867));
 sg13g2_buf_8 fanout6868 (.A(net6871),
    .X(net6868));
 sg13g2_buf_1 fanout6869 (.A(net6870),
    .X(net6869));
 sg13g2_buf_8 fanout6870 (.A(net6871),
    .X(net6870));
 sg13g2_buf_8 fanout6871 (.A(net6890),
    .X(net6871));
 sg13g2_buf_8 fanout6872 (.A(net6873),
    .X(net6872));
 sg13g2_buf_8 fanout6873 (.A(net6875),
    .X(net6873));
 sg13g2_buf_8 fanout6874 (.A(net6875),
    .X(net6874));
 sg13g2_buf_8 fanout6875 (.A(net6879),
    .X(net6875));
 sg13g2_buf_8 fanout6876 (.A(net6879),
    .X(net6876));
 sg13g2_buf_1 fanout6877 (.A(net6879),
    .X(net6877));
 sg13g2_buf_8 fanout6878 (.A(net6879),
    .X(net6878));
 sg13g2_buf_8 fanout6879 (.A(net6890),
    .X(net6879));
 sg13g2_buf_8 fanout6880 (.A(net6883),
    .X(net6880));
 sg13g2_buf_8 fanout6881 (.A(net6883),
    .X(net6881));
 sg13g2_buf_8 fanout6882 (.A(net6883),
    .X(net6882));
 sg13g2_buf_8 fanout6883 (.A(net6890),
    .X(net6883));
 sg13g2_buf_8 fanout6884 (.A(net6885),
    .X(net6884));
 sg13g2_buf_8 fanout6885 (.A(net6888),
    .X(net6885));
 sg13g2_buf_8 fanout6886 (.A(net6888),
    .X(net6886));
 sg13g2_buf_8 fanout6887 (.A(net6888),
    .X(net6887));
 sg13g2_buf_8 fanout6888 (.A(net6889),
    .X(net6888));
 sg13g2_buf_8 fanout6889 (.A(net6890),
    .X(net6889));
 sg13g2_buf_8 fanout6890 (.A(_02347_),
    .X(net6890));
 sg13g2_buf_8 fanout6891 (.A(net6896),
    .X(net6891));
 sg13g2_buf_1 fanout6892 (.A(net6896),
    .X(net6892));
 sg13g2_buf_8 fanout6893 (.A(net6895),
    .X(net6893));
 sg13g2_buf_1 fanout6894 (.A(net6895),
    .X(net6894));
 sg13g2_buf_8 fanout6895 (.A(net6896),
    .X(net6895));
 sg13g2_buf_8 fanout6896 (.A(net6908),
    .X(net6896));
 sg13g2_buf_8 fanout6897 (.A(net6899),
    .X(net6897));
 sg13g2_buf_2 fanout6898 (.A(net6899),
    .X(net6898));
 sg13g2_buf_8 fanout6899 (.A(net6902),
    .X(net6899));
 sg13g2_buf_8 fanout6900 (.A(net6901),
    .X(net6900));
 sg13g2_buf_2 fanout6901 (.A(net6902),
    .X(net6901));
 sg13g2_buf_8 fanout6902 (.A(net6903),
    .X(net6902));
 sg13g2_buf_8 fanout6903 (.A(net6908),
    .X(net6903));
 sg13g2_buf_8 fanout6904 (.A(net6905),
    .X(net6904));
 sg13g2_buf_8 fanout6905 (.A(net6907),
    .X(net6905));
 sg13g2_buf_8 fanout6906 (.A(net6907),
    .X(net6906));
 sg13g2_buf_8 fanout6907 (.A(net6908),
    .X(net6907));
 sg13g2_buf_8 fanout6908 (.A(net6915),
    .X(net6908));
 sg13g2_buf_8 fanout6909 (.A(net6910),
    .X(net6909));
 sg13g2_buf_8 fanout6910 (.A(net6911),
    .X(net6910));
 sg13g2_buf_8 fanout6911 (.A(net6915),
    .X(net6911));
 sg13g2_buf_8 fanout6912 (.A(net6913),
    .X(net6912));
 sg13g2_buf_8 fanout6913 (.A(net6914),
    .X(net6913));
 sg13g2_buf_8 fanout6914 (.A(net6915),
    .X(net6914));
 sg13g2_buf_8 fanout6915 (.A(net6939),
    .X(net6915));
 sg13g2_buf_8 fanout6916 (.A(net6917),
    .X(net6916));
 sg13g2_buf_1 fanout6917 (.A(net6920),
    .X(net6917));
 sg13g2_buf_8 fanout6918 (.A(net6919),
    .X(net6918));
 sg13g2_buf_8 fanout6919 (.A(net6920),
    .X(net6919));
 sg13g2_buf_8 fanout6920 (.A(net6939),
    .X(net6920));
 sg13g2_buf_8 fanout6921 (.A(net6924),
    .X(net6921));
 sg13g2_buf_8 fanout6922 (.A(net6924),
    .X(net6922));
 sg13g2_buf_8 fanout6923 (.A(net6924),
    .X(net6923));
 sg13g2_buf_8 fanout6924 (.A(net6939),
    .X(net6924));
 sg13g2_buf_8 fanout6925 (.A(net6927),
    .X(net6925));
 sg13g2_buf_8 fanout6926 (.A(net6938),
    .X(net6926));
 sg13g2_buf_8 fanout6927 (.A(net6938),
    .X(net6927));
 sg13g2_buf_8 fanout6928 (.A(net6929),
    .X(net6928));
 sg13g2_buf_8 fanout6929 (.A(net6930),
    .X(net6929));
 sg13g2_buf_8 fanout6930 (.A(net6931),
    .X(net6930));
 sg13g2_buf_8 fanout6931 (.A(net6938),
    .X(net6931));
 sg13g2_buf_8 fanout6932 (.A(net6937),
    .X(net6932));
 sg13g2_buf_8 fanout6933 (.A(net6934),
    .X(net6933));
 sg13g2_buf_8 fanout6934 (.A(net6937),
    .X(net6934));
 sg13g2_buf_8 fanout6935 (.A(net6937),
    .X(net6935));
 sg13g2_buf_1 fanout6936 (.A(net6937),
    .X(net6936));
 sg13g2_buf_8 fanout6937 (.A(net6938),
    .X(net6937));
 sg13g2_buf_8 fanout6938 (.A(net6939),
    .X(net6938));
 sg13g2_buf_8 fanout6939 (.A(_18903_),
    .X(net6939));
 sg13g2_buf_8 fanout6940 (.A(net6941),
    .X(net6940));
 sg13g2_buf_8 fanout6941 (.A(net6943),
    .X(net6941));
 sg13g2_buf_8 fanout6942 (.A(net6943),
    .X(net6942));
 sg13g2_buf_8 fanout6943 (.A(_18902_),
    .X(net6943));
 sg13g2_buf_8 fanout6944 (.A(net6945),
    .X(net6944));
 sg13g2_buf_8 fanout6945 (.A(_18902_),
    .X(net6945));
 sg13g2_buf_8 fanout6946 (.A(net6947),
    .X(net6946));
 sg13g2_buf_8 fanout6947 (.A(net6950),
    .X(net6947));
 sg13g2_buf_8 fanout6948 (.A(net6950),
    .X(net6948));
 sg13g2_buf_8 fanout6949 (.A(net6950),
    .X(net6949));
 sg13g2_buf_8 fanout6950 (.A(net6957),
    .X(net6950));
 sg13g2_buf_8 fanout6951 (.A(net6957),
    .X(net6951));
 sg13g2_buf_1 fanout6952 (.A(net6957),
    .X(net6952));
 sg13g2_buf_8 fanout6953 (.A(net6957),
    .X(net6953));
 sg13g2_buf_8 fanout6954 (.A(net6957),
    .X(net6954));
 sg13g2_buf_8 fanout6955 (.A(net6956),
    .X(net6955));
 sg13g2_buf_8 fanout6956 (.A(net6957),
    .X(net6956));
 sg13g2_buf_8 fanout6957 (.A(net6967),
    .X(net6957));
 sg13g2_buf_8 fanout6958 (.A(net6961),
    .X(net6958));
 sg13g2_buf_8 fanout6959 (.A(net6961),
    .X(net6959));
 sg13g2_buf_8 fanout6960 (.A(net6961),
    .X(net6960));
 sg13g2_buf_8 fanout6961 (.A(net6967),
    .X(net6961));
 sg13g2_buf_8 fanout6962 (.A(net6964),
    .X(net6962));
 sg13g2_buf_8 fanout6963 (.A(net6964),
    .X(net6963));
 sg13g2_buf_8 fanout6964 (.A(net6967),
    .X(net6964));
 sg13g2_buf_8 fanout6965 (.A(net6966),
    .X(net6965));
 sg13g2_buf_8 fanout6966 (.A(net6967),
    .X(net6966));
 sg13g2_buf_8 fanout6967 (.A(net6992),
    .X(net6967));
 sg13g2_buf_8 fanout6968 (.A(net6969),
    .X(net6968));
 sg13g2_buf_8 fanout6969 (.A(net6971),
    .X(net6969));
 sg13g2_buf_8 fanout6970 (.A(net6971),
    .X(net6970));
 sg13g2_buf_8 fanout6971 (.A(net6972),
    .X(net6971));
 sg13g2_buf_8 fanout6972 (.A(net6992),
    .X(net6972));
 sg13g2_buf_8 fanout6973 (.A(net6974),
    .X(net6973));
 sg13g2_buf_8 fanout6974 (.A(net6975),
    .X(net6974));
 sg13g2_buf_8 fanout6975 (.A(net6976),
    .X(net6975));
 sg13g2_buf_8 fanout6976 (.A(net6992),
    .X(net6976));
 sg13g2_buf_8 fanout6977 (.A(net6981),
    .X(net6977));
 sg13g2_buf_8 fanout6978 (.A(net6980),
    .X(net6978));
 sg13g2_buf_8 fanout6979 (.A(net6980),
    .X(net6979));
 sg13g2_buf_8 fanout6980 (.A(net6981),
    .X(net6980));
 sg13g2_buf_8 fanout6981 (.A(net6991),
    .X(net6981));
 sg13g2_buf_8 fanout6982 (.A(net6983),
    .X(net6982));
 sg13g2_buf_8 fanout6983 (.A(net6984),
    .X(net6983));
 sg13g2_buf_8 fanout6984 (.A(net6991),
    .X(net6984));
 sg13g2_buf_8 fanout6985 (.A(net6987),
    .X(net6985));
 sg13g2_buf_8 fanout6986 (.A(net6987),
    .X(net6986));
 sg13g2_buf_8 fanout6987 (.A(net6991),
    .X(net6987));
 sg13g2_buf_8 fanout6988 (.A(net6990),
    .X(net6988));
 sg13g2_buf_8 fanout6989 (.A(net6991),
    .X(net6989));
 sg13g2_buf_8 fanout6990 (.A(net6991),
    .X(net6990));
 sg13g2_buf_8 fanout6991 (.A(net6992),
    .X(net6991));
 sg13g2_buf_8 fanout6992 (.A(_18638_),
    .X(net6992));
 sg13g2_buf_8 fanout6993 (.A(_18621_),
    .X(net6993));
 sg13g2_buf_8 fanout6994 (.A(_04521_),
    .X(net6994));
 sg13g2_buf_8 fanout6995 (.A(_04361_),
    .X(net6995));
 sg13g2_buf_8 fanout6996 (.A(net6997),
    .X(net6996));
 sg13g2_buf_8 fanout6997 (.A(net7007),
    .X(net6997));
 sg13g2_buf_8 fanout6998 (.A(net7002),
    .X(net6998));
 sg13g2_buf_1 fanout6999 (.A(net7002),
    .X(net6999));
 sg13g2_buf_8 fanout7000 (.A(net7002),
    .X(net7000));
 sg13g2_buf_1 fanout7001 (.A(net7002),
    .X(net7001));
 sg13g2_buf_8 fanout7002 (.A(net7007),
    .X(net7002));
 sg13g2_buf_8 fanout7003 (.A(net7005),
    .X(net7003));
 sg13g2_buf_8 fanout7004 (.A(net7005),
    .X(net7004));
 sg13g2_buf_8 fanout7005 (.A(net7007),
    .X(net7005));
 sg13g2_buf_8 fanout7006 (.A(net7007),
    .X(net7006));
 sg13g2_buf_8 fanout7007 (.A(net7023),
    .X(net7007));
 sg13g2_buf_8 fanout7008 (.A(net7010),
    .X(net7008));
 sg13g2_buf_8 fanout7009 (.A(net7010),
    .X(net7009));
 sg13g2_buf_8 fanout7010 (.A(net7015),
    .X(net7010));
 sg13g2_buf_8 fanout7011 (.A(net7015),
    .X(net7011));
 sg13g2_buf_1 fanout7012 (.A(net7015),
    .X(net7012));
 sg13g2_buf_8 fanout7013 (.A(net7014),
    .X(net7013));
 sg13g2_buf_8 fanout7014 (.A(net7015),
    .X(net7014));
 sg13g2_buf_8 fanout7015 (.A(net7016),
    .X(net7015));
 sg13g2_buf_8 fanout7016 (.A(net7023),
    .X(net7016));
 sg13g2_buf_8 fanout7017 (.A(net7022),
    .X(net7017));
 sg13g2_buf_2 fanout7018 (.A(net7019),
    .X(net7018));
 sg13g2_buf_8 fanout7019 (.A(net7022),
    .X(net7019));
 sg13g2_buf_8 fanout7020 (.A(net7021),
    .X(net7020));
 sg13g2_buf_8 fanout7021 (.A(net7022),
    .X(net7021));
 sg13g2_buf_8 fanout7022 (.A(net7023),
    .X(net7022));
 sg13g2_buf_8 fanout7023 (.A(_19807_),
    .X(net7023));
 sg13g2_buf_8 fanout7024 (.A(net7027),
    .X(net7024));
 sg13g2_buf_8 fanout7025 (.A(net7027),
    .X(net7025));
 sg13g2_buf_1 fanout7026 (.A(net7027),
    .X(net7026));
 sg13g2_buf_8 fanout7027 (.A(net7028),
    .X(net7027));
 sg13g2_buf_8 fanout7028 (.A(net7035),
    .X(net7028));
 sg13g2_buf_8 fanout7029 (.A(net7035),
    .X(net7029));
 sg13g2_buf_1 fanout7030 (.A(net7035),
    .X(net7030));
 sg13g2_buf_8 fanout7031 (.A(net7034),
    .X(net7031));
 sg13g2_buf_1 fanout7032 (.A(net7034),
    .X(net7032));
 sg13g2_buf_8 fanout7033 (.A(net7034),
    .X(net7033));
 sg13g2_buf_8 fanout7034 (.A(net7035),
    .X(net7034));
 sg13g2_buf_8 fanout7035 (.A(_19807_),
    .X(net7035));
 sg13g2_buf_8 fanout7036 (.A(net7037),
    .X(net7036));
 sg13g2_buf_8 fanout7037 (.A(net7038),
    .X(net7037));
 sg13g2_buf_8 fanout7038 (.A(net7044),
    .X(net7038));
 sg13g2_buf_8 fanout7039 (.A(net7040),
    .X(net7039));
 sg13g2_buf_8 fanout7040 (.A(net7044),
    .X(net7040));
 sg13g2_buf_1 fanout7041 (.A(net7044),
    .X(net7041));
 sg13g2_buf_8 fanout7042 (.A(net7043),
    .X(net7042));
 sg13g2_buf_8 fanout7043 (.A(net7044),
    .X(net7043));
 sg13g2_buf_8 fanout7044 (.A(net7077),
    .X(net7044));
 sg13g2_buf_8 fanout7045 (.A(net7047),
    .X(net7045));
 sg13g2_buf_8 fanout7046 (.A(net7047),
    .X(net7046));
 sg13g2_buf_8 fanout7047 (.A(net7077),
    .X(net7047));
 sg13g2_buf_8 fanout7048 (.A(net7052),
    .X(net7048));
 sg13g2_buf_8 fanout7049 (.A(net7052),
    .X(net7049));
 sg13g2_buf_8 fanout7050 (.A(net7051),
    .X(net7050));
 sg13g2_buf_8 fanout7051 (.A(net7052),
    .X(net7051));
 sg13g2_buf_8 fanout7052 (.A(net7077),
    .X(net7052));
 sg13g2_buf_8 fanout7053 (.A(net7063),
    .X(net7053));
 sg13g2_buf_8 fanout7054 (.A(net7063),
    .X(net7054));
 sg13g2_buf_8 fanout7055 (.A(net7057),
    .X(net7055));
 sg13g2_buf_8 fanout7056 (.A(net7057),
    .X(net7056));
 sg13g2_buf_8 fanout7057 (.A(net7063),
    .X(net7057));
 sg13g2_buf_8 fanout7058 (.A(net7062),
    .X(net7058));
 sg13g2_buf_1 fanout7059 (.A(net7062),
    .X(net7059));
 sg13g2_buf_8 fanout7060 (.A(net7062),
    .X(net7060));
 sg13g2_buf_1 fanout7061 (.A(net7062),
    .X(net7061));
 sg13g2_buf_8 fanout7062 (.A(net7063),
    .X(net7062));
 sg13g2_buf_8 fanout7063 (.A(net7064),
    .X(net7063));
 sg13g2_buf_2 fanout7064 (.A(net7077),
    .X(net7064));
 sg13g2_buf_8 fanout7065 (.A(net7066),
    .X(net7065));
 sg13g2_buf_8 fanout7066 (.A(net7067),
    .X(net7066));
 sg13g2_buf_8 fanout7067 (.A(net7076),
    .X(net7067));
 sg13g2_buf_8 fanout7068 (.A(net7071),
    .X(net7068));
 sg13g2_buf_1 fanout7069 (.A(net7071),
    .X(net7069));
 sg13g2_buf_8 fanout7070 (.A(net7071),
    .X(net7070));
 sg13g2_buf_8 fanout7071 (.A(net7076),
    .X(net7071));
 sg13g2_buf_8 fanout7072 (.A(net7075),
    .X(net7072));
 sg13g2_buf_8 fanout7073 (.A(net7075),
    .X(net7073));
 sg13g2_buf_1 fanout7074 (.A(net7075),
    .X(net7074));
 sg13g2_buf_8 fanout7075 (.A(net7076),
    .X(net7075));
 sg13g2_buf_8 fanout7076 (.A(net7077),
    .X(net7076));
 sg13g2_buf_8 fanout7077 (.A(_19807_),
    .X(net7077));
 sg13g2_buf_8 fanout7078 (.A(net7080),
    .X(net7078));
 sg13g2_buf_8 fanout7079 (.A(net7080),
    .X(net7079));
 sg13g2_buf_8 fanout7080 (.A(net7081),
    .X(net7080));
 sg13g2_buf_8 fanout7081 (.A(net7094),
    .X(net7081));
 sg13g2_buf_8 fanout7082 (.A(net7083),
    .X(net7082));
 sg13g2_buf_2 fanout7083 (.A(net7084),
    .X(net7083));
 sg13g2_buf_8 fanout7084 (.A(net7094),
    .X(net7084));
 sg13g2_buf_8 fanout7085 (.A(net7086),
    .X(net7085));
 sg13g2_buf_8 fanout7086 (.A(net7087),
    .X(net7086));
 sg13g2_buf_8 fanout7087 (.A(net7094),
    .X(net7087));
 sg13g2_buf_8 fanout7088 (.A(net7090),
    .X(net7088));
 sg13g2_buf_8 fanout7089 (.A(net7090),
    .X(net7089));
 sg13g2_buf_8 fanout7090 (.A(net7094),
    .X(net7090));
 sg13g2_buf_8 fanout7091 (.A(net7093),
    .X(net7091));
 sg13g2_buf_2 fanout7092 (.A(net7094),
    .X(net7092));
 sg13g2_buf_8 fanout7093 (.A(net7094),
    .X(net7093));
 sg13g2_buf_8 fanout7094 (.A(net7113),
    .X(net7094));
 sg13g2_buf_8 fanout7095 (.A(net7098),
    .X(net7095));
 sg13g2_buf_8 fanout7096 (.A(net7098),
    .X(net7096));
 sg13g2_buf_2 fanout7097 (.A(net7098),
    .X(net7097));
 sg13g2_buf_2 fanout7098 (.A(net7113),
    .X(net7098));
 sg13g2_buf_8 fanout7099 (.A(net7103),
    .X(net7099));
 sg13g2_buf_8 fanout7100 (.A(net7103),
    .X(net7100));
 sg13g2_buf_8 fanout7101 (.A(net7103),
    .X(net7101));
 sg13g2_buf_2 fanout7102 (.A(net7103),
    .X(net7102));
 sg13g2_buf_8 fanout7103 (.A(net7113),
    .X(net7103));
 sg13g2_buf_8 fanout7104 (.A(net7107),
    .X(net7104));
 sg13g2_buf_8 fanout7105 (.A(net7107),
    .X(net7105));
 sg13g2_buf_2 fanout7106 (.A(net7107),
    .X(net7106));
 sg13g2_buf_8 fanout7107 (.A(net7112),
    .X(net7107));
 sg13g2_buf_8 fanout7108 (.A(net7112),
    .X(net7108));
 sg13g2_buf_1 fanout7109 (.A(net7112),
    .X(net7109));
 sg13g2_buf_8 fanout7110 (.A(net7111),
    .X(net7110));
 sg13g2_buf_8 fanout7111 (.A(net7112),
    .X(net7111));
 sg13g2_buf_8 fanout7112 (.A(net7113),
    .X(net7112));
 sg13g2_buf_8 fanout7113 (.A(_19806_),
    .X(net7113));
 sg13g2_buf_8 fanout7114 (.A(net7120),
    .X(net7114));
 sg13g2_buf_2 fanout7115 (.A(net7120),
    .X(net7115));
 sg13g2_buf_8 fanout7116 (.A(net7117),
    .X(net7116));
 sg13g2_buf_8 fanout7117 (.A(net7120),
    .X(net7117));
 sg13g2_buf_8 fanout7118 (.A(net7120),
    .X(net7118));
 sg13g2_buf_8 fanout7119 (.A(net7120),
    .X(net7119));
 sg13g2_buf_8 fanout7120 (.A(net7148),
    .X(net7120));
 sg13g2_buf_8 fanout7121 (.A(net7123),
    .X(net7121));
 sg13g2_buf_1 fanout7122 (.A(net7123),
    .X(net7122));
 sg13g2_buf_8 fanout7123 (.A(net7124),
    .X(net7123));
 sg13g2_buf_8 fanout7124 (.A(net7148),
    .X(net7124));
 sg13g2_buf_8 fanout7125 (.A(net7127),
    .X(net7125));
 sg13g2_buf_8 fanout7126 (.A(net7127),
    .X(net7126));
 sg13g2_buf_8 fanout7127 (.A(net7128),
    .X(net7127));
 sg13g2_buf_8 fanout7128 (.A(net7148),
    .X(net7128));
 sg13g2_buf_8 fanout7129 (.A(net7130),
    .X(net7129));
 sg13g2_buf_8 fanout7130 (.A(net7147),
    .X(net7130));
 sg13g2_buf_8 fanout7131 (.A(net7133),
    .X(net7131));
 sg13g2_buf_1 fanout7132 (.A(net7133),
    .X(net7132));
 sg13g2_buf_8 fanout7133 (.A(net7147),
    .X(net7133));
 sg13g2_buf_8 fanout7134 (.A(net7136),
    .X(net7134));
 sg13g2_buf_8 fanout7135 (.A(net7136),
    .X(net7135));
 sg13g2_buf_8 fanout7136 (.A(net7137),
    .X(net7136));
 sg13g2_buf_8 fanout7137 (.A(net7147),
    .X(net7137));
 sg13g2_buf_8 fanout7138 (.A(net7139),
    .X(net7138));
 sg13g2_buf_8 fanout7139 (.A(net7140),
    .X(net7139));
 sg13g2_buf_8 fanout7140 (.A(net7147),
    .X(net7140));
 sg13g2_buf_8 fanout7141 (.A(net7147),
    .X(net7141));
 sg13g2_buf_8 fanout7142 (.A(net7146),
    .X(net7142));
 sg13g2_buf_8 fanout7143 (.A(net7144),
    .X(net7143));
 sg13g2_buf_8 fanout7144 (.A(net7145),
    .X(net7144));
 sg13g2_buf_8 fanout7145 (.A(net7146),
    .X(net7145));
 sg13g2_buf_8 fanout7146 (.A(net7147),
    .X(net7146));
 sg13g2_buf_8 fanout7147 (.A(net7148),
    .X(net7147));
 sg13g2_buf_8 fanout7148 (.A(_19806_),
    .X(net7148));
 sg13g2_buf_8 fanout7149 (.A(net7150),
    .X(net7149));
 sg13g2_buf_1 fanout7150 (.A(net7162),
    .X(net7150));
 sg13g2_buf_8 fanout7151 (.A(net7153),
    .X(net7151));
 sg13g2_buf_1 fanout7152 (.A(net7153),
    .X(net7152));
 sg13g2_buf_2 fanout7153 (.A(net7162),
    .X(net7153));
 sg13g2_buf_8 fanout7154 (.A(net7155),
    .X(net7154));
 sg13g2_buf_2 fanout7155 (.A(net7156),
    .X(net7155));
 sg13g2_buf_8 fanout7156 (.A(net7157),
    .X(net7156));
 sg13g2_buf_1 fanout7157 (.A(net7162),
    .X(net7157));
 sg13g2_buf_8 fanout7158 (.A(net7159),
    .X(net7158));
 sg13g2_buf_8 fanout7159 (.A(net7160),
    .X(net7159));
 sg13g2_buf_8 fanout7160 (.A(net7161),
    .X(net7160));
 sg13g2_buf_8 fanout7161 (.A(net7162),
    .X(net7161));
 sg13g2_buf_8 fanout7162 (.A(_18944_),
    .X(net7162));
 sg13g2_buf_8 fanout7163 (.A(net7164),
    .X(net7163));
 sg13g2_buf_8 fanout7164 (.A(net7176),
    .X(net7164));
 sg13g2_buf_8 fanout7165 (.A(net7168),
    .X(net7165));
 sg13g2_buf_8 fanout7166 (.A(net7168),
    .X(net7166));
 sg13g2_buf_8 fanout7167 (.A(net7168),
    .X(net7167));
 sg13g2_buf_8 fanout7168 (.A(net7176),
    .X(net7168));
 sg13g2_buf_8 fanout7169 (.A(net7170),
    .X(net7169));
 sg13g2_buf_8 fanout7170 (.A(net7171),
    .X(net7170));
 sg13g2_buf_8 fanout7171 (.A(net7175),
    .X(net7171));
 sg13g2_buf_8 fanout7172 (.A(net7175),
    .X(net7172));
 sg13g2_buf_8 fanout7173 (.A(net7175),
    .X(net7173));
 sg13g2_buf_8 fanout7174 (.A(net7175),
    .X(net7174));
 sg13g2_buf_8 fanout7175 (.A(net7176),
    .X(net7175));
 sg13g2_buf_8 fanout7176 (.A(_18254_),
    .X(net7176));
 sg13g2_buf_8 fanout7177 (.A(net7178),
    .X(net7177));
 sg13g2_buf_8 fanout7178 (.A(net7180),
    .X(net7178));
 sg13g2_buf_8 fanout7179 (.A(net7180),
    .X(net7179));
 sg13g2_buf_8 fanout7180 (.A(net7195),
    .X(net7180));
 sg13g2_buf_8 fanout7181 (.A(net7182),
    .X(net7181));
 sg13g2_buf_8 fanout7182 (.A(net7183),
    .X(net7182));
 sg13g2_buf_2 fanout7183 (.A(net7195),
    .X(net7183));
 sg13g2_buf_8 fanout7184 (.A(net7185),
    .X(net7184));
 sg13g2_buf_8 fanout7185 (.A(net7194),
    .X(net7185));
 sg13g2_buf_8 fanout7186 (.A(net7194),
    .X(net7186));
 sg13g2_buf_8 fanout7187 (.A(net7188),
    .X(net7187));
 sg13g2_buf_1 fanout7188 (.A(net7193),
    .X(net7188));
 sg13g2_buf_8 fanout7189 (.A(net7190),
    .X(net7189));
 sg13g2_buf_8 fanout7190 (.A(net7191),
    .X(net7190));
 sg13g2_buf_8 fanout7191 (.A(net7193),
    .X(net7191));
 sg13g2_buf_8 fanout7192 (.A(net7193),
    .X(net7192));
 sg13g2_buf_8 fanout7193 (.A(net7194),
    .X(net7193));
 sg13g2_buf_8 fanout7194 (.A(net7195),
    .X(net7194));
 sg13g2_buf_8 fanout7195 (.A(_18099_),
    .X(net7195));
 sg13g2_buf_8 fanout7196 (.A(net7210),
    .X(net7196));
 sg13g2_buf_8 fanout7197 (.A(net7210),
    .X(net7197));
 sg13g2_buf_8 fanout7198 (.A(net7199),
    .X(net7198));
 sg13g2_buf_8 fanout7199 (.A(net7202),
    .X(net7199));
 sg13g2_buf_8 fanout7200 (.A(net7201),
    .X(net7200));
 sg13g2_buf_8 fanout7201 (.A(net7202),
    .X(net7201));
 sg13g2_buf_8 fanout7202 (.A(net7210),
    .X(net7202));
 sg13g2_buf_8 fanout7203 (.A(net7204),
    .X(net7203));
 sg13g2_buf_8 fanout7204 (.A(net7209),
    .X(net7204));
 sg13g2_buf_8 fanout7205 (.A(net7206),
    .X(net7205));
 sg13g2_buf_8 fanout7206 (.A(net7209),
    .X(net7206));
 sg13g2_buf_8 fanout7207 (.A(net7208),
    .X(net7207));
 sg13g2_buf_8 fanout7208 (.A(net7209),
    .X(net7208));
 sg13g2_buf_8 fanout7209 (.A(net7210),
    .X(net7209));
 sg13g2_buf_8 fanout7210 (.A(_18099_),
    .X(net7210));
 sg13g2_buf_8 fanout7211 (.A(net7212),
    .X(net7211));
 sg13g2_buf_8 fanout7212 (.A(net7213),
    .X(net7212));
 sg13g2_buf_8 fanout7213 (.A(net7245),
    .X(net7213));
 sg13g2_buf_8 fanout7214 (.A(net7215),
    .X(net7214));
 sg13g2_buf_8 fanout7215 (.A(net7218),
    .X(net7215));
 sg13g2_buf_8 fanout7216 (.A(net7218),
    .X(net7216));
 sg13g2_buf_1 fanout7217 (.A(net7218),
    .X(net7217));
 sg13g2_buf_8 fanout7218 (.A(net7245),
    .X(net7218));
 sg13g2_buf_8 fanout7219 (.A(net7226),
    .X(net7219));
 sg13g2_buf_8 fanout7220 (.A(net7226),
    .X(net7220));
 sg13g2_buf_8 fanout7221 (.A(net7226),
    .X(net7221));
 sg13g2_buf_2 fanout7222 (.A(net7226),
    .X(net7222));
 sg13g2_buf_8 fanout7223 (.A(net7225),
    .X(net7223));
 sg13g2_buf_1 fanout7224 (.A(net7225),
    .X(net7224));
 sg13g2_buf_8 fanout7225 (.A(net7226),
    .X(net7225));
 sg13g2_buf_8 fanout7226 (.A(net7245),
    .X(net7226));
 sg13g2_buf_8 fanout7227 (.A(net7229),
    .X(net7227));
 sg13g2_buf_2 fanout7228 (.A(net7229),
    .X(net7228));
 sg13g2_buf_8 fanout7229 (.A(net7235),
    .X(net7229));
 sg13g2_buf_8 fanout7230 (.A(net7235),
    .X(net7230));
 sg13g2_buf_8 fanout7231 (.A(net7234),
    .X(net7231));
 sg13g2_buf_8 fanout7232 (.A(net7234),
    .X(net7232));
 sg13g2_buf_1 fanout7233 (.A(net7234),
    .X(net7233));
 sg13g2_buf_8 fanout7234 (.A(net7235),
    .X(net7234));
 sg13g2_buf_8 fanout7235 (.A(net7245),
    .X(net7235));
 sg13g2_buf_8 fanout7236 (.A(net7237),
    .X(net7236));
 sg13g2_buf_8 fanout7237 (.A(net7244),
    .X(net7237));
 sg13g2_buf_8 fanout7238 (.A(net7239),
    .X(net7238));
 sg13g2_buf_8 fanout7239 (.A(net7244),
    .X(net7239));
 sg13g2_buf_8 fanout7240 (.A(net7243),
    .X(net7240));
 sg13g2_buf_8 fanout7241 (.A(net7243),
    .X(net7241));
 sg13g2_buf_2 fanout7242 (.A(net7243),
    .X(net7242));
 sg13g2_buf_8 fanout7243 (.A(net7244),
    .X(net7243));
 sg13g2_buf_8 fanout7244 (.A(net7245),
    .X(net7244));
 sg13g2_buf_8 fanout7245 (.A(_18099_),
    .X(net7245));
 sg13g2_buf_8 fanout7246 (.A(net3757),
    .X(net7246));
 sg13g2_buf_8 fanout7247 (.A(net3749),
    .X(net7247));
 sg13g2_buf_8 fanout7248 (.A(net7249),
    .X(net7248));
 sg13g2_buf_1 fanout7249 (.A(net3760),
    .X(net7249));
 sg13g2_buf_8 fanout7250 (.A(\u_inv.counter[0] ),
    .X(net7250));
 sg13g2_buf_1 fanout7251 (.A(net3743),
    .X(net7251));
 sg13g2_buf_8 fanout7252 (.A(net7254),
    .X(net7252));
 sg13g2_buf_8 fanout7253 (.A(net7254),
    .X(net7253));
 sg13g2_buf_8 fanout7254 (.A(net7255),
    .X(net7254));
 sg13g2_buf_8 fanout7255 (.A(net7259),
    .X(net7255));
 sg13g2_buf_8 fanout7256 (.A(net7258),
    .X(net7256));
 sg13g2_buf_1 fanout7257 (.A(net7258),
    .X(net7257));
 sg13g2_buf_2 fanout7258 (.A(net7259),
    .X(net7258));
 sg13g2_buf_1 fanout7259 (.A(net7286),
    .X(net7259));
 sg13g2_buf_8 fanout7260 (.A(net7264),
    .X(net7260));
 sg13g2_buf_8 fanout7261 (.A(net7264),
    .X(net7261));
 sg13g2_buf_1 fanout7262 (.A(net7263),
    .X(net7262));
 sg13g2_buf_8 fanout7263 (.A(net7264),
    .X(net7263));
 sg13g2_buf_8 fanout7264 (.A(net7268),
    .X(net7264));
 sg13g2_buf_8 fanout7265 (.A(net7268),
    .X(net7265));
 sg13g2_buf_8 fanout7266 (.A(net7267),
    .X(net7266));
 sg13g2_buf_8 fanout7267 (.A(net7268),
    .X(net7267));
 sg13g2_buf_8 fanout7268 (.A(net7286),
    .X(net7268));
 sg13g2_buf_8 fanout7269 (.A(net7272),
    .X(net7269));
 sg13g2_buf_1 fanout7270 (.A(net7272),
    .X(net7270));
 sg13g2_buf_8 fanout7271 (.A(net7272),
    .X(net7271));
 sg13g2_buf_8 fanout7272 (.A(net7286),
    .X(net7272));
 sg13g2_buf_8 fanout7273 (.A(net7274),
    .X(net7273));
 sg13g2_buf_8 fanout7274 (.A(net7275),
    .X(net7274));
 sg13g2_buf_8 fanout7275 (.A(net7286),
    .X(net7275));
 sg13g2_buf_8 fanout7276 (.A(net7277),
    .X(net7276));
 sg13g2_buf_8 fanout7277 (.A(net7278),
    .X(net7277));
 sg13g2_buf_8 fanout7278 (.A(net7279),
    .X(net7278));
 sg13g2_buf_8 fanout7279 (.A(net7285),
    .X(net7279));
 sg13g2_buf_8 fanout7280 (.A(net7281),
    .X(net7280));
 sg13g2_buf_2 fanout7281 (.A(net7282),
    .X(net7281));
 sg13g2_buf_8 fanout7282 (.A(net7285),
    .X(net7282));
 sg13g2_buf_8 fanout7283 (.A(net7285),
    .X(net7283));
 sg13g2_buf_1 fanout7284 (.A(net7285),
    .X(net7284));
 sg13g2_buf_8 fanout7285 (.A(net7286),
    .X(net7285));
 sg13g2_buf_8 fanout7286 (.A(\u_inv.f_reg[256] ),
    .X(net7286));
 sg13g2_buf_8 fanout7287 (.A(\u_inv.d_reg[241] ),
    .X(net7287));
 sg13g2_buf_8 fanout7288 (.A(\u_inv.d_reg[240] ),
    .X(net7288));
 sg13g2_buf_8 fanout7289 (.A(\u_inv.d_reg[130] ),
    .X(net7289));
 sg13g2_buf_8 fanout7290 (.A(\u_inv.d_reg[81] ),
    .X(net7290));
 sg13g2_buf_8 fanout7291 (.A(\u_inv.d_reg[22] ),
    .X(net7291));
 sg13g2_buf_8 fanout7292 (.A(\u_inv.d_reg[10] ),
    .X(net7292));
 sg13g2_buf_8 fanout7293 (.A(\u_inv.d_reg[1] ),
    .X(net7293));
 sg13g2_buf_8 fanout7294 (.A(\u_inv.d_reg[0] ),
    .X(net7294));
 sg13g2_buf_8 fanout7295 (.A(net1191),
    .X(net7295));
 sg13g2_buf_8 fanout7296 (.A(\u_inv.d_next[130] ),
    .X(net7296));
 sg13g2_buf_8 fanout7297 (.A(net1867),
    .X(net7297));
 sg13g2_buf_8 fanout7298 (.A(net1238),
    .X(net7298));
 sg13g2_buf_8 fanout7299 (.A(net2381),
    .X(net7299));
 sg13g2_buf_8 fanout7300 (.A(\u_inv.f_next[19] ),
    .X(net7300));
 sg13g2_buf_8 fanout7301 (.A(net7302),
    .X(net7301));
 sg13g2_buf_1 fanout7302 (.A(net7303),
    .X(net7302));
 sg13g2_buf_8 fanout7303 (.A(net7313),
    .X(net7303));
 sg13g2_buf_8 fanout7304 (.A(net7305),
    .X(net7304));
 sg13g2_buf_8 fanout7305 (.A(net7306),
    .X(net7305));
 sg13g2_buf_8 fanout7306 (.A(net7313),
    .X(net7306));
 sg13g2_buf_8 fanout7307 (.A(net7308),
    .X(net7307));
 sg13g2_buf_8 fanout7308 (.A(net7313),
    .X(net7308));
 sg13g2_buf_8 fanout7309 (.A(net7310),
    .X(net7309));
 sg13g2_buf_8 fanout7310 (.A(net7313),
    .X(net7310));
 sg13g2_buf_8 fanout7311 (.A(net7312),
    .X(net7311));
 sg13g2_buf_8 fanout7312 (.A(net7313),
    .X(net7312));
 sg13g2_buf_8 fanout7313 (.A(net7352),
    .X(net7313));
 sg13g2_buf_8 fanout7314 (.A(net7315),
    .X(net7314));
 sg13g2_buf_8 fanout7315 (.A(net7316),
    .X(net7315));
 sg13g2_buf_8 fanout7316 (.A(net7319),
    .X(net7316));
 sg13g2_buf_8 fanout7317 (.A(net7319),
    .X(net7317));
 sg13g2_buf_8 fanout7318 (.A(net7319),
    .X(net7318));
 sg13g2_buf_8 fanout7319 (.A(net7352),
    .X(net7319));
 sg13g2_buf_8 fanout7320 (.A(net7321),
    .X(net7320));
 sg13g2_buf_8 fanout7321 (.A(net7322),
    .X(net7321));
 sg13g2_buf_8 fanout7322 (.A(net7323),
    .X(net7322));
 sg13g2_buf_8 fanout7323 (.A(net7352),
    .X(net7323));
 sg13g2_buf_8 fanout7324 (.A(net7326),
    .X(net7324));
 sg13g2_buf_8 fanout7325 (.A(net7326),
    .X(net7325));
 sg13g2_buf_8 fanout7326 (.A(net7327),
    .X(net7326));
 sg13g2_buf_1 fanout7327 (.A(net7351),
    .X(net7327));
 sg13g2_buf_8 fanout7328 (.A(net7332),
    .X(net7328));
 sg13g2_buf_1 fanout7329 (.A(net7332),
    .X(net7329));
 sg13g2_buf_8 fanout7330 (.A(net7332),
    .X(net7330));
 sg13g2_buf_1 fanout7331 (.A(net7332),
    .X(net7331));
 sg13g2_buf_8 fanout7332 (.A(net7351),
    .X(net7332));
 sg13g2_buf_8 fanout7333 (.A(net7334),
    .X(net7333));
 sg13g2_buf_8 fanout7334 (.A(net7338),
    .X(net7334));
 sg13g2_buf_8 fanout7335 (.A(net7337),
    .X(net7335));
 sg13g2_buf_1 fanout7336 (.A(net7337),
    .X(net7336));
 sg13g2_buf_8 fanout7337 (.A(net7338),
    .X(net7337));
 sg13g2_buf_8 fanout7338 (.A(net7351),
    .X(net7338));
 sg13g2_buf_8 fanout7339 (.A(net7342),
    .X(net7339));
 sg13g2_buf_1 fanout7340 (.A(net7342),
    .X(net7340));
 sg13g2_buf_8 fanout7341 (.A(net7342),
    .X(net7341));
 sg13g2_buf_8 fanout7342 (.A(net7351),
    .X(net7342));
 sg13g2_buf_8 fanout7343 (.A(net7345),
    .X(net7343));
 sg13g2_buf_8 fanout7344 (.A(net7345),
    .X(net7344));
 sg13g2_buf_8 fanout7345 (.A(net7351),
    .X(net7345));
 sg13g2_buf_8 fanout7346 (.A(net7350),
    .X(net7346));
 sg13g2_buf_1 fanout7347 (.A(net7350),
    .X(net7347));
 sg13g2_buf_8 fanout7348 (.A(net7350),
    .X(net7348));
 sg13g2_buf_1 fanout7349 (.A(net7350),
    .X(net7349));
 sg13g2_buf_8 fanout7350 (.A(net7351),
    .X(net7350));
 sg13g2_buf_8 fanout7351 (.A(net7352),
    .X(net7351));
 sg13g2_buf_8 fanout7352 (.A(\u_inv.f_next[0] ),
    .X(net7352));
 sg13g2_buf_8 fanout7353 (.A(net7354),
    .X(net7353));
 sg13g2_buf_8 fanout7354 (.A(net7362),
    .X(net7354));
 sg13g2_buf_8 fanout7355 (.A(net7356),
    .X(net7355));
 sg13g2_buf_8 fanout7356 (.A(net7362),
    .X(net7356));
 sg13g2_buf_8 fanout7357 (.A(net7359),
    .X(net7357));
 sg13g2_buf_8 fanout7358 (.A(net7359),
    .X(net7358));
 sg13g2_buf_8 fanout7359 (.A(net7362),
    .X(net7359));
 sg13g2_buf_8 fanout7360 (.A(net7362),
    .X(net7360));
 sg13g2_buf_2 fanout7361 (.A(net7362),
    .X(net7361));
 sg13g2_buf_8 fanout7362 (.A(net7377),
    .X(net7362));
 sg13g2_buf_8 fanout7363 (.A(net7377),
    .X(net7363));
 sg13g2_buf_1 fanout7364 (.A(net7377),
    .X(net7364));
 sg13g2_buf_8 fanout7365 (.A(net7366),
    .X(net7365));
 sg13g2_buf_8 fanout7366 (.A(net7368),
    .X(net7366));
 sg13g2_buf_8 fanout7367 (.A(net7368),
    .X(net7367));
 sg13g2_buf_8 fanout7368 (.A(net7377),
    .X(net7368));
 sg13g2_buf_8 fanout7369 (.A(net7370),
    .X(net7369));
 sg13g2_buf_8 fanout7370 (.A(net7372),
    .X(net7370));
 sg13g2_buf_8 fanout7371 (.A(net7372),
    .X(net7371));
 sg13g2_buf_8 fanout7372 (.A(net7377),
    .X(net7372));
 sg13g2_buf_8 fanout7373 (.A(net7374),
    .X(net7373));
 sg13g2_buf_8 fanout7374 (.A(net7376),
    .X(net7374));
 sg13g2_buf_8 fanout7375 (.A(net7376),
    .X(net7375));
 sg13g2_buf_8 fanout7376 (.A(net7377),
    .X(net7376));
 sg13g2_buf_8 fanout7377 (.A(\u_inv.f_next[0] ),
    .X(net7377));
 sg13g2_buf_8 fanout7378 (.A(net7383),
    .X(net7378));
 sg13g2_buf_1 fanout7379 (.A(net7383),
    .X(net7379));
 sg13g2_buf_8 fanout7380 (.A(net7383),
    .X(net7380));
 sg13g2_buf_8 fanout7381 (.A(net7382),
    .X(net7381));
 sg13g2_buf_8 fanout7382 (.A(net7383),
    .X(net7382));
 sg13g2_buf_8 fanout7383 (.A(net7411),
    .X(net7383));
 sg13g2_buf_8 fanout7384 (.A(net7389),
    .X(net7384));
 sg13g2_buf_1 fanout7385 (.A(net7389),
    .X(net7385));
 sg13g2_buf_8 fanout7386 (.A(net7389),
    .X(net7386));
 sg13g2_buf_8 fanout7387 (.A(net7389),
    .X(net7387));
 sg13g2_buf_8 fanout7388 (.A(net7389),
    .X(net7388));
 sg13g2_buf_8 fanout7389 (.A(net7411),
    .X(net7389));
 sg13g2_buf_8 fanout7390 (.A(net7391),
    .X(net7390));
 sg13g2_buf_8 fanout7391 (.A(net7394),
    .X(net7391));
 sg13g2_buf_8 fanout7392 (.A(net7394),
    .X(net7392));
 sg13g2_buf_8 fanout7393 (.A(net7394),
    .X(net7393));
 sg13g2_buf_8 fanout7394 (.A(net7411),
    .X(net7394));
 sg13g2_buf_8 fanout7395 (.A(net7396),
    .X(net7395));
 sg13g2_buf_1 fanout7396 (.A(net7410),
    .X(net7396));
 sg13g2_buf_8 fanout7397 (.A(net7401),
    .X(net7397));
 sg13g2_buf_8 fanout7398 (.A(net7401),
    .X(net7398));
 sg13g2_buf_1 fanout7399 (.A(net7401),
    .X(net7399));
 sg13g2_buf_8 fanout7400 (.A(net7401),
    .X(net7400));
 sg13g2_buf_8 fanout7401 (.A(net7410),
    .X(net7401));
 sg13g2_buf_8 fanout7402 (.A(net7403),
    .X(net7402));
 sg13g2_buf_8 fanout7403 (.A(net7404),
    .X(net7403));
 sg13g2_buf_2 fanout7404 (.A(net7410),
    .X(net7404));
 sg13g2_buf_8 fanout7405 (.A(net7410),
    .X(net7405));
 sg13g2_buf_1 fanout7406 (.A(net7410),
    .X(net7406));
 sg13g2_buf_8 fanout7407 (.A(net7409),
    .X(net7407));
 sg13g2_buf_1 fanout7408 (.A(net7409),
    .X(net7408));
 sg13g2_buf_8 fanout7409 (.A(net7410),
    .X(net7409));
 sg13g2_buf_8 fanout7410 (.A(net7411),
    .X(net7410));
 sg13g2_buf_8 fanout7411 (.A(\u_inv.f_next[0] ),
    .X(net7411));
 sg13g2_buf_8 fanout7412 (.A(\state[1] ),
    .X(net7412));
 sg13g2_buf_8 fanout7413 (.A(net3747),
    .X(net7413));
 sg13g2_buf_8 fanout7414 (.A(net7415),
    .X(net7414));
 sg13g2_buf_8 fanout7415 (.A(net7416),
    .X(net7415));
 sg13g2_buf_8 fanout7416 (.A(net7429),
    .X(net7416));
 sg13g2_buf_8 fanout7417 (.A(net7420),
    .X(net7417));
 sg13g2_buf_8 fanout7418 (.A(net7420),
    .X(net7418));
 sg13g2_buf_8 fanout7419 (.A(net7420),
    .X(net7419));
 sg13g2_buf_8 fanout7420 (.A(net7429),
    .X(net7420));
 sg13g2_buf_8 fanout7421 (.A(net7424),
    .X(net7421));
 sg13g2_buf_8 fanout7422 (.A(net7424),
    .X(net7422));
 sg13g2_buf_2 fanout7423 (.A(net7424),
    .X(net7423));
 sg13g2_buf_8 fanout7424 (.A(net7429),
    .X(net7424));
 sg13g2_buf_8 fanout7425 (.A(net7428),
    .X(net7425));
 sg13g2_buf_8 fanout7426 (.A(net7428),
    .X(net7426));
 sg13g2_buf_8 fanout7427 (.A(net7428),
    .X(net7427));
 sg13g2_buf_8 fanout7428 (.A(net7429),
    .X(net7428));
 sg13g2_buf_8 fanout7429 (.A(net7455),
    .X(net7429));
 sg13g2_buf_8 fanout7430 (.A(net7433),
    .X(net7430));
 sg13g2_buf_2 fanout7431 (.A(net7433),
    .X(net7431));
 sg13g2_buf_8 fanout7432 (.A(net7433),
    .X(net7432));
 sg13g2_buf_8 fanout7433 (.A(net7434),
    .X(net7433));
 sg13g2_buf_8 fanout7434 (.A(net7440),
    .X(net7434));
 sg13g2_buf_8 fanout7435 (.A(net7440),
    .X(net7435));
 sg13g2_buf_1 fanout7436 (.A(net7440),
    .X(net7436));
 sg13g2_buf_8 fanout7437 (.A(net7438),
    .X(net7437));
 sg13g2_buf_8 fanout7438 (.A(net7439),
    .X(net7438));
 sg13g2_buf_8 fanout7439 (.A(net7440),
    .X(net7439));
 sg13g2_buf_8 fanout7440 (.A(net7455),
    .X(net7440));
 sg13g2_buf_8 fanout7441 (.A(net7442),
    .X(net7441));
 sg13g2_buf_8 fanout7442 (.A(net7447),
    .X(net7442));
 sg13g2_buf_8 fanout7443 (.A(net7447),
    .X(net7443));
 sg13g2_buf_2 fanout7444 (.A(net7447),
    .X(net7444));
 sg13g2_buf_8 fanout7445 (.A(net7446),
    .X(net7445));
 sg13g2_buf_8 fanout7446 (.A(net7447),
    .X(net7446));
 sg13g2_buf_8 fanout7447 (.A(net7455),
    .X(net7447));
 sg13g2_buf_8 fanout7448 (.A(net7452),
    .X(net7448));
 sg13g2_buf_8 fanout7449 (.A(net7452),
    .X(net7449));
 sg13g2_buf_8 fanout7450 (.A(net7452),
    .X(net7450));
 sg13g2_buf_8 fanout7451 (.A(net7452),
    .X(net7451));
 sg13g2_buf_8 fanout7452 (.A(net7454),
    .X(net7452));
 sg13g2_buf_8 fanout7453 (.A(net7454),
    .X(net7453));
 sg13g2_buf_8 fanout7454 (.A(net7455),
    .X(net7454));
 sg13g2_buf_8 fanout7455 (.A(net7569),
    .X(net7455));
 sg13g2_buf_8 fanout7456 (.A(net7457),
    .X(net7456));
 sg13g2_buf_2 fanout7457 (.A(net7458),
    .X(net7457));
 sg13g2_buf_8 fanout7458 (.A(net7462),
    .X(net7458));
 sg13g2_buf_8 fanout7459 (.A(net7460),
    .X(net7459));
 sg13g2_buf_8 fanout7460 (.A(net7462),
    .X(net7460));
 sg13g2_buf_8 fanout7461 (.A(net7462),
    .X(net7461));
 sg13g2_buf_8 fanout7462 (.A(net7470),
    .X(net7462));
 sg13g2_buf_8 fanout7463 (.A(net7469),
    .X(net7463));
 sg13g2_buf_8 fanout7464 (.A(net7469),
    .X(net7464));
 sg13g2_buf_8 fanout7465 (.A(net7466),
    .X(net7465));
 sg13g2_buf_8 fanout7466 (.A(net7467),
    .X(net7466));
 sg13g2_buf_8 fanout7467 (.A(net7468),
    .X(net7467));
 sg13g2_buf_8 fanout7468 (.A(net7469),
    .X(net7468));
 sg13g2_buf_8 fanout7469 (.A(net7470),
    .X(net7469));
 sg13g2_buf_8 fanout7470 (.A(net7569),
    .X(net7470));
 sg13g2_buf_8 fanout7471 (.A(net7477),
    .X(net7471));
 sg13g2_buf_8 fanout7472 (.A(net7477),
    .X(net7472));
 sg13g2_buf_8 fanout7473 (.A(net7477),
    .X(net7473));
 sg13g2_buf_8 fanout7474 (.A(net7476),
    .X(net7474));
 sg13g2_buf_8 fanout7475 (.A(net7476),
    .X(net7475));
 sg13g2_buf_8 fanout7476 (.A(net7477),
    .X(net7476));
 sg13g2_buf_8 fanout7477 (.A(net7494),
    .X(net7477));
 sg13g2_buf_8 fanout7478 (.A(net7479),
    .X(net7478));
 sg13g2_buf_8 fanout7479 (.A(net7482),
    .X(net7479));
 sg13g2_buf_8 fanout7480 (.A(net7482),
    .X(net7480));
 sg13g2_buf_8 fanout7481 (.A(net7482),
    .X(net7481));
 sg13g2_buf_8 fanout7482 (.A(net7494),
    .X(net7482));
 sg13g2_buf_8 fanout7483 (.A(net7484),
    .X(net7483));
 sg13g2_buf_8 fanout7484 (.A(net7485),
    .X(net7484));
 sg13g2_buf_8 fanout7485 (.A(net7492),
    .X(net7485));
 sg13g2_buf_8 fanout7486 (.A(net7492),
    .X(net7486));
 sg13g2_buf_8 fanout7487 (.A(net7492),
    .X(net7487));
 sg13g2_buf_8 fanout7488 (.A(net7489),
    .X(net7488));
 sg13g2_buf_8 fanout7489 (.A(net7491),
    .X(net7489));
 sg13g2_buf_8 fanout7490 (.A(net7491),
    .X(net7490));
 sg13g2_buf_8 fanout7491 (.A(net7492),
    .X(net7491));
 sg13g2_buf_8 fanout7492 (.A(net7494),
    .X(net7492));
 sg13g2_buf_8 fanout7493 (.A(net7494),
    .X(net7493));
 sg13g2_buf_8 fanout7494 (.A(net7569),
    .X(net7494));
 sg13g2_buf_8 fanout7495 (.A(net7497),
    .X(net7495));
 sg13g2_buf_8 fanout7496 (.A(net7497),
    .X(net7496));
 sg13g2_buf_8 fanout7497 (.A(net7501),
    .X(net7497));
 sg13g2_buf_8 fanout7498 (.A(net7500),
    .X(net7498));
 sg13g2_buf_8 fanout7499 (.A(net7500),
    .X(net7499));
 sg13g2_buf_8 fanout7500 (.A(net7501),
    .X(net7500));
 sg13g2_buf_8 fanout7501 (.A(net7568),
    .X(net7501));
 sg13g2_buf_8 fanout7502 (.A(net7503),
    .X(net7502));
 sg13g2_buf_8 fanout7503 (.A(net7511),
    .X(net7503));
 sg13g2_buf_8 fanout7504 (.A(net7506),
    .X(net7504));
 sg13g2_buf_8 fanout7505 (.A(net7506),
    .X(net7505));
 sg13g2_buf_8 fanout7506 (.A(net7511),
    .X(net7506));
 sg13g2_buf_8 fanout7507 (.A(net7509),
    .X(net7507));
 sg13g2_buf_8 fanout7508 (.A(net7509),
    .X(net7508));
 sg13g2_buf_8 fanout7509 (.A(net7510),
    .X(net7509));
 sg13g2_buf_8 fanout7510 (.A(net7511),
    .X(net7510));
 sg13g2_buf_8 fanout7511 (.A(net7568),
    .X(net7511));
 sg13g2_buf_8 fanout7512 (.A(net7515),
    .X(net7512));
 sg13g2_buf_8 fanout7513 (.A(net7514),
    .X(net7513));
 sg13g2_buf_8 fanout7514 (.A(net7515),
    .X(net7514));
 sg13g2_buf_8 fanout7515 (.A(net7516),
    .X(net7515));
 sg13g2_buf_8 fanout7516 (.A(net7525),
    .X(net7516));
 sg13g2_buf_8 fanout7517 (.A(net7518),
    .X(net7517));
 sg13g2_buf_8 fanout7518 (.A(net7519),
    .X(net7518));
 sg13g2_buf_8 fanout7519 (.A(net7520),
    .X(net7519));
 sg13g2_buf_8 fanout7520 (.A(net7525),
    .X(net7520));
 sg13g2_buf_8 fanout7521 (.A(net7522),
    .X(net7521));
 sg13g2_buf_8 fanout7522 (.A(net7525),
    .X(net7522));
 sg13g2_buf_8 fanout7523 (.A(net7524),
    .X(net7523));
 sg13g2_buf_8 fanout7524 (.A(net7525),
    .X(net7524));
 sg13g2_buf_8 fanout7525 (.A(net7568),
    .X(net7525));
 sg13g2_buf_8 fanout7526 (.A(net7528),
    .X(net7526));
 sg13g2_buf_8 fanout7527 (.A(net7528),
    .X(net7527));
 sg13g2_buf_8 fanout7528 (.A(net7549),
    .X(net7528));
 sg13g2_buf_8 fanout7529 (.A(net7530),
    .X(net7529));
 sg13g2_buf_8 fanout7530 (.A(net7549),
    .X(net7530));
 sg13g2_buf_8 fanout7531 (.A(net7532),
    .X(net7531));
 sg13g2_buf_8 fanout7532 (.A(net7533),
    .X(net7532));
 sg13g2_buf_8 fanout7533 (.A(net7537),
    .X(net7533));
 sg13g2_buf_8 fanout7534 (.A(net7535),
    .X(net7534));
 sg13g2_buf_8 fanout7535 (.A(net7537),
    .X(net7535));
 sg13g2_buf_8 fanout7536 (.A(net7537),
    .X(net7536));
 sg13g2_buf_8 fanout7537 (.A(net7549),
    .X(net7537));
 sg13g2_buf_8 fanout7538 (.A(net7541),
    .X(net7538));
 sg13g2_buf_2 fanout7539 (.A(net7544),
    .X(net7539));
 sg13g2_buf_8 fanout7540 (.A(net7541),
    .X(net7540));
 sg13g2_buf_8 fanout7541 (.A(net7544),
    .X(net7541));
 sg13g2_buf_8 fanout7542 (.A(net7544),
    .X(net7542));
 sg13g2_buf_2 fanout7543 (.A(net7544),
    .X(net7543));
 sg13g2_buf_2 fanout7544 (.A(net7549),
    .X(net7544));
 sg13g2_buf_8 fanout7545 (.A(net7547),
    .X(net7545));
 sg13g2_buf_8 fanout7546 (.A(net7547),
    .X(net7546));
 sg13g2_buf_8 fanout7547 (.A(net7548),
    .X(net7547));
 sg13g2_buf_8 fanout7548 (.A(net7549),
    .X(net7548));
 sg13g2_buf_8 fanout7549 (.A(net7568),
    .X(net7549));
 sg13g2_buf_8 fanout7550 (.A(net7557),
    .X(net7550));
 sg13g2_buf_8 fanout7551 (.A(net7552),
    .X(net7551));
 sg13g2_buf_8 fanout7552 (.A(net7557),
    .X(net7552));
 sg13g2_buf_8 fanout7553 (.A(net7557),
    .X(net7553));
 sg13g2_buf_8 fanout7554 (.A(net7557),
    .X(net7554));
 sg13g2_buf_8 fanout7555 (.A(net7556),
    .X(net7555));
 sg13g2_buf_8 fanout7556 (.A(net7557),
    .X(net7556));
 sg13g2_buf_8 fanout7557 (.A(net7567),
    .X(net7557));
 sg13g2_buf_8 fanout7558 (.A(net7560),
    .X(net7558));
 sg13g2_buf_8 fanout7559 (.A(net7560),
    .X(net7559));
 sg13g2_buf_8 fanout7560 (.A(net7562),
    .X(net7560));
 sg13g2_buf_8 fanout7561 (.A(net7562),
    .X(net7561));
 sg13g2_buf_8 fanout7562 (.A(net7567),
    .X(net7562));
 sg13g2_buf_8 fanout7563 (.A(net7565),
    .X(net7563));
 sg13g2_buf_8 fanout7564 (.A(net7565),
    .X(net7564));
 sg13g2_buf_8 fanout7565 (.A(net7566),
    .X(net7565));
 sg13g2_buf_8 fanout7566 (.A(net7567),
    .X(net7566));
 sg13g2_buf_8 fanout7567 (.A(net7568),
    .X(net7567));
 sg13g2_buf_8 fanout7568 (.A(net7569),
    .X(net7568));
 sg13g2_buf_8 fanout7569 (.A(rst_n),
    .X(net7569));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[2]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[3]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[4]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[5]),
    .X(net13));
 sg13g2_tielo tt_um_corey_14 (.L_LO(net14));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_8 clkbuf_leaf_113_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_8 clkbuf_leaf_123_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_8 clkbuf_leaf_124_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_8 clkbuf_leaf_125_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_8 clkbuf_leaf_126_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_8 clkbuf_leaf_127_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_8 clkbuf_leaf_128_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_8 clkbuf_leaf_129_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_8 clkbuf_leaf_130_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_8 clkbuf_leaf_131_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_8 clkbuf_leaf_132_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_8 clkbuf_leaf_133_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_8 clkbuf_leaf_134_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_8 clkbuf_leaf_135_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_8 clkbuf_leaf_136_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_8 clkbuf_leaf_137_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_8 clkbuf_leaf_138_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_8 clkbuf_leaf_139_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_8 clkbuf_leaf_140_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_8 clkbuf_leaf_141_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_8 clkbuf_leaf_142_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_8 clkbuf_leaf_143_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_8 clkbuf_leaf_144_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_8 clkbuf_leaf_145_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_8 clkbuf_leaf_146_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_8 clkbuf_leaf_147_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_8 clkbuf_leaf_148_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_8 clkbuf_leaf_149_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_8 clkbuf_leaf_150_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_8 clkbuf_leaf_151_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_8 clkbuf_leaf_152_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_8 clkbuf_leaf_153_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_8 clkbuf_leaf_154_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_8 clkbuf_leaf_155_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_8 clkbuf_leaf_156_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_8 clkbuf_leaf_157_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_8 clkbuf_leaf_158_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_8 clkbuf_leaf_159_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_8 clkbuf_leaf_160_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_8 clkbuf_leaf_161_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_8 clkbuf_leaf_162_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_8 clkbuf_leaf_163_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_8 clkbuf_leaf_164_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_8 clkbuf_leaf_165_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_8 clkbuf_leaf_166_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_8 clkbuf_leaf_167_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_8 clkbuf_leaf_168_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_8 clkbuf_leaf_169_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_8 clkbuf_leaf_170_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_8 clkbuf_leaf_171_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_8 clkbuf_leaf_172_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_8 clkbuf_leaf_173_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_8 clkbuf_leaf_174_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_8 clkbuf_leaf_175_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_8 clkbuf_leaf_176_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_8 clkbuf_leaf_177_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_8 clkbuf_leaf_178_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_8 clkbuf_leaf_179_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_8 clkbuf_leaf_180_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_8 clkbuf_leaf_181_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_8 clkbuf_leaf_182_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_8 clkbuf_leaf_183_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_8 clkbuf_leaf_184_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_8 clkbuf_leaf_185_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_8 clkbuf_leaf_186_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_8 clkbuf_leaf_187_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_8 clkbuf_leaf_188_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_8 clkbuf_leaf_189_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_8 clkbuf_leaf_190_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_8 clkbuf_leaf_191_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_8 clkbuf_leaf_192_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_8 clkbuf_leaf_193_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_8 clkbuf_leaf_194_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_8 clkbuf_leaf_195_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_8 clkbuf_leaf_196_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_8 clkbuf_leaf_197_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_8 clkbuf_leaf_198_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_8 clkbuf_leaf_199_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_8 clkbuf_leaf_200_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_8 clkbuf_leaf_201_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_8 clkbuf_leaf_202_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_8 clkbuf_leaf_203_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_8 clkbuf_leaf_204_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_8 clkbuf_leaf_205_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_8 clkbuf_leaf_206_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_8 clkbuf_leaf_207_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_8 clkbuf_leaf_208_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_8 clkbuf_leaf_209_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_8 clkbuf_leaf_210_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_8 clkbuf_leaf_211_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_8 clkbuf_leaf_212_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_8 clkbuf_leaf_213_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_8 clkbuf_leaf_214_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_8 clkbuf_leaf_215_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_8 clkbuf_leaf_216_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_8 clkbuf_leaf_217_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_8 clkbuf_leaf_218_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_8 clkbuf_leaf_219_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_8 clkbuf_leaf_220_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_8 clkbuf_leaf_221_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_8 clkbuf_leaf_222_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_8 clkbuf_leaf_223_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_8 clkbuf_leaf_224_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_8 clkbuf_leaf_225_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_8 clkbuf_leaf_226_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_8 clkbuf_leaf_227_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_8 clkbuf_leaf_228_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_8 clkbuf_leaf_229_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_8 clkbuf_leaf_230_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_8 clkbuf_leaf_231_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_8 clkbuf_leaf_232_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_8 clkbuf_leaf_233_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_8 clkbuf_leaf_234_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_8 clkbuf_leaf_235_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_8 clkbuf_leaf_236_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_8 clkbuf_leaf_237_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_8 clkbuf_leaf_238_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_8 clkbuf_leaf_239_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_8 clkbuf_leaf_240_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_8 clkbuf_leaf_241_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_8 clkbuf_leaf_242_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_8 clkbuf_leaf_243_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_8 clkbuf_leaf_244_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .X(clknet_2_0_0_clk));
 sg13g2_buf_8 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .X(clknet_2_1_0_clk));
 sg13g2_buf_8 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .X(clknet_2_2_0_clk));
 sg13g2_buf_8 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .X(clknet_2_3_0_clk));
 sg13g2_buf_8 clkbuf_5_0_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_0_0_clk));
 sg13g2_buf_8 clkbuf_5_1_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_1_0_clk));
 sg13g2_buf_8 clkbuf_5_2_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_2_0_clk));
 sg13g2_buf_8 clkbuf_5_3_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_3_0_clk));
 sg13g2_buf_8 clkbuf_5_4_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_4_0_clk));
 sg13g2_buf_8 clkbuf_5_5_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_5_0_clk));
 sg13g2_buf_8 clkbuf_5_6_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_6_0_clk));
 sg13g2_buf_8 clkbuf_5_7_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_7_0_clk));
 sg13g2_buf_8 clkbuf_5_8_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_8_0_clk));
 sg13g2_buf_8 clkbuf_5_9_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_9_0_clk));
 sg13g2_buf_8 clkbuf_5_10_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_10_0_clk));
 sg13g2_buf_8 clkbuf_5_11_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_11_0_clk));
 sg13g2_buf_8 clkbuf_5_12_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_12_0_clk));
 sg13g2_buf_8 clkbuf_5_13_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_13_0_clk));
 sg13g2_buf_8 clkbuf_5_14_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_14_0_clk));
 sg13g2_buf_8 clkbuf_5_15_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_15_0_clk));
 sg13g2_buf_8 clkbuf_5_16_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_16_0_clk));
 sg13g2_buf_8 clkbuf_5_17_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_17_0_clk));
 sg13g2_buf_8 clkbuf_5_18_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_18_0_clk));
 sg13g2_buf_8 clkbuf_5_19_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_19_0_clk));
 sg13g2_buf_8 clkbuf_5_20_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_20_0_clk));
 sg13g2_buf_8 clkbuf_5_21_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_21_0_clk));
 sg13g2_buf_8 clkbuf_5_22_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_22_0_clk));
 sg13g2_buf_8 clkbuf_5_23_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_23_0_clk));
 sg13g2_buf_8 clkbuf_5_24_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_24_0_clk));
 sg13g2_buf_8 clkbuf_5_25_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_25_0_clk));
 sg13g2_buf_8 clkbuf_5_26_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_26_0_clk));
 sg13g2_buf_8 clkbuf_5_27_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_27_0_clk));
 sg13g2_buf_8 clkbuf_5_28_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_28_0_clk));
 sg13g2_buf_8 clkbuf_5_29_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_29_0_clk));
 sg13g2_buf_8 clkbuf_5_30_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_30_0_clk));
 sg13g2_buf_8 clkbuf_5_31_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_31_0_clk));
 sg13g2_buf_8 clkbuf_6_0__f_clk (.A(clknet_5_0_0_clk),
    .X(clknet_6_0__leaf_clk));
 sg13g2_buf_8 clkbuf_6_1__f_clk (.A(clknet_5_0_0_clk),
    .X(clknet_6_1__leaf_clk));
 sg13g2_buf_8 clkbuf_6_2__f_clk (.A(clknet_5_1_0_clk),
    .X(clknet_6_2__leaf_clk));
 sg13g2_buf_8 clkbuf_6_3__f_clk (.A(clknet_5_1_0_clk),
    .X(clknet_6_3__leaf_clk));
 sg13g2_buf_8 clkbuf_6_4__f_clk (.A(clknet_5_2_0_clk),
    .X(clknet_6_4__leaf_clk));
 sg13g2_buf_8 clkbuf_6_5__f_clk (.A(clknet_5_2_0_clk),
    .X(clknet_6_5__leaf_clk));
 sg13g2_buf_8 clkbuf_6_6__f_clk (.A(clknet_5_3_0_clk),
    .X(clknet_6_6__leaf_clk));
 sg13g2_buf_8 clkbuf_6_7__f_clk (.A(clknet_5_3_0_clk),
    .X(clknet_6_7__leaf_clk));
 sg13g2_buf_8 clkbuf_6_8__f_clk (.A(clknet_5_4_0_clk),
    .X(clknet_6_8__leaf_clk));
 sg13g2_buf_8 clkbuf_6_9__f_clk (.A(clknet_5_4_0_clk),
    .X(clknet_6_9__leaf_clk));
 sg13g2_buf_8 clkbuf_6_10__f_clk (.A(clknet_5_5_0_clk),
    .X(clknet_6_10__leaf_clk));
 sg13g2_buf_8 clkbuf_6_11__f_clk (.A(clknet_5_5_0_clk),
    .X(clknet_6_11__leaf_clk));
 sg13g2_buf_8 clkbuf_6_12__f_clk (.A(clknet_5_6_0_clk),
    .X(clknet_6_12__leaf_clk));
 sg13g2_buf_8 clkbuf_6_13__f_clk (.A(clknet_5_6_0_clk),
    .X(clknet_6_13__leaf_clk));
 sg13g2_buf_8 clkbuf_6_14__f_clk (.A(clknet_5_7_0_clk),
    .X(clknet_6_14__leaf_clk));
 sg13g2_buf_8 clkbuf_6_15__f_clk (.A(clknet_5_7_0_clk),
    .X(clknet_6_15__leaf_clk));
 sg13g2_buf_8 clkbuf_6_16__f_clk (.A(clknet_5_8_0_clk),
    .X(clknet_6_16__leaf_clk));
 sg13g2_buf_8 clkbuf_6_17__f_clk (.A(clknet_5_8_0_clk),
    .X(clknet_6_17__leaf_clk));
 sg13g2_buf_8 clkbuf_6_18__f_clk (.A(clknet_5_9_0_clk),
    .X(clknet_6_18__leaf_clk));
 sg13g2_buf_8 clkbuf_6_19__f_clk (.A(clknet_5_9_0_clk),
    .X(clknet_6_19__leaf_clk));
 sg13g2_buf_8 clkbuf_6_20__f_clk (.A(clknet_5_10_0_clk),
    .X(clknet_6_20__leaf_clk));
 sg13g2_buf_8 clkbuf_6_21__f_clk (.A(clknet_5_10_0_clk),
    .X(clknet_6_21__leaf_clk));
 sg13g2_buf_8 clkbuf_6_22__f_clk (.A(clknet_5_11_0_clk),
    .X(clknet_6_22__leaf_clk));
 sg13g2_buf_8 clkbuf_6_23__f_clk (.A(clknet_5_11_0_clk),
    .X(clknet_6_23__leaf_clk));
 sg13g2_buf_8 clkbuf_6_24__f_clk (.A(clknet_5_12_0_clk),
    .X(clknet_6_24__leaf_clk));
 sg13g2_buf_8 clkbuf_6_25__f_clk (.A(clknet_5_12_0_clk),
    .X(clknet_6_25__leaf_clk));
 sg13g2_buf_8 clkbuf_6_26__f_clk (.A(clknet_5_13_0_clk),
    .X(clknet_6_26__leaf_clk));
 sg13g2_buf_8 clkbuf_6_27__f_clk (.A(clknet_5_13_0_clk),
    .X(clknet_6_27__leaf_clk));
 sg13g2_buf_8 clkbuf_6_28__f_clk (.A(clknet_5_14_0_clk),
    .X(clknet_6_28__leaf_clk));
 sg13g2_buf_8 clkbuf_6_29__f_clk (.A(clknet_5_14_0_clk),
    .X(clknet_6_29__leaf_clk));
 sg13g2_buf_8 clkbuf_6_30__f_clk (.A(clknet_5_15_0_clk),
    .X(clknet_6_30__leaf_clk));
 sg13g2_buf_8 clkbuf_6_31__f_clk (.A(clknet_5_15_0_clk),
    .X(clknet_6_31__leaf_clk));
 sg13g2_buf_8 clkbuf_6_32__f_clk (.A(clknet_5_16_0_clk),
    .X(clknet_6_32__leaf_clk));
 sg13g2_buf_8 clkbuf_6_33__f_clk (.A(clknet_5_16_0_clk),
    .X(clknet_6_33__leaf_clk));
 sg13g2_buf_8 clkbuf_6_34__f_clk (.A(clknet_5_17_0_clk),
    .X(clknet_6_34__leaf_clk));
 sg13g2_buf_8 clkbuf_6_35__f_clk (.A(clknet_5_17_0_clk),
    .X(clknet_6_35__leaf_clk));
 sg13g2_buf_8 clkbuf_6_36__f_clk (.A(clknet_5_18_0_clk),
    .X(clknet_6_36__leaf_clk));
 sg13g2_buf_8 clkbuf_6_37__f_clk (.A(clknet_5_18_0_clk),
    .X(clknet_6_37__leaf_clk));
 sg13g2_buf_8 clkbuf_6_38__f_clk (.A(clknet_5_19_0_clk),
    .X(clknet_6_38__leaf_clk));
 sg13g2_buf_8 clkbuf_6_39__f_clk (.A(clknet_5_19_0_clk),
    .X(clknet_6_39__leaf_clk));
 sg13g2_buf_8 clkbuf_6_40__f_clk (.A(clknet_5_20_0_clk),
    .X(clknet_6_40__leaf_clk));
 sg13g2_buf_8 clkbuf_6_41__f_clk (.A(clknet_5_20_0_clk),
    .X(clknet_6_41__leaf_clk));
 sg13g2_buf_8 clkbuf_6_42__f_clk (.A(clknet_5_21_0_clk),
    .X(clknet_6_42__leaf_clk));
 sg13g2_buf_8 clkbuf_6_43__f_clk (.A(clknet_5_21_0_clk),
    .X(clknet_6_43__leaf_clk));
 sg13g2_buf_8 clkbuf_6_44__f_clk (.A(clknet_5_22_0_clk),
    .X(clknet_6_44__leaf_clk));
 sg13g2_buf_8 clkbuf_6_45__f_clk (.A(clknet_5_22_0_clk),
    .X(clknet_6_45__leaf_clk));
 sg13g2_buf_8 clkbuf_6_46__f_clk (.A(clknet_5_23_0_clk),
    .X(clknet_6_46__leaf_clk));
 sg13g2_buf_8 clkbuf_6_47__f_clk (.A(clknet_5_23_0_clk),
    .X(clknet_6_47__leaf_clk));
 sg13g2_buf_8 clkbuf_6_48__f_clk (.A(clknet_5_24_0_clk),
    .X(clknet_6_48__leaf_clk));
 sg13g2_buf_8 clkbuf_6_49__f_clk (.A(clknet_5_24_0_clk),
    .X(clknet_6_49__leaf_clk));
 sg13g2_buf_8 clkbuf_6_50__f_clk (.A(clknet_5_25_0_clk),
    .X(clknet_6_50__leaf_clk));
 sg13g2_buf_8 clkbuf_6_51__f_clk (.A(clknet_5_25_0_clk),
    .X(clknet_6_51__leaf_clk));
 sg13g2_buf_8 clkbuf_6_52__f_clk (.A(clknet_5_26_0_clk),
    .X(clknet_6_52__leaf_clk));
 sg13g2_buf_8 clkbuf_6_53__f_clk (.A(clknet_5_26_0_clk),
    .X(clknet_6_53__leaf_clk));
 sg13g2_buf_8 clkbuf_6_54__f_clk (.A(clknet_5_27_0_clk),
    .X(clknet_6_54__leaf_clk));
 sg13g2_buf_8 clkbuf_6_55__f_clk (.A(clknet_5_27_0_clk),
    .X(clknet_6_55__leaf_clk));
 sg13g2_buf_8 clkbuf_6_56__f_clk (.A(clknet_5_28_0_clk),
    .X(clknet_6_56__leaf_clk));
 sg13g2_buf_8 clkbuf_6_57__f_clk (.A(clknet_5_28_0_clk),
    .X(clknet_6_57__leaf_clk));
 sg13g2_buf_8 clkbuf_6_58__f_clk (.A(clknet_5_29_0_clk),
    .X(clknet_6_58__leaf_clk));
 sg13g2_buf_8 clkbuf_6_59__f_clk (.A(clknet_5_29_0_clk),
    .X(clknet_6_59__leaf_clk));
 sg13g2_buf_8 clkbuf_6_60__f_clk (.A(clknet_5_30_0_clk),
    .X(clknet_6_60__leaf_clk));
 sg13g2_buf_8 clkbuf_6_61__f_clk (.A(clknet_5_30_0_clk),
    .X(clknet_6_61__leaf_clk));
 sg13g2_buf_8 clkbuf_6_62__f_clk (.A(clknet_5_31_0_clk),
    .X(clknet_6_62__leaf_clk));
 sg13g2_buf_8 clkbuf_6_63__f_clk (.A(clknet_5_31_0_clk),
    .X(clknet_6_63__leaf_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_6_7__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_6_15__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_6_23__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_6_27__leaf_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_6_31__leaf_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_6_39__leaf_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_6_43__leaf_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_6_47__leaf_clk));
 sg13g2_buf_8 clkload8 (.A(clknet_6_55__leaf_clk));
 sg13g2_buf_8 clkload9 (.A(clknet_6_59__leaf_clk));
 sg13g2_buf_8 clkload10 (.A(clknet_6_63__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_leaf_244_clk));
 sg13g2_inv_2 clkload12 (.A(clknet_leaf_239_clk));
 sg13g2_buf_8 clkload13 (.A(clknet_leaf_210_clk));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_70_clk));
 sg13g2_inv_1 clkload15 (.A(clknet_leaf_27_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_46_clk));
 sg13g2_inv_8 clkload17 (.A(clknet_leaf_76_clk));
 sg13g2_inv_4 clkload18 (.A(clknet_leaf_71_clk));
 sg13g2_buf_8 clkload19 (.A(clknet_leaf_43_clk));
 sg13g2_inv_4 clkload20 (.A(clknet_leaf_79_clk));
 sg13g2_buf_8 clkload21 (.A(clknet_leaf_75_clk));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_105_clk));
 sg13g2_inv_1 clkload23 (.A(clknet_leaf_128_clk));
 sg13g2_inv_2 clkload24 (.A(clknet_leaf_131_clk));
 sg13g2_inv_4 clkload25 (.A(clknet_leaf_98_clk));
 sg13g2_inv_4 clkload26 (.A(clknet_leaf_99_clk));
 sg13g2_inv_2 clkload27 (.A(clknet_leaf_102_clk));
 sg13g2_inv_4 clkload28 (.A(clknet_leaf_129_clk));
 sg13g2_inv_1 clkload29 (.A(clknet_leaf_106_clk));
 sg13g2_inv_1 clkload30 (.A(clknet_leaf_113_clk));
 sg13g2_inv_1 clkload31 (.A(clknet_leaf_115_clk));
 sg13g2_inv_1 clkload32 (.A(clknet_leaf_110_clk));
 sg13g2_buf_8 rebuffer1 (.A(_12839_),
    .X(net1064));
 sg13g2_buf_8 rebuffer2 (.A(_15899_),
    .X(net1065));
 sg13g2_buf_2 rebuffer3 (.A(_09614_),
    .X(net1066));
 sg13g2_buf_1 rebuffer4 (.A(net1066),
    .X(net1067));
 sg13g2_buf_8 rebuffer5 (.A(_15145_),
    .X(net1068));
 sg13g2_buf_1 rebuffer6 (.A(net1068),
    .X(net1069));
 sg13g2_buf_8 rebuffer7 (.A(_04398_),
    .X(net1070));
 sg13g2_buf_1 rebuffer8 (.A(net1070),
    .X(net1071));
 sg13g2_buf_8 rebuffer9 (.A(_15052_),
    .X(net1072));
 sg13g2_buf_8 rebuffer10 (.A(_15101_),
    .X(net1073));
 sg13g2_buf_8 rebuffer11 (.A(_11788_),
    .X(net1074));
 sg13g2_buf_8 rebuffer12 (.A(_15085_),
    .X(net1075));
 sg13g2_buf_1 rebuffer13 (.A(_15168_),
    .X(net1076));
 sg13g2_buf_2 rebuffer14 (.A(_08557_),
    .X(net1077));
 sg13g2_buf_1 rebuffer15 (.A(net1077),
    .X(net1078));
 sg13g2_buf_2 rebuffer16 (.A(_15133_),
    .X(net1079));
 sg13g2_buf_2 rebuffer17 (.A(_04583_),
    .X(net1080));
 sg13g2_buf_1 rebuffer18 (.A(net1080),
    .X(net1081));
 sg13g2_buf_2 rebuffer19 (.A(_15076_),
    .X(net1082));
 sg13g2_buf_8 rebuffer20 (.A(_08117_),
    .X(net1083));
 sg13g2_buf_2 rebuffer21 (.A(_15050_),
    .X(net1084));
 sg13g2_buf_8 rebuffer22 (.A(_15121_),
    .X(net1085));
 sg13g2_buf_8 rebuffer23 (.A(_08514_),
    .X(net1086));
 sg13g2_buf_2 rebuffer24 (.A(_15093_),
    .X(net1087));
 sg13g2_buf_1 rebuffer25 (.A(_15045_),
    .X(net1088));
 sg13g2_buf_1 rebuffer26 (.A(_15045_),
    .X(net1089));
 sg13g2_buf_1 rebuffer27 (.A(_15045_),
    .X(net1090));
 sg13g2_buf_2 rebuffer28 (.A(_15043_),
    .X(net1091));
 sg13g2_buf_8 rebuffer29 (.A(_15089_),
    .X(net1092));
 sg13g2_buf_2 rebuffer30 (.A(_16470_),
    .X(net1093));
 sg13g2_buf_8 rebuffer31 (.A(_10184_),
    .X(net1094));
 sg13g2_buf_8 rebuffer32 (.A(_15070_),
    .X(net1095));
 sg13g2_buf_2 rebuffer33 (.A(_15021_),
    .X(net1096));
 sg13g2_buf_2 rebuffer34 (.A(_08138_),
    .X(net1097));
 sg13g2_buf_1 rebuffer35 (.A(net1097),
    .X(net1098));
 sg13g2_buf_1 rebuffer36 (.A(_15140_),
    .X(net1099));
 sg13g2_buf_2 rebuffer37 (.A(_15060_),
    .X(net1100));
 sg13g2_buf_2 rebuffer38 (.A(_16276_),
    .X(net1101));
 sg13g2_buf_1 rebuffer39 (.A(net1131),
    .X(net1102));
 sg13g2_buf_1 rebuffer40 (.A(_15079_),
    .X(net1103));
 sg13g2_buf_8 rebuffer41 (.A(_05147_),
    .X(net1104));
 sg13g2_buf_1 rebuffer42 (.A(net1131),
    .X(net1105));
 sg13g2_buf_1 rebuffer43 (.A(_15035_),
    .X(net1106));
 sg13g2_buf_2 rebuffer44 (.A(_15033_),
    .X(net1107));
 sg13g2_buf_2 rebuffer45 (.A(_16026_),
    .X(net1108));
 sg13g2_buf_8 rebuffer46 (.A(_04421_),
    .X(net1109));
 sg13g2_buf_1 rebuffer47 (.A(_15095_),
    .X(net1110));
 sg13g2_buf_2 rebuffer48 (.A(_16748_),
    .X(net1111));
 sg13g2_buf_1 rebuffer49 (.A(net1141),
    .X(net1112));
 sg13g2_buf_1 rebuffer50 (.A(_15019_),
    .X(net1113));
 sg13g2_buf_1 rebuffer51 (.A(_15019_),
    .X(net1114));
 sg13g2_buf_1 rebuffer52 (.A(_15124_),
    .X(net1115));
 sg13g2_buf_1 rebuffer53 (.A(_15011_),
    .X(net1116));
 sg13g2_buf_1 rebuffer54 (.A(net1118),
    .X(net1117));
 sg13g2_buf_1 rebuffer55 (.A(_15154_),
    .X(net1118));
 sg13g2_buf_1 rebuffer56 (.A(_15157_),
    .X(net1119));
 sg13g2_buf_1 rebuffer57 (.A(_15157_),
    .X(net1120));
 sg13g2_buf_2 rebuffer58 (.A(_14464_),
    .X(net1121));
 sg13g2_buf_1 rebuffer59 (.A(_15094_),
    .X(net1122));
 sg13g2_buf_8 rebuffer60 (.A(_15854_),
    .X(net1123));
 sg13g2_buf_1 rebuffer61 (.A(_15167_),
    .X(net1124));
 sg13g2_buf_1 rebuffer62 (.A(_15013_),
    .X(net1125));
 sg13g2_buf_1 rebuffer63 (.A(_15119_),
    .X(net1126));
 sg13g2_buf_1 rebuffer64 (.A(_15119_),
    .X(net1127));
 sg13g2_buf_1 rebuffer65 (.A(_15110_),
    .X(net1128));
 sg13g2_buf_1 rebuffer66 (.A(_15110_),
    .X(net1129));
 sg13g2_buf_1 rebuffer67 (.A(net1079),
    .X(net1130));
 sg13g2_buf_1 rebuffer68 (.A(_15158_),
    .X(net1131));
 sg13g2_buf_1 rebuffer69 (.A(_15023_),
    .X(net1132));
 sg13g2_buf_1 rebuffer70 (.A(net1087),
    .X(net1133));
 sg13g2_buf_1 rebuffer71 (.A(net5357),
    .X(net1134));
 sg13g2_buf_1 rebuffer72 (.A(_15163_),
    .X(net1135));
 sg13g2_buf_1 rebuffer73 (.A(_15163_),
    .X(net1136));
 sg13g2_buf_1 rebuffer74 (.A(net1107),
    .X(net1137));
 sg13g2_buf_2 rebuffer75 (.A(_16850_),
    .X(net1138));
 sg13g2_buf_16 rebuffer76 (.X(net1139),
    .A(net5190));
 sg13g2_buf_1 rebuffer77 (.A(net5314),
    .X(net1140));
 sg13g2_buf_2 rebuffer79 (.A(_16068_),
    .X(net1142));
 sg13g2_buf_2 rebuffer80 (.A(_11793_),
    .X(net1143));
 sg13g2_buf_1 rebuffer81 (.A(net1143),
    .X(net1144));
 sg13g2_buf_1 rebuffer82 (.A(_15165_),
    .X(net1145));
 sg13g2_dlygate4sd3_1 hold83 (.A(\u_trng.entropy_ff1 ),
    .X(net1146));
 sg13g2_dlygate4sd3_1 hold84 (.A(\u_inv.load_input ),
    .X(net1147));
 sg13g2_dlygate4sd3_1 hold85 (.A(_00459_),
    .X(net1148));
 sg13g2_dlygate4sd3_1 hold86 (.A(\perf_double[9] ),
    .X(net1149));
 sg13g2_dlygate4sd3_1 hold88 (.A(\u_trng.bit_cnt[2] ),
    .X(net1151));
 sg13g2_dlygate4sd3_1 hold89 (.A(_00166_),
    .X(net1152));
 sg13g2_dlygate4sd3_1 hold90 (.A(\byte_cnt[3] ),
    .X(net1153));
 sg13g2_dlygate4sd3_1 hold91 (.A(_00172_),
    .X(net1154));
 sg13g2_dlygate4sd3_1 hold92 (.A(\perf_total[5] ),
    .X(net1155));
 sg13g2_dlygate4sd3_1 hold93 (.A(_00732_),
    .X(net1156));
 sg13g2_dlygate4sd3_1 hold94 (.A(\perf_double[2] ),
    .X(net1157));
 sg13g2_dlygate4sd3_1 hold96 (.A(inv_go),
    .X(net1159));
 sg13g2_dlygate4sd3_1 hold97 (.A(_00163_),
    .X(net1160));
 sg13g2_dlygate4sd3_1 hold98 (.A(\perf_total[3] ),
    .X(net1161));
 sg13g2_dlygate4sd3_1 hold99 (.A(_00730_),
    .X(net1162));
 sg13g2_dlygate4sd3_1 hold100 (.A(\perf_triple[2] ),
    .X(net1163));
 sg13g2_dlygate4sd3_1 hold101 (.A(\perf_double[3] ),
    .X(net1164));
 sg13g2_dlygate4sd3_1 hold103 (.A(\byte_cnt[1] ),
    .X(net1166));
 sg13g2_dlygate4sd3_1 hold104 (.A(_18918_),
    .X(net1167));
 sg13g2_dlygate4sd3_1 hold105 (.A(_00170_),
    .X(net1168));
 sg13g2_dlygate4sd3_1 hold106 (.A(\perf_double[7] ),
    .X(net1169));
 sg13g2_dlygate4sd3_1 hold108 (.A(\u_inv.delta_reg[6] ),
    .X(net1171));
 sg13g2_dlygate4sd3_1 hold109 (.A(_01782_),
    .X(net1172));
 sg13g2_dlygate4sd3_1 hold110 (.A(\u_trng.bit_cnt[0] ),
    .X(net1173));
 sg13g2_dlygate4sd3_1 hold111 (.A(\byte_cnt[4] ),
    .X(net1174));
 sg13g2_dlygate4sd3_1 hold112 (.A(_18922_),
    .X(net1175));
 sg13g2_dlygate4sd3_1 hold113 (.A(\u_trng.have_prev ),
    .X(net1176));
 sg13g2_dlygate4sd3_1 hold114 (.A(_00457_),
    .X(net1177));
 sg13g2_dlygate4sd3_1 hold115 (.A(\inv_result[144] ),
    .X(net1178));
 sg13g2_dlygate4sd3_1 hold116 (.A(next_loaded),
    .X(net1179));
 sg13g2_dlygate4sd3_1 hold117 (.A(_19802_),
    .X(net1180));
 sg13g2_dlygate4sd3_1 hold118 (.A(_00447_),
    .X(net1181));
 sg13g2_dlygate4sd3_1 hold119 (.A(\inv_result[228] ),
    .X(net1182));
 sg13g2_dlygate4sd3_1 hold120 (.A(\perf_total[6] ),
    .X(net1183));
 sg13g2_dlygate4sd3_1 hold121 (.A(_03332_),
    .X(net1184));
 sg13g2_dlygate4sd3_1 hold122 (.A(\u_inv.f_reg[183] ),
    .X(net1185));
 sg13g2_dlygate4sd3_1 hold123 (.A(_01690_),
    .X(net1186));
 sg13g2_dlygate4sd3_1 hold124 (.A(\perf_total[0] ),
    .X(net1187));
 sg13g2_dlygate4sd3_1 hold125 (.A(\inv_cycles[5] ),
    .X(net1188));
 sg13g2_dlygate4sd3_1 hold126 (.A(_01792_),
    .X(net1189));
 sg13g2_dlygate4sd3_1 hold127 (.A(\inv_result[24] ),
    .X(net1190));
 sg13g2_dlygate4sd3_1 hold128 (.A(\u_inv.d_next[245] ),
    .X(net1191));
 sg13g2_dlygate4sd3_1 hold129 (.A(\shift_reg[7] ),
    .X(net1192));
 sg13g2_dlygate4sd3_1 hold130 (.A(\perf_total[4] ),
    .X(net1193));
 sg13g2_dlygate4sd3_1 hold131 (.A(_03328_),
    .X(net1194));
 sg13g2_dlygate4sd3_1 hold132 (.A(_00731_),
    .X(net1195));
 sg13g2_dlygate4sd3_1 hold133 (.A(\inv_result[34] ),
    .X(net1196));
 sg13g2_dlygate4sd3_1 hold134 (.A(\inv_result[172] ),
    .X(net1197));
 sg13g2_dlygate4sd3_1 hold135 (.A(\inv_result[198] ),
    .X(net1198));
 sg13g2_dlygate4sd3_1 hold136 (.A(\shift_reg[13] ),
    .X(net1199));
 sg13g2_dlygate4sd3_1 hold137 (.A(_00188_),
    .X(net1200));
 sg13g2_dlygate4sd3_1 hold138 (.A(\inv_result[18] ),
    .X(net1201));
 sg13g2_dlygate4sd3_1 hold139 (.A(\inv_result[98] ),
    .X(net1202));
 sg13g2_dlygate4sd3_1 hold140 (.A(\inv_cycles[4] ),
    .X(net1203));
 sg13g2_dlygate4sd3_1 hold141 (.A(_01791_),
    .X(net1204));
 sg13g2_dlygate4sd3_1 hold142 (.A(\inv_result[188] ),
    .X(net1205));
 sg13g2_dlygate4sd3_1 hold144 (.A(\inv_result[76] ),
    .X(net1207));
 sg13g2_dlygate4sd3_1 hold145 (.A(\inv_result[92] ),
    .X(net1208));
 sg13g2_dlygate4sd3_1 hold146 (.A(\inv_result[104] ),
    .X(net1209));
 sg13g2_dlygate4sd3_1 hold147 (.A(\inv_result[156] ),
    .X(net1210));
 sg13g2_dlygate4sd3_1 hold148 (.A(\u_inv.delta_reg[2] ),
    .X(net1211));
 sg13g2_dlygate4sd3_1 hold149 (.A(\inv_cycles[3] ),
    .X(net1212));
 sg13g2_dlygate4sd3_1 hold150 (.A(_01790_),
    .X(net1213));
 sg13g2_dlygate4sd3_1 hold151 (.A(\inv_result[116] ),
    .X(net1214));
 sg13g2_dlygate4sd3_1 hold152 (.A(\u_inv.delta_reg[3] ),
    .X(net1215));
 sg13g2_dlygate4sd3_1 hold153 (.A(\perf_triple[9] ),
    .X(net1216));
 sg13g2_dlygate4sd3_1 hold154 (.A(\u_inv.input_reg[211] ),
    .X(net1217));
 sg13g2_dlygate4sd3_1 hold155 (.A(_00118_),
    .X(net1218));
 sg13g2_dlygate4sd3_1 hold156 (.A(\inv_result[165] ),
    .X(net1219));
 sg13g2_dlygate4sd3_1 hold157 (.A(\inv_result[83] ),
    .X(net1220));
 sg13g2_dlygate4sd3_1 hold158 (.A(\perf_triple[1] ),
    .X(net1221));
 sg13g2_dlygate4sd3_1 hold159 (.A(\u_trng.bit_cnt[1] ),
    .X(net1222));
 sg13g2_dlygate4sd3_1 hold160 (.A(_00001_),
    .X(net1223));
 sg13g2_dlygate4sd3_1 hold161 (.A(\inv_result[219] ),
    .X(net1224));
 sg13g2_dlygate4sd3_1 hold162 (.A(\u_inv.delta_reg[5] ),
    .X(net1225));
 sg13g2_dlygate4sd3_1 hold163 (.A(\inv_result[226] ),
    .X(net1226));
 sg13g2_dlygate4sd3_1 hold164 (.A(\inv_result[155] ),
    .X(net1227));
 sg13g2_dlygate4sd3_1 hold165 (.A(\inv_result[187] ),
    .X(net1228));
 sg13g2_dlygate4sd3_1 hold166 (.A(_01181_),
    .X(net1229));
 sg13g2_dlygate4sd3_1 hold167 (.A(\inv_result[139] ),
    .X(net1230));
 sg13g2_dlygate4sd3_1 hold168 (.A(\inv_result[224] ),
    .X(net1231));
 sg13g2_dlygate4sd3_1 hold169 (.A(\inv_result[137] ),
    .X(net1232));
 sg13g2_dlygate4sd3_1 hold170 (.A(\inv_cycles[0] ),
    .X(net1233));
 sg13g2_dlygate4sd3_1 hold171 (.A(_01787_),
    .X(net1234));
 sg13g2_dlygate4sd3_1 hold172 (.A(\perf_double[4] ),
    .X(net1235));
 sg13g2_dlygate4sd3_1 hold174 (.A(\inv_result[205] ),
    .X(net1237));
 sg13g2_dlygate4sd3_1 hold175 (.A(\u_inv.d_next[50] ),
    .X(net1238));
 sg13g2_dlygate4sd3_1 hold176 (.A(_01300_),
    .X(net1239));
 sg13g2_dlygate4sd3_1 hold177 (.A(\inv_result[88] ),
    .X(net1240));
 sg13g2_dlygate4sd3_1 hold179 (.A(_17156_),
    .X(net1242));
 sg13g2_dlygate4sd3_1 hold180 (.A(_01380_),
    .X(net1243));
 sg13g2_dlygate4sd3_1 hold181 (.A(\inv_result[102] ),
    .X(net1244));
 sg13g2_dlygate4sd3_1 hold182 (.A(\inv_result[101] ),
    .X(net1245));
 sg13g2_dlygate4sd3_1 hold183 (.A(\inv_result[216] ),
    .X(net1246));
 sg13g2_dlygate4sd3_1 hold184 (.A(\inv_result[182] ),
    .X(net1247));
 sg13g2_dlygate4sd3_1 hold185 (.A(\inv_result[213] ),
    .X(net1248));
 sg13g2_dlygate4sd3_1 hold186 (.A(\u_inv.delta_reg[9] ),
    .X(net1249));
 sg13g2_dlygate4sd3_1 hold187 (.A(_01785_),
    .X(net1250));
 sg13g2_dlygate4sd3_1 hold188 (.A(\perf_double[5] ),
    .X(net1251));
 sg13g2_dlygate4sd3_1 hold189 (.A(\u_inv.f_reg[163] ),
    .X(net1252));
 sg13g2_dlygate4sd3_1 hold190 (.A(_01670_),
    .X(net1253));
 sg13g2_dlygate4sd3_1 hold191 (.A(\inv_result[107] ),
    .X(net1254));
 sg13g2_dlygate4sd3_1 hold192 (.A(\perf_double[6] ),
    .X(net1255));
 sg13g2_dlygate4sd3_1 hold193 (.A(\u_inv.input_reg[35] ),
    .X(net1256));
 sg13g2_dlygate4sd3_1 hold194 (.A(_01841_),
    .X(net1257));
 sg13g2_dlygate4sd3_1 hold195 (.A(\u_inv.input_reg[123] ),
    .X(net1258));
 sg13g2_dlygate4sd3_1 hold196 (.A(_00030_),
    .X(net1259));
 sg13g2_dlygate4sd3_1 hold197 (.A(\inv_result[149] ),
    .X(net1260));
 sg13g2_dlygate4sd3_1 hold198 (.A(\inv_result[163] ),
    .X(net1261));
 sg13g2_dlygate4sd3_1 hold199 (.A(\u_inv.input_reg[48] ),
    .X(net1262));
 sg13g2_dlygate4sd3_1 hold200 (.A(_01854_),
    .X(net1263));
 sg13g2_dlygate4sd3_1 hold201 (.A(\u_inv.input_reg[36] ),
    .X(net1264));
 sg13g2_dlygate4sd3_1 hold202 (.A(_01842_),
    .X(net1265));
 sg13g2_dlygate4sd3_1 hold203 (.A(\perf_total[2] ),
    .X(net1266));
 sg13g2_dlygate4sd3_1 hold204 (.A(_00729_),
    .X(net1267));
 sg13g2_dlygate4sd3_1 hold205 (.A(\u_inv.input_reg[32] ),
    .X(net1268));
 sg13g2_dlygate4sd3_1 hold206 (.A(_01838_),
    .X(net1269));
 sg13g2_dlygate4sd3_1 hold207 (.A(\inv_result[125] ),
    .X(net1270));
 sg13g2_dlygate4sd3_1 hold208 (.A(\u_inv.input_reg[132] ),
    .X(net1271));
 sg13g2_dlygate4sd3_1 hold209 (.A(_00039_),
    .X(net1272));
 sg13g2_dlygate4sd3_1 hold210 (.A(\inv_result[133] ),
    .X(net1273));
 sg13g2_dlygate4sd3_1 hold211 (.A(\u_inv.input_reg[12] ),
    .X(net1274));
 sg13g2_dlygate4sd3_1 hold212 (.A(_01818_),
    .X(net1275));
 sg13g2_dlygate4sd3_1 hold213 (.A(\u_inv.input_reg[107] ),
    .X(net1276));
 sg13g2_dlygate4sd3_1 hold214 (.A(_00014_),
    .X(net1277));
 sg13g2_dlygate4sd3_1 hold215 (.A(\inv_result[243] ),
    .X(net1278));
 sg13g2_dlygate4sd3_1 hold216 (.A(\perf_total[7] ),
    .X(net1279));
 sg13g2_dlygate4sd3_1 hold217 (.A(_03336_),
    .X(net1280));
 sg13g2_dlygate4sd3_1 hold218 (.A(_00736_),
    .X(net1281));
 sg13g2_dlygate4sd3_1 hold219 (.A(\u_inv.input_reg[192] ),
    .X(net1282));
 sg13g2_dlygate4sd3_1 hold220 (.A(_00099_),
    .X(net1283));
 sg13g2_dlygate4sd3_1 hold221 (.A(\u_inv.f_next[45] ),
    .X(net1284));
 sg13g2_dlygate4sd3_1 hold222 (.A(_00505_),
    .X(net1285));
 sg13g2_dlygate4sd3_1 hold223 (.A(\perf_double[8] ),
    .X(net1286));
 sg13g2_dlygate4sd3_1 hold224 (.A(\u_inv.input_reg[173] ),
    .X(net1287));
 sg13g2_dlygate4sd3_1 hold225 (.A(_00080_),
    .X(net1288));
 sg13g2_dlygate4sd3_1 hold226 (.A(\u_inv.input_reg[237] ),
    .X(net1289));
 sg13g2_dlygate4sd3_1 hold227 (.A(_00144_),
    .X(net1290));
 sg13g2_dlygate4sd3_1 hold228 (.A(\inv_result[208] ),
    .X(net1291));
 sg13g2_dlygate4sd3_1 hold229 (.A(\inv_result[173] ),
    .X(net1292));
 sg13g2_dlygate4sd3_1 hold230 (.A(\u_inv.input_reg[8] ),
    .X(net1293));
 sg13g2_dlygate4sd3_1 hold231 (.A(_01814_),
    .X(net1294));
 sg13g2_dlygate4sd3_1 hold232 (.A(\u_inv.input_reg[4] ),
    .X(net1295));
 sg13g2_dlygate4sd3_1 hold233 (.A(_01810_),
    .X(net1296));
 sg13g2_dlygate4sd3_1 hold234 (.A(\inv_result[147] ),
    .X(net1297));
 sg13g2_dlygate4sd3_1 hold235 (.A(\inv_result[77] ),
    .X(net1298));
 sg13g2_dlygate4sd3_1 hold236 (.A(\u_inv.input_reg[29] ),
    .X(net1299));
 sg13g2_dlygate4sd3_1 hold237 (.A(_01835_),
    .X(net1300));
 sg13g2_dlygate4sd3_1 hold238 (.A(\inv_result[232] ),
    .X(net1301));
 sg13g2_dlygate4sd3_1 hold239 (.A(\u_inv.input_reg[14] ),
    .X(net1302));
 sg13g2_dlygate4sd3_1 hold240 (.A(_01820_),
    .X(net1303));
 sg13g2_dlygate4sd3_1 hold241 (.A(\u_inv.input_reg[39] ),
    .X(net1304));
 sg13g2_dlygate4sd3_1 hold242 (.A(_01845_),
    .X(net1305));
 sg13g2_dlygate4sd3_1 hold243 (.A(\u_inv.input_reg[0] ),
    .X(net1306));
 sg13g2_dlygate4sd3_1 hold244 (.A(_01806_),
    .X(net1307));
 sg13g2_dlygate4sd3_1 hold245 (.A(\u_inv.input_reg[247] ),
    .X(net1308));
 sg13g2_dlygate4sd3_1 hold246 (.A(_00154_),
    .X(net1309));
 sg13g2_dlygate4sd3_1 hold247 (.A(\u_inv.input_reg[217] ),
    .X(net1310));
 sg13g2_dlygate4sd3_1 hold248 (.A(_00124_),
    .X(net1311));
 sg13g2_dlygate4sd3_1 hold249 (.A(\u_inv.input_reg[220] ),
    .X(net1312));
 sg13g2_dlygate4sd3_1 hold250 (.A(_00127_),
    .X(net1313));
 sg13g2_dlygate4sd3_1 hold251 (.A(\u_inv.input_reg[253] ),
    .X(net1314));
 sg13g2_dlygate4sd3_1 hold252 (.A(_00160_),
    .X(net1315));
 sg13g2_dlygate4sd3_1 hold253 (.A(\u_inv.input_reg[120] ),
    .X(net1316));
 sg13g2_dlygate4sd3_1 hold254 (.A(_00027_),
    .X(net1317));
 sg13g2_dlygate4sd3_1 hold255 (.A(\u_inv.input_reg[27] ),
    .X(net1318));
 sg13g2_dlygate4sd3_1 hold256 (.A(_01833_),
    .X(net1319));
 sg13g2_dlygate4sd3_1 hold257 (.A(\u_inv.input_reg[241] ),
    .X(net1320));
 sg13g2_dlygate4sd3_1 hold258 (.A(_00148_),
    .X(net1321));
 sg13g2_dlygate4sd3_1 hold259 (.A(\u_inv.input_reg[99] ),
    .X(net1322));
 sg13g2_dlygate4sd3_1 hold260 (.A(_00006_),
    .X(net1323));
 sg13g2_dlygate4sd3_1 hold261 (.A(\shift_reg[9] ),
    .X(net1324));
 sg13g2_dlygate4sd3_1 hold262 (.A(_00184_),
    .X(net1325));
 sg13g2_dlygate4sd3_1 hold263 (.A(\inv_result[93] ),
    .X(net1326));
 sg13g2_dlygate4sd3_1 hold264 (.A(\u_inv.input_reg[240] ),
    .X(net1327));
 sg13g2_dlygate4sd3_1 hold265 (.A(_00147_),
    .X(net1328));
 sg13g2_dlygate4sd3_1 hold266 (.A(\u_inv.input_reg[172] ),
    .X(net1329));
 sg13g2_dlygate4sd3_1 hold267 (.A(_00079_),
    .X(net1330));
 sg13g2_dlygate4sd3_1 hold268 (.A(\u_inv.input_reg[10] ),
    .X(net1331));
 sg13g2_dlygate4sd3_1 hold269 (.A(_01816_),
    .X(net1332));
 sg13g2_dlygate4sd3_1 hold270 (.A(\u_inv.input_reg[239] ),
    .X(net1333));
 sg13g2_dlygate4sd3_1 hold271 (.A(_00146_),
    .X(net1334));
 sg13g2_dlygate4sd3_1 hold272 (.A(\u_inv.input_reg[23] ),
    .X(net1335));
 sg13g2_dlygate4sd3_1 hold273 (.A(_01829_),
    .X(net1336));
 sg13g2_dlygate4sd3_1 hold274 (.A(\u_inv.input_reg[143] ),
    .X(net1337));
 sg13g2_dlygate4sd3_1 hold275 (.A(_00050_),
    .X(net1338));
 sg13g2_dlygate4sd3_1 hold276 (.A(\inv_result[128] ),
    .X(net1339));
 sg13g2_dlygate4sd3_1 hold277 (.A(\u_inv.input_reg[200] ),
    .X(net1340));
 sg13g2_dlygate4sd3_1 hold278 (.A(_00107_),
    .X(net1341));
 sg13g2_dlygate4sd3_1 hold279 (.A(\u_inv.delta_reg[8] ),
    .X(net1342));
 sg13g2_dlygate4sd3_1 hold280 (.A(\u_inv.input_reg[26] ),
    .X(net1343));
 sg13g2_dlygate4sd3_1 hold281 (.A(_01832_),
    .X(net1344));
 sg13g2_dlygate4sd3_1 hold282 (.A(\u_inv.input_reg[34] ),
    .X(net1345));
 sg13g2_dlygate4sd3_1 hold283 (.A(_01840_),
    .X(net1346));
 sg13g2_dlygate4sd3_1 hold284 (.A(\u_inv.f_reg[2] ),
    .X(net1347));
 sg13g2_dlygate4sd3_1 hold285 (.A(_01509_),
    .X(net1348));
 sg13g2_dlygate4sd3_1 hold286 (.A(\u_inv.input_reg[46] ),
    .X(net1349));
 sg13g2_dlygate4sd3_1 hold287 (.A(_01852_),
    .X(net1350));
 sg13g2_dlygate4sd3_1 hold288 (.A(\u_inv.input_reg[38] ),
    .X(net1351));
 sg13g2_dlygate4sd3_1 hold289 (.A(_01844_),
    .X(net1352));
 sg13g2_dlygate4sd3_1 hold290 (.A(\u_inv.f_reg[37] ),
    .X(net1353));
 sg13g2_dlygate4sd3_1 hold291 (.A(_01544_),
    .X(net1354));
 sg13g2_dlygate4sd3_1 hold292 (.A(\inv_result[185] ),
    .X(net1355));
 sg13g2_dlygate4sd3_1 hold293 (.A(\u_inv.input_reg[166] ),
    .X(net1356));
 sg13g2_dlygate4sd3_1 hold294 (.A(_00073_),
    .X(net1357));
 sg13g2_dlygate4sd3_1 hold295 (.A(\u_inv.input_reg[84] ),
    .X(net1358));
 sg13g2_dlygate4sd3_1 hold296 (.A(_01890_),
    .X(net1359));
 sg13g2_dlygate4sd3_1 hold297 (.A(\inv_result[68] ),
    .X(net1360));
 sg13g2_dlygate4sd3_1 hold298 (.A(\trng_data[7] ),
    .X(net1361));
 sg13g2_dlygate4sd3_1 hold299 (.A(_00456_),
    .X(net1362));
 sg13g2_dlygate4sd3_1 hold300 (.A(\u_inv.input_reg[105] ),
    .X(net1363));
 sg13g2_dlygate4sd3_1 hold301 (.A(_00012_),
    .X(net1364));
 sg13g2_dlygate4sd3_1 hold302 (.A(\u_inv.input_reg[97] ),
    .X(net1365));
 sg13g2_dlygate4sd3_1 hold303 (.A(_00004_),
    .X(net1366));
 sg13g2_dlygate4sd3_1 hold304 (.A(\u_inv.input_reg[246] ),
    .X(net1367));
 sg13g2_dlygate4sd3_1 hold305 (.A(_00153_),
    .X(net1368));
 sg13g2_dlygate4sd3_1 hold306 (.A(\u_inv.input_reg[18] ),
    .X(net1369));
 sg13g2_dlygate4sd3_1 hold307 (.A(_01824_),
    .X(net1370));
 sg13g2_dlygate4sd3_1 hold308 (.A(\u_inv.input_reg[87] ),
    .X(net1371));
 sg13g2_dlygate4sd3_1 hold309 (.A(_01893_),
    .X(net1372));
 sg13g2_dlygate4sd3_1 hold310 (.A(\u_inv.input_reg[56] ),
    .X(net1373));
 sg13g2_dlygate4sd3_1 hold311 (.A(_01862_),
    .X(net1374));
 sg13g2_dlygate4sd3_1 hold312 (.A(\u_inv.input_reg[20] ),
    .X(net1375));
 sg13g2_dlygate4sd3_1 hold313 (.A(_01826_),
    .X(net1376));
 sg13g2_dlygate4sd3_1 hold314 (.A(\u_inv.input_reg[233] ),
    .X(net1377));
 sg13g2_dlygate4sd3_1 hold315 (.A(_00140_),
    .X(net1378));
 sg13g2_dlygate4sd3_1 hold316 (.A(\u_inv.input_reg[28] ),
    .X(net1379));
 sg13g2_dlygate4sd3_1 hold317 (.A(_01834_),
    .X(net1380));
 sg13g2_dlygate4sd3_1 hold318 (.A(\u_inv.input_reg[131] ),
    .X(net1381));
 sg13g2_dlygate4sd3_1 hold319 (.A(_00038_),
    .X(net1382));
 sg13g2_dlygate4sd3_1 hold320 (.A(\inv_result[7] ),
    .X(net1383));
 sg13g2_dlygate4sd3_1 hold321 (.A(\inv_result[234] ),
    .X(net1384));
 sg13g2_dlygate4sd3_1 hold322 (.A(\u_inv.input_reg[232] ),
    .X(net1385));
 sg13g2_dlygate4sd3_1 hold323 (.A(_00139_),
    .X(net1386));
 sg13g2_dlygate4sd3_1 hold324 (.A(\perf_double[1] ),
    .X(net1387));
 sg13g2_dlygate4sd3_1 hold326 (.A(\u_inv.d_next[11] ),
    .X(net1389));
 sg13g2_dlygate4sd3_1 hold327 (.A(_01261_),
    .X(net1390));
 sg13g2_dlygate4sd3_1 hold328 (.A(\u_inv.input_reg[9] ),
    .X(net1391));
 sg13g2_dlygate4sd3_1 hold329 (.A(_01815_),
    .X(net1392));
 sg13g2_dlygate4sd3_1 hold330 (.A(\u_inv.input_reg[181] ),
    .X(net1393));
 sg13g2_dlygate4sd3_1 hold331 (.A(_00088_),
    .X(net1394));
 sg13g2_dlygate4sd3_1 hold332 (.A(\u_inv.input_reg[226] ),
    .X(net1395));
 sg13g2_dlygate4sd3_1 hold333 (.A(_00133_),
    .X(net1396));
 sg13g2_dlygate4sd3_1 hold334 (.A(\u_inv.input_reg[112] ),
    .X(net1397));
 sg13g2_dlygate4sd3_1 hold335 (.A(_00019_),
    .X(net1398));
 sg13g2_dlygate4sd3_1 hold336 (.A(\u_inv.input_reg[224] ),
    .X(net1399));
 sg13g2_dlygate4sd3_1 hold337 (.A(_00131_),
    .X(net1400));
 sg13g2_dlygate4sd3_1 hold338 (.A(\u_inv.input_reg[230] ),
    .X(net1401));
 sg13g2_dlygate4sd3_1 hold339 (.A(_00137_),
    .X(net1402));
 sg13g2_dlygate4sd3_1 hold340 (.A(\inv_result[109] ),
    .X(net1403));
 sg13g2_dlygate4sd3_1 hold341 (.A(\u_inv.input_reg[178] ),
    .X(net1404));
 sg13g2_dlygate4sd3_1 hold342 (.A(_00085_),
    .X(net1405));
 sg13g2_dlygate4sd3_1 hold343 (.A(\inv_result[72] ),
    .X(net1406));
 sg13g2_dlygate4sd3_1 hold344 (.A(\inv_result[43] ),
    .X(net1407));
 sg13g2_dlygate4sd3_1 hold346 (.A(\u_inv.input_reg[103] ),
    .X(net1409));
 sg13g2_dlygate4sd3_1 hold347 (.A(_00010_),
    .X(net1410));
 sg13g2_dlygate4sd3_1 hold348 (.A(\u_inv.input_reg[44] ),
    .X(net1411));
 sg13g2_dlygate4sd3_1 hold349 (.A(_01850_),
    .X(net1412));
 sg13g2_dlygate4sd3_1 hold350 (.A(\u_inv.input_reg[156] ),
    .X(net1413));
 sg13g2_dlygate4sd3_1 hold351 (.A(_00063_),
    .X(net1414));
 sg13g2_dlygate4sd3_1 hold352 (.A(\inv_cycles[9] ),
    .X(net1415));
 sg13g2_dlygate4sd3_1 hold353 (.A(_01796_),
    .X(net1416));
 sg13g2_dlygate4sd3_1 hold354 (.A(\u_inv.input_reg[63] ),
    .X(net1417));
 sg13g2_dlygate4sd3_1 hold355 (.A(_01869_),
    .X(net1418));
 sg13g2_dlygate4sd3_1 hold356 (.A(\u_inv.f_next[105] ),
    .X(net1419));
 sg13g2_dlygate4sd3_1 hold357 (.A(\u_inv.input_reg[33] ),
    .X(net1420));
 sg13g2_dlygate4sd3_1 hold358 (.A(_01839_),
    .X(net1421));
 sg13g2_dlygate4sd3_1 hold359 (.A(\inv_result[231] ),
    .X(net1422));
 sg13g2_dlygate4sd3_1 hold360 (.A(\u_inv.input_reg[83] ),
    .X(net1423));
 sg13g2_dlygate4sd3_1 hold361 (.A(_01889_),
    .X(net1424));
 sg13g2_dlygate4sd3_1 hold362 (.A(\u_inv.input_reg[199] ),
    .X(net1425));
 sg13g2_dlygate4sd3_1 hold363 (.A(_00106_),
    .X(net1426));
 sg13g2_dlygate4sd3_1 hold364 (.A(\u_inv.input_reg[243] ),
    .X(net1427));
 sg13g2_dlygate4sd3_1 hold365 (.A(_00150_),
    .X(net1428));
 sg13g2_dlygate4sd3_1 hold366 (.A(\u_inv.input_reg[117] ),
    .X(net1429));
 sg13g2_dlygate4sd3_1 hold367 (.A(_00024_),
    .X(net1430));
 sg13g2_dlygate4sd3_1 hold368 (.A(\u_inv.f_reg[109] ),
    .X(net1431));
 sg13g2_dlygate4sd3_1 hold369 (.A(_01616_),
    .X(net1432));
 sg13g2_dlygate4sd3_1 hold370 (.A(\u_inv.f_reg[118] ),
    .X(net1433));
 sg13g2_dlygate4sd3_1 hold371 (.A(_01625_),
    .X(net1434));
 sg13g2_dlygate4sd3_1 hold372 (.A(\u_inv.input_reg[89] ),
    .X(net1435));
 sg13g2_dlygate4sd3_1 hold373 (.A(_01895_),
    .X(net1436));
 sg13g2_dlygate4sd3_1 hold374 (.A(\inv_result[148] ),
    .X(net1437));
 sg13g2_dlygate4sd3_1 hold375 (.A(\u_inv.input_reg[236] ),
    .X(net1438));
 sg13g2_dlygate4sd3_1 hold376 (.A(_00143_),
    .X(net1439));
 sg13g2_dlygate4sd3_1 hold377 (.A(\inv_result[164] ),
    .X(net1440));
 sg13g2_dlygate4sd3_1 hold378 (.A(\inv_result[143] ),
    .X(net1441));
 sg13g2_dlygate4sd3_1 hold379 (.A(\u_inv.f_reg[5] ),
    .X(net1442));
 sg13g2_dlygate4sd3_1 hold380 (.A(_01512_),
    .X(net1443));
 sg13g2_dlygate4sd3_1 hold381 (.A(\u_inv.f_reg[44] ),
    .X(net1444));
 sg13g2_dlygate4sd3_1 hold382 (.A(_01551_),
    .X(net1445));
 sg13g2_dlygate4sd3_1 hold383 (.A(\u_inv.f_next[37] ),
    .X(net1446));
 sg13g2_dlygate4sd3_1 hold384 (.A(_00497_),
    .X(net1447));
 sg13g2_dlygate4sd3_1 hold385 (.A(\u_inv.input_reg[11] ),
    .X(net1448));
 sg13g2_dlygate4sd3_1 hold386 (.A(_01817_),
    .X(net1449));
 sg13g2_dlygate4sd3_1 hold387 (.A(\u_inv.input_reg[24] ),
    .X(net1450));
 sg13g2_dlygate4sd3_1 hold388 (.A(_01830_),
    .X(net1451));
 sg13g2_dlygate4sd3_1 hold389 (.A(\u_inv.input_reg[17] ),
    .X(net1452));
 sg13g2_dlygate4sd3_1 hold390 (.A(_01823_),
    .X(net1453));
 sg13g2_dlygate4sd3_1 hold391 (.A(\u_inv.input_reg[162] ),
    .X(net1454));
 sg13g2_dlygate4sd3_1 hold392 (.A(_00069_),
    .X(net1455));
 sg13g2_dlygate4sd3_1 hold393 (.A(\u_inv.input_reg[198] ),
    .X(net1456));
 sg13g2_dlygate4sd3_1 hold394 (.A(_00105_),
    .X(net1457));
 sg13g2_dlygate4sd3_1 hold395 (.A(\inv_result[141] ),
    .X(net1458));
 sg13g2_dlygate4sd3_1 hold396 (.A(\inv_result[159] ),
    .X(net1459));
 sg13g2_dlygate4sd3_1 hold397 (.A(\u_inv.input_reg[88] ),
    .X(net1460));
 sg13g2_dlygate4sd3_1 hold398 (.A(_01894_),
    .X(net1461));
 sg13g2_dlygate4sd3_1 hold399 (.A(\u_inv.input_reg[191] ),
    .X(net1462));
 sg13g2_dlygate4sd3_1 hold400 (.A(_00098_),
    .X(net1463));
 sg13g2_dlygate4sd3_1 hold401 (.A(\inv_result[189] ),
    .X(net1464));
 sg13g2_dlygate4sd3_1 hold402 (.A(\u_inv.input_reg[59] ),
    .X(net1465));
 sg13g2_dlygate4sd3_1 hold403 (.A(_01865_),
    .X(net1466));
 sg13g2_dlygate4sd3_1 hold404 (.A(\u_inv.input_reg[54] ),
    .X(net1467));
 sg13g2_dlygate4sd3_1 hold405 (.A(_01860_),
    .X(net1468));
 sg13g2_dlygate4sd3_1 hold406 (.A(\u_inv.input_reg[218] ),
    .X(net1469));
 sg13g2_dlygate4sd3_1 hold407 (.A(_00125_),
    .X(net1470));
 sg13g2_dlygate4sd3_1 hold408 (.A(\u_inv.input_reg[73] ),
    .X(net1471));
 sg13g2_dlygate4sd3_1 hold409 (.A(_01879_),
    .X(net1472));
 sg13g2_dlygate4sd3_1 hold410 (.A(\u_inv.f_next[145] ),
    .X(net1473));
 sg13g2_dlygate4sd3_1 hold411 (.A(_00605_),
    .X(net1474));
 sg13g2_dlygate4sd3_1 hold412 (.A(\u_inv.input_reg[242] ),
    .X(net1475));
 sg13g2_dlygate4sd3_1 hold413 (.A(_00149_),
    .X(net1476));
 sg13g2_dlygate4sd3_1 hold414 (.A(\u_inv.input_reg[49] ),
    .X(net1477));
 sg13g2_dlygate4sd3_1 hold415 (.A(_01855_),
    .X(net1478));
 sg13g2_dlygate4sd3_1 hold416 (.A(\inv_result[157] ),
    .X(net1479));
 sg13g2_dlygate4sd3_1 hold418 (.A(\u_inv.input_reg[208] ),
    .X(net1481));
 sg13g2_dlygate4sd3_1 hold419 (.A(_00115_),
    .X(net1482));
 sg13g2_dlygate4sd3_1 hold420 (.A(\u_inv.d_next[187] ),
    .X(net1483));
 sg13g2_dlygate4sd3_1 hold421 (.A(_01437_),
    .X(net1484));
 sg13g2_dlygate4sd3_1 hold422 (.A(\inv_result[15] ),
    .X(net1485));
 sg13g2_dlygate4sd3_1 hold423 (.A(\u_inv.f_reg[34] ),
    .X(net1486));
 sg13g2_dlygate4sd3_1 hold424 (.A(_01541_),
    .X(net1487));
 sg13g2_dlygate4sd3_1 hold425 (.A(\inv_result[2] ),
    .X(net1488));
 sg13g2_dlygate4sd3_1 hold426 (.A(_00996_),
    .X(net1489));
 sg13g2_dlygate4sd3_1 hold427 (.A(\u_inv.input_reg[51] ),
    .X(net1490));
 sg13g2_dlygate4sd3_1 hold428 (.A(_01857_),
    .X(net1491));
 sg13g2_dlygate4sd3_1 hold429 (.A(\u_inv.input_reg[50] ),
    .X(net1492));
 sg13g2_dlygate4sd3_1 hold430 (.A(_01856_),
    .X(net1493));
 sg13g2_dlygate4sd3_1 hold431 (.A(\shift_reg[8] ),
    .X(net1494));
 sg13g2_dlygate4sd3_1 hold432 (.A(_00183_),
    .X(net1495));
 sg13g2_dlygate4sd3_1 hold433 (.A(\u_inv.d_next[163] ),
    .X(net1496));
 sg13g2_dlygate4sd3_1 hold434 (.A(_01413_),
    .X(net1497));
 sg13g2_dlygate4sd3_1 hold435 (.A(\u_inv.input_reg[152] ),
    .X(net1498));
 sg13g2_dlygate4sd3_1 hold436 (.A(_00059_),
    .X(net1499));
 sg13g2_dlygate4sd3_1 hold437 (.A(\u_inv.input_reg[31] ),
    .X(net1500));
 sg13g2_dlygate4sd3_1 hold438 (.A(_01837_),
    .X(net1501));
 sg13g2_dlygate4sd3_1 hold439 (.A(\u_inv.input_reg[158] ),
    .X(net1502));
 sg13g2_dlygate4sd3_1 hold440 (.A(_00065_),
    .X(net1503));
 sg13g2_dlygate4sd3_1 hold441 (.A(\u_inv.f_reg[145] ),
    .X(net1504));
 sg13g2_dlygate4sd3_1 hold442 (.A(\inv_result[229] ),
    .X(net1505));
 sg13g2_dlygate4sd3_1 hold443 (.A(\u_inv.f_reg[48] ),
    .X(net1506));
 sg13g2_dlygate4sd3_1 hold444 (.A(_01555_),
    .X(net1507));
 sg13g2_dlygate4sd3_1 hold445 (.A(\inv_result[255] ),
    .X(net1508));
 sg13g2_dlygate4sd3_1 hold446 (.A(\u_inv.input_reg[22] ),
    .X(net1509));
 sg13g2_dlygate4sd3_1 hold447 (.A(_01828_),
    .X(net1510));
 sg13g2_dlygate4sd3_1 hold448 (.A(\u_inv.f_next[165] ),
    .X(net1511));
 sg13g2_dlygate4sd3_1 hold449 (.A(_00625_),
    .X(net1512));
 sg13g2_dlygate4sd3_1 hold450 (.A(\inv_result[16] ),
    .X(net1513));
 sg13g2_dlygate4sd3_1 hold451 (.A(\u_inv.input_reg[234] ),
    .X(net1514));
 sg13g2_dlygate4sd3_1 hold452 (.A(_00141_),
    .X(net1515));
 sg13g2_dlygate4sd3_1 hold453 (.A(\u_inv.input_reg[167] ),
    .X(net1516));
 sg13g2_dlygate4sd3_1 hold454 (.A(_00074_),
    .X(net1517));
 sg13g2_dlygate4sd3_1 hold455 (.A(\inv_result[230] ),
    .X(net1518));
 sg13g2_dlygate4sd3_1 hold456 (.A(\u_inv.input_reg[171] ),
    .X(net1519));
 sg13g2_dlygate4sd3_1 hold457 (.A(_00078_),
    .X(net1520));
 sg13g2_dlygate4sd3_1 hold458 (.A(\shift_reg[2] ),
    .X(net1521));
 sg13g2_dlygate4sd3_1 hold459 (.A(_00177_),
    .X(net1522));
 sg13g2_dlygate4sd3_1 hold460 (.A(\u_inv.input_reg[47] ),
    .X(net1523));
 sg13g2_dlygate4sd3_1 hold461 (.A(_01853_),
    .X(net1524));
 sg13g2_dlygate4sd3_1 hold462 (.A(\inv_result[35] ),
    .X(net1525));
 sg13g2_dlygate4sd3_1 hold463 (.A(\u_inv.input_reg[91] ),
    .X(net1526));
 sg13g2_dlygate4sd3_1 hold464 (.A(_01897_),
    .X(net1527));
 sg13g2_dlygate4sd3_1 hold465 (.A(\u_inv.input_reg[210] ),
    .X(net1528));
 sg13g2_dlygate4sd3_1 hold466 (.A(_00117_),
    .X(net1529));
 sg13g2_dlygate4sd3_1 hold467 (.A(\inv_result[176] ),
    .X(net1530));
 sg13g2_dlygate4sd3_1 hold468 (.A(\u_inv.input_reg[133] ),
    .X(net1531));
 sg13g2_dlygate4sd3_1 hold469 (.A(_00040_),
    .X(net1532));
 sg13g2_dlygate4sd3_1 hold470 (.A(\u_inv.input_reg[92] ),
    .X(net1533));
 sg13g2_dlygate4sd3_1 hold471 (.A(_01898_),
    .X(net1534));
 sg13g2_dlygate4sd3_1 hold472 (.A(\u_inv.input_reg[113] ),
    .X(net1535));
 sg13g2_dlygate4sd3_1 hold473 (.A(_00020_),
    .X(net1536));
 sg13g2_dlygate4sd3_1 hold474 (.A(\u_inv.input_reg[2] ),
    .X(net1537));
 sg13g2_dlygate4sd3_1 hold475 (.A(_01808_),
    .X(net1538));
 sg13g2_dlygate4sd3_1 hold476 (.A(\u_inv.d_next[165] ),
    .X(net1539));
 sg13g2_dlygate4sd3_1 hold477 (.A(_01415_),
    .X(net1540));
 sg13g2_dlygate4sd3_1 hold478 (.A(\u_inv.input_reg[52] ),
    .X(net1541));
 sg13g2_dlygate4sd3_1 hold479 (.A(_01858_),
    .X(net1542));
 sg13g2_dlygate4sd3_1 hold480 (.A(\inv_result[217] ),
    .X(net1543));
 sg13g2_dlygate4sd3_1 hold481 (.A(\u_inv.input_reg[180] ),
    .X(net1544));
 sg13g2_dlygate4sd3_1 hold482 (.A(_00087_),
    .X(net1545));
 sg13g2_dlygate4sd3_1 hold483 (.A(\u_inv.input_reg[96] ),
    .X(net1546));
 sg13g2_dlygate4sd3_1 hold484 (.A(_00003_),
    .X(net1547));
 sg13g2_dlygate4sd3_1 hold485 (.A(\inv_result[33] ),
    .X(net1548));
 sg13g2_dlygate4sd3_1 hold486 (.A(\u_inv.f_reg[8] ),
    .X(net1549));
 sg13g2_dlygate4sd3_1 hold487 (.A(_01515_),
    .X(net1550));
 sg13g2_dlygate4sd3_1 hold488 (.A(\u_inv.input_reg[176] ),
    .X(net1551));
 sg13g2_dlygate4sd3_1 hold489 (.A(_00083_),
    .X(net1552));
 sg13g2_dlygate4sd3_1 hold490 (.A(\u_inv.input_reg[79] ),
    .X(net1553));
 sg13g2_dlygate4sd3_1 hold491 (.A(_01885_),
    .X(net1554));
 sg13g2_dlygate4sd3_1 hold492 (.A(\u_inv.input_reg[153] ),
    .X(net1555));
 sg13g2_dlygate4sd3_1 hold493 (.A(_00060_),
    .X(net1556));
 sg13g2_dlygate4sd3_1 hold494 (.A(\u_inv.input_reg[25] ),
    .X(net1557));
 sg13g2_dlygate4sd3_1 hold495 (.A(_01831_),
    .X(net1558));
 sg13g2_dlygate4sd3_1 hold496 (.A(\u_inv.input_reg[228] ),
    .X(net1559));
 sg13g2_dlygate4sd3_1 hold497 (.A(_00135_),
    .X(net1560));
 sg13g2_dlygate4sd3_1 hold498 (.A(\u_inv.input_reg[161] ),
    .X(net1561));
 sg13g2_dlygate4sd3_1 hold499 (.A(_00068_),
    .X(net1562));
 sg13g2_dlygate4sd3_1 hold500 (.A(\inv_result[36] ),
    .X(net1563));
 sg13g2_dlygate4sd3_1 hold501 (.A(\u_inv.input_reg[245] ),
    .X(net1564));
 sg13g2_dlygate4sd3_1 hold502 (.A(_00152_),
    .X(net1565));
 sg13g2_dlygate4sd3_1 hold503 (.A(\inv_result[90] ),
    .X(net1566));
 sg13g2_dlygate4sd3_1 hold504 (.A(\u_inv.input_reg[6] ),
    .X(net1567));
 sg13g2_dlygate4sd3_1 hold505 (.A(_01812_),
    .X(net1568));
 sg13g2_dlygate4sd3_1 hold506 (.A(\inv_result[126] ),
    .X(net1569));
 sg13g2_dlygate4sd3_1 hold507 (.A(\u_inv.input_reg[177] ),
    .X(net1570));
 sg13g2_dlygate4sd3_1 hold508 (.A(_00084_),
    .X(net1571));
 sg13g2_dlygate4sd3_1 hold509 (.A(\u_inv.input_reg[58] ),
    .X(net1572));
 sg13g2_dlygate4sd3_1 hold510 (.A(_01864_),
    .X(net1573));
 sg13g2_dlygate4sd3_1 hold511 (.A(\shift_reg[3] ),
    .X(net1574));
 sg13g2_dlygate4sd3_1 hold512 (.A(_00178_),
    .X(net1575));
 sg13g2_dlygate4sd3_1 hold513 (.A(\u_inv.f_next[87] ),
    .X(net1576));
 sg13g2_dlygate4sd3_1 hold514 (.A(\u_inv.f_reg[224] ),
    .X(net1577));
 sg13g2_dlygate4sd3_1 hold515 (.A(_01731_),
    .X(net1578));
 sg13g2_dlygate4sd3_1 hold516 (.A(\u_inv.f_reg[36] ),
    .X(net1579));
 sg13g2_dlygate4sd3_1 hold517 (.A(_01543_),
    .X(net1580));
 sg13g2_dlygate4sd3_1 hold518 (.A(\u_inv.input_reg[179] ),
    .X(net1581));
 sg13g2_dlygate4sd3_1 hold519 (.A(_00086_),
    .X(net1582));
 sg13g2_dlygate4sd3_1 hold520 (.A(\inv_result[150] ),
    .X(net1583));
 sg13g2_dlygate4sd3_1 hold521 (.A(\u_inv.input_reg[71] ),
    .X(net1584));
 sg13g2_dlygate4sd3_1 hold522 (.A(_01877_),
    .X(net1585));
 sg13g2_dlygate4sd3_1 hold523 (.A(\u_inv.f_reg[72] ),
    .X(net1586));
 sg13g2_dlygate4sd3_1 hold524 (.A(_01579_),
    .X(net1587));
 sg13g2_dlygate4sd3_1 hold525 (.A(\u_inv.f_reg[26] ),
    .X(net1588));
 sg13g2_dlygate4sd3_1 hold526 (.A(_01533_),
    .X(net1589));
 sg13g2_dlygate4sd3_1 hold527 (.A(\u_inv.input_reg[40] ),
    .X(net1590));
 sg13g2_dlygate4sd3_1 hold528 (.A(_01846_),
    .X(net1591));
 sg13g2_dlygate4sd3_1 hold529 (.A(\u_inv.input_reg[110] ),
    .X(net1592));
 sg13g2_dlygate4sd3_1 hold530 (.A(_00017_),
    .X(net1593));
 sg13g2_dlygate4sd3_1 hold531 (.A(\u_inv.input_reg[61] ),
    .X(net1594));
 sg13g2_dlygate4sd3_1 hold532 (.A(_01867_),
    .X(net1595));
 sg13g2_dlygate4sd3_1 hold533 (.A(\inv_result[38] ),
    .X(net1596));
 sg13g2_dlygate4sd3_1 hold534 (.A(\u_inv.input_reg[57] ),
    .X(net1597));
 sg13g2_dlygate4sd3_1 hold535 (.A(_01863_),
    .X(net1598));
 sg13g2_dlygate4sd3_1 hold536 (.A(\u_inv.input_reg[43] ),
    .X(net1599));
 sg13g2_dlygate4sd3_1 hold537 (.A(_01849_),
    .X(net1600));
 sg13g2_dlygate4sd3_1 hold538 (.A(\u_inv.input_reg[66] ),
    .X(net1601));
 sg13g2_dlygate4sd3_1 hold539 (.A(_01872_),
    .X(net1602));
 sg13g2_dlygate4sd3_1 hold540 (.A(\inv_result[115] ),
    .X(net1603));
 sg13g2_dlygate4sd3_1 hold541 (.A(\u_inv.input_reg[238] ),
    .X(net1604));
 sg13g2_dlygate4sd3_1 hold542 (.A(_00145_),
    .X(net1605));
 sg13g2_dlygate4sd3_1 hold543 (.A(\inv_result[222] ),
    .X(net1606));
 sg13g2_dlygate4sd3_1 hold544 (.A(\inv_result[108] ),
    .X(net1607));
 sg13g2_dlygate4sd3_1 hold545 (.A(\u_inv.input_reg[94] ),
    .X(net1608));
 sg13g2_dlygate4sd3_1 hold546 (.A(_01900_),
    .X(net1609));
 sg13g2_dlygate4sd3_1 hold547 (.A(\u_inv.input_reg[229] ),
    .X(net1610));
 sg13g2_dlygate4sd3_1 hold548 (.A(_00136_),
    .X(net1611));
 sg13g2_dlygate4sd3_1 hold549 (.A(\u_inv.input_reg[15] ),
    .X(net1612));
 sg13g2_dlygate4sd3_1 hold550 (.A(_01821_),
    .X(net1613));
 sg13g2_dlygate4sd3_1 hold551 (.A(\u_inv.input_reg[86] ),
    .X(net1614));
 sg13g2_dlygate4sd3_1 hold552 (.A(_01892_),
    .X(net1615));
 sg13g2_dlygate4sd3_1 hold553 (.A(\u_inv.input_reg[64] ),
    .X(net1616));
 sg13g2_dlygate4sd3_1 hold554 (.A(_01870_),
    .X(net1617));
 sg13g2_dlygate4sd3_1 hold555 (.A(\u_inv.counter[3] ),
    .X(net1618));
 sg13g2_dlygate4sd3_1 hold556 (.A(_01799_),
    .X(net1619));
 sg13g2_dlygate4sd3_1 hold557 (.A(\inv_result[142] ),
    .X(net1620));
 sg13g2_dlygate4sd3_1 hold558 (.A(\u_inv.f_reg[138] ),
    .X(net1621));
 sg13g2_dlygate4sd3_1 hold559 (.A(_01645_),
    .X(net1622));
 sg13g2_dlygate4sd3_1 hold560 (.A(\u_inv.f_reg[130] ),
    .X(net1623));
 sg13g2_dlygate4sd3_1 hold561 (.A(_01637_),
    .X(net1624));
 sg13g2_dlygate4sd3_1 hold562 (.A(\u_inv.input_reg[216] ),
    .X(net1625));
 sg13g2_dlygate4sd3_1 hold563 (.A(_00123_),
    .X(net1626));
 sg13g2_dlygate4sd3_1 hold564 (.A(\inv_result[78] ),
    .X(net1627));
 sg13g2_dlygate4sd3_1 hold565 (.A(\u_inv.input_reg[215] ),
    .X(net1628));
 sg13g2_dlygate4sd3_1 hold566 (.A(_00122_),
    .X(net1629));
 sg13g2_dlygate4sd3_1 hold567 (.A(\u_inv.input_reg[174] ),
    .X(net1630));
 sg13g2_dlygate4sd3_1 hold568 (.A(_00081_),
    .X(net1631));
 sg13g2_dlygate4sd3_1 hold569 (.A(\u_inv.f_reg[92] ),
    .X(net1632));
 sg13g2_dlygate4sd3_1 hold570 (.A(_01599_),
    .X(net1633));
 sg13g2_dlygate4sd3_1 hold571 (.A(\u_inv.f_reg[156] ),
    .X(net1634));
 sg13g2_dlygate4sd3_1 hold572 (.A(_01663_),
    .X(net1635));
 sg13g2_dlygate4sd3_1 hold573 (.A(\u_inv.f_reg[6] ),
    .X(net1636));
 sg13g2_dlygate4sd3_1 hold574 (.A(_01513_),
    .X(net1637));
 sg13g2_dlygate4sd3_1 hold575 (.A(\u_inv.d_next[91] ),
    .X(net1638));
 sg13g2_dlygate4sd3_1 hold576 (.A(_01341_),
    .X(net1639));
 sg13g2_dlygate4sd3_1 hold577 (.A(\u_inv.input_reg[129] ),
    .X(net1640));
 sg13g2_dlygate4sd3_1 hold578 (.A(_00036_),
    .X(net1641));
 sg13g2_dlygate4sd3_1 hold579 (.A(\u_inv.f_reg[104] ),
    .X(net1642));
 sg13g2_dlygate4sd3_1 hold580 (.A(_01611_),
    .X(net1643));
 sg13g2_dlygate4sd3_1 hold581 (.A(\inv_result[250] ),
    .X(net1644));
 sg13g2_dlygate4sd3_1 hold582 (.A(\inv_result[94] ),
    .X(net1645));
 sg13g2_dlygate4sd3_1 hold583 (.A(\u_inv.f_reg[16] ),
    .X(net1646));
 sg13g2_dlygate4sd3_1 hold584 (.A(_01523_),
    .X(net1647));
 sg13g2_dlygate4sd3_1 hold585 (.A(\u_inv.input_reg[3] ),
    .X(net1648));
 sg13g2_dlygate4sd3_1 hold586 (.A(_01809_),
    .X(net1649));
 sg13g2_dlygate4sd3_1 hold587 (.A(\u_inv.f_reg[184] ),
    .X(net1650));
 sg13g2_dlygate4sd3_1 hold588 (.A(_01691_),
    .X(net1651));
 sg13g2_dlygate4sd3_1 hold589 (.A(\u_inv.input_reg[227] ),
    .X(net1652));
 sg13g2_dlygate4sd3_1 hold590 (.A(_00134_),
    .X(net1653));
 sg13g2_dlygate4sd3_1 hold591 (.A(\u_inv.f_reg[38] ),
    .X(net1654));
 sg13g2_dlygate4sd3_1 hold592 (.A(_01545_),
    .X(net1655));
 sg13g2_dlygate4sd3_1 hold593 (.A(\u_inv.input_reg[122] ),
    .X(net1656));
 sg13g2_dlygate4sd3_1 hold594 (.A(_00029_),
    .X(net1657));
 sg13g2_dlygate4sd3_1 hold595 (.A(\u_inv.input_reg[98] ),
    .X(net1658));
 sg13g2_dlygate4sd3_1 hold596 (.A(_00005_),
    .X(net1659));
 sg13g2_dlygate4sd3_1 hold597 (.A(\u_inv.input_reg[202] ),
    .X(net1660));
 sg13g2_dlygate4sd3_1 hold598 (.A(_00109_),
    .X(net1661));
 sg13g2_dlygate4sd3_1 hold599 (.A(\inv_result[178] ),
    .X(net1662));
 sg13g2_dlygate4sd3_1 hold600 (.A(\inv_result[223] ),
    .X(net1663));
 sg13g2_dlygate4sd3_1 hold601 (.A(\inv_result[227] ),
    .X(net1664));
 sg13g2_dlygate4sd3_1 hold602 (.A(\u_inv.f_reg[77] ),
    .X(net1665));
 sg13g2_dlygate4sd3_1 hold603 (.A(_01584_),
    .X(net1666));
 sg13g2_dlygate4sd3_1 hold604 (.A(\u_inv.f_reg[146] ),
    .X(net1667));
 sg13g2_dlygate4sd3_1 hold605 (.A(_01653_),
    .X(net1668));
 sg13g2_dlygate4sd3_1 hold606 (.A(\u_inv.f_next[49] ),
    .X(net1669));
 sg13g2_dlygate4sd3_1 hold607 (.A(\u_inv.input_reg[60] ),
    .X(net1670));
 sg13g2_dlygate4sd3_1 hold608 (.A(_01866_),
    .X(net1671));
 sg13g2_dlygate4sd3_1 hold609 (.A(\u_inv.delta_reg[4] ),
    .X(net1672));
 sg13g2_dlygate4sd3_1 hold610 (.A(\inv_result[130] ),
    .X(net1673));
 sg13g2_dlygate4sd3_1 hold611 (.A(\inv_result[195] ),
    .X(net1674));
 sg13g2_dlygate4sd3_1 hold612 (.A(\u_inv.input_reg[75] ),
    .X(net1675));
 sg13g2_dlygate4sd3_1 hold613 (.A(_01881_),
    .X(net1676));
 sg13g2_dlygate4sd3_1 hold614 (.A(\inv_result[183] ),
    .X(net1677));
 sg13g2_dlygate4sd3_1 hold615 (.A(pipe_pending),
    .X(net1678));
 sg13g2_dlygate4sd3_1 hold616 (.A(_19804_),
    .X(net1679));
 sg13g2_dlygate4sd3_1 hold617 (.A(\u_inv.d_next[1] ),
    .X(net1680));
 sg13g2_dlygate4sd3_1 hold618 (.A(\inv_result[239] ),
    .X(net1681));
 sg13g2_dlygate4sd3_1 hold619 (.A(\u_inv.input_reg[104] ),
    .X(net1682));
 sg13g2_dlygate4sd3_1 hold620 (.A(_00011_),
    .X(net1683));
 sg13g2_dlygate4sd3_1 hold621 (.A(\u_inv.f_next[11] ),
    .X(net1684));
 sg13g2_dlygate4sd3_1 hold622 (.A(\u_inv.input_reg[134] ),
    .X(net1685));
 sg13g2_dlygate4sd3_1 hold623 (.A(_00041_),
    .X(net1686));
 sg13g2_dlygate4sd3_1 hold624 (.A(\u_inv.f_reg[60] ),
    .X(net1687));
 sg13g2_dlygate4sd3_1 hold625 (.A(_01567_),
    .X(net1688));
 sg13g2_dlygate4sd3_1 hold626 (.A(\u_inv.input_reg[108] ),
    .X(net1689));
 sg13g2_dlygate4sd3_1 hold627 (.A(_00015_),
    .X(net1690));
 sg13g2_dlygate4sd3_1 hold628 (.A(\u_inv.f_next[243] ),
    .X(net1691));
 sg13g2_dlygate4sd3_1 hold629 (.A(\u_inv.input_reg[21] ),
    .X(net1692));
 sg13g2_dlygate4sd3_1 hold630 (.A(_01827_),
    .X(net1693));
 sg13g2_dlygate4sd3_1 hold631 (.A(\u_inv.input_reg[13] ),
    .X(net1694));
 sg13g2_dlygate4sd3_1 hold632 (.A(_01819_),
    .X(net1695));
 sg13g2_dlygate4sd3_1 hold633 (.A(\u_inv.f_reg[12] ),
    .X(net1696));
 sg13g2_dlygate4sd3_1 hold634 (.A(_01519_),
    .X(net1697));
 sg13g2_dlygate4sd3_1 hold635 (.A(\inv_result[54] ),
    .X(net1698));
 sg13g2_dlygate4sd3_1 hold636 (.A(\u_inv.input_reg[212] ),
    .X(net1699));
 sg13g2_dlygate4sd3_1 hold637 (.A(_00119_),
    .X(net1700));
 sg13g2_dlygate4sd3_1 hold638 (.A(\u_inv.d_next[100] ),
    .X(net1701));
 sg13g2_dlygate4sd3_1 hold639 (.A(_01350_),
    .X(net1702));
 sg13g2_dlygate4sd3_1 hold640 (.A(\inv_result[146] ),
    .X(net1703));
 sg13g2_dlygate4sd3_1 hold641 (.A(\u_inv.input_reg[196] ),
    .X(net1704));
 sg13g2_dlygate4sd3_1 hold642 (.A(_00103_),
    .X(net1705));
 sg13g2_dlygate4sd3_1 hold643 (.A(\u_inv.input_reg[244] ),
    .X(net1706));
 sg13g2_dlygate4sd3_1 hold644 (.A(_00151_),
    .X(net1707));
 sg13g2_dlygate4sd3_1 hold645 (.A(\u_inv.f_reg[30] ),
    .X(net1708));
 sg13g2_dlygate4sd3_1 hold646 (.A(_01537_),
    .X(net1709));
 sg13g2_dlygate4sd3_1 hold647 (.A(\inv_result[181] ),
    .X(net1710));
 sg13g2_dlygate4sd3_1 hold648 (.A(\u_inv.f_reg[83] ),
    .X(net1711));
 sg13g2_dlygate4sd3_1 hold649 (.A(_01590_),
    .X(net1712));
 sg13g2_dlygate4sd3_1 hold650 (.A(\u_inv.input_reg[194] ),
    .X(net1713));
 sg13g2_dlygate4sd3_1 hold651 (.A(_00101_),
    .X(net1714));
 sg13g2_dlygate4sd3_1 hold652 (.A(\u_inv.input_reg[248] ),
    .X(net1715));
 sg13g2_dlygate4sd3_1 hold653 (.A(_00155_),
    .X(net1716));
 sg13g2_dlygate4sd3_1 hold654 (.A(\u_inv.f_reg[17] ),
    .X(net1717));
 sg13g2_dlygate4sd3_1 hold655 (.A(_01524_),
    .X(net1718));
 sg13g2_dlygate4sd3_1 hold656 (.A(\u_inv.input_reg[90] ),
    .X(net1719));
 sg13g2_dlygate4sd3_1 hold657 (.A(_01896_),
    .X(net1720));
 sg13g2_dlygate4sd3_1 hold658 (.A(\inv_result[99] ),
    .X(net1721));
 sg13g2_dlygate4sd3_1 hold659 (.A(\u_inv.f_reg[3] ),
    .X(net1722));
 sg13g2_dlygate4sd3_1 hold660 (.A(_01510_),
    .X(net1723));
 sg13g2_dlygate4sd3_1 hold661 (.A(\u_inv.d_next[42] ),
    .X(net1724));
 sg13g2_dlygate4sd3_1 hold662 (.A(_01292_),
    .X(net1725));
 sg13g2_dlygate4sd3_1 hold663 (.A(\u_inv.f_next[219] ),
    .X(net1726));
 sg13g2_dlygate4sd3_1 hold664 (.A(_00679_),
    .X(net1727));
 sg13g2_dlygate4sd3_1 hold665 (.A(\u_inv.input_reg[118] ),
    .X(net1728));
 sg13g2_dlygate4sd3_1 hold666 (.A(_00025_),
    .X(net1729));
 sg13g2_dlygate4sd3_1 hold667 (.A(\shift_reg[0] ),
    .X(net1730));
 sg13g2_dlygate4sd3_1 hold668 (.A(_00175_),
    .X(net1731));
 sg13g2_dlygate4sd3_1 hold669 (.A(\inv_result[26] ),
    .X(net1732));
 sg13g2_dlygate4sd3_1 hold670 (.A(\u_inv.input_reg[111] ),
    .X(net1733));
 sg13g2_dlygate4sd3_1 hold671 (.A(_00018_),
    .X(net1734));
 sg13g2_dlygate4sd3_1 hold672 (.A(\inv_cycles[8] ),
    .X(net1735));
 sg13g2_dlygate4sd3_1 hold673 (.A(_01795_),
    .X(net1736));
 sg13g2_dlygate4sd3_1 hold674 (.A(\u_inv.input_reg[65] ),
    .X(net1737));
 sg13g2_dlygate4sd3_1 hold675 (.A(_01871_),
    .X(net1738));
 sg13g2_dlygate4sd3_1 hold676 (.A(\u_inv.f_reg[121] ),
    .X(net1739));
 sg13g2_dlygate4sd3_1 hold677 (.A(_01628_),
    .X(net1740));
 sg13g2_dlygate4sd3_1 hold678 (.A(\inv_result[138] ),
    .X(net1741));
 sg13g2_dlygate4sd3_1 hold679 (.A(\u_inv.d_next[31] ),
    .X(net1742));
 sg13g2_dlygate4sd3_1 hold680 (.A(_01281_),
    .X(net1743));
 sg13g2_dlygate4sd3_1 hold681 (.A(\u_inv.input_reg[30] ),
    .X(net1744));
 sg13g2_dlygate4sd3_1 hold682 (.A(_01836_),
    .X(net1745));
 sg13g2_dlygate4sd3_1 hold683 (.A(\u_inv.f_reg[226] ),
    .X(net1746));
 sg13g2_dlygate4sd3_1 hold684 (.A(_01733_),
    .X(net1747));
 sg13g2_dlygate4sd3_1 hold685 (.A(\u_inv.input_reg[114] ),
    .X(net1748));
 sg13g2_dlygate4sd3_1 hold686 (.A(_00021_),
    .X(net1749));
 sg13g2_dlygate4sd3_1 hold687 (.A(\u_inv.f_reg[20] ),
    .X(net1750));
 sg13g2_dlygate4sd3_1 hold688 (.A(_01527_),
    .X(net1751));
 sg13g2_dlygate4sd3_1 hold689 (.A(\inv_result[103] ),
    .X(net1752));
 sg13g2_dlygate4sd3_1 hold690 (.A(\u_inv.f_next[4] ),
    .X(net1753));
 sg13g2_dlygate4sd3_1 hold691 (.A(_01511_),
    .X(net1754));
 sg13g2_dlygate4sd3_1 hold692 (.A(\u_inv.input_reg[42] ),
    .X(net1755));
 sg13g2_dlygate4sd3_1 hold693 (.A(_01848_),
    .X(net1756));
 sg13g2_dlygate4sd3_1 hold694 (.A(\u_inv.input_reg[67] ),
    .X(net1757));
 sg13g2_dlygate4sd3_1 hold695 (.A(_01873_),
    .X(net1758));
 sg13g2_dlygate4sd3_1 hold696 (.A(\inv_result[154] ),
    .X(net1759));
 sg13g2_dlygate4sd3_1 hold697 (.A(\u_inv.input_reg[7] ),
    .X(net1760));
 sg13g2_dlygate4sd3_1 hold698 (.A(_01813_),
    .X(net1761));
 sg13g2_dlygate4sd3_1 hold699 (.A(\u_inv.input_reg[109] ),
    .X(net1762));
 sg13g2_dlygate4sd3_1 hold700 (.A(_00016_),
    .X(net1763));
 sg13g2_dlygate4sd3_1 hold701 (.A(\shift_reg[45] ),
    .X(net1764));
 sg13g2_dlygate4sd3_1 hold702 (.A(_00220_),
    .X(net1765));
 sg13g2_dlygate4sd3_1 hold703 (.A(\inv_cycles[7] ),
    .X(net1766));
 sg13g2_dlygate4sd3_1 hold704 (.A(_01794_),
    .X(net1767));
 sg13g2_dlygate4sd3_1 hold705 (.A(\u_inv.state[1] ),
    .X(net1768));
 sg13g2_dlygate4sd3_1 hold706 (.A(_18623_),
    .X(net1769));
 sg13g2_dlygate4sd3_1 hold707 (.A(_00000_),
    .X(net1770));
 sg13g2_dlygate4sd3_1 hold708 (.A(\u_inv.input_reg[82] ),
    .X(net1771));
 sg13g2_dlygate4sd3_1 hold709 (.A(_01888_),
    .X(net1772));
 sg13g2_dlygate4sd3_1 hold710 (.A(\u_inv.f_reg[205] ),
    .X(net1773));
 sg13g2_dlygate4sd3_1 hold711 (.A(_01712_),
    .X(net1774));
 sg13g2_dlygate4sd3_1 hold712 (.A(\u_inv.input_reg[254] ),
    .X(net1775));
 sg13g2_dlygate4sd3_1 hold713 (.A(_00161_),
    .X(net1776));
 sg13g2_dlygate4sd3_1 hold714 (.A(\u_inv.f_reg[174] ),
    .X(net1777));
 sg13g2_dlygate4sd3_1 hold715 (.A(_01681_),
    .X(net1778));
 sg13g2_dlygate4sd3_1 hold716 (.A(\u_inv.f_next[60] ),
    .X(net1779));
 sg13g2_dlygate4sd3_1 hold717 (.A(\u_inv.input_reg[69] ),
    .X(net1780));
 sg13g2_dlygate4sd3_1 hold718 (.A(_01875_),
    .X(net1781));
 sg13g2_dlygate4sd3_1 hold719 (.A(\u_inv.d_next[174] ),
    .X(net1782));
 sg13g2_dlygate4sd3_1 hold720 (.A(\u_inv.input_reg[195] ),
    .X(net1783));
 sg13g2_dlygate4sd3_1 hold721 (.A(_00102_),
    .X(net1784));
 sg13g2_dlygate4sd3_1 hold722 (.A(\u_inv.f_reg[55] ),
    .X(net1785));
 sg13g2_dlygate4sd3_1 hold723 (.A(_01562_),
    .X(net1786));
 sg13g2_dlygate4sd3_1 hold724 (.A(\u_inv.f_reg[154] ),
    .X(net1787));
 sg13g2_dlygate4sd3_1 hold725 (.A(_01661_),
    .X(net1788));
 sg13g2_dlygate4sd3_1 hold726 (.A(\u_inv.f_reg[173] ),
    .X(net1789));
 sg13g2_dlygate4sd3_1 hold727 (.A(_01680_),
    .X(net1790));
 sg13g2_dlygate4sd3_1 hold728 (.A(\u_inv.input_reg[80] ),
    .X(net1791));
 sg13g2_dlygate4sd3_1 hold729 (.A(_01886_),
    .X(net1792));
 sg13g2_dlygate4sd3_1 hold730 (.A(\inv_result[11] ),
    .X(net1793));
 sg13g2_dlygate4sd3_1 hold731 (.A(\inv_result[210] ),
    .X(net1794));
 sg13g2_dlygate4sd3_1 hold732 (.A(\u_inv.input_reg[222] ),
    .X(net1795));
 sg13g2_dlygate4sd3_1 hold733 (.A(_00129_),
    .X(net1796));
 sg13g2_dlygate4sd3_1 hold734 (.A(\u_inv.input_reg[95] ),
    .X(net1797));
 sg13g2_dlygate4sd3_1 hold735 (.A(_00002_),
    .X(net1798));
 sg13g2_dlygate4sd3_1 hold736 (.A(\inv_result[135] ),
    .X(net1799));
 sg13g2_dlygate4sd3_1 hold737 (.A(\u_inv.input_reg[101] ),
    .X(net1800));
 sg13g2_dlygate4sd3_1 hold738 (.A(_00008_),
    .X(net1801));
 sg13g2_dlygate4sd3_1 hold739 (.A(\u_inv.input_reg[255] ),
    .X(net1802));
 sg13g2_dlygate4sd3_1 hold740 (.A(_00162_),
    .X(net1803));
 sg13g2_dlygate4sd3_1 hold741 (.A(\u_inv.input_reg[150] ),
    .X(net1804));
 sg13g2_dlygate4sd3_1 hold742 (.A(_00057_),
    .X(net1805));
 sg13g2_dlygate4sd3_1 hold743 (.A(\u_inv.input_reg[193] ),
    .X(net1806));
 sg13g2_dlygate4sd3_1 hold744 (.A(_00100_),
    .X(net1807));
 sg13g2_dlygate4sd3_1 hold745 (.A(\u_inv.input_reg[37] ),
    .X(net1808));
 sg13g2_dlygate4sd3_1 hold746 (.A(_01843_),
    .X(net1809));
 sg13g2_dlygate4sd3_1 hold747 (.A(\u_inv.f_reg[202] ),
    .X(net1810));
 sg13g2_dlygate4sd3_1 hold748 (.A(_01709_),
    .X(net1811));
 sg13g2_dlygate4sd3_1 hold749 (.A(\u_inv.input_reg[184] ),
    .X(net1812));
 sg13g2_dlygate4sd3_1 hold750 (.A(_00091_),
    .X(net1813));
 sg13g2_dlygate4sd3_1 hold751 (.A(\shift_reg[11] ),
    .X(net1814));
 sg13g2_dlygate4sd3_1 hold752 (.A(\u_inv.input_reg[81] ),
    .X(net1815));
 sg13g2_dlygate4sd3_1 hold753 (.A(_01887_),
    .X(net1816));
 sg13g2_dlygate4sd3_1 hold754 (.A(\u_inv.input_reg[185] ),
    .X(net1817));
 sg13g2_dlygate4sd3_1 hold755 (.A(_00092_),
    .X(net1818));
 sg13g2_dlygate4sd3_1 hold756 (.A(\inv_result[166] ),
    .X(net1819));
 sg13g2_dlygate4sd3_1 hold757 (.A(\u_inv.f_reg[150] ),
    .X(net1820));
 sg13g2_dlygate4sd3_1 hold758 (.A(_01657_),
    .X(net1821));
 sg13g2_dlygate4sd3_1 hold759 (.A(\inv_result[52] ),
    .X(net1822));
 sg13g2_dlygate4sd3_1 hold760 (.A(\u_inv.d_next[8] ),
    .X(net1823));
 sg13g2_dlygate4sd3_1 hold761 (.A(_01258_),
    .X(net1824));
 sg13g2_dlygate4sd3_1 hold762 (.A(\u_inv.input_reg[62] ),
    .X(net1825));
 sg13g2_dlygate4sd3_1 hold763 (.A(_01868_),
    .X(net1826));
 sg13g2_dlygate4sd3_1 hold764 (.A(\u_inv.input_reg[77] ),
    .X(net1827));
 sg13g2_dlygate4sd3_1 hold765 (.A(_01883_),
    .X(net1828));
 sg13g2_dlygate4sd3_1 hold766 (.A(\u_inv.input_reg[70] ),
    .X(net1829));
 sg13g2_dlygate4sd3_1 hold767 (.A(_01876_),
    .X(net1830));
 sg13g2_dlygate4sd3_1 hold768 (.A(\u_inv.f_reg[14] ),
    .X(net1831));
 sg13g2_dlygate4sd3_1 hold769 (.A(_01521_),
    .X(net1832));
 sg13g2_dlygate4sd3_1 hold770 (.A(\u_inv.input_reg[197] ),
    .X(net1833));
 sg13g2_dlygate4sd3_1 hold771 (.A(_00104_),
    .X(net1834));
 sg13g2_dlygate4sd3_1 hold772 (.A(\u_inv.input_reg[182] ),
    .X(net1835));
 sg13g2_dlygate4sd3_1 hold773 (.A(_00089_),
    .X(net1836));
 sg13g2_dlygate4sd3_1 hold774 (.A(\inv_result[110] ),
    .X(net1837));
 sg13g2_dlygate4sd3_1 hold775 (.A(\u_inv.input_reg[225] ),
    .X(net1838));
 sg13g2_dlygate4sd3_1 hold776 (.A(_00132_),
    .X(net1839));
 sg13g2_dlygate4sd3_1 hold777 (.A(\byte_cnt[2] ),
    .X(net1840));
 sg13g2_dlygate4sd3_1 hold778 (.A(_18919_),
    .X(net1841));
 sg13g2_dlygate4sd3_1 hold779 (.A(\u_inv.f_reg[229] ),
    .X(net1842));
 sg13g2_dlygate4sd3_1 hold780 (.A(_01736_),
    .X(net1843));
 sg13g2_dlygate4sd3_1 hold781 (.A(\u_inv.f_reg[162] ),
    .X(net1844));
 sg13g2_dlygate4sd3_1 hold782 (.A(_01669_),
    .X(net1845));
 sg13g2_dlygate4sd3_1 hold783 (.A(\inv_result[158] ),
    .X(net1846));
 sg13g2_dlygate4sd3_1 hold784 (.A(\inv_result[136] ),
    .X(net1847));
 sg13g2_dlygate4sd3_1 hold785 (.A(\inv_result[12] ),
    .X(net1848));
 sg13g2_dlygate4sd3_1 hold786 (.A(\u_inv.d_next[77] ),
    .X(net1849));
 sg13g2_dlygate4sd3_1 hold787 (.A(_01327_),
    .X(net1850));
 sg13g2_dlygate4sd3_1 hold788 (.A(\shift_reg[239] ),
    .X(net1851));
 sg13g2_dlygate4sd3_1 hold789 (.A(_00414_),
    .X(net1852));
 sg13g2_dlygate4sd3_1 hold790 (.A(\inv_result[186] ),
    .X(net1853));
 sg13g2_dlygate4sd3_1 hold791 (.A(\u_inv.f_reg[107] ),
    .X(net1854));
 sg13g2_dlygate4sd3_1 hold792 (.A(_01614_),
    .X(net1855));
 sg13g2_dlygate4sd3_1 hold793 (.A(\inv_result[160] ),
    .X(net1856));
 sg13g2_dlygate4sd3_1 hold794 (.A(\u_inv.f_reg[64] ),
    .X(net1857));
 sg13g2_dlygate4sd3_1 hold795 (.A(_01571_),
    .X(net1858));
 sg13g2_dlygate4sd3_1 hold796 (.A(\inv_result[196] ),
    .X(net1859));
 sg13g2_dlygate4sd3_1 hold797 (.A(\u_inv.f_reg[144] ),
    .X(net1860));
 sg13g2_dlygate4sd3_1 hold798 (.A(_01651_),
    .X(net1861));
 sg13g2_dlygate4sd3_1 hold799 (.A(\inv_result[114] ),
    .X(net1862));
 sg13g2_dlygate4sd3_1 hold800 (.A(\u_inv.input_reg[102] ),
    .X(net1863));
 sg13g2_dlygate4sd3_1 hold801 (.A(_00009_),
    .X(net1864));
 sg13g2_dlygate4sd3_1 hold802 (.A(\u_inv.f_reg[59] ),
    .X(net1865));
 sg13g2_dlygate4sd3_1 hold803 (.A(_01566_),
    .X(net1866));
 sg13g2_dlygate4sd3_1 hold804 (.A(\u_inv.d_next[70] ),
    .X(net1867));
 sg13g2_dlygate4sd3_1 hold805 (.A(\u_inv.input_reg[221] ),
    .X(net1868));
 sg13g2_dlygate4sd3_1 hold806 (.A(_00128_),
    .X(net1869));
 sg13g2_dlygate4sd3_1 hold807 (.A(\u_inv.input_reg[16] ),
    .X(net1870));
 sg13g2_dlygate4sd3_1 hold808 (.A(_01822_),
    .X(net1871));
 sg13g2_dlygate4sd3_1 hold809 (.A(\u_inv.input_reg[188] ),
    .X(net1872));
 sg13g2_dlygate4sd3_1 hold810 (.A(_00095_),
    .X(net1873));
 sg13g2_dlygate4sd3_1 hold811 (.A(\u_inv.f_reg[110] ),
    .X(net1874));
 sg13g2_dlygate4sd3_1 hold812 (.A(_01617_),
    .X(net1875));
 sg13g2_dlygate4sd3_1 hold813 (.A(\u_inv.input_reg[45] ),
    .X(net1876));
 sg13g2_dlygate4sd3_1 hold814 (.A(_01851_),
    .X(net1877));
 sg13g2_dlygate4sd3_1 hold815 (.A(\inv_cycles[6] ),
    .X(net1878));
 sg13g2_dlygate4sd3_1 hold816 (.A(_01793_),
    .X(net1879));
 sg13g2_dlygate4sd3_1 hold817 (.A(\inv_result[242] ),
    .X(net1880));
 sg13g2_dlygate4sd3_1 hold818 (.A(\inv_result[132] ),
    .X(net1881));
 sg13g2_dlygate4sd3_1 hold819 (.A(\inv_result[180] ),
    .X(net1882));
 sg13g2_dlygate4sd3_1 hold820 (.A(\u_inv.input_reg[165] ),
    .X(net1883));
 sg13g2_dlygate4sd3_1 hold821 (.A(_00072_),
    .X(net1884));
 sg13g2_dlygate4sd3_1 hold822 (.A(\u_inv.input_reg[148] ),
    .X(net1885));
 sg13g2_dlygate4sd3_1 hold823 (.A(_00055_),
    .X(net1886));
 sg13g2_dlygate4sd3_1 hold824 (.A(\inv_result[175] ),
    .X(net1887));
 sg13g2_dlygate4sd3_1 hold825 (.A(\u_inv.input_reg[5] ),
    .X(net1888));
 sg13g2_dlygate4sd3_1 hold826 (.A(_01811_),
    .X(net1889));
 sg13g2_dlygate4sd3_1 hold827 (.A(\u_inv.input_reg[53] ),
    .X(net1890));
 sg13g2_dlygate4sd3_1 hold828 (.A(_01859_),
    .X(net1891));
 sg13g2_dlygate4sd3_1 hold829 (.A(\inv_result[169] ),
    .X(net1892));
 sg13g2_dlygate4sd3_1 hold830 (.A(\inv_result[124] ),
    .X(net1893));
 sg13g2_dlygate4sd3_1 hold831 (.A(\u_inv.f_reg[50] ),
    .X(net1894));
 sg13g2_dlygate4sd3_1 hold832 (.A(_01557_),
    .X(net1895));
 sg13g2_dlygate4sd3_1 hold833 (.A(\inv_result[31] ),
    .X(net1896));
 sg13g2_dlygate4sd3_1 hold834 (.A(\u_inv.f_reg[123] ),
    .X(net1897));
 sg13g2_dlygate4sd3_1 hold835 (.A(_01630_),
    .X(net1898));
 sg13g2_dlygate4sd3_1 hold836 (.A(\inv_result[218] ),
    .X(net1899));
 sg13g2_dlygate4sd3_1 hold837 (.A(\u_inv.f_reg[70] ),
    .X(net1900));
 sg13g2_dlygate4sd3_1 hold838 (.A(_01577_),
    .X(net1901));
 sg13g2_dlygate4sd3_1 hold839 (.A(\u_inv.d_next[149] ),
    .X(net1902));
 sg13g2_dlygate4sd3_1 hold840 (.A(_01399_),
    .X(net1903));
 sg13g2_dlygate4sd3_1 hold841 (.A(\inv_result[241] ),
    .X(net1904));
 sg13g2_dlygate4sd3_1 hold842 (.A(\inv_result[127] ),
    .X(net1905));
 sg13g2_dlygate4sd3_1 hold843 (.A(\u_inv.input_reg[127] ),
    .X(net1906));
 sg13g2_dlygate4sd3_1 hold844 (.A(_00034_),
    .X(net1907));
 sg13g2_dlygate4sd3_1 hold845 (.A(\u_inv.f_reg[119] ),
    .X(net1908));
 sg13g2_dlygate4sd3_1 hold846 (.A(_01626_),
    .X(net1909));
 sg13g2_dlygate4sd3_1 hold847 (.A(\inv_result[14] ),
    .X(net1910));
 sg13g2_dlygate4sd3_1 hold848 (.A(\u_inv.input_reg[140] ),
    .X(net1911));
 sg13g2_dlygate4sd3_1 hold849 (.A(_00047_),
    .X(net1912));
 sg13g2_dlygate4sd3_1 hold850 (.A(\u_inv.f_reg[246] ),
    .X(net1913));
 sg13g2_dlygate4sd3_1 hold851 (.A(_01753_),
    .X(net1914));
 sg13g2_dlygate4sd3_1 hold852 (.A(\u_inv.d_next[29] ),
    .X(net1915));
 sg13g2_dlygate4sd3_1 hold853 (.A(_01279_),
    .X(net1916));
 sg13g2_dlygate4sd3_1 hold854 (.A(\trng_data[5] ),
    .X(net1917));
 sg13g2_dlygate4sd3_1 hold855 (.A(_00455_),
    .X(net1918));
 sg13g2_dlygate4sd3_1 hold856 (.A(\inv_result[211] ),
    .X(net1919));
 sg13g2_dlygate4sd3_1 hold857 (.A(\u_inv.f_reg[27] ),
    .X(net1920));
 sg13g2_dlygate4sd3_1 hold858 (.A(_01534_),
    .X(net1921));
 sg13g2_dlygate4sd3_1 hold859 (.A(\inv_result[168] ),
    .X(net1922));
 sg13g2_dlygate4sd3_1 hold860 (.A(\inv_result[70] ),
    .X(net1923));
 sg13g2_dlygate4sd3_1 hold861 (.A(\u_inv.input_reg[1] ),
    .X(net1924));
 sg13g2_dlygate4sd3_1 hold862 (.A(_01807_),
    .X(net1925));
 sg13g2_dlygate4sd3_1 hold863 (.A(\u_inv.f_next[205] ),
    .X(net1926));
 sg13g2_dlygate4sd3_1 hold864 (.A(_00665_),
    .X(net1927));
 sg13g2_dlygate4sd3_1 hold865 (.A(\u_inv.input_reg[206] ),
    .X(net1928));
 sg13g2_dlygate4sd3_1 hold866 (.A(_00113_),
    .X(net1929));
 sg13g2_dlygate4sd3_1 hold867 (.A(\u_inv.input_reg[170] ),
    .X(net1930));
 sg13g2_dlygate4sd3_1 hold868 (.A(_00077_),
    .X(net1931));
 sg13g2_dlygate4sd3_1 hold869 (.A(\inv_result[202] ),
    .X(net1932));
 sg13g2_dlygate4sd3_1 hold870 (.A(\inv_result[240] ),
    .X(net1933));
 sg13g2_dlygate4sd3_1 hold871 (.A(\u_inv.input_reg[85] ),
    .X(net1934));
 sg13g2_dlygate4sd3_1 hold872 (.A(_01891_),
    .X(net1935));
 sg13g2_dlygate4sd3_1 hold873 (.A(\shift_reg[127] ),
    .X(net1936));
 sg13g2_dlygate4sd3_1 hold874 (.A(_00302_),
    .X(net1937));
 sg13g2_dlygate4sd3_1 hold875 (.A(\inv_result[184] ),
    .X(net1938));
 sg13g2_dlygate4sd3_1 hold877 (.A(\u_inv.f_reg[238] ),
    .X(net1940));
 sg13g2_dlygate4sd3_1 hold878 (.A(_01745_),
    .X(net1941));
 sg13g2_dlygate4sd3_1 hold879 (.A(\u_inv.input_reg[235] ),
    .X(net1942));
 sg13g2_dlygate4sd3_1 hold880 (.A(_00142_),
    .X(net1943));
 sg13g2_dlygate4sd3_1 hold881 (.A(\inv_result[111] ),
    .X(net1944));
 sg13g2_dlygate4sd3_1 hold882 (.A(\u_inv.input_reg[100] ),
    .X(net1945));
 sg13g2_dlygate4sd3_1 hold883 (.A(_00007_),
    .X(net1946));
 sg13g2_dlygate4sd3_1 hold884 (.A(\u_inv.f_reg[73] ),
    .X(net1947));
 sg13g2_dlygate4sd3_1 hold885 (.A(_01580_),
    .X(net1948));
 sg13g2_dlygate4sd3_1 hold886 (.A(\u_inv.f_reg[62] ),
    .X(net1949));
 sg13g2_dlygate4sd3_1 hold887 (.A(_01569_),
    .X(net1950));
 sg13g2_dlygate4sd3_1 hold888 (.A(\u_inv.input_reg[68] ),
    .X(net1951));
 sg13g2_dlygate4sd3_1 hold889 (.A(_01874_),
    .X(net1952));
 sg13g2_dlygate4sd3_1 hold890 (.A(\u_inv.f_reg[198] ),
    .X(net1953));
 sg13g2_dlygate4sd3_1 hold891 (.A(_01705_),
    .X(net1954));
 sg13g2_dlygate4sd3_1 hold892 (.A(\u_inv.d_next[34] ),
    .X(net1955));
 sg13g2_dlygate4sd3_1 hold893 (.A(_01284_),
    .X(net1956));
 sg13g2_dlygate4sd3_1 hold894 (.A(\u_inv.f_reg[188] ),
    .X(net1957));
 sg13g2_dlygate4sd3_1 hold895 (.A(_01695_),
    .X(net1958));
 sg13g2_dlygate4sd3_1 hold896 (.A(\inv_result[161] ),
    .X(net1959));
 sg13g2_dlygate4sd3_1 hold897 (.A(\u_inv.input_reg[142] ),
    .X(net1960));
 sg13g2_dlygate4sd3_1 hold898 (.A(_00049_),
    .X(net1961));
 sg13g2_dlygate4sd3_1 hold899 (.A(\trng_data[4] ),
    .X(net1962));
 sg13g2_dlygate4sd3_1 hold900 (.A(\u_inv.input_reg[251] ),
    .X(net1963));
 sg13g2_dlygate4sd3_1 hold901 (.A(_00158_),
    .X(net1964));
 sg13g2_dlygate4sd3_1 hold902 (.A(\inv_result[252] ),
    .X(net1965));
 sg13g2_dlygate4sd3_1 hold903 (.A(\u_inv.input_reg[55] ),
    .X(net1966));
 sg13g2_dlygate4sd3_1 hold904 (.A(_01861_),
    .X(net1967));
 sg13g2_dlygate4sd3_1 hold905 (.A(\inv_result[21] ),
    .X(net1968));
 sg13g2_dlygate4sd3_1 hold906 (.A(\shift_reg[1] ),
    .X(net1969));
 sg13g2_dlygate4sd3_1 hold907 (.A(_00176_),
    .X(net1970));
 sg13g2_dlygate4sd3_1 hold908 (.A(\u_inv.f_next[44] ),
    .X(net1971));
 sg13g2_dlygate4sd3_1 hold909 (.A(\u_inv.f_reg[137] ),
    .X(net1972));
 sg13g2_dlygate4sd3_1 hold910 (.A(_01644_),
    .X(net1973));
 sg13g2_dlygate4sd3_1 hold911 (.A(\shift_reg[136] ),
    .X(net1974));
 sg13g2_dlygate4sd3_1 hold912 (.A(_00311_),
    .X(net1975));
 sg13g2_dlygate4sd3_1 hold913 (.A(\shift_reg[123] ),
    .X(net1976));
 sg13g2_dlygate4sd3_1 hold914 (.A(_00298_),
    .X(net1977));
 sg13g2_dlygate4sd3_1 hold915 (.A(\u_inv.input_reg[175] ),
    .X(net1978));
 sg13g2_dlygate4sd3_1 hold916 (.A(_00082_),
    .X(net1979));
 sg13g2_dlygate4sd3_1 hold917 (.A(\u_inv.input_reg[164] ),
    .X(net1980));
 sg13g2_dlygate4sd3_1 hold918 (.A(_00071_),
    .X(net1981));
 sg13g2_dlygate4sd3_1 hold919 (.A(\u_inv.d_next[181] ),
    .X(net1982));
 sg13g2_dlygate4sd3_1 hold920 (.A(_01431_),
    .X(net1983));
 sg13g2_dlygate4sd3_1 hold921 (.A(\inv_result[209] ),
    .X(net1984));
 sg13g2_dlygate4sd3_1 hold922 (.A(\inv_result[191] ),
    .X(net1985));
 sg13g2_dlygate4sd3_1 hold923 (.A(\inv_result[39] ),
    .X(net1986));
 sg13g2_dlygate4sd3_1 hold924 (.A(\u_inv.d_next[220] ),
    .X(net1987));
 sg13g2_dlygate4sd3_1 hold925 (.A(_01470_),
    .X(net1988));
 sg13g2_dlygate4sd3_1 hold926 (.A(\u_inv.input_reg[249] ),
    .X(net1989));
 sg13g2_dlygate4sd3_1 hold927 (.A(_00156_),
    .X(net1990));
 sg13g2_dlygate4sd3_1 hold928 (.A(\inv_result[79] ),
    .X(net1991));
 sg13g2_dlygate4sd3_1 hold929 (.A(\u_inv.f_reg[120] ),
    .X(net1992));
 sg13g2_dlygate4sd3_1 hold930 (.A(_01627_),
    .X(net1993));
 sg13g2_dlygate4sd3_1 hold931 (.A(\inv_result[42] ),
    .X(net1994));
 sg13g2_dlygate4sd3_1 hold932 (.A(\inv_result[106] ),
    .X(net1995));
 sg13g2_dlygate4sd3_1 hold933 (.A(\u_inv.f_reg[189] ),
    .X(net1996));
 sg13g2_dlygate4sd3_1 hold934 (.A(_01696_),
    .X(net1997));
 sg13g2_dlygate4sd3_1 hold935 (.A(\inv_result[22] ),
    .X(net1998));
 sg13g2_dlygate4sd3_1 hold936 (.A(\u_inv.input_reg[190] ),
    .X(net1999));
 sg13g2_dlygate4sd3_1 hold937 (.A(_00097_),
    .X(net2000));
 sg13g2_dlygate4sd3_1 hold938 (.A(\inv_result[197] ),
    .X(net2001));
 sg13g2_dlygate4sd3_1 hold939 (.A(\inv_result[249] ),
    .X(net2002));
 sg13g2_dlygate4sd3_1 hold940 (.A(\u_inv.input_reg[78] ),
    .X(net2003));
 sg13g2_dlygate4sd3_1 hold941 (.A(_01884_),
    .X(net2004));
 sg13g2_dlygate4sd3_1 hold942 (.A(\inv_result[23] ),
    .X(net2005));
 sg13g2_dlygate4sd3_1 hold943 (.A(\u_inv.d_next[162] ),
    .X(net2006));
 sg13g2_dlygate4sd3_1 hold944 (.A(\u_inv.f_reg[22] ),
    .X(net2007));
 sg13g2_dlygate4sd3_1 hold945 (.A(_01529_),
    .X(net2008));
 sg13g2_dlygate4sd3_1 hold946 (.A(\u_inv.f_reg[113] ),
    .X(net2009));
 sg13g2_dlygate4sd3_1 hold947 (.A(_01620_),
    .X(net2010));
 sg13g2_dlygate4sd3_1 hold948 (.A(\inv_result[170] ),
    .X(net2011));
 sg13g2_dlygate4sd3_1 hold949 (.A(\inv_result[177] ),
    .X(net2012));
 sg13g2_dlygate4sd3_1 hold950 (.A(\inv_result[199] ),
    .X(net2013));
 sg13g2_dlygate4sd3_1 hold951 (.A(_01193_),
    .X(net2014));
 sg13g2_dlygate4sd3_1 hold952 (.A(\u_inv.input_reg[115] ),
    .X(net2015));
 sg13g2_dlygate4sd3_1 hold953 (.A(_00022_),
    .X(net2016));
 sg13g2_dlygate4sd3_1 hold954 (.A(\u_inv.f_reg[170] ),
    .X(net2017));
 sg13g2_dlygate4sd3_1 hold955 (.A(_01677_),
    .X(net2018));
 sg13g2_dlygate4sd3_1 hold956 (.A(\shift_reg[128] ),
    .X(net2019));
 sg13g2_dlygate4sd3_1 hold957 (.A(_00303_),
    .X(net2020));
 sg13g2_dlygate4sd3_1 hold958 (.A(\u_inv.input_reg[157] ),
    .X(net2021));
 sg13g2_dlygate4sd3_1 hold959 (.A(_00064_),
    .X(net2022));
 sg13g2_dlygate4sd3_1 hold960 (.A(\u_inv.f_reg[90] ),
    .X(net2023));
 sg13g2_dlygate4sd3_1 hold961 (.A(_01597_),
    .X(net2024));
 sg13g2_dlygate4sd3_1 hold962 (.A(\u_inv.f_reg[10] ),
    .X(net2025));
 sg13g2_dlygate4sd3_1 hold963 (.A(_01517_),
    .X(net2026));
 sg13g2_dlygate4sd3_1 hold964 (.A(\u_inv.f_reg[93] ),
    .X(net2027));
 sg13g2_dlygate4sd3_1 hold965 (.A(_01600_),
    .X(net2028));
 sg13g2_dlygate4sd3_1 hold966 (.A(\inv_result[220] ),
    .X(net2029));
 sg13g2_dlygate4sd3_1 hold967 (.A(\u_inv.f_reg[49] ),
    .X(net2030));
 sg13g2_dlygate4sd3_1 hold968 (.A(\u_inv.d_next[180] ),
    .X(net2031));
 sg13g2_dlygate4sd3_1 hold969 (.A(_01430_),
    .X(net2032));
 sg13g2_dlygate4sd3_1 hold970 (.A(\u_inv.d_next[222] ),
    .X(net2033));
 sg13g2_dlygate4sd3_1 hold971 (.A(_01472_),
    .X(net2034));
 sg13g2_dlygate4sd3_1 hold972 (.A(\u_inv.f_reg[39] ),
    .X(net2035));
 sg13g2_dlygate4sd3_1 hold973 (.A(_01546_),
    .X(net2036));
 sg13g2_dlygate4sd3_1 hold974 (.A(\inv_result[30] ),
    .X(net2037));
 sg13g2_dlygate4sd3_1 hold975 (.A(\u_inv.d_next[27] ),
    .X(net2038));
 sg13g2_dlygate4sd3_1 hold976 (.A(_01277_),
    .X(net2039));
 sg13g2_dlygate4sd3_1 hold977 (.A(\inv_result[40] ),
    .X(net2040));
 sg13g2_dlygate4sd3_1 hold978 (.A(\u_inv.input_reg[154] ),
    .X(net2041));
 sg13g2_dlygate4sd3_1 hold979 (.A(_00061_),
    .X(net2042));
 sg13g2_dlygate4sd3_1 hold980 (.A(\u_inv.f_reg[132] ),
    .X(net2043));
 sg13g2_dlygate4sd3_1 hold981 (.A(_01639_),
    .X(net2044));
 sg13g2_dlygate4sd3_1 hold982 (.A(\u_inv.f_reg[165] ),
    .X(net2045));
 sg13g2_dlygate4sd3_1 hold983 (.A(\inv_result[82] ),
    .X(net2046));
 sg13g2_dlygate4sd3_1 hold984 (.A(\inv_result[119] ),
    .X(net2047));
 sg13g2_dlygate4sd3_1 hold985 (.A(\u_inv.input_reg[159] ),
    .X(net2048));
 sg13g2_dlygate4sd3_1 hold986 (.A(_00066_),
    .X(net2049));
 sg13g2_dlygate4sd3_1 hold987 (.A(\u_inv.f_reg[87] ),
    .X(net2050));
 sg13g2_dlygate4sd3_1 hold988 (.A(\inv_result[194] ),
    .X(net2051));
 sg13g2_dlygate4sd3_1 hold989 (.A(\u_inv.f_next[216] ),
    .X(net2052));
 sg13g2_dlygate4sd3_1 hold990 (.A(\u_inv.input_reg[19] ),
    .X(net2053));
 sg13g2_dlygate4sd3_1 hold991 (.A(_01825_),
    .X(net2054));
 sg13g2_dlygate4sd3_1 hold992 (.A(\u_inv.f_reg[33] ),
    .X(net2055));
 sg13g2_dlygate4sd3_1 hold993 (.A(_01540_),
    .X(net2056));
 sg13g2_dlygate4sd3_1 hold994 (.A(\inv_result[122] ),
    .X(net2057));
 sg13g2_dlygate4sd3_1 hold995 (.A(\inv_result[28] ),
    .X(net2058));
 sg13g2_dlygate4sd3_1 hold996 (.A(\u_inv.input_reg[186] ),
    .X(net2059));
 sg13g2_dlygate4sd3_1 hold997 (.A(_00093_),
    .X(net2060));
 sg13g2_dlygate4sd3_1 hold998 (.A(\inv_result[96] ),
    .X(net2061));
 sg13g2_dlygate4sd3_1 hold999 (.A(\trng_data[3] ),
    .X(net2062));
 sg13g2_dlygate4sd3_1 hold1000 (.A(_00452_),
    .X(net2063));
 sg13g2_dlygate4sd3_1 hold1001 (.A(\u_inv.f_next[177] ),
    .X(net2064));
 sg13g2_dlygate4sd3_1 hold1002 (.A(\inv_result[167] ),
    .X(net2065));
 sg13g2_dlygate4sd3_1 hold1003 (.A(\inv_result[44] ),
    .X(net2066));
 sg13g2_dlygate4sd3_1 hold1004 (.A(\inv_result[151] ),
    .X(net2067));
 sg13g2_dlygate4sd3_1 hold1005 (.A(\inv_result[60] ),
    .X(net2068));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\perf_total[8] ),
    .X(net2069));
 sg13g2_dlygate4sd3_1 hold1007 (.A(\u_inv.f_reg[35] ),
    .X(net2070));
 sg13g2_dlygate4sd3_1 hold1008 (.A(_01542_),
    .X(net2071));
 sg13g2_dlygate4sd3_1 hold1009 (.A(\u_inv.f_reg[97] ),
    .X(net2072));
 sg13g2_dlygate4sd3_1 hold1010 (.A(_01604_),
    .X(net2073));
 sg13g2_dlygate4sd3_1 hold1011 (.A(\u_inv.d_next[178] ),
    .X(net2074));
 sg13g2_dlygate4sd3_1 hold1012 (.A(_01428_),
    .X(net2075));
 sg13g2_dlygate4sd3_1 hold1013 (.A(\u_inv.f_reg[24] ),
    .X(net2076));
 sg13g2_dlygate4sd3_1 hold1014 (.A(_01531_),
    .X(net2077));
 sg13g2_dlygate4sd3_1 hold1015 (.A(\inv_result[212] ),
    .X(net2078));
 sg13g2_dlygate4sd3_1 hold1016 (.A(\u_inv.f_reg[46] ),
    .X(net2079));
 sg13g2_dlygate4sd3_1 hold1017 (.A(_01553_),
    .X(net2080));
 sg13g2_dlygate4sd3_1 hold1018 (.A(\inv_result[56] ),
    .X(net2081));
 sg13g2_dlygate4sd3_1 hold1019 (.A(\u_inv.d_next[138] ),
    .X(net2082));
 sg13g2_dlygate4sd3_1 hold1020 (.A(\u_inv.d_next[94] ),
    .X(net2083));
 sg13g2_dlygate4sd3_1 hold1021 (.A(_01344_),
    .X(net2084));
 sg13g2_dlygate4sd3_1 hold1022 (.A(\u_inv.input_reg[72] ),
    .X(net2085));
 sg13g2_dlygate4sd3_1 hold1023 (.A(_01878_),
    .X(net2086));
 sg13g2_dlygate4sd3_1 hold1024 (.A(\u_inv.input_reg[93] ),
    .X(net2087));
 sg13g2_dlygate4sd3_1 hold1025 (.A(_01899_),
    .X(net2088));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\u_inv.input_reg[155] ),
    .X(net2089));
 sg13g2_dlygate4sd3_1 hold1027 (.A(_00062_),
    .X(net2090));
 sg13g2_dlygate4sd3_1 hold1028 (.A(\u_inv.f_reg[88] ),
    .X(net2091));
 sg13g2_dlygate4sd3_1 hold1029 (.A(_01595_),
    .X(net2092));
 sg13g2_dlygate4sd3_1 hold1030 (.A(\u_inv.input_reg[231] ),
    .X(net2093));
 sg13g2_dlygate4sd3_1 hold1031 (.A(_00138_),
    .X(net2094));
 sg13g2_dlygate4sd3_1 hold1032 (.A(\u_inv.d_next[182] ),
    .X(net2095));
 sg13g2_dlygate4sd3_1 hold1033 (.A(\inv_result[204] ),
    .X(net2096));
 sg13g2_dlygate4sd3_1 hold1035 (.A(\inv_result[246] ),
    .X(net2098));
 sg13g2_dlygate4sd3_1 hold1036 (.A(\inv_result[8] ),
    .X(net2099));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\u_inv.d_next[32] ),
    .X(net2100));
 sg13g2_dlygate4sd3_1 hold1038 (.A(_01282_),
    .X(net2101));
 sg13g2_dlygate4sd3_1 hold1039 (.A(\u_inv.f_reg[136] ),
    .X(net2102));
 sg13g2_dlygate4sd3_1 hold1040 (.A(_01643_),
    .X(net2103));
 sg13g2_dlygate4sd3_1 hold1041 (.A(\u_inv.f_reg[181] ),
    .X(net2104));
 sg13g2_dlygate4sd3_1 hold1042 (.A(_01688_),
    .X(net2105));
 sg13g2_dlygate4sd3_1 hold1043 (.A(\inv_result[29] ),
    .X(net2106));
 sg13g2_dlygate4sd3_1 hold1044 (.A(\u_inv.f_reg[82] ),
    .X(net2107));
 sg13g2_dlygate4sd3_1 hold1045 (.A(_01589_),
    .X(net2108));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\shift_reg[262] ),
    .X(net2109));
 sg13g2_dlygate4sd3_1 hold1047 (.A(_00437_),
    .X(net2110));
 sg13g2_dlygate4sd3_1 hold1048 (.A(\inv_result[5] ),
    .X(net2111));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\inv_result[233] ),
    .X(net2112));
 sg13g2_dlygate4sd3_1 hold1050 (.A(\u_inv.f_reg[67] ),
    .X(net2113));
 sg13g2_dlygate4sd3_1 hold1051 (.A(_01574_),
    .X(net2114));
 sg13g2_dlygate4sd3_1 hold1052 (.A(\shift_reg[117] ),
    .X(net2115));
 sg13g2_dlygate4sd3_1 hold1053 (.A(_00292_),
    .X(net2116));
 sg13g2_dlygate4sd3_1 hold1054 (.A(\u_inv.f_reg[40] ),
    .X(net2117));
 sg13g2_dlygate4sd3_1 hold1055 (.A(_01547_),
    .X(net2118));
 sg13g2_dlygate4sd3_1 hold1056 (.A(\u_inv.d_next[85] ),
    .X(net2119));
 sg13g2_dlygate4sd3_1 hold1057 (.A(\u_inv.d_next[60] ),
    .X(net2120));
 sg13g2_dlygate4sd3_1 hold1058 (.A(_01310_),
    .X(net2121));
 sg13g2_dlygate4sd3_1 hold1059 (.A(\u_inv.d_next[219] ),
    .X(net2122));
 sg13g2_dlygate4sd3_1 hold1060 (.A(_01469_),
    .X(net2123));
 sg13g2_dlygate4sd3_1 hold1061 (.A(\u_inv.f_next[15] ),
    .X(net2124));
 sg13g2_dlygate4sd3_1 hold1062 (.A(\inv_result[190] ),
    .X(net2125));
 sg13g2_dlygate4sd3_1 hold1063 (.A(\u_inv.d_next[237] ),
    .X(net2126));
 sg13g2_dlygate4sd3_1 hold1064 (.A(_01487_),
    .X(net2127));
 sg13g2_dlygate4sd3_1 hold1065 (.A(\inv_result[25] ),
    .X(net2128));
 sg13g2_dlygate4sd3_1 hold1066 (.A(\u_inv.f_reg[80] ),
    .X(net2129));
 sg13g2_dlygate4sd3_1 hold1067 (.A(_01587_),
    .X(net2130));
 sg13g2_dlygate4sd3_1 hold1068 (.A(\inv_result[84] ),
    .X(net2131));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\u_inv.f_next[7] ),
    .X(net2132));
 sg13g2_dlygate4sd3_1 hold1070 (.A(_01514_),
    .X(net2133));
 sg13g2_dlygate4sd3_1 hold1071 (.A(\u_inv.d_next[110] ),
    .X(net2134));
 sg13g2_dlygate4sd3_1 hold1072 (.A(\inv_result[80] ),
    .X(net2135));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\inv_result[13] ),
    .X(net2136));
 sg13g2_dlygate4sd3_1 hold1074 (.A(\u_inv.f_reg[45] ),
    .X(net2137));
 sg13g2_dlygate4sd3_1 hold1075 (.A(\shift_reg[244] ),
    .X(net2138));
 sg13g2_dlygate4sd3_1 hold1076 (.A(_00419_),
    .X(net2139));
 sg13g2_dlygate4sd3_1 hold1077 (.A(\u_inv.f_reg[237] ),
    .X(net2140));
 sg13g2_dlygate4sd3_1 hold1078 (.A(_01744_),
    .X(net2141));
 sg13g2_dlygate4sd3_1 hold1079 (.A(\u_inv.d_reg[182] ),
    .X(net2142));
 sg13g2_dlygate4sd3_1 hold1080 (.A(\u_inv.f_next[116] ),
    .X(net2143));
 sg13g2_dlygate4sd3_1 hold1081 (.A(_00576_),
    .X(net2144));
 sg13g2_dlygate4sd3_1 hold1082 (.A(\inv_result[123] ),
    .X(net2145));
 sg13g2_dlygate4sd3_1 hold1083 (.A(\u_inv.f_reg[235] ),
    .X(net2146));
 sg13g2_dlygate4sd3_1 hold1084 (.A(_01742_),
    .X(net2147));
 sg13g2_dlygate4sd3_1 hold1085 (.A(\inv_result[236] ),
    .X(net2148));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\u_inv.f_reg[131] ),
    .X(net2149));
 sg13g2_dlygate4sd3_1 hold1087 (.A(_01638_),
    .X(net2150));
 sg13g2_dlygate4sd3_1 hold1088 (.A(\u_inv.input_reg[41] ),
    .X(net2151));
 sg13g2_dlygate4sd3_1 hold1089 (.A(_01847_),
    .X(net2152));
 sg13g2_dlygate4sd3_1 hold1090 (.A(\u_inv.input_reg[74] ),
    .X(net2153));
 sg13g2_dlygate4sd3_1 hold1091 (.A(_01880_),
    .X(net2154));
 sg13g2_dlygate4sd3_1 hold1092 (.A(\inv_result[20] ),
    .X(net2155));
 sg13g2_dlygate4sd3_1 hold1093 (.A(\shift_reg[258] ),
    .X(net2156));
 sg13g2_dlygate4sd3_1 hold1094 (.A(_00433_),
    .X(net2157));
 sg13g2_dlygate4sd3_1 hold1095 (.A(\shift_reg[259] ),
    .X(net2158));
 sg13g2_dlygate4sd3_1 hold1096 (.A(_00434_),
    .X(net2159));
 sg13g2_dlygate4sd3_1 hold1097 (.A(\u_inv.f_reg[219] ),
    .X(net2160));
 sg13g2_dlygate4sd3_1 hold1098 (.A(\inv_result[75] ),
    .X(net2161));
 sg13g2_dlygate4sd3_1 hold1099 (.A(\inv_result[95] ),
    .X(net2162));
 sg13g2_dlygate4sd3_1 hold1100 (.A(\u_inv.f_reg[207] ),
    .X(net2163));
 sg13g2_dlygate4sd3_1 hold1101 (.A(_01714_),
    .X(net2164));
 sg13g2_dlygate4sd3_1 hold1102 (.A(\u_inv.f_reg[250] ),
    .X(net2165));
 sg13g2_dlygate4sd3_1 hold1103 (.A(_01757_),
    .X(net2166));
 sg13g2_dlygate4sd3_1 hold1104 (.A(\u_inv.f_reg[227] ),
    .X(net2167));
 sg13g2_dlygate4sd3_1 hold1105 (.A(_01734_),
    .X(net2168));
 sg13g2_dlygate4sd3_1 hold1106 (.A(\u_inv.f_reg[21] ),
    .X(net2169));
 sg13g2_dlygate4sd3_1 hold1107 (.A(_01528_),
    .X(net2170));
 sg13g2_dlygate4sd3_1 hold1108 (.A(\shift_reg[217] ),
    .X(net2171));
 sg13g2_dlygate4sd3_1 hold1109 (.A(_00392_),
    .X(net2172));
 sg13g2_dlygate4sd3_1 hold1110 (.A(\u_inv.f_reg[116] ),
    .X(net2173));
 sg13g2_dlygate4sd3_1 hold1111 (.A(\shift_reg[233] ),
    .X(net2174));
 sg13g2_dlygate4sd3_1 hold1112 (.A(_00408_),
    .X(net2175));
 sg13g2_dlygate4sd3_1 hold1113 (.A(\inv_result[162] ),
    .X(net2176));
 sg13g2_dlygate4sd3_1 hold1114 (.A(\u_inv.f_reg[155] ),
    .X(net2177));
 sg13g2_dlygate4sd3_1 hold1115 (.A(_01662_),
    .X(net2178));
 sg13g2_dlygate4sd3_1 hold1116 (.A(\inv_result[1] ),
    .X(net2179));
 sg13g2_dlygate4sd3_1 hold1117 (.A(_00995_),
    .X(net2180));
 sg13g2_dlygate4sd3_1 hold1118 (.A(\u_inv.f_reg[1] ),
    .X(net2181));
 sg13g2_dlygate4sd3_1 hold1119 (.A(_01508_),
    .X(net2182));
 sg13g2_dlygate4sd3_1 hold1120 (.A(\inv_result[112] ),
    .X(net2183));
 sg13g2_dlygate4sd3_1 hold1121 (.A(\inv_result[152] ),
    .X(net2184));
 sg13g2_dlygate4sd3_1 hold1122 (.A(\u_inv.f_reg[167] ),
    .X(net2185));
 sg13g2_dlygate4sd3_1 hold1123 (.A(_01674_),
    .X(net2186));
 sg13g2_dlygate4sd3_1 hold1124 (.A(\inv_result[200] ),
    .X(net2187));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\u_inv.input_reg[76] ),
    .X(net2188));
 sg13g2_dlygate4sd3_1 hold1126 (.A(_01882_),
    .X(net2189));
 sg13g2_dlygate4sd3_1 hold1127 (.A(\inv_result[118] ),
    .X(net2190));
 sg13g2_dlygate4sd3_1 hold1128 (.A(\u_inv.d_next[173] ),
    .X(net2191));
 sg13g2_dlygate4sd3_1 hold1129 (.A(_01423_),
    .X(net2192));
 sg13g2_dlygate4sd3_1 hold1130 (.A(\inv_result[254] ),
    .X(net2193));
 sg13g2_dlygate4sd3_1 hold1131 (.A(\u_inv.f_reg[78] ),
    .X(net2194));
 sg13g2_dlygate4sd3_1 hold1132 (.A(_01585_),
    .X(net2195));
 sg13g2_dlygate4sd3_1 hold1133 (.A(\u_inv.d_next[171] ),
    .X(net2196));
 sg13g2_dlygate4sd3_1 hold1134 (.A(_01421_),
    .X(net2197));
 sg13g2_dlygate4sd3_1 hold1135 (.A(\u_inv.f_reg[61] ),
    .X(net2198));
 sg13g2_dlygate4sd3_1 hold1136 (.A(_01568_),
    .X(net2199));
 sg13g2_dlygate4sd3_1 hold1137 (.A(\u_inv.f_reg[100] ),
    .X(net2200));
 sg13g2_dlygate4sd3_1 hold1138 (.A(_01607_),
    .X(net2201));
 sg13g2_dlygate4sd3_1 hold1139 (.A(\inv_cycles[1] ),
    .X(net2202));
 sg13g2_dlygate4sd3_1 hold1140 (.A(_01788_),
    .X(net2203));
 sg13g2_dlygate4sd3_1 hold1141 (.A(\u_inv.f_reg[190] ),
    .X(net2204));
 sg13g2_dlygate4sd3_1 hold1142 (.A(_01697_),
    .X(net2205));
 sg13g2_dlygate4sd3_1 hold1143 (.A(\u_inv.f_reg[223] ),
    .X(net2206));
 sg13g2_dlygate4sd3_1 hold1144 (.A(_01730_),
    .X(net2207));
 sg13g2_dlygate4sd3_1 hold1145 (.A(\shift_reg[257] ),
    .X(net2208));
 sg13g2_dlygate4sd3_1 hold1146 (.A(_00432_),
    .X(net2209));
 sg13g2_dlygate4sd3_1 hold1147 (.A(\inv_result[45] ),
    .X(net2210));
 sg13g2_dlygate4sd3_1 hold1148 (.A(\shift_reg[193] ),
    .X(net2211));
 sg13g2_dlygate4sd3_1 hold1149 (.A(_00368_),
    .X(net2212));
 sg13g2_dlygate4sd3_1 hold1150 (.A(\inv_result[193] ),
    .X(net2213));
 sg13g2_dlygate4sd3_1 hold1151 (.A(\u_inv.f_reg[95] ),
    .X(net2214));
 sg13g2_dlygate4sd3_1 hold1152 (.A(_01602_),
    .X(net2215));
 sg13g2_dlygate4sd3_1 hold1153 (.A(\u_inv.f_next[39] ),
    .X(net2216));
 sg13g2_dlygate4sd3_1 hold1154 (.A(\inv_result[46] ),
    .X(net2217));
 sg13g2_dlygate4sd3_1 hold1155 (.A(\inv_result[50] ),
    .X(net2218));
 sg13g2_dlygate4sd3_1 hold1156 (.A(\inv_result[41] ),
    .X(net2219));
 sg13g2_dlygate4sd3_1 hold1157 (.A(\u_inv.f_reg[94] ),
    .X(net2220));
 sg13g2_dlygate4sd3_1 hold1158 (.A(_01601_),
    .X(net2221));
 sg13g2_dlygate4sd3_1 hold1159 (.A(\u_inv.f_reg[99] ),
    .X(net2222));
 sg13g2_dlygate4sd3_1 hold1160 (.A(_01606_),
    .X(net2223));
 sg13g2_dlygate4sd3_1 hold1161 (.A(\u_inv.f_reg[11] ),
    .X(net2224));
 sg13g2_dlygate4sd3_1 hold1162 (.A(\u_inv.d_next[120] ),
    .X(net2225));
 sg13g2_dlygate4sd3_1 hold1163 (.A(_01370_),
    .X(net2226));
 sg13g2_dlygate4sd3_1 hold1164 (.A(\u_inv.f_reg[125] ),
    .X(net2227));
 sg13g2_dlygate4sd3_1 hold1165 (.A(_01632_),
    .X(net2228));
 sg13g2_dlygate4sd3_1 hold1166 (.A(\u_inv.input_reg[138] ),
    .X(net2229));
 sg13g2_dlygate4sd3_1 hold1167 (.A(_00045_),
    .X(net2230));
 sg13g2_dlygate4sd3_1 hold1168 (.A(\u_inv.f_reg[245] ),
    .X(net2231));
 sg13g2_dlygate4sd3_1 hold1169 (.A(_01752_),
    .X(net2232));
 sg13g2_dlygate4sd3_1 hold1170 (.A(\shift_reg[190] ),
    .X(net2233));
 sg13g2_dlygate4sd3_1 hold1171 (.A(_00365_),
    .X(net2234));
 sg13g2_dlygate4sd3_1 hold1172 (.A(\u_inv.d_next[239] ),
    .X(net2235));
 sg13g2_dlygate4sd3_1 hold1173 (.A(\inv_result[9] ),
    .X(net2236));
 sg13g2_dlygate4sd3_1 hold1174 (.A(\inv_result[48] ),
    .X(net2237));
 sg13g2_dlygate4sd3_1 hold1175 (.A(\u_inv.input_reg[151] ),
    .X(net2238));
 sg13g2_dlygate4sd3_1 hold1176 (.A(_00058_),
    .X(net2239));
 sg13g2_dlygate4sd3_1 hold1177 (.A(\u_inv.d_next[179] ),
    .X(net2240));
 sg13g2_dlygate4sd3_1 hold1178 (.A(\u_inv.f_reg[101] ),
    .X(net2241));
 sg13g2_dlygate4sd3_1 hold1179 (.A(_01608_),
    .X(net2242));
 sg13g2_dlygate4sd3_1 hold1180 (.A(\u_inv.f_reg[15] ),
    .X(net2243));
 sg13g2_dlygate4sd3_1 hold1181 (.A(\u_inv.f_reg[28] ),
    .X(net2244));
 sg13g2_dlygate4sd3_1 hold1182 (.A(_01535_),
    .X(net2245));
 sg13g2_dlygate4sd3_1 hold1183 (.A(\shift_reg[236] ),
    .X(net2246));
 sg13g2_dlygate4sd3_1 hold1184 (.A(_00411_),
    .X(net2247));
 sg13g2_dlygate4sd3_1 hold1185 (.A(\shift_reg[205] ),
    .X(net2248));
 sg13g2_dlygate4sd3_1 hold1186 (.A(_00380_),
    .X(net2249));
 sg13g2_dlygate4sd3_1 hold1187 (.A(\inv_result[67] ),
    .X(net2250));
 sg13g2_dlygate4sd3_1 hold1188 (.A(\shift_reg[39] ),
    .X(net2251));
 sg13g2_dlygate4sd3_1 hold1189 (.A(_00214_),
    .X(net2252));
 sg13g2_dlygate4sd3_1 hold1190 (.A(\u_inv.d_next[64] ),
    .X(net2253));
 sg13g2_dlygate4sd3_1 hold1191 (.A(_01314_),
    .X(net2254));
 sg13g2_dlygate4sd3_1 hold1192 (.A(\inv_result[174] ),
    .X(net2255));
 sg13g2_dlygate4sd3_1 hold1193 (.A(\u_trng.have_prev ),
    .X(net2256));
 sg13g2_dlygate4sd3_1 hold1194 (.A(_18632_),
    .X(net2257));
 sg13g2_dlygate4sd3_1 hold1195 (.A(\inv_result[97] ),
    .X(net2258));
 sg13g2_dlygate4sd3_1 hold1196 (.A(\inv_result[244] ),
    .X(net2259));
 sg13g2_dlygate4sd3_1 hold1197 (.A(\u_inv.input_reg[205] ),
    .X(net2260));
 sg13g2_dlygate4sd3_1 hold1198 (.A(_00112_),
    .X(net2261));
 sg13g2_dlygate4sd3_1 hold1199 (.A(\u_inv.input_reg[141] ),
    .X(net2262));
 sg13g2_dlygate4sd3_1 hold1200 (.A(_00048_),
    .X(net2263));
 sg13g2_dlygate4sd3_1 hold1201 (.A(\trng_data[2] ),
    .X(net2264));
 sg13g2_dlygate4sd3_1 hold1202 (.A(_00451_),
    .X(net2265));
 sg13g2_dlygate4sd3_1 hold1203 (.A(\u_inv.d_next[161] ),
    .X(net2266));
 sg13g2_dlygate4sd3_1 hold1204 (.A(_01411_),
    .X(net2267));
 sg13g2_dlygate4sd3_1 hold1205 (.A(\u_inv.d_next[28] ),
    .X(net2268));
 sg13g2_dlygate4sd3_1 hold1206 (.A(_01278_),
    .X(net2269));
 sg13g2_dlygate4sd3_1 hold1207 (.A(\shift_reg[247] ),
    .X(net2270));
 sg13g2_dlygate4sd3_1 hold1208 (.A(_00422_),
    .X(net2271));
 sg13g2_dlygate4sd3_1 hold1209 (.A(\u_inv.input_reg[214] ),
    .X(net2272));
 sg13g2_dlygate4sd3_1 hold1210 (.A(_00121_),
    .X(net2273));
 sg13g2_dlygate4sd3_1 hold1211 (.A(\u_inv.f_reg[142] ),
    .X(net2274));
 sg13g2_dlygate4sd3_1 hold1212 (.A(_01649_),
    .X(net2275));
 sg13g2_dlygate4sd3_1 hold1213 (.A(\inv_result[238] ),
    .X(net2276));
 sg13g2_dlygate4sd3_1 hold1214 (.A(\shift_reg[203] ),
    .X(net2277));
 sg13g2_dlygate4sd3_1 hold1215 (.A(_00378_),
    .X(net2278));
 sg13g2_dlygate4sd3_1 hold1216 (.A(\trng_data[1] ),
    .X(net2279));
 sg13g2_dlygate4sd3_1 hold1217 (.A(_00450_),
    .X(net2280));
 sg13g2_dlygate4sd3_1 hold1218 (.A(\inv_result[113] ),
    .X(net2281));
 sg13g2_dlygate4sd3_1 hold1219 (.A(\shift_reg[185] ),
    .X(net2282));
 sg13g2_dlygate4sd3_1 hold1220 (.A(\u_inv.d_next[212] ),
    .X(net2283));
 sg13g2_dlygate4sd3_1 hold1221 (.A(_01462_),
    .X(net2284));
 sg13g2_dlygate4sd3_1 hold1222 (.A(\inv_result[192] ),
    .X(net2285));
 sg13g2_dlygate4sd3_1 hold1223 (.A(\shift_reg[131] ),
    .X(net2286));
 sg13g2_dlygate4sd3_1 hold1224 (.A(\shift_reg[263] ),
    .X(net2287));
 sg13g2_dlygate4sd3_1 hold1225 (.A(_00438_),
    .X(net2288));
 sg13g2_dlygate4sd3_1 hold1226 (.A(\u_inv.input_reg[183] ),
    .X(net2289));
 sg13g2_dlygate4sd3_1 hold1227 (.A(_00090_),
    .X(net2290));
 sg13g2_dlygate4sd3_1 hold1228 (.A(\shift_reg[137] ),
    .X(net2291));
 sg13g2_dlygate4sd3_1 hold1229 (.A(_00312_),
    .X(net2292));
 sg13g2_dlygate4sd3_1 hold1230 (.A(\shift_reg[187] ),
    .X(net2293));
 sg13g2_dlygate4sd3_1 hold1231 (.A(_00362_),
    .X(net2294));
 sg13g2_dlygate4sd3_1 hold1232 (.A(\u_inv.f_reg[65] ),
    .X(net2295));
 sg13g2_dlygate4sd3_1 hold1233 (.A(_01572_),
    .X(net2296));
 sg13g2_dlygate4sd3_1 hold1234 (.A(\inv_result[19] ),
    .X(net2297));
 sg13g2_dlygate4sd3_1 hold1235 (.A(\u_inv.d_next[216] ),
    .X(net2298));
 sg13g2_dlygate4sd3_1 hold1236 (.A(_01466_),
    .X(net2299));
 sg13g2_dlygate4sd3_1 hold1237 (.A(\u_inv.f_next[55] ),
    .X(net2300));
 sg13g2_dlygate4sd3_1 hold1238 (.A(\u_inv.input_reg[209] ),
    .X(net2301));
 sg13g2_dlygate4sd3_1 hold1239 (.A(_00116_),
    .X(net2302));
 sg13g2_dlygate4sd3_1 hold1240 (.A(\shift_reg[135] ),
    .X(net2303));
 sg13g2_dlygate4sd3_1 hold1241 (.A(\inv_cycles[2] ),
    .X(net2304));
 sg13g2_dlygate4sd3_1 hold1242 (.A(_01789_),
    .X(net2305));
 sg13g2_dlygate4sd3_1 hold1243 (.A(\u_inv.f_reg[117] ),
    .X(net2306));
 sg13g2_dlygate4sd3_1 hold1244 (.A(_01624_),
    .X(net2307));
 sg13g2_dlygate4sd3_1 hold1245 (.A(\u_inv.f_reg[209] ),
    .X(net2308));
 sg13g2_dlygate4sd3_1 hold1246 (.A(_01716_),
    .X(net2309));
 sg13g2_dlygate4sd3_1 hold1247 (.A(\u_inv.d_next[243] ),
    .X(net2310));
 sg13g2_dlygate4sd3_1 hold1248 (.A(_01493_),
    .X(net2311));
 sg13g2_dlygate4sd3_1 hold1249 (.A(\u_inv.input_reg[187] ),
    .X(net2312));
 sg13g2_dlygate4sd3_1 hold1250 (.A(\inv_result[37] ),
    .X(net2313));
 sg13g2_dlygate4sd3_1 hold1251 (.A(\u_inv.d_next[184] ),
    .X(net2314));
 sg13g2_dlygate4sd3_1 hold1252 (.A(\inv_result[87] ),
    .X(net2315));
 sg13g2_dlygate4sd3_1 hold1253 (.A(\u_inv.d_next[90] ),
    .X(net2316));
 sg13g2_dlygate4sd3_1 hold1254 (.A(\u_inv.input_reg[128] ),
    .X(net2317));
 sg13g2_dlygate4sd3_1 hold1255 (.A(_00035_),
    .X(net2318));
 sg13g2_dlygate4sd3_1 hold1256 (.A(\u_inv.d_next[96] ),
    .X(net2319));
 sg13g2_dlygate4sd3_1 hold1257 (.A(_01346_),
    .X(net2320));
 sg13g2_dlygate4sd3_1 hold1258 (.A(\shift_reg[194] ),
    .X(net2321));
 sg13g2_dlygate4sd3_1 hold1259 (.A(_00369_),
    .X(net2322));
 sg13g2_dlygate4sd3_1 hold1260 (.A(\u_inv.input_reg[250] ),
    .X(net2323));
 sg13g2_dlygate4sd3_1 hold1261 (.A(_00157_),
    .X(net2324));
 sg13g2_dlygate4sd3_1 hold1262 (.A(\u_inv.d_next[79] ),
    .X(net2325));
 sg13g2_dlygate4sd3_1 hold1263 (.A(_01329_),
    .X(net2326));
 sg13g2_dlygate4sd3_1 hold1264 (.A(\u_inv.f_next[5] ),
    .X(net2327));
 sg13g2_dlygate4sd3_1 hold1265 (.A(\u_inv.d_next[115] ),
    .X(net2328));
 sg13g2_dlygate4sd3_1 hold1266 (.A(_01365_),
    .X(net2329));
 sg13g2_dlygate4sd3_1 hold1267 (.A(\shift_reg[238] ),
    .X(net2330));
 sg13g2_dlygate4sd3_1 hold1268 (.A(_00413_),
    .X(net2331));
 sg13g2_dlygate4sd3_1 hold1269 (.A(\u_inv.f_reg[241] ),
    .X(net2332));
 sg13g2_dlygate4sd3_1 hold1270 (.A(_01748_),
    .X(net2333));
 sg13g2_dlygate4sd3_1 hold1271 (.A(\shift_reg[120] ),
    .X(net2334));
 sg13g2_dlygate4sd3_1 hold1272 (.A(_00295_),
    .X(net2335));
 sg13g2_dlygate4sd3_1 hold1273 (.A(\inv_result[3] ),
    .X(net2336));
 sg13g2_dlygate4sd3_1 hold1274 (.A(_00997_),
    .X(net2337));
 sg13g2_dlygate4sd3_1 hold1275 (.A(\inv_result[120] ),
    .X(net2338));
 sg13g2_dlygate4sd3_1 hold1276 (.A(\u_inv.f_reg[112] ),
    .X(net2339));
 sg13g2_dlygate4sd3_1 hold1277 (.A(_01619_),
    .X(net2340));
 sg13g2_dlygate4sd3_1 hold1278 (.A(\u_inv.f_reg[66] ),
    .X(net2341));
 sg13g2_dlygate4sd3_1 hold1279 (.A(_01573_),
    .X(net2342));
 sg13g2_dlygate4sd3_1 hold1280 (.A(\inv_result[201] ),
    .X(net2343));
 sg13g2_dlygate4sd3_1 hold1281 (.A(\u_inv.f_reg[51] ),
    .X(net2344));
 sg13g2_dlygate4sd3_1 hold1282 (.A(_01558_),
    .X(net2345));
 sg13g2_dlygate4sd3_1 hold1283 (.A(\u_inv.input_reg[121] ),
    .X(net2346));
 sg13g2_dlygate4sd3_1 hold1284 (.A(\shift_reg[124] ),
    .X(net2347));
 sg13g2_dlygate4sd3_1 hold1285 (.A(_00299_),
    .X(net2348));
 sg13g2_dlygate4sd3_1 hold1286 (.A(\u_inv.f_reg[204] ),
    .X(net2349));
 sg13g2_dlygate4sd3_1 hold1287 (.A(_01711_),
    .X(net2350));
 sg13g2_dlygate4sd3_1 hold1288 (.A(\shift_reg[195] ),
    .X(net2351));
 sg13g2_dlygate4sd3_1 hold1289 (.A(_00370_),
    .X(net2352));
 sg13g2_dlygate4sd3_1 hold1290 (.A(\u_inv.input_reg[168] ),
    .X(net2353));
 sg13g2_dlygate4sd3_1 hold1291 (.A(_00075_),
    .X(net2354));
 sg13g2_dlygate4sd3_1 hold1292 (.A(\u_inv.f_reg[159] ),
    .X(net2355));
 sg13g2_dlygate4sd3_1 hold1293 (.A(_01666_),
    .X(net2356));
 sg13g2_dlygate4sd3_1 hold1294 (.A(\u_inv.input_reg[145] ),
    .X(net2357));
 sg13g2_dlygate4sd3_1 hold1295 (.A(_00052_),
    .X(net2358));
 sg13g2_dlygate4sd3_1 hold1296 (.A(\u_inv.f_reg[91] ),
    .X(net2359));
 sg13g2_dlygate4sd3_1 hold1297 (.A(_01598_),
    .X(net2360));
 sg13g2_dlygate4sd3_1 hold1298 (.A(\u_inv.d_next[118] ),
    .X(net2361));
 sg13g2_dlygate4sd3_1 hold1299 (.A(\u_inv.input_reg[144] ),
    .X(net2362));
 sg13g2_dlygate4sd3_1 hold1300 (.A(_00051_),
    .X(net2363));
 sg13g2_dlygate4sd3_1 hold1301 (.A(\u_inv.f_reg[79] ),
    .X(net2364));
 sg13g2_dlygate4sd3_1 hold1302 (.A(_01586_),
    .X(net2365));
 sg13g2_dlygate4sd3_1 hold1303 (.A(\u_inv.d_next[80] ),
    .X(net2366));
 sg13g2_dlygate4sd3_1 hold1304 (.A(_01330_),
    .X(net2367));
 sg13g2_dlygate4sd3_1 hold1305 (.A(\u_inv.d_next[218] ),
    .X(net2368));
 sg13g2_dlygate4sd3_1 hold1306 (.A(_01468_),
    .X(net2369));
 sg13g2_dlygate4sd3_1 hold1307 (.A(\u_inv.input_reg[106] ),
    .X(net2370));
 sg13g2_dlygate4sd3_1 hold1308 (.A(_00013_),
    .X(net2371));
 sg13g2_dlygate4sd3_1 hold1309 (.A(\u_inv.f_next[181] ),
    .X(net2372));
 sg13g2_dlygate4sd3_1 hold1310 (.A(\inv_result[74] ),
    .X(net2373));
 sg13g2_dlygate4sd3_1 hold1311 (.A(\u_inv.f_reg[140] ),
    .X(net2374));
 sg13g2_dlygate4sd3_1 hold1312 (.A(_01647_),
    .X(net2375));
 sg13g2_dlygate4sd3_1 hold1313 (.A(\u_inv.d_next[236] ),
    .X(net2376));
 sg13g2_dlygate4sd3_1 hold1314 (.A(\u_inv.f_reg[166] ),
    .X(net2377));
 sg13g2_dlygate4sd3_1 hold1315 (.A(_01673_),
    .X(net2378));
 sg13g2_dlygate4sd3_1 hold1316 (.A(\inv_result[47] ),
    .X(net2379));
 sg13g2_dlygate4sd3_1 hold1317 (.A(\u_inv.f_next[199] ),
    .X(net2380));
 sg13g2_dlygate4sd3_1 hold1318 (.A(\u_inv.d_next[18] ),
    .X(net2381));
 sg13g2_dlygate4sd3_1 hold1319 (.A(\u_inv.input_reg[189] ),
    .X(net2382));
 sg13g2_dlygate4sd3_1 hold1320 (.A(\u_inv.d_reg[110] ),
    .X(net2383));
 sg13g2_dlygate4sd3_1 hold1321 (.A(\u_inv.f_reg[199] ),
    .X(net2384));
 sg13g2_dlygate4sd3_1 hold1322 (.A(\u_inv.f_reg[194] ),
    .X(net2385));
 sg13g2_dlygate4sd3_1 hold1323 (.A(_01701_),
    .X(net2386));
 sg13g2_dlygate4sd3_1 hold1324 (.A(\u_inv.f_reg[216] ),
    .X(net2387));
 sg13g2_dlygate4sd3_1 hold1325 (.A(\u_inv.f_reg[58] ),
    .X(net2388));
 sg13g2_dlygate4sd3_1 hold1326 (.A(_01565_),
    .X(net2389));
 sg13g2_dlygate4sd3_1 hold1327 (.A(\inv_result[105] ),
    .X(net2390));
 sg13g2_dlygate4sd3_1 hold1328 (.A(\shift_reg[246] ),
    .X(net2391));
 sg13g2_dlygate4sd3_1 hold1329 (.A(_00421_),
    .X(net2392));
 sg13g2_dlygate4sd3_1 hold1330 (.A(\u_inv.f_reg[31] ),
    .X(net2393));
 sg13g2_dlygate4sd3_1 hold1331 (.A(_01538_),
    .X(net2394));
 sg13g2_dlygate4sd3_1 hold1332 (.A(\u_inv.f_reg[85] ),
    .X(net2395));
 sg13g2_dlygate4sd3_1 hold1333 (.A(_01592_),
    .X(net2396));
 sg13g2_dlygate4sd3_1 hold1334 (.A(\u_inv.d_next[123] ),
    .X(net2397));
 sg13g2_dlygate4sd3_1 hold1335 (.A(_01373_),
    .X(net2398));
 sg13g2_dlygate4sd3_1 hold1336 (.A(\u_inv.input_reg[130] ),
    .X(net2399));
 sg13g2_dlygate4sd3_1 hold1337 (.A(_00037_),
    .X(net2400));
 sg13g2_dlygate4sd3_1 hold1338 (.A(\u_inv.d_next[126] ),
    .X(net2401));
 sg13g2_dlygate4sd3_1 hold1339 (.A(_01376_),
    .X(net2402));
 sg13g2_dlygate4sd3_1 hold1340 (.A(\shift_reg[243] ),
    .X(net2403));
 sg13g2_dlygate4sd3_1 hold1341 (.A(_00418_),
    .X(net2404));
 sg13g2_dlygate4sd3_1 hold1342 (.A(\u_inv.f_reg[102] ),
    .X(net2405));
 sg13g2_dlygate4sd3_1 hold1343 (.A(_01609_),
    .X(net2406));
 sg13g2_dlygate4sd3_1 hold1344 (.A(\u_inv.f_next[131] ),
    .X(net2407));
 sg13g2_dlygate4sd3_1 hold1345 (.A(\u_inv.f_reg[201] ),
    .X(net2408));
 sg13g2_dlygate4sd3_1 hold1346 (.A(_01708_),
    .X(net2409));
 sg13g2_dlygate4sd3_1 hold1347 (.A(\shift_reg[88] ),
    .X(net2410));
 sg13g2_dlygate4sd3_1 hold1348 (.A(_00263_),
    .X(net2411));
 sg13g2_dlygate4sd3_1 hold1349 (.A(\inv_result[17] ),
    .X(net2412));
 sg13g2_dlygate4sd3_1 hold1350 (.A(\u_inv.f_reg[114] ),
    .X(net2413));
 sg13g2_dlygate4sd3_1 hold1351 (.A(_01621_),
    .X(net2414));
 sg13g2_dlygate4sd3_1 hold1352 (.A(\u_inv.f_reg[76] ),
    .X(net2415));
 sg13g2_dlygate4sd3_1 hold1353 (.A(_01583_),
    .X(net2416));
 sg13g2_dlygate4sd3_1 hold1354 (.A(\u_inv.d_next[221] ),
    .X(net2417));
 sg13g2_dlygate4sd3_1 hold1355 (.A(_01471_),
    .X(net2418));
 sg13g2_dlygate4sd3_1 hold1356 (.A(\u_inv.f_reg[193] ),
    .X(net2419));
 sg13g2_dlygate4sd3_1 hold1357 (.A(_01700_),
    .X(net2420));
 sg13g2_dlygate4sd3_1 hold1358 (.A(\perf_triple[6] ),
    .X(net2421));
 sg13g2_dlygate4sd3_1 hold1359 (.A(\u_inv.f_next[26] ),
    .X(net2422));
 sg13g2_dlygate4sd3_1 hold1360 (.A(\shift_reg[121] ),
    .X(net2423));
 sg13g2_dlygate4sd3_1 hold1361 (.A(_00296_),
    .X(net2424));
 sg13g2_dlygate4sd3_1 hold1362 (.A(\u_inv.f_reg[56] ),
    .X(net2425));
 sg13g2_dlygate4sd3_1 hold1363 (.A(_01563_),
    .X(net2426));
 sg13g2_dlygate4sd3_1 hold1364 (.A(\u_inv.d_next[170] ),
    .X(net2427));
 sg13g2_dlygate4sd3_1 hold1365 (.A(\shift_reg[134] ),
    .X(net2428));
 sg13g2_dlygate4sd3_1 hold1366 (.A(_00309_),
    .X(net2429));
 sg13g2_dlygate4sd3_1 hold1367 (.A(\shift_reg[271] ),
    .X(net2430));
 sg13g2_dlygate4sd3_1 hold1368 (.A(_00446_),
    .X(net2431));
 sg13g2_dlygate4sd3_1 hold1369 (.A(\u_inv.f_reg[169] ),
    .X(net2432));
 sg13g2_dlygate4sd3_1 hold1370 (.A(_01676_),
    .X(net2433));
 sg13g2_dlygate4sd3_1 hold1371 (.A(\shift_reg[83] ),
    .X(net2434));
 sg13g2_dlygate4sd3_1 hold1372 (.A(_00258_),
    .X(net2435));
 sg13g2_dlygate4sd3_1 hold1373 (.A(\u_inv.d_next[62] ),
    .X(net2436));
 sg13g2_dlygate4sd3_1 hold1374 (.A(\u_inv.d_next[124] ),
    .X(net2437));
 sg13g2_dlygate4sd3_1 hold1375 (.A(_01374_),
    .X(net2438));
 sg13g2_dlygate4sd3_1 hold1376 (.A(\u_inv.f_next[41] ),
    .X(net2439));
 sg13g2_dlygate4sd3_1 hold1377 (.A(\u_inv.d_next[186] ),
    .X(net2440));
 sg13g2_dlygate4sd3_1 hold1378 (.A(_01436_),
    .X(net2441));
 sg13g2_dlygate4sd3_1 hold1379 (.A(\shift_reg[184] ),
    .X(net2442));
 sg13g2_dlygate4sd3_1 hold1380 (.A(\u_inv.d_reg[57] ),
    .X(net2443));
 sg13g2_dlygate4sd3_1 hold1381 (.A(_01307_),
    .X(net2444));
 sg13g2_dlygate4sd3_1 hold1382 (.A(\u_inv.f_reg[215] ),
    .X(net2445));
 sg13g2_dlygate4sd3_1 hold1383 (.A(_01722_),
    .X(net2446));
 sg13g2_dlygate4sd3_1 hold1384 (.A(\u_inv.d_next[194] ),
    .X(net2447));
 sg13g2_dlygate4sd3_1 hold1385 (.A(_01444_),
    .X(net2448));
 sg13g2_dlygate4sd3_1 hold1386 (.A(\inv_result[86] ),
    .X(net2449));
 sg13g2_dlygate4sd3_1 hold1387 (.A(\u_inv.d_next[246] ),
    .X(net2450));
 sg13g2_dlygate4sd3_1 hold1388 (.A(\shift_reg[122] ),
    .X(net2451));
 sg13g2_dlygate4sd3_1 hold1389 (.A(_00297_),
    .X(net2452));
 sg13g2_dlygate4sd3_1 hold1390 (.A(\u_inv.f_reg[52] ),
    .X(net2453));
 sg13g2_dlygate4sd3_1 hold1391 (.A(_01559_),
    .X(net2454));
 sg13g2_dlygate4sd3_1 hold1392 (.A(\u_inv.d_reg[179] ),
    .X(net2455));
 sg13g2_dlygate4sd3_1 hold1393 (.A(\u_inv.d_next[204] ),
    .X(net2456));
 sg13g2_dlygate4sd3_1 hold1394 (.A(\u_inv.input_reg[213] ),
    .X(net2457));
 sg13g2_dlygate4sd3_1 hold1395 (.A(_00120_),
    .X(net2458));
 sg13g2_dlygate4sd3_1 hold1396 (.A(\shift_reg[125] ),
    .X(net2459));
 sg13g2_dlygate4sd3_1 hold1397 (.A(\u_inv.f_reg[81] ),
    .X(net2460));
 sg13g2_dlygate4sd3_1 hold1398 (.A(_01588_),
    .X(net2461));
 sg13g2_dlygate4sd3_1 hold1399 (.A(\u_inv.f_reg[211] ),
    .X(net2462));
 sg13g2_dlygate4sd3_1 hold1400 (.A(_01718_),
    .X(net2463));
 sg13g2_dlygate4sd3_1 hold1401 (.A(\u_inv.d_next[5] ),
    .X(net2464));
 sg13g2_dlygate4sd3_1 hold1402 (.A(_01255_),
    .X(net2465));
 sg13g2_dlygate4sd3_1 hold1403 (.A(\shift_reg[12] ),
    .X(net2466));
 sg13g2_dlygate4sd3_1 hold1404 (.A(_00187_),
    .X(net2467));
 sg13g2_dlygate4sd3_1 hold1405 (.A(\u_inv.f_reg[177] ),
    .X(net2468));
 sg13g2_dlygate4sd3_1 hold1406 (.A(\inv_result[4] ),
    .X(net2469));
 sg13g2_dlygate4sd3_1 hold1407 (.A(_00998_),
    .X(net2470));
 sg13g2_dlygate4sd3_1 hold1408 (.A(\u_inv.d_next[158] ),
    .X(net2471));
 sg13g2_dlygate4sd3_1 hold1409 (.A(_01408_),
    .X(net2472));
 sg13g2_dlygate4sd3_1 hold1410 (.A(\u_inv.input_reg[139] ),
    .X(net2473));
 sg13g2_dlygate4sd3_1 hold1411 (.A(_00046_),
    .X(net2474));
 sg13g2_dlygate4sd3_1 hold1412 (.A(\u_inv.d_next[92] ),
    .X(net2475));
 sg13g2_dlygate4sd3_1 hold1413 (.A(_01342_),
    .X(net2476));
 sg13g2_dlygate4sd3_1 hold1414 (.A(\u_inv.input_reg[160] ),
    .X(net2477));
 sg13g2_dlygate4sd3_1 hold1415 (.A(_00067_),
    .X(net2478));
 sg13g2_dlygate4sd3_1 hold1416 (.A(\shift_reg[266] ),
    .X(net2479));
 sg13g2_dlygate4sd3_1 hold1417 (.A(\u_inv.d_next[48] ),
    .X(net2480));
 sg13g2_dlygate4sd3_1 hold1418 (.A(_01298_),
    .X(net2481));
 sg13g2_dlygate4sd3_1 hold1419 (.A(\u_inv.d_next[13] ),
    .X(net2482));
 sg13g2_dlygate4sd3_1 hold1420 (.A(\u_inv.d_next[55] ),
    .X(net2483));
 sg13g2_dlygate4sd3_1 hold1421 (.A(\u_inv.input_reg[204] ),
    .X(net2484));
 sg13g2_dlygate4sd3_1 hold1422 (.A(_00111_),
    .X(net2485));
 sg13g2_dlygate4sd3_1 hold1423 (.A(\byte_cnt[5] ),
    .X(net2486));
 sg13g2_dlygate4sd3_1 hold1424 (.A(_00174_),
    .X(net2487));
 sg13g2_dlygate4sd3_1 hold1425 (.A(\u_inv.f_reg[141] ),
    .X(net2488));
 sg13g2_dlygate4sd3_1 hold1426 (.A(_01648_),
    .X(net2489));
 sg13g2_dlygate4sd3_1 hold1427 (.A(\u_inv.d_next[153] ),
    .X(net2490));
 sg13g2_dlygate4sd3_1 hold1428 (.A(\u_inv.f_reg[96] ),
    .X(net2491));
 sg13g2_dlygate4sd3_1 hold1429 (.A(_01603_),
    .X(net2492));
 sg13g2_dlygate4sd3_1 hold1430 (.A(\u_inv.f_next[175] ),
    .X(net2493));
 sg13g2_dlygate4sd3_1 hold1431 (.A(\u_inv.f_next[65] ),
    .X(net2494));
 sg13g2_dlygate4sd3_1 hold1432 (.A(\u_inv.input_reg[147] ),
    .X(net2495));
 sg13g2_dlygate4sd3_1 hold1433 (.A(_00054_),
    .X(net2496));
 sg13g2_dlygate4sd3_1 hold1434 (.A(\u_inv.f_reg[0] ),
    .X(net2497));
 sg13g2_dlygate4sd3_1 hold1435 (.A(\u_inv.f_next[224] ),
    .X(net2498));
 sg13g2_dlygate4sd3_1 hold1436 (.A(\inv_result[55] ),
    .X(net2499));
 sg13g2_dlygate4sd3_1 hold1438 (.A(\u_inv.f_reg[68] ),
    .X(net2501));
 sg13g2_dlygate4sd3_1 hold1439 (.A(_01575_),
    .X(net2502));
 sg13g2_dlygate4sd3_1 hold1440 (.A(\u_inv.f_reg[129] ),
    .X(net2503));
 sg13g2_dlygate4sd3_1 hold1441 (.A(_01636_),
    .X(net2504));
 sg13g2_dlygate4sd3_1 hold1442 (.A(\u_inv.input_reg[252] ),
    .X(net2505));
 sg13g2_dlygate4sd3_1 hold1443 (.A(_00159_),
    .X(net2506));
 sg13g2_dlygate4sd3_1 hold1444 (.A(\shift_reg[206] ),
    .X(net2507));
 sg13g2_dlygate4sd3_1 hold1445 (.A(_00381_),
    .X(net2508));
 sg13g2_dlygate4sd3_1 hold1446 (.A(\shift_reg[252] ),
    .X(net2509));
 sg13g2_dlygate4sd3_1 hold1447 (.A(_00427_),
    .X(net2510));
 sg13g2_dlygate4sd3_1 hold1448 (.A(\inv_result[51] ),
    .X(net2511));
 sg13g2_dlygate4sd3_1 hold1449 (.A(\u_inv.input_reg[116] ),
    .X(net2512));
 sg13g2_dlygate4sd3_1 hold1450 (.A(_00023_),
    .X(net2513));
 sg13g2_dlygate4sd3_1 hold1451 (.A(\u_inv.d_next[2] ),
    .X(net2514));
 sg13g2_dlygate4sd3_1 hold1452 (.A(_01252_),
    .X(net2515));
 sg13g2_dlygate4sd3_1 hold1453 (.A(\u_inv.f_reg[214] ),
    .X(net2516));
 sg13g2_dlygate4sd3_1 hold1454 (.A(_01721_),
    .X(net2517));
 sg13g2_dlygate4sd3_1 hold1455 (.A(\inv_result[207] ),
    .X(net2518));
 sg13g2_dlygate4sd3_1 hold1456 (.A(\shift_reg[232] ),
    .X(net2519));
 sg13g2_dlygate4sd3_1 hold1457 (.A(_00407_),
    .X(net2520));
 sg13g2_dlygate4sd3_1 hold1458 (.A(\u_inv.d_next[66] ),
    .X(net2521));
 sg13g2_dlygate4sd3_1 hold1459 (.A(_01316_),
    .X(net2522));
 sg13g2_dlygate4sd3_1 hold1460 (.A(\u_inv.input_reg[219] ),
    .X(net2523));
 sg13g2_dlygate4sd3_1 hold1461 (.A(_00126_),
    .X(net2524));
 sg13g2_dlygate4sd3_1 hold1462 (.A(\shift_reg[240] ),
    .X(net2525));
 sg13g2_dlygate4sd3_1 hold1463 (.A(\u_inv.f_reg[252] ),
    .X(net2526));
 sg13g2_dlygate4sd3_1 hold1464 (.A(_01759_),
    .X(net2527));
 sg13g2_dlygate4sd3_1 hold1465 (.A(\u_inv.f_next[96] ),
    .X(net2528));
 sg13g2_dlygate4sd3_1 hold1466 (.A(\u_inv.f_next[88] ),
    .X(net2529));
 sg13g2_dlygate4sd3_1 hold1467 (.A(\inv_result[237] ),
    .X(net2530));
 sg13g2_dlygate4sd3_1 hold1468 (.A(\u_inv.f_reg[206] ),
    .X(net2531));
 sg13g2_dlygate4sd3_1 hold1469 (.A(_01713_),
    .X(net2532));
 sg13g2_dlygate4sd3_1 hold1470 (.A(\u_inv.d_next[225] ),
    .X(net2533));
 sg13g2_dlygate4sd3_1 hold1471 (.A(\u_inv.f_next[52] ),
    .X(net2534));
 sg13g2_dlygate4sd3_1 hold1472 (.A(\shift_reg[197] ),
    .X(net2535));
 sg13g2_dlygate4sd3_1 hold1473 (.A(_00372_),
    .X(net2536));
 sg13g2_dlygate4sd3_1 hold1474 (.A(\u_inv.d_next[24] ),
    .X(net2537));
 sg13g2_dlygate4sd3_1 hold1475 (.A(\u_inv.d_next[88] ),
    .X(net2538));
 sg13g2_dlygate4sd3_1 hold1476 (.A(_01338_),
    .X(net2539));
 sg13g2_dlygate4sd3_1 hold1477 (.A(\u_inv.f_reg[158] ),
    .X(net2540));
 sg13g2_dlygate4sd3_1 hold1478 (.A(_01665_),
    .X(net2541));
 sg13g2_dlygate4sd3_1 hold1479 (.A(\u_trng.prev_sample ),
    .X(net2542));
 sg13g2_dlygate4sd3_1 hold1480 (.A(_00458_),
    .X(net2543));
 sg13g2_dlygate4sd3_1 hold1481 (.A(\inv_result[100] ),
    .X(net2544));
 sg13g2_dlygate4sd3_1 hold1482 (.A(\u_inv.f_next[95] ),
    .X(net2545));
 sg13g2_dlygate4sd3_1 hold1483 (.A(\shift_reg[209] ),
    .X(net2546));
 sg13g2_dlygate4sd3_1 hold1484 (.A(_00384_),
    .X(net2547));
 sg13g2_dlygate4sd3_1 hold1485 (.A(\u_inv.d_next[190] ),
    .X(net2548));
 sg13g2_dlygate4sd3_1 hold1486 (.A(\shift_reg[241] ),
    .X(net2549));
 sg13g2_dlygate4sd3_1 hold1487 (.A(_00416_),
    .X(net2550));
 sg13g2_dlygate4sd3_1 hold1488 (.A(\inv_result[6] ),
    .X(net2551));
 sg13g2_dlygate4sd3_1 hold1489 (.A(\u_inv.input_reg[135] ),
    .X(net2552));
 sg13g2_dlygate4sd3_1 hold1490 (.A(_00042_),
    .X(net2553));
 sg13g2_dlygate4sd3_1 hold1491 (.A(\shift_reg[112] ),
    .X(net2554));
 sg13g2_dlygate4sd3_1 hold1492 (.A(_00287_),
    .X(net2555));
 sg13g2_dlygate4sd3_1 hold1493 (.A(\shift_reg[199] ),
    .X(net2556));
 sg13g2_dlygate4sd3_1 hold1494 (.A(_00374_),
    .X(net2557));
 sg13g2_dlygate4sd3_1 hold1495 (.A(\inv_result[63] ),
    .X(net2558));
 sg13g2_dlygate4sd3_1 hold1496 (.A(\u_inv.f_reg[186] ),
    .X(net2559));
 sg13g2_dlygate4sd3_1 hold1497 (.A(_01693_),
    .X(net2560));
 sg13g2_dlygate4sd3_1 hold1498 (.A(\u_inv.d_next[198] ),
    .X(net2561));
 sg13g2_dlygate4sd3_1 hold1499 (.A(net7293),
    .X(net2562));
 sg13g2_dlygate4sd3_1 hold1500 (.A(\u_inv.f_next[112] ),
    .X(net2563));
 sg13g2_dlygate4sd3_1 hold1501 (.A(\shift_reg[250] ),
    .X(net2564));
 sg13g2_dlygate4sd3_1 hold1502 (.A(_00425_),
    .X(net2565));
 sg13g2_dlygate4sd3_1 hold1503 (.A(\inv_result[62] ),
    .X(net2566));
 sg13g2_dlygate4sd3_1 hold1504 (.A(\u_inv.f_reg[195] ),
    .X(net2567));
 sg13g2_dlygate4sd3_1 hold1505 (.A(_01702_),
    .X(net2568));
 sg13g2_dlygate4sd3_1 hold1506 (.A(\u_inv.input_reg[119] ),
    .X(net2569));
 sg13g2_dlygate4sd3_1 hold1507 (.A(\shift_reg[270] ),
    .X(net2570));
 sg13g2_dlygate4sd3_1 hold1508 (.A(\shift_reg[99] ),
    .X(net2571));
 sg13g2_dlygate4sd3_1 hold1509 (.A(_00274_),
    .X(net2572));
 sg13g2_dlygate4sd3_1 hold1510 (.A(\u_inv.f_reg[105] ),
    .X(net2573));
 sg13g2_dlygate4sd3_1 hold1511 (.A(\shift_reg[268] ),
    .X(net2574));
 sg13g2_dlygate4sd3_1 hold1512 (.A(_00443_),
    .X(net2575));
 sg13g2_dlygate4sd3_1 hold1513 (.A(\shift_reg[133] ),
    .X(net2576));
 sg13g2_dlygate4sd3_1 hold1514 (.A(_00308_),
    .X(net2577));
 sg13g2_dlygate4sd3_1 hold1515 (.A(\u_inv.d_next[175] ),
    .X(net2578));
 sg13g2_dlygate4sd3_1 hold1516 (.A(_01425_),
    .X(net2579));
 sg13g2_dlygate4sd3_1 hold1517 (.A(\u_inv.f_next[104] ),
    .X(net2580));
 sg13g2_dlygate4sd3_1 hold1518 (.A(\u_inv.d_next[150] ),
    .X(net2581));
 sg13g2_dlygate4sd3_1 hold1519 (.A(\inv_result[134] ),
    .X(net2582));
 sg13g2_dlygate4sd3_1 hold1520 (.A(\u_inv.d_reg[13] ),
    .X(net2583));
 sg13g2_dlygate4sd3_1 hold1521 (.A(\shift_reg[255] ),
    .X(net2584));
 sg13g2_dlygate4sd3_1 hold1522 (.A(\u_inv.d_next[76] ),
    .X(net2585));
 sg13g2_dlygate4sd3_1 hold1523 (.A(_01326_),
    .X(net2586));
 sg13g2_dlygate4sd3_1 hold1524 (.A(\u_inv.d_next[128] ),
    .X(net2587));
 sg13g2_dlygate4sd3_1 hold1525 (.A(_01378_),
    .X(net2588));
 sg13g2_dlygate4sd3_1 hold1526 (.A(\u_inv.d_next[152] ),
    .X(net2589));
 sg13g2_dlygate4sd3_1 hold1527 (.A(_01402_),
    .X(net2590));
 sg13g2_dlygate4sd3_1 hold1528 (.A(\u_inv.d_next[226] ),
    .X(net2591));
 sg13g2_dlygate4sd3_1 hold1529 (.A(\perf_triple[7] ),
    .X(net2592));
 sg13g2_dlygate4sd3_1 hold1530 (.A(\u_inv.f_reg[187] ),
    .X(net2593));
 sg13g2_dlygate4sd3_1 hold1531 (.A(_01694_),
    .X(net2594));
 sg13g2_dlygate4sd3_1 hold1532 (.A(\u_inv.f_next[140] ),
    .X(net2595));
 sg13g2_dlygate4sd3_1 hold1533 (.A(\shift_reg[32] ),
    .X(net2596));
 sg13g2_dlygate4sd3_1 hold1534 (.A(_00207_),
    .X(net2597));
 sg13g2_dlygate4sd3_1 hold1535 (.A(\u_inv.f_reg[47] ),
    .X(net2598));
 sg13g2_dlygate4sd3_1 hold1536 (.A(_01554_),
    .X(net2599));
 sg13g2_dlygate4sd3_1 hold1537 (.A(\u_inv.input_reg[136] ),
    .X(net2600));
 sg13g2_dlygate4sd3_1 hold1538 (.A(_00043_),
    .X(net2601));
 sg13g2_dlygate4sd3_1 hold1539 (.A(\u_inv.f_reg[164] ),
    .X(net2602));
 sg13g2_dlygate4sd3_1 hold1540 (.A(_01671_),
    .X(net2603));
 sg13g2_dlygate4sd3_1 hold1541 (.A(\shift_reg[196] ),
    .X(net2604));
 sg13g2_dlygate4sd3_1 hold1542 (.A(_00371_),
    .X(net2605));
 sg13g2_dlygate4sd3_1 hold1543 (.A(\u_inv.d_next[140] ),
    .X(net2606));
 sg13g2_dlygate4sd3_1 hold1544 (.A(_01390_),
    .X(net2607));
 sg13g2_dlygate4sd3_1 hold1545 (.A(\shift_reg[245] ),
    .X(net2608));
 sg13g2_dlygate4sd3_1 hold1546 (.A(_00420_),
    .X(net2609));
 sg13g2_dlygate4sd3_1 hold1547 (.A(wr_prev),
    .X(net2610));
 sg13g2_dlygate4sd3_1 hold1548 (.A(_18620_),
    .X(net2611));
 sg13g2_dlygate4sd3_1 hold1549 (.A(_24690_[0]),
    .X(net2612));
 sg13g2_dlygate4sd3_1 hold1550 (.A(\u_inv.d_reg[153] ),
    .X(net2613));
 sg13g2_dlygate4sd3_1 hold1551 (.A(\u_inv.d_next[58] ),
    .X(net2614));
 sg13g2_dlygate4sd3_1 hold1552 (.A(_01308_),
    .X(net2615));
 sg13g2_dlygate4sd3_1 hold1553 (.A(\u_inv.f_reg[172] ),
    .X(net2616));
 sg13g2_dlygate4sd3_1 hold1554 (.A(_01679_),
    .X(net2617));
 sg13g2_dlygate4sd3_1 hold1555 (.A(\shift_reg[254] ),
    .X(net2618));
 sg13g2_dlygate4sd3_1 hold1556 (.A(\shift_reg[265] ),
    .X(net2619));
 sg13g2_dlygate4sd3_1 hold1557 (.A(\u_inv.d_next[234] ),
    .X(net2620));
 sg13g2_dlygate4sd3_1 hold1558 (.A(\shift_reg[69] ),
    .X(net2621));
 sg13g2_dlygate4sd3_1 hold1559 (.A(_00244_),
    .X(net2622));
 sg13g2_dlygate4sd3_1 hold1560 (.A(\u_inv.f_reg[251] ),
    .X(net2623));
 sg13g2_dlygate4sd3_1 hold1561 (.A(_01758_),
    .X(net2624));
 sg13g2_dlygate4sd3_1 hold1562 (.A(\shift_reg[198] ),
    .X(net2625));
 sg13g2_dlygate4sd3_1 hold1563 (.A(\shift_reg[264] ),
    .X(net2626));
 sg13g2_dlygate4sd3_1 hold1564 (.A(_00439_),
    .X(net2627));
 sg13g2_dlygate4sd3_1 hold1565 (.A(\u_inv.f_reg[9] ),
    .X(net2628));
 sg13g2_dlygate4sd3_1 hold1566 (.A(_01516_),
    .X(net2629));
 sg13g2_dlygate4sd3_1 hold1567 (.A(\inv_result[71] ),
    .X(net2630));
 sg13g2_dlygate4sd3_1 hold1568 (.A(\shift_reg[230] ),
    .X(net2631));
 sg13g2_dlygate4sd3_1 hold1569 (.A(_00405_),
    .X(net2632));
 sg13g2_dlygate4sd3_1 hold1570 (.A(\u_inv.d_next[244] ),
    .X(net2633));
 sg13g2_dlygate4sd3_1 hold1571 (.A(\u_inv.f_next[217] ),
    .X(net2634));
 sg13g2_dlygate4sd3_1 hold1572 (.A(\u_inv.f_next[16] ),
    .X(net2635));
 sg13g2_dlygate4sd3_1 hold1573 (.A(\shift_reg[249] ),
    .X(net2636));
 sg13g2_dlygate4sd3_1 hold1574 (.A(\u_inv.d_reg[118] ),
    .X(net2637));
 sg13g2_dlygate4sd3_1 hold1575 (.A(\inv_result[53] ),
    .X(net2638));
 sg13g2_dlygate4sd3_1 hold1576 (.A(\u_inv.input_reg[169] ),
    .X(net2639));
 sg13g2_dlygate4sd3_1 hold1577 (.A(\u_inv.f_reg[160] ),
    .X(net2640));
 sg13g2_dlygate4sd3_1 hold1578 (.A(_01667_),
    .X(net2641));
 sg13g2_dlygate4sd3_1 hold1579 (.A(\u_inv.f_reg[240] ),
    .X(net2642));
 sg13g2_dlygate4sd3_1 hold1580 (.A(_01747_),
    .X(net2643));
 sg13g2_dlygate4sd3_1 hold1581 (.A(\inv_result[89] ),
    .X(net2644));
 sg13g2_dlygate4sd3_1 hold1582 (.A(\shift_reg[129] ),
    .X(net2645));
 sg13g2_dlygate4sd3_1 hold1583 (.A(\u_inv.d_next[35] ),
    .X(net2646));
 sg13g2_dlygate4sd3_1 hold1584 (.A(_01285_),
    .X(net2647));
 sg13g2_dlygate4sd3_1 hold1585 (.A(\inv_result[32] ),
    .X(net2648));
 sg13g2_dlygate4sd3_1 hold1586 (.A(\shift_reg[256] ),
    .X(net2649));
 sg13g2_dlygate4sd3_1 hold1587 (.A(_00431_),
    .X(net2650));
 sg13g2_dlygate4sd3_1 hold1588 (.A(\shift_reg[113] ),
    .X(net2651));
 sg13g2_dlygate4sd3_1 hold1589 (.A(_00288_),
    .X(net2652));
 sg13g2_dlygate4sd3_1 hold1590 (.A(\u_inv.f_next[51] ),
    .X(net2653));
 sg13g2_dlygate4sd3_1 hold1591 (.A(\u_inv.d_next[183] ),
    .X(net2654));
 sg13g2_dlygate4sd3_1 hold1592 (.A(_01433_),
    .X(net2655));
 sg13g2_dlygate4sd3_1 hold1593 (.A(\u_inv.f_reg[18] ),
    .X(net2656));
 sg13g2_dlygate4sd3_1 hold1594 (.A(_01525_),
    .X(net2657));
 sg13g2_dlygate4sd3_1 hold1595 (.A(\shift_reg[10] ),
    .X(net2658));
 sg13g2_dlygate4sd3_1 hold1596 (.A(\u_inv.f_reg[41] ),
    .X(net2659));
 sg13g2_dlygate4sd3_1 hold1597 (.A(\u_inv.f_reg[254] ),
    .X(net2660));
 sg13g2_dlygate4sd3_1 hold1598 (.A(_01761_),
    .X(net2661));
 sg13g2_dlygate4sd3_1 hold1599 (.A(\u_inv.d_next[46] ),
    .X(net2662));
 sg13g2_dlygate4sd3_1 hold1600 (.A(\u_inv.d_next[106] ),
    .X(net2663));
 sg13g2_dlygate4sd3_1 hold1601 (.A(_01356_),
    .X(net2664));
 sg13g2_dlygate4sd3_1 hold1602 (.A(\u_inv.d_next[109] ),
    .X(net2665));
 sg13g2_dlygate4sd3_1 hold1603 (.A(_01359_),
    .X(net2666));
 sg13g2_dlygate4sd3_1 hold1604 (.A(\u_inv.f_reg[127] ),
    .X(net2667));
 sg13g2_dlygate4sd3_1 hold1605 (.A(_01634_),
    .X(net2668));
 sg13g2_dlygate4sd3_1 hold1606 (.A(\u_inv.d_next[156] ),
    .X(net2669));
 sg13g2_dlygate4sd3_1 hold1607 (.A(_01406_),
    .X(net2670));
 sg13g2_dlygate4sd3_1 hold1608 (.A(\u_inv.d_next[238] ),
    .X(net2671));
 sg13g2_dlygate4sd3_1 hold1609 (.A(\perf_triple[4] ),
    .X(net2672));
 sg13g2_dlygate4sd3_1 hold1610 (.A(\u_inv.input_reg[223] ),
    .X(net2673));
 sg13g2_dlygate4sd3_1 hold1612 (.A(_18476_),
    .X(net2675));
 sg13g2_dlygate4sd3_1 hold1613 (.A(\u_inv.f_reg[191] ),
    .X(net2676));
 sg13g2_dlygate4sd3_1 hold1614 (.A(_01698_),
    .X(net2677));
 sg13g2_dlygate4sd3_1 hold1615 (.A(\shift_reg[186] ),
    .X(net2678));
 sg13g2_dlygate4sd3_1 hold1616 (.A(_00361_),
    .X(net2679));
 sg13g2_dlygate4sd3_1 hold1617 (.A(\u_inv.f_reg[244] ),
    .X(net2680));
 sg13g2_dlygate4sd3_1 hold1618 (.A(_01751_),
    .X(net2681));
 sg13g2_dlygate4sd3_1 hold1619 (.A(\shift_reg[253] ),
    .X(net2682));
 sg13g2_dlygate4sd3_1 hold1620 (.A(\u_inv.f_reg[98] ),
    .X(net2683));
 sg13g2_dlygate4sd3_1 hold1621 (.A(_01605_),
    .X(net2684));
 sg13g2_dlygate4sd3_1 hold1622 (.A(\u_inv.f_reg[42] ),
    .X(net2685));
 sg13g2_dlygate4sd3_1 hold1623 (.A(_01549_),
    .X(net2686));
 sg13g2_dlygate4sd3_1 hold1624 (.A(\u_inv.d_next[188] ),
    .X(net2687));
 sg13g2_dlygate4sd3_1 hold1625 (.A(\u_inv.f_reg[248] ),
    .X(net2688));
 sg13g2_dlygate4sd3_1 hold1626 (.A(_01755_),
    .X(net2689));
 sg13g2_dlygate4sd3_1 hold1627 (.A(\shift_reg[248] ),
    .X(net2690));
 sg13g2_dlygate4sd3_1 hold1628 (.A(\u_inv.d_next[200] ),
    .X(net2691));
 sg13g2_dlygate4sd3_1 hold1629 (.A(_01450_),
    .X(net2692));
 sg13g2_dlygate4sd3_1 hold1630 (.A(\u_inv.d_next[202] ),
    .X(net2693));
 sg13g2_dlygate4sd3_1 hold1631 (.A(\u_inv.d_next[146] ),
    .X(net2694));
 sg13g2_dlygate4sd3_1 hold1632 (.A(\u_inv.f_reg[222] ),
    .X(net2695));
 sg13g2_dlygate4sd3_1 hold1633 (.A(_01729_),
    .X(net2696));
 sg13g2_dlygate4sd3_1 hold1634 (.A(\u_inv.f_reg[243] ),
    .X(net2697));
 sg13g2_dlygate4sd3_1 hold1635 (.A(\shift_reg[214] ),
    .X(net2698));
 sg13g2_dlygate4sd3_1 hold1636 (.A(\u_inv.f_reg[218] ),
    .X(net2699));
 sg13g2_dlygate4sd3_1 hold1637 (.A(_01725_),
    .X(net2700));
 sg13g2_dlygate4sd3_1 hold1638 (.A(\shift_reg[80] ),
    .X(net2701));
 sg13g2_dlygate4sd3_1 hold1639 (.A(_00255_),
    .X(net2702));
 sg13g2_dlygate4sd3_1 hold1640 (.A(\u_inv.d_next[0] ),
    .X(net2703));
 sg13g2_dlygate4sd3_1 hold1641 (.A(_01250_),
    .X(net2704));
 sg13g2_dlygate4sd3_1 hold1642 (.A(\u_inv.d_next[36] ),
    .X(net2705));
 sg13g2_dlygate4sd3_1 hold1643 (.A(_01286_),
    .X(net2706));
 sg13g2_dlygate4sd3_1 hold1644 (.A(\u_inv.d_next[177] ),
    .X(net2707));
 sg13g2_dlygate4sd3_1 hold1645 (.A(_01427_),
    .X(net2708));
 sg13g2_dlygate4sd3_1 hold1646 (.A(\u_inv.f_reg[108] ),
    .X(net2709));
 sg13g2_dlygate4sd3_1 hold1647 (.A(_01615_),
    .X(net2710));
 sg13g2_dlygate4sd3_1 hold1648 (.A(\inv_result[65] ),
    .X(net2711));
 sg13g2_dlygate4sd3_1 hold1649 (.A(\u_inv.d_next[164] ),
    .X(net2712));
 sg13g2_dlygate4sd3_1 hold1650 (.A(_01414_),
    .X(net2713));
 sg13g2_dlygate4sd3_1 hold1651 (.A(\u_inv.f_reg[134] ),
    .X(net2714));
 sg13g2_dlygate4sd3_1 hold1652 (.A(_01641_),
    .X(net2715));
 sg13g2_dlygate4sd3_1 hold1653 (.A(\u_inv.f_next[180] ),
    .X(net2716));
 sg13g2_dlygate4sd3_1 hold1654 (.A(\inv_result[140] ),
    .X(net2717));
 sg13g2_dlygate4sd3_1 hold1655 (.A(\u_inv.input_reg[207] ),
    .X(net2718));
 sg13g2_dlygate4sd3_1 hold1656 (.A(_00114_),
    .X(net2719));
 sg13g2_dlygate4sd3_1 hold1657 (.A(\u_inv.d_reg[170] ),
    .X(net2720));
 sg13g2_dlygate4sd3_1 hold1658 (.A(\u_inv.d_next[207] ),
    .X(net2721));
 sg13g2_dlygate4sd3_1 hold1659 (.A(_01457_),
    .X(net2722));
 sg13g2_dlygate4sd3_1 hold1660 (.A(\inv_result[248] ),
    .X(net2723));
 sg13g2_dlygate4sd3_1 hold1661 (.A(\u_inv.f_reg[242] ),
    .X(net2724));
 sg13g2_dlygate4sd3_1 hold1662 (.A(_01749_),
    .X(net2725));
 sg13g2_dlygate4sd3_1 hold1663 (.A(\u_inv.d_next[144] ),
    .X(net2726));
 sg13g2_dlygate4sd3_1 hold1664 (.A(_01394_),
    .X(net2727));
 sg13g2_dlygate4sd3_1 hold1665 (.A(\shift_reg[219] ),
    .X(net2728));
 sg13g2_dlygate4sd3_1 hold1666 (.A(_00394_),
    .X(net2729));
 sg13g2_dlygate4sd3_1 hold1667 (.A(\u_inv.f_next[256] ),
    .X(net2730));
 sg13g2_dlygate4sd3_1 hold1668 (.A(\u_inv.d_reg[81] ),
    .X(net2731));
 sg13g2_dlygate4sd3_1 hold1669 (.A(_01331_),
    .X(net2732));
 sg13g2_dlygate4sd3_1 hold1670 (.A(\shift_reg[50] ),
    .X(net2733));
 sg13g2_dlygate4sd3_1 hold1671 (.A(_00225_),
    .X(net2734));
 sg13g2_dlygate4sd3_1 hold1672 (.A(\u_inv.f_next[98] ),
    .X(net2735));
 sg13g2_dlygate4sd3_1 hold1673 (.A(\u_inv.d_next[7] ),
    .X(net2736));
 sg13g2_dlygate4sd3_1 hold1674 (.A(_01257_),
    .X(net2737));
 sg13g2_dlygate4sd3_1 hold1675 (.A(\u_inv.f_reg[74] ),
    .X(net2738));
 sg13g2_dlygate4sd3_1 hold1676 (.A(_01581_),
    .X(net2739));
 sg13g2_dlygate4sd3_1 hold1677 (.A(\u_inv.f_reg[86] ),
    .X(net2740));
 sg13g2_dlygate4sd3_1 hold1678 (.A(_01593_),
    .X(net2741));
 sg13g2_dlygate4sd3_1 hold1679 (.A(\shift_reg[234] ),
    .X(net2742));
 sg13g2_dlygate4sd3_1 hold1680 (.A(_00409_),
    .X(net2743));
 sg13g2_dlygate4sd3_1 hold1681 (.A(\u_inv.d_next[142] ),
    .X(net2744));
 sg13g2_dlygate4sd3_1 hold1682 (.A(\u_inv.d_reg[225] ),
    .X(net2745));
 sg13g2_dlygate4sd3_1 hold1683 (.A(\u_inv.d_next[82] ),
    .X(net2746));
 sg13g2_dlygate4sd3_1 hold1684 (.A(_01332_),
    .X(net2747));
 sg13g2_dlygate4sd3_1 hold1685 (.A(\u_inv.f_reg[152] ),
    .X(net2748));
 sg13g2_dlygate4sd3_1 hold1686 (.A(_01659_),
    .X(net2749));
 sg13g2_dlygate4sd3_1 hold1687 (.A(\shift_reg[155] ),
    .X(net2750));
 sg13g2_dlygate4sd3_1 hold1688 (.A(_00330_),
    .X(net2751));
 sg13g2_dlygate4sd3_1 hold1689 (.A(\inv_result[59] ),
    .X(net2752));
 sg13g2_dlygate4sd3_1 hold1690 (.A(\u_inv.f_reg[213] ),
    .X(net2753));
 sg13g2_dlygate4sd3_1 hold1691 (.A(_01720_),
    .X(net2754));
 sg13g2_dlygate4sd3_1 hold1692 (.A(\shift_reg[207] ),
    .X(net2755));
 sg13g2_dlygate4sd3_1 hold1693 (.A(\u_inv.f_next[209] ),
    .X(net2756));
 sg13g2_dlygate4sd3_1 hold1694 (.A(\inv_result[206] ),
    .X(net2757));
 sg13g2_dlygate4sd3_1 hold1695 (.A(\u_inv.f_next[129] ),
    .X(net2758));
 sg13g2_dlygate4sd3_1 hold1696 (.A(\u_inv.input_reg[201] ),
    .X(net2759));
 sg13g2_dlygate4sd3_1 hold1697 (.A(\u_inv.f_next[32] ),
    .X(net2760));
 sg13g2_dlygate4sd3_1 hold1698 (.A(_01539_),
    .X(net2761));
 sg13g2_dlygate4sd3_1 hold1699 (.A(\u_inv.d_next[38] ),
    .X(net2762));
 sg13g2_dlygate4sd3_1 hold1700 (.A(_01288_),
    .X(net2763));
 sg13g2_dlygate4sd3_1 hold1701 (.A(\u_inv.d_next[37] ),
    .X(net2764));
 sg13g2_dlygate4sd3_1 hold1702 (.A(_01287_),
    .X(net2765));
 sg13g2_dlygate4sd3_1 hold1703 (.A(\u_inv.f_reg[128] ),
    .X(net2766));
 sg13g2_dlygate4sd3_1 hold1704 (.A(_01635_),
    .X(net2767));
 sg13g2_dlygate4sd3_1 hold1705 (.A(\u_inv.f_reg[148] ),
    .X(net2768));
 sg13g2_dlygate4sd3_1 hold1706 (.A(_01655_),
    .X(net2769));
 sg13g2_dlygate4sd3_1 hold1707 (.A(\shift_reg[57] ),
    .X(net2770));
 sg13g2_dlygate4sd3_1 hold1708 (.A(_00232_),
    .X(net2771));
 sg13g2_dlygate4sd3_1 hold1709 (.A(\u_inv.d_next[201] ),
    .X(net2772));
 sg13g2_dlygate4sd3_1 hold1710 (.A(_01451_),
    .X(net2773));
 sg13g2_dlygate4sd3_1 hold1711 (.A(\u_inv.f_next[6] ),
    .X(net2774));
 sg13g2_dlygate4sd3_1 hold1712 (.A(\u_inv.d_reg[55] ),
    .X(net2775));
 sg13g2_dlygate4sd3_1 hold1713 (.A(\u_inv.f_reg[71] ),
    .X(net2776));
 sg13g2_dlygate4sd3_1 hold1714 (.A(_01578_),
    .X(net2777));
 sg13g2_dlygate4sd3_1 hold1715 (.A(\shift_reg[23] ),
    .X(net2778));
 sg13g2_dlygate4sd3_1 hold1716 (.A(_00198_),
    .X(net2779));
 sg13g2_dlygate4sd3_1 hold1717 (.A(\u_inv.f_next[21] ),
    .X(net2780));
 sg13g2_dlygate4sd3_1 hold1718 (.A(\shift_reg[44] ),
    .X(net2781));
 sg13g2_dlygate4sd3_1 hold1719 (.A(_00219_),
    .X(net2782));
 sg13g2_dlygate4sd3_1 hold1720 (.A(\u_inv.f_next[40] ),
    .X(net2783));
 sg13g2_dlygate4sd3_1 hold1721 (.A(\shift_reg[201] ),
    .X(net2784));
 sg13g2_dlygate4sd3_1 hold1722 (.A(\u_inv.input_reg[203] ),
    .X(net2785));
 sg13g2_dlygate4sd3_1 hold1723 (.A(\u_inv.d_next[230] ),
    .X(net2786));
 sg13g2_dlygate4sd3_1 hold1724 (.A(\u_inv.d_next[211] ),
    .X(net2787));
 sg13g2_dlygate4sd3_1 hold1725 (.A(_01461_),
    .X(net2788));
 sg13g2_dlygate4sd3_1 hold1726 (.A(\u_inv.f_reg[178] ),
    .X(net2789));
 sg13g2_dlygate4sd3_1 hold1727 (.A(_01685_),
    .X(net2790));
 sg13g2_dlygate4sd3_1 hold1728 (.A(\u_inv.input_reg[146] ),
    .X(net2791));
 sg13g2_dlygate4sd3_1 hold1729 (.A(_00053_),
    .X(net2792));
 sg13g2_dlygate4sd3_1 hold1730 (.A(\shift_reg[179] ),
    .X(net2793));
 sg13g2_dlygate4sd3_1 hold1731 (.A(_00354_),
    .X(net2794));
 sg13g2_dlygate4sd3_1 hold1732 (.A(\u_inv.f_reg[182] ),
    .X(net2795));
 sg13g2_dlygate4sd3_1 hold1733 (.A(_01689_),
    .X(net2796));
 sg13g2_dlygate4sd3_1 hold1734 (.A(\u_inv.d_next[15] ),
    .X(net2797));
 sg13g2_dlygate4sd3_1 hold1735 (.A(_01265_),
    .X(net2798));
 sg13g2_dlygate4sd3_1 hold1736 (.A(\shift_reg[260] ),
    .X(net2799));
 sg13g2_dlygate4sd3_1 hold1737 (.A(\shift_reg[235] ),
    .X(net2800));
 sg13g2_dlygate4sd3_1 hold1738 (.A(_00410_),
    .X(net2801));
 sg13g2_dlygate4sd3_1 hold1739 (.A(\shift_reg[33] ),
    .X(net2802));
 sg13g2_dlygate4sd3_1 hold1740 (.A(_00208_),
    .X(net2803));
 sg13g2_dlygate4sd3_1 hold1741 (.A(\u_inv.d_next[71] ),
    .X(net2804));
 sg13g2_dlygate4sd3_1 hold1742 (.A(\u_inv.d_next[6] ),
    .X(net2805));
 sg13g2_dlygate4sd3_1 hold1743 (.A(_01256_),
    .X(net2806));
 sg13g2_dlygate4sd3_1 hold1744 (.A(\u_inv.d_next[12] ),
    .X(net2807));
 sg13g2_dlygate4sd3_1 hold1745 (.A(_01262_),
    .X(net2808));
 sg13g2_dlygate4sd3_1 hold1746 (.A(\u_inv.d_next[251] ),
    .X(net2809));
 sg13g2_dlygate4sd3_1 hold1747 (.A(\u_inv.f_reg[63] ),
    .X(net2810));
 sg13g2_dlygate4sd3_1 hold1748 (.A(_01570_),
    .X(net2811));
 sg13g2_dlygate4sd3_1 hold1749 (.A(\u_inv.f_reg[103] ),
    .X(net2812));
 sg13g2_dlygate4sd3_1 hold1750 (.A(_01610_),
    .X(net2813));
 sg13g2_dlygate4sd3_1 hold1751 (.A(\u_inv.d_next[65] ),
    .X(net2814));
 sg13g2_dlygate4sd3_1 hold1752 (.A(_01315_),
    .X(net2815));
 sg13g2_dlygate4sd3_1 hold1753 (.A(\shift_reg[82] ),
    .X(net2816));
 sg13g2_dlygate4sd3_1 hold1754 (.A(_00257_),
    .X(net2817));
 sg13g2_dlygate4sd3_1 hold1755 (.A(\u_inv.f_next[233] ),
    .X(net2818));
 sg13g2_dlygate4sd3_1 hold1756 (.A(\u_inv.d_next[4] ),
    .X(net2819));
 sg13g2_dlygate4sd3_1 hold1757 (.A(_01254_),
    .X(net2820));
 sg13g2_dlygate4sd3_1 hold1758 (.A(\u_inv.f_next[101] ),
    .X(net2821));
 sg13g2_dlygate4sd3_1 hold1759 (.A(\shift_reg[48] ),
    .X(net2822));
 sg13g2_dlygate4sd3_1 hold1760 (.A(_00223_),
    .X(net2823));
 sg13g2_dlygate4sd3_1 hold1761 (.A(\u_inv.d_next[205] ),
    .X(net2824));
 sg13g2_dlygate4sd3_1 hold1762 (.A(_01455_),
    .X(net2825));
 sg13g2_dlygate4sd3_1 hold1763 (.A(\u_inv.d_next[136] ),
    .X(net2826));
 sg13g2_dlygate4sd3_1 hold1764 (.A(_01386_),
    .X(net2827));
 sg13g2_dlygate4sd3_1 hold1765 (.A(\shift_reg[14] ),
    .X(net2828));
 sg13g2_dlygate4sd3_1 hold1766 (.A(_00189_),
    .X(net2829));
 sg13g2_dlygate4sd3_1 hold1767 (.A(\u_inv.f_next[179] ),
    .X(net2830));
 sg13g2_dlygate4sd3_1 hold1768 (.A(\u_inv.f_reg[180] ),
    .X(net2831));
 sg13g2_dlygate4sd3_1 hold1769 (.A(\u_inv.f_next[33] ),
    .X(net2832));
 sg13g2_dlygate4sd3_1 hold1770 (.A(\u_inv.d_reg[204] ),
    .X(net2833));
 sg13g2_dlygate4sd3_1 hold1771 (.A(\u_inv.d_reg[190] ),
    .X(net2834));
 sg13g2_dlygate4sd3_1 hold1772 (.A(\u_inv.d_next[145] ),
    .X(net2835));
 sg13g2_dlygate4sd3_1 hold1773 (.A(_01395_),
    .X(net2836));
 sg13g2_dlygate4sd3_1 hold1774 (.A(\u_inv.d_reg[174] ),
    .X(net2837));
 sg13g2_dlygate4sd3_1 hold1775 (.A(\inv_result[57] ),
    .X(net2838));
 sg13g2_dlygate4sd3_1 hold1776 (.A(\u_inv.f_reg[13] ),
    .X(net2839));
 sg13g2_dlygate4sd3_1 hold1777 (.A(_01520_),
    .X(net2840));
 sg13g2_dlygate4sd3_1 hold1778 (.A(\u_inv.f_reg[53] ),
    .X(net2841));
 sg13g2_dlygate4sd3_1 hold1779 (.A(_01560_),
    .X(net2842));
 sg13g2_dlygate4sd3_1 hold1780 (.A(\u_inv.f_next[207] ),
    .X(net2843));
 sg13g2_dlygate4sd3_1 hold1781 (.A(\u_inv.f_next[121] ),
    .X(net2844));
 sg13g2_dlygate4sd3_1 hold1782 (.A(\u_inv.f_next[17] ),
    .X(net2845));
 sg13g2_dlygate4sd3_1 hold1783 (.A(\u_inv.f_next[93] ),
    .X(net2846));
 sg13g2_dlygate4sd3_1 hold1784 (.A(\shift_reg[192] ),
    .X(net2847));
 sg13g2_dlygate4sd3_1 hold1785 (.A(\u_inv.f_next[167] ),
    .X(net2848));
 sg13g2_dlygate4sd3_1 hold1786 (.A(\shift_reg[200] ),
    .X(net2849));
 sg13g2_dlygate4sd3_1 hold1787 (.A(\u_inv.f_next[183] ),
    .X(net2850));
 sg13g2_dlygate4sd3_1 hold1788 (.A(\trng_data[0] ),
    .X(net2851));
 sg13g2_dlygate4sd3_1 hold1789 (.A(_00449_),
    .X(net2852));
 sg13g2_dlygate4sd3_1 hold1790 (.A(\shift_reg[100] ),
    .X(net2853));
 sg13g2_dlygate4sd3_1 hold1791 (.A(_00275_),
    .X(net2854));
 sg13g2_dlygate4sd3_1 hold1792 (.A(\u_inv.f_reg[230] ),
    .X(net2855));
 sg13g2_dlygate4sd3_1 hold1793 (.A(_01737_),
    .X(net2856));
 sg13g2_dlygate4sd3_1 hold1794 (.A(\u_inv.f_reg[249] ),
    .X(net2857));
 sg13g2_dlygate4sd3_1 hold1795 (.A(_01756_),
    .X(net2858));
 sg13g2_dlygate4sd3_1 hold1796 (.A(\inv_result[66] ),
    .X(net2859));
 sg13g2_dlygate4sd3_1 hold1797 (.A(\shift_reg[267] ),
    .X(net2860));
 sg13g2_dlygate4sd3_1 hold1798 (.A(_00442_),
    .X(net2861));
 sg13g2_dlygate4sd3_1 hold1799 (.A(\u_inv.d_next[104] ),
    .X(net2862));
 sg13g2_dlygate4sd3_1 hold1800 (.A(_01354_),
    .X(net2863));
 sg13g2_dlygate4sd3_1 hold1801 (.A(\u_inv.f_reg[168] ),
    .X(net2864));
 sg13g2_dlygate4sd3_1 hold1802 (.A(_01675_),
    .X(net2865));
 sg13g2_dlygate4sd3_1 hold1803 (.A(\u_inv.f_reg[197] ),
    .X(net2866));
 sg13g2_dlygate4sd3_1 hold1804 (.A(_01704_),
    .X(net2867));
 sg13g2_dlygate4sd3_1 hold1805 (.A(\inv_result[247] ),
    .X(net2868));
 sg13g2_dlygate4sd3_1 hold1806 (.A(\u_inv.d_next[107] ),
    .X(net2869));
 sg13g2_dlygate4sd3_1 hold1807 (.A(_01357_),
    .X(net2870));
 sg13g2_dlygate4sd3_1 hold1808 (.A(\u_inv.d_next[210] ),
    .X(net2871));
 sg13g2_dlygate4sd3_1 hold1809 (.A(_01460_),
    .X(net2872));
 sg13g2_dlygate4sd3_1 hold1810 (.A(\inv_result[58] ),
    .X(net2873));
 sg13g2_dlygate4sd3_1 hold1811 (.A(\u_inv.f_next[235] ),
    .X(net2874));
 sg13g2_dlygate4sd3_1 hold1812 (.A(\u_inv.f_reg[54] ),
    .X(net2875));
 sg13g2_dlygate4sd3_1 hold1813 (.A(_01561_),
    .X(net2876));
 sg13g2_dlygate4sd3_1 hold1814 (.A(\u_inv.d_next[117] ),
    .X(net2877));
 sg13g2_dlygate4sd3_1 hold1815 (.A(_01367_),
    .X(net2878));
 sg13g2_dlygate4sd3_1 hold1816 (.A(\u_inv.f_next[56] ),
    .X(net2879));
 sg13g2_dlygate4sd3_1 hold1817 (.A(\u_inv.d_next[250] ),
    .X(net2880));
 sg13g2_dlygate4sd3_1 hold1818 (.A(\u_inv.f_reg[153] ),
    .X(net2881));
 sg13g2_dlygate4sd3_1 hold1819 (.A(_01660_),
    .X(net2882));
 sg13g2_dlygate4sd3_1 hold1820 (.A(\u_inv.f_next[184] ),
    .X(net2883));
 sg13g2_dlygate4sd3_1 hold1821 (.A(\u_inv.f_reg[232] ),
    .X(net2884));
 sg13g2_dlygate4sd3_1 hold1822 (.A(_01739_),
    .X(net2885));
 sg13g2_dlygate4sd3_1 hold1823 (.A(\u_inv.d_next[154] ),
    .X(net2886));
 sg13g2_dlygate4sd3_1 hold1824 (.A(_01404_),
    .X(net2887));
 sg13g2_dlygate4sd3_1 hold1825 (.A(\u_inv.d_next[254] ),
    .X(net2888));
 sg13g2_dlygate4sd3_1 hold1826 (.A(_01504_),
    .X(net2889));
 sg13g2_dlygate4sd3_1 hold1827 (.A(\u_inv.d_next[119] ),
    .X(net2890));
 sg13g2_dlygate4sd3_1 hold1828 (.A(_01369_),
    .X(net2891));
 sg13g2_dlygate4sd3_1 hold1829 (.A(\u_inv.input_reg[149] ),
    .X(net2892));
 sg13g2_dlygate4sd3_1 hold1830 (.A(_00056_),
    .X(net2893));
 sg13g2_dlygate4sd3_1 hold1831 (.A(\u_inv.d_reg[250] ),
    .X(net2894));
 sg13g2_dlygate4sd3_1 hold1832 (.A(\u_inv.d_reg[85] ),
    .X(net2895));
 sg13g2_dlygate4sd3_1 hold1833 (.A(\u_inv.f_reg[23] ),
    .X(net2896));
 sg13g2_dlygate4sd3_1 hold1834 (.A(_01530_),
    .X(net2897));
 sg13g2_dlygate4sd3_1 hold1835 (.A(\shift_reg[157] ),
    .X(net2898));
 sg13g2_dlygate4sd3_1 hold1836 (.A(_00332_),
    .X(net2899));
 sg13g2_dlygate4sd3_1 hold1837 (.A(\shift_reg[65] ),
    .X(net2900));
 sg13g2_dlygate4sd3_1 hold1838 (.A(_00240_),
    .X(net2901));
 sg13g2_dlygate4sd3_1 hold1839 (.A(\u_inv.f_reg[228] ),
    .X(net2902));
 sg13g2_dlygate4sd3_1 hold1840 (.A(_01735_),
    .X(net2903));
 sg13g2_dlygate4sd3_1 hold1841 (.A(\u_inv.f_reg[149] ),
    .X(net2904));
 sg13g2_dlygate4sd3_1 hold1842 (.A(_01656_),
    .X(net2905));
 sg13g2_dlygate4sd3_1 hold1843 (.A(\u_inv.f_reg[161] ),
    .X(net2906));
 sg13g2_dlygate4sd3_1 hold1844 (.A(_01668_),
    .X(net2907));
 sg13g2_dlygate4sd3_1 hold1845 (.A(\u_inv.f_reg[239] ),
    .X(net2908));
 sg13g2_dlygate4sd3_1 hold1846 (.A(_01746_),
    .X(net2909));
 sg13g2_dlygate4sd3_1 hold1847 (.A(\u_inv.d_next[54] ),
    .X(net2910));
 sg13g2_dlygate4sd3_1 hold1848 (.A(_01304_),
    .X(net2911));
 sg13g2_dlygate4sd3_1 hold1849 (.A(\shift_reg[84] ),
    .X(net2912));
 sg13g2_dlygate4sd3_1 hold1850 (.A(_00259_),
    .X(net2913));
 sg13g2_dlygate4sd3_1 hold1851 (.A(\shift_reg[114] ),
    .X(net2914));
 sg13g2_dlygate4sd3_1 hold1852 (.A(_00289_),
    .X(net2915));
 sg13g2_dlygate4sd3_1 hold1853 (.A(\u_inv.d_next[49] ),
    .X(net2916));
 sg13g2_dlygate4sd3_1 hold1854 (.A(\u_inv.f_reg[106] ),
    .X(net2917));
 sg13g2_dlygate4sd3_1 hold1855 (.A(_01613_),
    .X(net2918));
 sg13g2_dlygate4sd3_1 hold1856 (.A(\u_inv.f_reg[233] ),
    .X(net2919));
 sg13g2_dlygate4sd3_1 hold1857 (.A(\u_inv.d_next[214] ),
    .X(net2920));
 sg13g2_dlygate4sd3_1 hold1858 (.A(_01464_),
    .X(net2921));
 sg13g2_dlygate4sd3_1 hold1859 (.A(\u_inv.d_next[206] ),
    .X(net2922));
 sg13g2_dlygate4sd3_1 hold1860 (.A(\shift_reg[118] ),
    .X(net2923));
 sg13g2_dlygate4sd3_1 hold1861 (.A(_00293_),
    .X(net2924));
 sg13g2_dlygate4sd3_1 hold1862 (.A(\u_inv.d_next[192] ),
    .X(net2925));
 sg13g2_dlygate4sd3_1 hold1863 (.A(_01442_),
    .X(net2926));
 sg13g2_dlygate4sd3_1 hold1864 (.A(\u_inv.f_next[171] ),
    .X(net2927));
 sg13g2_dlygate4sd3_1 hold1865 (.A(\shift_reg[269] ),
    .X(net2928));
 sg13g2_dlygate4sd3_1 hold1866 (.A(_00444_),
    .X(net2929));
 sg13g2_dlygate4sd3_1 hold1867 (.A(\shift_reg[36] ),
    .X(net2930));
 sg13g2_dlygate4sd3_1 hold1868 (.A(_00211_),
    .X(net2931));
 sg13g2_dlygate4sd3_1 hold1869 (.A(\u_inv.d_reg[188] ),
    .X(net2932));
 sg13g2_dlygate4sd3_1 hold1870 (.A(\shift_reg[58] ),
    .X(net2933));
 sg13g2_dlygate4sd3_1 hold1871 (.A(\shift_reg[101] ),
    .X(net2934));
 sg13g2_dlygate4sd3_1 hold1872 (.A(_00276_),
    .X(net2935));
 sg13g2_dlygate4sd3_1 hold1873 (.A(\inv_result[81] ),
    .X(net2936));
 sg13g2_dlygate4sd3_1 hold1874 (.A(\u_inv.f_next[218] ),
    .X(net2937));
 sg13g2_dlygate4sd3_1 hold1875 (.A(\u_inv.f_next[119] ),
    .X(net2938));
 sg13g2_dlygate4sd3_1 hold1876 (.A(\u_inv.f_next[90] ),
    .X(net2939));
 sg13g2_dlygate4sd3_1 hold1877 (.A(\u_inv.d_reg[184] ),
    .X(net2940));
 sg13g2_dlygate4sd3_1 hold1878 (.A(\u_inv.f_reg[43] ),
    .X(net2941));
 sg13g2_dlygate4sd3_1 hold1879 (.A(_01550_),
    .X(net2942));
 sg13g2_dlygate4sd3_1 hold1880 (.A(\u_inv.f_reg[212] ),
    .X(net2943));
 sg13g2_dlygate4sd3_1 hold1881 (.A(_01719_),
    .X(net2944));
 sg13g2_dlygate4sd3_1 hold1882 (.A(\u_inv.d_next[14] ),
    .X(net2945));
 sg13g2_dlygate4sd3_1 hold1883 (.A(_01264_),
    .X(net2946));
 sg13g2_dlygate4sd3_1 hold1884 (.A(\u_inv.f_next[227] ),
    .X(net2947));
 sg13g2_dlygate4sd3_1 hold1885 (.A(\u_inv.d_next[25] ),
    .X(net2948));
 sg13g2_dlygate4sd3_1 hold1886 (.A(_01275_),
    .X(net2949));
 sg13g2_dlygate4sd3_1 hold1887 (.A(\u_inv.d_next[155] ),
    .X(net2950));
 sg13g2_dlygate4sd3_1 hold1888 (.A(_01405_),
    .X(net2951));
 sg13g2_dlygate4sd3_1 hold1889 (.A(\u_inv.f_reg[175] ),
    .X(net2952));
 sg13g2_dlygate4sd3_1 hold1890 (.A(\shift_reg[51] ),
    .X(net2953));
 sg13g2_dlygate4sd3_1 hold1891 (.A(_00226_),
    .X(net2954));
 sg13g2_dlygate4sd3_1 hold1892 (.A(\u_inv.f_reg[122] ),
    .X(net2955));
 sg13g2_dlygate4sd3_1 hold1893 (.A(_01629_),
    .X(net2956));
 sg13g2_dlygate4sd3_1 hold1894 (.A(\shift_reg[202] ),
    .X(net2957));
 sg13g2_dlygate4sd3_1 hold1895 (.A(\u_inv.f_reg[200] ),
    .X(net2958));
 sg13g2_dlygate4sd3_1 hold1896 (.A(_01707_),
    .X(net2959));
 sg13g2_dlygate4sd3_1 hold1897 (.A(\u_inv.f_reg[217] ),
    .X(net2960));
 sg13g2_dlygate4sd3_1 hold1898 (.A(\shift_reg[220] ),
    .X(net2961));
 sg13g2_dlygate4sd3_1 hold1899 (.A(_00395_),
    .X(net2962));
 sg13g2_dlygate4sd3_1 hold1900 (.A(\u_inv.d_reg[234] ),
    .X(net2963));
 sg13g2_dlygate4sd3_1 hold1901 (.A(\u_inv.f_next[97] ),
    .X(net2964));
 sg13g2_dlygate4sd3_1 hold1902 (.A(\shift_reg[130] ),
    .X(net2965));
 sg13g2_dlygate4sd3_1 hold1903 (.A(\u_inv.f_reg[220] ),
    .X(net2966));
 sg13g2_dlygate4sd3_1 hold1904 (.A(_01727_),
    .X(net2967));
 sg13g2_dlygate4sd3_1 hold1905 (.A(\u_inv.d_next[17] ),
    .X(net2968));
 sg13g2_dlygate4sd3_1 hold1906 (.A(\u_inv.input_reg[137] ),
    .X(net2969));
 sg13g2_dlygate4sd3_1 hold1907 (.A(_00044_),
    .X(net2970));
 sg13g2_dlygate4sd3_1 hold1908 (.A(\u_inv.d_reg[46] ),
    .X(net2971));
 sg13g2_dlygate4sd3_1 hold1909 (.A(\u_inv.d_next[98] ),
    .X(net2972));
 sg13g2_dlygate4sd3_1 hold1910 (.A(_01348_),
    .X(net2973));
 sg13g2_dlygate4sd3_1 hold1911 (.A(\u_inv.d_next[3] ),
    .X(net2974));
 sg13g2_dlygate4sd3_1 hold1912 (.A(_01253_),
    .X(net2975));
 sg13g2_dlygate4sd3_1 hold1913 (.A(\byte_cnt[0] ),
    .X(net2976));
 sg13g2_dlygate4sd3_1 hold1914 (.A(\u_inv.d_next[10] ),
    .X(net2977));
 sg13g2_dlygate4sd3_1 hold1915 (.A(_01260_),
    .X(net2978));
 sg13g2_dlygate4sd3_1 hold1916 (.A(\u_inv.d_next[59] ),
    .X(net2979));
 sg13g2_dlygate4sd3_1 hold1917 (.A(\u_inv.d_next[116] ),
    .X(net2980));
 sg13g2_dlygate4sd3_1 hold1918 (.A(_01366_),
    .X(net2981));
 sg13g2_dlygate4sd3_1 hold1919 (.A(\shift_reg[261] ),
    .X(net2982));
 sg13g2_dlygate4sd3_1 hold1920 (.A(_00436_),
    .X(net2983));
 sg13g2_dlygate4sd3_1 hold1921 (.A(\u_inv.f_reg[203] ),
    .X(net2984));
 sg13g2_dlygate4sd3_1 hold1922 (.A(_01710_),
    .X(net2985));
 sg13g2_dlygate4sd3_1 hold1923 (.A(\u_inv.d_next[105] ),
    .X(net2986));
 sg13g2_dlygate4sd3_1 hold1924 (.A(_01355_),
    .X(net2987));
 sg13g2_dlygate4sd3_1 hold1925 (.A(\u_inv.d_next[256] ),
    .X(net2988));
 sg13g2_dlygate4sd3_1 hold1926 (.A(\u_inv.d_next[224] ),
    .X(net2989));
 sg13g2_dlygate4sd3_1 hold1927 (.A(_01474_),
    .X(net2990));
 sg13g2_dlygate4sd3_1 hold1928 (.A(\u_inv.d_next[166] ),
    .X(net2991));
 sg13g2_dlygate4sd3_1 hold1929 (.A(\u_inv.d_next[102] ),
    .X(net2992));
 sg13g2_dlygate4sd3_1 hold1930 (.A(\shift_reg[91] ),
    .X(net2993));
 sg13g2_dlygate4sd3_1 hold1931 (.A(\shift_reg[81] ),
    .X(net2994));
 sg13g2_dlygate4sd3_1 hold1932 (.A(_00256_),
    .X(net2995));
 sg13g2_dlygate4sd3_1 hold1933 (.A(\u_inv.f_reg[157] ),
    .X(net2996));
 sg13g2_dlygate4sd3_1 hold1934 (.A(_01664_),
    .X(net2997));
 sg13g2_dlygate4sd3_1 hold1935 (.A(\u_inv.input_reg[126] ),
    .X(net2998));
 sg13g2_dlygate4sd3_1 hold1936 (.A(_00033_),
    .X(net2999));
 sg13g2_dlygate4sd3_1 hold1937 (.A(\u_inv.f_next[156] ),
    .X(net3000));
 sg13g2_dlygate4sd3_1 hold1938 (.A(\shift_reg[132] ),
    .X(net3001));
 sg13g2_dlygate4sd3_1 hold1939 (.A(\shift_reg[212] ),
    .X(net3002));
 sg13g2_dlygate4sd3_1 hold1940 (.A(_00387_),
    .X(net3003));
 sg13g2_dlygate4sd3_1 hold1941 (.A(\u_inv.f_reg[75] ),
    .X(net3004));
 sg13g2_dlygate4sd3_1 hold1942 (.A(_01582_),
    .X(net3005));
 sg13g2_dlygate4sd3_1 hold1943 (.A(\u_inv.f_next[163] ),
    .X(net3006));
 sg13g2_dlygate4sd3_1 hold1944 (.A(_00623_),
    .X(net3007));
 sg13g2_dlygate4sd3_1 hold1945 (.A(\u_inv.d_reg[162] ),
    .X(net3008));
 sg13g2_dlygate4sd3_1 hold1946 (.A(\u_inv.d_next[63] ),
    .X(net3009));
 sg13g2_dlygate4sd3_1 hold1947 (.A(_01313_),
    .X(net3010));
 sg13g2_dlygate4sd3_1 hold1948 (.A(\u_inv.d_next[43] ),
    .X(net3011));
 sg13g2_dlygate4sd3_1 hold1949 (.A(_01293_),
    .X(net3012));
 sg13g2_dlygate4sd3_1 hold1950 (.A(\u_inv.f_reg[143] ),
    .X(net3013));
 sg13g2_dlygate4sd3_1 hold1951 (.A(_01650_),
    .X(net3014));
 sg13g2_dlygate4sd3_1 hold1952 (.A(\shift_reg[37] ),
    .X(net3015));
 sg13g2_dlygate4sd3_1 hold1953 (.A(_00212_),
    .X(net3016));
 sg13g2_dlygate4sd3_1 hold1954 (.A(\u_inv.d_next[247] ),
    .X(net3017));
 sg13g2_dlygate4sd3_1 hold1955 (.A(_01497_),
    .X(net3018));
 sg13g2_dlygate4sd3_1 hold1956 (.A(\u_inv.input_reg[163] ),
    .X(net3019));
 sg13g2_dlygate4sd3_1 hold1957 (.A(\shift_reg[251] ),
    .X(net3020));
 sg13g2_dlygate4sd3_1 hold1958 (.A(_00426_),
    .X(net3021));
 sg13g2_dlygate4sd3_1 hold1959 (.A(\u_inv.f_next[12] ),
    .X(net3022));
 sg13g2_dlygate4sd3_1 hold1960 (.A(\u_inv.f_next[103] ),
    .X(net3023));
 sg13g2_dlygate4sd3_1 hold1961 (.A(\shift_reg[211] ),
    .X(net3024));
 sg13g2_dlygate4sd3_1 hold1962 (.A(\u_inv.d_reg[239] ),
    .X(net3025));
 sg13g2_dlygate4sd3_1 hold1963 (.A(\shift_reg[208] ),
    .X(net3026));
 sg13g2_dlygate4sd3_1 hold1964 (.A(\u_inv.d_next[199] ),
    .X(net3027));
 sg13g2_dlygate4sd3_1 hold1965 (.A(_01449_),
    .X(net3028));
 sg13g2_dlygate4sd3_1 hold1966 (.A(\u_inv.f_reg[236] ),
    .X(net3029));
 sg13g2_dlygate4sd3_1 hold1967 (.A(_01743_),
    .X(net3030));
 sg13g2_dlygate4sd3_1 hold1968 (.A(\shift_reg[73] ),
    .X(net3031));
 sg13g2_dlygate4sd3_1 hold1969 (.A(\u_inv.f_reg[176] ),
    .X(net3032));
 sg13g2_dlygate4sd3_1 hold1970 (.A(_01683_),
    .X(net3033));
 sg13g2_dlygate4sd3_1 hold1971 (.A(\u_inv.f_reg[221] ),
    .X(net3034));
 sg13g2_dlygate4sd3_1 hold1972 (.A(_01728_),
    .X(net3035));
 sg13g2_dlygate4sd3_1 hold1973 (.A(\u_inv.f_next[100] ),
    .X(net3036));
 sg13g2_dlygate4sd3_1 hold1974 (.A(\u_inv.f_next[120] ),
    .X(net3037));
 sg13g2_dlygate4sd3_1 hold1975 (.A(\u_inv.d_reg[206] ),
    .X(net3038));
 sg13g2_dlygate4sd3_1 hold1976 (.A(\u_inv.d_reg[24] ),
    .X(net3039));
 sg13g2_dlygate4sd3_1 hold1977 (.A(\shift_reg[55] ),
    .X(net3040));
 sg13g2_dlygate4sd3_1 hold1978 (.A(_00230_),
    .X(net3041));
 sg13g2_dlygate4sd3_1 hold1979 (.A(\u_inv.f_reg[29] ),
    .X(net3042));
 sg13g2_dlygate4sd3_1 hold1980 (.A(_01536_),
    .X(net3043));
 sg13g2_dlygate4sd3_1 hold1981 (.A(\u_inv.d_reg[246] ),
    .X(net3044));
 sg13g2_dlygate4sd3_1 hold1982 (.A(\u_inv.d_next[47] ),
    .X(net3045));
 sg13g2_dlygate4sd3_1 hold1983 (.A(_01297_),
    .X(net3046));
 sg13g2_dlygate4sd3_1 hold1984 (.A(\u_inv.f_next[14] ),
    .X(net3047));
 sg13g2_dlygate4sd3_1 hold1985 (.A(\shift_reg[95] ),
    .X(net3048));
 sg13g2_dlygate4sd3_1 hold1986 (.A(_00270_),
    .X(net3049));
 sg13g2_dlygate4sd3_1 hold1987 (.A(\u_inv.f_reg[115] ),
    .X(net3050));
 sg13g2_dlygate4sd3_1 hold1988 (.A(_01622_),
    .X(net3051));
 sg13g2_dlygate4sd3_1 hold1989 (.A(\u_inv.d_next[113] ),
    .X(net3052));
 sg13g2_dlygate4sd3_1 hold1990 (.A(_01363_),
    .X(net3053));
 sg13g2_dlygate4sd3_1 hold1991 (.A(\u_inv.f_next[109] ),
    .X(net3054));
 sg13g2_dlygate4sd3_1 hold1992 (.A(\u_inv.f_reg[247] ),
    .X(net3055));
 sg13g2_dlygate4sd3_1 hold1993 (.A(_01754_),
    .X(net3056));
 sg13g2_dlygate4sd3_1 hold1994 (.A(\inv_result[69] ),
    .X(net3057));
 sg13g2_dlygate4sd3_1 hold1995 (.A(\u_inv.d_next[168] ),
    .X(net3058));
 sg13g2_dlygate4sd3_1 hold1996 (.A(_01418_),
    .X(net3059));
 sg13g2_dlygate4sd3_1 hold1997 (.A(\shift_reg[53] ),
    .X(net3060));
 sg13g2_dlygate4sd3_1 hold1998 (.A(\shift_reg[96] ),
    .X(net3061));
 sg13g2_dlygate4sd3_1 hold1999 (.A(\shift_reg[242] ),
    .X(net3062));
 sg13g2_dlygate4sd3_1 hold2000 (.A(_00417_),
    .X(net3063));
 sg13g2_dlygate4sd3_1 hold2001 (.A(\u_inv.d_reg[251] ),
    .X(net3064));
 sg13g2_dlygate4sd3_1 hold2002 (.A(\u_inv.d_next[172] ),
    .X(net3065));
 sg13g2_dlygate4sd3_1 hold2003 (.A(_01422_),
    .X(net3066));
 sg13g2_dlygate4sd3_1 hold2004 (.A(\inv_result[131] ),
    .X(net3067));
 sg13g2_dlygate4sd3_1 hold2005 (.A(\u_inv.f_reg[89] ),
    .X(net3068));
 sg13g2_dlygate4sd3_1 hold2006 (.A(_01596_),
    .X(net3069));
 sg13g2_dlygate4sd3_1 hold2007 (.A(\u_inv.d_next[223] ),
    .X(net3070));
 sg13g2_dlygate4sd3_1 hold2008 (.A(_01473_),
    .X(net3071));
 sg13g2_dlygate4sd3_1 hold2009 (.A(\u_inv.f_reg[253] ),
    .X(net3072));
 sg13g2_dlygate4sd3_1 hold2010 (.A(_01760_),
    .X(net3073));
 sg13g2_dlygate4sd3_1 hold2011 (.A(\u_inv.d_next[61] ),
    .X(net3074));
 sg13g2_dlygate4sd3_1 hold2012 (.A(_01311_),
    .X(net3075));
 sg13g2_dlygate4sd3_1 hold2013 (.A(\shift_reg[227] ),
    .X(net3076));
 sg13g2_dlygate4sd3_1 hold2014 (.A(\u_inv.f_next[71] ),
    .X(net3077));
 sg13g2_dlygate4sd3_1 hold2015 (.A(\u_inv.d_next[16] ),
    .X(net3078));
 sg13g2_dlygate4sd3_1 hold2016 (.A(_01266_),
    .X(net3079));
 sg13g2_dlygate4sd3_1 hold2017 (.A(\u_inv.d_next[21] ),
    .X(net3080));
 sg13g2_dlygate4sd3_1 hold2018 (.A(_01271_),
    .X(net3081));
 sg13g2_dlygate4sd3_1 hold2019 (.A(\shift_reg[56] ),
    .X(net3082));
 sg13g2_dlygate4sd3_1 hold2020 (.A(\u_inv.f_next[36] ),
    .X(net3083));
 sg13g2_dlygate4sd3_1 hold2021 (.A(\u_inv.f_reg[133] ),
    .X(net3084));
 sg13g2_dlygate4sd3_1 hold2022 (.A(_01640_),
    .X(net3085));
 sg13g2_dlygate4sd3_1 hold2023 (.A(\shift_reg[93] ),
    .X(net3086));
 sg13g2_dlygate4sd3_1 hold2024 (.A(_00268_),
    .X(net3087));
 sg13g2_dlygate4sd3_1 hold2025 (.A(\shift_reg[86] ),
    .X(net3088));
 sg13g2_dlygate4sd3_1 hold2026 (.A(_00261_),
    .X(net3089));
 sg13g2_dlygate4sd3_1 hold2027 (.A(\u_inv.f_reg[192] ),
    .X(net3090));
 sg13g2_dlygate4sd3_1 hold2028 (.A(_01699_),
    .X(net3091));
 sg13g2_dlygate4sd3_1 hold2029 (.A(\shift_reg[126] ),
    .X(net3092));
 sg13g2_dlygate4sd3_1 hold2030 (.A(\u_inv.f_reg[84] ),
    .X(net3093));
 sg13g2_dlygate4sd3_1 hold2031 (.A(_01591_),
    .X(net3094));
 sg13g2_dlygate4sd3_1 hold2032 (.A(\u_inv.delta_reg[7] ),
    .X(net3095));
 sg13g2_dlygate4sd3_1 hold2033 (.A(\u_inv.d_next[33] ),
    .X(net3096));
 sg13g2_dlygate4sd3_1 hold2034 (.A(_01283_),
    .X(net3097));
 sg13g2_dlygate4sd3_1 hold2035 (.A(\shift_reg[153] ),
    .X(net3098));
 sg13g2_dlygate4sd3_1 hold2036 (.A(_00328_),
    .X(net3099));
 sg13g2_dlygate4sd3_1 hold2037 (.A(\shift_reg[49] ),
    .X(net3100));
 sg13g2_dlygate4sd3_1 hold2038 (.A(_00224_),
    .X(net3101));
 sg13g2_dlygate4sd3_1 hold2039 (.A(\shift_reg[204] ),
    .X(net3102));
 sg13g2_dlygate4sd3_1 hold2040 (.A(\u_inv.f_reg[135] ),
    .X(net3103));
 sg13g2_dlygate4sd3_1 hold2041 (.A(_01642_),
    .X(net3104));
 sg13g2_dlygate4sd3_1 hold2042 (.A(\u_inv.d_next[160] ),
    .X(net3105));
 sg13g2_dlygate4sd3_1 hold2043 (.A(_01410_),
    .X(net3106));
 sg13g2_dlygate4sd3_1 hold2044 (.A(\shift_reg[164] ),
    .X(net3107));
 sg13g2_dlygate4sd3_1 hold2045 (.A(_00339_),
    .X(net3108));
 sg13g2_dlygate4sd3_1 hold2046 (.A(\u_inv.f_reg[57] ),
    .X(net3109));
 sg13g2_dlygate4sd3_1 hold2047 (.A(_01564_),
    .X(net3110));
 sg13g2_dlygate4sd3_1 hold2048 (.A(\u_inv.d_next[176] ),
    .X(net3111));
 sg13g2_dlygate4sd3_1 hold2049 (.A(_01426_),
    .X(net3112));
 sg13g2_dlygate4sd3_1 hold2050 (.A(\u_inv.f_reg[147] ),
    .X(net3113));
 sg13g2_dlygate4sd3_1 hold2051 (.A(_01654_),
    .X(net3114));
 sg13g2_dlygate4sd3_1 hold2052 (.A(\shift_reg[215] ),
    .X(net3115));
 sg13g2_dlygate4sd3_1 hold2053 (.A(\shift_reg[47] ),
    .X(net3116));
 sg13g2_dlygate4sd3_1 hold2054 (.A(\shift_reg[66] ),
    .X(net3117));
 sg13g2_dlygate4sd3_1 hold2055 (.A(\shift_reg[92] ),
    .X(net3118));
 sg13g2_dlygate4sd3_1 hold2056 (.A(\u_inv.d_next[101] ),
    .X(net3119));
 sg13g2_dlygate4sd3_1 hold2057 (.A(_01351_),
    .X(net3120));
 sg13g2_dlygate4sd3_1 hold2058 (.A(\perf_triple[3] ),
    .X(net3121));
 sg13g2_dlygate4sd3_1 hold2059 (.A(\shift_reg[98] ),
    .X(net3122));
 sg13g2_dlygate4sd3_1 hold2060 (.A(_00273_),
    .X(net3123));
 sg13g2_dlygate4sd3_1 hold2061 (.A(\u_inv.d_next[44] ),
    .X(net3124));
 sg13g2_dlygate4sd3_1 hold2062 (.A(_01294_),
    .X(net3125));
 sg13g2_dlygate4sd3_1 hold2063 (.A(\shift_reg[85] ),
    .X(net3126));
 sg13g2_dlygate4sd3_1 hold2064 (.A(_00260_),
    .X(net3127));
 sg13g2_dlygate4sd3_1 hold2065 (.A(\u_inv.d_next[121] ),
    .X(net3128));
 sg13g2_dlygate4sd3_1 hold2066 (.A(_01371_),
    .X(net3129));
 sg13g2_dlygate4sd3_1 hold2067 (.A(\u_inv.f_next[231] ),
    .X(net3130));
 sg13g2_dlygate4sd3_1 hold2068 (.A(\u_inv.f_reg[210] ),
    .X(net3131));
 sg13g2_dlygate4sd3_1 hold2069 (.A(_01717_),
    .X(net3132));
 sg13g2_dlygate4sd3_1 hold2070 (.A(\u_inv.d_next[26] ),
    .X(net3133));
 sg13g2_dlygate4sd3_1 hold2071 (.A(_01276_),
    .X(net3134));
 sg13g2_dlygate4sd3_1 hold2072 (.A(\u_inv.f_next[48] ),
    .X(net3135));
 sg13g2_dlygate4sd3_1 hold2073 (.A(\u_inv.f_reg[185] ),
    .X(net3136));
 sg13g2_dlygate4sd3_1 hold2074 (.A(_01692_),
    .X(net3137));
 sg13g2_dlygate4sd3_1 hold2075 (.A(\u_inv.d_reg[244] ),
    .X(net3138));
 sg13g2_dlygate4sd3_1 hold2076 (.A(\shift_reg[67] ),
    .X(net3139));
 sg13g2_dlygate4sd3_1 hold2077 (.A(_00242_),
    .X(net3140));
 sg13g2_dlygate4sd3_1 hold2078 (.A(\u_inv.f_next[10] ),
    .X(net3141));
 sg13g2_dlygate4sd3_1 hold2079 (.A(\u_inv.d_next[23] ),
    .X(net3142));
 sg13g2_dlygate4sd3_1 hold2080 (.A(_01273_),
    .X(net3143));
 sg13g2_dlygate4sd3_1 hold2081 (.A(\u_inv.d_reg[202] ),
    .X(net3144));
 sg13g2_dlygate4sd3_1 hold2082 (.A(\u_inv.d_next[9] ),
    .X(net3145));
 sg13g2_dlygate4sd3_1 hold2083 (.A(_01259_),
    .X(net3146));
 sg13g2_dlygate4sd3_1 hold2084 (.A(\shift_reg[115] ),
    .X(net3147));
 sg13g2_dlygate4sd3_1 hold2085 (.A(_00290_),
    .X(net3148));
 sg13g2_dlygate4sd3_1 hold2086 (.A(\u_inv.d_next[231] ),
    .X(net3149));
 sg13g2_dlygate4sd3_1 hold2087 (.A(_01481_),
    .X(net3150));
 sg13g2_dlygate4sd3_1 hold2088 (.A(\u_inv.f_next[143] ),
    .X(net3151));
 sg13g2_dlygate4sd3_1 hold2089 (.A(\shift_reg[103] ),
    .X(net3152));
 sg13g2_dlygate4sd3_1 hold2090 (.A(\u_inv.f_reg[124] ),
    .X(net3153));
 sg13g2_dlygate4sd3_1 hold2091 (.A(_01631_),
    .X(net3154));
 sg13g2_dlygate4sd3_1 hold2092 (.A(\u_inv.f_reg[196] ),
    .X(net3155));
 sg13g2_dlygate4sd3_1 hold2093 (.A(_01703_),
    .X(net3156));
 sg13g2_dlygate4sd3_1 hold2094 (.A(\u_inv.d_next[122] ),
    .X(net3157));
 sg13g2_dlygate4sd3_1 hold2095 (.A(_01372_),
    .X(net3158));
 sg13g2_dlygate4sd3_1 hold2096 (.A(\u_inv.f_reg[139] ),
    .X(net3159));
 sg13g2_dlygate4sd3_1 hold2097 (.A(_01646_),
    .X(net3160));
 sg13g2_dlygate4sd3_1 hold2098 (.A(\u_inv.d_next[233] ),
    .X(net3161));
 sg13g2_dlygate4sd3_1 hold2099 (.A(_01483_),
    .X(net3162));
 sg13g2_dlygate4sd3_1 hold2100 (.A(\u_inv.d_next[39] ),
    .X(net3163));
 sg13g2_dlygate4sd3_1 hold2101 (.A(_01289_),
    .X(net3164));
 sg13g2_dlygate4sd3_1 hold2102 (.A(\u_inv.input_reg[125] ),
    .X(net3165));
 sg13g2_dlygate4sd3_1 hold2103 (.A(_00032_),
    .X(net3166));
 sg13g2_dlygate4sd3_1 hold2104 (.A(\u_inv.f_next[127] ),
    .X(net3167));
 sg13g2_dlygate4sd3_1 hold2105 (.A(\shift_reg[87] ),
    .X(net3168));
 sg13g2_dlygate4sd3_1 hold2106 (.A(_00262_),
    .X(net3169));
 sg13g2_dlygate4sd3_1 hold2107 (.A(\u_inv.input_reg[124] ),
    .X(net3170));
 sg13g2_dlygate4sd3_1 hold2108 (.A(_00031_),
    .X(net3171));
 sg13g2_dlygate4sd3_1 hold2109 (.A(\inv_result[215] ),
    .X(net3172));
 sg13g2_dlygate4sd3_1 hold2110 (.A(\inv_result[27] ),
    .X(net3173));
 sg13g2_dlygate4sd3_1 hold2111 (.A(\inv_result[73] ),
    .X(net3174));
 sg13g2_dlygate4sd3_1 hold2112 (.A(\u_inv.d_next[93] ),
    .X(net3175));
 sg13g2_dlygate4sd3_1 hold2113 (.A(_01343_),
    .X(net3176));
 sg13g2_dlygate4sd3_1 hold2114 (.A(\shift_reg[183] ),
    .X(net3177));
 sg13g2_dlygate4sd3_1 hold2115 (.A(_00358_),
    .X(net3178));
 sg13g2_dlygate4sd3_1 hold2116 (.A(\u_inv.d_reg[49] ),
    .X(net3179));
 sg13g2_dlygate4sd3_1 hold2117 (.A(\inv_result[49] ),
    .X(net3180));
 sg13g2_dlygate4sd3_1 hold2118 (.A(\u_inv.d_next[167] ),
    .X(net3181));
 sg13g2_dlygate4sd3_1 hold2119 (.A(_01417_),
    .X(net3182));
 sg13g2_dlygate4sd3_1 hold2120 (.A(\shift_reg[116] ),
    .X(net3183));
 sg13g2_dlygate4sd3_1 hold2121 (.A(_00291_),
    .X(net3184));
 sg13g2_dlygate4sd3_1 hold2122 (.A(\u_inv.f_next[81] ),
    .X(net3185));
 sg13g2_dlygate4sd3_1 hold2123 (.A(\inv_result[245] ),
    .X(net3186));
 sg13g2_dlygate4sd3_1 hold2124 (.A(\u_inv.f_next[130] ),
    .X(net3187));
 sg13g2_dlygate4sd3_1 hold2125 (.A(\u_inv.f_next[74] ),
    .X(net3188));
 sg13g2_dlygate4sd3_1 hold2126 (.A(\inv_result[64] ),
    .X(net3189));
 sg13g2_dlygate4sd3_1 hold2127 (.A(\u_inv.f_reg[179] ),
    .X(net3190));
 sg13g2_dlygate4sd3_1 hold2128 (.A(\shift_reg[34] ),
    .X(net3191));
 sg13g2_dlygate4sd3_1 hold2129 (.A(_00209_),
    .X(net3192));
 sg13g2_dlygate4sd3_1 hold2130 (.A(\shift_reg[102] ),
    .X(net3193));
 sg13g2_dlygate4sd3_1 hold2131 (.A(_00277_),
    .X(net3194));
 sg13g2_dlygate4sd3_1 hold2132 (.A(\u_inv.f_next[232] ),
    .X(net3195));
 sg13g2_dlygate4sd3_1 hold2133 (.A(\u_inv.f_reg[231] ),
    .X(net3196));
 sg13g2_dlygate4sd3_1 hold2134 (.A(\u_inv.f_reg[19] ),
    .X(net3197));
 sg13g2_dlygate4sd3_1 hold2135 (.A(_01526_),
    .X(net3198));
 sg13g2_dlygate4sd3_1 hold2136 (.A(\u_inv.d_next[67] ),
    .X(net3199));
 sg13g2_dlygate4sd3_1 hold2137 (.A(_01317_),
    .X(net3200));
 sg13g2_dlygate4sd3_1 hold2138 (.A(\u_inv.d_reg[238] ),
    .X(net3201));
 sg13g2_dlygate4sd3_1 hold2139 (.A(\shift_reg[210] ),
    .X(net3202));
 sg13g2_dlygate4sd3_1 hold2140 (.A(\u_inv.f_reg[225] ),
    .X(net3203));
 sg13g2_dlygate4sd3_1 hold2141 (.A(_01732_),
    .X(net3204));
 sg13g2_dlygate4sd3_1 hold2142 (.A(\u_inv.f_next[34] ),
    .X(net3205));
 sg13g2_dlygate4sd3_1 hold2143 (.A(\shift_reg[30] ),
    .X(net3206));
 sg13g2_dlygate4sd3_1 hold2144 (.A(_00205_),
    .X(net3207));
 sg13g2_dlygate4sd3_1 hold2145 (.A(\u_inv.f_reg[111] ),
    .X(net3208));
 sg13g2_dlygate4sd3_1 hold2146 (.A(_01618_),
    .X(net3209));
 sg13g2_dlygate4sd3_1 hold2147 (.A(\u_inv.d_next[22] ),
    .X(net3210));
 sg13g2_dlygate4sd3_1 hold2148 (.A(_01272_),
    .X(net3211));
 sg13g2_dlygate4sd3_1 hold2149 (.A(\inv_result[145] ),
    .X(net3212));
 sg13g2_dlygate4sd3_1 hold2150 (.A(\u_inv.d_reg[198] ),
    .X(net3213));
 sg13g2_dlygate4sd3_1 hold2151 (.A(\u_inv.f_reg[255] ),
    .X(net3214));
 sg13g2_dlygate4sd3_1 hold2152 (.A(_01762_),
    .X(net3215));
 sg13g2_dlygate4sd3_1 hold2153 (.A(\shift_reg[111] ),
    .X(net3216));
 sg13g2_dlygate4sd3_1 hold2154 (.A(\u_inv.f_next[173] ),
    .X(net3217));
 sg13g2_dlygate4sd3_1 hold2155 (.A(\shift_reg[71] ),
    .X(net3218));
 sg13g2_dlygate4sd3_1 hold2156 (.A(_00246_),
    .X(net3219));
 sg13g2_dlygate4sd3_1 hold2157 (.A(\u_inv.d_next[157] ),
    .X(net3220));
 sg13g2_dlygate4sd3_1 hold2158 (.A(_01407_),
    .X(net3221));
 sg13g2_dlygate4sd3_1 hold2159 (.A(\inv_result[203] ),
    .X(net3222));
 sg13g2_dlygate4sd3_1 hold2160 (.A(\shift_reg[182] ),
    .X(net3223));
 sg13g2_dlygate4sd3_1 hold2161 (.A(_00357_),
    .X(net3224));
 sg13g2_dlygate4sd3_1 hold2162 (.A(\u_inv.d_next[134] ),
    .X(net3225));
 sg13g2_dlygate4sd3_1 hold2163 (.A(\shift_reg[64] ),
    .X(net3226));
 sg13g2_dlygate4sd3_1 hold2164 (.A(\shift_reg[63] ),
    .X(net3227));
 sg13g2_dlygate4sd3_1 hold2165 (.A(\shift_reg[226] ),
    .X(net3228));
 sg13g2_dlygate4sd3_1 hold2166 (.A(_00401_),
    .X(net3229));
 sg13g2_dlygate4sd3_1 hold2167 (.A(\u_inv.f_next[151] ),
    .X(net3230));
 sg13g2_dlygate4sd3_1 hold2168 (.A(\u_inv.d_next[228] ),
    .X(net3231));
 sg13g2_dlygate4sd3_1 hold2169 (.A(\u_inv.f_reg[126] ),
    .X(net3232));
 sg13g2_dlygate4sd3_1 hold2170 (.A(_01633_),
    .X(net3233));
 sg13g2_dlygate4sd3_1 hold2171 (.A(\shift_reg[221] ),
    .X(net3234));
 sg13g2_dlygate4sd3_1 hold2172 (.A(_00396_),
    .X(net3235));
 sg13g2_dlygate4sd3_1 hold2173 (.A(\u_inv.d_next[53] ),
    .X(net3236));
 sg13g2_dlygate4sd3_1 hold2174 (.A(_01303_),
    .X(net3237));
 sg13g2_dlygate4sd3_1 hold2175 (.A(\u_inv.f_next[91] ),
    .X(net3238));
 sg13g2_dlygate4sd3_1 hold2176 (.A(\u_inv.d_next[69] ),
    .X(net3239));
 sg13g2_dlygate4sd3_1 hold2177 (.A(_01319_),
    .X(net3240));
 sg13g2_dlygate4sd3_1 hold2178 (.A(\u_inv.f_reg[171] ),
    .X(net3241));
 sg13g2_dlygate4sd3_1 hold2179 (.A(\shift_reg[167] ),
    .X(net3242));
 sg13g2_dlygate4sd3_1 hold2180 (.A(_00342_),
    .X(net3243));
 sg13g2_dlygate4sd3_1 hold2181 (.A(\u_inv.f_reg[208] ),
    .X(net3244));
 sg13g2_dlygate4sd3_1 hold2182 (.A(_01715_),
    .X(net3245));
 sg13g2_dlygate4sd3_1 hold2183 (.A(\shift_reg[29] ),
    .X(net3246));
 sg13g2_dlygate4sd3_1 hold2184 (.A(_00204_),
    .X(net3247));
 sg13g2_dlygate4sd3_1 hold2185 (.A(\shift_reg[162] ),
    .X(net3248));
 sg13g2_dlygate4sd3_1 hold2186 (.A(_00337_),
    .X(net3249));
 sg13g2_dlygate4sd3_1 hold2187 (.A(\shift_reg[59] ),
    .X(net3250));
 sg13g2_dlygate4sd3_1 hold2188 (.A(\shift_reg[94] ),
    .X(net3251));
 sg13g2_dlygate4sd3_1 hold2189 (.A(\u_inv.d_next[114] ),
    .X(net3252));
 sg13g2_dlygate4sd3_1 hold2190 (.A(\u_inv.d_next[141] ),
    .X(net3253));
 sg13g2_dlygate4sd3_1 hold2191 (.A(_01391_),
    .X(net3254));
 sg13g2_dlygate4sd3_1 hold2192 (.A(\u_inv.d_reg[102] ),
    .X(net3255));
 sg13g2_dlygate4sd3_1 hold2193 (.A(\shift_reg[152] ),
    .X(net3256));
 sg13g2_dlygate4sd3_1 hold2194 (.A(_00327_),
    .X(net3257));
 sg13g2_dlygate4sd3_1 hold2195 (.A(\u_inv.d_reg[59] ),
    .X(net3258));
 sg13g2_dlygate4sd3_1 hold2196 (.A(\u_inv.f_next[250] ),
    .X(net3259));
 sg13g2_dlygate4sd3_1 hold2197 (.A(\u_inv.d_next[73] ),
    .X(net3260));
 sg13g2_dlygate4sd3_1 hold2198 (.A(\shift_reg[31] ),
    .X(net3261));
 sg13g2_dlygate4sd3_1 hold2199 (.A(\shift_reg[237] ),
    .X(net3262));
 sg13g2_dlygate4sd3_1 hold2200 (.A(_00412_),
    .X(net3263));
 sg13g2_dlygate4sd3_1 hold2201 (.A(\u_inv.d_reg[114] ),
    .X(net3264));
 sg13g2_dlygate4sd3_1 hold2202 (.A(\shift_reg[21] ),
    .X(net3265));
 sg13g2_dlygate4sd3_1 hold2203 (.A(\u_inv.f_next[113] ),
    .X(net3266));
 sg13g2_dlygate4sd3_1 hold2204 (.A(\u_inv.f_next[43] ),
    .X(net3267));
 sg13g2_dlygate4sd3_1 hold2205 (.A(\shift_reg[68] ),
    .X(net3268));
 sg13g2_dlygate4sd3_1 hold2206 (.A(_00243_),
    .X(net3269));
 sg13g2_dlygate4sd3_1 hold2207 (.A(\u_inv.f_reg[151] ),
    .X(net3270));
 sg13g2_dlygate4sd3_1 hold2208 (.A(\u_inv.d_next[209] ),
    .X(net3271));
 sg13g2_dlygate4sd3_1 hold2209 (.A(_01459_),
    .X(net3272));
 sg13g2_dlygate4sd3_1 hold2210 (.A(\u_inv.d_next[232] ),
    .X(net3273));
 sg13g2_dlygate4sd3_1 hold2211 (.A(\u_inv.d_next[78] ),
    .X(net3274));
 sg13g2_dlygate4sd3_1 hold2212 (.A(_01328_),
    .X(net3275));
 sg13g2_dlygate4sd3_1 hold2213 (.A(\u_inv.f_reg[234] ),
    .X(net3276));
 sg13g2_dlygate4sd3_1 hold2214 (.A(_01741_),
    .X(net3277));
 sg13g2_dlygate4sd3_1 hold2215 (.A(\shift_reg[35] ),
    .X(net3278));
 sg13g2_dlygate4sd3_1 hold2216 (.A(_00210_),
    .X(net3279));
 sg13g2_dlygate4sd3_1 hold2217 (.A(\u_inv.d_reg[90] ),
    .X(net3280));
 sg13g2_dlygate4sd3_1 hold2218 (.A(\shift_reg[177] ),
    .X(net3281));
 sg13g2_dlygate4sd3_1 hold2219 (.A(_00352_),
    .X(net3282));
 sg13g2_dlygate4sd3_1 hold2220 (.A(\inv_result[129] ),
    .X(net3283));
 sg13g2_dlygate4sd3_1 hold2221 (.A(\perf_triple[5] ),
    .X(net3284));
 sg13g2_dlygate4sd3_1 hold2222 (.A(\u_inv.d_next[151] ),
    .X(net3285));
 sg13g2_dlygate4sd3_1 hold2223 (.A(\shift_reg[40] ),
    .X(net3286));
 sg13g2_dlygate4sd3_1 hold2224 (.A(\u_inv.d_reg[62] ),
    .X(net3287));
 sg13g2_dlygate4sd3_1 hold2225 (.A(\shift_reg[161] ),
    .X(net3288));
 sg13g2_dlygate4sd3_1 hold2226 (.A(\u_inv.f_reg[25] ),
    .X(net3289));
 sg13g2_dlygate4sd3_1 hold2227 (.A(_01532_),
    .X(net3290));
 sg13g2_dlygate4sd3_1 hold2228 (.A(\u_inv.d_reg[226] ),
    .X(net3291));
 sg13g2_dlygate4sd3_1 hold2229 (.A(\u_inv.f_next[102] ),
    .X(net3292));
 sg13g2_dlygate4sd3_1 hold2230 (.A(\u_inv.d_next[20] ),
    .X(net3293));
 sg13g2_dlygate4sd3_1 hold2231 (.A(_01270_),
    .X(net3294));
 sg13g2_dlygate4sd3_1 hold2232 (.A(\shift_reg[52] ),
    .X(net3295));
 sg13g2_dlygate4sd3_1 hold2233 (.A(\u_inv.d_next[133] ),
    .X(net3296));
 sg13g2_dlygate4sd3_1 hold2234 (.A(\shift_reg[89] ),
    .X(net3297));
 sg13g2_dlygate4sd3_1 hold2235 (.A(\u_inv.f_next[110] ),
    .X(net3298));
 sg13g2_dlygate4sd3_1 hold2236 (.A(\u_inv.d_next[129] ),
    .X(net3299));
 sg13g2_dlygate4sd3_1 hold2237 (.A(_01379_),
    .X(net3300));
 sg13g2_dlygate4sd3_1 hold2238 (.A(\shift_reg[158] ),
    .X(net3301));
 sg13g2_dlygate4sd3_1 hold2239 (.A(_00333_),
    .X(net3302));
 sg13g2_dlygate4sd3_1 hold2240 (.A(\u_inv.f_next[23] ),
    .X(net3303));
 sg13g2_dlygate4sd3_1 hold2241 (.A(\inv_result[253] ),
    .X(net3304));
 sg13g2_dlygate4sd3_1 hold2242 (.A(\inv_result[214] ),
    .X(net3305));
 sg13g2_dlygate4sd3_1 hold2244 (.A(\u_inv.d_next[137] ),
    .X(net3307));
 sg13g2_dlygate4sd3_1 hold2245 (.A(_01387_),
    .X(net3308));
 sg13g2_dlygate4sd3_1 hold2246 (.A(\u_inv.d_reg[232] ),
    .X(net3309));
 sg13g2_dlygate4sd3_1 hold2247 (.A(\shift_reg[180] ),
    .X(net3310));
 sg13g2_dlygate4sd3_1 hold2248 (.A(_00355_),
    .X(net3311));
 sg13g2_dlygate4sd3_1 hold2249 (.A(\u_inv.f_next[35] ),
    .X(net3312));
 sg13g2_dlygate4sd3_1 hold2250 (.A(\u_inv.f_next[202] ),
    .X(net3313));
 sg13g2_dlygate4sd3_1 hold2251 (.A(\u_inv.d_next[159] ),
    .X(net3314));
 sg13g2_dlygate4sd3_1 hold2252 (.A(_01409_),
    .X(net3315));
 sg13g2_dlygate4sd3_1 hold2253 (.A(\inv_result[85] ),
    .X(net3316));
 sg13g2_dlygate4sd3_1 hold2254 (.A(\u_inv.f_next[75] ),
    .X(net3317));
 sg13g2_dlygate4sd3_1 hold2255 (.A(\shift_reg[231] ),
    .X(net3318));
 sg13g2_dlygate4sd3_1 hold2256 (.A(_00406_),
    .X(net3319));
 sg13g2_dlygate4sd3_1 hold2257 (.A(\inv_result[121] ),
    .X(net3320));
 sg13g2_dlygate4sd3_1 hold2258 (.A(\u_inv.d_next[108] ),
    .X(net3321));
 sg13g2_dlygate4sd3_1 hold2259 (.A(_01358_),
    .X(net3322));
 sg13g2_dlygate4sd3_1 hold2260 (.A(\u_inv.d_next[40] ),
    .X(net3323));
 sg13g2_dlygate4sd3_1 hold2261 (.A(_01290_),
    .X(net3324));
 sg13g2_dlygate4sd3_1 hold2262 (.A(\shift_reg[119] ),
    .X(net3325));
 sg13g2_dlygate4sd3_1 hold2263 (.A(\u_inv.f_next[213] ),
    .X(net3326));
 sg13g2_dlygate4sd3_1 hold2264 (.A(\u_inv.d_next[112] ),
    .X(net3327));
 sg13g2_dlygate4sd3_1 hold2265 (.A(\inv_result[10] ),
    .X(net3328));
 sg13g2_dlygate4sd3_1 hold2266 (.A(\shift_reg[159] ),
    .X(net3329));
 sg13g2_dlygate4sd3_1 hold2267 (.A(_00334_),
    .X(net3330));
 sg13g2_dlygate4sd3_1 hold2268 (.A(\u_inv.f_next[2] ),
    .X(net3331));
 sg13g2_dlygate4sd3_1 hold2269 (.A(\shift_reg[154] ),
    .X(net3332));
 sg13g2_dlygate4sd3_1 hold2270 (.A(_00329_),
    .X(net3333));
 sg13g2_dlygate4sd3_1 hold2271 (.A(\u_inv.d_next[84] ),
    .X(net3334));
 sg13g2_dlygate4sd3_1 hold2272 (.A(_01334_),
    .X(net3335));
 sg13g2_dlygate4sd3_1 hold2273 (.A(\shift_reg[26] ),
    .X(net3336));
 sg13g2_dlygate4sd3_1 hold2274 (.A(_00201_),
    .X(net3337));
 sg13g2_dlygate4sd3_1 hold2275 (.A(\u_inv.d_reg[146] ),
    .X(net3338));
 sg13g2_dlygate4sd3_1 hold2276 (.A(\shift_reg[165] ),
    .X(net3339));
 sg13g2_dlygate4sd3_1 hold2277 (.A(\u_inv.d_next[68] ),
    .X(net3340));
 sg13g2_dlygate4sd3_1 hold2278 (.A(_01318_),
    .X(net3341));
 sg13g2_dlygate4sd3_1 hold2279 (.A(\u_inv.d_next[103] ),
    .X(net3342));
 sg13g2_dlygate4sd3_1 hold2280 (.A(_01353_),
    .X(net3343));
 sg13g2_dlygate4sd3_1 hold2281 (.A(\u_inv.f_reg[69] ),
    .X(net3344));
 sg13g2_dlygate4sd3_1 hold2282 (.A(_01576_),
    .X(net3345));
 sg13g2_dlygate4sd3_1 hold2283 (.A(\shift_reg[90] ),
    .X(net3346));
 sg13g2_dlygate4sd3_1 hold2284 (.A(\u_inv.d_next[252] ),
    .X(net3347));
 sg13g2_dlygate4sd3_1 hold2285 (.A(\u_inv.f_next[174] ),
    .X(net3348));
 sg13g2_dlygate4sd3_1 hold2286 (.A(\u_inv.f_next[135] ),
    .X(net3349));
 sg13g2_dlygate4sd3_1 hold2287 (.A(\u_inv.f_next[188] ),
    .X(net3350));
 sg13g2_dlygate4sd3_1 hold2288 (.A(\shift_reg[171] ),
    .X(net3351));
 sg13g2_dlygate4sd3_1 hold2289 (.A(_00346_),
    .X(net3352));
 sg13g2_dlygate4sd3_1 hold2290 (.A(\u_inv.d_next[45] ),
    .X(net3353));
 sg13g2_dlygate4sd3_1 hold2291 (.A(_01295_),
    .X(net3354));
 sg13g2_dlygate4sd3_1 hold2292 (.A(\u_inv.f_next[191] ),
    .X(net3355));
 sg13g2_dlygate4sd3_1 hold2293 (.A(\perf_triple[8] ),
    .X(net3356));
 sg13g2_dlygate4sd3_1 hold2294 (.A(\shift_reg[141] ),
    .X(net3357));
 sg13g2_dlygate4sd3_1 hold2295 (.A(\u_inv.f_next[153] ),
    .X(net3358));
 sg13g2_dlygate4sd3_1 hold2296 (.A(\u_inv.f_next[85] ),
    .X(net3359));
 sg13g2_dlygate4sd3_1 hold2297 (.A(\u_inv.d_next[125] ),
    .X(net3360));
 sg13g2_dlygate4sd3_1 hold2298 (.A(_01375_),
    .X(net3361));
 sg13g2_dlygate4sd3_1 hold2299 (.A(\inv_result[171] ),
    .X(net3362));
 sg13g2_dlygate4sd3_1 hold2300 (.A(\u_inv.d_next[131] ),
    .X(net3363));
 sg13g2_dlygate4sd3_1 hold2301 (.A(_01381_),
    .X(net3364));
 sg13g2_dlygate4sd3_1 hold2302 (.A(\inv_result[221] ),
    .X(net3365));
 sg13g2_dlygate4sd3_1 hold2303 (.A(\u_inv.d_next[148] ),
    .X(net3366));
 sg13g2_dlygate4sd3_1 hold2304 (.A(_01398_),
    .X(net3367));
 sg13g2_dlygate4sd3_1 hold2305 (.A(\u_inv.f_next[251] ),
    .X(net3368));
 sg13g2_dlygate4sd3_1 hold2306 (.A(\u_inv.f_next[226] ),
    .X(net3369));
 sg13g2_dlygate4sd3_1 hold2307 (.A(\inv_result[91] ),
    .X(net3370));
 sg13g2_dlygate4sd3_1 hold2308 (.A(\inv_result[251] ),
    .X(net3371));
 sg13g2_dlygate4sd3_1 hold2309 (.A(\u_inv.f_next[67] ),
    .X(net3372));
 sg13g2_dlygate4sd3_1 hold2310 (.A(\shift_reg[108] ),
    .X(net3373));
 sg13g2_dlygate4sd3_1 hold2311 (.A(\u_inv.d_next[185] ),
    .X(net3374));
 sg13g2_dlygate4sd3_1 hold2312 (.A(_01435_),
    .X(net3375));
 sg13g2_dlygate4sd3_1 hold2313 (.A(\u_inv.d_next[227] ),
    .X(net3376));
 sg13g2_dlygate4sd3_1 hold2314 (.A(_01477_),
    .X(net3377));
 sg13g2_dlygate4sd3_1 hold2315 (.A(\u_inv.f_next[53] ),
    .X(net3378));
 sg13g2_dlygate4sd3_1 hold2316 (.A(\shift_reg[138] ),
    .X(net3379));
 sg13g2_dlygate4sd3_1 hold2317 (.A(\shift_reg[60] ),
    .X(net3380));
 sg13g2_dlygate4sd3_1 hold2318 (.A(\shift_reg[156] ),
    .X(net3381));
 sg13g2_dlygate4sd3_1 hold2319 (.A(_00331_),
    .X(net3382));
 sg13g2_dlygate4sd3_1 hold2320 (.A(\u_inv.d_next[19] ),
    .X(net3383));
 sg13g2_dlygate4sd3_1 hold2321 (.A(_01269_),
    .X(net3384));
 sg13g2_dlygate4sd3_1 hold2322 (.A(\shift_reg[20] ),
    .X(net3385));
 sg13g2_dlygate4sd3_1 hold2323 (.A(\u_inv.f_next[144] ),
    .X(net3386));
 sg13g2_dlygate4sd3_1 hold2324 (.A(\shift_reg[61] ),
    .X(net3387));
 sg13g2_dlygate4sd3_1 hold2325 (.A(\u_inv.d_reg[256] ),
    .X(net3388));
 sg13g2_dlygate4sd3_1 hold2326 (.A(\u_inv.d_next[195] ),
    .X(net3389));
 sg13g2_dlygate4sd3_1 hold2327 (.A(_01445_),
    .X(net3390));
 sg13g2_dlygate4sd3_1 hold2328 (.A(\u_inv.f_next[157] ),
    .X(net3391));
 sg13g2_dlygate4sd3_1 hold2329 (.A(\u_inv.f_next[82] ),
    .X(net3392));
 sg13g2_dlygate4sd3_1 hold2330 (.A(\u_inv.d_next[75] ),
    .X(net3393));
 sg13g2_dlygate4sd3_1 hold2331 (.A(_01325_),
    .X(net3394));
 sg13g2_dlygate4sd3_1 hold2332 (.A(\shift_reg[223] ),
    .X(net3395));
 sg13g2_dlygate4sd3_1 hold2333 (.A(\u_inv.d_next[143] ),
    .X(net3396));
 sg13g2_dlygate4sd3_1 hold2334 (.A(_01393_),
    .X(net3397));
 sg13g2_dlygate4sd3_1 hold2335 (.A(\shift_reg[143] ),
    .X(net3398));
 sg13g2_dlygate4sd3_1 hold2336 (.A(\shift_reg[27] ),
    .X(net3399));
 sg13g2_dlygate4sd3_1 hold2337 (.A(_00202_),
    .X(net3400));
 sg13g2_dlygate4sd3_1 hold2338 (.A(\u_inv.f_next[245] ),
    .X(net3401));
 sg13g2_dlygate4sd3_1 hold2339 (.A(\shift_reg[4] ),
    .X(net3402));
 sg13g2_dlygate4sd3_1 hold2340 (.A(_00179_),
    .X(net3403));
 sg13g2_dlygate4sd3_1 hold2341 (.A(\u_inv.d_reg[236] ),
    .X(net3404));
 sg13g2_dlygate4sd3_1 hold2342 (.A(\u_inv.d_next[255] ),
    .X(net3405));
 sg13g2_dlygate4sd3_1 hold2343 (.A(_01505_),
    .X(net3406));
 sg13g2_dlygate4sd3_1 hold2344 (.A(\u_inv.f_next[253] ),
    .X(net3407));
 sg13g2_dlygate4sd3_1 hold2345 (.A(\u_inv.d_next[52] ),
    .X(net3408));
 sg13g2_dlygate4sd3_1 hold2346 (.A(\u_inv.f_next[249] ),
    .X(net3409));
 sg13g2_dlygate4sd3_1 hold2347 (.A(\shift_reg[213] ),
    .X(net3410));
 sg13g2_dlygate4sd3_1 hold2348 (.A(\u_inv.f_next[31] ),
    .X(net3411));
 sg13g2_dlygate4sd3_1 hold2349 (.A(\perf_triple[0] ),
    .X(net3412));
 sg13g2_dlygate4sd3_1 hold2350 (.A(\u_inv.d_next[132] ),
    .X(net3413));
 sg13g2_dlygate4sd3_1 hold2351 (.A(_01382_),
    .X(net3414));
 sg13g2_dlygate4sd3_1 hold2352 (.A(\shift_reg[172] ),
    .X(net3415));
 sg13g2_dlygate4sd3_1 hold2353 (.A(\u_inv.d_next[41] ),
    .X(net3416));
 sg13g2_dlygate4sd3_1 hold2354 (.A(_01291_),
    .X(net3417));
 sg13g2_dlygate4sd3_1 hold2355 (.A(\u_inv.f_next[252] ),
    .X(net3418));
 sg13g2_dlygate4sd3_1 hold2356 (.A(\u_inv.f_next[203] ),
    .X(net3419));
 sg13g2_dlygate4sd3_1 hold2357 (.A(\u_inv.delta_reg[1] ),
    .X(net3420));
 sg13g2_dlygate4sd3_1 hold2358 (.A(\inv_result[179] ),
    .X(net3421));
 sg13g2_dlygate4sd3_1 hold2359 (.A(\u_inv.d_reg[150] ),
    .X(net3422));
 sg13g2_dlygate4sd3_1 hold2360 (.A(\shift_reg[97] ),
    .X(net3423));
 sg13g2_dlygate4sd3_1 hold2361 (.A(\shift_reg[38] ),
    .X(net3424));
 sg13g2_dlygate4sd3_1 hold2362 (.A(\u_inv.d_next[208] ),
    .X(net3425));
 sg13g2_dlygate4sd3_1 hold2363 (.A(_01458_),
    .X(net3426));
 sg13g2_dlygate4sd3_1 hold2364 (.A(\shift_reg[78] ),
    .X(net3427));
 sg13g2_dlygate4sd3_1 hold2365 (.A(_00253_),
    .X(net3428));
 sg13g2_dlygate4sd3_1 hold2366 (.A(\shift_reg[140] ),
    .X(net3429));
 sg13g2_dlygate4sd3_1 hold2367 (.A(\shift_reg[70] ),
    .X(net3430));
 sg13g2_dlygate4sd3_1 hold2368 (.A(_00245_),
    .X(net3431));
 sg13g2_dlygate4sd3_1 hold2369 (.A(\shift_reg[224] ),
    .X(net3432));
 sg13g2_dlygate4sd3_1 hold2370 (.A(_00399_),
    .X(net3433));
 sg13g2_dlygate4sd3_1 hold2371 (.A(\u_inv.f_next[78] ),
    .X(net3434));
 sg13g2_dlygate4sd3_1 hold2372 (.A(\u_inv.f_next[142] ),
    .X(net3435));
 sg13g2_dlygate4sd3_1 hold2373 (.A(\u_inv.f_next[38] ),
    .X(net3436));
 sg13g2_dlygate4sd3_1 hold2374 (.A(\shift_reg[163] ),
    .X(net3437));
 sg13g2_dlygate4sd3_1 hold2375 (.A(\u_inv.d_next[197] ),
    .X(net3438));
 sg13g2_dlygate4sd3_1 hold2376 (.A(\shift_reg[72] ),
    .X(net3439));
 sg13g2_dlygate4sd3_1 hold2377 (.A(\shift_reg[79] ),
    .X(net3440));
 sg13g2_dlygate4sd3_1 hold2378 (.A(\shift_reg[105] ),
    .X(net3441));
 sg13g2_dlygate4sd3_1 hold2379 (.A(\shift_reg[76] ),
    .X(net3442));
 sg13g2_dlygate4sd3_1 hold2380 (.A(\shift_reg[77] ),
    .X(net3443));
 sg13g2_dlygate4sd3_1 hold2381 (.A(_00252_),
    .X(net3444));
 sg13g2_dlygate4sd3_1 hold2382 (.A(\u_inv.d_next[229] ),
    .X(net3445));
 sg13g2_dlygate4sd3_1 hold2383 (.A(_01479_),
    .X(net3446));
 sg13g2_dlygate4sd3_1 hold2384 (.A(\shift_reg[160] ),
    .X(net3447));
 sg13g2_dlygate4sd3_1 hold2385 (.A(\u_inv.f_next[160] ),
    .X(net3448));
 sg13g2_dlygate4sd3_1 hold2386 (.A(\shift_reg[142] ),
    .X(net3449));
 sg13g2_dlygate4sd3_1 hold2387 (.A(\shift_reg[6] ),
    .X(net3450));
 sg13g2_dlygate4sd3_1 hold2388 (.A(_00181_),
    .X(net3451));
 sg13g2_dlygate4sd3_1 hold2389 (.A(\shift_reg[62] ),
    .X(net3452));
 sg13g2_dlygate4sd3_1 hold2390 (.A(_00237_),
    .X(net3453));
 sg13g2_dlygate4sd3_1 hold2391 (.A(\inv_result[117] ),
    .X(net3454));
 sg13g2_dlygate4sd3_1 hold2392 (.A(\u_inv.d_next[203] ),
    .X(net3455));
 sg13g2_dlygate4sd3_1 hold2393 (.A(_01453_),
    .X(net3456));
 sg13g2_dlygate4sd3_1 hold2394 (.A(\u_inv.f_next[164] ),
    .X(net3457));
 sg13g2_dlygate4sd3_1 hold2395 (.A(\shift_reg[22] ),
    .X(net3458));
 sg13g2_dlygate4sd3_1 hold2396 (.A(\u_inv.f_next[133] ),
    .X(net3459));
 sg13g2_dlygate4sd3_1 hold2397 (.A(\u_inv.f_next[166] ),
    .X(net3460));
 sg13g2_dlygate4sd3_1 hold2398 (.A(\shift_reg[75] ),
    .X(net3461));
 sg13g2_dlygate4sd3_1 hold2399 (.A(\u_inv.d_next[83] ),
    .X(net3462));
 sg13g2_dlygate4sd3_1 hold2400 (.A(_01333_),
    .X(net3463));
 sg13g2_dlygate4sd3_1 hold2401 (.A(\shift_reg[110] ),
    .X(net3464));
 sg13g2_dlygate4sd3_1 hold2402 (.A(\u_inv.d_reg[189] ),
    .X(net3465));
 sg13g2_dlygate4sd3_1 hold2403 (.A(_01439_),
    .X(net3466));
 sg13g2_dlygate4sd3_1 hold2404 (.A(\shift_reg[54] ),
    .X(net3467));
 sg13g2_dlygate4sd3_1 hold2405 (.A(_00229_),
    .X(net3468));
 sg13g2_dlygate4sd3_1 hold2406 (.A(\u_inv.f_next[246] ),
    .X(net3469));
 sg13g2_dlygate4sd3_1 hold2407 (.A(\shift_reg[216] ),
    .X(net3470));
 sg13g2_dlygate4sd3_1 hold2408 (.A(\u_inv.d_next[30] ),
    .X(net3471));
 sg13g2_dlygate4sd3_1 hold2409 (.A(_01280_),
    .X(net3472));
 sg13g2_dlygate4sd3_1 hold2410 (.A(\u_inv.f_next[117] ),
    .X(net3473));
 sg13g2_dlygate4sd3_1 hold2411 (.A(\shift_reg[19] ),
    .X(net3474));
 sg13g2_dlygate4sd3_1 hold2412 (.A(\u_inv.d_next[135] ),
    .X(net3475));
 sg13g2_dlygate4sd3_1 hold2413 (.A(_01385_),
    .X(net3476));
 sg13g2_dlygate4sd3_1 hold2414 (.A(\u_inv.d_next[74] ),
    .X(net3477));
 sg13g2_dlygate4sd3_1 hold2415 (.A(_01324_),
    .X(net3478));
 sg13g2_dlygate4sd3_1 hold2416 (.A(\shift_reg[148] ),
    .X(net3479));
 sg13g2_dlygate4sd3_1 hold2417 (.A(\u_inv.d_reg[71] ),
    .X(net3480));
 sg13g2_dlygate4sd3_1 hold2418 (.A(\u_inv.f_next[86] ),
    .X(net3481));
 sg13g2_dlygate4sd3_1 hold2419 (.A(\u_inv.f_next[19] ),
    .X(net3482));
 sg13g2_dlygate4sd3_1 hold2420 (.A(\u_inv.d_reg[230] ),
    .X(net3483));
 sg13g2_dlygate4sd3_1 hold2421 (.A(\shift_reg[222] ),
    .X(net3484));
 sg13g2_dlygate4sd3_1 hold2422 (.A(\u_inv.f_next[50] ),
    .X(net3485));
 sg13g2_dlygate4sd3_1 hold2423 (.A(\inv_result[153] ),
    .X(net3486));
 sg13g2_dlygate4sd3_1 hold2424 (.A(\shift_reg[139] ),
    .X(net3487));
 sg13g2_dlygate4sd3_1 hold2425 (.A(\u_inv.f_next[63] ),
    .X(net3488));
 sg13g2_dlygate4sd3_1 hold2426 (.A(\shift_reg[170] ),
    .X(net3489));
 sg13g2_dlygate4sd3_1 hold2427 (.A(\inv_result[61] ),
    .X(net3490));
 sg13g2_dlygate4sd3_1 hold2428 (.A(\u_inv.f_next[229] ),
    .X(net3491));
 sg13g2_dlygate4sd3_1 hold2429 (.A(\shift_reg[43] ),
    .X(net3492));
 sg13g2_dlygate4sd3_1 hold2430 (.A(\u_inv.d_next[253] ),
    .X(net3493));
 sg13g2_dlygate4sd3_1 hold2431 (.A(\u_inv.d_next[87] ),
    .X(net3494));
 sg13g2_dlygate4sd3_1 hold2432 (.A(_01337_),
    .X(net3495));
 sg13g2_dlygate4sd3_1 hold2433 (.A(\u_inv.f_next[99] ),
    .X(net3496));
 sg13g2_dlygate4sd3_1 hold2434 (.A(\inv_result[225] ),
    .X(net3497));
 sg13g2_dlygate4sd3_1 hold2435 (.A(\shift_reg[181] ),
    .X(net3498));
 sg13g2_dlygate4sd3_1 hold2436 (.A(_00356_),
    .X(net3499));
 sg13g2_dlygate4sd3_1 hold2437 (.A(\shift_reg[106] ),
    .X(net3500));
 sg13g2_dlygate4sd3_1 hold2438 (.A(\u_inv.f_next[241] ),
    .X(net3501));
 sg13g2_dlygate4sd3_1 hold2439 (.A(\u_inv.f_next[187] ),
    .X(net3502));
 sg13g2_dlygate4sd3_1 hold2440 (.A(\shift_reg[228] ),
    .X(net3503));
 sg13g2_dlygate4sd3_1 hold2441 (.A(\u_inv.d_next[249] ),
    .X(net3504));
 sg13g2_dlygate4sd3_1 hold2442 (.A(_01499_),
    .X(net3505));
 sg13g2_dlygate4sd3_1 hold2443 (.A(\u_inv.d_next[217] ),
    .X(net3506));
 sg13g2_dlygate4sd3_1 hold2444 (.A(_01467_),
    .X(net3507));
 sg13g2_dlygate4sd3_1 hold2445 (.A(\shift_reg[145] ),
    .X(net3508));
 sg13g2_dlygate4sd3_1 hold2446 (.A(\u_inv.f_next[114] ),
    .X(net3509));
 sg13g2_dlygate4sd3_1 hold2447 (.A(\u_inv.d_next[86] ),
    .X(net3510));
 sg13g2_dlygate4sd3_1 hold2448 (.A(_01336_),
    .X(net3511));
 sg13g2_dlygate4sd3_1 hold2449 (.A(\shift_reg[191] ),
    .X(net3512));
 sg13g2_dlygate4sd3_1 hold2450 (.A(\u_inv.f_next[186] ),
    .X(net3513));
 sg13g2_dlygate4sd3_1 hold2451 (.A(\u_trng.prev_sample ),
    .X(net3514));
 sg13g2_dlygate4sd3_1 hold2452 (.A(\u_inv.d_reg[73] ),
    .X(net3515));
 sg13g2_dlygate4sd3_1 hold2453 (.A(\shift_reg[150] ),
    .X(net3516));
 sg13g2_dlygate4sd3_1 hold2454 (.A(\shift_reg[109] ),
    .X(net3517));
 sg13g2_dlygate4sd3_1 hold2455 (.A(\shift_reg[188] ),
    .X(net3518));
 sg13g2_dlygate4sd3_1 hold2456 (.A(\shift_reg[218] ),
    .X(net3519));
 sg13g2_dlygate4sd3_1 hold2457 (.A(\u_inv.f_next[18] ),
    .X(net3520));
 sg13g2_dlygate4sd3_1 hold2458 (.A(\shift_reg[176] ),
    .X(net3521));
 sg13g2_dlygate4sd3_1 hold2459 (.A(_00351_),
    .X(net3522));
 sg13g2_dlygate4sd3_1 hold2460 (.A(\u_inv.d_next[72] ),
    .X(net3523));
 sg13g2_dlygate4sd3_1 hold2461 (.A(_01322_),
    .X(net3524));
 sg13g2_dlygate4sd3_1 hold2462 (.A(\u_inv.d_reg[253] ),
    .X(net3525));
 sg13g2_dlygate4sd3_1 hold2463 (.A(\shift_reg[24] ),
    .X(net3526));
 sg13g2_dlygate4sd3_1 hold2464 (.A(_00199_),
    .X(net3527));
 sg13g2_dlygate4sd3_1 hold2465 (.A(\shift_reg[42] ),
    .X(net3528));
 sg13g2_dlygate4sd3_1 hold2466 (.A(\shift_reg[169] ),
    .X(net3529));
 sg13g2_dlygate4sd3_1 hold2467 (.A(\shift_reg[17] ),
    .X(net3530));
 sg13g2_dlygate4sd3_1 hold2468 (.A(\u_inv.f_next[198] ),
    .X(net3531));
 sg13g2_dlygate4sd3_1 hold2469 (.A(\u_inv.f_next[29] ),
    .X(net3532));
 sg13g2_dlygate4sd3_1 hold2470 (.A(\u_inv.d_reg[166] ),
    .X(net3533));
 sg13g2_dlygate4sd3_1 hold2471 (.A(\shift_reg[46] ),
    .X(net3534));
 sg13g2_dlygate4sd3_1 hold2472 (.A(\u_inv.f_next[236] ),
    .X(net3535));
 sg13g2_dlygate4sd3_1 hold2473 (.A(\u_inv.d_reg[52] ),
    .X(net3536));
 sg13g2_dlygate4sd3_1 hold2474 (.A(\u_inv.f_next[159] ),
    .X(net3537));
 sg13g2_dlygate4sd3_1 hold2475 (.A(\shift_reg[28] ),
    .X(net3538));
 sg13g2_dlygate4sd3_1 hold2476 (.A(\u_inv.d_next[191] ),
    .X(net3539));
 sg13g2_dlygate4sd3_1 hold2477 (.A(_01441_),
    .X(net3540));
 sg13g2_dlygate4sd3_1 hold2478 (.A(\shift_reg[166] ),
    .X(net3541));
 sg13g2_dlygate4sd3_1 hold2479 (.A(\u_inv.d_reg[228] ),
    .X(net3542));
 sg13g2_dlygate4sd3_1 hold2480 (.A(\u_inv.d_next[248] ),
    .X(net3543));
 sg13g2_dlygate4sd3_1 hold2481 (.A(_01498_),
    .X(net3544));
 sg13g2_dlygate4sd3_1 hold2482 (.A(\shift_reg[173] ),
    .X(net3545));
 sg13g2_dlygate4sd3_1 hold2483 (.A(\u_inv.f_next[193] ),
    .X(net3546));
 sg13g2_dlygate4sd3_1 hold2484 (.A(\u_inv.d_next[193] ),
    .X(net3547));
 sg13g2_dlygate4sd3_1 hold2485 (.A(\shift_reg[189] ),
    .X(net3548));
 sg13g2_dlygate4sd3_1 hold2486 (.A(\u_inv.d_next[196] ),
    .X(net3549));
 sg13g2_dlygate4sd3_1 hold2487 (.A(_01446_),
    .X(net3550));
 sg13g2_dlygate4sd3_1 hold2488 (.A(\u_inv.d_reg[17] ),
    .X(net3551));
 sg13g2_dlygate4sd3_1 hold2489 (.A(\shift_reg[147] ),
    .X(net3552));
 sg13g2_dlygate4sd3_1 hold2490 (.A(\u_inv.f_next[107] ),
    .X(net3553));
 sg13g2_dlygate4sd3_1 hold2491 (.A(\u_inv.f_next[152] ),
    .X(net3554));
 sg13g2_dlygate4sd3_1 hold2493 (.A(_18481_),
    .X(net3556));
 sg13g2_dlygate4sd3_1 hold2494 (.A(\shift_reg[178] ),
    .X(net3557));
 sg13g2_dlygate4sd3_1 hold2495 (.A(\shift_reg[25] ),
    .X(net3558));
 sg13g2_dlygate4sd3_1 hold2496 (.A(\shift_reg[168] ),
    .X(net3559));
 sg13g2_dlygate4sd3_1 hold2497 (.A(\u_inv.f_next[66] ),
    .X(net3560));
 sg13g2_dlygate4sd3_1 hold2498 (.A(\u_inv.d_next[169] ),
    .X(net3561));
 sg13g2_dlygate4sd3_1 hold2499 (.A(_01419_),
    .X(net3562));
 sg13g2_dlygate4sd3_1 hold2500 (.A(\u_inv.f_next[150] ),
    .X(net3563));
 sg13g2_dlygate4sd3_1 hold2501 (.A(\u_inv.f_next[1] ),
    .X(net3564));
 sg13g2_dlygate4sd3_1 hold2502 (.A(\shift_reg[41] ),
    .X(net3565));
 sg13g2_dlygate4sd3_1 hold2503 (.A(\u_inv.d_next[89] ),
    .X(net3566));
 sg13g2_dlygate4sd3_1 hold2504 (.A(_01339_),
    .X(net3567));
 sg13g2_dlygate4sd3_1 hold2505 (.A(\u_inv.d_next[139] ),
    .X(net3568));
 sg13g2_dlygate4sd3_1 hold2506 (.A(_01389_),
    .X(net3569));
 sg13g2_dlygate4sd3_1 hold2507 (.A(\shift_reg[144] ),
    .X(net3570));
 sg13g2_dlygate4sd3_1 hold2508 (.A(\u_inv.d_reg[134] ),
    .X(net3571));
 sg13g2_dlygate4sd3_1 hold2509 (.A(\shift_reg[151] ),
    .X(net3572));
 sg13g2_dlygate4sd3_1 hold2510 (.A(\shift_reg[149] ),
    .X(net3573));
 sg13g2_dlygate4sd3_1 hold2511 (.A(\u_inv.d_reg[252] ),
    .X(net3574));
 sg13g2_dlygate4sd3_1 hold2512 (.A(\u_inv.d_next[241] ),
    .X(net3575));
 sg13g2_dlygate4sd3_1 hold2513 (.A(_01491_),
    .X(net3576));
 sg13g2_dlygate4sd3_1 hold2514 (.A(\shift_reg[74] ),
    .X(net3577));
 sg13g2_dlygate4sd3_1 hold2515 (.A(\perf_double[0] ),
    .X(net3578));
 sg13g2_dlygate4sd3_1 hold2516 (.A(\u_inv.d_next[51] ),
    .X(net3579));
 sg13g2_dlygate4sd3_1 hold2517 (.A(_01301_),
    .X(net3580));
 sg13g2_dlygate4sd3_1 hold2518 (.A(\u_inv.d_next[215] ),
    .X(net3581));
 sg13g2_dlygate4sd3_1 hold2519 (.A(_01465_),
    .X(net3582));
 sg13g2_dlygate4sd3_1 hold2520 (.A(\u_inv.d_next[56] ),
    .X(net3583));
 sg13g2_dlygate4sd3_1 hold2521 (.A(_01306_),
    .X(net3584));
 sg13g2_dlygate4sd3_1 hold2522 (.A(\u_inv.d_next[127] ),
    .X(net3585));
 sg13g2_dlygate4sd3_1 hold2523 (.A(\u_inv.f_next[212] ),
    .X(net3586));
 sg13g2_dlygate4sd3_1 hold2524 (.A(\u_inv.f_next[168] ),
    .X(net3587));
 sg13g2_dlygate4sd3_1 hold2525 (.A(\u_inv.f_next[47] ),
    .X(net3588));
 sg13g2_dlygate4sd3_1 hold2526 (.A(\u_inv.f_next[57] ),
    .X(net3589));
 sg13g2_dlygate4sd3_1 hold2527 (.A(\u_inv.d_reg[197] ),
    .X(net3590));
 sg13g2_dlygate4sd3_1 hold2528 (.A(\inv_result[0] ),
    .X(net3591));
 sg13g2_dlygate4sd3_1 hold2529 (.A(_00994_),
    .X(net3592));
 sg13g2_dlygate4sd3_1 hold2530 (.A(\u_inv.d_next[235] ),
    .X(net3593));
 sg13g2_dlygate4sd3_1 hold2531 (.A(_01485_),
    .X(net3594));
 sg13g2_dlygate4sd3_1 hold2532 (.A(\u_inv.f_next[22] ),
    .X(net3595));
 sg13g2_dlygate4sd3_1 hold2533 (.A(\u_inv.f_next[201] ),
    .X(net3596));
 sg13g2_dlygate4sd3_1 hold2534 (.A(\shift_reg[174] ),
    .X(net3597));
 sg13g2_dlygate4sd3_1 hold2535 (.A(\u_inv.d_reg[18] ),
    .X(net3598));
 sg13g2_dlygate4sd3_1 hold2536 (.A(\u_inv.f_next[123] ),
    .X(net3599));
 sg13g2_dlygate4sd3_1 hold2537 (.A(\shift_reg[104] ),
    .X(net3600));
 sg13g2_dlygate4sd3_1 hold2538 (.A(\u_inv.d_next[242] ),
    .X(net3601));
 sg13g2_dlygate4sd3_1 hold2539 (.A(\u_inv.delta_double[0] ),
    .X(net3602));
 sg13g2_dlygate4sd3_1 hold2540 (.A(\u_inv.f_next[122] ),
    .X(net3603));
 sg13g2_dlygate4sd3_1 hold2541 (.A(\u_inv.d_reg[111] ),
    .X(net3604));
 sg13g2_dlygate4sd3_1 hold2542 (.A(_01361_),
    .X(net3605));
 sg13g2_dlygate4sd3_1 hold2543 (.A(\u_inv.d_next[240] ),
    .X(net3606));
 sg13g2_dlygate4sd3_1 hold2544 (.A(_01490_),
    .X(net3607));
 sg13g2_dlygate4sd3_1 hold2545 (.A(\u_inv.d_reg[151] ),
    .X(net3608));
 sg13g2_dlygate4sd3_1 hold2546 (.A(\u_inv.f_next[222] ),
    .X(net3609));
 sg13g2_dlygate4sd3_1 hold2547 (.A(\u_inv.d_reg[193] ),
    .X(net3610));
 sg13g2_dlygate4sd3_1 hold2548 (.A(\u_inv.d_reg[242] ),
    .X(net3611));
 sg13g2_dlygate4sd3_1 hold2549 (.A(\u_inv.f_next[195] ),
    .X(net3612));
 sg13g2_dlygate4sd3_1 hold2550 (.A(\u_inv.f_next[223] ),
    .X(net3613));
 sg13g2_dlygate4sd3_1 hold2551 (.A(\u_inv.f_next[73] ),
    .X(net3614));
 sg13g2_dlygate4sd3_1 hold2552 (.A(\shift_reg[146] ),
    .X(net3615));
 sg13g2_dlygate4sd3_1 hold2553 (.A(\u_inv.d_reg[127] ),
    .X(net3616));
 sg13g2_dlygate4sd3_1 hold2554 (.A(\u_inv.f_next[137] ),
    .X(net3617));
 sg13g2_dlygate4sd3_1 hold2555 (.A(\u_inv.d_reg[142] ),
    .X(net3618));
 sg13g2_dlygate4sd3_1 hold2556 (.A(\u_inv.f_next[162] ),
    .X(net3619));
 sg13g2_dlygate4sd3_1 hold2557 (.A(\u_inv.d_next[213] ),
    .X(net3620));
 sg13g2_dlygate4sd3_1 hold2558 (.A(_01463_),
    .X(net3621));
 sg13g2_dlygate4sd3_1 hold2559 (.A(\shift_reg[229] ),
    .X(net3622));
 sg13g2_dlygate4sd3_1 hold2560 (.A(\shift_reg[175] ),
    .X(net3623));
 sg13g2_dlygate4sd3_1 hold2561 (.A(\u_inv.f_next[155] ),
    .X(net3624));
 sg13g2_dlygate4sd3_1 hold2562 (.A(\u_inv.d_next[147] ),
    .X(net3625));
 sg13g2_dlygate4sd3_1 hold2563 (.A(_01397_),
    .X(net3626));
 sg13g2_dlygate4sd3_1 hold2564 (.A(\u_inv.f_next[80] ),
    .X(net3627));
 sg13g2_dlygate4sd3_1 hold2565 (.A(\u_inv.f_next[20] ),
    .X(net3628));
 sg13g2_dlygate4sd3_1 hold2566 (.A(\shift_reg[18] ),
    .X(net3629));
 sg13g2_dlygate4sd3_1 hold2567 (.A(\u_inv.f_next[138] ),
    .X(net3630));
 sg13g2_dlygate4sd3_1 hold2568 (.A(\u_inv.f_next[169] ),
    .X(net3631));
 sg13g2_dlygate4sd3_1 hold2569 (.A(\u_inv.f_next[27] ),
    .X(net3632));
 sg13g2_dlygate4sd3_1 hold2570 (.A(\u_inv.f_next[254] ),
    .X(net3633));
 sg13g2_dlygate4sd3_1 hold2571 (.A(\u_inv.f_next[215] ),
    .X(net3634));
 sg13g2_dlygate4sd3_1 hold2572 (.A(\inv_result[235] ),
    .X(net3635));
 sg13g2_dlygate4sd3_1 hold2573 (.A(\u_inv.counter[4] ),
    .X(net3636));
 sg13g2_dlygate4sd3_1 hold2574 (.A(\u_inv.f_next[132] ),
    .X(net3637));
 sg13g2_dlygate4sd3_1 hold2575 (.A(\u_inv.f_next[189] ),
    .X(net3638));
 sg13g2_dlygate4sd3_1 hold2576 (.A(\u_inv.counter[5] ),
    .X(net3639));
 sg13g2_dlygate4sd3_1 hold2577 (.A(\u_inv.d_reg[95] ),
    .X(net3640));
 sg13g2_dlygate4sd3_1 hold2578 (.A(_01345_),
    .X(net3641));
 sg13g2_dlygate4sd3_1 hold2579 (.A(\u_inv.f_next[24] ),
    .X(net3642));
 sg13g2_dlygate4sd3_1 hold2580 (.A(\shift_reg[225] ),
    .X(net3643));
 sg13g2_dlygate4sd3_1 hold2581 (.A(\u_inv.f_next[8] ),
    .X(net3644));
 sg13g2_dlygate4sd3_1 hold2582 (.A(\u_inv.f_next[141] ),
    .X(net3645));
 sg13g2_dlygate4sd3_1 hold2583 (.A(\u_inv.f_next[125] ),
    .X(net3646));
 sg13g2_dlygate4sd3_1 hold2584 (.A(\u_inv.f_next[72] ),
    .X(net3647));
 sg13g2_dlygate4sd3_1 hold2585 (.A(\u_inv.f_next[146] ),
    .X(net3648));
 sg13g2_dlygate4sd3_1 hold2586 (.A(\u_inv.f_next[61] ),
    .X(net3649));
 sg13g2_dlygate4sd3_1 hold2587 (.A(\u_inv.f_next[79] ),
    .X(net3650));
 sg13g2_dlygate4sd3_1 hold2588 (.A(\u_inv.f_next[70] ),
    .X(net3651));
 sg13g2_dlygate4sd3_1 hold2589 (.A(\u_inv.d_next[97] ),
    .X(net3652));
 sg13g2_dlygate4sd3_1 hold2590 (.A(_01347_),
    .X(net3653));
 sg13g2_dlygate4sd3_1 hold2591 (.A(\u_inv.f_next[83] ),
    .X(net3654));
 sg13g2_dlygate4sd3_1 hold2592 (.A(\u_inv.f_next[211] ),
    .X(net3655));
 sg13g2_dlygate4sd3_1 hold2593 (.A(\u_inv.f_next[111] ),
    .X(net3656));
 sg13g2_dlygate4sd3_1 hold2594 (.A(\u_inv.f_next[64] ),
    .X(net3657));
 sg13g2_dlygate4sd3_1 hold2595 (.A(\u_inv.f_next[69] ),
    .X(net3658));
 sg13g2_dlygate4sd3_1 hold2596 (.A(\u_inv.d_next[81] ),
    .X(net3659));
 sg13g2_dlygate4sd3_1 hold2597 (.A(\shift_reg[16] ),
    .X(net3660));
 sg13g2_dlygate4sd3_1 hold2598 (.A(\shift_reg[107] ),
    .X(net3661));
 sg13g2_dlygate4sd3_1 hold2599 (.A(\u_inv.f_next[197] ),
    .X(net3662));
 sg13g2_dlygate4sd3_1 hold2600 (.A(\u_inv.f_next[46] ),
    .X(net3663));
 sg13g2_dlygate4sd3_1 hold2601 (.A(\u_inv.d_next[99] ),
    .X(net3664));
 sg13g2_dlygate4sd3_1 hold2602 (.A(_01349_),
    .X(net3665));
 sg13g2_dlygate4sd3_1 hold2603 (.A(\u_inv.f_next[62] ),
    .X(net3666));
 sg13g2_dlygate4sd3_1 hold2604 (.A(\u_inv.f_next[54] ),
    .X(net3667));
 sg13g2_dlygate4sd3_1 hold2605 (.A(inv_done),
    .X(net3668));
 sg13g2_dlygate4sd3_1 hold2606 (.A(_18627_),
    .X(net3669));
 sg13g2_dlygate4sd3_1 hold2607 (.A(\u_inv.f_next[196] ),
    .X(net3670));
 sg13g2_dlygate4sd3_1 hold2608 (.A(\shift_reg[5] ),
    .X(net3671));
 sg13g2_dlygate4sd3_1 hold2609 (.A(_00180_),
    .X(net3672));
 sg13g2_dlygate4sd3_1 hold2610 (.A(\u_inv.d_reg[70] ),
    .X(net3673));
 sg13g2_dlygate4sd3_1 hold2611 (.A(\u_inv.f_next[244] ),
    .X(net3674));
 sg13g2_dlygate4sd3_1 hold2612 (.A(\u_inv.d_reg[245] ),
    .X(net3675));
 sg13g2_dlygate4sd3_1 hold2613 (.A(\u_inv.f_next[220] ),
    .X(net3676));
 sg13g2_dlygate4sd3_1 hold2614 (.A(\u_inv.f_next[255] ),
    .X(net3677));
 sg13g2_dlygate4sd3_1 hold2615 (.A(\u_inv.f_next[92] ),
    .X(net3678));
 sg13g2_dlygate4sd3_1 hold2616 (.A(\u_inv.f_next[126] ),
    .X(net3679));
 sg13g2_dlygate4sd3_1 hold2617 (.A(\u_inv.d_reg[112] ),
    .X(net3680));
 sg13g2_dlygate4sd3_1 hold2618 (.A(\u_inv.d_next[57] ),
    .X(net3681));
 sg13g2_dlygate4sd3_1 hold2619 (.A(\u_inv.f_next[192] ),
    .X(net3682));
 sg13g2_dlygate4sd3_1 hold2620 (.A(\u_inv.f_next[247] ),
    .X(net3683));
 sg13g2_dlygate4sd3_1 hold2621 (.A(\u_inv.f_next[106] ),
    .X(net3684));
 sg13g2_dlygate4sd3_1 hold2622 (.A(\u_inv.f_next[134] ),
    .X(net3685));
 sg13g2_dlygate4sd3_1 hold2623 (.A(\u_inv.f_next[124] ),
    .X(net3686));
 sg13g2_dlygate4sd3_1 hold2624 (.A(\u_inv.f_next[108] ),
    .X(net3687));
 sg13g2_dlygate4sd3_1 hold2625 (.A(\u_inv.f_next[154] ),
    .X(net3688));
 sg13g2_dlygate4sd3_1 hold2626 (.A(\u_inv.f_next[149] ),
    .X(net3689));
 sg13g2_dlygate4sd3_1 hold2627 (.A(\u_inv.f_next[3] ),
    .X(net3690));
 sg13g2_dlygate4sd3_1 hold2628 (.A(\u_inv.f_next[248] ),
    .X(net3691));
 sg13g2_dlygate4sd3_1 hold2629 (.A(\u_inv.counter[1] ),
    .X(net3692));
 sg13g2_dlygate4sd3_1 hold2630 (.A(\perf_total[1] ),
    .X(net3693));
 sg13g2_dlygate4sd3_1 hold2631 (.A(\u_inv.f_next[161] ),
    .X(net3694));
 sg13g2_dlygate4sd3_1 hold2632 (.A(\u_inv.f_next[178] ),
    .X(net3695));
 sg13g2_dlygate4sd3_1 hold2633 (.A(\u_inv.f_next[58] ),
    .X(net3696));
 sg13g2_dlygate4sd3_1 hold2634 (.A(_02579_),
    .X(net3697));
 sg13g2_dlygate4sd3_1 hold2635 (.A(\u_inv.f_next[185] ),
    .X(net3698));
 sg13g2_dlygate4sd3_1 hold2636 (.A(\u_inv.f_next[200] ),
    .X(net3699));
 sg13g2_dlygate4sd3_1 hold2637 (.A(\u_inv.f_next[190] ),
    .X(net3700));
 sg13g2_dlygate4sd3_1 hold2638 (.A(\u_inv.f_next[89] ),
    .X(net3701));
 sg13g2_dlygate4sd3_1 hold2639 (.A(\u_inv.f_next[221] ),
    .X(net3702));
 sg13g2_dlygate4sd3_1 hold2640 (.A(\u_inv.f_next[208] ),
    .X(net3703));
 sg13g2_dlygate4sd3_1 hold2641 (.A(\u_inv.f_next[28] ),
    .X(net3704));
 sg13g2_dlygate4sd3_1 hold2642 (.A(\u_inv.f_next[230] ),
    .X(net3705));
 sg13g2_dlygate4sd3_1 hold2643 (.A(\u_inv.f_next[147] ),
    .X(net3706));
 sg13g2_dlygate4sd3_1 hold2644 (.A(\u_inv.f_next[194] ),
    .X(net3707));
 sg13g2_dlygate4sd3_1 hold2645 (.A(\u_inv.f_next[170] ),
    .X(net3708));
 sg13g2_dlygate4sd3_1 hold2646 (.A(\u_inv.f_next[13] ),
    .X(net3709));
 sg13g2_dlygate4sd3_1 hold2647 (.A(\u_inv.f_next[172] ),
    .X(net3710));
 sg13g2_dlygate4sd3_1 hold2648 (.A(\u_inv.f_next[206] ),
    .X(net3711));
 sg13g2_dlygate4sd3_1 hold2649 (.A(\u_inv.f_next[128] ),
    .X(net3712));
 sg13g2_dlygate4sd3_1 hold2650 (.A(\u_inv.f_next[30] ),
    .X(net3713));
 sg13g2_dlygate4sd3_1 hold2651 (.A(\u_inv.f_next[76] ),
    .X(net3714));
 sg13g2_dlygate4sd3_1 hold2652 (.A(\u_inv.f_next[59] ),
    .X(net3715));
 sg13g2_dlygate4sd3_1 hold2653 (.A(\u_inv.f_next[238] ),
    .X(net3716));
 sg13g2_dlygate4sd3_1 hold2654 (.A(\u_inv.f_next[68] ),
    .X(net3717));
 sg13g2_dlygate4sd3_1 hold2655 (.A(\u_inv.f_next[77] ),
    .X(net3718));
 sg13g2_dlygate4sd3_1 hold2656 (.A(\u_inv.f_next[25] ),
    .X(net3719));
 sg13g2_dlygate4sd3_1 hold2657 (.A(\u_inv.f_next[136] ),
    .X(net3720));
 sg13g2_dlygate4sd3_1 hold2658 (.A(\u_inv.f_next[210] ),
    .X(net3721));
 sg13g2_dlygate4sd3_1 hold2659 (.A(\u_inv.f_next[242] ),
    .X(net3722));
 sg13g2_dlygate4sd3_1 hold2660 (.A(\u_inv.d_next[95] ),
    .X(net3723));
 sg13g2_dlygate4sd3_1 hold2661 (.A(\u_inv.f_next[94] ),
    .X(net3724));
 sg13g2_dlygate4sd3_1 hold2662 (.A(\u_inv.f_next[214] ),
    .X(net3725));
 sg13g2_dlygate4sd3_1 hold2663 (.A(\u_inv.f_next[84] ),
    .X(net3726));
 sg13g2_dlygate4sd3_1 hold2664 (.A(\u_inv.f_next[158] ),
    .X(net3727));
 sg13g2_dlygate4sd3_1 hold2665 (.A(\u_inv.f_next[115] ),
    .X(net3728));
 sg13g2_dlygate4sd3_1 hold2666 (.A(\u_inv.f_next[176] ),
    .X(net3729));
 sg13g2_dlygate4sd3_1 hold2667 (.A(\u_inv.f_next[239] ),
    .X(net3730));
 sg13g2_dlygate4sd3_1 hold2668 (.A(\u_inv.f_next[182] ),
    .X(net3731));
 sg13g2_dlygate4sd3_1 hold2669 (.A(\u_inv.f_next[228] ),
    .X(net3732));
 sg13g2_dlygate4sd3_1 hold2670 (.A(\u_inv.f_next[237] ),
    .X(net3733));
 sg13g2_dlygate4sd3_1 hold2671 (.A(\u_inv.f_next[148] ),
    .X(net3734));
 sg13g2_dlygate4sd3_1 hold2672 (.A(\u_inv.f_next[240] ),
    .X(net3735));
 sg13g2_dlygate4sd3_1 hold2673 (.A(\u_inv.f_next[204] ),
    .X(net3736));
 sg13g2_dlygate4sd3_1 hold2674 (.A(\u_inv.f_next[139] ),
    .X(net3737));
 sg13g2_dlygate4sd3_1 hold2675 (.A(\u_inv.f_next[42] ),
    .X(net3738));
 sg13g2_dlygate4sd3_1 hold2676 (.A(\u_inv.d_next[111] ),
    .X(net3739));
 sg13g2_dlygate4sd3_1 hold2677 (.A(\u_inv.f_next[9] ),
    .X(net3740));
 sg13g2_dlygate4sd3_1 hold2678 (.A(\u_inv.counter[9] ),
    .X(net3741));
 sg13g2_dlygate4sd3_1 hold2679 (.A(_17960_),
    .X(net3742));
 sg13g2_dlygate4sd3_1 hold2680 (.A(\u_inv.counter[0] ),
    .X(net3743));
 sg13g2_dlygate4sd3_1 hold2681 (.A(_01786_),
    .X(net3744));
 sg13g2_dlygate4sd3_1 hold2682 (.A(\u_inv.f_next[118] ),
    .X(net3745));
 sg13g2_dlygate4sd3_1 hold2683 (.A(\u_inv.f_next[234] ),
    .X(net3746));
 sg13g2_dlygate4sd3_1 hold2684 (.A(\state[0] ),
    .X(net3747));
 sg13g2_dlygate4sd3_1 hold2685 (.A(_00167_),
    .X(net3748));
 sg13g2_dlygate4sd3_1 hold2686 (.A(\u_inv.counter[7] ),
    .X(net3749));
 sg13g2_dlygate4sd3_1 hold2688 (.A(net7296),
    .X(net3751));
 sg13g2_dlygate4sd3_1 hold2689 (.A(\u_inv.f_next[225] ),
    .X(net3752));
 sg13g2_dlygate4sd3_1 hold2690 (.A(\shift_reg[15] ),
    .X(net3753));
 sg13g2_dlygate4sd3_1 hold2691 (.A(\u_inv.d_next[189] ),
    .X(net3754));
 sg13g2_dlygate4sd3_1 hold2692 (.A(\state[1] ),
    .X(net3755));
 sg13g2_dlygate4sd3_1 hold2693 (.A(\u_inv.counter[2] ),
    .X(net3756));
 sg13g2_dlygate4sd3_1 hold2694 (.A(\u_inv.counter[8] ),
    .X(net3757));
 sg13g2_dlygate4sd3_1 hold2695 (.A(_17951_),
    .X(net3758));
 sg13g2_dlygate4sd3_1 hold2696 (.A(_01804_),
    .X(net3759));
 sg13g2_dlygate4sd3_1 hold2697 (.A(\u_inv.counter[6] ),
    .X(net3760));
 sg13g2_dlygate4sd3_1 hold2698 (.A(\u_inv.d_reg[137] ),
    .X(net3761));
 sg13g2_dlygate4sd3_1 hold2699 (.A(\u_inv.d_reg[157] ),
    .X(net3762));
 sg13g2_dlygate4sd3_1 hold2700 (.A(\u_inv.d_reg[201] ),
    .X(net3763));
 sg13g2_dlygate4sd3_1 hold2701 (.A(\u_inv.d_reg[123] ),
    .X(net3764));
 sg13g2_dlygate4sd3_1 hold2702 (.A(\u_inv.d_reg[43] ),
    .X(net3765));
 sg13g2_dlygate4sd3_1 hold2703 (.A(\u_inv.d_reg[87] ),
    .X(net3766));
 sg13g2_dlygate4sd3_1 hold2704 (.A(\u_inv.d_reg[207] ),
    .X(net3767));
 sg13g2_dlygate4sd3_1 hold2705 (.A(\u_inv.d_reg[195] ),
    .X(net3768));
 sg13g2_dlygate4sd3_1 hold2706 (.A(\byte_cnt[0] ),
    .X(net3769));
 sg13g2_dlygate4sd3_1 hold2707 (.A(\u_inv.d_reg[138] ),
    .X(net3770));
 sg13g2_dlygate4sd3_1 hold2708 (.A(\u_inv.d_reg[214] ),
    .X(net3771));
 sg13g2_dlygate4sd3_1 hold2709 (.A(\u_inv.d_reg[194] ),
    .X(net3772));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_4 FILLER_0_119 ();
 sg13g2_fill_1 FILLER_0_123 ();
 sg13g2_decap_8 FILLER_0_132 ();
 sg13g2_fill_2 FILLER_0_139 ();
 sg13g2_decap_8 FILLER_0_157 ();
 sg13g2_decap_8 FILLER_0_164 ();
 sg13g2_decap_8 FILLER_0_171 ();
 sg13g2_decap_8 FILLER_0_178 ();
 sg13g2_decap_8 FILLER_0_185 ();
 sg13g2_decap_8 FILLER_0_192 ();
 sg13g2_decap_8 FILLER_0_199 ();
 sg13g2_decap_8 FILLER_0_206 ();
 sg13g2_decap_8 FILLER_0_213 ();
 sg13g2_decap_8 FILLER_0_220 ();
 sg13g2_decap_8 FILLER_0_227 ();
 sg13g2_decap_8 FILLER_0_234 ();
 sg13g2_decap_8 FILLER_0_241 ();
 sg13g2_decap_8 FILLER_0_248 ();
 sg13g2_decap_8 FILLER_0_255 ();
 sg13g2_decap_8 FILLER_0_262 ();
 sg13g2_decap_8 FILLER_0_269 ();
 sg13g2_decap_8 FILLER_0_276 ();
 sg13g2_decap_8 FILLER_0_283 ();
 sg13g2_decap_8 FILLER_0_290 ();
 sg13g2_decap_8 FILLER_0_297 ();
 sg13g2_decap_4 FILLER_0_304 ();
 sg13g2_fill_2 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_323 ();
 sg13g2_decap_8 FILLER_0_330 ();
 sg13g2_decap_4 FILLER_0_337 ();
 sg13g2_fill_1 FILLER_0_341 ();
 sg13g2_decap_8 FILLER_0_360 ();
 sg13g2_fill_2 FILLER_0_367 ();
 sg13g2_fill_1 FILLER_0_369 ();
 sg13g2_decap_8 FILLER_0_374 ();
 sg13g2_decap_8 FILLER_0_381 ();
 sg13g2_decap_8 FILLER_0_388 ();
 sg13g2_decap_4 FILLER_0_395 ();
 sg13g2_fill_2 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_423 ();
 sg13g2_decap_4 FILLER_0_442 ();
 sg13g2_fill_1 FILLER_0_446 ();
 sg13g2_fill_1 FILLER_0_456 ();
 sg13g2_decap_8 FILLER_0_493 ();
 sg13g2_decap_8 FILLER_0_500 ();
 sg13g2_decap_8 FILLER_0_507 ();
 sg13g2_decap_8 FILLER_0_514 ();
 sg13g2_decap_8 FILLER_0_521 ();
 sg13g2_decap_8 FILLER_0_528 ();
 sg13g2_decap_8 FILLER_0_535 ();
 sg13g2_decap_4 FILLER_0_542 ();
 sg13g2_decap_8 FILLER_0_550 ();
 sg13g2_decap_8 FILLER_0_557 ();
 sg13g2_decap_8 FILLER_0_564 ();
 sg13g2_decap_8 FILLER_0_571 ();
 sg13g2_decap_8 FILLER_0_578 ();
 sg13g2_decap_8 FILLER_0_585 ();
 sg13g2_decap_8 FILLER_0_592 ();
 sg13g2_decap_8 FILLER_0_599 ();
 sg13g2_decap_8 FILLER_0_606 ();
 sg13g2_decap_8 FILLER_0_613 ();
 sg13g2_decap_8 FILLER_0_620 ();
 sg13g2_decap_8 FILLER_0_627 ();
 sg13g2_decap_8 FILLER_0_634 ();
 sg13g2_decap_8 FILLER_0_641 ();
 sg13g2_decap_8 FILLER_0_648 ();
 sg13g2_decap_8 FILLER_0_655 ();
 sg13g2_decap_8 FILLER_0_662 ();
 sg13g2_decap_8 FILLER_0_669 ();
 sg13g2_decap_8 FILLER_0_676 ();
 sg13g2_decap_8 FILLER_0_683 ();
 sg13g2_decap_8 FILLER_0_690 ();
 sg13g2_decap_8 FILLER_0_697 ();
 sg13g2_decap_8 FILLER_0_704 ();
 sg13g2_decap_8 FILLER_0_711 ();
 sg13g2_decap_8 FILLER_0_718 ();
 sg13g2_decap_8 FILLER_0_725 ();
 sg13g2_decap_8 FILLER_0_732 ();
 sg13g2_decap_8 FILLER_0_739 ();
 sg13g2_decap_8 FILLER_0_746 ();
 sg13g2_decap_8 FILLER_0_753 ();
 sg13g2_decap_8 FILLER_0_760 ();
 sg13g2_decap_8 FILLER_0_767 ();
 sg13g2_decap_8 FILLER_0_774 ();
 sg13g2_decap_8 FILLER_0_781 ();
 sg13g2_decap_8 FILLER_0_788 ();
 sg13g2_decap_8 FILLER_0_795 ();
 sg13g2_decap_8 FILLER_0_802 ();
 sg13g2_decap_8 FILLER_0_809 ();
 sg13g2_decap_8 FILLER_0_816 ();
 sg13g2_decap_8 FILLER_0_823 ();
 sg13g2_decap_8 FILLER_0_830 ();
 sg13g2_fill_1 FILLER_0_837 ();
 sg13g2_decap_8 FILLER_0_842 ();
 sg13g2_decap_8 FILLER_0_849 ();
 sg13g2_decap_4 FILLER_0_856 ();
 sg13g2_fill_2 FILLER_0_860 ();
 sg13g2_decap_8 FILLER_0_871 ();
 sg13g2_fill_1 FILLER_0_878 ();
 sg13g2_decap_4 FILLER_0_907 ();
 sg13g2_fill_1 FILLER_0_911 ();
 sg13g2_decap_8 FILLER_0_916 ();
 sg13g2_decap_8 FILLER_0_923 ();
 sg13g2_decap_8 FILLER_0_930 ();
 sg13g2_decap_8 FILLER_0_937 ();
 sg13g2_decap_8 FILLER_0_944 ();
 sg13g2_decap_8 FILLER_0_951 ();
 sg13g2_decap_8 FILLER_0_958 ();
 sg13g2_fill_2 FILLER_0_965 ();
 sg13g2_decap_8 FILLER_0_975 ();
 sg13g2_decap_4 FILLER_0_982 ();
 sg13g2_fill_2 FILLER_0_986 ();
 sg13g2_fill_1 FILLER_0_992 ();
 sg13g2_decap_8 FILLER_0_1001 ();
 sg13g2_fill_2 FILLER_0_1008 ();
 sg13g2_decap_8 FILLER_0_1046 ();
 sg13g2_decap_4 FILLER_0_1053 ();
 sg13g2_fill_2 FILLER_0_1057 ();
 sg13g2_fill_2 FILLER_0_1090 ();
 sg13g2_fill_1 FILLER_0_1092 ();
 sg13g2_decap_8 FILLER_0_1097 ();
 sg13g2_decap_4 FILLER_0_1104 ();
 sg13g2_fill_1 FILLER_0_1108 ();
 sg13g2_decap_8 FILLER_0_1141 ();
 sg13g2_decap_8 FILLER_0_1148 ();
 sg13g2_decap_8 FILLER_0_1155 ();
 sg13g2_decap_4 FILLER_0_1162 ();
 sg13g2_fill_2 FILLER_0_1166 ();
 sg13g2_decap_8 FILLER_0_1172 ();
 sg13g2_decap_4 FILLER_0_1179 ();
 sg13g2_fill_2 FILLER_0_1183 ();
 sg13g2_decap_4 FILLER_0_1189 ();
 sg13g2_decap_8 FILLER_0_1197 ();
 sg13g2_decap_8 FILLER_0_1204 ();
 sg13g2_decap_8 FILLER_0_1211 ();
 sg13g2_fill_1 FILLER_0_1218 ();
 sg13g2_fill_2 FILLER_0_1247 ();
 sg13g2_fill_1 FILLER_0_1249 ();
 sg13g2_fill_2 FILLER_0_1254 ();
 sg13g2_fill_2 FILLER_0_1283 ();
 sg13g2_fill_1 FILLER_0_1285 ();
 sg13g2_decap_4 FILLER_0_1296 ();
 sg13g2_decap_8 FILLER_0_1303 ();
 sg13g2_decap_8 FILLER_0_1310 ();
 sg13g2_decap_4 FILLER_0_1317 ();
 sg13g2_fill_1 FILLER_0_1321 ();
 sg13g2_decap_8 FILLER_0_1354 ();
 sg13g2_fill_1 FILLER_0_1361 ();
 sg13g2_decap_8 FILLER_0_1412 ();
 sg13g2_decap_8 FILLER_0_1419 ();
 sg13g2_fill_1 FILLER_0_1426 ();
 sg13g2_fill_1 FILLER_0_1461 ();
 sg13g2_fill_2 FILLER_0_1507 ();
 sg13g2_fill_1 FILLER_0_1509 ();
 sg13g2_fill_2 FILLER_0_1538 ();
 sg13g2_fill_1 FILLER_0_1540 ();
 sg13g2_fill_1 FILLER_0_1545 ();
 sg13g2_decap_8 FILLER_0_1550 ();
 sg13g2_decap_4 FILLER_0_1557 ();
 sg13g2_fill_2 FILLER_0_1561 ();
 sg13g2_decap_8 FILLER_0_1576 ();
 sg13g2_decap_8 FILLER_0_1583 ();
 sg13g2_decap_8 FILLER_0_1590 ();
 sg13g2_fill_2 FILLER_0_1597 ();
 sg13g2_fill_2 FILLER_0_1607 ();
 sg13g2_fill_2 FILLER_0_1631 ();
 sg13g2_fill_2 FILLER_0_1642 ();
 sg13g2_decap_8 FILLER_0_1671 ();
 sg13g2_decap_8 FILLER_0_1678 ();
 sg13g2_decap_8 FILLER_0_1685 ();
 sg13g2_fill_2 FILLER_0_1692 ();
 sg13g2_decap_4 FILLER_0_1706 ();
 sg13g2_fill_1 FILLER_0_1710 ();
 sg13g2_decap_8 FILLER_0_1715 ();
 sg13g2_decap_8 FILLER_0_1722 ();
 sg13g2_decap_8 FILLER_0_1729 ();
 sg13g2_decap_8 FILLER_0_1736 ();
 sg13g2_decap_8 FILLER_0_1743 ();
 sg13g2_decap_4 FILLER_0_1750 ();
 sg13g2_fill_2 FILLER_0_1754 ();
 sg13g2_fill_2 FILLER_0_1760 ();
 sg13g2_fill_1 FILLER_0_1762 ();
 sg13g2_decap_8 FILLER_0_1767 ();
 sg13g2_decap_8 FILLER_0_1774 ();
 sg13g2_decap_8 FILLER_0_1781 ();
 sg13g2_decap_4 FILLER_0_1788 ();
 sg13g2_fill_2 FILLER_0_1792 ();
 sg13g2_fill_2 FILLER_0_1826 ();
 sg13g2_fill_1 FILLER_0_1861 ();
 sg13g2_fill_1 FILLER_0_1889 ();
 sg13g2_fill_1 FILLER_0_1899 ();
 sg13g2_fill_2 FILLER_0_1914 ();
 sg13g2_decap_8 FILLER_0_1945 ();
 sg13g2_fill_2 FILLER_0_1952 ();
 sg13g2_decap_8 FILLER_0_1958 ();
 sg13g2_decap_8 FILLER_0_1965 ();
 sg13g2_decap_4 FILLER_0_1972 ();
 sg13g2_fill_2 FILLER_0_2002 ();
 sg13g2_fill_1 FILLER_0_2031 ();
 sg13g2_decap_8 FILLER_0_2058 ();
 sg13g2_decap_8 FILLER_0_2065 ();
 sg13g2_decap_4 FILLER_0_2072 ();
 sg13g2_fill_2 FILLER_0_2080 ();
 sg13g2_fill_1 FILLER_0_2082 ();
 sg13g2_decap_4 FILLER_0_2101 ();
 sg13g2_fill_2 FILLER_0_2133 ();
 sg13g2_fill_1 FILLER_0_2144 ();
 sg13g2_fill_2 FILLER_0_2191 ();
 sg13g2_fill_1 FILLER_0_2193 ();
 sg13g2_decap_8 FILLER_0_2198 ();
 sg13g2_decap_8 FILLER_0_2205 ();
 sg13g2_decap_8 FILLER_0_2212 ();
 sg13g2_decap_8 FILLER_0_2219 ();
 sg13g2_decap_4 FILLER_0_2226 ();
 sg13g2_fill_1 FILLER_0_2230 ();
 sg13g2_decap_8 FILLER_0_2263 ();
 sg13g2_fill_1 FILLER_0_2270 ();
 sg13g2_fill_1 FILLER_0_2299 ();
 sg13g2_decap_8 FILLER_0_2327 ();
 sg13g2_fill_2 FILLER_0_2361 ();
 sg13g2_decap_8 FILLER_0_2389 ();
 sg13g2_fill_2 FILLER_0_2396 ();
 sg13g2_decap_4 FILLER_0_2403 ();
 sg13g2_fill_1 FILLER_0_2407 ();
 sg13g2_fill_1 FILLER_0_2412 ();
 sg13g2_fill_2 FILLER_0_2444 ();
 sg13g2_fill_1 FILLER_0_2446 ();
 sg13g2_decap_8 FILLER_0_2464 ();
 sg13g2_decap_8 FILLER_0_2471 ();
 sg13g2_decap_8 FILLER_0_2478 ();
 sg13g2_fill_2 FILLER_0_2485 ();
 sg13g2_decap_8 FILLER_0_2491 ();
 sg13g2_decap_8 FILLER_0_2498 ();
 sg13g2_fill_2 FILLER_0_2505 ();
 sg13g2_fill_2 FILLER_0_2542 ();
 sg13g2_fill_2 FILLER_0_2566 ();
 sg13g2_fill_2 FILLER_0_2605 ();
 sg13g2_fill_2 FILLER_0_2625 ();
 sg13g2_fill_1 FILLER_0_2636 ();
 sg13g2_decap_8 FILLER_0_2654 ();
 sg13g2_decap_8 FILLER_0_2661 ();
 sg13g2_decap_8 FILLER_0_2668 ();
 sg13g2_decap_8 FILLER_0_2675 ();
 sg13g2_decap_8 FILLER_0_2682 ();
 sg13g2_fill_2 FILLER_0_2689 ();
 sg13g2_decap_8 FILLER_0_2699 ();
 sg13g2_decap_8 FILLER_0_2706 ();
 sg13g2_decap_8 FILLER_0_2713 ();
 sg13g2_decap_8 FILLER_0_2720 ();
 sg13g2_decap_8 FILLER_0_2727 ();
 sg13g2_fill_1 FILLER_0_2762 ();
 sg13g2_decap_4 FILLER_0_2771 ();
 sg13g2_decap_4 FILLER_0_2831 ();
 sg13g2_fill_2 FILLER_0_2835 ();
 sg13g2_decap_4 FILLER_0_2864 ();
 sg13g2_fill_1 FILLER_0_2872 ();
 sg13g2_fill_2 FILLER_0_2909 ();
 sg13g2_fill_1 FILLER_0_2911 ();
 sg13g2_fill_2 FILLER_0_2955 ();
 sg13g2_decap_8 FILLER_0_2999 ();
 sg13g2_fill_2 FILLER_0_3006 ();
 sg13g2_fill_1 FILLER_0_3008 ();
 sg13g2_decap_8 FILLER_0_3013 ();
 sg13g2_fill_2 FILLER_0_3024 ();
 sg13g2_fill_2 FILLER_0_3048 ();
 sg13g2_fill_1 FILLER_0_3059 ();
 sg13g2_fill_2 FILLER_0_3074 ();
 sg13g2_fill_1 FILLER_0_3076 ();
 sg13g2_fill_1 FILLER_0_3123 ();
 sg13g2_fill_2 FILLER_0_3133 ();
 sg13g2_fill_2 FILLER_0_3149 ();
 sg13g2_fill_1 FILLER_0_3151 ();
 sg13g2_fill_2 FILLER_0_3161 ();
 sg13g2_fill_1 FILLER_0_3163 ();
 sg13g2_fill_2 FILLER_0_3178 ();
 sg13g2_fill_2 FILLER_0_3220 ();
 sg13g2_fill_2 FILLER_0_3226 ();
 sg13g2_fill_1 FILLER_0_3228 ();
 sg13g2_decap_4 FILLER_0_3310 ();
 sg13g2_fill_1 FILLER_0_3314 ();
 sg13g2_decap_8 FILLER_0_3347 ();
 sg13g2_fill_2 FILLER_0_3354 ();
 sg13g2_fill_1 FILLER_0_3397 ();
 sg13g2_fill_2 FILLER_0_3402 ();
 sg13g2_fill_2 FILLER_0_3441 ();
 sg13g2_fill_1 FILLER_0_3443 ();
 sg13g2_fill_1 FILLER_0_3485 ();
 sg13g2_fill_2 FILLER_0_3495 ();
 sg13g2_fill_1 FILLER_0_3497 ();
 sg13g2_decap_8 FILLER_0_3515 ();
 sg13g2_decap_8 FILLER_0_3522 ();
 sg13g2_decap_8 FILLER_0_3529 ();
 sg13g2_decap_8 FILLER_0_3536 ();
 sg13g2_decap_8 FILLER_0_3543 ();
 sg13g2_decap_8 FILLER_0_3550 ();
 sg13g2_decap_8 FILLER_0_3557 ();
 sg13g2_decap_8 FILLER_0_3564 ();
 sg13g2_decap_8 FILLER_0_3571 ();
 sg13g2_fill_2 FILLER_0_3578 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_60 ();
 sg13g2_decap_8 FILLER_1_67 ();
 sg13g2_decap_8 FILLER_1_74 ();
 sg13g2_decap_8 FILLER_1_81 ();
 sg13g2_decap_8 FILLER_1_88 ();
 sg13g2_decap_8 FILLER_1_95 ();
 sg13g2_decap_4 FILLER_1_102 ();
 sg13g2_fill_1 FILLER_1_106 ();
 sg13g2_fill_2 FILLER_1_111 ();
 sg13g2_fill_2 FILLER_1_126 ();
 sg13g2_fill_1 FILLER_1_128 ();
 sg13g2_decap_8 FILLER_1_162 ();
 sg13g2_decap_8 FILLER_1_169 ();
 sg13g2_decap_8 FILLER_1_176 ();
 sg13g2_decap_8 FILLER_1_183 ();
 sg13g2_decap_8 FILLER_1_190 ();
 sg13g2_decap_8 FILLER_1_197 ();
 sg13g2_decap_8 FILLER_1_204 ();
 sg13g2_decap_8 FILLER_1_211 ();
 sg13g2_decap_8 FILLER_1_218 ();
 sg13g2_decap_8 FILLER_1_225 ();
 sg13g2_decap_8 FILLER_1_232 ();
 sg13g2_decap_8 FILLER_1_239 ();
 sg13g2_decap_8 FILLER_1_246 ();
 sg13g2_decap_8 FILLER_1_253 ();
 sg13g2_decap_8 FILLER_1_260 ();
 sg13g2_decap_8 FILLER_1_267 ();
 sg13g2_decap_8 FILLER_1_274 ();
 sg13g2_decap_8 FILLER_1_281 ();
 sg13g2_fill_2 FILLER_1_288 ();
 sg13g2_fill_1 FILLER_1_308 ();
 sg13g2_fill_2 FILLER_1_393 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_fill_1 FILLER_1_407 ();
 sg13g2_fill_1 FILLER_1_464 ();
 sg13g2_fill_2 FILLER_1_474 ();
 sg13g2_fill_2 FILLER_1_485 ();
 sg13g2_fill_1 FILLER_1_487 ();
 sg13g2_decap_8 FILLER_1_501 ();
 sg13g2_decap_8 FILLER_1_508 ();
 sg13g2_decap_8 FILLER_1_515 ();
 sg13g2_fill_1 FILLER_1_522 ();
 sg13g2_decap_8 FILLER_1_559 ();
 sg13g2_decap_8 FILLER_1_566 ();
 sg13g2_decap_8 FILLER_1_573 ();
 sg13g2_decap_8 FILLER_1_580 ();
 sg13g2_decap_8 FILLER_1_587 ();
 sg13g2_decap_8 FILLER_1_594 ();
 sg13g2_decap_8 FILLER_1_601 ();
 sg13g2_decap_8 FILLER_1_608 ();
 sg13g2_decap_8 FILLER_1_615 ();
 sg13g2_decap_8 FILLER_1_622 ();
 sg13g2_decap_8 FILLER_1_629 ();
 sg13g2_decap_8 FILLER_1_636 ();
 sg13g2_decap_8 FILLER_1_643 ();
 sg13g2_decap_8 FILLER_1_650 ();
 sg13g2_decap_8 FILLER_1_657 ();
 sg13g2_fill_2 FILLER_1_664 ();
 sg13g2_decap_8 FILLER_1_670 ();
 sg13g2_decap_8 FILLER_1_677 ();
 sg13g2_decap_8 FILLER_1_684 ();
 sg13g2_decap_8 FILLER_1_691 ();
 sg13g2_decap_8 FILLER_1_698 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_fill_2 FILLER_1_861 ();
 sg13g2_fill_1 FILLER_1_863 ();
 sg13g2_fill_1 FILLER_1_873 ();
 sg13g2_fill_2 FILLER_1_896 ();
 sg13g2_decap_8 FILLER_1_935 ();
 sg13g2_fill_1 FILLER_1_942 ();
 sg13g2_decap_4 FILLER_1_947 ();
 sg13g2_fill_1 FILLER_1_951 ();
 sg13g2_fill_1 FILLER_1_956 ();
 sg13g2_fill_2 FILLER_1_1062 ();
 sg13g2_fill_2 FILLER_1_1078 ();
 sg13g2_decap_8 FILLER_1_1142 ();
 sg13g2_decap_4 FILLER_1_1149 ();
 sg13g2_fill_2 FILLER_1_1156 ();
 sg13g2_fill_1 FILLER_1_1158 ();
 sg13g2_fill_2 FILLER_1_1187 ();
 sg13g2_fill_1 FILLER_1_1189 ();
 sg13g2_fill_2 FILLER_1_1195 ();
 sg13g2_decap_4 FILLER_1_1208 ();
 sg13g2_fill_2 FILLER_1_1212 ();
 sg13g2_fill_1 FILLER_1_1244 ();
 sg13g2_fill_2 FILLER_1_1259 ();
 sg13g2_decap_4 FILLER_1_1265 ();
 sg13g2_decap_4 FILLER_1_1292 ();
 sg13g2_decap_4 FILLER_1_1309 ();
 sg13g2_fill_2 FILLER_1_1313 ();
 sg13g2_fill_2 FILLER_1_1323 ();
 sg13g2_fill_1 FILLER_1_1325 ();
 sg13g2_fill_2 FILLER_1_1335 ();
 sg13g2_fill_1 FILLER_1_1337 ();
 sg13g2_fill_1 FILLER_1_1351 ();
 sg13g2_fill_2 FILLER_1_1386 ();
 sg13g2_fill_1 FILLER_1_1388 ();
 sg13g2_fill_2 FILLER_1_1393 ();
 sg13g2_fill_2 FILLER_1_1404 ();
 sg13g2_fill_1 FILLER_1_1419 ();
 sg13g2_fill_1 FILLER_1_1476 ();
 sg13g2_fill_2 FILLER_1_1655 ();
 sg13g2_fill_1 FILLER_1_1657 ();
 sg13g2_fill_1 FILLER_1_1667 ();
 sg13g2_fill_1 FILLER_1_1695 ();
 sg13g2_decap_8 FILLER_1_1729 ();
 sg13g2_decap_8 FILLER_1_1736 ();
 sg13g2_decap_8 FILLER_1_1743 ();
 sg13g2_fill_1 FILLER_1_1750 ();
 sg13g2_fill_2 FILLER_1_1816 ();
 sg13g2_fill_2 FILLER_1_1835 ();
 sg13g2_fill_1 FILLER_1_1837 ();
 sg13g2_fill_1 FILLER_1_1869 ();
 sg13g2_decap_4 FILLER_1_2066 ();
 sg13g2_fill_1 FILLER_1_2070 ();
 sg13g2_decap_8 FILLER_1_2116 ();
 sg13g2_decap_8 FILLER_1_2181 ();
 sg13g2_fill_1 FILLER_1_2188 ();
 sg13g2_fill_2 FILLER_1_2217 ();
 sg13g2_fill_1 FILLER_1_2219 ();
 sg13g2_fill_2 FILLER_1_2242 ();
 sg13g2_fill_2 FILLER_1_2266 ();
 sg13g2_fill_1 FILLER_1_2268 ();
 sg13g2_fill_1 FILLER_1_2291 ();
 sg13g2_fill_1 FILLER_1_2301 ();
 sg13g2_decap_8 FILLER_1_2329 ();
 sg13g2_fill_2 FILLER_1_2336 ();
 sg13g2_fill_2 FILLER_1_2366 ();
 sg13g2_fill_2 FILLER_1_2401 ();
 sg13g2_fill_1 FILLER_1_2431 ();
 sg13g2_decap_4 FILLER_1_2460 ();
 sg13g2_fill_2 FILLER_1_2464 ();
 sg13g2_decap_8 FILLER_1_2470 ();
 sg13g2_decap_4 FILLER_1_2477 ();
 sg13g2_fill_1 FILLER_1_2481 ();
 sg13g2_fill_2 FILLER_1_2528 ();
 sg13g2_fill_1 FILLER_1_2543 ();
 sg13g2_fill_2 FILLER_1_2576 ();
 sg13g2_fill_1 FILLER_1_2578 ();
 sg13g2_fill_2 FILLER_1_2672 ();
 sg13g2_fill_1 FILLER_1_2674 ();
 sg13g2_decap_8 FILLER_1_2716 ();
 sg13g2_decap_4 FILLER_1_2723 ();
 sg13g2_fill_1 FILLER_1_2727 ();
 sg13g2_fill_2 FILLER_1_2750 ();
 sg13g2_fill_1 FILLER_1_2770 ();
 sg13g2_fill_2 FILLER_1_2776 ();
 sg13g2_fill_1 FILLER_1_2791 ();
 sg13g2_fill_1 FILLER_1_2818 ();
 sg13g2_fill_1 FILLER_1_2832 ();
 sg13g2_fill_1 FILLER_1_2838 ();
 sg13g2_fill_1 FILLER_1_2861 ();
 sg13g2_fill_2 FILLER_1_2875 ();
 sg13g2_fill_1 FILLER_1_2886 ();
 sg13g2_fill_2 FILLER_1_2920 ();
 sg13g2_fill_1 FILLER_1_2931 ();
 sg13g2_fill_1 FILLER_1_2986 ();
 sg13g2_decap_4 FILLER_1_3000 ();
 sg13g2_fill_2 FILLER_1_3088 ();
 sg13g2_fill_1 FILLER_1_3378 ();
 sg13g2_fill_2 FILLER_1_3407 ();
 sg13g2_fill_2 FILLER_1_3441 ();
 sg13g2_decap_8 FILLER_1_3530 ();
 sg13g2_fill_1 FILLER_1_3537 ();
 sg13g2_fill_1 FILLER_1_3542 ();
 sg13g2_decap_8 FILLER_1_3569 ();
 sg13g2_decap_4 FILLER_1_3576 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_4 FILLER_2_35 ();
 sg13g2_fill_2 FILLER_2_39 ();
 sg13g2_fill_2 FILLER_2_59 ();
 sg13g2_fill_1 FILLER_2_61 ();
 sg13g2_decap_8 FILLER_2_71 ();
 sg13g2_decap_8 FILLER_2_78 ();
 sg13g2_decap_8 FILLER_2_85 ();
 sg13g2_decap_8 FILLER_2_92 ();
 sg13g2_fill_2 FILLER_2_99 ();
 sg13g2_fill_1 FILLER_2_101 ();
 sg13g2_fill_2 FILLER_2_130 ();
 sg13g2_fill_2 FILLER_2_160 ();
 sg13g2_fill_2 FILLER_2_172 ();
 sg13g2_fill_1 FILLER_2_174 ();
 sg13g2_decap_8 FILLER_2_180 ();
 sg13g2_decap_8 FILLER_2_187 ();
 sg13g2_decap_8 FILLER_2_194 ();
 sg13g2_decap_8 FILLER_2_201 ();
 sg13g2_decap_8 FILLER_2_208 ();
 sg13g2_decap_8 FILLER_2_215 ();
 sg13g2_decap_8 FILLER_2_222 ();
 sg13g2_decap_8 FILLER_2_229 ();
 sg13g2_decap_8 FILLER_2_236 ();
 sg13g2_decap_8 FILLER_2_243 ();
 sg13g2_decap_8 FILLER_2_250 ();
 sg13g2_decap_8 FILLER_2_257 ();
 sg13g2_decap_8 FILLER_2_264 ();
 sg13g2_decap_4 FILLER_2_271 ();
 sg13g2_fill_2 FILLER_2_312 ();
 sg13g2_fill_1 FILLER_2_314 ();
 sg13g2_fill_2 FILLER_2_324 ();
 sg13g2_fill_1 FILLER_2_339 ();
 sg13g2_decap_4 FILLER_2_365 ();
 sg13g2_fill_1 FILLER_2_369 ();
 sg13g2_fill_1 FILLER_2_373 ();
 sg13g2_fill_1 FILLER_2_389 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_fill_1 FILLER_2_444 ();
 sg13g2_fill_2 FILLER_2_458 ();
 sg13g2_fill_2 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_503 ();
 sg13g2_decap_8 FILLER_2_510 ();
 sg13g2_fill_1 FILLER_2_517 ();
 sg13g2_fill_1 FILLER_2_523 ();
 sg13g2_fill_2 FILLER_2_547 ();
 sg13g2_fill_2 FILLER_2_558 ();
 sg13g2_decap_8 FILLER_2_564 ();
 sg13g2_decap_8 FILLER_2_571 ();
 sg13g2_fill_1 FILLER_2_582 ();
 sg13g2_fill_2 FILLER_2_611 ();
 sg13g2_decap_8 FILLER_2_617 ();
 sg13g2_decap_4 FILLER_2_624 ();
 sg13g2_fill_2 FILLER_2_628 ();
 sg13g2_decap_8 FILLER_2_634 ();
 sg13g2_decap_8 FILLER_2_641 ();
 sg13g2_decap_8 FILLER_2_648 ();
 sg13g2_decap_4 FILLER_2_655 ();
 sg13g2_fill_1 FILLER_2_659 ();
 sg13g2_decap_8 FILLER_2_724 ();
 sg13g2_decap_8 FILLER_2_731 ();
 sg13g2_fill_2 FILLER_2_738 ();
 sg13g2_decap_4 FILLER_2_744 ();
 sg13g2_fill_1 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_766 ();
 sg13g2_decap_8 FILLER_2_773 ();
 sg13g2_decap_8 FILLER_2_780 ();
 sg13g2_decap_8 FILLER_2_787 ();
 sg13g2_decap_8 FILLER_2_794 ();
 sg13g2_decap_8 FILLER_2_801 ();
 sg13g2_decap_8 FILLER_2_808 ();
 sg13g2_decap_8 FILLER_2_815 ();
 sg13g2_decap_8 FILLER_2_822 ();
 sg13g2_decap_8 FILLER_2_829 ();
 sg13g2_fill_2 FILLER_2_836 ();
 sg13g2_decap_8 FILLER_2_874 ();
 sg13g2_fill_2 FILLER_2_898 ();
 sg13g2_fill_2 FILLER_2_922 ();
 sg13g2_fill_1 FILLER_2_924 ();
 sg13g2_fill_2 FILLER_2_953 ();
 sg13g2_fill_1 FILLER_2_955 ();
 sg13g2_fill_1 FILLER_2_987 ();
 sg13g2_fill_1 FILLER_2_1002 ();
 sg13g2_fill_1 FILLER_2_1017 ();
 sg13g2_fill_1 FILLER_2_1040 ();
 sg13g2_decap_4 FILLER_2_1046 ();
 sg13g2_fill_2 FILLER_2_1050 ();
 sg13g2_fill_2 FILLER_2_1057 ();
 sg13g2_fill_1 FILLER_2_1059 ();
 sg13g2_fill_2 FILLER_2_1086 ();
 sg13g2_fill_1 FILLER_2_1088 ();
 sg13g2_decap_8 FILLER_2_1098 ();
 sg13g2_fill_2 FILLER_2_1105 ();
 sg13g2_fill_1 FILLER_2_1107 ();
 sg13g2_fill_1 FILLER_2_1121 ();
 sg13g2_fill_2 FILLER_2_1153 ();
 sg13g2_fill_2 FILLER_2_1169 ();
 sg13g2_fill_1 FILLER_2_1171 ();
 sg13g2_fill_1 FILLER_2_1185 ();
 sg13g2_decap_8 FILLER_2_1215 ();
 sg13g2_decap_4 FILLER_2_1257 ();
 sg13g2_fill_1 FILLER_2_1261 ();
 sg13g2_fill_1 FILLER_2_1275 ();
 sg13g2_fill_2 FILLER_2_1280 ();
 sg13g2_fill_2 FILLER_2_1290 ();
 sg13g2_fill_1 FILLER_2_1306 ();
 sg13g2_decap_4 FILLER_2_1316 ();
 sg13g2_fill_2 FILLER_2_1361 ();
 sg13g2_fill_1 FILLER_2_1363 ();
 sg13g2_fill_2 FILLER_2_1440 ();
 sg13g2_fill_1 FILLER_2_1442 ();
 sg13g2_fill_2 FILLER_2_1452 ();
 sg13g2_fill_1 FILLER_2_1454 ();
 sg13g2_fill_2 FILLER_2_1463 ();
 sg13g2_fill_1 FILLER_2_1477 ();
 sg13g2_fill_1 FILLER_2_1515 ();
 sg13g2_fill_1 FILLER_2_1549 ();
 sg13g2_fill_2 FILLER_2_1614 ();
 sg13g2_decap_8 FILLER_2_1630 ();
 sg13g2_fill_1 FILLER_2_1637 ();
 sg13g2_fill_1 FILLER_2_1651 ();
 sg13g2_decap_4 FILLER_2_1661 ();
 sg13g2_fill_1 FILLER_2_1665 ();
 sg13g2_fill_2 FILLER_2_1697 ();
 sg13g2_fill_1 FILLER_2_1699 ();
 sg13g2_fill_2 FILLER_2_1714 ();
 sg13g2_fill_2 FILLER_2_1725 ();
 sg13g2_fill_1 FILLER_2_1727 ();
 sg13g2_fill_2 FILLER_2_1819 ();
 sg13g2_fill_1 FILLER_2_1821 ();
 sg13g2_fill_2 FILLER_2_1850 ();
 sg13g2_fill_2 FILLER_2_1874 ();
 sg13g2_fill_1 FILLER_2_1876 ();
 sg13g2_fill_2 FILLER_2_1913 ();
 sg13g2_decap_4 FILLER_2_1961 ();
 sg13g2_fill_1 FILLER_2_1965 ();
 sg13g2_fill_2 FILLER_2_1979 ();
 sg13g2_fill_1 FILLER_2_1981 ();
 sg13g2_fill_2 FILLER_2_2013 ();
 sg13g2_fill_1 FILLER_2_2015 ();
 sg13g2_fill_2 FILLER_2_2034 ();
 sg13g2_fill_1 FILLER_2_2036 ();
 sg13g2_decap_8 FILLER_2_2075 ();
 sg13g2_fill_2 FILLER_2_2082 ();
 sg13g2_fill_1 FILLER_2_2084 ();
 sg13g2_decap_4 FILLER_2_2108 ();
 sg13g2_fill_2 FILLER_2_2122 ();
 sg13g2_fill_1 FILLER_2_2129 ();
 sg13g2_fill_2 FILLER_2_2169 ();
 sg13g2_fill_1 FILLER_2_2171 ();
 sg13g2_decap_8 FILLER_2_2176 ();
 sg13g2_decap_8 FILLER_2_2188 ();
 sg13g2_decap_4 FILLER_2_2195 ();
 sg13g2_decap_4 FILLER_2_2216 ();
 sg13g2_fill_2 FILLER_2_2220 ();
 sg13g2_fill_2 FILLER_2_2281 ();
 sg13g2_fill_1 FILLER_2_2283 ();
 sg13g2_fill_2 FILLER_2_2292 ();
 sg13g2_fill_1 FILLER_2_2312 ();
 sg13g2_fill_2 FILLER_2_2367 ();
 sg13g2_fill_1 FILLER_2_2426 ();
 sg13g2_fill_2 FILLER_2_2448 ();
 sg13g2_fill_1 FILLER_2_2459 ();
 sg13g2_fill_2 FILLER_2_2514 ();
 sg13g2_decap_8 FILLER_2_2542 ();
 sg13g2_decap_4 FILLER_2_2549 ();
 sg13g2_fill_1 FILLER_2_2583 ();
 sg13g2_fill_2 FILLER_2_2612 ();
 sg13g2_fill_2 FILLER_2_2623 ();
 sg13g2_fill_1 FILLER_2_2625 ();
 sg13g2_fill_1 FILLER_2_2638 ();
 sg13g2_fill_1 FILLER_2_2653 ();
 sg13g2_decap_4 FILLER_2_2721 ();
 sg13g2_fill_1 FILLER_2_2725 ();
 sg13g2_fill_2 FILLER_2_2742 ();
 sg13g2_decap_8 FILLER_2_2766 ();
 sg13g2_fill_1 FILLER_2_2773 ();
 sg13g2_fill_2 FILLER_2_2787 ();
 sg13g2_decap_4 FILLER_2_2806 ();
 sg13g2_decap_8 FILLER_2_2847 ();
 sg13g2_fill_1 FILLER_2_2854 ();
 sg13g2_fill_1 FILLER_2_2954 ();
 sg13g2_decap_8 FILLER_2_2972 ();
 sg13g2_fill_2 FILLER_2_2979 ();
 sg13g2_fill_2 FILLER_2_3036 ();
 sg13g2_fill_1 FILLER_2_3038 ();
 sg13g2_fill_1 FILLER_2_3043 ();
 sg13g2_decap_4 FILLER_2_3052 ();
 sg13g2_fill_1 FILLER_2_3056 ();
 sg13g2_fill_2 FILLER_2_3077 ();
 sg13g2_fill_1 FILLER_2_3079 ();
 sg13g2_fill_2 FILLER_2_3093 ();
 sg13g2_fill_1 FILLER_2_3095 ();
 sg13g2_decap_4 FILLER_2_3121 ();
 sg13g2_fill_2 FILLER_2_3130 ();
 sg13g2_fill_1 FILLER_2_3132 ();
 sg13g2_fill_2 FILLER_2_3141 ();
 sg13g2_fill_2 FILLER_2_3147 ();
 sg13g2_decap_8 FILLER_2_3153 ();
 sg13g2_fill_2 FILLER_2_3160 ();
 sg13g2_fill_2 FILLER_2_3174 ();
 sg13g2_fill_1 FILLER_2_3198 ();
 sg13g2_fill_2 FILLER_2_3270 ();
 sg13g2_fill_1 FILLER_2_3272 ();
 sg13g2_fill_1 FILLER_2_3291 ();
 sg13g2_fill_2 FILLER_2_3335 ();
 sg13g2_fill_1 FILLER_2_3337 ();
 sg13g2_fill_2 FILLER_2_3351 ();
 sg13g2_fill_1 FILLER_2_3353 ();
 sg13g2_fill_1 FILLER_2_3380 ();
 sg13g2_fill_1 FILLER_2_3413 ();
 sg13g2_fill_1 FILLER_2_3460 ();
 sg13g2_fill_1 FILLER_2_3492 ();
 sg13g2_fill_2 FILLER_2_3540 ();
 sg13g2_decap_4 FILLER_2_3575 ();
 sg13g2_fill_1 FILLER_2_3579 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_fill_1 FILLER_3_21 ();
 sg13g2_fill_2 FILLER_3_31 ();
 sg13g2_decap_4 FILLER_3_38 ();
 sg13g2_fill_1 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_75 ();
 sg13g2_fill_1 FILLER_3_124 ();
 sg13g2_fill_1 FILLER_3_142 ();
 sg13g2_fill_2 FILLER_3_185 ();
 sg13g2_decap_8 FILLER_3_200 ();
 sg13g2_decap_8 FILLER_3_207 ();
 sg13g2_decap_4 FILLER_3_214 ();
 sg13g2_fill_2 FILLER_3_218 ();
 sg13g2_decap_8 FILLER_3_228 ();
 sg13g2_decap_8 FILLER_3_235 ();
 sg13g2_decap_8 FILLER_3_242 ();
 sg13g2_decap_8 FILLER_3_249 ();
 sg13g2_decap_8 FILLER_3_256 ();
 sg13g2_decap_8 FILLER_3_263 ();
 sg13g2_decap_8 FILLER_3_270 ();
 sg13g2_fill_2 FILLER_3_277 ();
 sg13g2_fill_1 FILLER_3_279 ();
 sg13g2_decap_8 FILLER_3_284 ();
 sg13g2_decap_4 FILLER_3_291 ();
 sg13g2_fill_1 FILLER_3_295 ();
 sg13g2_decap_4 FILLER_3_300 ();
 sg13g2_fill_1 FILLER_3_304 ();
 sg13g2_fill_2 FILLER_3_313 ();
 sg13g2_fill_1 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_338 ();
 sg13g2_decap_4 FILLER_3_345 ();
 sg13g2_fill_1 FILLER_3_349 ();
 sg13g2_fill_1 FILLER_3_365 ();
 sg13g2_fill_1 FILLER_3_381 ();
 sg13g2_decap_8 FILLER_3_403 ();
 sg13g2_decap_4 FILLER_3_410 ();
 sg13g2_fill_2 FILLER_3_451 ();
 sg13g2_fill_1 FILLER_3_453 ();
 sg13g2_decap_4 FILLER_3_485 ();
 sg13g2_fill_1 FILLER_3_489 ();
 sg13g2_fill_1 FILLER_3_508 ();
 sg13g2_fill_1 FILLER_3_541 ();
 sg13g2_fill_2 FILLER_3_583 ();
 sg13g2_fill_1 FILLER_3_585 ();
 sg13g2_fill_2 FILLER_3_664 ();
 sg13g2_fill_2 FILLER_3_684 ();
 sg13g2_fill_1 FILLER_3_686 ();
 sg13g2_fill_2 FILLER_3_696 ();
 sg13g2_fill_1 FILLER_3_698 ();
 sg13g2_fill_2 FILLER_3_708 ();
 sg13g2_fill_1 FILLER_3_710 ();
 sg13g2_fill_2 FILLER_3_729 ();
 sg13g2_fill_2 FILLER_3_772 ();
 sg13g2_fill_1 FILLER_3_774 ();
 sg13g2_fill_1 FILLER_3_784 ();
 sg13g2_fill_2 FILLER_3_794 ();
 sg13g2_fill_1 FILLER_3_796 ();
 sg13g2_decap_8 FILLER_3_801 ();
 sg13g2_decap_8 FILLER_3_808 ();
 sg13g2_decap_8 FILLER_3_815 ();
 sg13g2_decap_8 FILLER_3_822 ();
 sg13g2_fill_1 FILLER_3_829 ();
 sg13g2_fill_2 FILLER_3_843 ();
 sg13g2_fill_1 FILLER_3_863 ();
 sg13g2_fill_2 FILLER_3_881 ();
 sg13g2_fill_1 FILLER_3_890 ();
 sg13g2_fill_2 FILLER_3_936 ();
 sg13g2_fill_2 FILLER_3_966 ();
 sg13g2_fill_1 FILLER_3_968 ();
 sg13g2_fill_2 FILLER_3_986 ();
 sg13g2_fill_1 FILLER_3_1009 ();
 sg13g2_fill_2 FILLER_3_1035 ();
 sg13g2_fill_2 FILLER_3_1069 ();
 sg13g2_decap_8 FILLER_3_1105 ();
 sg13g2_decap_8 FILLER_3_1112 ();
 sg13g2_decap_8 FILLER_3_1146 ();
 sg13g2_decap_8 FILLER_3_1153 ();
 sg13g2_fill_2 FILLER_3_1160 ();
 sg13g2_fill_1 FILLER_3_1162 ();
 sg13g2_fill_2 FILLER_3_1168 ();
 sg13g2_fill_1 FILLER_3_1170 ();
 sg13g2_fill_2 FILLER_3_1189 ();
 sg13g2_fill_1 FILLER_3_1191 ();
 sg13g2_fill_1 FILLER_3_1204 ();
 sg13g2_fill_2 FILLER_3_1216 ();
 sg13g2_decap_4 FILLER_3_1222 ();
 sg13g2_decap_4 FILLER_3_1231 ();
 sg13g2_fill_2 FILLER_3_1235 ();
 sg13g2_decap_4 FILLER_3_1296 ();
 sg13g2_fill_1 FILLER_3_1300 ();
 sg13g2_decap_4 FILLER_3_1346 ();
 sg13g2_fill_2 FILLER_3_1350 ();
 sg13g2_decap_4 FILLER_3_1361 ();
 sg13g2_fill_2 FILLER_3_1378 ();
 sg13g2_fill_1 FILLER_3_1393 ();
 sg13g2_decap_4 FILLER_3_1421 ();
 sg13g2_fill_2 FILLER_3_1425 ();
 sg13g2_fill_1 FILLER_3_1440 ();
 sg13g2_fill_2 FILLER_3_1492 ();
 sg13g2_fill_1 FILLER_3_1494 ();
 sg13g2_fill_2 FILLER_3_1500 ();
 sg13g2_fill_2 FILLER_3_1555 ();
 sg13g2_fill_1 FILLER_3_1557 ();
 sg13g2_fill_2 FILLER_3_1609 ();
 sg13g2_fill_1 FILLER_3_1611 ();
 sg13g2_fill_2 FILLER_3_1633 ();
 sg13g2_fill_1 FILLER_3_1635 ();
 sg13g2_decap_8 FILLER_3_1666 ();
 sg13g2_decap_4 FILLER_3_1673 ();
 sg13g2_fill_2 FILLER_3_1677 ();
 sg13g2_fill_2 FILLER_3_1683 ();
 sg13g2_fill_1 FILLER_3_1712 ();
 sg13g2_decap_4 FILLER_3_1721 ();
 sg13g2_fill_2 FILLER_3_1725 ();
 sg13g2_fill_1 FILLER_3_1753 ();
 sg13g2_fill_2 FILLER_3_1776 ();
 sg13g2_fill_1 FILLER_3_1778 ();
 sg13g2_fill_2 FILLER_3_1796 ();
 sg13g2_fill_1 FILLER_3_1798 ();
 sg13g2_fill_1 FILLER_3_1804 ();
 sg13g2_fill_2 FILLER_3_1822 ();
 sg13g2_fill_2 FILLER_3_1849 ();
 sg13g2_fill_1 FILLER_3_1851 ();
 sg13g2_fill_2 FILLER_3_1917 ();
 sg13g2_fill_2 FILLER_3_1961 ();
 sg13g2_fill_2 FILLER_3_1991 ();
 sg13g2_fill_1 FILLER_3_1993 ();
 sg13g2_fill_1 FILLER_3_1999 ();
 sg13g2_fill_1 FILLER_3_2008 ();
 sg13g2_fill_1 FILLER_3_2039 ();
 sg13g2_decap_4 FILLER_3_2060 ();
 sg13g2_fill_1 FILLER_3_2108 ();
 sg13g2_fill_2 FILLER_3_2144 ();
 sg13g2_fill_2 FILLER_3_2158 ();
 sg13g2_decap_4 FILLER_3_2192 ();
 sg13g2_fill_1 FILLER_3_2218 ();
 sg13g2_fill_1 FILLER_3_2270 ();
 sg13g2_decap_4 FILLER_3_2278 ();
 sg13g2_fill_2 FILLER_3_2297 ();
 sg13g2_fill_1 FILLER_3_2299 ();
 sg13g2_fill_1 FILLER_3_2329 ();
 sg13g2_fill_2 FILLER_3_2348 ();
 sg13g2_fill_1 FILLER_3_2350 ();
 sg13g2_fill_2 FILLER_3_2364 ();
 sg13g2_fill_1 FILLER_3_2383 ();
 sg13g2_fill_1 FILLER_3_2389 ();
 sg13g2_fill_2 FILLER_3_2422 ();
 sg13g2_fill_1 FILLER_3_2432 ();
 sg13g2_fill_2 FILLER_3_2464 ();
 sg13g2_decap_8 FILLER_3_2482 ();
 sg13g2_fill_2 FILLER_3_2522 ();
 sg13g2_fill_1 FILLER_3_2524 ();
 sg13g2_fill_2 FILLER_3_2530 ();
 sg13g2_fill_1 FILLER_3_2541 ();
 sg13g2_fill_2 FILLER_3_2569 ();
 sg13g2_fill_1 FILLER_3_2571 ();
 sg13g2_fill_2 FILLER_3_2577 ();
 sg13g2_fill_1 FILLER_3_2584 ();
 sg13g2_fill_1 FILLER_3_2590 ();
 sg13g2_fill_1 FILLER_3_2608 ();
 sg13g2_decap_8 FILLER_3_2622 ();
 sg13g2_fill_2 FILLER_3_2629 ();
 sg13g2_fill_2 FILLER_3_2640 ();
 sg13g2_fill_1 FILLER_3_2659 ();
 sg13g2_fill_2 FILLER_3_2665 ();
 sg13g2_fill_1 FILLER_3_2700 ();
 sg13g2_fill_2 FILLER_3_2734 ();
 sg13g2_fill_2 FILLER_3_2744 ();
 sg13g2_fill_1 FILLER_3_2746 ();
 sg13g2_decap_8 FILLER_3_2759 ();
 sg13g2_fill_2 FILLER_3_2766 ();
 sg13g2_fill_2 FILLER_3_2776 ();
 sg13g2_fill_1 FILLER_3_2778 ();
 sg13g2_fill_2 FILLER_3_2789 ();
 sg13g2_decap_4 FILLER_3_2813 ();
 sg13g2_fill_2 FILLER_3_2817 ();
 sg13g2_fill_2 FILLER_3_2822 ();
 sg13g2_decap_8 FILLER_3_2828 ();
 sg13g2_fill_2 FILLER_3_2844 ();
 sg13g2_fill_1 FILLER_3_2846 ();
 sg13g2_decap_4 FILLER_3_2866 ();
 sg13g2_decap_4 FILLER_3_2875 ();
 sg13g2_fill_2 FILLER_3_2887 ();
 sg13g2_fill_1 FILLER_3_2889 ();
 sg13g2_fill_1 FILLER_3_2943 ();
 sg13g2_decap_8 FILLER_3_2960 ();
 sg13g2_fill_2 FILLER_3_2975 ();
 sg13g2_fill_2 FILLER_3_3004 ();
 sg13g2_fill_2 FILLER_3_3033 ();
 sg13g2_fill_1 FILLER_3_3035 ();
 sg13g2_decap_4 FILLER_3_3053 ();
 sg13g2_fill_1 FILLER_3_3057 ();
 sg13g2_decap_8 FILLER_3_3079 ();
 sg13g2_fill_2 FILLER_3_3086 ();
 sg13g2_decap_4 FILLER_3_3099 ();
 sg13g2_fill_1 FILLER_3_3103 ();
 sg13g2_fill_2 FILLER_3_3121 ();
 sg13g2_fill_2 FILLER_3_3141 ();
 sg13g2_fill_1 FILLER_3_3143 ();
 sg13g2_decap_4 FILLER_3_3172 ();
 sg13g2_fill_1 FILLER_3_3176 ();
 sg13g2_fill_2 FILLER_3_3205 ();
 sg13g2_fill_2 FILLER_3_3212 ();
 sg13g2_fill_2 FILLER_3_3243 ();
 sg13g2_fill_2 FILLER_3_3258 ();
 sg13g2_fill_1 FILLER_3_3276 ();
 sg13g2_fill_2 FILLER_3_3290 ();
 sg13g2_fill_1 FILLER_3_3292 ();
 sg13g2_fill_2 FILLER_3_3318 ();
 sg13g2_fill_1 FILLER_3_3320 ();
 sg13g2_fill_1 FILLER_3_3342 ();
 sg13g2_fill_2 FILLER_3_3351 ();
 sg13g2_fill_1 FILLER_3_3353 ();
 sg13g2_fill_2 FILLER_3_3377 ();
 sg13g2_fill_1 FILLER_3_3403 ();
 sg13g2_fill_2 FILLER_3_3428 ();
 sg13g2_fill_1 FILLER_3_3430 ();
 sg13g2_fill_1 FILLER_3_3448 ();
 sg13g2_decap_4 FILLER_3_3486 ();
 sg13g2_fill_1 FILLER_3_3490 ();
 sg13g2_fill_2 FILLER_3_3503 ();
 sg13g2_fill_2 FILLER_3_3536 ();
 sg13g2_fill_1 FILLER_3_3538 ();
 sg13g2_decap_4 FILLER_3_3552 ();
 sg13g2_fill_2 FILLER_3_3556 ();
 sg13g2_decap_8 FILLER_3_3571 ();
 sg13g2_fill_2 FILLER_3_3578 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_fill_2 FILLER_4_7 ();
 sg13g2_decap_4 FILLER_4_71 ();
 sg13g2_fill_1 FILLER_4_75 ();
 sg13g2_decap_4 FILLER_4_81 ();
 sg13g2_fill_2 FILLER_4_85 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_fill_1 FILLER_4_98 ();
 sg13g2_fill_2 FILLER_4_136 ();
 sg13g2_fill_1 FILLER_4_138 ();
 sg13g2_fill_2 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_176 ();
 sg13g2_fill_2 FILLER_4_193 ();
 sg13g2_fill_1 FILLER_4_195 ();
 sg13g2_decap_4 FILLER_4_201 ();
 sg13g2_fill_1 FILLER_4_205 ();
 sg13g2_decap_8 FILLER_4_211 ();
 sg13g2_fill_2 FILLER_4_218 ();
 sg13g2_fill_1 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_247 ();
 sg13g2_decap_8 FILLER_4_254 ();
 sg13g2_decap_8 FILLER_4_261 ();
 sg13g2_fill_2 FILLER_4_268 ();
 sg13g2_fill_1 FILLER_4_298 ();
 sg13g2_fill_1 FILLER_4_309 ();
 sg13g2_decap_8 FILLER_4_324 ();
 sg13g2_decap_4 FILLER_4_331 ();
 sg13g2_fill_2 FILLER_4_352 ();
 sg13g2_fill_1 FILLER_4_359 ();
 sg13g2_decap_4 FILLER_4_368 ();
 sg13g2_fill_2 FILLER_4_372 ();
 sg13g2_fill_2 FILLER_4_377 ();
 sg13g2_fill_1 FILLER_4_379 ();
 sg13g2_decap_4 FILLER_4_413 ();
 sg13g2_fill_2 FILLER_4_417 ();
 sg13g2_fill_2 FILLER_4_423 ();
 sg13g2_fill_1 FILLER_4_451 ();
 sg13g2_fill_2 FILLER_4_470 ();
 sg13g2_fill_1 FILLER_4_472 ();
 sg13g2_decap_4 FILLER_4_486 ();
 sg13g2_fill_1 FILLER_4_490 ();
 sg13g2_decap_4 FILLER_4_532 ();
 sg13g2_fill_1 FILLER_4_536 ();
 sg13g2_fill_2 FILLER_4_541 ();
 sg13g2_fill_1 FILLER_4_543 ();
 sg13g2_decap_4 FILLER_4_572 ();
 sg13g2_fill_1 FILLER_4_576 ();
 sg13g2_decap_4 FILLER_4_594 ();
 sg13g2_fill_1 FILLER_4_598 ();
 sg13g2_fill_1 FILLER_4_693 ();
 sg13g2_fill_2 FILLER_4_707 ();
 sg13g2_fill_1 FILLER_4_709 ();
 sg13g2_fill_2 FILLER_4_738 ();
 sg13g2_fill_2 FILLER_4_754 ();
 sg13g2_fill_2 FILLER_4_820 ();
 sg13g2_fill_2 FILLER_4_855 ();
 sg13g2_fill_1 FILLER_4_857 ();
 sg13g2_fill_1 FILLER_4_877 ();
 sg13g2_fill_2 FILLER_4_896 ();
 sg13g2_fill_1 FILLER_4_898 ();
 sg13g2_fill_1 FILLER_4_923 ();
 sg13g2_fill_1 FILLER_4_939 ();
 sg13g2_fill_1 FILLER_4_1016 ();
 sg13g2_fill_2 FILLER_4_1033 ();
 sg13g2_fill_1 FILLER_4_1035 ();
 sg13g2_decap_8 FILLER_4_1045 ();
 sg13g2_fill_2 FILLER_4_1052 ();
 sg13g2_fill_1 FILLER_4_1060 ();
 sg13g2_fill_2 FILLER_4_1066 ();
 sg13g2_fill_1 FILLER_4_1068 ();
 sg13g2_fill_1 FILLER_4_1089 ();
 sg13g2_fill_2 FILLER_4_1095 ();
 sg13g2_fill_1 FILLER_4_1097 ();
 sg13g2_decap_4 FILLER_4_1103 ();
 sg13g2_fill_1 FILLER_4_1107 ();
 sg13g2_fill_2 FILLER_4_1136 ();
 sg13g2_fill_1 FILLER_4_1252 ();
 sg13g2_decap_8 FILLER_4_1294 ();
 sg13g2_fill_1 FILLER_4_1301 ();
 sg13g2_fill_2 FILLER_4_1312 ();
 sg13g2_fill_2 FILLER_4_1366 ();
 sg13g2_fill_1 FILLER_4_1368 ();
 sg13g2_decap_4 FILLER_4_1373 ();
 sg13g2_fill_2 FILLER_4_1377 ();
 sg13g2_fill_2 FILLER_4_1415 ();
 sg13g2_fill_2 FILLER_4_1430 ();
 sg13g2_decap_4 FILLER_4_1437 ();
 sg13g2_fill_2 FILLER_4_1454 ();
 sg13g2_fill_2 FILLER_4_1470 ();
 sg13g2_decap_4 FILLER_4_1478 ();
 sg13g2_fill_1 FILLER_4_1482 ();
 sg13g2_fill_2 FILLER_4_1499 ();
 sg13g2_fill_2 FILLER_4_1544 ();
 sg13g2_fill_1 FILLER_4_1555 ();
 sg13g2_decap_8 FILLER_4_1566 ();
 sg13g2_decap_8 FILLER_4_1573 ();
 sg13g2_fill_1 FILLER_4_1580 ();
 sg13g2_fill_2 FILLER_4_1622 ();
 sg13g2_fill_1 FILLER_4_1624 ();
 sg13g2_decap_4 FILLER_4_1650 ();
 sg13g2_decap_8 FILLER_4_1659 ();
 sg13g2_decap_4 FILLER_4_1666 ();
 sg13g2_fill_2 FILLER_4_1670 ();
 sg13g2_decap_4 FILLER_4_1682 ();
 sg13g2_fill_1 FILLER_4_1694 ();
 sg13g2_fill_1 FILLER_4_1700 ();
 sg13g2_decap_4 FILLER_4_1729 ();
 sg13g2_fill_1 FILLER_4_1733 ();
 sg13g2_fill_2 FILLER_4_1737 ();
 sg13g2_fill_1 FILLER_4_1739 ();
 sg13g2_fill_1 FILLER_4_1753 ();
 sg13g2_fill_1 FILLER_4_1774 ();
 sg13g2_fill_2 FILLER_4_1780 ();
 sg13g2_fill_1 FILLER_4_1789 ();
 sg13g2_fill_2 FILLER_4_1799 ();
 sg13g2_decap_8 FILLER_4_1817 ();
 sg13g2_fill_1 FILLER_4_1824 ();
 sg13g2_fill_1 FILLER_4_1846 ();
 sg13g2_fill_2 FILLER_4_1855 ();
 sg13g2_fill_1 FILLER_4_1865 ();
 sg13g2_fill_2 FILLER_4_1878 ();
 sg13g2_fill_1 FILLER_4_1880 ();
 sg13g2_fill_2 FILLER_4_1895 ();
 sg13g2_fill_1 FILLER_4_1897 ();
 sg13g2_decap_8 FILLER_4_1908 ();
 sg13g2_fill_1 FILLER_4_1915 ();
 sg13g2_fill_2 FILLER_4_1936 ();
 sg13g2_decap_8 FILLER_4_1952 ();
 sg13g2_fill_1 FILLER_4_1959 ();
 sg13g2_fill_2 FILLER_4_1965 ();
 sg13g2_fill_1 FILLER_4_1967 ();
 sg13g2_fill_1 FILLER_4_1990 ();
 sg13g2_fill_2 FILLER_4_2000 ();
 sg13g2_fill_2 FILLER_4_2018 ();
 sg13g2_fill_2 FILLER_4_2029 ();
 sg13g2_fill_1 FILLER_4_2031 ();
 sg13g2_fill_1 FILLER_4_2040 ();
 sg13g2_decap_8 FILLER_4_2059 ();
 sg13g2_decap_4 FILLER_4_2076 ();
 sg13g2_fill_2 FILLER_4_2080 ();
 sg13g2_fill_1 FILLER_4_2092 ();
 sg13g2_decap_4 FILLER_4_2107 ();
 sg13g2_decap_8 FILLER_4_2130 ();
 sg13g2_fill_2 FILLER_4_2137 ();
 sg13g2_fill_1 FILLER_4_2139 ();
 sg13g2_fill_2 FILLER_4_2156 ();
 sg13g2_fill_2 FILLER_4_2175 ();
 sg13g2_fill_1 FILLER_4_2177 ();
 sg13g2_fill_2 FILLER_4_2202 ();
 sg13g2_decap_4 FILLER_4_2243 ();
 sg13g2_fill_2 FILLER_4_2271 ();
 sg13g2_fill_1 FILLER_4_2273 ();
 sg13g2_fill_2 FILLER_4_2288 ();
 sg13g2_fill_1 FILLER_4_2290 ();
 sg13g2_decap_4 FILLER_4_2304 ();
 sg13g2_fill_2 FILLER_4_2313 ();
 sg13g2_fill_1 FILLER_4_2315 ();
 sg13g2_fill_1 FILLER_4_2356 ();
 sg13g2_fill_2 FILLER_4_2366 ();
 sg13g2_fill_1 FILLER_4_2389 ();
 sg13g2_decap_4 FILLER_4_2400 ();
 sg13g2_fill_1 FILLER_4_2404 ();
 sg13g2_fill_2 FILLER_4_2431 ();
 sg13g2_fill_1 FILLER_4_2433 ();
 sg13g2_fill_2 FILLER_4_2451 ();
 sg13g2_fill_2 FILLER_4_2485 ();
 sg13g2_fill_2 FILLER_4_2525 ();
 sg13g2_fill_1 FILLER_4_2527 ();
 sg13g2_decap_8 FILLER_4_2541 ();
 sg13g2_decap_8 FILLER_4_2548 ();
 sg13g2_fill_1 FILLER_4_2555 ();
 sg13g2_fill_2 FILLER_4_2573 ();
 sg13g2_fill_1 FILLER_4_2575 ();
 sg13g2_decap_8 FILLER_4_2595 ();
 sg13g2_fill_1 FILLER_4_2602 ();
 sg13g2_decap_4 FILLER_4_2628 ();
 sg13g2_fill_1 FILLER_4_2632 ();
 sg13g2_fill_1 FILLER_4_2649 ();
 sg13g2_decap_8 FILLER_4_2655 ();
 sg13g2_fill_2 FILLER_4_2672 ();
 sg13g2_fill_2 FILLER_4_2688 ();
 sg13g2_decap_4 FILLER_4_2711 ();
 sg13g2_fill_1 FILLER_4_2715 ();
 sg13g2_decap_8 FILLER_4_2728 ();
 sg13g2_fill_1 FILLER_4_2735 ();
 sg13g2_decap_4 FILLER_4_2759 ();
 sg13g2_fill_2 FILLER_4_2787 ();
 sg13g2_fill_1 FILLER_4_2789 ();
 sg13g2_fill_2 FILLER_4_2809 ();
 sg13g2_fill_1 FILLER_4_2811 ();
 sg13g2_decap_4 FILLER_4_2831 ();
 sg13g2_fill_1 FILLER_4_2844 ();
 sg13g2_fill_1 FILLER_4_2850 ();
 sg13g2_fill_2 FILLER_4_2860 ();
 sg13g2_decap_4 FILLER_4_2871 ();
 sg13g2_fill_1 FILLER_4_2912 ();
 sg13g2_fill_2 FILLER_4_2934 ();
 sg13g2_fill_1 FILLER_4_2936 ();
 sg13g2_fill_1 FILLER_4_2956 ();
 sg13g2_decap_4 FILLER_4_2962 ();
 sg13g2_fill_2 FILLER_4_2974 ();
 sg13g2_fill_1 FILLER_4_2976 ();
 sg13g2_fill_1 FILLER_4_3001 ();
 sg13g2_decap_4 FILLER_4_3006 ();
 sg13g2_fill_2 FILLER_4_3027 ();
 sg13g2_fill_2 FILLER_4_3042 ();
 sg13g2_fill_1 FILLER_4_3044 ();
 sg13g2_fill_1 FILLER_4_3091 ();
 sg13g2_fill_1 FILLER_4_3105 ();
 sg13g2_fill_2 FILLER_4_3119 ();
 sg13g2_fill_2 FILLER_4_3152 ();
 sg13g2_decap_4 FILLER_4_3164 ();
 sg13g2_fill_2 FILLER_4_3168 ();
 sg13g2_fill_1 FILLER_4_3181 ();
 sg13g2_fill_1 FILLER_4_3187 ();
 sg13g2_fill_2 FILLER_4_3192 ();
 sg13g2_fill_2 FILLER_4_3220 ();
 sg13g2_fill_2 FILLER_4_3230 ();
 sg13g2_fill_2 FILLER_4_3284 ();
 sg13g2_fill_2 FILLER_4_3326 ();
 sg13g2_decap_4 FILLER_4_3332 ();
 sg13g2_fill_2 FILLER_4_3336 ();
 sg13g2_decap_4 FILLER_4_3420 ();
 sg13g2_fill_2 FILLER_4_3424 ();
 sg13g2_fill_2 FILLER_4_3483 ();
 sg13g2_fill_1 FILLER_4_3532 ();
 sg13g2_decap_4 FILLER_4_3552 ();
 sg13g2_fill_2 FILLER_4_3556 ();
 sg13g2_decap_8 FILLER_4_3562 ();
 sg13g2_decap_8 FILLER_4_3569 ();
 sg13g2_decap_4 FILLER_4_3576 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_18 ();
 sg13g2_fill_1 FILLER_5_25 ();
 sg13g2_fill_2 FILLER_5_43 ();
 sg13g2_fill_1 FILLER_5_58 ();
 sg13g2_fill_1 FILLER_5_76 ();
 sg13g2_fill_2 FILLER_5_97 ();
 sg13g2_fill_1 FILLER_5_99 ();
 sg13g2_fill_2 FILLER_5_109 ();
 sg13g2_fill_1 FILLER_5_111 ();
 sg13g2_fill_1 FILLER_5_130 ();
 sg13g2_decap_4 FILLER_5_144 ();
 sg13g2_fill_2 FILLER_5_167 ();
 sg13g2_decap_4 FILLER_5_179 ();
 sg13g2_fill_2 FILLER_5_188 ();
 sg13g2_fill_2 FILLER_5_219 ();
 sg13g2_fill_1 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_256 ();
 sg13g2_decap_8 FILLER_5_263 ();
 sg13g2_fill_2 FILLER_5_270 ();
 sg13g2_fill_1 FILLER_5_280 ();
 sg13g2_fill_2 FILLER_5_294 ();
 sg13g2_fill_1 FILLER_5_305 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_fill_2 FILLER_5_335 ();
 sg13g2_fill_1 FILLER_5_352 ();
 sg13g2_fill_1 FILLER_5_360 ();
 sg13g2_fill_2 FILLER_5_366 ();
 sg13g2_fill_2 FILLER_5_381 ();
 sg13g2_fill_1 FILLER_5_383 ();
 sg13g2_fill_1 FILLER_5_388 ();
 sg13g2_decap_8 FILLER_5_403 ();
 sg13g2_decap_4 FILLER_5_410 ();
 sg13g2_fill_1 FILLER_5_418 ();
 sg13g2_fill_1 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_451 ();
 sg13g2_fill_1 FILLER_5_458 ();
 sg13g2_fill_2 FILLER_5_495 ();
 sg13g2_fill_1 FILLER_5_497 ();
 sg13g2_fill_1 FILLER_5_526 ();
 sg13g2_decap_4 FILLER_5_535 ();
 sg13g2_fill_1 FILLER_5_539 ();
 sg13g2_decap_4 FILLER_5_562 ();
 sg13g2_decap_4 FILLER_5_569 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_4 FILLER_5_595 ();
 sg13g2_fill_1 FILLER_5_599 ();
 sg13g2_fill_2 FILLER_5_628 ();
 sg13g2_fill_1 FILLER_5_630 ();
 sg13g2_fill_2 FILLER_5_657 ();
 sg13g2_fill_1 FILLER_5_695 ();
 sg13g2_fill_2 FILLER_5_705 ();
 sg13g2_fill_2 FILLER_5_717 ();
 sg13g2_fill_2 FILLER_5_732 ();
 sg13g2_fill_1 FILLER_5_766 ();
 sg13g2_fill_2 FILLER_5_848 ();
 sg13g2_fill_2 FILLER_5_895 ();
 sg13g2_fill_1 FILLER_5_897 ();
 sg13g2_decap_4 FILLER_5_920 ();
 sg13g2_fill_1 FILLER_5_955 ();
 sg13g2_fill_2 FILLER_5_1008 ();
 sg13g2_decap_8 FILLER_5_1015 ();
 sg13g2_decap_8 FILLER_5_1027 ();
 sg13g2_decap_8 FILLER_5_1034 ();
 sg13g2_decap_4 FILLER_5_1041 ();
 sg13g2_fill_1 FILLER_5_1045 ();
 sg13g2_fill_2 FILLER_5_1102 ();
 sg13g2_fill_1 FILLER_5_1104 ();
 sg13g2_decap_4 FILLER_5_1119 ();
 sg13g2_fill_1 FILLER_5_1123 ();
 sg13g2_fill_2 FILLER_5_1137 ();
 sg13g2_fill_1 FILLER_5_1139 ();
 sg13g2_fill_1 FILLER_5_1145 ();
 sg13g2_fill_2 FILLER_5_1154 ();
 sg13g2_fill_1 FILLER_5_1156 ();
 sg13g2_fill_2 FILLER_5_1166 ();
 sg13g2_fill_1 FILLER_5_1168 ();
 sg13g2_decap_8 FILLER_5_1195 ();
 sg13g2_decap_8 FILLER_5_1202 ();
 sg13g2_decap_4 FILLER_5_1209 ();
 sg13g2_decap_4 FILLER_5_1222 ();
 sg13g2_fill_2 FILLER_5_1226 ();
 sg13g2_fill_2 FILLER_5_1277 ();
 sg13g2_fill_1 FILLER_5_1279 ();
 sg13g2_fill_1 FILLER_5_1383 ();
 sg13g2_fill_2 FILLER_5_1397 ();
 sg13g2_fill_1 FILLER_5_1399 ();
 sg13g2_fill_1 FILLER_5_1405 ();
 sg13g2_fill_2 FILLER_5_1416 ();
 sg13g2_fill_1 FILLER_5_1418 ();
 sg13g2_decap_8 FILLER_5_1439 ();
 sg13g2_fill_2 FILLER_5_1446 ();
 sg13g2_decap_4 FILLER_5_1456 ();
 sg13g2_fill_2 FILLER_5_1495 ();
 sg13g2_fill_1 FILLER_5_1497 ();
 sg13g2_decap_8 FILLER_5_1509 ();
 sg13g2_fill_2 FILLER_5_1516 ();
 sg13g2_fill_2 FILLER_5_1550 ();
 sg13g2_decap_8 FILLER_5_1632 ();
 sg13g2_decap_4 FILLER_5_1662 ();
 sg13g2_fill_2 FILLER_5_1666 ();
 sg13g2_fill_1 FILLER_5_1694 ();
 sg13g2_fill_2 FILLER_5_1700 ();
 sg13g2_fill_1 FILLER_5_1702 ();
 sg13g2_decap_4 FILLER_5_1724 ();
 sg13g2_fill_1 FILLER_5_1746 ();
 sg13g2_fill_1 FILLER_5_1759 ();
 sg13g2_fill_1 FILLER_5_1765 ();
 sg13g2_fill_1 FILLER_5_1771 ();
 sg13g2_decap_8 FILLER_5_1778 ();
 sg13g2_fill_1 FILLER_5_1785 ();
 sg13g2_fill_2 FILLER_5_1791 ();
 sg13g2_fill_2 FILLER_5_1797 ();
 sg13g2_fill_2 FILLER_5_1811 ();
 sg13g2_fill_1 FILLER_5_1813 ();
 sg13g2_decap_8 FILLER_5_1822 ();
 sg13g2_decap_4 FILLER_5_1829 ();
 sg13g2_fill_2 FILLER_5_1837 ();
 sg13g2_fill_2 FILLER_5_1858 ();
 sg13g2_fill_1 FILLER_5_1860 ();
 sg13g2_fill_2 FILLER_5_1876 ();
 sg13g2_fill_1 FILLER_5_1878 ();
 sg13g2_fill_2 FILLER_5_1892 ();
 sg13g2_decap_8 FILLER_5_1916 ();
 sg13g2_fill_2 FILLER_5_1923 ();
 sg13g2_fill_1 FILLER_5_1925 ();
 sg13g2_fill_1 FILLER_5_1931 ();
 sg13g2_fill_2 FILLER_5_1940 ();
 sg13g2_fill_2 FILLER_5_1950 ();
 sg13g2_fill_2 FILLER_5_1980 ();
 sg13g2_fill_1 FILLER_5_1991 ();
 sg13g2_fill_1 FILLER_5_2004 ();
 sg13g2_fill_2 FILLER_5_2010 ();
 sg13g2_fill_1 FILLER_5_2033 ();
 sg13g2_fill_1 FILLER_5_2052 ();
 sg13g2_fill_1 FILLER_5_2063 ();
 sg13g2_fill_2 FILLER_5_2080 ();
 sg13g2_decap_4 FILLER_5_2105 ();
 sg13g2_fill_2 FILLER_5_2109 ();
 sg13g2_fill_1 FILLER_5_2135 ();
 sg13g2_fill_2 FILLER_5_2144 ();
 sg13g2_fill_1 FILLER_5_2146 ();
 sg13g2_fill_2 FILLER_5_2160 ();
 sg13g2_decap_4 FILLER_5_2166 ();
 sg13g2_fill_1 FILLER_5_2170 ();
 sg13g2_fill_2 FILLER_5_2188 ();
 sg13g2_decap_8 FILLER_5_2214 ();
 sg13g2_decap_4 FILLER_5_2221 ();
 sg13g2_decap_8 FILLER_5_2239 ();
 sg13g2_decap_8 FILLER_5_2246 ();
 sg13g2_fill_1 FILLER_5_2253 ();
 sg13g2_decap_8 FILLER_5_2259 ();
 sg13g2_decap_8 FILLER_5_2266 ();
 sg13g2_decap_8 FILLER_5_2273 ();
 sg13g2_fill_2 FILLER_5_2280 ();
 sg13g2_fill_1 FILLER_5_2336 ();
 sg13g2_fill_2 FILLER_5_2352 ();
 sg13g2_fill_1 FILLER_5_2354 ();
 sg13g2_decap_8 FILLER_5_2380 ();
 sg13g2_fill_1 FILLER_5_2387 ();
 sg13g2_fill_1 FILLER_5_2419 ();
 sg13g2_fill_1 FILLER_5_2435 ();
 sg13g2_decap_4 FILLER_5_2440 ();
 sg13g2_fill_2 FILLER_5_2444 ();
 sg13g2_fill_1 FILLER_5_2506 ();
 sg13g2_fill_2 FILLER_5_2522 ();
 sg13g2_fill_1 FILLER_5_2541 ();
 sg13g2_fill_1 FILLER_5_2570 ();
 sg13g2_decap_4 FILLER_5_2597 ();
 sg13g2_fill_2 FILLER_5_2601 ();
 sg13g2_fill_1 FILLER_5_2631 ();
 sg13g2_decap_8 FILLER_5_2652 ();
 sg13g2_decap_4 FILLER_5_2659 ();
 sg13g2_fill_2 FILLER_5_2676 ();
 sg13g2_fill_1 FILLER_5_2678 ();
 sg13g2_fill_2 FILLER_5_2692 ();
 sg13g2_fill_1 FILLER_5_2719 ();
 sg13g2_fill_1 FILLER_5_2724 ();
 sg13g2_fill_2 FILLER_5_2757 ();
 sg13g2_fill_1 FILLER_5_2759 ();
 sg13g2_decap_4 FILLER_5_2770 ();
 sg13g2_decap_4 FILLER_5_2789 ();
 sg13g2_fill_1 FILLER_5_2793 ();
 sg13g2_fill_2 FILLER_5_2822 ();
 sg13g2_fill_2 FILLER_5_2834 ();
 sg13g2_fill_1 FILLER_5_2836 ();
 sg13g2_fill_1 FILLER_5_2853 ();
 sg13g2_fill_1 FILLER_5_2859 ();
 sg13g2_decap_8 FILLER_5_2873 ();
 sg13g2_fill_2 FILLER_5_2904 ();
 sg13g2_fill_2 FILLER_5_2919 ();
 sg13g2_fill_1 FILLER_5_2921 ();
 sg13g2_fill_2 FILLER_5_2934 ();
 sg13g2_fill_1 FILLER_5_2936 ();
 sg13g2_fill_2 FILLER_5_2960 ();
 sg13g2_decap_4 FILLER_5_2977 ();
 sg13g2_decap_8 FILLER_5_3000 ();
 sg13g2_fill_2 FILLER_5_3007 ();
 sg13g2_fill_1 FILLER_5_3032 ();
 sg13g2_fill_2 FILLER_5_3038 ();
 sg13g2_decap_4 FILLER_5_3053 ();
 sg13g2_fill_1 FILLER_5_3057 ();
 sg13g2_fill_2 FILLER_5_3080 ();
 sg13g2_fill_2 FILLER_5_3103 ();
 sg13g2_fill_1 FILLER_5_3105 ();
 sg13g2_fill_2 FILLER_5_3124 ();
 sg13g2_fill_1 FILLER_5_3126 ();
 sg13g2_fill_1 FILLER_5_3141 ();
 sg13g2_fill_2 FILLER_5_3146 ();
 sg13g2_fill_1 FILLER_5_3178 ();
 sg13g2_fill_1 FILLER_5_3184 ();
 sg13g2_fill_1 FILLER_5_3227 ();
 sg13g2_fill_1 FILLER_5_3232 ();
 sg13g2_decap_8 FILLER_5_3243 ();
 sg13g2_decap_4 FILLER_5_3250 ();
 sg13g2_fill_2 FILLER_5_3254 ();
 sg13g2_fill_2 FILLER_5_3272 ();
 sg13g2_fill_1 FILLER_5_3274 ();
 sg13g2_fill_2 FILLER_5_3283 ();
 sg13g2_fill_1 FILLER_5_3322 ();
 sg13g2_decap_4 FILLER_5_3332 ();
 sg13g2_fill_1 FILLER_5_3336 ();
 sg13g2_fill_1 FILLER_5_3340 ();
 sg13g2_fill_2 FILLER_5_3349 ();
 sg13g2_decap_4 FILLER_5_3360 ();
 sg13g2_fill_2 FILLER_5_3364 ();
 sg13g2_fill_2 FILLER_5_3375 ();
 sg13g2_fill_1 FILLER_5_3384 ();
 sg13g2_fill_2 FILLER_5_3390 ();
 sg13g2_fill_2 FILLER_5_3397 ();
 sg13g2_fill_2 FILLER_5_3408 ();
 sg13g2_fill_1 FILLER_5_3410 ();
 sg13g2_decap_8 FILLER_5_3437 ();
 sg13g2_decap_4 FILLER_5_3444 ();
 sg13g2_fill_2 FILLER_5_3448 ();
 sg13g2_fill_1 FILLER_5_3474 ();
 sg13g2_decap_4 FILLER_5_3488 ();
 sg13g2_fill_1 FILLER_5_3492 ();
 sg13g2_fill_1 FILLER_5_3526 ();
 sg13g2_fill_2 FILLER_5_3545 ();
 sg13g2_fill_1 FILLER_5_3547 ();
 sg13g2_decap_8 FILLER_5_3571 ();
 sg13g2_fill_2 FILLER_5_3578 ();
 sg13g2_decap_4 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_4 ();
 sg13g2_fill_2 FILLER_6_34 ();
 sg13g2_fill_1 FILLER_6_52 ();
 sg13g2_fill_2 FILLER_6_75 ();
 sg13g2_fill_2 FILLER_6_90 ();
 sg13g2_fill_1 FILLER_6_102 ();
 sg13g2_fill_1 FILLER_6_124 ();
 sg13g2_fill_2 FILLER_6_134 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_4 FILLER_6_147 ();
 sg13g2_fill_1 FILLER_6_151 ();
 sg13g2_fill_2 FILLER_6_162 ();
 sg13g2_fill_2 FILLER_6_213 ();
 sg13g2_fill_1 FILLER_6_215 ();
 sg13g2_fill_1 FILLER_6_228 ();
 sg13g2_fill_2 FILLER_6_239 ();
 sg13g2_fill_2 FILLER_6_244 ();
 sg13g2_fill_2 FILLER_6_250 ();
 sg13g2_fill_2 FILLER_6_263 ();
 sg13g2_fill_1 FILLER_6_265 ();
 sg13g2_decap_4 FILLER_6_285 ();
 sg13g2_fill_2 FILLER_6_289 ();
 sg13g2_decap_8 FILLER_6_360 ();
 sg13g2_decap_4 FILLER_6_375 ();
 sg13g2_fill_1 FILLER_6_379 ();
 sg13g2_fill_1 FILLER_6_393 ();
 sg13g2_decap_4 FILLER_6_407 ();
 sg13g2_fill_2 FILLER_6_411 ();
 sg13g2_decap_4 FILLER_6_426 ();
 sg13g2_fill_2 FILLER_6_430 ();
 sg13g2_fill_1 FILLER_6_443 ();
 sg13g2_fill_1 FILLER_6_474 ();
 sg13g2_fill_2 FILLER_6_484 ();
 sg13g2_fill_1 FILLER_6_486 ();
 sg13g2_fill_1 FILLER_6_495 ();
 sg13g2_decap_4 FILLER_6_500 ();
 sg13g2_fill_1 FILLER_6_507 ();
 sg13g2_fill_1 FILLER_6_528 ();
 sg13g2_fill_2 FILLER_6_548 ();
 sg13g2_fill_1 FILLER_6_550 ();
 sg13g2_fill_2 FILLER_6_568 ();
 sg13g2_fill_1 FILLER_6_570 ();
 sg13g2_decap_4 FILLER_6_610 ();
 sg13g2_fill_1 FILLER_6_637 ();
 sg13g2_fill_2 FILLER_6_679 ();
 sg13g2_fill_1 FILLER_6_681 ();
 sg13g2_decap_4 FILLER_6_694 ();
 sg13g2_fill_2 FILLER_6_698 ();
 sg13g2_decap_4 FILLER_6_724 ();
 sg13g2_fill_1 FILLER_6_728 ();
 sg13g2_fill_2 FILLER_6_742 ();
 sg13g2_fill_1 FILLER_6_744 ();
 sg13g2_fill_2 FILLER_6_824 ();
 sg13g2_decap_8 FILLER_6_839 ();
 sg13g2_decap_8 FILLER_6_864 ();
 sg13g2_decap_8 FILLER_6_871 ();
 sg13g2_fill_2 FILLER_6_878 ();
 sg13g2_fill_1 FILLER_6_880 ();
 sg13g2_fill_2 FILLER_6_906 ();
 sg13g2_decap_8 FILLER_6_912 ();
 sg13g2_fill_2 FILLER_6_919 ();
 sg13g2_fill_1 FILLER_6_921 ();
 sg13g2_fill_2 FILLER_6_974 ();
 sg13g2_fill_1 FILLER_6_976 ();
 sg13g2_fill_2 FILLER_6_982 ();
 sg13g2_fill_1 FILLER_6_984 ();
 sg13g2_fill_2 FILLER_6_1035 ();
 sg13g2_fill_2 FILLER_6_1065 ();
 sg13g2_decap_4 FILLER_6_1168 ();
 sg13g2_decap_4 FILLER_6_1175 ();
 sg13g2_fill_1 FILLER_6_1179 ();
 sg13g2_fill_1 FILLER_6_1184 ();
 sg13g2_fill_2 FILLER_6_1190 ();
 sg13g2_fill_1 FILLER_6_1192 ();
 sg13g2_fill_2 FILLER_6_1289 ();
 sg13g2_decap_4 FILLER_6_1313 ();
 sg13g2_fill_1 FILLER_6_1317 ();
 sg13g2_fill_2 FILLER_6_1377 ();
 sg13g2_fill_2 FILLER_6_1392 ();
 sg13g2_decap_4 FILLER_6_1419 ();
 sg13g2_fill_2 FILLER_6_1423 ();
 sg13g2_decap_8 FILLER_6_1433 ();
 sg13g2_fill_2 FILLER_6_1440 ();
 sg13g2_fill_1 FILLER_6_1442 ();
 sg13g2_decap_8 FILLER_6_1467 ();
 sg13g2_fill_2 FILLER_6_1505 ();
 sg13g2_fill_2 FILLER_6_1515 ();
 sg13g2_decap_4 FILLER_6_1527 ();
 sg13g2_fill_2 FILLER_6_1536 ();
 sg13g2_fill_1 FILLER_6_1538 ();
 sg13g2_fill_2 FILLER_6_1553 ();
 sg13g2_fill_1 FILLER_6_1568 ();
 sg13g2_decap_8 FILLER_6_1578 ();
 sg13g2_fill_2 FILLER_6_1589 ();
 sg13g2_fill_1 FILLER_6_1591 ();
 sg13g2_decap_8 FILLER_6_1612 ();
 sg13g2_decap_4 FILLER_6_1619 ();
 sg13g2_fill_1 FILLER_6_1623 ();
 sg13g2_fill_2 FILLER_6_1637 ();
 sg13g2_fill_2 FILLER_6_1649 ();
 sg13g2_decap_8 FILLER_6_1659 ();
 sg13g2_decap_8 FILLER_6_1666 ();
 sg13g2_decap_4 FILLER_6_1673 ();
 sg13g2_decap_4 FILLER_6_1687 ();
 sg13g2_fill_2 FILLER_6_1691 ();
 sg13g2_fill_2 FILLER_6_1722 ();
 sg13g2_fill_1 FILLER_6_1724 ();
 sg13g2_fill_2 FILLER_6_1765 ();
 sg13g2_fill_1 FILLER_6_1767 ();
 sg13g2_fill_2 FILLER_6_1773 ();
 sg13g2_fill_2 FILLER_6_1795 ();
 sg13g2_fill_1 FILLER_6_1817 ();
 sg13g2_decap_8 FILLER_6_1828 ();
 sg13g2_decap_4 FILLER_6_1835 ();
 sg13g2_fill_1 FILLER_6_1839 ();
 sg13g2_fill_2 FILLER_6_1868 ();
 sg13g2_fill_1 FILLER_6_1870 ();
 sg13g2_fill_2 FILLER_6_1876 ();
 sg13g2_fill_2 FILLER_6_1888 ();
 sg13g2_fill_1 FILLER_6_1890 ();
 sg13g2_fill_2 FILLER_6_1904 ();
 sg13g2_fill_1 FILLER_6_1906 ();
 sg13g2_fill_1 FILLER_6_1916 ();
 sg13g2_decap_8 FILLER_6_1936 ();
 sg13g2_fill_1 FILLER_6_1961 ();
 sg13g2_fill_1 FILLER_6_1980 ();
 sg13g2_fill_1 FILLER_6_1990 ();
 sg13g2_fill_1 FILLER_6_2013 ();
 sg13g2_fill_1 FILLER_6_2019 ();
 sg13g2_fill_2 FILLER_6_2030 ();
 sg13g2_fill_1 FILLER_6_2032 ();
 sg13g2_fill_1 FILLER_6_2064 ();
 sg13g2_fill_2 FILLER_6_2081 ();
 sg13g2_fill_1 FILLER_6_2095 ();
 sg13g2_fill_1 FILLER_6_2106 ();
 sg13g2_fill_2 FILLER_6_2189 ();
 sg13g2_fill_1 FILLER_6_2191 ();
 sg13g2_fill_2 FILLER_6_2208 ();
 sg13g2_fill_1 FILLER_6_2210 ();
 sg13g2_decap_4 FILLER_6_2216 ();
 sg13g2_decap_4 FILLER_6_2244 ();
 sg13g2_fill_1 FILLER_6_2248 ();
 sg13g2_decap_8 FILLER_6_2286 ();
 sg13g2_fill_2 FILLER_6_2293 ();
 sg13g2_fill_2 FILLER_6_2340 ();
 sg13g2_fill_1 FILLER_6_2348 ();
 sg13g2_fill_2 FILLER_6_2363 ();
 sg13g2_decap_4 FILLER_6_2379 ();
 sg13g2_fill_2 FILLER_6_2383 ();
 sg13g2_fill_2 FILLER_6_2413 ();
 sg13g2_fill_1 FILLER_6_2415 ();
 sg13g2_fill_2 FILLER_6_2439 ();
 sg13g2_fill_2 FILLER_6_2497 ();
 sg13g2_fill_2 FILLER_6_2520 ();
 sg13g2_fill_1 FILLER_6_2522 ();
 sg13g2_fill_1 FILLER_6_2528 ();
 sg13g2_fill_2 FILLER_6_2533 ();
 sg13g2_decap_4 FILLER_6_2543 ();
 sg13g2_decap_8 FILLER_6_2555 ();
 sg13g2_fill_1 FILLER_6_2590 ();
 sg13g2_fill_1 FILLER_6_2609 ();
 sg13g2_fill_2 FILLER_6_2615 ();
 sg13g2_decap_4 FILLER_6_2654 ();
 sg13g2_fill_2 FILLER_6_2658 ();
 sg13g2_decap_4 FILLER_6_2680 ();
 sg13g2_fill_2 FILLER_6_2684 ();
 sg13g2_decap_4 FILLER_6_2699 ();
 sg13g2_decap_4 FILLER_6_2720 ();
 sg13g2_decap_4 FILLER_6_2734 ();
 sg13g2_decap_4 FILLER_6_2757 ();
 sg13g2_fill_2 FILLER_6_2776 ();
 sg13g2_decap_8 FILLER_6_2790 ();
 sg13g2_decap_8 FILLER_6_2797 ();
 sg13g2_fill_2 FILLER_6_2804 ();
 sg13g2_fill_1 FILLER_6_2806 ();
 sg13g2_decap_8 FILLER_6_2815 ();
 sg13g2_fill_2 FILLER_6_2832 ();
 sg13g2_decap_4 FILLER_6_2874 ();
 sg13g2_fill_1 FILLER_6_2878 ();
 sg13g2_decap_4 FILLER_6_2923 ();
 sg13g2_decap_4 FILLER_6_2932 ();
 sg13g2_fill_1 FILLER_6_2967 ();
 sg13g2_fill_1 FILLER_6_2978 ();
 sg13g2_decap_4 FILLER_6_2996 ();
 sg13g2_decap_4 FILLER_6_3013 ();
 sg13g2_fill_1 FILLER_6_3017 ();
 sg13g2_fill_2 FILLER_6_3042 ();
 sg13g2_fill_1 FILLER_6_3044 ();
 sg13g2_fill_2 FILLER_6_3050 ();
 sg13g2_fill_1 FILLER_6_3052 ();
 sg13g2_decap_8 FILLER_6_3074 ();
 sg13g2_fill_2 FILLER_6_3081 ();
 sg13g2_fill_1 FILLER_6_3083 ();
 sg13g2_fill_2 FILLER_6_3102 ();
 sg13g2_fill_1 FILLER_6_3104 ();
 sg13g2_fill_2 FILLER_6_3154 ();
 sg13g2_decap_4 FILLER_6_3192 ();
 sg13g2_fill_2 FILLER_6_3196 ();
 sg13g2_decap_4 FILLER_6_3206 ();
 sg13g2_fill_2 FILLER_6_3210 ();
 sg13g2_fill_2 FILLER_6_3216 ();
 sg13g2_fill_1 FILLER_6_3218 ();
 sg13g2_decap_4 FILLER_6_3222 ();
 sg13g2_decap_4 FILLER_6_3243 ();
 sg13g2_fill_1 FILLER_6_3247 ();
 sg13g2_decap_4 FILLER_6_3251 ();
 sg13g2_fill_1 FILLER_6_3255 ();
 sg13g2_fill_1 FILLER_6_3260 ();
 sg13g2_fill_2 FILLER_6_3276 ();
 sg13g2_fill_2 FILLER_6_3285 ();
 sg13g2_fill_2 FILLER_6_3334 ();
 sg13g2_fill_2 FILLER_6_3357 ();
 sg13g2_fill_1 FILLER_6_3364 ();
 sg13g2_fill_1 FILLER_6_3375 ();
 sg13g2_fill_2 FILLER_6_3381 ();
 sg13g2_fill_2 FILLER_6_3409 ();
 sg13g2_fill_1 FILLER_6_3411 ();
 sg13g2_fill_1 FILLER_6_3420 ();
 sg13g2_fill_2 FILLER_6_3425 ();
 sg13g2_fill_1 FILLER_6_3427 ();
 sg13g2_fill_1 FILLER_6_3437 ();
 sg13g2_fill_2 FILLER_6_3441 ();
 sg13g2_fill_2 FILLER_6_3461 ();
 sg13g2_fill_1 FILLER_6_3463 ();
 sg13g2_fill_1 FILLER_6_3477 ();
 sg13g2_decap_4 FILLER_6_3495 ();
 sg13g2_fill_1 FILLER_6_3499 ();
 sg13g2_decap_8 FILLER_6_3523 ();
 sg13g2_fill_1 FILLER_6_3534 ();
 sg13g2_fill_2 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_2 ();
 sg13g2_fill_1 FILLER_7_10 ();
 sg13g2_decap_8 FILLER_7_15 ();
 sg13g2_decap_4 FILLER_7_22 ();
 sg13g2_fill_2 FILLER_7_26 ();
 sg13g2_fill_1 FILLER_7_45 ();
 sg13g2_fill_2 FILLER_7_54 ();
 sg13g2_fill_2 FILLER_7_90 ();
 sg13g2_fill_1 FILLER_7_102 ();
 sg13g2_fill_2 FILLER_7_171 ();
 sg13g2_fill_1 FILLER_7_173 ();
 sg13g2_fill_1 FILLER_7_179 ();
 sg13g2_fill_2 FILLER_7_184 ();
 sg13g2_decap_4 FILLER_7_232 ();
 sg13g2_fill_1 FILLER_7_266 ();
 sg13g2_fill_1 FILLER_7_304 ();
 sg13g2_fill_2 FILLER_7_320 ();
 sg13g2_fill_2 FILLER_7_350 ();
 sg13g2_fill_1 FILLER_7_364 ();
 sg13g2_decap_4 FILLER_7_368 ();
 sg13g2_fill_1 FILLER_7_372 ();
 sg13g2_fill_2 FILLER_7_386 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_439 ();
 sg13g2_decap_4 FILLER_7_448 ();
 sg13g2_fill_1 FILLER_7_452 ();
 sg13g2_fill_2 FILLER_7_462 ();
 sg13g2_fill_1 FILLER_7_473 ();
 sg13g2_fill_2 FILLER_7_499 ();
 sg13g2_fill_2 FILLER_7_509 ();
 sg13g2_fill_1 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_522 ();
 sg13g2_decap_8 FILLER_7_529 ();
 sg13g2_decap_4 FILLER_7_536 ();
 sg13g2_fill_2 FILLER_7_567 ();
 sg13g2_fill_1 FILLER_7_569 ();
 sg13g2_fill_1 FILLER_7_583 ();
 sg13g2_fill_2 FILLER_7_632 ();
 sg13g2_decap_8 FILLER_7_646 ();
 sg13g2_decap_4 FILLER_7_653 ();
 sg13g2_fill_1 FILLER_7_666 ();
 sg13g2_fill_2 FILLER_7_672 ();
 sg13g2_fill_2 FILLER_7_684 ();
 sg13g2_decap_4 FILLER_7_721 ();
 sg13g2_fill_1 FILLER_7_725 ();
 sg13g2_fill_2 FILLER_7_737 ();
 sg13g2_fill_1 FILLER_7_739 ();
 sg13g2_fill_2 FILLER_7_814 ();
 sg13g2_fill_1 FILLER_7_829 ();
 sg13g2_fill_2 FILLER_7_874 ();
 sg13g2_fill_1 FILLER_7_876 ();
 sg13g2_decap_8 FILLER_7_894 ();
 sg13g2_fill_1 FILLER_7_901 ();
 sg13g2_decap_4 FILLER_7_938 ();
 sg13g2_fill_1 FILLER_7_942 ();
 sg13g2_decap_4 FILLER_7_947 ();
 sg13g2_fill_2 FILLER_7_956 ();
 sg13g2_fill_1 FILLER_7_958 ();
 sg13g2_fill_1 FILLER_7_971 ();
 sg13g2_decap_8 FILLER_7_1021 ();
 sg13g2_decap_8 FILLER_7_1028 ();
 sg13g2_fill_2 FILLER_7_1035 ();
 sg13g2_fill_2 FILLER_7_1058 ();
 sg13g2_decap_8 FILLER_7_1111 ();
 sg13g2_decap_8 FILLER_7_1118 ();
 sg13g2_decap_8 FILLER_7_1125 ();
 sg13g2_fill_2 FILLER_7_1132 ();
 sg13g2_fill_1 FILLER_7_1134 ();
 sg13g2_fill_2 FILLER_7_1147 ();
 sg13g2_fill_1 FILLER_7_1149 ();
 sg13g2_fill_2 FILLER_7_1155 ();
 sg13g2_fill_1 FILLER_7_1157 ();
 sg13g2_fill_1 FILLER_7_1174 ();
 sg13g2_fill_2 FILLER_7_1181 ();
 sg13g2_fill_1 FILLER_7_1183 ();
 sg13g2_fill_1 FILLER_7_1197 ();
 sg13g2_decap_4 FILLER_7_1202 ();
 sg13g2_decap_8 FILLER_7_1211 ();
 sg13g2_fill_2 FILLER_7_1257 ();
 sg13g2_fill_2 FILLER_7_1272 ();
 sg13g2_fill_1 FILLER_7_1274 ();
 sg13g2_fill_1 FILLER_7_1284 ();
 sg13g2_fill_2 FILLER_7_1298 ();
 sg13g2_fill_1 FILLER_7_1322 ();
 sg13g2_decap_8 FILLER_7_1378 ();
 sg13g2_fill_1 FILLER_7_1385 ();
 sg13g2_fill_1 FILLER_7_1397 ();
 sg13g2_decap_8 FILLER_7_1421 ();
 sg13g2_decap_4 FILLER_7_1428 ();
 sg13g2_decap_4 FILLER_7_1453 ();
 sg13g2_fill_2 FILLER_7_1457 ();
 sg13g2_fill_2 FILLER_7_1466 ();
 sg13g2_decap_4 FILLER_7_1476 ();
 sg13g2_fill_1 FILLER_7_1480 ();
 sg13g2_decap_4 FILLER_7_1487 ();
 sg13g2_fill_2 FILLER_7_1491 ();
 sg13g2_fill_2 FILLER_7_1502 ();
 sg13g2_fill_2 FILLER_7_1514 ();
 sg13g2_fill_2 FILLER_7_1538 ();
 sg13g2_decap_4 FILLER_7_1585 ();
 sg13g2_fill_1 FILLER_7_1589 ();
 sg13g2_decap_4 FILLER_7_1662 ();
 sg13g2_fill_1 FILLER_7_1666 ();
 sg13g2_fill_2 FILLER_7_1671 ();
 sg13g2_fill_1 FILLER_7_1706 ();
 sg13g2_decap_8 FILLER_7_1717 ();
 sg13g2_fill_2 FILLER_7_1724 ();
 sg13g2_decap_8 FILLER_7_1744 ();
 sg13g2_decap_4 FILLER_7_1751 ();
 sg13g2_fill_2 FILLER_7_1755 ();
 sg13g2_decap_8 FILLER_7_1772 ();
 sg13g2_fill_1 FILLER_7_1785 ();
 sg13g2_fill_1 FILLER_7_1795 ();
 sg13g2_fill_1 FILLER_7_1811 ();
 sg13g2_decap_8 FILLER_7_1830 ();
 sg13g2_decap_8 FILLER_7_1857 ();
 sg13g2_decap_4 FILLER_7_1898 ();
 sg13g2_fill_1 FILLER_7_1919 ();
 sg13g2_decap_8 FILLER_7_1940 ();
 sg13g2_fill_1 FILLER_7_1975 ();
 sg13g2_fill_1 FILLER_7_1984 ();
 sg13g2_fill_2 FILLER_7_1995 ();
 sg13g2_decap_8 FILLER_7_2028 ();
 sg13g2_decap_8 FILLER_7_2035 ();
 sg13g2_fill_2 FILLER_7_2042 ();
 sg13g2_fill_1 FILLER_7_2044 ();
 sg13g2_decap_8 FILLER_7_2049 ();
 sg13g2_decap_8 FILLER_7_2056 ();
 sg13g2_decap_4 FILLER_7_2063 ();
 sg13g2_fill_2 FILLER_7_2067 ();
 sg13g2_fill_2 FILLER_7_2082 ();
 sg13g2_fill_1 FILLER_7_2108 ();
 sg13g2_fill_1 FILLER_7_2123 ();
 sg13g2_fill_2 FILLER_7_2138 ();
 sg13g2_fill_1 FILLER_7_2140 ();
 sg13g2_fill_2 FILLER_7_2150 ();
 sg13g2_decap_4 FILLER_7_2175 ();
 sg13g2_fill_2 FILLER_7_2193 ();
 sg13g2_fill_1 FILLER_7_2195 ();
 sg13g2_fill_2 FILLER_7_2201 ();
 sg13g2_decap_8 FILLER_7_2216 ();
 sg13g2_fill_1 FILLER_7_2223 ();
 sg13g2_fill_2 FILLER_7_2233 ();
 sg13g2_fill_2 FILLER_7_2239 ();
 sg13g2_fill_1 FILLER_7_2241 ();
 sg13g2_fill_2 FILLER_7_2287 ();
 sg13g2_fill_1 FILLER_7_2289 ();
 sg13g2_fill_1 FILLER_7_2299 ();
 sg13g2_fill_1 FILLER_7_2319 ();
 sg13g2_fill_2 FILLER_7_2337 ();
 sg13g2_fill_1 FILLER_7_2339 ();
 sg13g2_fill_1 FILLER_7_2376 ();
 sg13g2_fill_1 FILLER_7_2471 ();
 sg13g2_fill_1 FILLER_7_2547 ();
 sg13g2_fill_2 FILLER_7_2606 ();
 sg13g2_fill_1 FILLER_7_2608 ();
 sg13g2_fill_2 FILLER_7_2625 ();
 sg13g2_fill_1 FILLER_7_2627 ();
 sg13g2_fill_2 FILLER_7_2637 ();
 sg13g2_decap_8 FILLER_7_2654 ();
 sg13g2_decap_8 FILLER_7_2661 ();
 sg13g2_decap_8 FILLER_7_2678 ();
 sg13g2_fill_1 FILLER_7_2685 ();
 sg13g2_fill_1 FILLER_7_2689 ();
 sg13g2_fill_2 FILLER_7_2718 ();
 sg13g2_decap_8 FILLER_7_2755 ();
 sg13g2_fill_1 FILLER_7_2762 ();
 sg13g2_fill_2 FILLER_7_2780 ();
 sg13g2_decap_4 FILLER_7_2804 ();
 sg13g2_fill_2 FILLER_7_2839 ();
 sg13g2_fill_1 FILLER_7_2850 ();
 sg13g2_fill_2 FILLER_7_2864 ();
 sg13g2_decap_4 FILLER_7_2881 ();
 sg13g2_fill_1 FILLER_7_2885 ();
 sg13g2_fill_1 FILLER_7_2909 ();
 sg13g2_decap_4 FILLER_7_2923 ();
 sg13g2_fill_2 FILLER_7_2927 ();
 sg13g2_fill_2 FILLER_7_2933 ();
 sg13g2_decap_8 FILLER_7_2945 ();
 sg13g2_decap_8 FILLER_7_2952 ();
 sg13g2_fill_2 FILLER_7_2959 ();
 sg13g2_fill_1 FILLER_7_2961 ();
 sg13g2_fill_2 FILLER_7_2966 ();
 sg13g2_decap_8 FILLER_7_2972 ();
 sg13g2_decap_8 FILLER_7_2979 ();
 sg13g2_fill_2 FILLER_7_2996 ();
 sg13g2_fill_1 FILLER_7_2998 ();
 sg13g2_fill_1 FILLER_7_3022 ();
 sg13g2_decap_4 FILLER_7_3028 ();
 sg13g2_fill_1 FILLER_7_3052 ();
 sg13g2_fill_2 FILLER_7_3065 ();
 sg13g2_decap_8 FILLER_7_3082 ();
 sg13g2_fill_2 FILLER_7_3102 ();
 sg13g2_fill_1 FILLER_7_3104 ();
 sg13g2_decap_4 FILLER_7_3110 ();
 sg13g2_fill_2 FILLER_7_3127 ();
 sg13g2_fill_1 FILLER_7_3149 ();
 sg13g2_fill_1 FILLER_7_3196 ();
 sg13g2_fill_1 FILLER_7_3207 ();
 sg13g2_fill_2 FILLER_7_3225 ();
 sg13g2_fill_1 FILLER_7_3227 ();
 sg13g2_decap_8 FILLER_7_3250 ();
 sg13g2_fill_2 FILLER_7_3257 ();
 sg13g2_fill_1 FILLER_7_3299 ();
 sg13g2_fill_2 FILLER_7_3305 ();
 sg13g2_fill_1 FILLER_7_3354 ();
 sg13g2_fill_1 FILLER_7_3365 ();
 sg13g2_fill_1 FILLER_7_3378 ();
 sg13g2_fill_2 FILLER_7_3401 ();
 sg13g2_fill_1 FILLER_7_3403 ();
 sg13g2_fill_2 FILLER_7_3428 ();
 sg13g2_fill_1 FILLER_7_3430 ();
 sg13g2_fill_1 FILLER_7_3445 ();
 sg13g2_fill_2 FILLER_7_3466 ();
 sg13g2_fill_1 FILLER_7_3481 ();
 sg13g2_decap_8 FILLER_7_3502 ();
 sg13g2_fill_1 FILLER_7_3509 ();
 sg13g2_fill_2 FILLER_7_3515 ();
 sg13g2_fill_2 FILLER_7_3522 ();
 sg13g2_fill_1 FILLER_7_3524 ();
 sg13g2_fill_2 FILLER_7_3530 ();
 sg13g2_decap_8 FILLER_7_3553 ();
 sg13g2_decap_8 FILLER_7_3560 ();
 sg13g2_decap_8 FILLER_7_3567 ();
 sg13g2_decap_4 FILLER_7_3574 ();
 sg13g2_fill_2 FILLER_7_3578 ();
 sg13g2_fill_1 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_52 ();
 sg13g2_fill_1 FILLER_8_59 ();
 sg13g2_fill_2 FILLER_8_79 ();
 sg13g2_fill_1 FILLER_8_81 ();
 sg13g2_fill_1 FILLER_8_92 ();
 sg13g2_decap_8 FILLER_8_188 ();
 sg13g2_fill_1 FILLER_8_195 ();
 sg13g2_decap_4 FILLER_8_200 ();
 sg13g2_fill_1 FILLER_8_204 ();
 sg13g2_fill_2 FILLER_8_242 ();
 sg13g2_decap_8 FILLER_8_260 ();
 sg13g2_fill_2 FILLER_8_267 ();
 sg13g2_decap_4 FILLER_8_311 ();
 sg13g2_fill_1 FILLER_8_315 ();
 sg13g2_fill_2 FILLER_8_329 ();
 sg13g2_fill_1 FILLER_8_331 ();
 sg13g2_decap_4 FILLER_8_340 ();
 sg13g2_fill_2 FILLER_8_354 ();
 sg13g2_decap_8 FILLER_8_373 ();
 sg13g2_fill_2 FILLER_8_392 ();
 sg13g2_fill_1 FILLER_8_394 ();
 sg13g2_decap_8 FILLER_8_403 ();
 sg13g2_decap_8 FILLER_8_410 ();
 sg13g2_fill_2 FILLER_8_417 ();
 sg13g2_fill_2 FILLER_8_432 ();
 sg13g2_decap_8 FILLER_8_438 ();
 sg13g2_fill_2 FILLER_8_445 ();
 sg13g2_fill_2 FILLER_8_457 ();
 sg13g2_fill_1 FILLER_8_459 ();
 sg13g2_decap_4 FILLER_8_481 ();
 sg13g2_fill_2 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_fill_1 FILLER_8_518 ();
 sg13g2_fill_1 FILLER_8_532 ();
 sg13g2_fill_1 FILLER_8_569 ();
 sg13g2_fill_2 FILLER_8_588 ();
 sg13g2_fill_1 FILLER_8_590 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_fill_2 FILLER_8_625 ();
 sg13g2_fill_1 FILLER_8_627 ();
 sg13g2_decap_8 FILLER_8_640 ();
 sg13g2_fill_2 FILLER_8_647 ();
 sg13g2_fill_1 FILLER_8_649 ();
 sg13g2_decap_8 FILLER_8_654 ();
 sg13g2_decap_8 FILLER_8_661 ();
 sg13g2_fill_1 FILLER_8_675 ();
 sg13g2_fill_2 FILLER_8_693 ();
 sg13g2_fill_2 FILLER_8_699 ();
 sg13g2_fill_1 FILLER_8_701 ();
 sg13g2_fill_1 FILLER_8_711 ();
 sg13g2_decap_4 FILLER_8_726 ();
 sg13g2_fill_1 FILLER_8_730 ();
 sg13g2_decap_4 FILLER_8_747 ();
 sg13g2_fill_2 FILLER_8_754 ();
 sg13g2_decap_4 FILLER_8_772 ();
 sg13g2_fill_2 FILLER_8_781 ();
 sg13g2_fill_2 FILLER_8_801 ();
 sg13g2_fill_2 FILLER_8_811 ();
 sg13g2_fill_1 FILLER_8_834 ();
 sg13g2_decap_4 FILLER_8_839 ();
 sg13g2_fill_2 FILLER_8_846 ();
 sg13g2_decap_8 FILLER_8_888 ();
 sg13g2_fill_2 FILLER_8_895 ();
 sg13g2_fill_1 FILLER_8_897 ();
 sg13g2_decap_8 FILLER_8_921 ();
 sg13g2_decap_8 FILLER_8_937 ();
 sg13g2_fill_2 FILLER_8_954 ();
 sg13g2_fill_1 FILLER_8_956 ();
 sg13g2_fill_2 FILLER_8_962 ();
 sg13g2_fill_1 FILLER_8_969 ();
 sg13g2_decap_4 FILLER_8_975 ();
 sg13g2_fill_1 FILLER_8_979 ();
 sg13g2_fill_1 FILLER_8_989 ();
 sg13g2_decap_4 FILLER_8_998 ();
 sg13g2_decap_8 FILLER_8_1007 ();
 sg13g2_decap_4 FILLER_8_1014 ();
 sg13g2_fill_1 FILLER_8_1018 ();
 sg13g2_decap_4 FILLER_8_1084 ();
 sg13g2_fill_2 FILLER_8_1093 ();
 sg13g2_decap_8 FILLER_8_1115 ();
 sg13g2_fill_2 FILLER_8_1122 ();
 sg13g2_fill_1 FILLER_8_1124 ();
 sg13g2_fill_2 FILLER_8_1134 ();
 sg13g2_fill_1 FILLER_8_1161 ();
 sg13g2_fill_2 FILLER_8_1180 ();
 sg13g2_fill_1 FILLER_8_1182 ();
 sg13g2_decap_4 FILLER_8_1217 ();
 sg13g2_fill_2 FILLER_8_1262 ();
 sg13g2_fill_1 FILLER_8_1264 ();
 sg13g2_fill_2 FILLER_8_1293 ();
 sg13g2_fill_1 FILLER_8_1295 ();
 sg13g2_fill_2 FILLER_8_1333 ();
 sg13g2_fill_1 FILLER_8_1346 ();
 sg13g2_fill_1 FILLER_8_1352 ();
 sg13g2_decap_4 FILLER_8_1375 ();
 sg13g2_fill_2 FILLER_8_1404 ();
 sg13g2_fill_1 FILLER_8_1412 ();
 sg13g2_fill_1 FILLER_8_1447 ();
 sg13g2_fill_2 FILLER_8_1452 ();
 sg13g2_fill_1 FILLER_8_1480 ();
 sg13g2_fill_1 FILLER_8_1493 ();
 sg13g2_fill_1 FILLER_8_1539 ();
 sg13g2_fill_1 FILLER_8_1559 ();
 sg13g2_fill_2 FILLER_8_1586 ();
 sg13g2_fill_1 FILLER_8_1603 ();
 sg13g2_fill_2 FILLER_8_1671 ();
 sg13g2_fill_1 FILLER_8_1673 ();
 sg13g2_decap_4 FILLER_8_1688 ();
 sg13g2_decap_8 FILLER_8_1701 ();
 sg13g2_decap_4 FILLER_8_1708 ();
 sg13g2_fill_2 FILLER_8_1712 ();
 sg13g2_fill_1 FILLER_8_1758 ();
 sg13g2_decap_8 FILLER_8_1775 ();
 sg13g2_fill_1 FILLER_8_1782 ();
 sg13g2_decap_4 FILLER_8_1811 ();
 sg13g2_decap_8 FILLER_8_1821 ();
 sg13g2_decap_4 FILLER_8_1828 ();
 sg13g2_fill_1 FILLER_8_1832 ();
 sg13g2_fill_1 FILLER_8_1837 ();
 sg13g2_fill_2 FILLER_8_1850 ();
 sg13g2_fill_1 FILLER_8_1852 ();
 sg13g2_fill_1 FILLER_8_1872 ();
 sg13g2_decap_4 FILLER_8_1879 ();
 sg13g2_decap_4 FILLER_8_1902 ();
 sg13g2_decap_8 FILLER_8_1910 ();
 sg13g2_decap_8 FILLER_8_1917 ();
 sg13g2_decap_4 FILLER_8_1924 ();
 sg13g2_fill_1 FILLER_8_1928 ();
 sg13g2_decap_4 FILLER_8_1933 ();
 sg13g2_fill_2 FILLER_8_1937 ();
 sg13g2_fill_1 FILLER_8_1999 ();
 sg13g2_decap_4 FILLER_8_2022 ();
 sg13g2_fill_1 FILLER_8_2030 ();
 sg13g2_fill_1 FILLER_8_2039 ();
 sg13g2_fill_1 FILLER_8_2096 ();
 sg13g2_fill_2 FILLER_8_2110 ();
 sg13g2_decap_4 FILLER_8_2156 ();
 sg13g2_fill_2 FILLER_8_2160 ();
 sg13g2_decap_4 FILLER_8_2188 ();
 sg13g2_fill_2 FILLER_8_2192 ();
 sg13g2_decap_8 FILLER_8_2220 ();
 sg13g2_fill_1 FILLER_8_2231 ();
 sg13g2_fill_1 FILLER_8_2236 ();
 sg13g2_decap_4 FILLER_8_2278 ();
 sg13g2_fill_2 FILLER_8_2347 ();
 sg13g2_fill_2 FILLER_8_2422 ();
 sg13g2_fill_1 FILLER_8_2424 ();
 sg13g2_fill_2 FILLER_8_2462 ();
 sg13g2_fill_1 FILLER_8_2464 ();
 sg13g2_fill_2 FILLER_8_2478 ();
 sg13g2_fill_1 FILLER_8_2480 ();
 sg13g2_fill_1 FILLER_8_2509 ();
 sg13g2_decap_4 FILLER_8_2556 ();
 sg13g2_fill_1 FILLER_8_2560 ();
 sg13g2_fill_2 FILLER_8_2612 ();
 sg13g2_fill_1 FILLER_8_2641 ();
 sg13g2_fill_1 FILLER_8_2670 ();
 sg13g2_fill_1 FILLER_8_2720 ();
 sg13g2_fill_2 FILLER_8_2736 ();
 sg13g2_fill_1 FILLER_8_2738 ();
 sg13g2_fill_1 FILLER_8_2752 ();
 sg13g2_decap_4 FILLER_8_2757 ();
 sg13g2_fill_1 FILLER_8_2816 ();
 sg13g2_fill_2 FILLER_8_2849 ();
 sg13g2_fill_1 FILLER_8_2878 ();
 sg13g2_fill_1 FILLER_8_2897 ();
 sg13g2_decap_4 FILLER_8_2911 ();
 sg13g2_decap_4 FILLER_8_2919 ();
 sg13g2_fill_1 FILLER_8_2923 ();
 sg13g2_fill_2 FILLER_8_2952 ();
 sg13g2_fill_1 FILLER_8_2954 ();
 sg13g2_fill_1 FILLER_8_2995 ();
 sg13g2_decap_8 FILLER_8_3030 ();
 sg13g2_decap_8 FILLER_8_3083 ();
 sg13g2_decap_4 FILLER_8_3090 ();
 sg13g2_fill_2 FILLER_8_3098 ();
 sg13g2_fill_1 FILLER_8_3100 ();
 sg13g2_fill_2 FILLER_8_3130 ();
 sg13g2_fill_1 FILLER_8_3132 ();
 sg13g2_fill_2 FILLER_8_3141 ();
 sg13g2_fill_1 FILLER_8_3143 ();
 sg13g2_fill_1 FILLER_8_3164 ();
 sg13g2_decap_8 FILLER_8_3173 ();
 sg13g2_fill_1 FILLER_8_3180 ();
 sg13g2_decap_4 FILLER_8_3194 ();
 sg13g2_decap_4 FILLER_8_3214 ();
 sg13g2_fill_1 FILLER_8_3218 ();
 sg13g2_fill_2 FILLER_8_3227 ();
 sg13g2_fill_2 FILLER_8_3234 ();
 sg13g2_decap_4 FILLER_8_3248 ();
 sg13g2_fill_1 FILLER_8_3252 ();
 sg13g2_fill_1 FILLER_8_3298 ();
 sg13g2_fill_2 FILLER_8_3304 ();
 sg13g2_fill_2 FILLER_8_3311 ();
 sg13g2_fill_1 FILLER_8_3341 ();
 sg13g2_fill_2 FILLER_8_3370 ();
 sg13g2_fill_1 FILLER_8_3372 ();
 sg13g2_decap_8 FILLER_8_3404 ();
 sg13g2_fill_2 FILLER_8_3411 ();
 sg13g2_fill_1 FILLER_8_3413 ();
 sg13g2_decap_4 FILLER_8_3419 ();
 sg13g2_fill_2 FILLER_8_3423 ();
 sg13g2_fill_2 FILLER_8_3461 ();
 sg13g2_fill_1 FILLER_8_3463 ();
 sg13g2_fill_1 FILLER_8_3477 ();
 sg13g2_fill_2 FILLER_8_3491 ();
 sg13g2_fill_1 FILLER_8_3493 ();
 sg13g2_fill_2 FILLER_8_3505 ();
 sg13g2_decap_8 FILLER_8_3530 ();
 sg13g2_fill_2 FILLER_8_3537 ();
 sg13g2_fill_2 FILLER_8_3549 ();
 sg13g2_fill_1 FILLER_8_3551 ();
 sg13g2_decap_4 FILLER_8_3556 ();
 sg13g2_fill_1 FILLER_8_3560 ();
 sg13g2_decap_8 FILLER_8_3570 ();
 sg13g2_fill_2 FILLER_8_3577 ();
 sg13g2_fill_1 FILLER_8_3579 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_2 ();
 sg13g2_fill_2 FILLER_9_21 ();
 sg13g2_fill_2 FILLER_9_32 ();
 sg13g2_fill_1 FILLER_9_50 ();
 sg13g2_fill_1 FILLER_9_56 ();
 sg13g2_fill_2 FILLER_9_65 ();
 sg13g2_fill_1 FILLER_9_67 ();
 sg13g2_fill_1 FILLER_9_73 ();
 sg13g2_fill_2 FILLER_9_99 ();
 sg13g2_fill_1 FILLER_9_101 ();
 sg13g2_fill_1 FILLER_9_112 ();
 sg13g2_fill_2 FILLER_9_141 ();
 sg13g2_fill_1 FILLER_9_143 ();
 sg13g2_fill_1 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_193 ();
 sg13g2_decap_8 FILLER_9_200 ();
 sg13g2_fill_1 FILLER_9_207 ();
 sg13g2_fill_1 FILLER_9_225 ();
 sg13g2_fill_2 FILLER_9_240 ();
 sg13g2_fill_2 FILLER_9_253 ();
 sg13g2_decap_8 FILLER_9_264 ();
 sg13g2_decap_4 FILLER_9_271 ();
 sg13g2_fill_2 FILLER_9_298 ();
 sg13g2_fill_2 FILLER_9_305 ();
 sg13g2_fill_1 FILLER_9_330 ();
 sg13g2_decap_4 FILLER_9_362 ();
 sg13g2_fill_2 FILLER_9_366 ();
 sg13g2_fill_2 FILLER_9_373 ();
 sg13g2_decap_8 FILLER_9_403 ();
 sg13g2_fill_2 FILLER_9_410 ();
 sg13g2_fill_2 FILLER_9_446 ();
 sg13g2_fill_1 FILLER_9_448 ();
 sg13g2_fill_1 FILLER_9_460 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_fill_2 FILLER_9_543 ();
 sg13g2_fill_1 FILLER_9_545 ();
 sg13g2_fill_2 FILLER_9_550 ();
 sg13g2_fill_1 FILLER_9_552 ();
 sg13g2_fill_2 FILLER_9_570 ();
 sg13g2_fill_1 FILLER_9_572 ();
 sg13g2_fill_2 FILLER_9_588 ();
 sg13g2_fill_1 FILLER_9_590 ();
 sg13g2_fill_2 FILLER_9_606 ();
 sg13g2_fill_1 FILLER_9_608 ();
 sg13g2_fill_1 FILLER_9_614 ();
 sg13g2_fill_2 FILLER_9_642 ();
 sg13g2_fill_1 FILLER_9_644 ();
 sg13g2_fill_2 FILLER_9_689 ();
 sg13g2_decap_8 FILLER_9_709 ();
 sg13g2_fill_2 FILLER_9_716 ();
 sg13g2_fill_1 FILLER_9_718 ();
 sg13g2_fill_2 FILLER_9_736 ();
 sg13g2_fill_1 FILLER_9_738 ();
 sg13g2_fill_2 FILLER_9_756 ();
 sg13g2_decap_4 FILLER_9_782 ();
 sg13g2_fill_1 FILLER_9_786 ();
 sg13g2_fill_2 FILLER_9_811 ();
 sg13g2_fill_2 FILLER_9_838 ();
 sg13g2_fill_2 FILLER_9_844 ();
 sg13g2_fill_1 FILLER_9_870 ();
 sg13g2_decap_8 FILLER_9_875 ();
 sg13g2_fill_1 FILLER_9_882 ();
 sg13g2_decap_8 FILLER_9_888 ();
 sg13g2_decap_4 FILLER_9_895 ();
 sg13g2_fill_1 FILLER_9_899 ();
 sg13g2_fill_2 FILLER_9_952 ();
 sg13g2_fill_1 FILLER_9_954 ();
 sg13g2_fill_1 FILLER_9_973 ();
 sg13g2_fill_1 FILLER_9_982 ();
 sg13g2_fill_1 FILLER_9_988 ();
 sg13g2_fill_2 FILLER_9_1041 ();
 sg13g2_fill_2 FILLER_9_1060 ();
 sg13g2_decap_4 FILLER_9_1086 ();
 sg13g2_fill_1 FILLER_9_1090 ();
 sg13g2_fill_1 FILLER_9_1096 ();
 sg13g2_fill_2 FILLER_9_1107 ();
 sg13g2_fill_1 FILLER_9_1109 ();
 sg13g2_fill_1 FILLER_9_1123 ();
 sg13g2_fill_1 FILLER_9_1137 ();
 sg13g2_fill_2 FILLER_9_1168 ();
 sg13g2_fill_2 FILLER_9_1185 ();
 sg13g2_fill_1 FILLER_9_1187 ();
 sg13g2_fill_1 FILLER_9_1197 ();
 sg13g2_fill_2 FILLER_9_1222 ();
 sg13g2_fill_1 FILLER_9_1242 ();
 sg13g2_fill_2 FILLER_9_1264 ();
 sg13g2_fill_1 FILLER_9_1266 ();
 sg13g2_fill_1 FILLER_9_1299 ();
 sg13g2_decap_4 FILLER_9_1321 ();
 sg13g2_fill_1 FILLER_9_1325 ();
 sg13g2_fill_2 FILLER_9_1344 ();
 sg13g2_fill_1 FILLER_9_1346 ();
 sg13g2_decap_8 FILLER_9_1385 ();
 sg13g2_decap_4 FILLER_9_1392 ();
 sg13g2_decap_4 FILLER_9_1418 ();
 sg13g2_fill_1 FILLER_9_1422 ();
 sg13g2_decap_4 FILLER_9_1443 ();
 sg13g2_fill_2 FILLER_9_1447 ();
 sg13g2_fill_2 FILLER_9_1480 ();
 sg13g2_fill_2 FILLER_9_1518 ();
 sg13g2_fill_1 FILLER_9_1520 ();
 sg13g2_fill_1 FILLER_9_1559 ();
 sg13g2_fill_2 FILLER_9_1577 ();
 sg13g2_fill_1 FILLER_9_1579 ();
 sg13g2_decap_4 FILLER_9_1593 ();
 sg13g2_decap_8 FILLER_9_1614 ();
 sg13g2_fill_1 FILLER_9_1621 ();
 sg13g2_fill_1 FILLER_9_1638 ();
 sg13g2_fill_2 FILLER_9_1669 ();
 sg13g2_fill_2 FILLER_9_1731 ();
 sg13g2_fill_1 FILLER_9_1733 ();
 sg13g2_fill_1 FILLER_9_1747 ();
 sg13g2_fill_2 FILLER_9_1785 ();
 sg13g2_fill_1 FILLER_9_1787 ();
 sg13g2_decap_4 FILLER_9_1824 ();
 sg13g2_fill_2 FILLER_9_1861 ();
 sg13g2_fill_1 FILLER_9_1863 ();
 sg13g2_fill_2 FILLER_9_1876 ();
 sg13g2_fill_1 FILLER_9_1878 ();
 sg13g2_fill_1 FILLER_9_1937 ();
 sg13g2_fill_2 FILLER_9_1969 ();
 sg13g2_fill_1 FILLER_9_1971 ();
 sg13g2_fill_2 FILLER_9_2009 ();
 sg13g2_fill_1 FILLER_9_2049 ();
 sg13g2_decap_8 FILLER_9_2081 ();
 sg13g2_decap_8 FILLER_9_2102 ();
 sg13g2_fill_2 FILLER_9_2109 ();
 sg13g2_fill_1 FILLER_9_2111 ();
 sg13g2_decap_4 FILLER_9_2117 ();
 sg13g2_fill_1 FILLER_9_2121 ();
 sg13g2_fill_1 FILLER_9_2125 ();
 sg13g2_decap_8 FILLER_9_2137 ();
 sg13g2_decap_8 FILLER_9_2144 ();
 sg13g2_fill_1 FILLER_9_2164 ();
 sg13g2_fill_1 FILLER_9_2178 ();
 sg13g2_fill_1 FILLER_9_2184 ();
 sg13g2_decap_4 FILLER_9_2193 ();
 sg13g2_fill_1 FILLER_9_2197 ();
 sg13g2_fill_1 FILLER_9_2201 ();
 sg13g2_decap_4 FILLER_9_2211 ();
 sg13g2_fill_2 FILLER_9_2215 ();
 sg13g2_decap_4 FILLER_9_2254 ();
 sg13g2_fill_2 FILLER_9_2295 ();
 sg13g2_fill_2 FILLER_9_2302 ();
 sg13g2_fill_1 FILLER_9_2304 ();
 sg13g2_fill_2 FILLER_9_2314 ();
 sg13g2_fill_2 FILLER_9_2353 ();
 sg13g2_fill_2 FILLER_9_2387 ();
 sg13g2_fill_1 FILLER_9_2389 ();
 sg13g2_fill_2 FILLER_9_2403 ();
 sg13g2_fill_1 FILLER_9_2422 ();
 sg13g2_fill_1 FILLER_9_2428 ();
 sg13g2_fill_2 FILLER_9_2439 ();
 sg13g2_fill_2 FILLER_9_2496 ();
 sg13g2_fill_1 FILLER_9_2498 ();
 sg13g2_fill_2 FILLER_9_2539 ();
 sg13g2_fill_1 FILLER_9_2541 ();
 sg13g2_fill_1 FILLER_9_2629 ();
 sg13g2_fill_1 FILLER_9_2657 ();
 sg13g2_decap_4 FILLER_9_2685 ();
 sg13g2_fill_2 FILLER_9_2689 ();
 sg13g2_decap_4 FILLER_9_2709 ();
 sg13g2_fill_1 FILLER_9_2726 ();
 sg13g2_fill_1 FILLER_9_2793 ();
 sg13g2_decap_4 FILLER_9_2815 ();
 sg13g2_fill_1 FILLER_9_2819 ();
 sg13g2_fill_2 FILLER_9_2873 ();
 sg13g2_fill_1 FILLER_9_2875 ();
 sg13g2_fill_1 FILLER_9_2909 ();
 sg13g2_fill_1 FILLER_9_3004 ();
 sg13g2_fill_2 FILLER_9_3038 ();
 sg13g2_fill_2 FILLER_9_3063 ();
 sg13g2_fill_2 FILLER_9_3158 ();
 sg13g2_decap_4 FILLER_9_3193 ();
 sg13g2_decap_8 FILLER_9_3202 ();
 sg13g2_fill_1 FILLER_9_3209 ();
 sg13g2_fill_1 FILLER_9_3231 ();
 sg13g2_fill_2 FILLER_9_3239 ();
 sg13g2_fill_2 FILLER_9_3250 ();
 sg13g2_fill_2 FILLER_9_3266 ();
 sg13g2_fill_1 FILLER_9_3268 ();
 sg13g2_fill_1 FILLER_9_3290 ();
 sg13g2_fill_1 FILLER_9_3332 ();
 sg13g2_fill_1 FILLER_9_3359 ();
 sg13g2_fill_2 FILLER_9_3366 ();
 sg13g2_decap_8 FILLER_9_3391 ();
 sg13g2_fill_2 FILLER_9_3398 ();
 sg13g2_fill_1 FILLER_9_3400 ();
 sg13g2_fill_2 FILLER_9_3429 ();
 sg13g2_decap_8 FILLER_9_3448 ();
 sg13g2_decap_8 FILLER_9_3455 ();
 sg13g2_decap_8 FILLER_9_3462 ();
 sg13g2_fill_1 FILLER_9_3469 ();
 sg13g2_fill_2 FILLER_9_3483 ();
 sg13g2_fill_1 FILLER_9_3485 ();
 sg13g2_decap_4 FILLER_9_3490 ();
 sg13g2_fill_2 FILLER_9_3499 ();
 sg13g2_fill_1 FILLER_9_3524 ();
 sg13g2_decap_8 FILLER_9_3569 ();
 sg13g2_decap_4 FILLER_9_3576 ();
 sg13g2_fill_2 FILLER_10_22 ();
 sg13g2_fill_1 FILLER_10_24 ();
 sg13g2_fill_2 FILLER_10_34 ();
 sg13g2_decap_8 FILLER_10_72 ();
 sg13g2_decap_4 FILLER_10_79 ();
 sg13g2_fill_2 FILLER_10_83 ();
 sg13g2_fill_2 FILLER_10_94 ();
 sg13g2_fill_1 FILLER_10_96 ();
 sg13g2_fill_1 FILLER_10_123 ();
 sg13g2_fill_1 FILLER_10_140 ();
 sg13g2_fill_2 FILLER_10_154 ();
 sg13g2_fill_1 FILLER_10_156 ();
 sg13g2_fill_1 FILLER_10_185 ();
 sg13g2_fill_2 FILLER_10_211 ();
 sg13g2_fill_1 FILLER_10_256 ();
 sg13g2_decap_4 FILLER_10_265 ();
 sg13g2_fill_2 FILLER_10_269 ();
 sg13g2_fill_1 FILLER_10_280 ();
 sg13g2_decap_4 FILLER_10_285 ();
 sg13g2_fill_2 FILLER_10_325 ();
 sg13g2_fill_1 FILLER_10_327 ();
 sg13g2_fill_2 FILLER_10_332 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_365 ();
 sg13g2_fill_2 FILLER_10_395 ();
 sg13g2_decap_4 FILLER_10_430 ();
 sg13g2_fill_2 FILLER_10_438 ();
 sg13g2_fill_2 FILLER_10_461 ();
 sg13g2_fill_2 FILLER_10_476 ();
 sg13g2_fill_1 FILLER_10_478 ();
 sg13g2_fill_2 FILLER_10_528 ();
 sg13g2_decap_4 FILLER_10_535 ();
 sg13g2_fill_1 FILLER_10_539 ();
 sg13g2_fill_2 FILLER_10_544 ();
 sg13g2_fill_1 FILLER_10_576 ();
 sg13g2_fill_2 FILLER_10_592 ();
 sg13g2_fill_1 FILLER_10_594 ();
 sg13g2_fill_2 FILLER_10_600 ();
 sg13g2_fill_2 FILLER_10_611 ();
 sg13g2_fill_1 FILLER_10_613 ();
 sg13g2_fill_1 FILLER_10_636 ();
 sg13g2_fill_2 FILLER_10_646 ();
 sg13g2_fill_2 FILLER_10_653 ();
 sg13g2_decap_4 FILLER_10_674 ();
 sg13g2_decap_4 FILLER_10_713 ();
 sg13g2_fill_2 FILLER_10_725 ();
 sg13g2_fill_1 FILLER_10_737 ();
 sg13g2_fill_2 FILLER_10_752 ();
 sg13g2_fill_1 FILLER_10_754 ();
 sg13g2_fill_2 FILLER_10_792 ();
 sg13g2_fill_1 FILLER_10_804 ();
 sg13g2_decap_4 FILLER_10_821 ();
 sg13g2_fill_2 FILLER_10_833 ();
 sg13g2_fill_2 FILLER_10_843 ();
 sg13g2_fill_1 FILLER_10_890 ();
 sg13g2_fill_2 FILLER_10_900 ();
 sg13g2_fill_1 FILLER_10_902 ();
 sg13g2_decap_4 FILLER_10_920 ();
 sg13g2_fill_1 FILLER_10_924 ();
 sg13g2_decap_4 FILLER_10_940 ();
 sg13g2_fill_2 FILLER_10_944 ();
 sg13g2_fill_2 FILLER_10_957 ();
 sg13g2_fill_1 FILLER_10_959 ();
 sg13g2_decap_8 FILLER_10_964 ();
 sg13g2_decap_8 FILLER_10_971 ();
 sg13g2_decap_8 FILLER_10_978 ();
 sg13g2_decap_4 FILLER_10_988 ();
 sg13g2_fill_2 FILLER_10_1006 ();
 sg13g2_fill_1 FILLER_10_1008 ();
 sg13g2_fill_1 FILLER_10_1052 ();
 sg13g2_fill_2 FILLER_10_1062 ();
 sg13g2_fill_2 FILLER_10_1076 ();
 sg13g2_decap_8 FILLER_10_1087 ();
 sg13g2_fill_2 FILLER_10_1094 ();
 sg13g2_fill_1 FILLER_10_1096 ();
 sg13g2_decap_4 FILLER_10_1101 ();
 sg13g2_fill_2 FILLER_10_1105 ();
 sg13g2_fill_2 FILLER_10_1135 ();
 sg13g2_fill_1 FILLER_10_1137 ();
 sg13g2_fill_2 FILLER_10_1165 ();
 sg13g2_fill_2 FILLER_10_1248 ();
 sg13g2_fill_1 FILLER_10_1250 ();
 sg13g2_fill_2 FILLER_10_1266 ();
 sg13g2_fill_1 FILLER_10_1268 ();
 sg13g2_fill_1 FILLER_10_1278 ();
 sg13g2_fill_1 FILLER_10_1288 ();
 sg13g2_fill_2 FILLER_10_1300 ();
 sg13g2_fill_1 FILLER_10_1302 ();
 sg13g2_fill_1 FILLER_10_1358 ();
 sg13g2_decap_4 FILLER_10_1388 ();
 sg13g2_decap_8 FILLER_10_1410 ();
 sg13g2_decap_8 FILLER_10_1417 ();
 sg13g2_decap_4 FILLER_10_1424 ();
 sg13g2_fill_2 FILLER_10_1428 ();
 sg13g2_fill_1 FILLER_10_1434 ();
 sg13g2_decap_8 FILLER_10_1440 ();
 sg13g2_decap_4 FILLER_10_1447 ();
 sg13g2_fill_1 FILLER_10_1451 ();
 sg13g2_fill_1 FILLER_10_1511 ();
 sg13g2_fill_2 FILLER_10_1533 ();
 sg13g2_fill_1 FILLER_10_1563 ();
 sg13g2_fill_2 FILLER_10_1585 ();
 sg13g2_fill_1 FILLER_10_1587 ();
 sg13g2_fill_2 FILLER_10_1597 ();
 sg13g2_decap_4 FILLER_10_1613 ();
 sg13g2_fill_1 FILLER_10_1626 ();
 sg13g2_fill_2 FILLER_10_1641 ();
 sg13g2_fill_1 FILLER_10_1671 ();
 sg13g2_fill_1 FILLER_10_1690 ();
 sg13g2_fill_1 FILLER_10_1714 ();
 sg13g2_fill_1 FILLER_10_1759 ();
 sg13g2_fill_1 FILLER_10_1765 ();
 sg13g2_fill_1 FILLER_10_1774 ();
 sg13g2_fill_2 FILLER_10_1784 ();
 sg13g2_decap_8 FILLER_10_1803 ();
 sg13g2_fill_1 FILLER_10_1810 ();
 sg13g2_decap_4 FILLER_10_1872 ();
 sg13g2_fill_2 FILLER_10_1896 ();
 sg13g2_fill_1 FILLER_10_1898 ();
 sg13g2_fill_1 FILLER_10_1941 ();
 sg13g2_decap_4 FILLER_10_1959 ();
 sg13g2_fill_2 FILLER_10_1963 ();
 sg13g2_fill_1 FILLER_10_2045 ();
 sg13g2_fill_1 FILLER_10_2088 ();
 sg13g2_fill_2 FILLER_10_2099 ();
 sg13g2_fill_1 FILLER_10_2101 ();
 sg13g2_fill_2 FILLER_10_2129 ();
 sg13g2_fill_1 FILLER_10_2356 ();
 sg13g2_fill_1 FILLER_10_2468 ();
 sg13g2_fill_1 FILLER_10_2478 ();
 sg13g2_fill_1 FILLER_10_2510 ();
 sg13g2_fill_2 FILLER_10_2516 ();
 sg13g2_fill_2 FILLER_10_2522 ();
 sg13g2_fill_1 FILLER_10_2524 ();
 sg13g2_decap_4 FILLER_10_2538 ();
 sg13g2_fill_2 FILLER_10_2555 ();
 sg13g2_fill_2 FILLER_10_2594 ();
 sg13g2_fill_2 FILLER_10_2636 ();
 sg13g2_decap_4 FILLER_10_2684 ();
 sg13g2_fill_2 FILLER_10_2688 ();
 sg13g2_fill_2 FILLER_10_2717 ();
 sg13g2_fill_1 FILLER_10_2734 ();
 sg13g2_fill_2 FILLER_10_2753 ();
 sg13g2_fill_1 FILLER_10_2755 ();
 sg13g2_fill_1 FILLER_10_2765 ();
 sg13g2_fill_2 FILLER_10_2820 ();
 sg13g2_fill_2 FILLER_10_2861 ();
 sg13g2_fill_2 FILLER_10_2900 ();
 sg13g2_decap_8 FILLER_10_2976 ();
 sg13g2_fill_2 FILLER_10_2983 ();
 sg13g2_fill_1 FILLER_10_2985 ();
 sg13g2_fill_1 FILLER_10_3034 ();
 sg13g2_fill_2 FILLER_10_3057 ();
 sg13g2_fill_1 FILLER_10_3108 ();
 sg13g2_fill_1 FILLER_10_3126 ();
 sg13g2_fill_2 FILLER_10_3162 ();
 sg13g2_fill_1 FILLER_10_3164 ();
 sg13g2_decap_4 FILLER_10_3187 ();
 sg13g2_decap_4 FILLER_10_3201 ();
 sg13g2_fill_2 FILLER_10_3288 ();
 sg13g2_fill_1 FILLER_10_3290 ();
 sg13g2_fill_1 FILLER_10_3315 ();
 sg13g2_fill_1 FILLER_10_3358 ();
 sg13g2_fill_1 FILLER_10_3378 ();
 sg13g2_fill_2 FILLER_10_3405 ();
 sg13g2_fill_2 FILLER_10_3413 ();
 sg13g2_decap_4 FILLER_10_3452 ();
 sg13g2_decap_8 FILLER_10_3484 ();
 sg13g2_fill_2 FILLER_10_3491 ();
 sg13g2_fill_2 FILLER_10_3510 ();
 sg13g2_fill_2 FILLER_10_3541 ();
 sg13g2_fill_1 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_42 ();
 sg13g2_fill_1 FILLER_11_44 ();
 sg13g2_fill_2 FILLER_11_50 ();
 sg13g2_fill_1 FILLER_11_52 ();
 sg13g2_fill_1 FILLER_11_118 ();
 sg13g2_fill_1 FILLER_11_193 ();
 sg13g2_decap_4 FILLER_11_234 ();
 sg13g2_fill_1 FILLER_11_238 ();
 sg13g2_fill_2 FILLER_11_285 ();
 sg13g2_fill_2 FILLER_11_314 ();
 sg13g2_fill_1 FILLER_11_316 ();
 sg13g2_fill_2 FILLER_11_350 ();
 sg13g2_fill_1 FILLER_11_352 ();
 sg13g2_fill_1 FILLER_11_381 ();
 sg13g2_fill_1 FILLER_11_395 ();
 sg13g2_fill_1 FILLER_11_434 ();
 sg13g2_fill_2 FILLER_11_448 ();
 sg13g2_fill_2 FILLER_11_459 ();
 sg13g2_fill_2 FILLER_11_473 ();
 sg13g2_fill_1 FILLER_11_475 ();
 sg13g2_fill_1 FILLER_11_481 ();
 sg13g2_fill_1 FILLER_11_543 ();
 sg13g2_decap_8 FILLER_11_564 ();
 sg13g2_decap_4 FILLER_11_571 ();
 sg13g2_fill_1 FILLER_11_575 ();
 sg13g2_fill_1 FILLER_11_584 ();
 sg13g2_fill_2 FILLER_11_594 ();
 sg13g2_fill_1 FILLER_11_596 ();
 sg13g2_fill_2 FILLER_11_607 ();
 sg13g2_fill_2 FILLER_11_614 ();
 sg13g2_fill_1 FILLER_11_616 ();
 sg13g2_fill_2 FILLER_11_643 ();
 sg13g2_fill_1 FILLER_11_645 ();
 sg13g2_fill_2 FILLER_11_662 ();
 sg13g2_fill_1 FILLER_11_664 ();
 sg13g2_fill_1 FILLER_11_686 ();
 sg13g2_fill_1 FILLER_11_707 ();
 sg13g2_fill_2 FILLER_11_752 ();
 sg13g2_fill_1 FILLER_11_768 ();
 sg13g2_decap_8 FILLER_11_785 ();
 sg13g2_fill_2 FILLER_11_792 ();
 sg13g2_fill_2 FILLER_11_814 ();
 sg13g2_fill_2 FILLER_11_820 ();
 sg13g2_fill_1 FILLER_11_822 ();
 sg13g2_fill_1 FILLER_11_832 ();
 sg13g2_decap_8 FILLER_11_862 ();
 sg13g2_decap_4 FILLER_11_882 ();
 sg13g2_fill_1 FILLER_11_906 ();
 sg13g2_decap_8 FILLER_11_915 ();
 sg13g2_fill_2 FILLER_11_932 ();
 sg13g2_fill_1 FILLER_11_934 ();
 sg13g2_fill_2 FILLER_11_960 ();
 sg13g2_fill_2 FILLER_11_970 ();
 sg13g2_fill_1 FILLER_11_985 ();
 sg13g2_fill_1 FILLER_11_994 ();
 sg13g2_decap_4 FILLER_11_1008 ();
 sg13g2_fill_1 FILLER_11_1056 ();
 sg13g2_fill_2 FILLER_11_1069 ();
 sg13g2_fill_1 FILLER_11_1071 ();
 sg13g2_decap_8 FILLER_11_1085 ();
 sg13g2_fill_2 FILLER_11_1096 ();
 sg13g2_fill_1 FILLER_11_1098 ();
 sg13g2_fill_1 FILLER_11_1109 ();
 sg13g2_fill_2 FILLER_11_1126 ();
 sg13g2_fill_1 FILLER_11_1128 ();
 sg13g2_fill_2 FILLER_11_1148 ();
 sg13g2_fill_1 FILLER_11_1150 ();
 sg13g2_decap_4 FILLER_11_1171 ();
 sg13g2_fill_2 FILLER_11_1175 ();
 sg13g2_fill_2 FILLER_11_1190 ();
 sg13g2_fill_1 FILLER_11_1192 ();
 sg13g2_decap_8 FILLER_11_1196 ();
 sg13g2_fill_2 FILLER_11_1203 ();
 sg13g2_fill_1 FILLER_11_1205 ();
 sg13g2_fill_2 FILLER_11_1219 ();
 sg13g2_fill_2 FILLER_11_1259 ();
 sg13g2_fill_2 FILLER_11_1294 ();
 sg13g2_fill_1 FILLER_11_1296 ();
 sg13g2_fill_2 FILLER_11_1310 ();
 sg13g2_fill_1 FILLER_11_1312 ();
 sg13g2_fill_2 FILLER_11_1326 ();
 sg13g2_fill_2 FILLER_11_1352 ();
 sg13g2_fill_2 FILLER_11_1357 ();
 sg13g2_decap_8 FILLER_11_1362 ();
 sg13g2_fill_1 FILLER_11_1369 ();
 sg13g2_decap_8 FILLER_11_1391 ();
 sg13g2_decap_8 FILLER_11_1398 ();
 sg13g2_fill_1 FILLER_11_1405 ();
 sg13g2_fill_2 FILLER_11_1410 ();
 sg13g2_fill_1 FILLER_11_1412 ();
 sg13g2_fill_2 FILLER_11_1453 ();
 sg13g2_fill_2 FILLER_11_1481 ();
 sg13g2_fill_1 FILLER_11_1491 ();
 sg13g2_fill_1 FILLER_11_1537 ();
 sg13g2_fill_2 FILLER_11_1554 ();
 sg13g2_fill_1 FILLER_11_1586 ();
 sg13g2_fill_2 FILLER_11_1592 ();
 sg13g2_fill_1 FILLER_11_1594 ();
 sg13g2_fill_2 FILLER_11_1620 ();
 sg13g2_fill_1 FILLER_11_1622 ();
 sg13g2_fill_2 FILLER_11_1662 ();
 sg13g2_fill_1 FILLER_11_1664 ();
 sg13g2_fill_2 FILLER_11_1695 ();
 sg13g2_fill_2 FILLER_11_1710 ();
 sg13g2_fill_1 FILLER_11_1712 ();
 sg13g2_decap_4 FILLER_11_1745 ();
 sg13g2_fill_1 FILLER_11_1749 ();
 sg13g2_decap_4 FILLER_11_1794 ();
 sg13g2_fill_1 FILLER_11_1825 ();
 sg13g2_fill_2 FILLER_11_1830 ();
 sg13g2_fill_1 FILLER_11_1832 ();
 sg13g2_fill_2 FILLER_11_1863 ();
 sg13g2_decap_4 FILLER_11_1875 ();
 sg13g2_fill_2 FILLER_11_1889 ();
 sg13g2_fill_2 FILLER_11_1899 ();
 sg13g2_fill_1 FILLER_11_1901 ();
 sg13g2_fill_1 FILLER_11_1933 ();
 sg13g2_decap_4 FILLER_11_1985 ();
 sg13g2_fill_1 FILLER_11_1989 ();
 sg13g2_fill_2 FILLER_11_2026 ();
 sg13g2_fill_1 FILLER_11_2028 ();
 sg13g2_fill_2 FILLER_11_2038 ();
 sg13g2_fill_1 FILLER_11_2058 ();
 sg13g2_fill_2 FILLER_11_2082 ();
 sg13g2_fill_2 FILLER_11_2113 ();
 sg13g2_fill_1 FILLER_11_2318 ();
 sg13g2_fill_1 FILLER_11_2419 ();
 sg13g2_fill_2 FILLER_11_2481 ();
 sg13g2_fill_2 FILLER_11_2541 ();
 sg13g2_fill_1 FILLER_11_2543 ();
 sg13g2_fill_2 FILLER_11_2571 ();
 sg13g2_fill_2 FILLER_11_2592 ();
 sg13g2_fill_1 FILLER_11_2607 ();
 sg13g2_fill_2 FILLER_11_2718 ();
 sg13g2_fill_2 FILLER_11_2762 ();
 sg13g2_fill_1 FILLER_11_2764 ();
 sg13g2_fill_2 FILLER_11_2784 ();
 sg13g2_fill_1 FILLER_11_2786 ();
 sg13g2_fill_1 FILLER_11_2830 ();
 sg13g2_fill_2 FILLER_11_2910 ();
 sg13g2_fill_1 FILLER_11_2925 ();
 sg13g2_fill_1 FILLER_11_2945 ();
 sg13g2_fill_2 FILLER_11_2964 ();
 sg13g2_fill_1 FILLER_11_2966 ();
 sg13g2_fill_2 FILLER_11_3053 ();
 sg13g2_fill_1 FILLER_11_3055 ();
 sg13g2_fill_2 FILLER_11_3090 ();
 sg13g2_fill_1 FILLER_11_3097 ();
 sg13g2_fill_2 FILLER_11_3150 ();
 sg13g2_fill_2 FILLER_11_3166 ();
 sg13g2_fill_1 FILLER_11_3168 ();
 sg13g2_fill_2 FILLER_11_3182 ();
 sg13g2_fill_1 FILLER_11_3190 ();
 sg13g2_fill_2 FILLER_11_3209 ();
 sg13g2_fill_1 FILLER_11_3228 ();
 sg13g2_fill_1 FILLER_11_3249 ();
 sg13g2_fill_2 FILLER_11_3387 ();
 sg13g2_fill_1 FILLER_11_3389 ();
 sg13g2_fill_2 FILLER_11_3403 ();
 sg13g2_fill_1 FILLER_11_3427 ();
 sg13g2_decap_4 FILLER_11_3475 ();
 sg13g2_fill_2 FILLER_11_3479 ();
 sg13g2_fill_2 FILLER_11_3505 ();
 sg13g2_fill_1 FILLER_11_3535 ();
 sg13g2_fill_2 FILLER_11_3547 ();
 sg13g2_fill_2 FILLER_11_3567 ();
 sg13g2_fill_2 FILLER_11_3578 ();
 sg13g2_decap_4 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_4 ();
 sg13g2_fill_2 FILLER_12_10 ();
 sg13g2_fill_1 FILLER_12_12 ();
 sg13g2_fill_1 FILLER_12_22 ();
 sg13g2_fill_2 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_38 ();
 sg13g2_fill_1 FILLER_12_45 ();
 sg13g2_decap_4 FILLER_12_69 ();
 sg13g2_fill_2 FILLER_12_93 ();
 sg13g2_fill_1 FILLER_12_95 ();
 sg13g2_fill_2 FILLER_12_118 ();
 sg13g2_fill_1 FILLER_12_126 ();
 sg13g2_fill_1 FILLER_12_136 ();
 sg13g2_fill_2 FILLER_12_151 ();
 sg13g2_fill_2 FILLER_12_158 ();
 sg13g2_fill_1 FILLER_12_173 ();
 sg13g2_fill_1 FILLER_12_189 ();
 sg13g2_fill_1 FILLER_12_202 ();
 sg13g2_fill_1 FILLER_12_208 ();
 sg13g2_fill_2 FILLER_12_235 ();
 sg13g2_fill_2 FILLER_12_261 ();
 sg13g2_fill_2 FILLER_12_321 ();
 sg13g2_fill_1 FILLER_12_323 ();
 sg13g2_fill_2 FILLER_12_338 ();
 sg13g2_fill_1 FILLER_12_340 ();
 sg13g2_fill_2 FILLER_12_417 ();
 sg13g2_fill_1 FILLER_12_419 ();
 sg13g2_fill_1 FILLER_12_476 ();
 sg13g2_fill_2 FILLER_12_490 ();
 sg13g2_fill_1 FILLER_12_492 ();
 sg13g2_fill_2 FILLER_12_498 ();
 sg13g2_fill_1 FILLER_12_500 ();
 sg13g2_fill_2 FILLER_12_524 ();
 sg13g2_fill_1 FILLER_12_588 ();
 sg13g2_decap_4 FILLER_12_601 ();
 sg13g2_decap_8 FILLER_12_617 ();
 sg13g2_fill_2 FILLER_12_624 ();
 sg13g2_fill_1 FILLER_12_626 ();
 sg13g2_decap_4 FILLER_12_643 ();
 sg13g2_decap_8 FILLER_12_659 ();
 sg13g2_decap_4 FILLER_12_666 ();
 sg13g2_fill_2 FILLER_12_696 ();
 sg13g2_fill_1 FILLER_12_698 ();
 sg13g2_fill_1 FILLER_12_723 ();
 sg13g2_fill_1 FILLER_12_742 ();
 sg13g2_fill_1 FILLER_12_766 ();
 sg13g2_decap_4 FILLER_12_773 ();
 sg13g2_fill_2 FILLER_12_783 ();
 sg13g2_fill_1 FILLER_12_789 ();
 sg13g2_fill_2 FILLER_12_797 ();
 sg13g2_fill_1 FILLER_12_799 ();
 sg13g2_fill_2 FILLER_12_809 ();
 sg13g2_fill_2 FILLER_12_848 ();
 sg13g2_fill_2 FILLER_12_862 ();
 sg13g2_fill_2 FILLER_12_908 ();
 sg13g2_fill_1 FILLER_12_910 ();
 sg13g2_fill_1 FILLER_12_919 ();
 sg13g2_fill_1 FILLER_12_940 ();
 sg13g2_decap_4 FILLER_12_961 ();
 sg13g2_fill_1 FILLER_12_965 ();
 sg13g2_fill_2 FILLER_12_1004 ();
 sg13g2_fill_1 FILLER_12_1006 ();
 sg13g2_fill_1 FILLER_12_1014 ();
 sg13g2_fill_2 FILLER_12_1044 ();
 sg13g2_fill_2 FILLER_12_1060 ();
 sg13g2_fill_2 FILLER_12_1083 ();
 sg13g2_fill_1 FILLER_12_1085 ();
 sg13g2_fill_2 FILLER_12_1101 ();
 sg13g2_fill_1 FILLER_12_1103 ();
 sg13g2_fill_1 FILLER_12_1121 ();
 sg13g2_fill_2 FILLER_12_1153 ();
 sg13g2_fill_1 FILLER_12_1187 ();
 sg13g2_fill_2 FILLER_12_1250 ();
 sg13g2_fill_1 FILLER_12_1252 ();
 sg13g2_fill_2 FILLER_12_1274 ();
 sg13g2_fill_1 FILLER_12_1276 ();
 sg13g2_fill_1 FILLER_12_1291 ();
 sg13g2_fill_2 FILLER_12_1309 ();
 sg13g2_fill_1 FILLER_12_1311 ();
 sg13g2_decap_8 FILLER_12_1347 ();
 sg13g2_fill_2 FILLER_12_1354 ();
 sg13g2_fill_1 FILLER_12_1374 ();
 sg13g2_fill_2 FILLER_12_1379 ();
 sg13g2_fill_1 FILLER_12_1381 ();
 sg13g2_decap_8 FILLER_12_1385 ();
 sg13g2_fill_2 FILLER_12_1392 ();
 sg13g2_fill_2 FILLER_12_1435 ();
 sg13g2_fill_1 FILLER_12_1437 ();
 sg13g2_fill_2 FILLER_12_1453 ();
 sg13g2_fill_2 FILLER_12_1461 ();
 sg13g2_fill_1 FILLER_12_1463 ();
 sg13g2_fill_1 FILLER_12_1483 ();
 sg13g2_fill_1 FILLER_12_1498 ();
 sg13g2_fill_2 FILLER_12_1512 ();
 sg13g2_fill_2 FILLER_12_1581 ();
 sg13g2_fill_1 FILLER_12_1617 ();
 sg13g2_fill_2 FILLER_12_1627 ();
 sg13g2_fill_1 FILLER_12_1629 ();
 sg13g2_fill_1 FILLER_12_1685 ();
 sg13g2_fill_2 FILLER_12_1705 ();
 sg13g2_fill_1 FILLER_12_1722 ();
 sg13g2_fill_1 FILLER_12_1733 ();
 sg13g2_fill_2 FILLER_12_1743 ();
 sg13g2_fill_2 FILLER_12_1771 ();
 sg13g2_decap_4 FILLER_12_1792 ();
 sg13g2_decap_4 FILLER_12_1823 ();
 sg13g2_fill_2 FILLER_12_1827 ();
 sg13g2_decap_4 FILLER_12_1883 ();
 sg13g2_fill_1 FILLER_12_1915 ();
 sg13g2_fill_1 FILLER_12_1929 ();
 sg13g2_fill_2 FILLER_12_1980 ();
 sg13g2_fill_1 FILLER_12_1982 ();
 sg13g2_fill_2 FILLER_12_2011 ();
 sg13g2_fill_2 FILLER_12_2058 ();
 sg13g2_fill_1 FILLER_12_2082 ();
 sg13g2_fill_1 FILLER_12_2106 ();
 sg13g2_decap_8 FILLER_12_2133 ();
 sg13g2_fill_2 FILLER_12_2153 ();
 sg13g2_fill_1 FILLER_12_2160 ();
 sg13g2_fill_1 FILLER_12_2174 ();
 sg13g2_fill_1 FILLER_12_2197 ();
 sg13g2_fill_2 FILLER_12_2220 ();
 sg13g2_fill_1 FILLER_12_2222 ();
 sg13g2_fill_1 FILLER_12_2236 ();
 sg13g2_fill_2 FILLER_12_2245 ();
 sg13g2_fill_1 FILLER_12_2247 ();
 sg13g2_fill_2 FILLER_12_2267 ();
 sg13g2_fill_1 FILLER_12_2269 ();
 sg13g2_fill_2 FILLER_12_2294 ();
 sg13g2_fill_2 FILLER_12_2341 ();
 sg13g2_fill_1 FILLER_12_2343 ();
 sg13g2_fill_2 FILLER_12_2388 ();
 sg13g2_fill_1 FILLER_12_2390 ();
 sg13g2_fill_2 FILLER_12_2400 ();
 sg13g2_fill_1 FILLER_12_2408 ();
 sg13g2_fill_1 FILLER_12_2477 ();
 sg13g2_fill_2 FILLER_12_2494 ();
 sg13g2_fill_2 FILLER_12_2529 ();
 sg13g2_fill_1 FILLER_12_2531 ();
 sg13g2_fill_2 FILLER_12_2646 ();
 sg13g2_fill_1 FILLER_12_2683 ();
 sg13g2_fill_1 FILLER_12_2719 ();
 sg13g2_fill_1 FILLER_12_2810 ();
 sg13g2_fill_2 FILLER_12_2839 ();
 sg13g2_fill_1 FILLER_12_2841 ();
 sg13g2_fill_2 FILLER_12_2884 ();
 sg13g2_decap_4 FILLER_12_2926 ();
 sg13g2_fill_2 FILLER_12_2935 ();
 sg13g2_fill_1 FILLER_12_2943 ();
 sg13g2_fill_1 FILLER_12_2954 ();
 sg13g2_decap_4 FILLER_12_2968 ();
 sg13g2_fill_1 FILLER_12_2972 ();
 sg13g2_fill_2 FILLER_12_3008 ();
 sg13g2_fill_1 FILLER_12_3010 ();
 sg13g2_fill_2 FILLER_12_3088 ();
 sg13g2_fill_1 FILLER_12_3090 ();
 sg13g2_fill_2 FILLER_12_3096 ();
 sg13g2_fill_2 FILLER_12_3140 ();
 sg13g2_fill_2 FILLER_12_3155 ();
 sg13g2_fill_2 FILLER_12_3204 ();
 sg13g2_fill_1 FILLER_12_3206 ();
 sg13g2_fill_1 FILLER_12_3321 ();
 sg13g2_fill_1 FILLER_12_3380 ();
 sg13g2_fill_1 FILLER_12_3399 ();
 sg13g2_fill_2 FILLER_12_3413 ();
 sg13g2_decap_4 FILLER_12_3432 ();
 sg13g2_decap_4 FILLER_12_3446 ();
 sg13g2_fill_1 FILLER_12_3458 ();
 sg13g2_fill_2 FILLER_12_3472 ();
 sg13g2_fill_2 FILLER_12_3484 ();
 sg13g2_fill_2 FILLER_12_3496 ();
 sg13g2_decap_8 FILLER_12_3509 ();
 sg13g2_fill_2 FILLER_12_3537 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_29 ();
 sg13g2_decap_8 FILLER_13_43 ();
 sg13g2_decap_4 FILLER_13_50 ();
 sg13g2_decap_8 FILLER_13_64 ();
 sg13g2_decap_8 FILLER_13_71 ();
 sg13g2_fill_1 FILLER_13_78 ();
 sg13g2_fill_2 FILLER_13_98 ();
 sg13g2_fill_1 FILLER_13_167 ();
 sg13g2_decap_8 FILLER_13_187 ();
 sg13g2_fill_1 FILLER_13_235 ();
 sg13g2_fill_1 FILLER_13_248 ();
 sg13g2_decap_4 FILLER_13_287 ();
 sg13g2_decap_4 FILLER_13_327 ();
 sg13g2_fill_1 FILLER_13_336 ();
 sg13g2_fill_1 FILLER_13_350 ();
 sg13g2_fill_1 FILLER_13_365 ();
 sg13g2_fill_1 FILLER_13_392 ();
 sg13g2_fill_1 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_412 ();
 sg13g2_fill_1 FILLER_13_484 ();
 sg13g2_fill_1 FILLER_13_521 ();
 sg13g2_fill_2 FILLER_13_530 ();
 sg13g2_fill_1 FILLER_13_532 ();
 sg13g2_fill_2 FILLER_13_543 ();
 sg13g2_fill_2 FILLER_13_558 ();
 sg13g2_fill_1 FILLER_13_560 ();
 sg13g2_decap_4 FILLER_13_593 ();
 sg13g2_fill_1 FILLER_13_597 ();
 sg13g2_fill_1 FILLER_13_608 ();
 sg13g2_decap_4 FILLER_13_613 ();
 sg13g2_fill_1 FILLER_13_617 ();
 sg13g2_fill_2 FILLER_13_656 ();
 sg13g2_decap_4 FILLER_13_697 ();
 sg13g2_fill_1 FILLER_13_701 ();
 sg13g2_fill_2 FILLER_13_761 ();
 sg13g2_fill_1 FILLER_13_772 ();
 sg13g2_fill_1 FILLER_13_779 ();
 sg13g2_fill_1 FILLER_13_852 ();
 sg13g2_fill_2 FILLER_13_863 ();
 sg13g2_fill_1 FILLER_13_865 ();
 sg13g2_decap_8 FILLER_13_874 ();
 sg13g2_decap_8 FILLER_13_881 ();
 sg13g2_fill_2 FILLER_13_919 ();
 sg13g2_fill_2 FILLER_13_953 ();
 sg13g2_fill_1 FILLER_13_964 ();
 sg13g2_fill_2 FILLER_13_984 ();
 sg13g2_fill_1 FILLER_13_986 ();
 sg13g2_fill_1 FILLER_13_1059 ();
 sg13g2_fill_2 FILLER_13_1065 ();
 sg13g2_fill_1 FILLER_13_1080 ();
 sg13g2_fill_2 FILLER_13_1089 ();
 sg13g2_fill_1 FILLER_13_1091 ();
 sg13g2_decap_8 FILLER_13_1110 ();
 sg13g2_fill_1 FILLER_13_1117 ();
 sg13g2_fill_2 FILLER_13_1127 ();
 sg13g2_fill_1 FILLER_13_1129 ();
 sg13g2_fill_1 FILLER_13_1162 ();
 sg13g2_fill_1 FILLER_13_1255 ();
 sg13g2_fill_2 FILLER_13_1261 ();
 sg13g2_fill_2 FILLER_13_1274 ();
 sg13g2_decap_4 FILLER_13_1285 ();
 sg13g2_fill_1 FILLER_13_1289 ();
 sg13g2_decap_8 FILLER_13_1347 ();
 sg13g2_fill_1 FILLER_13_1382 ();
 sg13g2_decap_4 FILLER_13_1410 ();
 sg13g2_fill_1 FILLER_13_1414 ();
 sg13g2_fill_1 FILLER_13_1448 ();
 sg13g2_fill_2 FILLER_13_1482 ();
 sg13g2_fill_2 FILLER_13_1570 ();
 sg13g2_fill_1 FILLER_13_1572 ();
 sg13g2_fill_2 FILLER_13_1608 ();
 sg13g2_fill_2 FILLER_13_1638 ();
 sg13g2_fill_2 FILLER_13_1683 ();
 sg13g2_decap_8 FILLER_13_1785 ();
 sg13g2_fill_2 FILLER_13_1792 ();
 sg13g2_fill_1 FILLER_13_1794 ();
 sg13g2_decap_4 FILLER_13_1840 ();
 sg13g2_fill_2 FILLER_13_1844 ();
 sg13g2_fill_1 FILLER_13_1864 ();
 sg13g2_fill_2 FILLER_13_1882 ();
 sg13g2_fill_1 FILLER_13_1884 ();
 sg13g2_fill_2 FILLER_13_1919 ();
 sg13g2_decap_4 FILLER_13_1934 ();
 sg13g2_fill_1 FILLER_13_1938 ();
 sg13g2_fill_2 FILLER_13_1963 ();
 sg13g2_fill_2 FILLER_13_1974 ();
 sg13g2_fill_2 FILLER_13_2042 ();
 sg13g2_fill_1 FILLER_13_2044 ();
 sg13g2_fill_2 FILLER_13_2073 ();
 sg13g2_fill_2 FILLER_13_2119 ();
 sg13g2_fill_1 FILLER_13_2180 ();
 sg13g2_fill_1 FILLER_13_2190 ();
 sg13g2_fill_2 FILLER_13_2300 ();
 sg13g2_fill_2 FILLER_13_2311 ();
 sg13g2_fill_2 FILLER_13_2361 ();
 sg13g2_fill_1 FILLER_13_2399 ();
 sg13g2_fill_2 FILLER_13_2427 ();
 sg13g2_fill_1 FILLER_13_2470 ();
 sg13g2_fill_2 FILLER_13_2496 ();
 sg13g2_fill_2 FILLER_13_2512 ();
 sg13g2_fill_1 FILLER_13_2514 ();
 sg13g2_fill_2 FILLER_13_2548 ();
 sg13g2_fill_1 FILLER_13_2550 ();
 sg13g2_fill_1 FILLER_13_2613 ();
 sg13g2_fill_2 FILLER_13_2632 ();
 sg13g2_fill_2 FILLER_13_2662 ();
 sg13g2_fill_1 FILLER_13_2664 ();
 sg13g2_fill_2 FILLER_13_2764 ();
 sg13g2_fill_1 FILLER_13_2766 ();
 sg13g2_fill_2 FILLER_13_2892 ();
 sg13g2_fill_2 FILLER_13_2939 ();
 sg13g2_fill_2 FILLER_13_2954 ();
 sg13g2_fill_1 FILLER_13_3033 ();
 sg13g2_fill_2 FILLER_13_3052 ();
 sg13g2_fill_1 FILLER_13_3054 ();
 sg13g2_fill_1 FILLER_13_3088 ();
 sg13g2_fill_2 FILLER_13_3099 ();
 sg13g2_fill_2 FILLER_13_3123 ();
 sg13g2_fill_1 FILLER_13_3125 ();
 sg13g2_fill_2 FILLER_13_3163 ();
 sg13g2_fill_1 FILLER_13_3165 ();
 sg13g2_fill_1 FILLER_13_3236 ();
 sg13g2_fill_2 FILLER_13_3259 ();
 sg13g2_fill_1 FILLER_13_3261 ();
 sg13g2_fill_1 FILLER_13_3289 ();
 sg13g2_fill_2 FILLER_13_3300 ();
 sg13g2_fill_1 FILLER_13_3302 ();
 sg13g2_fill_2 FILLER_13_3363 ();
 sg13g2_fill_1 FILLER_13_3381 ();
 sg13g2_fill_2 FILLER_13_3395 ();
 sg13g2_fill_1 FILLER_13_3397 ();
 sg13g2_decap_4 FILLER_13_3418 ();
 sg13g2_fill_1 FILLER_13_3422 ();
 sg13g2_decap_4 FILLER_13_3435 ();
 sg13g2_fill_2 FILLER_13_3489 ();
 sg13g2_fill_1 FILLER_13_3491 ();
 sg13g2_fill_2 FILLER_13_3496 ();
 sg13g2_fill_1 FILLER_13_3498 ();
 sg13g2_fill_1 FILLER_13_3515 ();
 sg13g2_fill_1 FILLER_13_3542 ();
 sg13g2_decap_4 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_4 ();
 sg13g2_decap_8 FILLER_14_10 ();
 sg13g2_fill_1 FILLER_14_17 ();
 sg13g2_fill_2 FILLER_14_27 ();
 sg13g2_fill_2 FILLER_14_43 ();
 sg13g2_fill_1 FILLER_14_63 ();
 sg13g2_fill_2 FILLER_14_74 ();
 sg13g2_fill_2 FILLER_14_81 ();
 sg13g2_fill_1 FILLER_14_83 ();
 sg13g2_fill_2 FILLER_14_99 ();
 sg13g2_fill_1 FILLER_14_101 ();
 sg13g2_fill_2 FILLER_14_115 ();
 sg13g2_fill_2 FILLER_14_177 ();
 sg13g2_decap_4 FILLER_14_187 ();
 sg13g2_fill_2 FILLER_14_201 ();
 sg13g2_fill_2 FILLER_14_213 ();
 sg13g2_decap_8 FILLER_14_220 ();
 sg13g2_fill_2 FILLER_14_227 ();
 sg13g2_fill_1 FILLER_14_248 ();
 sg13g2_fill_1 FILLER_14_318 ();
 sg13g2_fill_2 FILLER_14_340 ();
 sg13g2_fill_1 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_422 ();
 sg13g2_fill_2 FILLER_14_495 ();
 sg13g2_fill_1 FILLER_14_502 ();
 sg13g2_fill_1 FILLER_14_517 ();
 sg13g2_fill_2 FILLER_14_536 ();
 sg13g2_fill_2 FILLER_14_607 ();
 sg13g2_fill_1 FILLER_14_609 ();
 sg13g2_fill_2 FILLER_14_620 ();
 sg13g2_fill_1 FILLER_14_622 ();
 sg13g2_fill_1 FILLER_14_661 ();
 sg13g2_fill_2 FILLER_14_690 ();
 sg13g2_fill_2 FILLER_14_713 ();
 sg13g2_fill_2 FILLER_14_731 ();
 sg13g2_fill_1 FILLER_14_744 ();
 sg13g2_fill_2 FILLER_14_787 ();
 sg13g2_fill_1 FILLER_14_789 ();
 sg13g2_fill_1 FILLER_14_850 ();
 sg13g2_fill_1 FILLER_14_856 ();
 sg13g2_fill_2 FILLER_14_864 ();
 sg13g2_fill_1 FILLER_14_881 ();
 sg13g2_fill_1 FILLER_14_957 ();
 sg13g2_fill_1 FILLER_14_963 ();
 sg13g2_fill_2 FILLER_14_998 ();
 sg13g2_fill_1 FILLER_14_1000 ();
 sg13g2_fill_1 FILLER_14_1015 ();
 sg13g2_fill_2 FILLER_14_1030 ();
 sg13g2_fill_1 FILLER_14_1091 ();
 sg13g2_decap_4 FILLER_14_1104 ();
 sg13g2_fill_1 FILLER_14_1180 ();
 sg13g2_fill_1 FILLER_14_1263 ();
 sg13g2_fill_1 FILLER_14_1304 ();
 sg13g2_fill_2 FILLER_14_1318 ();
 sg13g2_fill_1 FILLER_14_1320 ();
 sg13g2_decap_4 FILLER_14_1330 ();
 sg13g2_fill_2 FILLER_14_1334 ();
 sg13g2_decap_8 FILLER_14_1354 ();
 sg13g2_fill_1 FILLER_14_1361 ();
 sg13g2_fill_2 FILLER_14_1371 ();
 sg13g2_fill_1 FILLER_14_1373 ();
 sg13g2_fill_1 FILLER_14_1424 ();
 sg13g2_fill_1 FILLER_14_1438 ();
 sg13g2_fill_1 FILLER_14_1453 ();
 sg13g2_fill_1 FILLER_14_1463 ();
 sg13g2_fill_1 FILLER_14_1477 ();
 sg13g2_fill_2 FILLER_14_1502 ();
 sg13g2_fill_2 FILLER_14_1523 ();
 sg13g2_fill_2 FILLER_14_1592 ();
 sg13g2_fill_2 FILLER_14_1598 ();
 sg13g2_fill_2 FILLER_14_1618 ();
 sg13g2_fill_2 FILLER_14_1657 ();
 sg13g2_fill_2 FILLER_14_1708 ();
 sg13g2_fill_1 FILLER_14_1710 ();
 sg13g2_fill_1 FILLER_14_1814 ();
 sg13g2_decap_8 FILLER_14_1824 ();
 sg13g2_fill_2 FILLER_14_1831 ();
 sg13g2_decap_4 FILLER_14_1841 ();
 sg13g2_decap_4 FILLER_14_1882 ();
 sg13g2_fill_2 FILLER_14_1886 ();
 sg13g2_fill_2 FILLER_14_1948 ();
 sg13g2_fill_1 FILLER_14_1950 ();
 sg13g2_fill_2 FILLER_14_1984 ();
 sg13g2_fill_1 FILLER_14_2000 ();
 sg13g2_fill_2 FILLER_14_2015 ();
 sg13g2_fill_1 FILLER_14_2085 ();
 sg13g2_fill_2 FILLER_14_2123 ();
 sg13g2_fill_1 FILLER_14_2125 ();
 sg13g2_fill_2 FILLER_14_2139 ();
 sg13g2_fill_1 FILLER_14_2141 ();
 sg13g2_fill_2 FILLER_14_2225 ();
 sg13g2_fill_1 FILLER_14_2227 ();
 sg13g2_decap_4 FILLER_14_2233 ();
 sg13g2_fill_1 FILLER_14_2253 ();
 sg13g2_fill_1 FILLER_14_2277 ();
 sg13g2_fill_1 FILLER_14_2327 ();
 sg13g2_fill_2 FILLER_14_2333 ();
 sg13g2_fill_2 FILLER_14_2365 ();
 sg13g2_fill_1 FILLER_14_2367 ();
 sg13g2_fill_2 FILLER_14_2420 ();
 sg13g2_decap_8 FILLER_14_2544 ();
 sg13g2_fill_2 FILLER_14_2555 ();
 sg13g2_fill_1 FILLER_14_2578 ();
 sg13g2_fill_1 FILLER_14_2604 ();
 sg13g2_fill_1 FILLER_14_2613 ();
 sg13g2_fill_2 FILLER_14_2666 ();
 sg13g2_fill_1 FILLER_14_2668 ();
 sg13g2_fill_1 FILLER_14_2710 ();
 sg13g2_fill_2 FILLER_14_2733 ();
 sg13g2_fill_1 FILLER_14_2773 ();
 sg13g2_fill_1 FILLER_14_2903 ();
 sg13g2_fill_1 FILLER_14_2913 ();
 sg13g2_fill_1 FILLER_14_2927 ();
 sg13g2_fill_2 FILLER_14_3001 ();
 sg13g2_fill_1 FILLER_14_3003 ();
 sg13g2_fill_2 FILLER_14_3059 ();
 sg13g2_decap_4 FILLER_14_3092 ();
 sg13g2_fill_2 FILLER_14_3150 ();
 sg13g2_decap_4 FILLER_14_3165 ();
 sg13g2_fill_1 FILLER_14_3169 ();
 sg13g2_fill_2 FILLER_14_3237 ();
 sg13g2_fill_1 FILLER_14_3264 ();
 sg13g2_fill_2 FILLER_14_3292 ();
 sg13g2_fill_1 FILLER_14_3294 ();
 sg13g2_fill_1 FILLER_14_3341 ();
 sg13g2_fill_2 FILLER_14_3360 ();
 sg13g2_fill_1 FILLER_14_3362 ();
 sg13g2_fill_1 FILLER_14_3438 ();
 sg13g2_fill_2 FILLER_14_3454 ();
 sg13g2_fill_1 FILLER_14_3456 ();
 sg13g2_decap_4 FILLER_14_3489 ();
 sg13g2_fill_1 FILLER_14_3493 ();
 sg13g2_decap_4 FILLER_14_3499 ();
 sg13g2_fill_1 FILLER_14_3520 ();
 sg13g2_fill_2 FILLER_14_3524 ();
 sg13g2_fill_1 FILLER_14_3567 ();
 sg13g2_fill_2 FILLER_14_3577 ();
 sg13g2_fill_1 FILLER_14_3579 ();
 sg13g2_fill_1 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_29 ();
 sg13g2_fill_2 FILLER_15_43 ();
 sg13g2_fill_2 FILLER_15_65 ();
 sg13g2_fill_2 FILLER_15_82 ();
 sg13g2_fill_1 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_107 ();
 sg13g2_decap_4 FILLER_15_114 ();
 sg13g2_decap_4 FILLER_15_121 ();
 sg13g2_fill_1 FILLER_15_125 ();
 sg13g2_fill_2 FILLER_15_139 ();
 sg13g2_fill_1 FILLER_15_141 ();
 sg13g2_decap_8 FILLER_15_146 ();
 sg13g2_fill_2 FILLER_15_237 ();
 sg13g2_fill_2 FILLER_15_258 ();
 sg13g2_fill_1 FILLER_15_300 ();
 sg13g2_fill_2 FILLER_15_335 ();
 sg13g2_fill_1 FILLER_15_337 ();
 sg13g2_decap_4 FILLER_15_369 ();
 sg13g2_fill_2 FILLER_15_440 ();
 sg13g2_fill_1 FILLER_15_442 ();
 sg13g2_fill_2 FILLER_15_509 ();
 sg13g2_fill_1 FILLER_15_511 ();
 sg13g2_fill_1 FILLER_15_538 ();
 sg13g2_fill_1 FILLER_15_569 ();
 sg13g2_fill_2 FILLER_15_579 ();
 sg13g2_fill_2 FILLER_15_593 ();
 sg13g2_fill_2 FILLER_15_608 ();
 sg13g2_fill_1 FILLER_15_610 ();
 sg13g2_fill_2 FILLER_15_633 ();
 sg13g2_fill_1 FILLER_15_648 ();
 sg13g2_fill_2 FILLER_15_671 ();
 sg13g2_fill_2 FILLER_15_724 ();
 sg13g2_fill_2 FILLER_15_753 ();
 sg13g2_fill_1 FILLER_15_755 ();
 sg13g2_fill_1 FILLER_15_766 ();
 sg13g2_fill_1 FILLER_15_783 ();
 sg13g2_fill_1 FILLER_15_825 ();
 sg13g2_decap_8 FILLER_15_870 ();
 sg13g2_decap_8 FILLER_15_877 ();
 sg13g2_fill_1 FILLER_15_884 ();
 sg13g2_decap_4 FILLER_15_894 ();
 sg13g2_fill_2 FILLER_15_919 ();
 sg13g2_fill_1 FILLER_15_925 ();
 sg13g2_decap_4 FILLER_15_939 ();
 sg13g2_fill_1 FILLER_15_943 ();
 sg13g2_fill_1 FILLER_15_948 ();
 sg13g2_fill_2 FILLER_15_959 ();
 sg13g2_fill_2 FILLER_15_969 ();
 sg13g2_fill_1 FILLER_15_998 ();
 sg13g2_fill_1 FILLER_15_1034 ();
 sg13g2_fill_2 FILLER_15_1074 ();
 sg13g2_fill_2 FILLER_15_1089 ();
 sg13g2_fill_2 FILLER_15_1132 ();
 sg13g2_fill_1 FILLER_15_1177 ();
 sg13g2_fill_1 FILLER_15_1184 ();
 sg13g2_fill_1 FILLER_15_1260 ();
 sg13g2_fill_1 FILLER_15_1475 ();
 sg13g2_fill_2 FILLER_15_1565 ();
 sg13g2_fill_2 FILLER_15_1626 ();
 sg13g2_fill_1 FILLER_15_1633 ();
 sg13g2_fill_2 FILLER_15_1765 ();
 sg13g2_decap_8 FILLER_15_1776 ();
 sg13g2_fill_1 FILLER_15_1783 ();
 sg13g2_decap_4 FILLER_15_1825 ();
 sg13g2_fill_2 FILLER_15_1870 ();
 sg13g2_fill_1 FILLER_15_1872 ();
 sg13g2_fill_2 FILLER_15_1878 ();
 sg13g2_fill_1 FILLER_15_1880 ();
 sg13g2_decap_4 FILLER_15_1909 ();
 sg13g2_fill_1 FILLER_15_1960 ();
 sg13g2_fill_2 FILLER_15_1976 ();
 sg13g2_fill_1 FILLER_15_2047 ();
 sg13g2_fill_1 FILLER_15_2057 ();
 sg13g2_fill_2 FILLER_15_2116 ();
 sg13g2_decap_4 FILLER_15_2142 ();
 sg13g2_fill_1 FILLER_15_2146 ();
 sg13g2_decap_4 FILLER_15_2151 ();
 sg13g2_fill_1 FILLER_15_2227 ();
 sg13g2_decap_4 FILLER_15_2241 ();
 sg13g2_decap_8 FILLER_15_2253 ();
 sg13g2_fill_1 FILLER_15_2260 ();
 sg13g2_fill_2 FILLER_15_2269 ();
 sg13g2_fill_2 FILLER_15_2287 ();
 sg13g2_fill_1 FILLER_15_2294 ();
 sg13g2_fill_2 FILLER_15_2303 ();
 sg13g2_fill_2 FILLER_15_2315 ();
 sg13g2_fill_1 FILLER_15_2317 ();
 sg13g2_fill_2 FILLER_15_2474 ();
 sg13g2_fill_1 FILLER_15_2476 ();
 sg13g2_decap_4 FILLER_15_2516 ();
 sg13g2_fill_2 FILLER_15_2520 ();
 sg13g2_fill_2 FILLER_15_2544 ();
 sg13g2_fill_2 FILLER_15_2583 ();
 sg13g2_fill_1 FILLER_15_2585 ();
 sg13g2_fill_1 FILLER_15_2599 ();
 sg13g2_decap_4 FILLER_15_2621 ();
 sg13g2_fill_2 FILLER_15_2633 ();
 sg13g2_fill_1 FILLER_15_2663 ();
 sg13g2_fill_1 FILLER_15_2682 ();
 sg13g2_fill_2 FILLER_15_2716 ();
 sg13g2_fill_1 FILLER_15_2718 ();
 sg13g2_fill_1 FILLER_15_2733 ();
 sg13g2_fill_2 FILLER_15_2756 ();
 sg13g2_fill_1 FILLER_15_2758 ();
 sg13g2_fill_1 FILLER_15_2800 ();
 sg13g2_fill_1 FILLER_15_2829 ();
 sg13g2_fill_2 FILLER_15_2853 ();
 sg13g2_fill_1 FILLER_15_2877 ();
 sg13g2_fill_1 FILLER_15_2918 ();
 sg13g2_fill_2 FILLER_15_2935 ();
 sg13g2_fill_1 FILLER_15_2937 ();
 sg13g2_fill_1 FILLER_15_2947 ();
 sg13g2_fill_1 FILLER_15_2957 ();
 sg13g2_fill_1 FILLER_15_3018 ();
 sg13g2_fill_1 FILLER_15_3032 ();
 sg13g2_fill_1 FILLER_15_3072 ();
 sg13g2_fill_2 FILLER_15_3105 ();
 sg13g2_fill_1 FILLER_15_3122 ();
 sg13g2_fill_2 FILLER_15_3136 ();
 sg13g2_fill_1 FILLER_15_3151 ();
 sg13g2_fill_2 FILLER_15_3204 ();
 sg13g2_fill_1 FILLER_15_3206 ();
 sg13g2_fill_1 FILLER_15_3252 ();
 sg13g2_fill_1 FILLER_15_3299 ();
 sg13g2_fill_2 FILLER_15_3347 ();
 sg13g2_fill_1 FILLER_15_3349 ();
 sg13g2_decap_4 FILLER_15_3360 ();
 sg13g2_fill_2 FILLER_15_3364 ();
 sg13g2_fill_1 FILLER_15_3435 ();
 sg13g2_fill_2 FILLER_15_3441 ();
 sg13g2_fill_1 FILLER_15_3461 ();
 sg13g2_fill_2 FILLER_15_3489 ();
 sg13g2_fill_2 FILLER_15_3529 ();
 sg13g2_decap_8 FILLER_15_3535 ();
 sg13g2_fill_2 FILLER_15_3542 ();
 sg13g2_fill_2 FILLER_15_3578 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_11 ();
 sg13g2_fill_2 FILLER_16_34 ();
 sg13g2_fill_1 FILLER_16_36 ();
 sg13g2_fill_2 FILLER_16_50 ();
 sg13g2_fill_2 FILLER_16_64 ();
 sg13g2_fill_1 FILLER_16_66 ();
 sg13g2_decap_8 FILLER_16_72 ();
 sg13g2_fill_1 FILLER_16_79 ();
 sg13g2_fill_2 FILLER_16_90 ();
 sg13g2_fill_1 FILLER_16_92 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_4 FILLER_16_112 ();
 sg13g2_fill_1 FILLER_16_144 ();
 sg13g2_fill_1 FILLER_16_166 ();
 sg13g2_fill_1 FILLER_16_206 ();
 sg13g2_fill_2 FILLER_16_217 ();
 sg13g2_fill_1 FILLER_16_219 ();
 sg13g2_fill_1 FILLER_16_280 ();
 sg13g2_fill_1 FILLER_16_376 ();
 sg13g2_fill_1 FILLER_16_451 ();
 sg13g2_fill_2 FILLER_16_520 ();
 sg13g2_fill_1 FILLER_16_522 ();
 sg13g2_fill_1 FILLER_16_602 ();
 sg13g2_decap_4 FILLER_16_644 ();
 sg13g2_fill_1 FILLER_16_648 ();
 sg13g2_fill_1 FILLER_16_721 ();
 sg13g2_fill_2 FILLER_16_781 ();
 sg13g2_fill_2 FILLER_16_873 ();
 sg13g2_fill_1 FILLER_16_875 ();
 sg13g2_fill_2 FILLER_16_889 ();
 sg13g2_fill_2 FILLER_16_919 ();
 sg13g2_fill_2 FILLER_16_1025 ();
 sg13g2_fill_1 FILLER_16_1027 ();
 sg13g2_fill_2 FILLER_16_1066 ();
 sg13g2_fill_2 FILLER_16_1087 ();
 sg13g2_fill_2 FILLER_16_1122 ();
 sg13g2_fill_1 FILLER_16_1124 ();
 sg13g2_fill_2 FILLER_16_1157 ();
 sg13g2_fill_1 FILLER_16_1159 ();
 sg13g2_fill_1 FILLER_16_1169 ();
 sg13g2_fill_2 FILLER_16_1189 ();
 sg13g2_fill_1 FILLER_16_1191 ();
 sg13g2_fill_2 FILLER_16_1205 ();
 sg13g2_fill_1 FILLER_16_1290 ();
 sg13g2_fill_2 FILLER_16_1331 ();
 sg13g2_fill_1 FILLER_16_1333 ();
 sg13g2_fill_2 FILLER_16_1338 ();
 sg13g2_fill_1 FILLER_16_1340 ();
 sg13g2_decap_4 FILLER_16_1354 ();
 sg13g2_decap_8 FILLER_16_1414 ();
 sg13g2_decap_4 FILLER_16_1430 ();
 sg13g2_fill_1 FILLER_16_1434 ();
 sg13g2_fill_1 FILLER_16_1489 ();
 sg13g2_fill_1 FILLER_16_1530 ();
 sg13g2_fill_2 FILLER_16_1550 ();
 sg13g2_fill_1 FILLER_16_1552 ();
 sg13g2_fill_1 FILLER_16_1601 ();
 sg13g2_fill_1 FILLER_16_1694 ();
 sg13g2_fill_2 FILLER_16_1724 ();
 sg13g2_fill_1 FILLER_16_1726 ();
 sg13g2_fill_1 FILLER_16_1765 ();
 sg13g2_decap_4 FILLER_16_1793 ();
 sg13g2_fill_1 FILLER_16_1797 ();
 sg13g2_fill_2 FILLER_16_1833 ();
 sg13g2_fill_1 FILLER_16_1835 ();
 sg13g2_fill_2 FILLER_16_1840 ();
 sg13g2_fill_2 FILLER_16_1859 ();
 sg13g2_fill_1 FILLER_16_1861 ();
 sg13g2_fill_1 FILLER_16_1881 ();
 sg13g2_fill_2 FILLER_16_1945 ();
 sg13g2_fill_1 FILLER_16_1947 ();
 sg13g2_fill_1 FILLER_16_1987 ();
 sg13g2_fill_2 FILLER_16_2056 ();
 sg13g2_fill_1 FILLER_16_2058 ();
 sg13g2_fill_1 FILLER_16_2068 ();
 sg13g2_fill_2 FILLER_16_2090 ();
 sg13g2_fill_1 FILLER_16_2121 ();
 sg13g2_decap_4 FILLER_16_2168 ();
 sg13g2_fill_2 FILLER_16_2187 ();
 sg13g2_fill_1 FILLER_16_2189 ();
 sg13g2_decap_8 FILLER_16_2200 ();
 sg13g2_fill_2 FILLER_16_2207 ();
 sg13g2_fill_1 FILLER_16_2209 ();
 sg13g2_decap_8 FILLER_16_2223 ();
 sg13g2_fill_2 FILLER_16_2264 ();
 sg13g2_fill_1 FILLER_16_2266 ();
 sg13g2_decap_4 FILLER_16_2328 ();
 sg13g2_fill_2 FILLER_16_2332 ();
 sg13g2_fill_1 FILLER_16_2365 ();
 sg13g2_fill_2 FILLER_16_2402 ();
 sg13g2_fill_1 FILLER_16_2404 ();
 sg13g2_fill_2 FILLER_16_2433 ();
 sg13g2_fill_1 FILLER_16_2435 ();
 sg13g2_fill_2 FILLER_16_2457 ();
 sg13g2_fill_2 FILLER_16_2492 ();
 sg13g2_fill_1 FILLER_16_2494 ();
 sg13g2_decap_8 FILLER_16_2580 ();
 sg13g2_decap_8 FILLER_16_2622 ();
 sg13g2_fill_2 FILLER_16_2679 ();
 sg13g2_fill_1 FILLER_16_2681 ();
 sg13g2_fill_1 FILLER_16_2705 ();
 sg13g2_fill_2 FILLER_16_2715 ();
 sg13g2_fill_2 FILLER_16_2745 ();
 sg13g2_fill_2 FILLER_16_2784 ();
 sg13g2_fill_2 FILLER_16_2799 ();
 sg13g2_fill_1 FILLER_16_2819 ();
 sg13g2_fill_2 FILLER_16_2890 ();
 sg13g2_fill_1 FILLER_16_2900 ();
 sg13g2_fill_1 FILLER_16_2918 ();
 sg13g2_fill_1 FILLER_16_2944 ();
 sg13g2_fill_1 FILLER_16_2973 ();
 sg13g2_fill_2 FILLER_16_3069 ();
 sg13g2_fill_2 FILLER_16_3126 ();
 sg13g2_fill_2 FILLER_16_3202 ();
 sg13g2_fill_2 FILLER_16_3257 ();
 sg13g2_fill_2 FILLER_16_3357 ();
 sg13g2_fill_2 FILLER_16_3472 ();
 sg13g2_decap_8 FILLER_16_3506 ();
 sg13g2_decap_4 FILLER_16_3513 ();
 sg13g2_fill_1 FILLER_16_3517 ();
 sg13g2_fill_1 FILLER_16_3542 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_43 ();
 sg13g2_fill_1 FILLER_17_47 ();
 sg13g2_decap_8 FILLER_17_57 ();
 sg13g2_fill_2 FILLER_17_77 ();
 sg13g2_decap_4 FILLER_17_84 ();
 sg13g2_fill_2 FILLER_17_88 ();
 sg13g2_decap_4 FILLER_17_94 ();
 sg13g2_fill_1 FILLER_17_155 ();
 sg13g2_fill_2 FILLER_17_161 ();
 sg13g2_fill_2 FILLER_17_247 ();
 sg13g2_fill_2 FILLER_17_270 ();
 sg13g2_fill_1 FILLER_17_272 ();
 sg13g2_fill_2 FILLER_17_286 ();
 sg13g2_fill_2 FILLER_17_330 ();
 sg13g2_fill_2 FILLER_17_347 ();
 sg13g2_fill_1 FILLER_17_349 ();
 sg13g2_fill_1 FILLER_17_364 ();
 sg13g2_fill_2 FILLER_17_384 ();
 sg13g2_fill_2 FILLER_17_399 ();
 sg13g2_fill_1 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_415 ();
 sg13g2_fill_2 FILLER_17_479 ();
 sg13g2_fill_2 FILLER_17_500 ();
 sg13g2_fill_1 FILLER_17_502 ();
 sg13g2_fill_1 FILLER_17_571 ();
 sg13g2_decap_8 FILLER_17_636 ();
 sg13g2_fill_2 FILLER_17_652 ();
 sg13g2_fill_1 FILLER_17_654 ();
 sg13g2_fill_1 FILLER_17_685 ();
 sg13g2_fill_2 FILLER_17_740 ();
 sg13g2_fill_1 FILLER_17_760 ();
 sg13g2_fill_2 FILLER_17_785 ();
 sg13g2_fill_1 FILLER_17_787 ();
 sg13g2_fill_2 FILLER_17_797 ();
 sg13g2_fill_1 FILLER_17_799 ();
 sg13g2_fill_1 FILLER_17_826 ();
 sg13g2_fill_2 FILLER_17_905 ();
 sg13g2_fill_1 FILLER_17_907 ();
 sg13g2_decap_8 FILLER_17_933 ();
 sg13g2_decap_8 FILLER_17_940 ();
 sg13g2_fill_1 FILLER_17_1020 ();
 sg13g2_fill_1 FILLER_17_1032 ();
 sg13g2_fill_1 FILLER_17_1073 ();
 sg13g2_fill_2 FILLER_17_1091 ();
 sg13g2_fill_1 FILLER_17_1093 ();
 sg13g2_fill_1 FILLER_17_1121 ();
 sg13g2_fill_2 FILLER_17_1150 ();
 sg13g2_fill_1 FILLER_17_1152 ();
 sg13g2_fill_2 FILLER_17_1232 ();
 sg13g2_fill_2 FILLER_17_1330 ();
 sg13g2_fill_1 FILLER_17_1332 ();
 sg13g2_fill_2 FILLER_17_1371 ();
 sg13g2_fill_1 FILLER_17_1401 ();
 sg13g2_decap_8 FILLER_17_1435 ();
 sg13g2_fill_2 FILLER_17_1442 ();
 sg13g2_fill_2 FILLER_17_1579 ();
 sg13g2_fill_2 FILLER_17_1617 ();
 sg13g2_fill_2 FILLER_17_1641 ();
 sg13g2_fill_2 FILLER_17_1734 ();
 sg13g2_fill_1 FILLER_17_1736 ();
 sg13g2_fill_2 FILLER_17_1751 ();
 sg13g2_fill_1 FILLER_17_1764 ();
 sg13g2_fill_2 FILLER_17_1770 ();
 sg13g2_decap_4 FILLER_17_1790 ();
 sg13g2_fill_1 FILLER_17_1794 ();
 sg13g2_fill_1 FILLER_17_1852 ();
 sg13g2_fill_2 FILLER_17_1866 ();
 sg13g2_fill_2 FILLER_17_1930 ();
 sg13g2_fill_2 FILLER_17_1968 ();
 sg13g2_fill_2 FILLER_17_2018 ();
 sg13g2_fill_2 FILLER_17_2098 ();
 sg13g2_decap_4 FILLER_17_2123 ();
 sg13g2_fill_2 FILLER_17_2127 ();
 sg13g2_fill_1 FILLER_17_2146 ();
 sg13g2_fill_2 FILLER_17_2165 ();
 sg13g2_fill_2 FILLER_17_2182 ();
 sg13g2_fill_1 FILLER_17_2184 ();
 sg13g2_decap_4 FILLER_17_2193 ();
 sg13g2_fill_2 FILLER_17_2205 ();
 sg13g2_fill_1 FILLER_17_2207 ();
 sg13g2_fill_1 FILLER_17_2236 ();
 sg13g2_fill_1 FILLER_17_2258 ();
 sg13g2_fill_1 FILLER_17_2273 ();
 sg13g2_decap_8 FILLER_17_2335 ();
 sg13g2_decap_4 FILLER_17_2342 ();
 sg13g2_fill_1 FILLER_17_2346 ();
 sg13g2_fill_2 FILLER_17_2380 ();
 sg13g2_fill_1 FILLER_17_2382 ();
 sg13g2_fill_1 FILLER_17_2392 ();
 sg13g2_fill_1 FILLER_17_2439 ();
 sg13g2_fill_2 FILLER_17_2477 ();
 sg13g2_fill_2 FILLER_17_2534 ();
 sg13g2_fill_1 FILLER_17_2536 ();
 sg13g2_fill_1 FILLER_17_2587 ();
 sg13g2_fill_1 FILLER_17_2591 ();
 sg13g2_fill_1 FILLER_17_2618 ();
 sg13g2_fill_2 FILLER_17_2652 ();
 sg13g2_fill_1 FILLER_17_2654 ();
 sg13g2_fill_1 FILLER_17_2668 ();
 sg13g2_fill_2 FILLER_17_2734 ();
 sg13g2_fill_1 FILLER_17_2813 ();
 sg13g2_fill_2 FILLER_17_2852 ();
 sg13g2_fill_1 FILLER_17_2854 ();
 sg13g2_fill_2 FILLER_17_2896 ();
 sg13g2_fill_1 FILLER_17_2898 ();
 sg13g2_decap_4 FILLER_17_2932 ();
 sg13g2_fill_2 FILLER_17_2936 ();
 sg13g2_fill_2 FILLER_17_2951 ();
 sg13g2_fill_2 FILLER_17_3023 ();
 sg13g2_fill_1 FILLER_17_3025 ();
 sg13g2_fill_2 FILLER_17_3068 ();
 sg13g2_fill_1 FILLER_17_3070 ();
 sg13g2_fill_1 FILLER_17_3075 ();
 sg13g2_fill_2 FILLER_17_3080 ();
 sg13g2_fill_1 FILLER_17_3082 ();
 sg13g2_fill_2 FILLER_17_3101 ();
 sg13g2_fill_2 FILLER_17_3287 ();
 sg13g2_fill_1 FILLER_17_3289 ();
 sg13g2_fill_2 FILLER_17_3349 ();
 sg13g2_fill_1 FILLER_17_3351 ();
 sg13g2_fill_1 FILLER_17_3407 ();
 sg13g2_fill_2 FILLER_17_3428 ();
 sg13g2_fill_2 FILLER_17_3439 ();
 sg13g2_decap_4 FILLER_17_3450 ();
 sg13g2_fill_1 FILLER_17_3454 ();
 sg13g2_fill_2 FILLER_17_3459 ();
 sg13g2_fill_1 FILLER_17_3461 ();
 sg13g2_fill_1 FILLER_17_3466 ();
 sg13g2_fill_2 FILLER_17_3481 ();
 sg13g2_fill_1 FILLER_17_3483 ();
 sg13g2_decap_8 FILLER_17_3509 ();
 sg13g2_decap_8 FILLER_17_3536 ();
 sg13g2_fill_1 FILLER_17_3543 ();
 sg13g2_fill_2 FILLER_17_3561 ();
 sg13g2_fill_1 FILLER_17_3563 ();
 sg13g2_fill_2 FILLER_17_3577 ();
 sg13g2_fill_1 FILLER_17_3579 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_22 ();
 sg13g2_fill_2 FILLER_18_28 ();
 sg13g2_fill_2 FILLER_18_35 ();
 sg13g2_fill_2 FILLER_18_49 ();
 sg13g2_fill_1 FILLER_18_75 ();
 sg13g2_fill_2 FILLER_18_116 ();
 sg13g2_decap_4 FILLER_18_126 ();
 sg13g2_fill_2 FILLER_18_130 ();
 sg13g2_fill_1 FILLER_18_142 ();
 sg13g2_fill_1 FILLER_18_169 ();
 sg13g2_fill_2 FILLER_18_217 ();
 sg13g2_fill_1 FILLER_18_259 ();
 sg13g2_fill_1 FILLER_18_340 ();
 sg13g2_fill_1 FILLER_18_369 ();
 sg13g2_fill_1 FILLER_18_415 ();
 sg13g2_fill_2 FILLER_18_426 ();
 sg13g2_fill_1 FILLER_18_460 ();
 sg13g2_fill_1 FILLER_18_470 ();
 sg13g2_fill_1 FILLER_18_508 ();
 sg13g2_fill_1 FILLER_18_522 ();
 sg13g2_fill_1 FILLER_18_536 ();
 sg13g2_fill_1 FILLER_18_583 ();
 sg13g2_fill_1 FILLER_18_610 ();
 sg13g2_fill_1 FILLER_18_657 ();
 sg13g2_fill_2 FILLER_18_695 ();
 sg13g2_fill_2 FILLER_18_713 ();
 sg13g2_fill_1 FILLER_18_715 ();
 sg13g2_fill_2 FILLER_18_754 ();
 sg13g2_fill_1 FILLER_18_756 ();
 sg13g2_fill_2 FILLER_18_855 ();
 sg13g2_fill_1 FILLER_18_887 ();
 sg13g2_fill_1 FILLER_18_906 ();
 sg13g2_decap_8 FILLER_18_940 ();
 sg13g2_decap_8 FILLER_18_960 ();
 sg13g2_fill_2 FILLER_18_967 ();
 sg13g2_fill_1 FILLER_18_982 ();
 sg13g2_fill_2 FILLER_18_1111 ();
 sg13g2_fill_1 FILLER_18_1113 ();
 sg13g2_fill_2 FILLER_18_1183 ();
 sg13g2_fill_1 FILLER_18_1185 ();
 sg13g2_fill_1 FILLER_18_1244 ();
 sg13g2_fill_1 FILLER_18_1284 ();
 sg13g2_fill_2 FILLER_18_1315 ();
 sg13g2_decap_8 FILLER_18_1325 ();
 sg13g2_fill_1 FILLER_18_1345 ();
 sg13g2_fill_1 FILLER_18_1361 ();
 sg13g2_fill_2 FILLER_18_1386 ();
 sg13g2_fill_1 FILLER_18_1388 ();
 sg13g2_fill_1 FILLER_18_1415 ();
 sg13g2_fill_1 FILLER_18_1429 ();
 sg13g2_fill_1 FILLER_18_1463 ();
 sg13g2_fill_2 FILLER_18_1515 ();
 sg13g2_fill_1 FILLER_18_1517 ();
 sg13g2_fill_2 FILLER_18_1534 ();
 sg13g2_fill_2 FILLER_18_1549 ();
 sg13g2_fill_1 FILLER_18_1551 ();
 sg13g2_fill_2 FILLER_18_1606 ();
 sg13g2_fill_1 FILLER_18_1608 ();
 sg13g2_fill_1 FILLER_18_1615 ();
 sg13g2_fill_1 FILLER_18_1630 ();
 sg13g2_fill_2 FILLER_18_1698 ();
 sg13g2_fill_1 FILLER_18_1700 ();
 sg13g2_fill_2 FILLER_18_1765 ();
 sg13g2_decap_8 FILLER_18_1795 ();
 sg13g2_fill_1 FILLER_18_1802 ();
 sg13g2_fill_2 FILLER_18_1834 ();
 sg13g2_decap_4 FILLER_18_1849 ();
 sg13g2_fill_1 FILLER_18_1853 ();
 sg13g2_fill_2 FILLER_18_1885 ();
 sg13g2_fill_1 FILLER_18_1887 ();
 sg13g2_fill_1 FILLER_18_1933 ();
 sg13g2_fill_2 FILLER_18_2030 ();
 sg13g2_fill_2 FILLER_18_2056 ();
 sg13g2_fill_2 FILLER_18_2087 ();
 sg13g2_decap_4 FILLER_18_2121 ();
 sg13g2_fill_1 FILLER_18_2125 ();
 sg13g2_fill_2 FILLER_18_2138 ();
 sg13g2_fill_1 FILLER_18_2166 ();
 sg13g2_fill_2 FILLER_18_2194 ();
 sg13g2_fill_1 FILLER_18_2196 ();
 sg13g2_decap_4 FILLER_18_2221 ();
 sg13g2_fill_2 FILLER_18_2225 ();
 sg13g2_decap_8 FILLER_18_2287 ();
 sg13g2_decap_4 FILLER_18_2294 ();
 sg13g2_fill_1 FILLER_18_2298 ();
 sg13g2_fill_1 FILLER_18_2330 ();
 sg13g2_fill_2 FILLER_18_2361 ();
 sg13g2_fill_2 FILLER_18_2376 ();
 sg13g2_fill_2 FILLER_18_2450 ();
 sg13g2_fill_1 FILLER_18_2452 ();
 sg13g2_decap_8 FILLER_18_2516 ();
 sg13g2_fill_2 FILLER_18_2551 ();
 sg13g2_fill_1 FILLER_18_2580 ();
 sg13g2_fill_2 FILLER_18_2586 ();
 sg13g2_fill_2 FILLER_18_2597 ();
 sg13g2_fill_2 FILLER_18_2612 ();
 sg13g2_fill_1 FILLER_18_2614 ();
 sg13g2_fill_2 FILLER_18_2633 ();
 sg13g2_fill_2 FILLER_18_2657 ();
 sg13g2_fill_1 FILLER_18_2659 ();
 sg13g2_fill_2 FILLER_18_2669 ();
 sg13g2_fill_1 FILLER_18_2680 ();
 sg13g2_fill_1 FILLER_18_2709 ();
 sg13g2_fill_1 FILLER_18_2715 ();
 sg13g2_fill_2 FILLER_18_2728 ();
 sg13g2_fill_1 FILLER_18_2758 ();
 sg13g2_fill_2 FILLER_18_2787 ();
 sg13g2_fill_1 FILLER_18_2807 ();
 sg13g2_fill_1 FILLER_18_2830 ();
 sg13g2_decap_4 FILLER_18_2840 ();
 sg13g2_fill_1 FILLER_18_2844 ();
 sg13g2_fill_2 FILLER_18_2879 ();
 sg13g2_fill_1 FILLER_18_2940 ();
 sg13g2_fill_2 FILLER_18_3063 ();
 sg13g2_fill_2 FILLER_18_3162 ();
 sg13g2_fill_1 FILLER_18_3241 ();
 sg13g2_decap_4 FILLER_18_3372 ();
 sg13g2_fill_1 FILLER_18_3484 ();
 sg13g2_decap_4 FILLER_18_3490 ();
 sg13g2_fill_2 FILLER_18_3511 ();
 sg13g2_fill_1 FILLER_18_3513 ();
 sg13g2_decap_4 FILLER_18_3539 ();
 sg13g2_fill_1 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_44 ();
 sg13g2_fill_1 FILLER_19_46 ();
 sg13g2_decap_4 FILLER_19_94 ();
 sg13g2_fill_1 FILLER_19_98 ();
 sg13g2_fill_1 FILLER_19_104 ();
 sg13g2_fill_1 FILLER_19_141 ();
 sg13g2_fill_1 FILLER_19_150 ();
 sg13g2_fill_1 FILLER_19_160 ();
 sg13g2_fill_1 FILLER_19_229 ();
 sg13g2_fill_1 FILLER_19_312 ();
 sg13g2_fill_1 FILLER_19_331 ();
 sg13g2_decap_4 FILLER_19_389 ();
 sg13g2_fill_2 FILLER_19_469 ();
 sg13g2_decap_4 FILLER_19_488 ();
 sg13g2_fill_2 FILLER_19_492 ();
 sg13g2_fill_2 FILLER_19_503 ();
 sg13g2_fill_2 FILLER_19_550 ();
 sg13g2_fill_1 FILLER_19_552 ();
 sg13g2_fill_1 FILLER_19_593 ();
 sg13g2_fill_2 FILLER_19_635 ();
 sg13g2_fill_1 FILLER_19_637 ();
 sg13g2_fill_1 FILLER_19_666 ();
 sg13g2_fill_2 FILLER_19_705 ();
 sg13g2_fill_2 FILLER_19_734 ();
 sg13g2_fill_1 FILLER_19_777 ();
 sg13g2_fill_2 FILLER_19_788 ();
 sg13g2_fill_1 FILLER_19_790 ();
 sg13g2_fill_1 FILLER_19_823 ();
 sg13g2_fill_1 FILLER_19_851 ();
 sg13g2_decap_4 FILLER_19_920 ();
 sg13g2_fill_1 FILLER_19_1000 ();
 sg13g2_fill_1 FILLER_19_1017 ();
 sg13g2_fill_2 FILLER_19_1048 ();
 sg13g2_fill_1 FILLER_19_1138 ();
 sg13g2_fill_2 FILLER_19_1188 ();
 sg13g2_fill_2 FILLER_19_1230 ();
 sg13g2_fill_2 FILLER_19_1246 ();
 sg13g2_fill_1 FILLER_19_1248 ();
 sg13g2_fill_2 FILLER_19_1299 ();
 sg13g2_fill_1 FILLER_19_1314 ();
 sg13g2_fill_2 FILLER_19_1372 ();
 sg13g2_fill_2 FILLER_19_1400 ();
 sg13g2_fill_1 FILLER_19_1438 ();
 sg13g2_fill_2 FILLER_19_1467 ();
 sg13g2_fill_2 FILLER_19_1524 ();
 sg13g2_fill_2 FILLER_19_1554 ();
 sg13g2_fill_1 FILLER_19_1556 ();
 sg13g2_decap_4 FILLER_19_1583 ();
 sg13g2_fill_2 FILLER_19_1587 ();
 sg13g2_fill_1 FILLER_19_1608 ();
 sg13g2_fill_2 FILLER_19_1646 ();
 sg13g2_fill_2 FILLER_19_1652 ();
 sg13g2_fill_2 FILLER_19_1688 ();
 sg13g2_fill_2 FILLER_19_1712 ();
 sg13g2_decap_4 FILLER_19_1745 ();
 sg13g2_fill_2 FILLER_19_1749 ();
 sg13g2_fill_2 FILLER_19_1761 ();
 sg13g2_fill_2 FILLER_19_1776 ();
 sg13g2_fill_1 FILLER_19_1778 ();
 sg13g2_fill_1 FILLER_19_1834 ();
 sg13g2_decap_8 FILLER_19_1941 ();
 sg13g2_decap_4 FILLER_19_1948 ();
 sg13g2_fill_1 FILLER_19_1952 ();
 sg13g2_fill_2 FILLER_19_1979 ();
 sg13g2_fill_2 FILLER_19_1994 ();
 sg13g2_fill_1 FILLER_19_1996 ();
 sg13g2_fill_2 FILLER_19_2048 ();
 sg13g2_fill_1 FILLER_19_2059 ();
 sg13g2_fill_2 FILLER_19_2075 ();
 sg13g2_fill_1 FILLER_19_2077 ();
 sg13g2_fill_2 FILLER_19_2083 ();
 sg13g2_fill_1 FILLER_19_2085 ();
 sg13g2_fill_2 FILLER_19_2094 ();
 sg13g2_fill_1 FILLER_19_2101 ();
 sg13g2_decap_8 FILLER_19_2119 ();
 sg13g2_fill_1 FILLER_19_2139 ();
 sg13g2_fill_1 FILLER_19_2148 ();
 sg13g2_decap_4 FILLER_19_2162 ();
 sg13g2_fill_1 FILLER_19_2166 ();
 sg13g2_fill_2 FILLER_19_2172 ();
 sg13g2_fill_1 FILLER_19_2174 ();
 sg13g2_fill_1 FILLER_19_2216 ();
 sg13g2_fill_1 FILLER_19_2244 ();
 sg13g2_fill_1 FILLER_19_2254 ();
 sg13g2_decap_4 FILLER_19_2285 ();
 sg13g2_fill_2 FILLER_19_2289 ();
 sg13g2_fill_2 FILLER_19_2310 ();
 sg13g2_fill_2 FILLER_19_2320 ();
 sg13g2_fill_1 FILLER_19_2322 ();
 sg13g2_decap_4 FILLER_19_2358 ();
 sg13g2_fill_1 FILLER_19_2388 ();
 sg13g2_fill_1 FILLER_19_2397 ();
 sg13g2_fill_2 FILLER_19_2448 ();
 sg13g2_fill_2 FILLER_19_2460 ();
 sg13g2_fill_2 FILLER_19_2484 ();
 sg13g2_fill_2 FILLER_19_2527 ();
 sg13g2_fill_1 FILLER_19_2529 ();
 sg13g2_decap_8 FILLER_19_2594 ();
 sg13g2_fill_2 FILLER_19_2601 ();
 sg13g2_fill_1 FILLER_19_2603 ();
 sg13g2_fill_2 FILLER_19_2616 ();
 sg13g2_decap_4 FILLER_19_2622 ();
 sg13g2_fill_2 FILLER_19_2626 ();
 sg13g2_fill_2 FILLER_19_2659 ();
 sg13g2_fill_1 FILLER_19_2661 ();
 sg13g2_fill_1 FILLER_19_2672 ();
 sg13g2_fill_2 FILLER_19_2728 ();
 sg13g2_fill_2 FILLER_19_2748 ();
 sg13g2_fill_1 FILLER_19_2750 ();
 sg13g2_fill_2 FILLER_19_2760 ();
 sg13g2_fill_2 FILLER_19_2771 ();
 sg13g2_fill_1 FILLER_19_2798 ();
 sg13g2_decap_8 FILLER_19_2827 ();
 sg13g2_decap_4 FILLER_19_2834 ();
 sg13g2_decap_4 FILLER_19_2875 ();
 sg13g2_fill_1 FILLER_19_2879 ();
 sg13g2_fill_2 FILLER_19_2908 ();
 sg13g2_fill_1 FILLER_19_2910 ();
 sg13g2_fill_1 FILLER_19_2920 ();
 sg13g2_fill_1 FILLER_19_2930 ();
 sg13g2_fill_1 FILLER_19_2994 ();
 sg13g2_fill_1 FILLER_19_3027 ();
 sg13g2_fill_2 FILLER_19_3041 ();
 sg13g2_fill_1 FILLER_19_3043 ();
 sg13g2_fill_1 FILLER_19_3057 ();
 sg13g2_fill_2 FILLER_19_3087 ();
 sg13g2_fill_2 FILLER_19_3111 ();
 sg13g2_fill_2 FILLER_19_3145 ();
 sg13g2_fill_2 FILLER_19_3173 ();
 sg13g2_fill_2 FILLER_19_3196 ();
 sg13g2_fill_1 FILLER_19_3253 ();
 sg13g2_fill_2 FILLER_19_3330 ();
 sg13g2_fill_2 FILLER_19_3373 ();
 sg13g2_fill_1 FILLER_19_3375 ();
 sg13g2_decap_8 FILLER_19_3441 ();
 sg13g2_fill_1 FILLER_19_3448 ();
 sg13g2_decap_4 FILLER_19_3466 ();
 sg13g2_fill_1 FILLER_19_3518 ();
 sg13g2_decap_4 FILLER_19_3533 ();
 sg13g2_fill_2 FILLER_19_3537 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_4 ();
 sg13g2_decap_8 FILLER_20_10 ();
 sg13g2_fill_1 FILLER_20_17 ();
 sg13g2_fill_2 FILLER_20_47 ();
 sg13g2_fill_1 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_68 ();
 sg13g2_decap_4 FILLER_20_94 ();
 sg13g2_fill_2 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_104 ();
 sg13g2_fill_1 FILLER_20_111 ();
 sg13g2_fill_2 FILLER_20_180 ();
 sg13g2_fill_1 FILLER_20_182 ();
 sg13g2_fill_1 FILLER_20_192 ();
 sg13g2_fill_1 FILLER_20_216 ();
 sg13g2_fill_2 FILLER_20_236 ();
 sg13g2_fill_1 FILLER_20_313 ();
 sg13g2_fill_2 FILLER_20_342 ();
 sg13g2_fill_1 FILLER_20_344 ();
 sg13g2_fill_1 FILLER_20_414 ();
 sg13g2_fill_1 FILLER_20_482 ();
 sg13g2_fill_2 FILLER_20_500 ();
 sg13g2_fill_1 FILLER_20_502 ();
 sg13g2_fill_1 FILLER_20_532 ();
 sg13g2_fill_1 FILLER_20_542 ();
 sg13g2_fill_2 FILLER_20_564 ();
 sg13g2_fill_2 FILLER_20_609 ();
 sg13g2_fill_2 FILLER_20_634 ();
 sg13g2_decap_8 FILLER_20_650 ();
 sg13g2_fill_1 FILLER_20_657 ();
 sg13g2_fill_2 FILLER_20_686 ();
 sg13g2_fill_1 FILLER_20_697 ();
 sg13g2_fill_1 FILLER_20_753 ();
 sg13g2_fill_1 FILLER_20_781 ();
 sg13g2_fill_1 FILLER_20_802 ();
 sg13g2_fill_1 FILLER_20_853 ();
 sg13g2_fill_1 FILLER_20_862 ();
 sg13g2_fill_1 FILLER_20_912 ();
 sg13g2_fill_2 FILLER_20_926 ();
 sg13g2_fill_1 FILLER_20_928 ();
 sg13g2_decap_4 FILLER_20_955 ();
 sg13g2_decap_4 FILLER_20_981 ();
 sg13g2_fill_2 FILLER_20_1065 ();
 sg13g2_fill_2 FILLER_20_1137 ();
 sg13g2_fill_2 FILLER_20_1185 ();
 sg13g2_fill_2 FILLER_20_1254 ();
 sg13g2_decap_4 FILLER_20_1301 ();
 sg13g2_fill_1 FILLER_20_1351 ();
 sg13g2_fill_2 FILLER_20_1409 ();
 sg13g2_fill_2 FILLER_20_1451 ();
 sg13g2_fill_1 FILLER_20_1453 ();
 sg13g2_fill_2 FILLER_20_1492 ();
 sg13g2_fill_1 FILLER_20_1512 ();
 sg13g2_fill_2 FILLER_20_1537 ();
 sg13g2_fill_2 FILLER_20_1569 ();
 sg13g2_decap_4 FILLER_20_1638 ();
 sg13g2_fill_2 FILLER_20_1642 ();
 sg13g2_fill_2 FILLER_20_1653 ();
 sg13g2_fill_1 FILLER_20_1668 ();
 sg13g2_fill_1 FILLER_20_1682 ();
 sg13g2_fill_2 FILLER_20_1701 ();
 sg13g2_fill_2 FILLER_20_1711 ();
 sg13g2_fill_2 FILLER_20_1725 ();
 sg13g2_fill_1 FILLER_20_1727 ();
 sg13g2_fill_2 FILLER_20_1752 ();
 sg13g2_fill_1 FILLER_20_1754 ();
 sg13g2_decap_4 FILLER_20_1798 ();
 sg13g2_fill_2 FILLER_20_1802 ();
 sg13g2_decap_4 FILLER_20_1837 ();
 sg13g2_fill_1 FILLER_20_1841 ();
 sg13g2_fill_1 FILLER_20_1850 ();
 sg13g2_fill_1 FILLER_20_1863 ();
 sg13g2_fill_2 FILLER_20_1899 ();
 sg13g2_fill_1 FILLER_20_1901 ();
 sg13g2_decap_4 FILLER_20_1918 ();
 sg13g2_fill_1 FILLER_20_1922 ();
 sg13g2_decap_8 FILLER_20_1939 ();
 sg13g2_fill_2 FILLER_20_1946 ();
 sg13g2_fill_1 FILLER_20_1998 ();
 sg13g2_fill_2 FILLER_20_2012 ();
 sg13g2_fill_1 FILLER_20_2014 ();
 sg13g2_fill_1 FILLER_20_2024 ();
 sg13g2_fill_2 FILLER_20_2049 ();
 sg13g2_fill_2 FILLER_20_2073 ();
 sg13g2_fill_2 FILLER_20_2090 ();
 sg13g2_fill_1 FILLER_20_2092 ();
 sg13g2_decap_4 FILLER_20_2100 ();
 sg13g2_fill_2 FILLER_20_2130 ();
 sg13g2_fill_2 FILLER_20_2147 ();
 sg13g2_fill_1 FILLER_20_2149 ();
 sg13g2_decap_4 FILLER_20_2160 ();
 sg13g2_decap_8 FILLER_20_2188 ();
 sg13g2_decap_4 FILLER_20_2195 ();
 sg13g2_fill_2 FILLER_20_2209 ();
 sg13g2_decap_8 FILLER_20_2219 ();
 sg13g2_fill_2 FILLER_20_2226 ();
 sg13g2_fill_2 FILLER_20_2277 ();
 sg13g2_fill_2 FILLER_20_2300 ();
 sg13g2_fill_1 FILLER_20_2356 ();
 sg13g2_fill_2 FILLER_20_2365 ();
 sg13g2_fill_1 FILLER_20_2367 ();
 sg13g2_fill_1 FILLER_20_2373 ();
 sg13g2_fill_2 FILLER_20_2397 ();
 sg13g2_decap_8 FILLER_20_2407 ();
 sg13g2_fill_2 FILLER_20_2414 ();
 sg13g2_decap_4 FILLER_20_2421 ();
 sg13g2_fill_1 FILLER_20_2425 ();
 sg13g2_fill_2 FILLER_20_2444 ();
 sg13g2_decap_4 FILLER_20_2479 ();
 sg13g2_fill_2 FILLER_20_2496 ();
 sg13g2_fill_1 FILLER_20_2498 ();
 sg13g2_fill_1 FILLER_20_2540 ();
 sg13g2_decap_4 FILLER_20_2562 ();
 sg13g2_fill_2 FILLER_20_2588 ();
 sg13g2_fill_1 FILLER_20_2590 ();
 sg13g2_decap_8 FILLER_20_2623 ();
 sg13g2_fill_2 FILLER_20_2630 ();
 sg13g2_fill_1 FILLER_20_2632 ();
 sg13g2_fill_2 FILLER_20_2651 ();
 sg13g2_fill_1 FILLER_20_2670 ();
 sg13g2_fill_1 FILLER_20_2703 ();
 sg13g2_decap_8 FILLER_20_2725 ();
 sg13g2_decap_8 FILLER_20_2748 ();
 sg13g2_fill_2 FILLER_20_2811 ();
 sg13g2_decap_4 FILLER_20_2830 ();
 sg13g2_fill_1 FILLER_20_2922 ();
 sg13g2_fill_2 FILLER_20_2931 ();
 sg13g2_fill_1 FILLER_20_2933 ();
 sg13g2_fill_1 FILLER_20_2947 ();
 sg13g2_fill_2 FILLER_20_2957 ();
 sg13g2_fill_1 FILLER_20_2959 ();
 sg13g2_fill_2 FILLER_20_2970 ();
 sg13g2_fill_1 FILLER_20_2972 ();
 sg13g2_fill_2 FILLER_20_2981 ();
 sg13g2_fill_2 FILLER_20_3024 ();
 sg13g2_fill_1 FILLER_20_3039 ();
 sg13g2_fill_1 FILLER_20_3045 ();
 sg13g2_decap_4 FILLER_20_3074 ();
 sg13g2_decap_8 FILLER_20_3091 ();
 sg13g2_fill_2 FILLER_20_3115 ();
 sg13g2_fill_1 FILLER_20_3117 ();
 sg13g2_fill_1 FILLER_20_3136 ();
 sg13g2_fill_2 FILLER_20_3152 ();
 sg13g2_fill_1 FILLER_20_3154 ();
 sg13g2_fill_2 FILLER_20_3168 ();
 sg13g2_fill_2 FILLER_20_3183 ();
 sg13g2_fill_2 FILLER_20_3222 ();
 sg13g2_fill_1 FILLER_20_3224 ();
 sg13g2_fill_1 FILLER_20_3364 ();
 sg13g2_decap_8 FILLER_20_3385 ();
 sg13g2_fill_1 FILLER_20_3392 ();
 sg13g2_fill_2 FILLER_20_3447 ();
 sg13g2_decap_8 FILLER_20_3462 ();
 sg13g2_fill_2 FILLER_20_3469 ();
 sg13g2_decap_8 FILLER_20_3492 ();
 sg13g2_fill_1 FILLER_20_3503 ();
 sg13g2_decap_4 FILLER_20_3509 ();
 sg13g2_fill_2 FILLER_20_3527 ();
 sg13g2_fill_1 FILLER_20_3533 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_4 FILLER_21_70 ();
 sg13g2_fill_1 FILLER_21_74 ();
 sg13g2_fill_1 FILLER_21_98 ();
 sg13g2_fill_2 FILLER_21_107 ();
 sg13g2_fill_1 FILLER_21_168 ();
 sg13g2_fill_2 FILLER_21_242 ();
 sg13g2_fill_2 FILLER_21_419 ();
 sg13g2_fill_2 FILLER_21_466 ();
 sg13g2_fill_1 FILLER_21_468 ();
 sg13g2_fill_1 FILLER_21_478 ();
 sg13g2_fill_2 FILLER_21_520 ();
 sg13g2_fill_1 FILLER_21_522 ();
 sg13g2_fill_1 FILLER_21_580 ();
 sg13g2_fill_1 FILLER_21_633 ();
 sg13g2_fill_2 FILLER_21_654 ();
 sg13g2_decap_4 FILLER_21_682 ();
 sg13g2_fill_1 FILLER_21_714 ();
 sg13g2_fill_1 FILLER_21_724 ();
 sg13g2_fill_1 FILLER_21_734 ();
 sg13g2_fill_1 FILLER_21_776 ();
 sg13g2_fill_1 FILLER_21_791 ();
 sg13g2_fill_1 FILLER_21_801 ();
 sg13g2_fill_1 FILLER_21_820 ();
 sg13g2_fill_2 FILLER_21_843 ();
 sg13g2_fill_2 FILLER_21_857 ();
 sg13g2_fill_2 FILLER_21_886 ();
 sg13g2_fill_1 FILLER_21_943 ();
 sg13g2_fill_2 FILLER_21_971 ();
 sg13g2_decap_4 FILLER_21_993 ();
 sg13g2_fill_2 FILLER_21_1119 ();
 sg13g2_fill_1 FILLER_21_1121 ();
 sg13g2_fill_2 FILLER_21_1158 ();
 sg13g2_fill_2 FILLER_21_1245 ();
 sg13g2_decap_4 FILLER_21_1269 ();
 sg13g2_fill_1 FILLER_21_1273 ();
 sg13g2_fill_2 FILLER_21_1310 ();
 sg13g2_fill_1 FILLER_21_1312 ();
 sg13g2_fill_1 FILLER_21_1321 ();
 sg13g2_fill_2 FILLER_21_1330 ();
 sg13g2_fill_1 FILLER_21_1332 ();
 sg13g2_fill_2 FILLER_21_1366 ();
 sg13g2_fill_2 FILLER_21_1399 ();
 sg13g2_fill_2 FILLER_21_1407 ();
 sg13g2_decap_4 FILLER_21_1447 ();
 sg13g2_fill_1 FILLER_21_1478 ();
 sg13g2_decap_8 FILLER_21_1587 ();
 sg13g2_fill_1 FILLER_21_1598 ();
 sg13g2_decap_8 FILLER_21_1604 ();
 sg13g2_fill_2 FILLER_21_1611 ();
 sg13g2_decap_4 FILLER_21_1637 ();
 sg13g2_fill_2 FILLER_21_1653 ();
 sg13g2_fill_2 FILLER_21_1660 ();
 sg13g2_fill_1 FILLER_21_1670 ();
 sg13g2_decap_4 FILLER_21_1683 ();
 sg13g2_decap_8 FILLER_21_1723 ();
 sg13g2_fill_1 FILLER_21_1730 ();
 sg13g2_fill_1 FILLER_21_1749 ();
 sg13g2_decap_4 FILLER_21_1755 ();
 sg13g2_fill_2 FILLER_21_1759 ();
 sg13g2_fill_2 FILLER_21_1782 ();
 sg13g2_fill_1 FILLER_21_1808 ();
 sg13g2_fill_1 FILLER_21_1827 ();
 sg13g2_fill_1 FILLER_21_1844 ();
 sg13g2_decap_8 FILLER_21_1907 ();
 sg13g2_fill_1 FILLER_21_1914 ();
 sg13g2_decap_8 FILLER_21_1919 ();
 sg13g2_fill_2 FILLER_21_1934 ();
 sg13g2_fill_1 FILLER_21_1936 ();
 sg13g2_fill_1 FILLER_21_1953 ();
 sg13g2_decap_8 FILLER_21_1991 ();
 sg13g2_decap_4 FILLER_21_2059 ();
 sg13g2_fill_2 FILLER_21_2063 ();
 sg13g2_fill_2 FILLER_21_2078 ();
 sg13g2_fill_1 FILLER_21_2080 ();
 sg13g2_fill_2 FILLER_21_2092 ();
 sg13g2_decap_8 FILLER_21_2098 ();
 sg13g2_decap_4 FILLER_21_2105 ();
 sg13g2_fill_1 FILLER_21_2109 ();
 sg13g2_fill_2 FILLER_21_2126 ();
 sg13g2_fill_1 FILLER_21_2128 ();
 sg13g2_fill_1 FILLER_21_2141 ();
 sg13g2_decap_4 FILLER_21_2150 ();
 sg13g2_fill_2 FILLER_21_2164 ();
 sg13g2_decap_8 FILLER_21_2183 ();
 sg13g2_decap_4 FILLER_21_2190 ();
 sg13g2_fill_1 FILLER_21_2194 ();
 sg13g2_fill_2 FILLER_21_2213 ();
 sg13g2_fill_1 FILLER_21_2215 ();
 sg13g2_decap_4 FILLER_21_2243 ();
 sg13g2_fill_2 FILLER_21_2247 ();
 sg13g2_decap_4 FILLER_21_2294 ();
 sg13g2_fill_1 FILLER_21_2298 ();
 sg13g2_fill_1 FILLER_21_2321 ();
 sg13g2_decap_4 FILLER_21_2343 ();
 sg13g2_fill_1 FILLER_21_2347 ();
 sg13g2_fill_1 FILLER_21_2353 ();
 sg13g2_fill_2 FILLER_21_2371 ();
 sg13g2_fill_1 FILLER_21_2373 ();
 sg13g2_fill_1 FILLER_21_2441 ();
 sg13g2_fill_1 FILLER_21_2469 ();
 sg13g2_fill_1 FILLER_21_2483 ();
 sg13g2_decap_4 FILLER_21_2492 ();
 sg13g2_fill_1 FILLER_21_2496 ();
 sg13g2_decap_4 FILLER_21_2505 ();
 sg13g2_fill_2 FILLER_21_2509 ();
 sg13g2_fill_2 FILLER_21_2539 ();
 sg13g2_fill_2 FILLER_21_2564 ();
 sg13g2_fill_2 FILLER_21_2574 ();
 sg13g2_decap_8 FILLER_21_2589 ();
 sg13g2_fill_2 FILLER_21_2596 ();
 sg13g2_decap_4 FILLER_21_2630 ();
 sg13g2_fill_1 FILLER_21_2647 ();
 sg13g2_fill_1 FILLER_21_2653 ();
 sg13g2_fill_2 FILLER_21_2673 ();
 sg13g2_fill_1 FILLER_21_2675 ();
 sg13g2_fill_2 FILLER_21_2684 ();
 sg13g2_fill_2 FILLER_21_2703 ();
 sg13g2_fill_2 FILLER_21_2715 ();
 sg13g2_decap_8 FILLER_21_2727 ();
 sg13g2_fill_1 FILLER_21_2734 ();
 sg13g2_decap_4 FILLER_21_2741 ();
 sg13g2_fill_1 FILLER_21_2745 ();
 sg13g2_fill_2 FILLER_21_2782 ();
 sg13g2_decap_4 FILLER_21_2808 ();
 sg13g2_fill_2 FILLER_21_2812 ();
 sg13g2_decap_8 FILLER_21_2834 ();
 sg13g2_fill_2 FILLER_21_2841 ();
 sg13g2_fill_1 FILLER_21_2871 ();
 sg13g2_fill_2 FILLER_21_2913 ();
 sg13g2_fill_1 FILLER_21_2945 ();
 sg13g2_fill_1 FILLER_21_2961 ();
 sg13g2_decap_4 FILLER_21_3064 ();
 sg13g2_fill_2 FILLER_21_3068 ();
 sg13g2_fill_2 FILLER_21_3105 ();
 sg13g2_fill_1 FILLER_21_3107 ();
 sg13g2_fill_1 FILLER_21_3112 ();
 sg13g2_fill_1 FILLER_21_3184 ();
 sg13g2_fill_1 FILLER_21_3269 ();
 sg13g2_fill_2 FILLER_21_3435 ();
 sg13g2_fill_1 FILLER_21_3437 ();
 sg13g2_decap_4 FILLER_21_3447 ();
 sg13g2_fill_1 FILLER_21_3451 ();
 sg13g2_fill_1 FILLER_21_3492 ();
 sg13g2_decap_4 FILLER_21_3501 ();
 sg13g2_fill_2 FILLER_21_3505 ();
 sg13g2_fill_2 FILLER_21_3515 ();
 sg13g2_fill_1 FILLER_21_3517 ();
 sg13g2_fill_2 FILLER_21_3547 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_2 ();
 sg13g2_fill_1 FILLER_22_31 ();
 sg13g2_fill_2 FILLER_22_53 ();
 sg13g2_fill_1 FILLER_22_55 ();
 sg13g2_decap_4 FILLER_22_62 ();
 sg13g2_decap_8 FILLER_22_71 ();
 sg13g2_fill_1 FILLER_22_88 ();
 sg13g2_decap_8 FILLER_22_108 ();
 sg13g2_decap_4 FILLER_22_115 ();
 sg13g2_fill_1 FILLER_22_119 ();
 sg13g2_fill_2 FILLER_22_143 ();
 sg13g2_fill_1 FILLER_22_209 ();
 sg13g2_fill_1 FILLER_22_281 ();
 sg13g2_fill_1 FILLER_22_296 ();
 sg13g2_fill_1 FILLER_22_348 ();
 sg13g2_fill_2 FILLER_22_402 ();
 sg13g2_fill_1 FILLER_22_475 ();
 sg13g2_fill_1 FILLER_22_498 ();
 sg13g2_fill_2 FILLER_22_517 ();
 sg13g2_fill_1 FILLER_22_551 ();
 sg13g2_fill_1 FILLER_22_588 ();
 sg13g2_fill_1 FILLER_22_613 ();
 sg13g2_fill_2 FILLER_22_623 ();
 sg13g2_fill_1 FILLER_22_625 ();
 sg13g2_fill_1 FILLER_22_636 ();
 sg13g2_fill_2 FILLER_22_664 ();
 sg13g2_fill_2 FILLER_22_964 ();
 sg13g2_fill_1 FILLER_22_966 ();
 sg13g2_fill_2 FILLER_22_977 ();
 sg13g2_fill_1 FILLER_22_979 ();
 sg13g2_fill_2 FILLER_22_1007 ();
 sg13g2_fill_2 FILLER_22_1157 ();
 sg13g2_fill_2 FILLER_22_1212 ();
 sg13g2_fill_2 FILLER_22_1228 ();
 sg13g2_fill_2 FILLER_22_1244 ();
 sg13g2_decap_4 FILLER_22_1294 ();
 sg13g2_fill_1 FILLER_22_1298 ();
 sg13g2_fill_2 FILLER_22_1339 ();
 sg13g2_fill_1 FILLER_22_1341 ();
 sg13g2_fill_1 FILLER_22_1359 ();
 sg13g2_fill_1 FILLER_22_1398 ();
 sg13g2_decap_4 FILLER_22_1422 ();
 sg13g2_fill_1 FILLER_22_1426 ();
 sg13g2_fill_1 FILLER_22_1436 ();
 sg13g2_decap_8 FILLER_22_1461 ();
 sg13g2_fill_1 FILLER_22_1468 ();
 sg13g2_fill_1 FILLER_22_1473 ();
 sg13g2_fill_1 FILLER_22_1477 ();
 sg13g2_decap_4 FILLER_22_1509 ();
 sg13g2_fill_2 FILLER_22_1531 ();
 sg13g2_fill_1 FILLER_22_1533 ();
 sg13g2_decap_8 FILLER_22_1554 ();
 sg13g2_fill_2 FILLER_22_1561 ();
 sg13g2_fill_2 FILLER_22_1609 ();
 sg13g2_decap_4 FILLER_22_1623 ();
 sg13g2_decap_8 FILLER_22_1635 ();
 sg13g2_decap_4 FILLER_22_1642 ();
 sg13g2_decap_8 FILLER_22_1681 ();
 sg13g2_fill_2 FILLER_22_1688 ();
 sg13g2_fill_1 FILLER_22_1690 ();
 sg13g2_decap_8 FILLER_22_1699 ();
 sg13g2_fill_2 FILLER_22_1710 ();
 sg13g2_decap_8 FILLER_22_1716 ();
 sg13g2_fill_2 FILLER_22_1723 ();
 sg13g2_decap_8 FILLER_22_1757 ();
 sg13g2_decap_4 FILLER_22_1764 ();
 sg13g2_fill_1 FILLER_22_1772 ();
 sg13g2_decap_8 FILLER_22_1776 ();
 sg13g2_decap_4 FILLER_22_1790 ();
 sg13g2_fill_1 FILLER_22_1794 ();
 sg13g2_fill_2 FILLER_22_1800 ();
 sg13g2_fill_2 FILLER_22_1850 ();
 sg13g2_fill_2 FILLER_22_1893 ();
 sg13g2_fill_1 FILLER_22_1895 ();
 sg13g2_fill_2 FILLER_22_1914 ();
 sg13g2_decap_8 FILLER_22_1949 ();
 sg13g2_fill_2 FILLER_22_1956 ();
 sg13g2_fill_1 FILLER_22_1958 ();
 sg13g2_fill_2 FILLER_22_1972 ();
 sg13g2_fill_2 FILLER_22_2001 ();
 sg13g2_fill_2 FILLER_22_2029 ();
 sg13g2_fill_1 FILLER_22_2031 ();
 sg13g2_fill_2 FILLER_22_2042 ();
 sg13g2_fill_2 FILLER_22_2080 ();
 sg13g2_decap_4 FILLER_22_2106 ();
 sg13g2_fill_1 FILLER_22_2110 ();
 sg13g2_fill_1 FILLER_22_2116 ();
 sg13g2_decap_4 FILLER_22_2123 ();
 sg13g2_fill_1 FILLER_22_2190 ();
 sg13g2_fill_2 FILLER_22_2215 ();
 sg13g2_fill_1 FILLER_22_2217 ();
 sg13g2_decap_4 FILLER_22_2223 ();
 sg13g2_fill_1 FILLER_22_2232 ();
 sg13g2_fill_2 FILLER_22_2241 ();
 sg13g2_fill_1 FILLER_22_2243 ();
 sg13g2_fill_1 FILLER_22_2253 ();
 sg13g2_decap_8 FILLER_22_2258 ();
 sg13g2_decap_4 FILLER_22_2265 ();
 sg13g2_fill_2 FILLER_22_2269 ();
 sg13g2_fill_1 FILLER_22_2306 ();
 sg13g2_decap_8 FILLER_22_2316 ();
 sg13g2_decap_8 FILLER_22_2323 ();
 sg13g2_decap_8 FILLER_22_2330 ();
 sg13g2_decap_8 FILLER_22_2337 ();
 sg13g2_fill_2 FILLER_22_2344 ();
 sg13g2_fill_1 FILLER_22_2346 ();
 sg13g2_decap_8 FILLER_22_2382 ();
 sg13g2_decap_8 FILLER_22_2389 ();
 sg13g2_decap_8 FILLER_22_2396 ();
 sg13g2_decap_4 FILLER_22_2414 ();
 sg13g2_fill_2 FILLER_22_2441 ();
 sg13g2_fill_1 FILLER_22_2451 ();
 sg13g2_fill_1 FILLER_22_2466 ();
 sg13g2_decap_8 FILLER_22_2477 ();
 sg13g2_fill_2 FILLER_22_2484 ();
 sg13g2_decap_4 FILLER_22_2510 ();
 sg13g2_fill_2 FILLER_22_2514 ();
 sg13g2_decap_8 FILLER_22_2520 ();
 sg13g2_decap_8 FILLER_22_2527 ();
 sg13g2_fill_2 FILLER_22_2534 ();
 sg13g2_fill_2 FILLER_22_2571 ();
 sg13g2_fill_1 FILLER_22_2573 ();
 sg13g2_decap_4 FILLER_22_2597 ();
 sg13g2_fill_1 FILLER_22_2601 ();
 sg13g2_fill_2 FILLER_22_2616 ();
 sg13g2_fill_1 FILLER_22_2618 ();
 sg13g2_fill_2 FILLER_22_2624 ();
 sg13g2_fill_1 FILLER_22_2626 ();
 sg13g2_fill_1 FILLER_22_2632 ();
 sg13g2_fill_1 FILLER_22_2661 ();
 sg13g2_fill_1 FILLER_22_2699 ();
 sg13g2_decap_8 FILLER_22_2705 ();
 sg13g2_fill_1 FILLER_22_2712 ();
 sg13g2_fill_1 FILLER_22_2727 ();
 sg13g2_decap_8 FILLER_22_2745 ();
 sg13g2_fill_1 FILLER_22_2773 ();
 sg13g2_decap_4 FILLER_22_2803 ();
 sg13g2_fill_2 FILLER_22_2807 ();
 sg13g2_fill_1 FILLER_22_2813 ();
 sg13g2_fill_2 FILLER_22_2836 ();
 sg13g2_fill_1 FILLER_22_2838 ();
 sg13g2_fill_1 FILLER_22_2859 ();
 sg13g2_fill_2 FILLER_22_2865 ();
 sg13g2_fill_2 FILLER_22_2898 ();
 sg13g2_fill_1 FILLER_22_2912 ();
 sg13g2_decap_8 FILLER_22_2944 ();
 sg13g2_fill_2 FILLER_22_2955 ();
 sg13g2_fill_1 FILLER_22_2957 ();
 sg13g2_fill_1 FILLER_22_2963 ();
 sg13g2_fill_2 FILLER_22_2968 ();
 sg13g2_fill_1 FILLER_22_2970 ();
 sg13g2_fill_1 FILLER_22_3005 ();
 sg13g2_fill_1 FILLER_22_3018 ();
 sg13g2_fill_1 FILLER_22_3028 ();
 sg13g2_fill_2 FILLER_22_3043 ();
 sg13g2_fill_2 FILLER_22_3127 ();
 sg13g2_fill_1 FILLER_22_3129 ();
 sg13g2_fill_2 FILLER_22_3139 ();
 sg13g2_fill_2 FILLER_22_3150 ();
 sg13g2_fill_1 FILLER_22_3152 ();
 sg13g2_fill_1 FILLER_22_3195 ();
 sg13g2_fill_2 FILLER_22_3205 ();
 sg13g2_fill_1 FILLER_22_3212 ();
 sg13g2_fill_2 FILLER_22_3222 ();
 sg13g2_fill_1 FILLER_22_3224 ();
 sg13g2_fill_2 FILLER_22_3288 ();
 sg13g2_fill_1 FILLER_22_3290 ();
 sg13g2_fill_1 FILLER_22_3312 ();
 sg13g2_fill_2 FILLER_22_3374 ();
 sg13g2_decap_4 FILLER_22_3452 ();
 sg13g2_fill_2 FILLER_22_3471 ();
 sg13g2_fill_1 FILLER_22_3473 ();
 sg13g2_fill_2 FILLER_22_3494 ();
 sg13g2_fill_1 FILLER_22_3496 ();
 sg13g2_decap_4 FILLER_22_3512 ();
 sg13g2_fill_1 FILLER_22_3516 ();
 sg13g2_decap_4 FILLER_22_3532 ();
 sg13g2_fill_1 FILLER_22_3536 ();
 sg13g2_fill_1 FILLER_22_3545 ();
 sg13g2_fill_1 FILLER_22_3551 ();
 sg13g2_fill_2 FILLER_22_3565 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_29 ();
 sg13g2_fill_1 FILLER_23_47 ();
 sg13g2_decap_4 FILLER_23_57 ();
 sg13g2_fill_2 FILLER_23_61 ();
 sg13g2_decap_4 FILLER_23_68 ();
 sg13g2_fill_1 FILLER_23_85 ();
 sg13g2_fill_1 FILLER_23_275 ();
 sg13g2_fill_1 FILLER_23_406 ();
 sg13g2_fill_2 FILLER_23_438 ();
 sg13g2_fill_1 FILLER_23_518 ();
 sg13g2_fill_2 FILLER_23_554 ();
 sg13g2_fill_1 FILLER_23_556 ();
 sg13g2_fill_1 FILLER_23_580 ();
 sg13g2_fill_1 FILLER_23_653 ();
 sg13g2_fill_1 FILLER_23_664 ();
 sg13g2_fill_2 FILLER_23_724 ();
 sg13g2_fill_1 FILLER_23_726 ();
 sg13g2_fill_2 FILLER_23_748 ();
 sg13g2_fill_1 FILLER_23_750 ();
 sg13g2_fill_1 FILLER_23_808 ();
 sg13g2_fill_2 FILLER_23_953 ();
 sg13g2_fill_2 FILLER_23_965 ();
 sg13g2_fill_1 FILLER_23_967 ();
 sg13g2_fill_1 FILLER_23_1081 ();
 sg13g2_fill_2 FILLER_23_1109 ();
 sg13g2_fill_1 FILLER_23_1111 ();
 sg13g2_fill_1 FILLER_23_1148 ();
 sg13g2_decap_8 FILLER_23_1301 ();
 sg13g2_decap_8 FILLER_23_1308 ();
 sg13g2_decap_4 FILLER_23_1328 ();
 sg13g2_fill_2 FILLER_23_1363 ();
 sg13g2_fill_2 FILLER_23_1383 ();
 sg13g2_fill_1 FILLER_23_1385 ();
 sg13g2_fill_2 FILLER_23_1416 ();
 sg13g2_fill_2 FILLER_23_1426 ();
 sg13g2_fill_1 FILLER_23_1447 ();
 sg13g2_fill_2 FILLER_23_1458 ();
 sg13g2_fill_1 FILLER_23_1460 ();
 sg13g2_fill_2 FILLER_23_1469 ();
 sg13g2_fill_1 FILLER_23_1498 ();
 sg13g2_decap_4 FILLER_23_1514 ();
 sg13g2_decap_4 FILLER_23_1548 ();
 sg13g2_fill_1 FILLER_23_1552 ();
 sg13g2_decap_4 FILLER_23_1557 ();
 sg13g2_fill_1 FILLER_23_1561 ();
 sg13g2_fill_2 FILLER_23_1588 ();
 sg13g2_fill_1 FILLER_23_1590 ();
 sg13g2_fill_2 FILLER_23_1600 ();
 sg13g2_fill_1 FILLER_23_1602 ();
 sg13g2_decap_4 FILLER_23_1628 ();
 sg13g2_fill_1 FILLER_23_1632 ();
 sg13g2_fill_2 FILLER_23_1661 ();
 sg13g2_fill_2 FILLER_23_1676 ();
 sg13g2_fill_1 FILLER_23_1686 ();
 sg13g2_fill_1 FILLER_23_1732 ();
 sg13g2_decap_4 FILLER_23_1741 ();
 sg13g2_decap_4 FILLER_23_1749 ();
 sg13g2_fill_2 FILLER_23_1753 ();
 sg13g2_fill_2 FILLER_23_1791 ();
 sg13g2_fill_1 FILLER_23_1804 ();
 sg13g2_fill_1 FILLER_23_1810 ();
 sg13g2_fill_1 FILLER_23_1865 ();
 sg13g2_decap_4 FILLER_23_1882 ();
 sg13g2_fill_1 FILLER_23_1886 ();
 sg13g2_fill_1 FILLER_23_1891 ();
 sg13g2_decap_4 FILLER_23_1917 ();
 sg13g2_decap_8 FILLER_23_1945 ();
 sg13g2_fill_2 FILLER_23_1984 ();
 sg13g2_decap_8 FILLER_23_1999 ();
 sg13g2_decap_4 FILLER_23_2006 ();
 sg13g2_decap_4 FILLER_23_2023 ();
 sg13g2_fill_1 FILLER_23_2027 ();
 sg13g2_fill_1 FILLER_23_2056 ();
 sg13g2_fill_1 FILLER_23_2062 ();
 sg13g2_fill_1 FILLER_23_2080 ();
 sg13g2_fill_1 FILLER_23_2087 ();
 sg13g2_fill_2 FILLER_23_2199 ();
 sg13g2_fill_1 FILLER_23_2201 ();
 sg13g2_decap_4 FILLER_23_2220 ();
 sg13g2_decap_8 FILLER_23_2255 ();
 sg13g2_fill_2 FILLER_23_2280 ();
 sg13g2_fill_2 FILLER_23_2296 ();
 sg13g2_fill_1 FILLER_23_2298 ();
 sg13g2_decap_4 FILLER_23_2341 ();
 sg13g2_fill_2 FILLER_23_2378 ();
 sg13g2_fill_2 FILLER_23_2402 ();
 sg13g2_fill_1 FILLER_23_2404 ();
 sg13g2_fill_1 FILLER_23_2421 ();
 sg13g2_fill_1 FILLER_23_2456 ();
 sg13g2_fill_1 FILLER_23_2475 ();
 sg13g2_fill_2 FILLER_23_2485 ();
 sg13g2_decap_4 FILLER_23_2517 ();
 sg13g2_fill_2 FILLER_23_2521 ();
 sg13g2_decap_8 FILLER_23_2527 ();
 sg13g2_decap_8 FILLER_23_2534 ();
 sg13g2_fill_2 FILLER_23_2541 ();
 sg13g2_fill_1 FILLER_23_2543 ();
 sg13g2_decap_8 FILLER_23_2568 ();
 sg13g2_decap_4 FILLER_23_2575 ();
 sg13g2_decap_8 FILLER_23_2592 ();
 sg13g2_fill_2 FILLER_23_2599 ();
 sg13g2_fill_1 FILLER_23_2601 ();
 sg13g2_fill_1 FILLER_23_2642 ();
 sg13g2_fill_2 FILLER_23_2655 ();
 sg13g2_fill_1 FILLER_23_2657 ();
 sg13g2_fill_2 FILLER_23_2666 ();
 sg13g2_decap_8 FILLER_23_2672 ();
 sg13g2_decap_8 FILLER_23_2679 ();
 sg13g2_decap_8 FILLER_23_2686 ();
 sg13g2_fill_2 FILLER_23_2706 ();
 sg13g2_fill_2 FILLER_23_2723 ();
 sg13g2_fill_1 FILLER_23_2725 ();
 sg13g2_fill_2 FILLER_23_2748 ();
 sg13g2_fill_1 FILLER_23_2750 ();
 sg13g2_fill_2 FILLER_23_2759 ();
 sg13g2_fill_2 FILLER_23_2766 ();
 sg13g2_fill_2 FILLER_23_2771 ();
 sg13g2_fill_2 FILLER_23_2781 ();
 sg13g2_decap_4 FILLER_23_2800 ();
 sg13g2_fill_1 FILLER_23_2804 ();
 sg13g2_fill_2 FILLER_23_2831 ();
 sg13g2_fill_1 FILLER_23_2833 ();
 sg13g2_decap_4 FILLER_23_2884 ();
 sg13g2_fill_2 FILLER_23_2896 ();
 sg13g2_fill_1 FILLER_23_2898 ();
 sg13g2_fill_2 FILLER_23_2918 ();
 sg13g2_fill_1 FILLER_23_2920 ();
 sg13g2_fill_2 FILLER_23_2935 ();
 sg13g2_decap_4 FILLER_23_2948 ();
 sg13g2_fill_2 FILLER_23_2974 ();
 sg13g2_fill_1 FILLER_23_2976 ();
 sg13g2_fill_1 FILLER_23_3022 ();
 sg13g2_fill_2 FILLER_23_3056 ();
 sg13g2_fill_1 FILLER_23_3058 ();
 sg13g2_fill_2 FILLER_23_3067 ();
 sg13g2_fill_1 FILLER_23_3069 ();
 sg13g2_fill_1 FILLER_23_3093 ();
 sg13g2_fill_2 FILLER_23_3110 ();
 sg13g2_decap_8 FILLER_23_3125 ();
 sg13g2_fill_2 FILLER_23_3132 ();
 sg13g2_fill_1 FILLER_23_3134 ();
 sg13g2_decap_8 FILLER_23_3149 ();
 sg13g2_fill_2 FILLER_23_3156 ();
 sg13g2_fill_1 FILLER_23_3181 ();
 sg13g2_fill_1 FILLER_23_3191 ();
 sg13g2_fill_1 FILLER_23_3219 ();
 sg13g2_fill_2 FILLER_23_3239 ();
 sg13g2_fill_2 FILLER_23_3276 ();
 sg13g2_fill_1 FILLER_23_3278 ();
 sg13g2_fill_2 FILLER_23_3346 ();
 sg13g2_fill_1 FILLER_23_3406 ();
 sg13g2_fill_2 FILLER_23_3435 ();
 sg13g2_decap_8 FILLER_23_3445 ();
 sg13g2_fill_2 FILLER_23_3452 ();
 sg13g2_fill_2 FILLER_23_3479 ();
 sg13g2_fill_1 FILLER_23_3481 ();
 sg13g2_decap_4 FILLER_23_3503 ();
 sg13g2_fill_2 FILLER_23_3507 ();
 sg13g2_fill_1 FILLER_23_3518 ();
 sg13g2_fill_2 FILLER_23_3534 ();
 sg13g2_fill_1 FILLER_23_3536 ();
 sg13g2_fill_1 FILLER_23_3551 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_12 ();
 sg13g2_fill_2 FILLER_24_19 ();
 sg13g2_fill_1 FILLER_24_21 ();
 sg13g2_fill_1 FILLER_24_43 ();
 sg13g2_decap_8 FILLER_24_73 ();
 sg13g2_fill_1 FILLER_24_80 ();
 sg13g2_fill_2 FILLER_24_100 ();
 sg13g2_fill_1 FILLER_24_102 ();
 sg13g2_fill_1 FILLER_24_178 ();
 sg13g2_fill_1 FILLER_24_288 ();
 sg13g2_fill_1 FILLER_24_348 ();
 sg13g2_fill_1 FILLER_24_364 ();
 sg13g2_fill_1 FILLER_24_410 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_fill_2 FILLER_24_467 ();
 sg13g2_fill_1 FILLER_24_469 ();
 sg13g2_fill_2 FILLER_24_498 ();
 sg13g2_fill_1 FILLER_24_500 ();
 sg13g2_fill_2 FILLER_24_540 ();
 sg13g2_fill_1 FILLER_24_584 ();
 sg13g2_fill_1 FILLER_24_630 ();
 sg13g2_fill_2 FILLER_24_681 ();
 sg13g2_fill_2 FILLER_24_779 ();
 sg13g2_fill_2 FILLER_24_796 ();
 sg13g2_fill_1 FILLER_24_833 ();
 sg13g2_fill_1 FILLER_24_862 ();
 sg13g2_fill_2 FILLER_24_897 ();
 sg13g2_fill_1 FILLER_24_899 ();
 sg13g2_fill_2 FILLER_24_944 ();
 sg13g2_fill_1 FILLER_24_946 ();
 sg13g2_fill_1 FILLER_24_992 ();
 sg13g2_fill_1 FILLER_24_1006 ();
 sg13g2_fill_1 FILLER_24_1168 ();
 sg13g2_fill_2 FILLER_24_1178 ();
 sg13g2_fill_1 FILLER_24_1226 ();
 sg13g2_fill_2 FILLER_24_1268 ();
 sg13g2_fill_1 FILLER_24_1346 ();
 sg13g2_decap_8 FILLER_24_1366 ();
 sg13g2_fill_2 FILLER_24_1373 ();
 sg13g2_fill_1 FILLER_24_1375 ();
 sg13g2_fill_2 FILLER_24_1389 ();
 sg13g2_fill_1 FILLER_24_1401 ();
 sg13g2_fill_2 FILLER_24_1421 ();
 sg13g2_fill_2 FILLER_24_1469 ();
 sg13g2_fill_2 FILLER_24_1485 ();
 sg13g2_fill_1 FILLER_24_1487 ();
 sg13g2_fill_1 FILLER_24_1514 ();
 sg13g2_fill_1 FILLER_24_1576 ();
 sg13g2_fill_1 FILLER_24_1595 ();
 sg13g2_fill_2 FILLER_24_1629 ();
 sg13g2_fill_1 FILLER_24_1631 ();
 sg13g2_fill_1 FILLER_24_1663 ();
 sg13g2_fill_1 FILLER_24_1701 ();
 sg13g2_fill_2 FILLER_24_1716 ();
 sg13g2_fill_2 FILLER_24_1726 ();
 sg13g2_fill_2 FILLER_24_1747 ();
 sg13g2_fill_1 FILLER_24_1757 ();
 sg13g2_decap_8 FILLER_24_1777 ();
 sg13g2_fill_2 FILLER_24_1784 ();
 sg13g2_decap_8 FILLER_24_1840 ();
 sg13g2_fill_1 FILLER_24_1847 ();
 sg13g2_fill_2 FILLER_24_1858 ();
 sg13g2_fill_1 FILLER_24_1860 ();
 sg13g2_fill_2 FILLER_24_1866 ();
 sg13g2_fill_1 FILLER_24_1868 ();
 sg13g2_decap_4 FILLER_24_1878 ();
 sg13g2_fill_2 FILLER_24_1882 ();
 sg13g2_fill_2 FILLER_24_1925 ();
 sg13g2_fill_1 FILLER_24_1927 ();
 sg13g2_fill_2 FILLER_24_1956 ();
 sg13g2_fill_2 FILLER_24_2022 ();
 sg13g2_fill_1 FILLER_24_2024 ();
 sg13g2_decap_8 FILLER_24_2079 ();
 sg13g2_fill_2 FILLER_24_2100 ();
 sg13g2_decap_8 FILLER_24_2124 ();
 sg13g2_decap_8 FILLER_24_2131 ();
 sg13g2_fill_2 FILLER_24_2138 ();
 sg13g2_fill_1 FILLER_24_2140 ();
 sg13g2_decap_4 FILLER_24_2199 ();
 sg13g2_fill_2 FILLER_24_2203 ();
 sg13g2_fill_2 FILLER_24_2220 ();
 sg13g2_fill_1 FILLER_24_2222 ();
 sg13g2_fill_1 FILLER_24_2242 ();
 sg13g2_fill_1 FILLER_24_2313 ();
 sg13g2_fill_2 FILLER_24_2323 ();
 sg13g2_decap_4 FILLER_24_2334 ();
 sg13g2_fill_1 FILLER_24_2351 ();
 sg13g2_decap_4 FILLER_24_2358 ();
 sg13g2_fill_1 FILLER_24_2403 ();
 sg13g2_fill_1 FILLER_24_2425 ();
 sg13g2_fill_1 FILLER_24_2432 ();
 sg13g2_fill_2 FILLER_24_2446 ();
 sg13g2_fill_2 FILLER_24_2452 ();
 sg13g2_fill_1 FILLER_24_2465 ();
 sg13g2_fill_2 FILLER_24_2489 ();
 sg13g2_fill_1 FILLER_24_2491 ();
 sg13g2_decap_8 FILLER_24_2500 ();
 sg13g2_fill_1 FILLER_24_2507 ();
 sg13g2_decap_4 FILLER_24_2513 ();
 sg13g2_fill_1 FILLER_24_2517 ();
 sg13g2_fill_2 FILLER_24_2567 ();
 sg13g2_decap_4 FILLER_24_2579 ();
 sg13g2_decap_4 FILLER_24_2603 ();
 sg13g2_fill_2 FILLER_24_2628 ();
 sg13g2_fill_1 FILLER_24_2635 ();
 sg13g2_decap_8 FILLER_24_2663 ();
 sg13g2_fill_2 FILLER_24_2670 ();
 sg13g2_fill_1 FILLER_24_2672 ();
 sg13g2_decap_4 FILLER_24_2685 ();
 sg13g2_fill_1 FILLER_24_2689 ();
 sg13g2_decap_4 FILLER_24_2706 ();
 sg13g2_fill_2 FILLER_24_2715 ();
 sg13g2_fill_2 FILLER_24_2722 ();
 sg13g2_fill_2 FILLER_24_2732 ();
 sg13g2_fill_2 FILLER_24_2740 ();
 sg13g2_fill_1 FILLER_24_2742 ();
 sg13g2_decap_4 FILLER_24_2776 ();
 sg13g2_fill_1 FILLER_24_2780 ();
 sg13g2_decap_4 FILLER_24_2803 ();
 sg13g2_fill_1 FILLER_24_2807 ();
 sg13g2_decap_8 FILLER_24_2821 ();
 sg13g2_fill_2 FILLER_24_2828 ();
 sg13g2_fill_2 FILLER_24_2849 ();
 sg13g2_fill_1 FILLER_24_2851 ();
 sg13g2_decap_8 FILLER_24_2878 ();
 sg13g2_fill_1 FILLER_24_2885 ();
 sg13g2_fill_1 FILLER_24_2895 ();
 sg13g2_fill_2 FILLER_24_2919 ();
 sg13g2_fill_1 FILLER_24_2921 ();
 sg13g2_fill_1 FILLER_24_2930 ();
 sg13g2_fill_1 FILLER_24_2949 ();
 sg13g2_fill_2 FILLER_24_2959 ();
 sg13g2_fill_1 FILLER_24_2961 ();
 sg13g2_fill_1 FILLER_24_2976 ();
 sg13g2_fill_1 FILLER_24_3003 ();
 sg13g2_fill_1 FILLER_24_3024 ();
 sg13g2_fill_2 FILLER_24_3036 ();
 sg13g2_fill_1 FILLER_24_3038 ();
 sg13g2_fill_2 FILLER_24_3066 ();
 sg13g2_fill_1 FILLER_24_3068 ();
 sg13g2_fill_2 FILLER_24_3093 ();
 sg13g2_decap_8 FILLER_24_3099 ();
 sg13g2_fill_2 FILLER_24_3106 ();
 sg13g2_fill_2 FILLER_24_3112 ();
 sg13g2_fill_1 FILLER_24_3114 ();
 sg13g2_fill_1 FILLER_24_3120 ();
 sg13g2_fill_2 FILLER_24_3149 ();
 sg13g2_decap_4 FILLER_24_3185 ();
 sg13g2_fill_1 FILLER_24_3189 ();
 sg13g2_fill_2 FILLER_24_3198 ();
 sg13g2_fill_2 FILLER_24_3294 ();
 sg13g2_fill_1 FILLER_24_3296 ();
 sg13g2_fill_1 FILLER_24_3359 ();
 sg13g2_fill_1 FILLER_24_3387 ();
 sg13g2_fill_2 FILLER_24_3401 ();
 sg13g2_fill_1 FILLER_24_3403 ();
 sg13g2_fill_1 FILLER_24_3416 ();
 sg13g2_decap_4 FILLER_24_3502 ();
 sg13g2_fill_1 FILLER_24_3560 ();
 sg13g2_fill_1 FILLER_24_3579 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_2 ();
 sg13g2_fill_1 FILLER_25_38 ();
 sg13g2_decap_4 FILLER_25_57 ();
 sg13g2_fill_1 FILLER_25_61 ();
 sg13g2_fill_2 FILLER_25_89 ();
 sg13g2_fill_1 FILLER_25_91 ();
 sg13g2_fill_1 FILLER_25_106 ();
 sg13g2_fill_2 FILLER_25_115 ();
 sg13g2_fill_2 FILLER_25_125 ();
 sg13g2_fill_1 FILLER_25_127 ();
 sg13g2_fill_1 FILLER_25_230 ();
 sg13g2_fill_1 FILLER_25_297 ();
 sg13g2_fill_1 FILLER_25_394 ();
 sg13g2_fill_1 FILLER_25_431 ();
 sg13g2_fill_2 FILLER_25_486 ();
 sg13g2_fill_1 FILLER_25_564 ();
 sg13g2_fill_1 FILLER_25_570 ();
 sg13g2_fill_2 FILLER_25_597 ();
 sg13g2_fill_1 FILLER_25_599 ();
 sg13g2_fill_1 FILLER_25_687 ();
 sg13g2_fill_1 FILLER_25_693 ();
 sg13g2_fill_1 FILLER_25_703 ();
 sg13g2_fill_1 FILLER_25_750 ();
 sg13g2_fill_1 FILLER_25_852 ();
 sg13g2_fill_1 FILLER_25_895 ();
 sg13g2_fill_2 FILLER_25_933 ();
 sg13g2_fill_1 FILLER_25_935 ();
 sg13g2_fill_1 FILLER_25_964 ();
 sg13g2_fill_2 FILLER_25_993 ();
 sg13g2_fill_2 FILLER_25_1008 ();
 sg13g2_fill_2 FILLER_25_1044 ();
 sg13g2_fill_2 FILLER_25_1131 ();
 sg13g2_fill_2 FILLER_25_1189 ();
 sg13g2_fill_1 FILLER_25_1191 ();
 sg13g2_fill_2 FILLER_25_1254 ();
 sg13g2_fill_2 FILLER_25_1273 ();
 sg13g2_fill_2 FILLER_25_1284 ();
 sg13g2_fill_2 FILLER_25_1308 ();
 sg13g2_decap_8 FILLER_25_1319 ();
 sg13g2_fill_2 FILLER_25_1326 ();
 sg13g2_decap_8 FILLER_25_1341 ();
 sg13g2_fill_1 FILLER_25_1348 ();
 sg13g2_fill_1 FILLER_25_1389 ();
 sg13g2_fill_2 FILLER_25_1400 ();
 sg13g2_fill_1 FILLER_25_1402 ();
 sg13g2_decap_8 FILLER_25_1423 ();
 sg13g2_fill_1 FILLER_25_1439 ();
 sg13g2_fill_2 FILLER_25_1465 ();
 sg13g2_decap_4 FILLER_25_1490 ();
 sg13g2_fill_2 FILLER_25_1494 ();
 sg13g2_fill_2 FILLER_25_1514 ();
 sg13g2_fill_1 FILLER_25_1516 ();
 sg13g2_fill_2 FILLER_25_1535 ();
 sg13g2_fill_1 FILLER_25_1537 ();
 sg13g2_decap_4 FILLER_25_1543 ();
 sg13g2_fill_1 FILLER_25_1547 ();
 sg13g2_decap_4 FILLER_25_1561 ();
 sg13g2_fill_2 FILLER_25_1612 ();
 sg13g2_decap_4 FILLER_25_1622 ();
 sg13g2_fill_2 FILLER_25_1626 ();
 sg13g2_fill_1 FILLER_25_1641 ();
 sg13g2_fill_2 FILLER_25_1687 ();
 sg13g2_fill_1 FILLER_25_1689 ();
 sg13g2_fill_2 FILLER_25_1707 ();
 sg13g2_fill_1 FILLER_25_1709 ();
 sg13g2_fill_1 FILLER_25_1715 ();
 sg13g2_fill_2 FILLER_25_1778 ();
 sg13g2_fill_1 FILLER_25_1780 ();
 sg13g2_decap_8 FILLER_25_1786 ();
 sg13g2_fill_2 FILLER_25_1793 ();
 sg13g2_fill_1 FILLER_25_1795 ();
 sg13g2_decap_8 FILLER_25_1801 ();
 sg13g2_decap_4 FILLER_25_1858 ();
 sg13g2_fill_2 FILLER_25_1898 ();
 sg13g2_decap_8 FILLER_25_1909 ();
 sg13g2_fill_2 FILLER_25_1916 ();
 sg13g2_fill_1 FILLER_25_1918 ();
 sg13g2_fill_1 FILLER_25_1924 ();
 sg13g2_fill_1 FILLER_25_1947 ();
 sg13g2_fill_2 FILLER_25_1961 ();
 sg13g2_fill_1 FILLER_25_2046 ();
 sg13g2_decap_8 FILLER_25_2079 ();
 sg13g2_decap_4 FILLER_25_2086 ();
 sg13g2_fill_1 FILLER_25_2090 ();
 sg13g2_fill_2 FILLER_25_2110 ();
 sg13g2_fill_1 FILLER_25_2117 ();
 sg13g2_fill_2 FILLER_25_2154 ();
 sg13g2_fill_1 FILLER_25_2156 ();
 sg13g2_fill_2 FILLER_25_2170 ();
 sg13g2_fill_1 FILLER_25_2172 ();
 sg13g2_decap_4 FILLER_25_2186 ();
 sg13g2_fill_1 FILLER_25_2190 ();
 sg13g2_fill_1 FILLER_25_2249 ();
 sg13g2_fill_2 FILLER_25_2262 ();
 sg13g2_decap_4 FILLER_25_2269 ();
 sg13g2_fill_1 FILLER_25_2273 ();
 sg13g2_decap_8 FILLER_25_2279 ();
 sg13g2_decap_4 FILLER_25_2286 ();
 sg13g2_decap_8 FILLER_25_2294 ();
 sg13g2_fill_2 FILLER_25_2301 ();
 sg13g2_fill_1 FILLER_25_2308 ();
 sg13g2_fill_2 FILLER_25_2364 ();
 sg13g2_fill_1 FILLER_25_2375 ();
 sg13g2_fill_1 FILLER_25_2422 ();
 sg13g2_fill_2 FILLER_25_2462 ();
 sg13g2_fill_2 FILLER_25_2468 ();
 sg13g2_decap_8 FILLER_25_2490 ();
 sg13g2_decap_8 FILLER_25_2497 ();
 sg13g2_fill_1 FILLER_25_2504 ();
 sg13g2_decap_8 FILLER_25_2531 ();
 sg13g2_fill_1 FILLER_25_2568 ();
 sg13g2_fill_2 FILLER_25_2584 ();
 sg13g2_fill_1 FILLER_25_2586 ();
 sg13g2_decap_4 FILLER_25_2609 ();
 sg13g2_fill_2 FILLER_25_2623 ();
 sg13g2_fill_2 FILLER_25_2630 ();
 sg13g2_fill_1 FILLER_25_2632 ();
 sg13g2_fill_2 FILLER_25_2653 ();
 sg13g2_decap_4 FILLER_25_2662 ();
 sg13g2_fill_1 FILLER_25_2666 ();
 sg13g2_fill_2 FILLER_25_2675 ();
 sg13g2_decap_8 FILLER_25_2705 ();
 sg13g2_fill_2 FILLER_25_2712 ();
 sg13g2_fill_1 FILLER_25_2714 ();
 sg13g2_fill_2 FILLER_25_2772 ();
 sg13g2_fill_2 FILLER_25_2782 ();
 sg13g2_fill_2 FILLER_25_2799 ();
 sg13g2_decap_4 FILLER_25_2806 ();
 sg13g2_fill_1 FILLER_25_2823 ();
 sg13g2_fill_1 FILLER_25_2855 ();
 sg13g2_fill_1 FILLER_25_2883 ();
 sg13g2_fill_1 FILLER_25_2901 ();
 sg13g2_fill_2 FILLER_25_2910 ();
 sg13g2_fill_1 FILLER_25_2912 ();
 sg13g2_decap_8 FILLER_25_2925 ();
 sg13g2_fill_2 FILLER_25_2948 ();
 sg13g2_fill_1 FILLER_25_2950 ();
 sg13g2_fill_1 FILLER_25_2959 ();
 sg13g2_fill_2 FILLER_25_2973 ();
 sg13g2_fill_1 FILLER_25_3049 ();
 sg13g2_fill_1 FILLER_25_3078 ();
 sg13g2_decap_8 FILLER_25_3103 ();
 sg13g2_fill_2 FILLER_25_3136 ();
 sg13g2_fill_2 FILLER_25_3146 ();
 sg13g2_fill_1 FILLER_25_3148 ();
 sg13g2_fill_1 FILLER_25_3158 ();
 sg13g2_fill_2 FILLER_25_3164 ();
 sg13g2_fill_2 FILLER_25_3179 ();
 sg13g2_fill_1 FILLER_25_3181 ();
 sg13g2_fill_1 FILLER_25_3217 ();
 sg13g2_fill_1 FILLER_25_3244 ();
 sg13g2_fill_1 FILLER_25_3250 ();
 sg13g2_fill_1 FILLER_25_3281 ();
 sg13g2_fill_2 FILLER_25_3291 ();
 sg13g2_decap_8 FILLER_25_3441 ();
 sg13g2_decap_8 FILLER_25_3448 ();
 sg13g2_decap_4 FILLER_25_3475 ();
 sg13g2_fill_1 FILLER_25_3479 ();
 sg13g2_decap_8 FILLER_25_3495 ();
 sg13g2_fill_2 FILLER_25_3515 ();
 sg13g2_decap_4 FILLER_25_3529 ();
 sg13g2_fill_2 FILLER_25_3533 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_4 ();
 sg13g2_decap_8 FILLER_26_10 ();
 sg13g2_fill_2 FILLER_26_37 ();
 sg13g2_fill_1 FILLER_26_39 ();
 sg13g2_fill_2 FILLER_26_64 ();
 sg13g2_fill_2 FILLER_26_108 ();
 sg13g2_fill_1 FILLER_26_123 ();
 sg13g2_decap_8 FILLER_26_160 ();
 sg13g2_fill_1 FILLER_26_167 ();
 sg13g2_fill_1 FILLER_26_205 ();
 sg13g2_fill_1 FILLER_26_220 ();
 sg13g2_fill_1 FILLER_26_240 ();
 sg13g2_fill_1 FILLER_26_302 ();
 sg13g2_fill_1 FILLER_26_309 ();
 sg13g2_fill_2 FILLER_26_342 ();
 sg13g2_fill_1 FILLER_26_344 ();
 sg13g2_fill_2 FILLER_26_493 ();
 sg13g2_fill_2 FILLER_26_614 ();
 sg13g2_fill_1 FILLER_26_1042 ();
 sg13g2_fill_1 FILLER_26_1126 ();
 sg13g2_fill_2 FILLER_26_1142 ();
 sg13g2_fill_1 FILLER_26_1169 ();
 sg13g2_fill_1 FILLER_26_1267 ();
 sg13g2_fill_1 FILLER_26_1296 ();
 sg13g2_fill_2 FILLER_26_1325 ();
 sg13g2_fill_1 FILLER_26_1349 ();
 sg13g2_fill_1 FILLER_26_1372 ();
 sg13g2_fill_2 FILLER_26_1386 ();
 sg13g2_decap_4 FILLER_26_1425 ();
 sg13g2_fill_1 FILLER_26_1429 ();
 sg13g2_fill_2 FILLER_26_1446 ();
 sg13g2_fill_2 FILLER_26_1456 ();
 sg13g2_fill_1 FILLER_26_1472 ();
 sg13g2_fill_2 FILLER_26_1505 ();
 sg13g2_fill_1 FILLER_26_1507 ();
 sg13g2_fill_2 FILLER_26_1524 ();
 sg13g2_fill_1 FILLER_26_1539 ();
 sg13g2_decap_8 FILLER_26_1544 ();
 sg13g2_decap_8 FILLER_26_1551 ();
 sg13g2_fill_1 FILLER_26_1558 ();
 sg13g2_fill_2 FILLER_26_1593 ();
 sg13g2_fill_1 FILLER_26_1595 ();
 sg13g2_fill_2 FILLER_26_1614 ();
 sg13g2_decap_4 FILLER_26_1622 ();
 sg13g2_fill_1 FILLER_26_1626 ();
 sg13g2_decap_4 FILLER_26_1645 ();
 sg13g2_fill_1 FILLER_26_1658 ();
 sg13g2_fill_1 FILLER_26_1663 ();
 sg13g2_fill_2 FILLER_26_1753 ();
 sg13g2_fill_2 FILLER_26_1760 ();
 sg13g2_fill_1 FILLER_26_1773 ();
 sg13g2_fill_1 FILLER_26_1778 ();
 sg13g2_fill_1 FILLER_26_1820 ();
 sg13g2_decap_4 FILLER_26_1826 ();
 sg13g2_fill_1 FILLER_26_1830 ();
 sg13g2_decap_4 FILLER_26_1839 ();
 sg13g2_fill_2 FILLER_26_1843 ();
 sg13g2_fill_1 FILLER_26_1854 ();
 sg13g2_fill_2 FILLER_26_1860 ();
 sg13g2_fill_1 FILLER_26_1862 ();
 sg13g2_decap_8 FILLER_26_1906 ();
 sg13g2_decap_8 FILLER_26_1913 ();
 sg13g2_fill_2 FILLER_26_1920 ();
 sg13g2_fill_1 FILLER_26_1922 ();
 sg13g2_fill_1 FILLER_26_1994 ();
 sg13g2_fill_2 FILLER_26_2000 ();
 sg13g2_fill_1 FILLER_26_2011 ();
 sg13g2_fill_2 FILLER_26_2033 ();
 sg13g2_fill_2 FILLER_26_2079 ();
 sg13g2_fill_1 FILLER_26_2107 ();
 sg13g2_fill_2 FILLER_26_2144 ();
 sg13g2_fill_1 FILLER_26_2146 ();
 sg13g2_decap_8 FILLER_26_2160 ();
 sg13g2_fill_1 FILLER_26_2167 ();
 sg13g2_fill_1 FILLER_26_2213 ();
 sg13g2_decap_4 FILLER_26_2227 ();
 sg13g2_fill_2 FILLER_26_2231 ();
 sg13g2_decap_8 FILLER_26_2237 ();
 sg13g2_decap_8 FILLER_26_2244 ();
 sg13g2_fill_2 FILLER_26_2251 ();
 sg13g2_fill_2 FILLER_26_2294 ();
 sg13g2_fill_1 FILLER_26_2296 ();
 sg13g2_fill_1 FILLER_26_2305 ();
 sg13g2_fill_2 FILLER_26_2324 ();
 sg13g2_fill_1 FILLER_26_2347 ();
 sg13g2_fill_1 FILLER_26_2362 ();
 sg13g2_fill_2 FILLER_26_2398 ();
 sg13g2_fill_1 FILLER_26_2400 ();
 sg13g2_fill_2 FILLER_26_2414 ();
 sg13g2_fill_2 FILLER_26_2442 ();
 sg13g2_fill_2 FILLER_26_2466 ();
 sg13g2_fill_2 FILLER_26_2481 ();
 sg13g2_fill_1 FILLER_26_2516 ();
 sg13g2_fill_1 FILLER_26_2566 ();
 sg13g2_decap_8 FILLER_26_2575 ();
 sg13g2_fill_1 FILLER_26_2582 ();
 sg13g2_fill_2 FILLER_26_2588 ();
 sg13g2_fill_1 FILLER_26_2590 ();
 sg13g2_fill_2 FILLER_26_2599 ();
 sg13g2_fill_1 FILLER_26_2625 ();
 sg13g2_fill_1 FILLER_26_2639 ();
 sg13g2_decap_4 FILLER_26_2650 ();
 sg13g2_fill_1 FILLER_26_2660 ();
 sg13g2_fill_1 FILLER_26_2665 ();
 sg13g2_fill_2 FILLER_26_2692 ();
 sg13g2_fill_2 FILLER_26_2743 ();
 sg13g2_fill_2 FILLER_26_2779 ();
 sg13g2_fill_2 FILLER_26_2793 ();
 sg13g2_fill_1 FILLER_26_2814 ();
 sg13g2_fill_2 FILLER_26_2832 ();
 sg13g2_fill_1 FILLER_26_2834 ();
 sg13g2_fill_1 FILLER_26_2840 ();
 sg13g2_decap_8 FILLER_26_2848 ();
 sg13g2_fill_2 FILLER_26_2873 ();
 sg13g2_fill_1 FILLER_26_2875 ();
 sg13g2_fill_2 FILLER_26_2891 ();
 sg13g2_fill_2 FILLER_26_2927 ();
 sg13g2_decap_4 FILLER_26_2942 ();
 sg13g2_fill_2 FILLER_26_2974 ();
 sg13g2_fill_2 FILLER_26_3096 ();
 sg13g2_fill_1 FILLER_26_3098 ();
 sg13g2_decap_4 FILLER_26_3114 ();
 sg13g2_fill_1 FILLER_26_3118 ();
 sg13g2_fill_2 FILLER_26_3126 ();
 sg13g2_fill_1 FILLER_26_3128 ();
 sg13g2_fill_1 FILLER_26_3137 ();
 sg13g2_fill_1 FILLER_26_3171 ();
 sg13g2_fill_2 FILLER_26_3198 ();
 sg13g2_fill_2 FILLER_26_3245 ();
 sg13g2_fill_2 FILLER_26_3257 ();
 sg13g2_fill_1 FILLER_26_3259 ();
 sg13g2_fill_1 FILLER_26_3307 ();
 sg13g2_fill_1 FILLER_26_3331 ();
 sg13g2_fill_1 FILLER_26_3419 ();
 sg13g2_fill_1 FILLER_26_3453 ();
 sg13g2_fill_1 FILLER_26_3459 ();
 sg13g2_fill_2 FILLER_26_3477 ();
 sg13g2_fill_1 FILLER_26_3479 ();
 sg13g2_decap_4 FILLER_26_3493 ();
 sg13g2_fill_2 FILLER_26_3497 ();
 sg13g2_fill_2 FILLER_26_3517 ();
 sg13g2_decap_8 FILLER_26_3538 ();
 sg13g2_fill_1 FILLER_26_3545 ();
 sg13g2_fill_2 FILLER_26_3554 ();
 sg13g2_fill_2 FILLER_26_3577 ();
 sg13g2_fill_1 FILLER_26_3579 ();
 sg13g2_fill_1 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_42 ();
 sg13g2_decap_4 FILLER_27_60 ();
 sg13g2_fill_1 FILLER_27_115 ();
 sg13g2_fill_2 FILLER_27_199 ();
 sg13g2_fill_1 FILLER_27_201 ();
 sg13g2_fill_2 FILLER_27_240 ();
 sg13g2_fill_1 FILLER_27_282 ();
 sg13g2_fill_1 FILLER_27_313 ();
 sg13g2_fill_1 FILLER_27_385 ();
 sg13g2_decap_4 FILLER_27_442 ();
 sg13g2_fill_2 FILLER_27_446 ();
 sg13g2_fill_2 FILLER_27_456 ();
 sg13g2_fill_2 FILLER_27_492 ();
 sg13g2_fill_1 FILLER_27_494 ();
 sg13g2_fill_1 FILLER_27_517 ();
 sg13g2_fill_2 FILLER_27_634 ();
 sg13g2_decap_4 FILLER_27_646 ();
 sg13g2_fill_2 FILLER_27_650 ();
 sg13g2_fill_2 FILLER_27_791 ();
 sg13g2_fill_2 FILLER_27_909 ();
 sg13g2_fill_1 FILLER_27_917 ();
 sg13g2_fill_2 FILLER_27_924 ();
 sg13g2_fill_1 FILLER_27_926 ();
 sg13g2_fill_2 FILLER_27_1060 ();
 sg13g2_fill_1 FILLER_27_1062 ();
 sg13g2_fill_2 FILLER_27_1098 ();
 sg13g2_fill_1 FILLER_27_1100 ();
 sg13g2_fill_2 FILLER_27_1111 ();
 sg13g2_fill_1 FILLER_27_1113 ();
 sg13g2_fill_1 FILLER_27_1178 ();
 sg13g2_fill_2 FILLER_27_1191 ();
 sg13g2_fill_1 FILLER_27_1212 ();
 sg13g2_fill_1 FILLER_27_1241 ();
 sg13g2_fill_1 FILLER_27_1251 ();
 sg13g2_fill_2 FILLER_27_1287 ();
 sg13g2_fill_2 FILLER_27_1294 ();
 sg13g2_fill_2 FILLER_27_1308 ();
 sg13g2_decap_4 FILLER_27_1324 ();
 sg13g2_fill_1 FILLER_27_1328 ();
 sg13g2_fill_2 FILLER_27_1334 ();
 sg13g2_fill_1 FILLER_27_1336 ();
 sg13g2_fill_1 FILLER_27_1350 ();
 sg13g2_decap_4 FILLER_27_1361 ();
 sg13g2_fill_1 FILLER_27_1365 ();
 sg13g2_decap_4 FILLER_27_1378 ();
 sg13g2_fill_2 FILLER_27_1382 ();
 sg13g2_fill_2 FILLER_27_1392 ();
 sg13g2_fill_2 FILLER_27_1407 ();
 sg13g2_decap_8 FILLER_27_1427 ();
 sg13g2_fill_2 FILLER_27_1434 ();
 sg13g2_fill_1 FILLER_27_1436 ();
 sg13g2_fill_1 FILLER_27_1441 ();
 sg13g2_fill_2 FILLER_27_1447 ();
 sg13g2_fill_2 FILLER_27_1477 ();
 sg13g2_fill_1 FILLER_27_1479 ();
 sg13g2_fill_2 FILLER_27_1511 ();
 sg13g2_fill_2 FILLER_27_1521 ();
 sg13g2_fill_1 FILLER_27_1537 ();
 sg13g2_fill_2 FILLER_27_1558 ();
 sg13g2_fill_2 FILLER_27_1583 ();
 sg13g2_fill_2 FILLER_27_1593 ();
 sg13g2_decap_4 FILLER_27_1612 ();
 sg13g2_fill_2 FILLER_27_1616 ();
 sg13g2_decap_8 FILLER_27_1639 ();
 sg13g2_decap_8 FILLER_27_1646 ();
 sg13g2_fill_2 FILLER_27_1653 ();
 sg13g2_fill_2 FILLER_27_1660 ();
 sg13g2_decap_4 FILLER_27_1683 ();
 sg13g2_decap_4 FILLER_27_1691 ();
 sg13g2_decap_4 FILLER_27_1703 ();
 sg13g2_fill_1 FILLER_27_1707 ();
 sg13g2_fill_2 FILLER_27_1712 ();
 sg13g2_fill_1 FILLER_27_1714 ();
 sg13g2_fill_1 FILLER_27_1731 ();
 sg13g2_fill_1 FILLER_27_1736 ();
 sg13g2_fill_2 FILLER_27_1764 ();
 sg13g2_fill_1 FILLER_27_1766 ();
 sg13g2_fill_2 FILLER_27_1801 ();
 sg13g2_decap_4 FILLER_27_1816 ();
 sg13g2_decap_8 FILLER_27_1832 ();
 sg13g2_decap_4 FILLER_27_1839 ();
 sg13g2_fill_1 FILLER_27_1843 ();
 sg13g2_fill_2 FILLER_27_1884 ();
 sg13g2_decap_8 FILLER_27_1915 ();
 sg13g2_fill_2 FILLER_27_1922 ();
 sg13g2_fill_1 FILLER_27_1924 ();
 sg13g2_fill_2 FILLER_27_1940 ();
 sg13g2_fill_1 FILLER_27_1942 ();
 sg13g2_fill_1 FILLER_27_1957 ();
 sg13g2_fill_1 FILLER_27_1985 ();
 sg13g2_fill_1 FILLER_27_2021 ();
 sg13g2_fill_1 FILLER_27_2078 ();
 sg13g2_decap_4 FILLER_27_2120 ();
 sg13g2_fill_2 FILLER_27_2124 ();
 sg13g2_decap_4 FILLER_27_2139 ();
 sg13g2_fill_1 FILLER_27_2143 ();
 sg13g2_decap_4 FILLER_27_2165 ();
 sg13g2_fill_2 FILLER_27_2169 ();
 sg13g2_fill_2 FILLER_27_2191 ();
 sg13g2_fill_1 FILLER_27_2193 ();
 sg13g2_fill_1 FILLER_27_2211 ();
 sg13g2_fill_1 FILLER_27_2240 ();
 sg13g2_decap_4 FILLER_27_2249 ();
 sg13g2_fill_1 FILLER_27_2258 ();
 sg13g2_fill_2 FILLER_27_2267 ();
 sg13g2_decap_4 FILLER_27_2279 ();
 sg13g2_fill_1 FILLER_27_2283 ();
 sg13g2_fill_2 FILLER_27_2314 ();
 sg13g2_fill_1 FILLER_27_2316 ();
 sg13g2_fill_2 FILLER_27_2352 ();
 sg13g2_decap_4 FILLER_27_2396 ();
 sg13g2_fill_2 FILLER_27_2400 ();
 sg13g2_fill_1 FILLER_27_2437 ();
 sg13g2_fill_1 FILLER_27_2451 ();
 sg13g2_fill_1 FILLER_27_2462 ();
 sg13g2_fill_1 FILLER_27_2476 ();
 sg13g2_fill_1 FILLER_27_2487 ();
 sg13g2_fill_2 FILLER_27_2492 ();
 sg13g2_fill_1 FILLER_27_2494 ();
 sg13g2_decap_4 FILLER_27_2508 ();
 sg13g2_fill_1 FILLER_27_2512 ();
 sg13g2_fill_1 FILLER_27_2521 ();
 sg13g2_fill_2 FILLER_27_2526 ();
 sg13g2_fill_1 FILLER_27_2528 ();
 sg13g2_fill_1 FILLER_27_2538 ();
 sg13g2_fill_2 FILLER_27_2572 ();
 sg13g2_fill_1 FILLER_27_2574 ();
 sg13g2_fill_2 FILLER_27_2607 ();
 sg13g2_fill_2 FILLER_27_2632 ();
 sg13g2_fill_1 FILLER_27_2642 ();
 sg13g2_decap_4 FILLER_27_2663 ();
 sg13g2_fill_2 FILLER_27_2667 ();
 sg13g2_fill_1 FILLER_27_2679 ();
 sg13g2_fill_2 FILLER_27_2721 ();
 sg13g2_fill_1 FILLER_27_2774 ();
 sg13g2_fill_1 FILLER_27_2788 ();
 sg13g2_decap_8 FILLER_27_2803 ();
 sg13g2_fill_2 FILLER_27_2832 ();
 sg13g2_fill_1 FILLER_27_2834 ();
 sg13g2_fill_2 FILLER_27_2886 ();
 sg13g2_fill_1 FILLER_27_2888 ();
 sg13g2_fill_2 FILLER_27_2907 ();
 sg13g2_fill_1 FILLER_27_2909 ();
 sg13g2_fill_2 FILLER_27_2923 ();
 sg13g2_fill_2 FILLER_27_2983 ();
 sg13g2_fill_2 FILLER_27_2990 ();
 sg13g2_fill_1 FILLER_27_2992 ();
 sg13g2_fill_1 FILLER_27_2998 ();
 sg13g2_fill_2 FILLER_27_3018 ();
 sg13g2_fill_2 FILLER_27_3024 ();
 sg13g2_fill_1 FILLER_27_3057 ();
 sg13g2_fill_2 FILLER_27_3084 ();
 sg13g2_fill_1 FILLER_27_3086 ();
 sg13g2_fill_1 FILLER_27_3122 ();
 sg13g2_fill_2 FILLER_27_3145 ();
 sg13g2_fill_1 FILLER_27_3147 ();
 sg13g2_fill_2 FILLER_27_3156 ();
 sg13g2_fill_1 FILLER_27_3158 ();
 sg13g2_fill_2 FILLER_27_3173 ();
 sg13g2_fill_1 FILLER_27_3200 ();
 sg13g2_fill_1 FILLER_27_3244 ();
 sg13g2_fill_1 FILLER_27_3364 ();
 sg13g2_fill_2 FILLER_27_3389 ();
 sg13g2_fill_2 FILLER_27_3430 ();
 sg13g2_fill_1 FILLER_27_3432 ();
 sg13g2_fill_2 FILLER_27_3437 ();
 sg13g2_decap_4 FILLER_27_3453 ();
 sg13g2_decap_8 FILLER_27_3468 ();
 sg13g2_decap_4 FILLER_27_3475 ();
 sg13g2_fill_2 FILLER_27_3479 ();
 sg13g2_decap_4 FILLER_27_3486 ();
 sg13g2_fill_1 FILLER_27_3490 ();
 sg13g2_fill_1 FILLER_27_3501 ();
 sg13g2_decap_4 FILLER_27_3511 ();
 sg13g2_fill_1 FILLER_27_3541 ();
 sg13g2_fill_1 FILLER_27_3546 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_2 ();
 sg13g2_decap_4 FILLER_28_57 ();
 sg13g2_fill_2 FILLER_28_76 ();
 sg13g2_fill_1 FILLER_28_78 ();
 sg13g2_fill_1 FILLER_28_87 ();
 sg13g2_fill_2 FILLER_28_149 ();
 sg13g2_fill_1 FILLER_28_179 ();
 sg13g2_fill_1 FILLER_28_225 ();
 sg13g2_fill_2 FILLER_28_251 ();
 sg13g2_fill_1 FILLER_28_253 ();
 sg13g2_decap_4 FILLER_28_278 ();
 sg13g2_fill_1 FILLER_28_282 ();
 sg13g2_fill_1 FILLER_28_286 ();
 sg13g2_fill_2 FILLER_28_305 ();
 sg13g2_fill_2 FILLER_28_351 ();
 sg13g2_fill_2 FILLER_28_385 ();
 sg13g2_fill_1 FILLER_28_403 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_fill_1 FILLER_28_426 ();
 sg13g2_decap_4 FILLER_28_436 ();
 sg13g2_fill_1 FILLER_28_440 ();
 sg13g2_fill_1 FILLER_28_474 ();
 sg13g2_fill_2 FILLER_28_497 ();
 sg13g2_fill_1 FILLER_28_538 ();
 sg13g2_fill_2 FILLER_28_595 ();
 sg13g2_fill_2 FILLER_28_632 ();
 sg13g2_fill_1 FILLER_28_634 ();
 sg13g2_fill_2 FILLER_28_690 ();
 sg13g2_fill_2 FILLER_28_735 ();
 sg13g2_fill_2 FILLER_28_821 ();
 sg13g2_fill_2 FILLER_28_860 ();
 sg13g2_fill_2 FILLER_28_875 ();
 sg13g2_fill_1 FILLER_28_911 ();
 sg13g2_fill_1 FILLER_28_918 ();
 sg13g2_fill_1 FILLER_28_962 ();
 sg13g2_fill_1 FILLER_28_1014 ();
 sg13g2_fill_1 FILLER_28_1052 ();
 sg13g2_fill_2 FILLER_28_1062 ();
 sg13g2_fill_2 FILLER_28_1105 ();
 sg13g2_fill_1 FILLER_28_1152 ();
 sg13g2_fill_2 FILLER_28_1189 ();
 sg13g2_fill_2 FILLER_28_1288 ();
 sg13g2_fill_1 FILLER_28_1290 ();
 sg13g2_fill_2 FILLER_28_1297 ();
 sg13g2_fill_2 FILLER_28_1312 ();
 sg13g2_fill_2 FILLER_28_1319 ();
 sg13g2_fill_2 FILLER_28_1350 ();
 sg13g2_fill_1 FILLER_28_1392 ();
 sg13g2_decap_8 FILLER_28_1438 ();
 sg13g2_decap_8 FILLER_28_1445 ();
 sg13g2_fill_2 FILLER_28_1452 ();
 sg13g2_fill_1 FILLER_28_1520 ();
 sg13g2_decap_8 FILLER_28_1526 ();
 sg13g2_fill_2 FILLER_28_1533 ();
 sg13g2_fill_2 FILLER_28_1579 ();
 sg13g2_fill_2 FILLER_28_1586 ();
 sg13g2_fill_1 FILLER_28_1598 ();
 sg13g2_fill_2 FILLER_28_1612 ();
 sg13g2_fill_1 FILLER_28_1614 ();
 sg13g2_decap_8 FILLER_28_1635 ();
 sg13g2_fill_1 FILLER_28_1642 ();
 sg13g2_fill_1 FILLER_28_1679 ();
 sg13g2_decap_4 FILLER_28_1697 ();
 sg13g2_fill_1 FILLER_28_1701 ();
 sg13g2_fill_1 FILLER_28_1714 ();
 sg13g2_decap_4 FILLER_28_1742 ();
 sg13g2_fill_2 FILLER_28_1763 ();
 sg13g2_fill_2 FILLER_28_1770 ();
 sg13g2_fill_1 FILLER_28_1772 ();
 sg13g2_fill_2 FILLER_28_1801 ();
 sg13g2_fill_1 FILLER_28_1803 ();
 sg13g2_fill_1 FILLER_28_1814 ();
 sg13g2_fill_2 FILLER_28_1827 ();
 sg13g2_fill_1 FILLER_28_1829 ();
 sg13g2_fill_2 FILLER_28_1837 ();
 sg13g2_fill_1 FILLER_28_1839 ();
 sg13g2_fill_1 FILLER_28_1896 ();
 sg13g2_fill_1 FILLER_28_1912 ();
 sg13g2_fill_2 FILLER_28_1933 ();
 sg13g2_fill_2 FILLER_28_1939 ();
 sg13g2_fill_2 FILLER_28_1951 ();
 sg13g2_fill_1 FILLER_28_1953 ();
 sg13g2_fill_1 FILLER_28_1972 ();
 sg13g2_fill_2 FILLER_28_1981 ();
 sg13g2_fill_2 FILLER_28_1988 ();
 sg13g2_fill_1 FILLER_28_1990 ();
 sg13g2_fill_1 FILLER_28_2024 ();
 sg13g2_fill_1 FILLER_28_2034 ();
 sg13g2_fill_2 FILLER_28_2044 ();
 sg13g2_fill_1 FILLER_28_2096 ();
 sg13g2_fill_2 FILLER_28_2111 ();
 sg13g2_fill_2 FILLER_28_2173 ();
 sg13g2_fill_2 FILLER_28_2183 ();
 sg13g2_fill_1 FILLER_28_2185 ();
 sg13g2_fill_2 FILLER_28_2203 ();
 sg13g2_decap_8 FILLER_28_2223 ();
 sg13g2_fill_2 FILLER_28_2230 ();
 sg13g2_fill_2 FILLER_28_2252 ();
 sg13g2_fill_1 FILLER_28_2266 ();
 sg13g2_decap_8 FILLER_28_2274 ();
 sg13g2_decap_8 FILLER_28_2285 ();
 sg13g2_fill_2 FILLER_28_2292 ();
 sg13g2_fill_1 FILLER_28_2294 ();
 sg13g2_fill_2 FILLER_28_2308 ();
 sg13g2_decap_4 FILLER_28_2320 ();
 sg13g2_fill_2 FILLER_28_2324 ();
 sg13g2_decap_4 FILLER_28_2338 ();
 sg13g2_decap_8 FILLER_28_2354 ();
 sg13g2_decap_8 FILLER_28_2361 ();
 sg13g2_fill_1 FILLER_28_2368 ();
 sg13g2_fill_1 FILLER_28_2379 ();
 sg13g2_fill_2 FILLER_28_2405 ();
 sg13g2_fill_1 FILLER_28_2420 ();
 sg13g2_fill_2 FILLER_28_2453 ();
 sg13g2_fill_1 FILLER_28_2488 ();
 sg13g2_fill_1 FILLER_28_2516 ();
 sg13g2_decap_4 FILLER_28_2579 ();
 sg13g2_fill_2 FILLER_28_2583 ();
 sg13g2_fill_1 FILLER_28_2602 ();
 sg13g2_fill_1 FILLER_28_2623 ();
 sg13g2_fill_1 FILLER_28_2649 ();
 sg13g2_fill_2 FILLER_28_2691 ();
 sg13g2_fill_2 FILLER_28_2715 ();
 sg13g2_fill_2 FILLER_28_2726 ();
 sg13g2_fill_2 FILLER_28_2758 ();
 sg13g2_decap_4 FILLER_28_2809 ();
 sg13g2_fill_2 FILLER_28_2826 ();
 sg13g2_fill_1 FILLER_28_2841 ();
 sg13g2_fill_2 FILLER_28_2883 ();
 sg13g2_fill_2 FILLER_28_2926 ();
 sg13g2_fill_1 FILLER_28_2928 ();
 sg13g2_fill_2 FILLER_28_3018 ();
 sg13g2_fill_2 FILLER_28_3069 ();
 sg13g2_fill_1 FILLER_28_3071 ();
 sg13g2_fill_1 FILLER_28_3159 ();
 sg13g2_decap_8 FILLER_28_3188 ();
 sg13g2_fill_2 FILLER_28_3208 ();
 sg13g2_fill_1 FILLER_28_3210 ();
 sg13g2_fill_1 FILLER_28_3239 ();
 sg13g2_fill_2 FILLER_28_3318 ();
 sg13g2_fill_1 FILLER_28_3320 ();
 sg13g2_fill_1 FILLER_28_3383 ();
 sg13g2_fill_2 FILLER_28_3420 ();
 sg13g2_fill_1 FILLER_28_3434 ();
 sg13g2_decap_4 FILLER_28_3482 ();
 sg13g2_decap_8 FILLER_28_3513 ();
 sg13g2_fill_1 FILLER_28_3520 ();
 sg13g2_fill_1 FILLER_28_3526 ();
 sg13g2_decap_4 FILLER_28_3540 ();
 sg13g2_fill_1 FILLER_28_3570 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_38 ();
 sg13g2_fill_1 FILLER_29_40 ();
 sg13g2_fill_2 FILLER_29_59 ();
 sg13g2_fill_2 FILLER_29_80 ();
 sg13g2_fill_1 FILLER_29_82 ();
 sg13g2_fill_2 FILLER_29_96 ();
 sg13g2_fill_2 FILLER_29_103 ();
 sg13g2_fill_1 FILLER_29_105 ();
 sg13g2_fill_2 FILLER_29_156 ();
 sg13g2_fill_2 FILLER_29_176 ();
 sg13g2_fill_1 FILLER_29_178 ();
 sg13g2_fill_1 FILLER_29_269 ();
 sg13g2_fill_2 FILLER_29_280 ();
 sg13g2_fill_2 FILLER_29_285 ();
 sg13g2_fill_2 FILLER_29_291 ();
 sg13g2_fill_1 FILLER_29_293 ();
 sg13g2_decap_4 FILLER_29_302 ();
 sg13g2_decap_4 FILLER_29_309 ();
 sg13g2_fill_2 FILLER_29_351 ();
 sg13g2_fill_2 FILLER_29_362 ();
 sg13g2_fill_1 FILLER_29_394 ();
 sg13g2_fill_2 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_420 ();
 sg13g2_fill_1 FILLER_29_478 ();
 sg13g2_fill_1 FILLER_29_492 ();
 sg13g2_fill_2 FILLER_29_507 ();
 sg13g2_fill_2 FILLER_29_521 ();
 sg13g2_fill_2 FILLER_29_532 ();
 sg13g2_fill_2 FILLER_29_570 ();
 sg13g2_fill_1 FILLER_29_572 ();
 sg13g2_fill_1 FILLER_29_643 ();
 sg13g2_fill_2 FILLER_29_666 ();
 sg13g2_fill_1 FILLER_29_714 ();
 sg13g2_fill_2 FILLER_29_726 ();
 sg13g2_fill_1 FILLER_29_812 ();
 sg13g2_fill_1 FILLER_29_829 ();
 sg13g2_fill_2 FILLER_29_876 ();
 sg13g2_fill_1 FILLER_29_878 ();
 sg13g2_fill_1 FILLER_29_902 ();
 sg13g2_fill_1 FILLER_29_972 ();
 sg13g2_fill_1 FILLER_29_1070 ();
 sg13g2_decap_8 FILLER_29_1103 ();
 sg13g2_decap_4 FILLER_29_1110 ();
 sg13g2_fill_1 FILLER_29_1114 ();
 sg13g2_fill_1 FILLER_29_1119 ();
 sg13g2_fill_2 FILLER_29_1133 ();
 sg13g2_fill_2 FILLER_29_1176 ();
 sg13g2_decap_4 FILLER_29_1211 ();
 sg13g2_fill_2 FILLER_29_1228 ();
 sg13g2_fill_2 FILLER_29_1258 ();
 sg13g2_fill_2 FILLER_29_1289 ();
 sg13g2_fill_1 FILLER_29_1291 ();
 sg13g2_fill_2 FILLER_29_1297 ();
 sg13g2_fill_2 FILLER_29_1309 ();
 sg13g2_decap_8 FILLER_29_1320 ();
 sg13g2_fill_2 FILLER_29_1335 ();
 sg13g2_decap_8 FILLER_29_1369 ();
 sg13g2_decap_4 FILLER_29_1376 ();
 sg13g2_fill_2 FILLER_29_1380 ();
 sg13g2_decap_4 FILLER_29_1387 ();
 sg13g2_decap_8 FILLER_29_1396 ();
 sg13g2_fill_2 FILLER_29_1403 ();
 sg13g2_fill_1 FILLER_29_1405 ();
 sg13g2_fill_1 FILLER_29_1453 ();
 sg13g2_fill_2 FILLER_29_1486 ();
 sg13g2_decap_4 FILLER_29_1505 ();
 sg13g2_fill_2 FILLER_29_1517 ();
 sg13g2_fill_1 FILLER_29_1519 ();
 sg13g2_decap_8 FILLER_29_1525 ();
 sg13g2_decap_4 FILLER_29_1532 ();
 sg13g2_decap_8 FILLER_29_1554 ();
 sg13g2_fill_2 FILLER_29_1561 ();
 sg13g2_fill_2 FILLER_29_1587 ();
 sg13g2_fill_1 FILLER_29_1621 ();
 sg13g2_fill_2 FILLER_29_1635 ();
 sg13g2_fill_2 FILLER_29_1650 ();
 sg13g2_fill_2 FILLER_29_1689 ();
 sg13g2_fill_2 FILLER_29_1728 ();
 sg13g2_fill_1 FILLER_29_1730 ();
 sg13g2_fill_2 FILLER_29_1743 ();
 sg13g2_fill_1 FILLER_29_1745 ();
 sg13g2_fill_1 FILLER_29_1755 ();
 sg13g2_fill_2 FILLER_29_1780 ();
 sg13g2_fill_2 FILLER_29_1817 ();
 sg13g2_fill_1 FILLER_29_1819 ();
 sg13g2_decap_4 FILLER_29_1829 ();
 sg13g2_fill_2 FILLER_29_1846 ();
 sg13g2_decap_4 FILLER_29_1853 ();
 sg13g2_fill_2 FILLER_29_1874 ();
 sg13g2_decap_4 FILLER_29_1893 ();
 sg13g2_fill_2 FILLER_29_1915 ();
 sg13g2_fill_2 FILLER_29_1931 ();
 sg13g2_fill_2 FILLER_29_1946 ();
 sg13g2_fill_1 FILLER_29_1948 ();
 sg13g2_fill_2 FILLER_29_1968 ();
 sg13g2_decap_4 FILLER_29_1989 ();
 sg13g2_fill_1 FILLER_29_2037 ();
 sg13g2_fill_2 FILLER_29_2061 ();
 sg13g2_fill_1 FILLER_29_2063 ();
 sg13g2_fill_2 FILLER_29_2077 ();
 sg13g2_decap_8 FILLER_29_2092 ();
 sg13g2_fill_2 FILLER_29_2104 ();
 sg13g2_fill_2 FILLER_29_2119 ();
 sg13g2_fill_1 FILLER_29_2121 ();
 sg13g2_fill_1 FILLER_29_2148 ();
 sg13g2_fill_2 FILLER_29_2178 ();
 sg13g2_fill_2 FILLER_29_2201 ();
 sg13g2_fill_1 FILLER_29_2236 ();
 sg13g2_fill_1 FILLER_29_2253 ();
 sg13g2_decap_8 FILLER_29_2266 ();
 sg13g2_fill_2 FILLER_29_2273 ();
 sg13g2_fill_1 FILLER_29_2275 ();
 sg13g2_decap_4 FILLER_29_2304 ();
 sg13g2_decap_4 FILLER_29_2328 ();
 sg13g2_fill_2 FILLER_29_2332 ();
 sg13g2_decap_4 FILLER_29_2338 ();
 sg13g2_decap_8 FILLER_29_2359 ();
 sg13g2_decap_8 FILLER_29_2370 ();
 sg13g2_decap_4 FILLER_29_2382 ();
 sg13g2_decap_8 FILLER_29_2417 ();
 sg13g2_fill_1 FILLER_29_2424 ();
 sg13g2_fill_2 FILLER_29_2447 ();
 sg13g2_fill_2 FILLER_29_2459 ();
 sg13g2_fill_1 FILLER_29_2461 ();
 sg13g2_fill_2 FILLER_29_2515 ();
 sg13g2_fill_1 FILLER_29_2522 ();
 sg13g2_fill_2 FILLER_29_2551 ();
 sg13g2_fill_1 FILLER_29_2553 ();
 sg13g2_fill_1 FILLER_29_2582 ();
 sg13g2_fill_1 FILLER_29_2588 ();
 sg13g2_fill_1 FILLER_29_2601 ();
 sg13g2_fill_1 FILLER_29_2611 ();
 sg13g2_fill_1 FILLER_29_2667 ();
 sg13g2_decap_4 FILLER_29_2677 ();
 sg13g2_fill_2 FILLER_29_2681 ();
 sg13g2_fill_2 FILLER_29_2788 ();
 sg13g2_fill_2 FILLER_29_2850 ();
 sg13g2_fill_1 FILLER_29_2852 ();
 sg13g2_fill_1 FILLER_29_2883 ();
 sg13g2_fill_2 FILLER_29_2901 ();
 sg13g2_fill_1 FILLER_29_2912 ();
 sg13g2_fill_1 FILLER_29_2964 ();
 sg13g2_fill_2 FILLER_29_2987 ();
 sg13g2_fill_1 FILLER_29_2989 ();
 sg13g2_fill_1 FILLER_29_3003 ();
 sg13g2_fill_1 FILLER_29_3128 ();
 sg13g2_fill_1 FILLER_29_3164 ();
 sg13g2_fill_2 FILLER_29_3193 ();
 sg13g2_fill_2 FILLER_29_3208 ();
 sg13g2_fill_1 FILLER_29_3210 ();
 sg13g2_fill_1 FILLER_29_3229 ();
 sg13g2_fill_2 FILLER_29_3276 ();
 sg13g2_fill_1 FILLER_29_3328 ();
 sg13g2_fill_2 FILLER_29_3374 ();
 sg13g2_fill_1 FILLER_29_3445 ();
 sg13g2_fill_2 FILLER_29_3454 ();
 sg13g2_fill_1 FILLER_29_3456 ();
 sg13g2_decap_4 FILLER_29_3468 ();
 sg13g2_fill_1 FILLER_29_3472 ();
 sg13g2_fill_1 FILLER_29_3478 ();
 sg13g2_fill_2 FILLER_29_3489 ();
 sg13g2_decap_4 FILLER_29_3500 ();
 sg13g2_fill_1 FILLER_29_3504 ();
 sg13g2_decap_4 FILLER_29_3515 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_26 ();
 sg13g2_fill_2 FILLER_30_43 ();
 sg13g2_fill_1 FILLER_30_45 ();
 sg13g2_fill_2 FILLER_30_63 ();
 sg13g2_fill_1 FILLER_30_72 ();
 sg13g2_fill_2 FILLER_30_79 ();
 sg13g2_fill_2 FILLER_30_119 ();
 sg13g2_fill_1 FILLER_30_121 ();
 sg13g2_fill_2 FILLER_30_141 ();
 sg13g2_fill_1 FILLER_30_153 ();
 sg13g2_fill_2 FILLER_30_187 ();
 sg13g2_fill_2 FILLER_30_199 ();
 sg13g2_fill_1 FILLER_30_201 ();
 sg13g2_fill_1 FILLER_30_235 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_fill_2 FILLER_30_261 ();
 sg13g2_fill_1 FILLER_30_263 ();
 sg13g2_decap_4 FILLER_30_297 ();
 sg13g2_fill_1 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_357 ();
 sg13g2_fill_2 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_30_430 ();
 sg13g2_decap_4 FILLER_30_437 ();
 sg13g2_fill_1 FILLER_30_441 ();
 sg13g2_fill_2 FILLER_30_487 ();
 sg13g2_fill_2 FILLER_30_552 ();
 sg13g2_fill_1 FILLER_30_554 ();
 sg13g2_fill_2 FILLER_30_623 ();
 sg13g2_fill_1 FILLER_30_625 ();
 sg13g2_fill_1 FILLER_30_639 ();
 sg13g2_decap_4 FILLER_30_652 ();
 sg13g2_decap_4 FILLER_30_695 ();
 sg13g2_fill_2 FILLER_30_699 ();
 sg13g2_fill_1 FILLER_30_729 ();
 sg13g2_fill_2 FILLER_30_743 ();
 sg13g2_decap_4 FILLER_30_805 ();
 sg13g2_fill_2 FILLER_30_923 ();
 sg13g2_fill_1 FILLER_30_925 ();
 sg13g2_fill_2 FILLER_30_958 ();
 sg13g2_fill_1 FILLER_30_1002 ();
 sg13g2_fill_1 FILLER_30_1021 ();
 sg13g2_fill_2 FILLER_30_1057 ();
 sg13g2_fill_1 FILLER_30_1059 ();
 sg13g2_fill_2 FILLER_30_1082 ();
 sg13g2_fill_1 FILLER_30_1084 ();
 sg13g2_fill_2 FILLER_30_1093 ();
 sg13g2_decap_4 FILLER_30_1120 ();
 sg13g2_fill_2 FILLER_30_1124 ();
 sg13g2_decap_4 FILLER_30_1147 ();
 sg13g2_fill_2 FILLER_30_1185 ();
 sg13g2_fill_2 FILLER_30_1228 ();
 sg13g2_fill_1 FILLER_30_1244 ();
 sg13g2_fill_2 FILLER_30_1260 ();
 sg13g2_fill_1 FILLER_30_1279 ();
 sg13g2_fill_2 FILLER_30_1335 ();
 sg13g2_fill_2 FILLER_30_1378 ();
 sg13g2_decap_4 FILLER_30_1390 ();
 sg13g2_fill_1 FILLER_30_1394 ();
 sg13g2_fill_1 FILLER_30_1403 ();
 sg13g2_fill_2 FILLER_30_1417 ();
 sg13g2_fill_1 FILLER_30_1419 ();
 sg13g2_fill_2 FILLER_30_1434 ();
 sg13g2_fill_2 FILLER_30_1444 ();
 sg13g2_fill_2 FILLER_30_1467 ();
 sg13g2_decap_8 FILLER_30_1490 ();
 sg13g2_fill_1 FILLER_30_1510 ();
 sg13g2_fill_2 FILLER_30_1515 ();
 sg13g2_fill_1 FILLER_30_1517 ();
 sg13g2_fill_1 FILLER_30_1528 ();
 sg13g2_fill_2 FILLER_30_1561 ();
 sg13g2_fill_1 FILLER_30_1598 ();
 sg13g2_decap_8 FILLER_30_1627 ();
 sg13g2_fill_2 FILLER_30_1634 ();
 sg13g2_decap_8 FILLER_30_1670 ();
 sg13g2_decap_8 FILLER_30_1682 ();
 sg13g2_decap_4 FILLER_30_1689 ();
 sg13g2_decap_4 FILLER_30_1727 ();
 sg13g2_decap_8 FILLER_30_1736 ();
 sg13g2_fill_2 FILLER_30_1743 ();
 sg13g2_fill_2 FILLER_30_1760 ();
 sg13g2_fill_1 FILLER_30_1762 ();
 sg13g2_fill_2 FILLER_30_1775 ();
 sg13g2_fill_1 FILLER_30_1777 ();
 sg13g2_fill_1 FILLER_30_1791 ();
 sg13g2_fill_1 FILLER_30_1805 ();
 sg13g2_fill_2 FILLER_30_1814 ();
 sg13g2_fill_2 FILLER_30_1821 ();
 sg13g2_decap_4 FILLER_30_1830 ();
 sg13g2_fill_2 FILLER_30_1834 ();
 sg13g2_fill_2 FILLER_30_1849 ();
 sg13g2_fill_1 FILLER_30_1851 ();
 sg13g2_fill_1 FILLER_30_1878 ();
 sg13g2_decap_4 FILLER_30_1884 ();
 sg13g2_fill_2 FILLER_30_1888 ();
 sg13g2_fill_2 FILLER_30_1895 ();
 sg13g2_fill_1 FILLER_30_1897 ();
 sg13g2_decap_8 FILLER_30_1921 ();
 sg13g2_fill_1 FILLER_30_1928 ();
 sg13g2_fill_2 FILLER_30_1934 ();
 sg13g2_fill_1 FILLER_30_1936 ();
 sg13g2_fill_1 FILLER_30_1940 ();
 sg13g2_fill_2 FILLER_30_1946 ();
 sg13g2_decap_8 FILLER_30_1952 ();
 sg13g2_decap_8 FILLER_30_1959 ();
 sg13g2_decap_4 FILLER_30_1966 ();
 sg13g2_fill_2 FILLER_30_1978 ();
 sg13g2_fill_2 FILLER_30_1993 ();
 sg13g2_fill_1 FILLER_30_1995 ();
 sg13g2_fill_1 FILLER_30_2014 ();
 sg13g2_fill_2 FILLER_30_2078 ();
 sg13g2_fill_1 FILLER_30_2080 ();
 sg13g2_fill_1 FILLER_30_2094 ();
 sg13g2_fill_1 FILLER_30_2100 ();
 sg13g2_fill_2 FILLER_30_2153 ();
 sg13g2_fill_2 FILLER_30_2163 ();
 sg13g2_fill_1 FILLER_30_2261 ();
 sg13g2_fill_1 FILLER_30_2301 ();
 sg13g2_fill_1 FILLER_30_2327 ();
 sg13g2_fill_2 FILLER_30_2397 ();
 sg13g2_fill_1 FILLER_30_2399 ();
 sg13g2_decap_8 FILLER_30_2408 ();
 sg13g2_fill_2 FILLER_30_2415 ();
 sg13g2_decap_4 FILLER_30_2421 ();
 sg13g2_fill_2 FILLER_30_2425 ();
 sg13g2_fill_2 FILLER_30_2485 ();
 sg13g2_fill_1 FILLER_30_2487 ();
 sg13g2_decap_4 FILLER_30_2514 ();
 sg13g2_decap_8 FILLER_30_2540 ();
 sg13g2_decap_4 FILLER_30_2547 ();
 sg13g2_fill_1 FILLER_30_2568 ();
 sg13g2_fill_2 FILLER_30_2582 ();
 sg13g2_decap_4 FILLER_30_2638 ();
 sg13g2_fill_1 FILLER_30_2642 ();
 sg13g2_fill_2 FILLER_30_2674 ();
 sg13g2_fill_1 FILLER_30_2676 ();
 sg13g2_decap_8 FILLER_30_2719 ();
 sg13g2_fill_2 FILLER_30_2753 ();
 sg13g2_fill_1 FILLER_30_2755 ();
 sg13g2_fill_2 FILLER_30_2791 ();
 sg13g2_fill_1 FILLER_30_2798 ();
 sg13g2_fill_1 FILLER_30_2813 ();
 sg13g2_fill_1 FILLER_30_2853 ();
 sg13g2_fill_2 FILLER_30_2881 ();
 sg13g2_fill_2 FILLER_30_2925 ();
 sg13g2_fill_2 FILLER_30_2936 ();
 sg13g2_fill_1 FILLER_30_2938 ();
 sg13g2_fill_1 FILLER_30_2976 ();
 sg13g2_fill_2 FILLER_30_3012 ();
 sg13g2_fill_1 FILLER_30_3153 ();
 sg13g2_fill_2 FILLER_30_3183 ();
 sg13g2_fill_2 FILLER_30_3196 ();
 sg13g2_fill_1 FILLER_30_3198 ();
 sg13g2_fill_2 FILLER_30_3285 ();
 sg13g2_fill_2 FILLER_30_3299 ();
 sg13g2_fill_1 FILLER_30_3310 ();
 sg13g2_fill_1 FILLER_30_3320 ();
 sg13g2_fill_2 FILLER_30_3343 ();
 sg13g2_fill_2 FILLER_30_3414 ();
 sg13g2_decap_4 FILLER_30_3460 ();
 sg13g2_fill_2 FILLER_30_3487 ();
 sg13g2_decap_4 FILLER_30_3500 ();
 sg13g2_fill_2 FILLER_30_3504 ();
 sg13g2_fill_2 FILLER_30_3518 ();
 sg13g2_fill_2 FILLER_30_3535 ();
 sg13g2_fill_1 FILLER_30_3563 ();
 sg13g2_fill_2 FILLER_30_3577 ();
 sg13g2_fill_1 FILLER_30_3579 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_42 ();
 sg13g2_fill_2 FILLER_31_68 ();
 sg13g2_fill_2 FILLER_31_80 ();
 sg13g2_decap_4 FILLER_31_201 ();
 sg13g2_fill_2 FILLER_31_233 ();
 sg13g2_fill_1 FILLER_31_235 ();
 sg13g2_fill_1 FILLER_31_244 ();
 sg13g2_fill_2 FILLER_31_254 ();
 sg13g2_fill_1 FILLER_31_287 ();
 sg13g2_decap_4 FILLER_31_356 ();
 sg13g2_fill_1 FILLER_31_360 ();
 sg13g2_fill_1 FILLER_31_370 ();
 sg13g2_fill_1 FILLER_31_380 ();
 sg13g2_fill_1 FILLER_31_407 ();
 sg13g2_fill_2 FILLER_31_445 ();
 sg13g2_fill_2 FILLER_31_474 ();
 sg13g2_fill_2 FILLER_31_502 ();
 sg13g2_fill_1 FILLER_31_504 ();
 sg13g2_fill_2 FILLER_31_531 ();
 sg13g2_fill_2 FILLER_31_537 ();
 sg13g2_fill_1 FILLER_31_539 ();
 sg13g2_fill_1 FILLER_31_553 ();
 sg13g2_fill_2 FILLER_31_568 ();
 sg13g2_fill_1 FILLER_31_570 ();
 sg13g2_fill_1 FILLER_31_597 ();
 sg13g2_fill_2 FILLER_31_606 ();
 sg13g2_fill_1 FILLER_31_629 ();
 sg13g2_fill_2 FILLER_31_645 ();
 sg13g2_fill_1 FILLER_31_647 ();
 sg13g2_decap_4 FILLER_31_661 ();
 sg13g2_fill_2 FILLER_31_665 ();
 sg13g2_fill_2 FILLER_31_690 ();
 sg13g2_fill_2 FILLER_31_704 ();
 sg13g2_decap_8 FILLER_31_710 ();
 sg13g2_decap_8 FILLER_31_717 ();
 sg13g2_fill_2 FILLER_31_746 ();
 sg13g2_fill_1 FILLER_31_748 ();
 sg13g2_fill_2 FILLER_31_772 ();
 sg13g2_fill_1 FILLER_31_774 ();
 sg13g2_fill_2 FILLER_31_803 ();
 sg13g2_fill_2 FILLER_31_870 ();
 sg13g2_fill_1 FILLER_31_872 ();
 sg13g2_fill_1 FILLER_31_882 ();
 sg13g2_fill_2 FILLER_31_944 ();
 sg13g2_fill_1 FILLER_31_946 ();
 sg13g2_fill_2 FILLER_31_984 ();
 sg13g2_fill_1 FILLER_31_1010 ();
 sg13g2_fill_2 FILLER_31_1080 ();
 sg13g2_fill_2 FILLER_31_1126 ();
 sg13g2_fill_1 FILLER_31_1177 ();
 sg13g2_fill_2 FILLER_31_1199 ();
 sg13g2_fill_2 FILLER_31_1253 ();
 sg13g2_fill_1 FILLER_31_1266 ();
 sg13g2_fill_2 FILLER_31_1307 ();
 sg13g2_decap_4 FILLER_31_1318 ();
 sg13g2_fill_2 FILLER_31_1361 ();
 sg13g2_fill_2 FILLER_31_1368 ();
 sg13g2_decap_8 FILLER_31_1395 ();
 sg13g2_decap_4 FILLER_31_1402 ();
 sg13g2_fill_2 FILLER_31_1406 ();
 sg13g2_fill_1 FILLER_31_1413 ();
 sg13g2_fill_2 FILLER_31_1423 ();
 sg13g2_fill_1 FILLER_31_1425 ();
 sg13g2_decap_4 FILLER_31_1443 ();
 sg13g2_fill_1 FILLER_31_1447 ();
 sg13g2_fill_1 FILLER_31_1461 ();
 sg13g2_fill_2 FILLER_31_1475 ();
 sg13g2_decap_4 FILLER_31_1497 ();
 sg13g2_fill_2 FILLER_31_1511 ();
 sg13g2_decap_8 FILLER_31_1532 ();
 sg13g2_decap_8 FILLER_31_1552 ();
 sg13g2_decap_4 FILLER_31_1559 ();
 sg13g2_fill_1 FILLER_31_1563 ();
 sg13g2_fill_2 FILLER_31_1584 ();
 sg13g2_fill_1 FILLER_31_1586 ();
 sg13g2_fill_2 FILLER_31_1600 ();
 sg13g2_fill_1 FILLER_31_1602 ();
 sg13g2_fill_2 FILLER_31_1607 ();
 sg13g2_fill_1 FILLER_31_1609 ();
 sg13g2_decap_4 FILLER_31_1623 ();
 sg13g2_decap_8 FILLER_31_1663 ();
 sg13g2_decap_4 FILLER_31_1670 ();
 sg13g2_fill_1 FILLER_31_1674 ();
 sg13g2_decap_4 FILLER_31_1688 ();
 sg13g2_fill_1 FILLER_31_1692 ();
 sg13g2_fill_1 FILLER_31_1710 ();
 sg13g2_decap_8 FILLER_31_1728 ();
 sg13g2_decap_8 FILLER_31_1735 ();
 sg13g2_fill_2 FILLER_31_1742 ();
 sg13g2_fill_1 FILLER_31_1744 ();
 sg13g2_fill_2 FILLER_31_1758 ();
 sg13g2_decap_8 FILLER_31_1773 ();
 sg13g2_decap_8 FILLER_31_1785 ();
 sg13g2_decap_8 FILLER_31_1792 ();
 sg13g2_decap_8 FILLER_31_1799 ();
 sg13g2_fill_2 FILLER_31_1806 ();
 sg13g2_decap_8 FILLER_31_1812 ();
 sg13g2_fill_2 FILLER_31_1819 ();
 sg13g2_fill_1 FILLER_31_1837 ();
 sg13g2_decap_4 FILLER_31_1848 ();
 sg13g2_decap_8 FILLER_31_1870 ();
 sg13g2_decap_4 FILLER_31_1877 ();
 sg13g2_fill_2 FILLER_31_1888 ();
 sg13g2_fill_2 FILLER_31_1941 ();
 sg13g2_decap_4 FILLER_31_1971 ();
 sg13g2_fill_1 FILLER_31_1975 ();
 sg13g2_decap_8 FILLER_31_2013 ();
 sg13g2_fill_1 FILLER_31_2020 ();
 sg13g2_fill_1 FILLER_31_2110 ();
 sg13g2_decap_8 FILLER_31_2123 ();
 sg13g2_fill_2 FILLER_31_2171 ();
 sg13g2_fill_1 FILLER_31_2173 ();
 sg13g2_fill_2 FILLER_31_2197 ();
 sg13g2_fill_2 FILLER_31_2228 ();
 sg13g2_fill_1 FILLER_31_2230 ();
 sg13g2_decap_8 FILLER_31_2259 ();
 sg13g2_decap_8 FILLER_31_2266 ();
 sg13g2_fill_1 FILLER_31_2346 ();
 sg13g2_fill_2 FILLER_31_2352 ();
 sg13g2_fill_1 FILLER_31_2367 ();
 sg13g2_fill_2 FILLER_31_2381 ();
 sg13g2_fill_1 FILLER_31_2383 ();
 sg13g2_decap_4 FILLER_31_2390 ();
 sg13g2_fill_2 FILLER_31_2394 ();
 sg13g2_decap_4 FILLER_31_2401 ();
 sg13g2_fill_2 FILLER_31_2440 ();
 sg13g2_fill_1 FILLER_31_2442 ();
 sg13g2_fill_2 FILLER_31_2456 ();
 sg13g2_fill_1 FILLER_31_2458 ();
 sg13g2_fill_2 FILLER_31_2475 ();
 sg13g2_decap_4 FILLER_31_2514 ();
 sg13g2_fill_2 FILLER_31_2549 ();
 sg13g2_fill_1 FILLER_31_2551 ();
 sg13g2_fill_2 FILLER_31_2574 ();
 sg13g2_fill_1 FILLER_31_2589 ();
 sg13g2_fill_2 FILLER_31_2604 ();
 sg13g2_fill_1 FILLER_31_2606 ();
 sg13g2_decap_4 FILLER_31_2658 ();
 sg13g2_fill_2 FILLER_31_2699 ();
 sg13g2_decap_8 FILLER_31_2728 ();
 sg13g2_decap_4 FILLER_31_2748 ();
 sg13g2_fill_2 FILLER_31_2752 ();
 sg13g2_fill_1 FILLER_31_2782 ();
 sg13g2_fill_1 FILLER_31_2833 ();
 sg13g2_fill_1 FILLER_31_2903 ();
 sg13g2_fill_1 FILLER_31_2931 ();
 sg13g2_fill_1 FILLER_31_2977 ();
 sg13g2_fill_2 FILLER_31_3050 ();
 sg13g2_fill_2 FILLER_31_3086 ();
 sg13g2_fill_2 FILLER_31_3124 ();
 sg13g2_fill_1 FILLER_31_3126 ();
 sg13g2_fill_1 FILLER_31_3252 ();
 sg13g2_fill_1 FILLER_31_3265 ();
 sg13g2_fill_2 FILLER_31_3322 ();
 sg13g2_fill_2 FILLER_31_3332 ();
 sg13g2_fill_1 FILLER_31_3334 ();
 sg13g2_fill_2 FILLER_31_3367 ();
 sg13g2_fill_1 FILLER_31_3382 ();
 sg13g2_decap_8 FILLER_31_3415 ();
 sg13g2_fill_2 FILLER_31_3422 ();
 sg13g2_fill_1 FILLER_31_3428 ();
 sg13g2_fill_1 FILLER_31_3437 ();
 sg13g2_fill_2 FILLER_31_3516 ();
 sg13g2_fill_1 FILLER_31_3546 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_4 ();
 sg13g2_decap_4 FILLER_32_10 ();
 sg13g2_fill_2 FILLER_32_14 ();
 sg13g2_fill_1 FILLER_32_33 ();
 sg13g2_decap_4 FILLER_32_50 ();
 sg13g2_decap_4 FILLER_32_59 ();
 sg13g2_fill_1 FILLER_32_78 ();
 sg13g2_fill_2 FILLER_32_147 ();
 sg13g2_fill_2 FILLER_32_176 ();
 sg13g2_fill_1 FILLER_32_178 ();
 sg13g2_decap_4 FILLER_32_209 ();
 sg13g2_fill_2 FILLER_32_213 ();
 sg13g2_fill_2 FILLER_32_228 ();
 sg13g2_fill_1 FILLER_32_230 ();
 sg13g2_decap_8 FILLER_32_240 ();
 sg13g2_decap_4 FILLER_32_247 ();
 sg13g2_fill_1 FILLER_32_251 ();
 sg13g2_decap_8 FILLER_32_279 ();
 sg13g2_fill_1 FILLER_32_286 ();
 sg13g2_fill_2 FILLER_32_315 ();
 sg13g2_fill_1 FILLER_32_317 ();
 sg13g2_fill_1 FILLER_32_326 ();
 sg13g2_fill_2 FILLER_32_404 ();
 sg13g2_fill_2 FILLER_32_453 ();
 sg13g2_fill_2 FILLER_32_521 ();
 sg13g2_fill_1 FILLER_32_556 ();
 sg13g2_fill_1 FILLER_32_562 ();
 sg13g2_fill_2 FILLER_32_576 ();
 sg13g2_fill_2 FILLER_32_595 ();
 sg13g2_decap_4 FILLER_32_621 ();
 sg13g2_fill_2 FILLER_32_645 ();
 sg13g2_decap_4 FILLER_32_659 ();
 sg13g2_fill_1 FILLER_32_674 ();
 sg13g2_fill_2 FILLER_32_688 ();
 sg13g2_fill_1 FILLER_32_690 ();
 sg13g2_fill_1 FILLER_32_707 ();
 sg13g2_fill_2 FILLER_32_729 ();
 sg13g2_fill_1 FILLER_32_731 ();
 sg13g2_fill_2 FILLER_32_776 ();
 sg13g2_fill_1 FILLER_32_778 ();
 sg13g2_fill_1 FILLER_32_787 ();
 sg13g2_decap_8 FILLER_32_797 ();
 sg13g2_fill_1 FILLER_32_804 ();
 sg13g2_fill_2 FILLER_32_871 ();
 sg13g2_fill_2 FILLER_32_946 ();
 sg13g2_fill_1 FILLER_32_948 ();
 sg13g2_fill_1 FILLER_32_975 ();
 sg13g2_fill_1 FILLER_32_1060 ();
 sg13g2_decap_8 FILLER_32_1065 ();
 sg13g2_fill_2 FILLER_32_1072 ();
 sg13g2_decap_4 FILLER_32_1090 ();
 sg13g2_fill_2 FILLER_32_1144 ();
 sg13g2_fill_1 FILLER_32_1146 ();
 sg13g2_fill_1 FILLER_32_1160 ();
 sg13g2_fill_2 FILLER_32_1206 ();
 sg13g2_fill_2 FILLER_32_1212 ();
 sg13g2_fill_2 FILLER_32_1234 ();
 sg13g2_fill_1 FILLER_32_1236 ();
 sg13g2_fill_2 FILLER_32_1276 ();
 sg13g2_fill_1 FILLER_32_1278 ();
 sg13g2_fill_2 FILLER_32_1288 ();
 sg13g2_fill_2 FILLER_32_1294 ();
 sg13g2_fill_1 FILLER_32_1296 ();
 sg13g2_fill_2 FILLER_32_1322 ();
 sg13g2_decap_8 FILLER_32_1338 ();
 sg13g2_fill_2 FILLER_32_1361 ();
 sg13g2_fill_1 FILLER_32_1363 ();
 sg13g2_fill_1 FILLER_32_1391 ();
 sg13g2_fill_1 FILLER_32_1405 ();
 sg13g2_fill_2 FILLER_32_1539 ();
 sg13g2_decap_8 FILLER_32_1582 ();
 sg13g2_fill_1 FILLER_32_1630 ();
 sg13g2_fill_2 FILLER_32_1659 ();
 sg13g2_fill_2 FILLER_32_1689 ();
 sg13g2_fill_1 FILLER_32_1691 ();
 sg13g2_decap_8 FILLER_32_1696 ();
 sg13g2_decap_4 FILLER_32_1703 ();
 sg13g2_decap_4 FILLER_32_1720 ();
 sg13g2_fill_2 FILLER_32_1724 ();
 sg13g2_decap_8 FILLER_32_1736 ();
 sg13g2_fill_2 FILLER_32_1743 ();
 sg13g2_decap_8 FILLER_32_1820 ();
 sg13g2_decap_4 FILLER_32_1827 ();
 sg13g2_fill_1 FILLER_32_1831 ();
 sg13g2_decap_8 FILLER_32_1840 ();
 sg13g2_fill_2 FILLER_32_1856 ();
 sg13g2_decap_4 FILLER_32_1893 ();
 sg13g2_fill_2 FILLER_32_1897 ();
 sg13g2_decap_8 FILLER_32_1924 ();
 sg13g2_fill_2 FILLER_32_1931 ();
 sg13g2_decap_8 FILLER_32_1938 ();
 sg13g2_decap_8 FILLER_32_1945 ();
 sg13g2_fill_1 FILLER_32_1952 ();
 sg13g2_decap_4 FILLER_32_1981 ();
 sg13g2_fill_2 FILLER_32_1985 ();
 sg13g2_decap_4 FILLER_32_2009 ();
 sg13g2_decap_8 FILLER_32_2053 ();
 sg13g2_decap_8 FILLER_32_2126 ();
 sg13g2_fill_2 FILLER_32_2133 ();
 sg13g2_fill_2 FILLER_32_2140 ();
 sg13g2_fill_2 FILLER_32_2146 ();
 sg13g2_fill_1 FILLER_32_2148 ();
 sg13g2_decap_4 FILLER_32_2171 ();
 sg13g2_fill_1 FILLER_32_2198 ();
 sg13g2_fill_1 FILLER_32_2221 ();
 sg13g2_fill_2 FILLER_32_2234 ();
 sg13g2_decap_8 FILLER_32_2258 ();
 sg13g2_fill_1 FILLER_32_2265 ();
 sg13g2_fill_2 FILLER_32_2270 ();
 sg13g2_fill_2 FILLER_32_2326 ();
 sg13g2_decap_4 FILLER_32_2347 ();
 sg13g2_fill_2 FILLER_32_2356 ();
 sg13g2_fill_1 FILLER_32_2358 ();
 sg13g2_decap_4 FILLER_32_2368 ();
 sg13g2_fill_1 FILLER_32_2376 ();
 sg13g2_fill_1 FILLER_32_2389 ();
 sg13g2_fill_2 FILLER_32_2404 ();
 sg13g2_fill_1 FILLER_32_2414 ();
 sg13g2_fill_2 FILLER_32_2452 ();
 sg13g2_decap_4 FILLER_32_2498 ();
 sg13g2_fill_1 FILLER_32_2502 ();
 sg13g2_fill_1 FILLER_32_2513 ();
 sg13g2_fill_2 FILLER_32_2524 ();
 sg13g2_fill_2 FILLER_32_2554 ();
 sg13g2_fill_1 FILLER_32_2556 ();
 sg13g2_fill_1 FILLER_32_2613 ();
 sg13g2_fill_1 FILLER_32_2618 ();
 sg13g2_decap_4 FILLER_32_2647 ();
 sg13g2_fill_1 FILLER_32_2683 ();
 sg13g2_decap_4 FILLER_32_2711 ();
 sg13g2_fill_1 FILLER_32_2715 ();
 sg13g2_fill_1 FILLER_32_2766 ();
 sg13g2_fill_1 FILLER_32_2831 ();
 sg13g2_fill_1 FILLER_32_2853 ();
 sg13g2_fill_2 FILLER_32_2867 ();
 sg13g2_fill_2 FILLER_32_2884 ();
 sg13g2_fill_1 FILLER_32_2886 ();
 sg13g2_fill_1 FILLER_32_2913 ();
 sg13g2_fill_1 FILLER_32_2941 ();
 sg13g2_fill_2 FILLER_32_2982 ();
 sg13g2_fill_1 FILLER_32_2984 ();
 sg13g2_fill_1 FILLER_32_3008 ();
 sg13g2_fill_1 FILLER_32_3084 ();
 sg13g2_fill_1 FILLER_32_3124 ();
 sg13g2_fill_2 FILLER_32_3131 ();
 sg13g2_fill_2 FILLER_32_3155 ();
 sg13g2_fill_1 FILLER_32_3212 ();
 sg13g2_fill_1 FILLER_32_3222 ();
 sg13g2_fill_1 FILLER_32_3273 ();
 sg13g2_fill_2 FILLER_32_3291 ();
 sg13g2_fill_2 FILLER_32_3313 ();
 sg13g2_fill_1 FILLER_32_3319 ();
 sg13g2_fill_2 FILLER_32_3378 ();
 sg13g2_fill_2 FILLER_32_3408 ();
 sg13g2_fill_1 FILLER_32_3410 ();
 sg13g2_fill_1 FILLER_32_3473 ();
 sg13g2_fill_1 FILLER_32_3484 ();
 sg13g2_fill_2 FILLER_32_3490 ();
 sg13g2_decap_8 FILLER_32_3507 ();
 sg13g2_decap_8 FILLER_32_3514 ();
 sg13g2_fill_1 FILLER_32_3521 ();
 sg13g2_decap_4 FILLER_32_3535 ();
 sg13g2_fill_1 FILLER_32_3539 ();
 sg13g2_fill_1 FILLER_32_3562 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_43 ();
 sg13g2_decap_8 FILLER_33_58 ();
 sg13g2_fill_2 FILLER_33_93 ();
 sg13g2_fill_1 FILLER_33_95 ();
 sg13g2_decap_4 FILLER_33_102 ();
 sg13g2_decap_8 FILLER_33_117 ();
 sg13g2_fill_2 FILLER_33_124 ();
 sg13g2_fill_2 FILLER_33_171 ();
 sg13g2_fill_1 FILLER_33_173 ();
 sg13g2_fill_2 FILLER_33_230 ();
 sg13g2_fill_1 FILLER_33_232 ();
 sg13g2_fill_1 FILLER_33_238 ();
 sg13g2_fill_2 FILLER_33_266 ();
 sg13g2_fill_1 FILLER_33_268 ();
 sg13g2_fill_1 FILLER_33_295 ();
 sg13g2_fill_1 FILLER_33_314 ();
 sg13g2_fill_2 FILLER_33_329 ();
 sg13g2_fill_1 FILLER_33_331 ();
 sg13g2_decap_4 FILLER_33_359 ();
 sg13g2_fill_2 FILLER_33_363 ();
 sg13g2_fill_2 FILLER_33_382 ();
 sg13g2_fill_1 FILLER_33_384 ();
 sg13g2_fill_1 FILLER_33_390 ();
 sg13g2_fill_1 FILLER_33_399 ();
 sg13g2_fill_2 FILLER_33_405 ();
 sg13g2_fill_1 FILLER_33_407 ();
 sg13g2_fill_2 FILLER_33_420 ();
 sg13g2_fill_1 FILLER_33_422 ();
 sg13g2_decap_8 FILLER_33_428 ();
 sg13g2_decap_4 FILLER_33_435 ();
 sg13g2_fill_2 FILLER_33_504 ();
 sg13g2_fill_1 FILLER_33_506 ();
 sg13g2_fill_2 FILLER_33_524 ();
 sg13g2_decap_8 FILLER_33_554 ();
 sg13g2_fill_1 FILLER_33_561 ();
 sg13g2_fill_2 FILLER_33_583 ();
 sg13g2_fill_2 FILLER_33_590 ();
 sg13g2_fill_2 FILLER_33_597 ();
 sg13g2_fill_1 FILLER_33_599 ();
 sg13g2_fill_2 FILLER_33_605 ();
 sg13g2_fill_1 FILLER_33_607 ();
 sg13g2_fill_2 FILLER_33_645 ();
 sg13g2_decap_8 FILLER_33_657 ();
 sg13g2_decap_8 FILLER_33_664 ();
 sg13g2_fill_1 FILLER_33_671 ();
 sg13g2_fill_2 FILLER_33_676 ();
 sg13g2_fill_1 FILLER_33_678 ();
 sg13g2_fill_1 FILLER_33_699 ();
 sg13g2_decap_8 FILLER_33_705 ();
 sg13g2_fill_2 FILLER_33_712 ();
 sg13g2_fill_2 FILLER_33_728 ();
 sg13g2_fill_1 FILLER_33_730 ();
 sg13g2_fill_1 FILLER_33_739 ();
 sg13g2_fill_1 FILLER_33_787 ();
 sg13g2_fill_1 FILLER_33_792 ();
 sg13g2_decap_8 FILLER_33_862 ();
 sg13g2_decap_4 FILLER_33_869 ();
 sg13g2_fill_2 FILLER_33_873 ();
 sg13g2_fill_2 FILLER_33_914 ();
 sg13g2_fill_1 FILLER_33_916 ();
 sg13g2_fill_2 FILLER_33_930 ();
 sg13g2_fill_1 FILLER_33_932 ();
 sg13g2_fill_2 FILLER_33_998 ();
 sg13g2_fill_2 FILLER_33_1033 ();
 sg13g2_fill_1 FILLER_33_1035 ();
 sg13g2_fill_1 FILLER_33_1097 ();
 sg13g2_decap_4 FILLER_33_1156 ();
 sg13g2_fill_2 FILLER_33_1160 ();
 sg13g2_decap_4 FILLER_33_1261 ();
 sg13g2_fill_1 FILLER_33_1270 ();
 sg13g2_fill_2 FILLER_33_1294 ();
 sg13g2_fill_1 FILLER_33_1296 ();
 sg13g2_fill_2 FILLER_33_1320 ();
 sg13g2_fill_1 FILLER_33_1322 ();
 sg13g2_decap_4 FILLER_33_1339 ();
 sg13g2_fill_1 FILLER_33_1364 ();
 sg13g2_decap_8 FILLER_33_1401 ();
 sg13g2_fill_2 FILLER_33_1413 ();
 sg13g2_fill_1 FILLER_33_1420 ();
 sg13g2_decap_4 FILLER_33_1431 ();
 sg13g2_fill_1 FILLER_33_1435 ();
 sg13g2_fill_2 FILLER_33_1453 ();
 sg13g2_fill_2 FILLER_33_1474 ();
 sg13g2_decap_8 FILLER_33_1502 ();
 sg13g2_decap_4 FILLER_33_1509 ();
 sg13g2_fill_2 FILLER_33_1513 ();
 sg13g2_decap_8 FILLER_33_1551 ();
 sg13g2_fill_1 FILLER_33_1558 ();
 sg13g2_decap_4 FILLER_33_1563 ();
 sg13g2_fill_1 FILLER_33_1567 ();
 sg13g2_decap_4 FILLER_33_1581 ();
 sg13g2_decap_8 FILLER_33_1588 ();
 sg13g2_decap_4 FILLER_33_1598 ();
 sg13g2_fill_1 FILLER_33_1602 ();
 sg13g2_decap_8 FILLER_33_1620 ();
 sg13g2_decap_4 FILLER_33_1627 ();
 sg13g2_decap_4 FILLER_33_1646 ();
 sg13g2_fill_2 FILLER_33_1719 ();
 sg13g2_fill_2 FILLER_33_1770 ();
 sg13g2_fill_2 FILLER_33_1782 ();
 sg13g2_decap_8 FILLER_33_1788 ();
 sg13g2_fill_2 FILLER_33_1795 ();
 sg13g2_fill_1 FILLER_33_1797 ();
 sg13g2_decap_4 FILLER_33_1861 ();
 sg13g2_fill_1 FILLER_33_1865 ();
 sg13g2_decap_8 FILLER_33_1879 ();
 sg13g2_decap_8 FILLER_33_1886 ();
 sg13g2_fill_1 FILLER_33_1893 ();
 sg13g2_fill_2 FILLER_33_1905 ();
 sg13g2_fill_2 FILLER_33_1925 ();
 sg13g2_fill_1 FILLER_33_1927 ();
 sg13g2_fill_1 FILLER_33_1962 ();
 sg13g2_decap_8 FILLER_33_1972 ();
 sg13g2_fill_2 FILLER_33_1979 ();
 sg13g2_fill_2 FILLER_33_2072 ();
 sg13g2_fill_1 FILLER_33_2074 ();
 sg13g2_fill_2 FILLER_33_2114 ();
 sg13g2_fill_2 FILLER_33_2126 ();
 sg13g2_fill_2 FILLER_33_2153 ();
 sg13g2_decap_4 FILLER_33_2175 ();
 sg13g2_fill_2 FILLER_33_2188 ();
 sg13g2_fill_1 FILLER_33_2190 ();
 sg13g2_fill_1 FILLER_33_2205 ();
 sg13g2_fill_2 FILLER_33_2215 ();
 sg13g2_fill_1 FILLER_33_2217 ();
 sg13g2_fill_2 FILLER_33_2244 ();
 sg13g2_fill_1 FILLER_33_2246 ();
 sg13g2_decap_4 FILLER_33_2255 ();
 sg13g2_fill_2 FILLER_33_2259 ();
 sg13g2_fill_2 FILLER_33_2299 ();
 sg13g2_fill_1 FILLER_33_2301 ();
 sg13g2_fill_1 FILLER_33_2327 ();
 sg13g2_decap_4 FILLER_33_2396 ();
 sg13g2_fill_2 FILLER_33_2421 ();
 sg13g2_fill_1 FILLER_33_2423 ();
 sg13g2_fill_2 FILLER_33_2442 ();
 sg13g2_fill_1 FILLER_33_2456 ();
 sg13g2_fill_2 FILLER_33_2470 ();
 sg13g2_fill_2 FILLER_33_2485 ();
 sg13g2_fill_1 FILLER_33_2487 ();
 sg13g2_decap_8 FILLER_33_2501 ();
 sg13g2_fill_1 FILLER_33_2508 ();
 sg13g2_fill_2 FILLER_33_2576 ();
 sg13g2_fill_2 FILLER_33_2591 ();
 sg13g2_fill_1 FILLER_33_2593 ();
 sg13g2_fill_2 FILLER_33_2615 ();
 sg13g2_fill_1 FILLER_33_2617 ();
 sg13g2_fill_1 FILLER_33_2631 ();
 sg13g2_fill_1 FILLER_33_2641 ();
 sg13g2_fill_1 FILLER_33_2682 ();
 sg13g2_decap_8 FILLER_33_2711 ();
 sg13g2_fill_2 FILLER_33_2728 ();
 sg13g2_fill_1 FILLER_33_2730 ();
 sg13g2_fill_2 FILLER_33_2803 ();
 sg13g2_fill_2 FILLER_33_2916 ();
 sg13g2_fill_1 FILLER_33_2918 ();
 sg13g2_fill_2 FILLER_33_2932 ();
 sg13g2_decap_4 FILLER_33_2953 ();
 sg13g2_fill_2 FILLER_33_3011 ();
 sg13g2_fill_1 FILLER_33_3077 ();
 sg13g2_fill_1 FILLER_33_3091 ();
 sg13g2_fill_1 FILLER_33_3122 ();
 sg13g2_fill_2 FILLER_33_3131 ();
 sg13g2_fill_1 FILLER_33_3278 ();
 sg13g2_decap_8 FILLER_33_3288 ();
 sg13g2_fill_1 FILLER_33_3295 ();
 sg13g2_fill_2 FILLER_33_3300 ();
 sg13g2_fill_1 FILLER_33_3310 ();
 sg13g2_fill_2 FILLER_33_3349 ();
 sg13g2_fill_1 FILLER_33_3351 ();
 sg13g2_decap_8 FILLER_33_3439 ();
 sg13g2_fill_2 FILLER_33_3466 ();
 sg13g2_fill_1 FILLER_33_3493 ();
 sg13g2_decap_8 FILLER_33_3512 ();
 sg13g2_fill_1 FILLER_33_3519 ();
 sg13g2_fill_2 FILLER_33_3540 ();
 sg13g2_fill_1 FILLER_33_3542 ();
 sg13g2_fill_1 FILLER_33_3551 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_4 ();
 sg13g2_decap_8 FILLER_34_117 ();
 sg13g2_decap_8 FILLER_34_124 ();
 sg13g2_fill_1 FILLER_34_131 ();
 sg13g2_fill_2 FILLER_34_223 ();
 sg13g2_decap_8 FILLER_34_260 ();
 sg13g2_fill_1 FILLER_34_272 ();
 sg13g2_fill_2 FILLER_34_286 ();
 sg13g2_fill_2 FILLER_34_320 ();
 sg13g2_fill_1 FILLER_34_322 ();
 sg13g2_fill_2 FILLER_34_333 ();
 sg13g2_fill_2 FILLER_34_340 ();
 sg13g2_fill_1 FILLER_34_342 ();
 sg13g2_decap_4 FILLER_34_364 ();
 sg13g2_fill_1 FILLER_34_368 ();
 sg13g2_fill_1 FILLER_34_376 ();
 sg13g2_decap_8 FILLER_34_390 ();
 sg13g2_decap_8 FILLER_34_397 ();
 sg13g2_fill_1 FILLER_34_404 ();
 sg13g2_decap_4 FILLER_34_413 ();
 sg13g2_decap_4 FILLER_34_474 ();
 sg13g2_fill_2 FILLER_34_478 ();
 sg13g2_fill_2 FILLER_34_513 ();
 sg13g2_fill_1 FILLER_34_515 ();
 sg13g2_fill_2 FILLER_34_525 ();
 sg13g2_fill_1 FILLER_34_527 ();
 sg13g2_fill_1 FILLER_34_533 ();
 sg13g2_fill_1 FILLER_34_543 ();
 sg13g2_decap_4 FILLER_34_562 ();
 sg13g2_fill_2 FILLER_34_566 ();
 sg13g2_fill_1 FILLER_34_576 ();
 sg13g2_fill_1 FILLER_34_602 ();
 sg13g2_decap_4 FILLER_34_611 ();
 sg13g2_fill_2 FILLER_34_615 ();
 sg13g2_fill_1 FILLER_34_625 ();
 sg13g2_fill_2 FILLER_34_643 ();
 sg13g2_fill_1 FILLER_34_645 ();
 sg13g2_decap_4 FILLER_34_663 ();
 sg13g2_fill_2 FILLER_34_667 ();
 sg13g2_fill_1 FILLER_34_681 ();
 sg13g2_decap_4 FILLER_34_699 ();
 sg13g2_fill_2 FILLER_34_703 ();
 sg13g2_decap_8 FILLER_34_710 ();
 sg13g2_decap_8 FILLER_34_717 ();
 sg13g2_decap_4 FILLER_34_724 ();
 sg13g2_fill_1 FILLER_34_728 ();
 sg13g2_fill_1 FILLER_34_747 ();
 sg13g2_fill_2 FILLER_34_791 ();
 sg13g2_decap_8 FILLER_34_806 ();
 sg13g2_fill_2 FILLER_34_813 ();
 sg13g2_fill_1 FILLER_34_815 ();
 sg13g2_fill_1 FILLER_34_910 ();
 sg13g2_fill_1 FILLER_34_952 ();
 sg13g2_fill_2 FILLER_34_975 ();
 sg13g2_fill_1 FILLER_34_977 ();
 sg13g2_fill_2 FILLER_34_987 ();
 sg13g2_fill_1 FILLER_34_989 ();
 sg13g2_fill_2 FILLER_34_1003 ();
 sg13g2_fill_1 FILLER_34_1014 ();
 sg13g2_fill_2 FILLER_34_1037 ();
 sg13g2_fill_1 FILLER_34_1053 ();
 sg13g2_decap_4 FILLER_34_1072 ();
 sg13g2_fill_1 FILLER_34_1076 ();
 sg13g2_fill_2 FILLER_34_1128 ();
 sg13g2_fill_1 FILLER_34_1220 ();
 sg13g2_fill_1 FILLER_34_1234 ();
 sg13g2_decap_4 FILLER_34_1248 ();
 sg13g2_fill_2 FILLER_34_1252 ();
 sg13g2_decap_4 FILLER_34_1263 ();
 sg13g2_fill_2 FILLER_34_1267 ();
 sg13g2_fill_2 FILLER_34_1285 ();
 sg13g2_decap_4 FILLER_34_1312 ();
 sg13g2_decap_8 FILLER_34_1329 ();
 sg13g2_decap_8 FILLER_34_1336 ();
 sg13g2_fill_1 FILLER_34_1369 ();
 sg13g2_fill_2 FILLER_34_1397 ();
 sg13g2_decap_4 FILLER_34_1404 ();
 sg13g2_fill_2 FILLER_34_1421 ();
 sg13g2_fill_2 FILLER_34_1432 ();
 sg13g2_fill_1 FILLER_34_1434 ();
 sg13g2_fill_1 FILLER_34_1489 ();
 sg13g2_fill_2 FILLER_34_1502 ();
 sg13g2_fill_1 FILLER_34_1504 ();
 sg13g2_fill_1 FILLER_34_1510 ();
 sg13g2_decap_8 FILLER_34_1556 ();
 sg13g2_fill_2 FILLER_34_1563 ();
 sg13g2_fill_1 FILLER_34_1591 ();
 sg13g2_decap_4 FILLER_34_1625 ();
 sg13g2_decap_4 FILLER_34_1633 ();
 sg13g2_fill_1 FILLER_34_1673 ();
 sg13g2_decap_8 FILLER_34_1688 ();
 sg13g2_decap_4 FILLER_34_1695 ();
 sg13g2_fill_2 FILLER_34_1699 ();
 sg13g2_decap_4 FILLER_34_1726 ();
 sg13g2_fill_2 FILLER_34_1760 ();
 sg13g2_decap_4 FILLER_34_1815 ();
 sg13g2_fill_2 FILLER_34_1819 ();
 sg13g2_decap_4 FILLER_34_1860 ();
 sg13g2_fill_1 FILLER_34_1884 ();
 sg13g2_decap_4 FILLER_34_1923 ();
 sg13g2_decap_8 FILLER_34_1947 ();
 sg13g2_fill_2 FILLER_34_1954 ();
 sg13g2_decap_4 FILLER_34_1975 ();
 sg13g2_fill_2 FILLER_34_2000 ();
 sg13g2_decap_4 FILLER_34_2011 ();
 sg13g2_fill_1 FILLER_34_2015 ();
 sg13g2_decap_4 FILLER_34_2076 ();
 sg13g2_fill_2 FILLER_34_2114 ();
 sg13g2_fill_1 FILLER_34_2116 ();
 sg13g2_fill_2 FILLER_34_2135 ();
 sg13g2_fill_1 FILLER_34_2147 ();
 sg13g2_decap_8 FILLER_34_2168 ();
 sg13g2_fill_2 FILLER_34_2175 ();
 sg13g2_fill_1 FILLER_34_2177 ();
 sg13g2_decap_4 FILLER_34_2204 ();
 sg13g2_fill_1 FILLER_34_2213 ();
 sg13g2_decap_4 FILLER_34_2229 ();
 sg13g2_fill_1 FILLER_34_2263 ();
 sg13g2_decap_4 FILLER_34_2267 ();
 sg13g2_fill_2 FILLER_34_2275 ();
 sg13g2_decap_4 FILLER_34_2293 ();
 sg13g2_decap_4 FILLER_34_2322 ();
 sg13g2_fill_2 FILLER_34_2359 ();
 sg13g2_decap_4 FILLER_34_2395 ();
 sg13g2_fill_2 FILLER_34_2399 ();
 sg13g2_fill_1 FILLER_34_2414 ();
 sg13g2_fill_1 FILLER_34_2428 ();
 sg13g2_fill_1 FILLER_34_2449 ();
 sg13g2_fill_2 FILLER_34_2454 ();
 sg13g2_fill_2 FILLER_34_2472 ();
 sg13g2_fill_1 FILLER_34_2474 ();
 sg13g2_fill_1 FILLER_34_2508 ();
 sg13g2_fill_2 FILLER_34_2518 ();
 sg13g2_fill_2 FILLER_34_2533 ();
 sg13g2_fill_1 FILLER_34_2535 ();
 sg13g2_fill_2 FILLER_34_2579 ();
 sg13g2_fill_1 FILLER_34_2581 ();
 sg13g2_fill_1 FILLER_34_2586 ();
 sg13g2_fill_2 FILLER_34_2611 ();
 sg13g2_decap_4 FILLER_34_2650 ();
 sg13g2_fill_2 FILLER_34_2654 ();
 sg13g2_fill_2 FILLER_34_2665 ();
 sg13g2_fill_1 FILLER_34_2667 ();
 sg13g2_fill_2 FILLER_34_2719 ();
 sg13g2_fill_2 FILLER_34_2758 ();
 sg13g2_fill_1 FILLER_34_2760 ();
 sg13g2_fill_2 FILLER_34_2825 ();
 sg13g2_fill_1 FILLER_34_2827 ();
 sg13g2_fill_1 FILLER_34_2899 ();
 sg13g2_fill_1 FILLER_34_2909 ();
 sg13g2_fill_2 FILLER_34_2970 ();
 sg13g2_fill_1 FILLER_34_2972 ();
 sg13g2_fill_1 FILLER_34_3006 ();
 sg13g2_fill_2 FILLER_34_3149 ();
 sg13g2_fill_1 FILLER_34_3184 ();
 sg13g2_fill_1 FILLER_34_3202 ();
 sg13g2_fill_1 FILLER_34_3216 ();
 sg13g2_fill_2 FILLER_34_3272 ();
 sg13g2_fill_1 FILLER_34_3274 ();
 sg13g2_decap_4 FILLER_34_3437 ();
 sg13g2_fill_2 FILLER_34_3441 ();
 sg13g2_fill_2 FILLER_34_3460 ();
 sg13g2_fill_1 FILLER_34_3462 ();
 sg13g2_fill_2 FILLER_34_3486 ();
 sg13g2_fill_1 FILLER_34_3488 ();
 sg13g2_decap_4 FILLER_34_3516 ();
 sg13g2_decap_8 FILLER_34_3535 ();
 sg13g2_fill_2 FILLER_34_3542 ();
 sg13g2_fill_2 FILLER_34_3552 ();
 sg13g2_fill_1 FILLER_34_3554 ();
 sg13g2_decap_4 FILLER_34_3576 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_4 ();
 sg13g2_decap_4 FILLER_35_10 ();
 sg13g2_fill_1 FILLER_35_14 ();
 sg13g2_fill_1 FILLER_35_49 ();
 sg13g2_fill_2 FILLER_35_150 ();
 sg13g2_fill_1 FILLER_35_152 ();
 sg13g2_fill_2 FILLER_35_175 ();
 sg13g2_fill_1 FILLER_35_177 ();
 sg13g2_fill_2 FILLER_35_197 ();
 sg13g2_fill_2 FILLER_35_214 ();
 sg13g2_fill_1 FILLER_35_237 ();
 sg13g2_fill_2 FILLER_35_266 ();
 sg13g2_fill_1 FILLER_35_268 ();
 sg13g2_fill_2 FILLER_35_333 ();
 sg13g2_decap_4 FILLER_35_358 ();
 sg13g2_fill_2 FILLER_35_362 ();
 sg13g2_fill_1 FILLER_35_372 ();
 sg13g2_fill_2 FILLER_35_381 ();
 sg13g2_fill_2 FILLER_35_392 ();
 sg13g2_fill_1 FILLER_35_425 ();
 sg13g2_fill_2 FILLER_35_452 ();
 sg13g2_fill_1 FILLER_35_454 ();
 sg13g2_fill_2 FILLER_35_463 ();
 sg13g2_fill_1 FILLER_35_465 ();
 sg13g2_fill_2 FILLER_35_495 ();
 sg13g2_fill_2 FILLER_35_516 ();
 sg13g2_fill_2 FILLER_35_540 ();
 sg13g2_fill_2 FILLER_35_554 ();
 sg13g2_fill_1 FILLER_35_556 ();
 sg13g2_fill_2 FILLER_35_570 ();
 sg13g2_fill_1 FILLER_35_572 ();
 sg13g2_fill_2 FILLER_35_583 ();
 sg13g2_fill_1 FILLER_35_585 ();
 sg13g2_decap_4 FILLER_35_595 ();
 sg13g2_decap_4 FILLER_35_604 ();
 sg13g2_fill_2 FILLER_35_608 ();
 sg13g2_decap_8 FILLER_35_615 ();
 sg13g2_decap_4 FILLER_35_622 ();
 sg13g2_fill_1 FILLER_35_626 ();
 sg13g2_fill_2 FILLER_35_647 ();
 sg13g2_decap_4 FILLER_35_663 ();
 sg13g2_fill_2 FILLER_35_667 ();
 sg13g2_decap_4 FILLER_35_715 ();
 sg13g2_fill_1 FILLER_35_736 ();
 sg13g2_fill_2 FILLER_35_751 ();
 sg13g2_decap_4 FILLER_35_774 ();
 sg13g2_fill_1 FILLER_35_778 ();
 sg13g2_fill_1 FILLER_35_784 ();
 sg13g2_fill_2 FILLER_35_813 ();
 sg13g2_fill_1 FILLER_35_848 ();
 sg13g2_fill_2 FILLER_35_858 ();
 sg13g2_fill_1 FILLER_35_860 ();
 sg13g2_fill_2 FILLER_35_889 ();
 sg13g2_fill_2 FILLER_35_900 ();
 sg13g2_fill_1 FILLER_35_902 ();
 sg13g2_fill_2 FILLER_35_954 ();
 sg13g2_fill_1 FILLER_35_984 ();
 sg13g2_decap_4 FILLER_35_1080 ();
 sg13g2_fill_1 FILLER_35_1084 ();
 sg13g2_fill_2 FILLER_35_1088 ();
 sg13g2_fill_1 FILLER_35_1090 ();
 sg13g2_fill_2 FILLER_35_1100 ();
 sg13g2_fill_1 FILLER_35_1102 ();
 sg13g2_fill_1 FILLER_35_1117 ();
 sg13g2_fill_2 FILLER_35_1146 ();
 sg13g2_fill_1 FILLER_35_1263 ();
 sg13g2_fill_1 FILLER_35_1290 ();
 sg13g2_fill_2 FILLER_35_1338 ();
 sg13g2_decap_4 FILLER_35_1365 ();
 sg13g2_decap_4 FILLER_35_1373 ();
 sg13g2_fill_2 FILLER_35_1392 ();
 sg13g2_fill_1 FILLER_35_1394 ();
 sg13g2_fill_2 FILLER_35_1408 ();
 sg13g2_fill_1 FILLER_35_1410 ();
 sg13g2_decap_4 FILLER_35_1433 ();
 sg13g2_fill_1 FILLER_35_1437 ();
 sg13g2_decap_8 FILLER_35_1442 ();
 sg13g2_decap_8 FILLER_35_1449 ();
 sg13g2_fill_1 FILLER_35_1487 ();
 sg13g2_fill_1 FILLER_35_1500 ();
 sg13g2_fill_1 FILLER_35_1518 ();
 sg13g2_fill_2 FILLER_35_1544 ();
 sg13g2_fill_1 FILLER_35_1546 ();
 sg13g2_decap_8 FILLER_35_1551 ();
 sg13g2_fill_2 FILLER_35_1558 ();
 sg13g2_fill_2 FILLER_35_1573 ();
 sg13g2_fill_2 FILLER_35_1585 ();
 sg13g2_decap_8 FILLER_35_1591 ();
 sg13g2_decap_4 FILLER_35_1598 ();
 sg13g2_fill_2 FILLER_35_1602 ();
 sg13g2_fill_2 FILLER_35_1689 ();
 sg13g2_decap_4 FILLER_35_1727 ();
 sg13g2_fill_2 FILLER_35_1752 ();
 sg13g2_decap_8 FILLER_35_1782 ();
 sg13g2_fill_2 FILLER_35_1789 ();
 sg13g2_fill_1 FILLER_35_1791 ();
 sg13g2_fill_2 FILLER_35_1804 ();
 sg13g2_fill_1 FILLER_35_1806 ();
 sg13g2_fill_2 FILLER_35_1812 ();
 sg13g2_fill_1 FILLER_35_1823 ();
 sg13g2_fill_2 FILLER_35_1837 ();
 sg13g2_fill_2 FILLER_35_1856 ();
 sg13g2_fill_1 FILLER_35_1858 ();
 sg13g2_decap_8 FILLER_35_1881 ();
 sg13g2_decap_4 FILLER_35_1888 ();
 sg13g2_fill_2 FILLER_35_1892 ();
 sg13g2_decap_4 FILLER_35_1921 ();
 sg13g2_fill_1 FILLER_35_1925 ();
 sg13g2_fill_1 FILLER_35_1936 ();
 sg13g2_fill_2 FILLER_35_1948 ();
 sg13g2_fill_1 FILLER_35_1950 ();
 sg13g2_fill_1 FILLER_35_2019 ();
 sg13g2_fill_2 FILLER_35_2103 ();
 sg13g2_fill_2 FILLER_35_2119 ();
 sg13g2_fill_1 FILLER_35_2144 ();
 sg13g2_fill_2 FILLER_35_2158 ();
 sg13g2_decap_8 FILLER_35_2171 ();
 sg13g2_decap_4 FILLER_35_2178 ();
 sg13g2_fill_1 FILLER_35_2182 ();
 sg13g2_fill_2 FILLER_35_2214 ();
 sg13g2_fill_1 FILLER_35_2216 ();
 sg13g2_fill_2 FILLER_35_2231 ();
 sg13g2_fill_1 FILLER_35_2233 ();
 sg13g2_fill_1 FILLER_35_2258 ();
 sg13g2_fill_2 FILLER_35_2264 ();
 sg13g2_decap_8 FILLER_35_2290 ();
 sg13g2_decap_4 FILLER_35_2297 ();
 sg13g2_fill_2 FILLER_35_2301 ();
 sg13g2_fill_1 FILLER_35_2312 ();
 sg13g2_fill_2 FILLER_35_2331 ();
 sg13g2_fill_1 FILLER_35_2342 ();
 sg13g2_fill_1 FILLER_35_2348 ();
 sg13g2_fill_1 FILLER_35_2376 ();
 sg13g2_decap_8 FILLER_35_2393 ();
 sg13g2_decap_4 FILLER_35_2400 ();
 sg13g2_fill_1 FILLER_35_2404 ();
 sg13g2_fill_2 FILLER_35_2438 ();
 sg13g2_decap_4 FILLER_35_2467 ();
 sg13g2_fill_1 FILLER_35_2471 ();
 sg13g2_fill_2 FILLER_35_2489 ();
 sg13g2_fill_1 FILLER_35_2491 ();
 sg13g2_decap_4 FILLER_35_2511 ();
 sg13g2_fill_2 FILLER_35_2543 ();
 sg13g2_fill_1 FILLER_35_2545 ();
 sg13g2_fill_2 FILLER_35_2555 ();
 sg13g2_fill_1 FILLER_35_2593 ();
 sg13g2_fill_2 FILLER_35_2600 ();
 sg13g2_decap_4 FILLER_35_2610 ();
 sg13g2_fill_1 FILLER_35_2627 ();
 sg13g2_fill_1 FILLER_35_2765 ();
 sg13g2_fill_2 FILLER_35_2835 ();
 sg13g2_fill_1 FILLER_35_2846 ();
 sg13g2_fill_1 FILLER_35_2879 ();
 sg13g2_fill_2 FILLER_35_2913 ();
 sg13g2_fill_1 FILLER_35_2928 ();
 sg13g2_fill_2 FILLER_35_2951 ();
 sg13g2_fill_1 FILLER_35_2953 ();
 sg13g2_fill_2 FILLER_35_2988 ();
 sg13g2_fill_2 FILLER_35_3005 ();
 sg13g2_fill_2 FILLER_35_3054 ();
 sg13g2_fill_1 FILLER_35_3137 ();
 sg13g2_fill_2 FILLER_35_3142 ();
 sg13g2_decap_4 FILLER_35_3170 ();
 sg13g2_fill_2 FILLER_35_3174 ();
 sg13g2_fill_1 FILLER_35_3201 ();
 sg13g2_fill_2 FILLER_35_3294 ();
 sg13g2_fill_1 FILLER_35_3296 ();
 sg13g2_fill_2 FILLER_35_3379 ();
 sg13g2_fill_1 FILLER_35_3409 ();
 sg13g2_fill_2 FILLER_35_3423 ();
 sg13g2_fill_1 FILLER_35_3425 ();
 sg13g2_decap_8 FILLER_35_3454 ();
 sg13g2_decap_4 FILLER_35_3461 ();
 sg13g2_fill_2 FILLER_35_3465 ();
 sg13g2_fill_1 FILLER_35_3487 ();
 sg13g2_decap_4 FILLER_35_3520 ();
 sg13g2_fill_1 FILLER_35_3524 ();
 sg13g2_fill_1 FILLER_35_3546 ();
 sg13g2_fill_1 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_34 ();
 sg13g2_fill_2 FILLER_36_78 ();
 sg13g2_fill_1 FILLER_36_80 ();
 sg13g2_fill_2 FILLER_36_100 ();
 sg13g2_fill_2 FILLER_36_225 ();
 sg13g2_fill_2 FILLER_36_290 ();
 sg13g2_fill_1 FILLER_36_292 ();
 sg13g2_fill_1 FILLER_36_298 ();
 sg13g2_fill_2 FILLER_36_321 ();
 sg13g2_fill_1 FILLER_36_323 ();
 sg13g2_decap_8 FILLER_36_351 ();
 sg13g2_decap_4 FILLER_36_384 ();
 sg13g2_fill_1 FILLER_36_388 ();
 sg13g2_fill_2 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_433 ();
 sg13g2_fill_2 FILLER_36_445 ();
 sg13g2_decap_4 FILLER_36_455 ();
 sg13g2_fill_2 FILLER_36_464 ();
 sg13g2_fill_2 FILLER_36_485 ();
 sg13g2_fill_1 FILLER_36_499 ();
 sg13g2_fill_2 FILLER_36_588 ();
 sg13g2_decap_4 FILLER_36_601 ();
 sg13g2_fill_2 FILLER_36_620 ();
 sg13g2_fill_2 FILLER_36_657 ();
 sg13g2_fill_2 FILLER_36_685 ();
 sg13g2_fill_1 FILLER_36_687 ();
 sg13g2_fill_1 FILLER_36_713 ();
 sg13g2_fill_2 FILLER_36_727 ();
 sg13g2_fill_1 FILLER_36_729 ();
 sg13g2_decap_4 FILLER_36_740 ();
 sg13g2_fill_1 FILLER_36_744 ();
 sg13g2_decap_4 FILLER_36_753 ();
 sg13g2_fill_1 FILLER_36_757 ();
 sg13g2_decap_8 FILLER_36_766 ();
 sg13g2_fill_2 FILLER_36_773 ();
 sg13g2_fill_1 FILLER_36_775 ();
 sg13g2_fill_2 FILLER_36_781 ();
 sg13g2_decap_4 FILLER_36_787 ();
 sg13g2_fill_2 FILLER_36_795 ();
 sg13g2_fill_1 FILLER_36_797 ();
 sg13g2_fill_1 FILLER_36_807 ();
 sg13g2_fill_2 FILLER_36_838 ();
 sg13g2_fill_1 FILLER_36_840 ();
 sg13g2_fill_2 FILLER_36_853 ();
 sg13g2_fill_1 FILLER_36_855 ();
 sg13g2_fill_1 FILLER_36_862 ();
 sg13g2_fill_1 FILLER_36_884 ();
 sg13g2_fill_2 FILLER_36_898 ();
 sg13g2_decap_8 FILLER_36_912 ();
 sg13g2_decap_8 FILLER_36_919 ();
 sg13g2_decap_4 FILLER_36_926 ();
 sg13g2_decap_8 FILLER_36_944 ();
 sg13g2_fill_2 FILLER_36_951 ();
 sg13g2_fill_1 FILLER_36_953 ();
 sg13g2_fill_2 FILLER_36_1002 ();
 sg13g2_decap_4 FILLER_36_1016 ();
 sg13g2_fill_1 FILLER_36_1020 ();
 sg13g2_decap_4 FILLER_36_1046 ();
 sg13g2_fill_1 FILLER_36_1050 ();
 sg13g2_decap_4 FILLER_36_1055 ();
 sg13g2_fill_1 FILLER_36_1059 ();
 sg13g2_decap_4 FILLER_36_1074 ();
 sg13g2_fill_1 FILLER_36_1138 ();
 sg13g2_fill_2 FILLER_36_1165 ();
 sg13g2_fill_2 FILLER_36_1177 ();
 sg13g2_fill_1 FILLER_36_1179 ();
 sg13g2_fill_1 FILLER_36_1224 ();
 sg13g2_fill_2 FILLER_36_1303 ();
 sg13g2_fill_1 FILLER_36_1305 ();
 sg13g2_fill_1 FILLER_36_1319 ();
 sg13g2_decap_4 FILLER_36_1346 ();
 sg13g2_fill_2 FILLER_36_1378 ();
 sg13g2_decap_4 FILLER_36_1408 ();
 sg13g2_fill_2 FILLER_36_1412 ();
 sg13g2_fill_2 FILLER_36_1431 ();
 sg13g2_fill_1 FILLER_36_1466 ();
 sg13g2_fill_2 FILLER_36_1473 ();
 sg13g2_fill_1 FILLER_36_1475 ();
 sg13g2_decap_4 FILLER_36_1480 ();
 sg13g2_fill_1 FILLER_36_1505 ();
 sg13g2_decap_8 FILLER_36_1522 ();
 sg13g2_fill_1 FILLER_36_1546 ();
 sg13g2_decap_8 FILLER_36_1555 ();
 sg13g2_fill_2 FILLER_36_1562 ();
 sg13g2_fill_1 FILLER_36_1564 ();
 sg13g2_decap_8 FILLER_36_1596 ();
 sg13g2_fill_1 FILLER_36_1603 ();
 sg13g2_fill_2 FILLER_36_1619 ();
 sg13g2_fill_1 FILLER_36_1621 ();
 sg13g2_decap_4 FILLER_36_1626 ();
 sg13g2_fill_2 FILLER_36_1630 ();
 sg13g2_decap_4 FILLER_36_1637 ();
 sg13g2_fill_1 FILLER_36_1641 ();
 sg13g2_fill_2 FILLER_36_1655 ();
 sg13g2_decap_8 FILLER_36_1689 ();
 sg13g2_fill_1 FILLER_36_1701 ();
 sg13g2_fill_2 FILLER_36_1707 ();
 sg13g2_fill_1 FILLER_36_1709 ();
 sg13g2_decap_8 FILLER_36_1727 ();
 sg13g2_fill_1 FILLER_36_1734 ();
 sg13g2_fill_1 FILLER_36_1750 ();
 sg13g2_fill_2 FILLER_36_1768 ();
 sg13g2_fill_1 FILLER_36_1770 ();
 sg13g2_fill_2 FILLER_36_1776 ();
 sg13g2_decap_8 FILLER_36_1786 ();
 sg13g2_decap_4 FILLER_36_1793 ();
 sg13g2_fill_1 FILLER_36_1797 ();
 sg13g2_fill_2 FILLER_36_1815 ();
 sg13g2_fill_1 FILLER_36_1817 ();
 sg13g2_decap_4 FILLER_36_1831 ();
 sg13g2_fill_2 FILLER_36_1835 ();
 sg13g2_fill_2 FILLER_36_1865 ();
 sg13g2_fill_1 FILLER_36_1867 ();
 sg13g2_fill_2 FILLER_36_1874 ();
 sg13g2_fill_1 FILLER_36_1906 ();
 sg13g2_decap_8 FILLER_36_1920 ();
 sg13g2_decap_4 FILLER_36_1927 ();
 sg13g2_decap_8 FILLER_36_1951 ();
 sg13g2_decap_4 FILLER_36_1970 ();
 sg13g2_decap_8 FILLER_36_1978 ();
 sg13g2_fill_2 FILLER_36_1985 ();
 sg13g2_fill_1 FILLER_36_1987 ();
 sg13g2_decap_8 FILLER_36_1991 ();
 sg13g2_decap_8 FILLER_36_1998 ();
 sg13g2_decap_8 FILLER_36_2021 ();
 sg13g2_fill_1 FILLER_36_2028 ();
 sg13g2_fill_1 FILLER_36_2037 ();
 sg13g2_fill_2 FILLER_36_2051 ();
 sg13g2_fill_1 FILLER_36_2053 ();
 sg13g2_decap_8 FILLER_36_2082 ();
 sg13g2_fill_2 FILLER_36_2089 ();
 sg13g2_fill_1 FILLER_36_2091 ();
 sg13g2_fill_1 FILLER_36_2101 ();
 sg13g2_fill_1 FILLER_36_2110 ();
 sg13g2_fill_1 FILLER_36_2115 ();
 sg13g2_decap_8 FILLER_36_2144 ();
 sg13g2_decap_4 FILLER_36_2151 ();
 sg13g2_decap_8 FILLER_36_2200 ();
 sg13g2_decap_4 FILLER_36_2215 ();
 sg13g2_decap_4 FILLER_36_2231 ();
 sg13g2_fill_1 FILLER_36_2235 ();
 sg13g2_fill_2 FILLER_36_2251 ();
 sg13g2_fill_2 FILLER_36_2270 ();
 sg13g2_decap_4 FILLER_36_2295 ();
 sg13g2_fill_1 FILLER_36_2299 ();
 sg13g2_fill_1 FILLER_36_2303 ();
 sg13g2_fill_2 FILLER_36_2322 ();
 sg13g2_fill_1 FILLER_36_2332 ();
 sg13g2_fill_2 FILLER_36_2343 ();
 sg13g2_fill_1 FILLER_36_2345 ();
 sg13g2_fill_2 FILLER_36_2383 ();
 sg13g2_fill_1 FILLER_36_2385 ();
 sg13g2_decap_8 FILLER_36_2400 ();
 sg13g2_decap_8 FILLER_36_2407 ();
 sg13g2_fill_1 FILLER_36_2414 ();
 sg13g2_fill_2 FILLER_36_2424 ();
 sg13g2_fill_1 FILLER_36_2439 ();
 sg13g2_fill_2 FILLER_36_2473 ();
 sg13g2_fill_2 FILLER_36_2479 ();
 sg13g2_fill_1 FILLER_36_2481 ();
 sg13g2_fill_1 FILLER_36_2539 ();
 sg13g2_fill_2 FILLER_36_2584 ();
 sg13g2_fill_2 FILLER_36_2591 ();
 sg13g2_fill_1 FILLER_36_2613 ();
 sg13g2_fill_2 FILLER_36_2636 ();
 sg13g2_decap_4 FILLER_36_2651 ();
 sg13g2_decap_8 FILLER_36_2660 ();
 sg13g2_decap_4 FILLER_36_2667 ();
 sg13g2_fill_1 FILLER_36_2671 ();
 sg13g2_fill_1 FILLER_36_2718 ();
 sg13g2_fill_1 FILLER_36_2756 ();
 sg13g2_fill_1 FILLER_36_2843 ();
 sg13g2_fill_1 FILLER_36_2858 ();
 sg13g2_fill_2 FILLER_36_2894 ();
 sg13g2_fill_1 FILLER_36_2896 ();
 sg13g2_fill_2 FILLER_36_2928 ();
 sg13g2_fill_2 FILLER_36_2986 ();
 sg13g2_fill_1 FILLER_36_2996 ();
 sg13g2_fill_1 FILLER_36_3078 ();
 sg13g2_fill_1 FILLER_36_3116 ();
 sg13g2_fill_2 FILLER_36_3121 ();
 sg13g2_fill_1 FILLER_36_3123 ();
 sg13g2_fill_2 FILLER_36_3200 ();
 sg13g2_decap_8 FILLER_36_3207 ();
 sg13g2_decap_4 FILLER_36_3214 ();
 sg13g2_fill_1 FILLER_36_3218 ();
 sg13g2_decap_8 FILLER_36_3227 ();
 sg13g2_fill_2 FILLER_36_3256 ();
 sg13g2_fill_1 FILLER_36_3276 ();
 sg13g2_fill_2 FILLER_36_3321 ();
 sg13g2_fill_2 FILLER_36_3350 ();
 sg13g2_fill_1 FILLER_36_3352 ();
 sg13g2_fill_1 FILLER_36_3390 ();
 sg13g2_fill_1 FILLER_36_3436 ();
 sg13g2_decap_8 FILLER_36_3463 ();
 sg13g2_decap_8 FILLER_36_3486 ();
 sg13g2_fill_2 FILLER_36_3493 ();
 sg13g2_fill_1 FILLER_36_3495 ();
 sg13g2_fill_1 FILLER_36_3506 ();
 sg13g2_fill_2 FILLER_36_3549 ();
 sg13g2_fill_1 FILLER_36_3551 ();
 sg13g2_fill_2 FILLER_36_3565 ();
 sg13g2_fill_1 FILLER_36_3567 ();
 sg13g2_fill_2 FILLER_36_3577 ();
 sg13g2_fill_1 FILLER_36_3579 ();
 sg13g2_decap_4 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_4 ();
 sg13g2_fill_2 FILLER_37_39 ();
 sg13g2_fill_1 FILLER_37_41 ();
 sg13g2_fill_2 FILLER_37_50 ();
 sg13g2_fill_1 FILLER_37_52 ();
 sg13g2_decap_8 FILLER_37_58 ();
 sg13g2_fill_1 FILLER_37_65 ();
 sg13g2_decap_4 FILLER_37_71 ();
 sg13g2_fill_1 FILLER_37_75 ();
 sg13g2_fill_2 FILLER_37_79 ();
 sg13g2_fill_2 FILLER_37_109 ();
 sg13g2_fill_2 FILLER_37_167 ();
 sg13g2_fill_1 FILLER_37_169 ();
 sg13g2_fill_2 FILLER_37_179 ();
 sg13g2_fill_2 FILLER_37_190 ();
 sg13g2_fill_2 FILLER_37_210 ();
 sg13g2_fill_1 FILLER_37_212 ();
 sg13g2_fill_2 FILLER_37_244 ();
 sg13g2_fill_2 FILLER_37_319 ();
 sg13g2_fill_1 FILLER_37_350 ();
 sg13g2_decap_4 FILLER_37_359 ();
 sg13g2_fill_2 FILLER_37_400 ();
 sg13g2_decap_4 FILLER_37_427 ();
 sg13g2_fill_2 FILLER_37_431 ();
 sg13g2_fill_1 FILLER_37_456 ();
 sg13g2_decap_4 FILLER_37_460 ();
 sg13g2_fill_2 FILLER_37_464 ();
 sg13g2_decap_4 FILLER_37_490 ();
 sg13g2_fill_1 FILLER_37_512 ();
 sg13g2_decap_8 FILLER_37_517 ();
 sg13g2_decap_8 FILLER_37_524 ();
 sg13g2_fill_1 FILLER_37_536 ();
 sg13g2_fill_2 FILLER_37_558 ();
 sg13g2_decap_8 FILLER_37_568 ();
 sg13g2_fill_1 FILLER_37_575 ();
 sg13g2_fill_1 FILLER_37_590 ();
 sg13g2_fill_1 FILLER_37_596 ();
 sg13g2_fill_2 FILLER_37_609 ();
 sg13g2_decap_8 FILLER_37_623 ();
 sg13g2_fill_2 FILLER_37_630 ();
 sg13g2_fill_1 FILLER_37_636 ();
 sg13g2_decap_8 FILLER_37_642 ();
 sg13g2_decap_4 FILLER_37_649 ();
 sg13g2_fill_2 FILLER_37_653 ();
 sg13g2_decap_8 FILLER_37_664 ();
 sg13g2_fill_2 FILLER_37_671 ();
 sg13g2_fill_1 FILLER_37_673 ();
 sg13g2_fill_1 FILLER_37_687 ();
 sg13g2_fill_1 FILLER_37_708 ();
 sg13g2_fill_2 FILLER_37_723 ();
 sg13g2_fill_1 FILLER_37_725 ();
 sg13g2_decap_4 FILLER_37_751 ();
 sg13g2_fill_1 FILLER_37_770 ();
 sg13g2_fill_2 FILLER_37_776 ();
 sg13g2_fill_1 FILLER_37_778 ();
 sg13g2_fill_2 FILLER_37_783 ();
 sg13g2_fill_1 FILLER_37_785 ();
 sg13g2_fill_1 FILLER_37_814 ();
 sg13g2_fill_2 FILLER_37_837 ();
 sg13g2_fill_1 FILLER_37_839 ();
 sg13g2_fill_2 FILLER_37_853 ();
 sg13g2_decap_4 FILLER_37_871 ();
 sg13g2_fill_1 FILLER_37_891 ();
 sg13g2_fill_2 FILLER_37_908 ();
 sg13g2_fill_1 FILLER_37_910 ();
 sg13g2_decap_8 FILLER_37_921 ();
 sg13g2_fill_1 FILLER_37_928 ();
 sg13g2_fill_2 FILLER_37_950 ();
 sg13g2_fill_1 FILLER_37_952 ();
 sg13g2_fill_2 FILLER_37_988 ();
 sg13g2_fill_1 FILLER_37_990 ();
 sg13g2_fill_1 FILLER_37_1004 ();
 sg13g2_fill_2 FILLER_37_1011 ();
 sg13g2_decap_4 FILLER_37_1030 ();
 sg13g2_decap_8 FILLER_37_1046 ();
 sg13g2_fill_1 FILLER_37_1053 ();
 sg13g2_fill_2 FILLER_37_1058 ();
 sg13g2_fill_1 FILLER_37_1060 ();
 sg13g2_fill_1 FILLER_37_1089 ();
 sg13g2_fill_2 FILLER_37_1110 ();
 sg13g2_fill_1 FILLER_37_1128 ();
 sg13g2_fill_1 FILLER_37_1155 ();
 sg13g2_fill_2 FILLER_37_1162 ();
 sg13g2_fill_1 FILLER_37_1164 ();
 sg13g2_fill_2 FILLER_37_1196 ();
 sg13g2_fill_1 FILLER_37_1198 ();
 sg13g2_fill_2 FILLER_37_1216 ();
 sg13g2_fill_1 FILLER_37_1218 ();
 sg13g2_fill_1 FILLER_37_1224 ();
 sg13g2_fill_1 FILLER_37_1229 ();
 sg13g2_fill_1 FILLER_37_1253 ();
 sg13g2_fill_2 FILLER_37_1288 ();
 sg13g2_fill_1 FILLER_37_1290 ();
 sg13g2_fill_2 FILLER_37_1307 ();
 sg13g2_fill_2 FILLER_37_1322 ();
 sg13g2_fill_1 FILLER_37_1324 ();
 sg13g2_decap_4 FILLER_37_1342 ();
 sg13g2_fill_2 FILLER_37_1346 ();
 sg13g2_fill_2 FILLER_37_1370 ();
 sg13g2_fill_1 FILLER_37_1372 ();
 sg13g2_decap_8 FILLER_37_1399 ();
 sg13g2_fill_2 FILLER_37_1406 ();
 sg13g2_decap_8 FILLER_37_1431 ();
 sg13g2_decap_8 FILLER_37_1438 ();
 sg13g2_decap_4 FILLER_37_1445 ();
 sg13g2_fill_1 FILLER_37_1449 ();
 sg13g2_fill_2 FILLER_37_1468 ();
 sg13g2_fill_1 FILLER_37_1470 ();
 sg13g2_decap_8 FILLER_37_1502 ();
 sg13g2_decap_4 FILLER_37_1509 ();
 sg13g2_fill_1 FILLER_37_1520 ();
 sg13g2_decap_8 FILLER_37_1526 ();
 sg13g2_fill_2 FILLER_37_1533 ();
 sg13g2_fill_1 FILLER_37_1552 ();
 sg13g2_decap_4 FILLER_37_1561 ();
 sg13g2_fill_1 FILLER_37_1565 ();
 sg13g2_fill_2 FILLER_37_1579 ();
 sg13g2_decap_8 FILLER_37_1599 ();
 sg13g2_decap_4 FILLER_37_1606 ();
 sg13g2_fill_2 FILLER_37_1610 ();
 sg13g2_decap_8 FILLER_37_1629 ();
 sg13g2_fill_2 FILLER_37_1636 ();
 sg13g2_decap_8 FILLER_37_1646 ();
 sg13g2_decap_8 FILLER_37_1653 ();
 sg13g2_decap_4 FILLER_37_1690 ();
 sg13g2_fill_2 FILLER_37_1704 ();
 sg13g2_decap_8 FILLER_37_1714 ();
 sg13g2_decap_8 FILLER_37_1731 ();
 sg13g2_decap_4 FILLER_37_1743 ();
 sg13g2_fill_1 FILLER_37_1747 ();
 sg13g2_fill_2 FILLER_37_1761 ();
 sg13g2_fill_1 FILLER_37_1763 ();
 sg13g2_fill_1 FILLER_37_1777 ();
 sg13g2_decap_4 FILLER_37_1783 ();
 sg13g2_fill_1 FILLER_37_1787 ();
 sg13g2_decap_8 FILLER_37_1815 ();
 sg13g2_decap_4 FILLER_37_1822 ();
 sg13g2_decap_4 FILLER_37_1831 ();
 sg13g2_fill_2 FILLER_37_1844 ();
 sg13g2_decap_8 FILLER_37_1870 ();
 sg13g2_decap_4 FILLER_37_1877 ();
 sg13g2_decap_4 FILLER_37_1891 ();
 sg13g2_fill_1 FILLER_37_1895 ();
 sg13g2_fill_2 FILLER_37_1905 ();
 sg13g2_decap_8 FILLER_37_1919 ();
 sg13g2_decap_8 FILLER_37_1926 ();
 sg13g2_decap_8 FILLER_37_1933 ();
 sg13g2_fill_2 FILLER_37_1940 ();
 sg13g2_fill_1 FILLER_37_1942 ();
 sg13g2_fill_2 FILLER_37_1953 ();
 sg13g2_fill_1 FILLER_37_1959 ();
 sg13g2_decap_4 FILLER_37_1968 ();
 sg13g2_fill_1 FILLER_37_1972 ();
 sg13g2_decap_4 FILLER_37_1978 ();
 sg13g2_fill_1 FILLER_37_2024 ();
 sg13g2_decap_4 FILLER_37_2091 ();
 sg13g2_fill_2 FILLER_37_2095 ();
 sg13g2_fill_1 FILLER_37_2110 ();
 sg13g2_fill_2 FILLER_37_2157 ();
 sg13g2_fill_1 FILLER_37_2192 ();
 sg13g2_fill_2 FILLER_37_2219 ();
 sg13g2_decap_8 FILLER_37_2235 ();
 sg13g2_fill_2 FILLER_37_2242 ();
 sg13g2_fill_1 FILLER_37_2244 ();
 sg13g2_fill_2 FILLER_37_2293 ();
 sg13g2_fill_1 FILLER_37_2304 ();
 sg13g2_decap_8 FILLER_37_2315 ();
 sg13g2_decap_4 FILLER_37_2322 ();
 sg13g2_fill_2 FILLER_37_2326 ();
 sg13g2_fill_2 FILLER_37_2345 ();
 sg13g2_fill_1 FILLER_37_2347 ();
 sg13g2_fill_1 FILLER_37_2364 ();
 sg13g2_fill_2 FILLER_37_2370 ();
 sg13g2_fill_1 FILLER_37_2385 ();
 sg13g2_decap_8 FILLER_37_2399 ();
 sg13g2_decap_4 FILLER_37_2406 ();
 sg13g2_fill_1 FILLER_37_2410 ();
 sg13g2_fill_1 FILLER_37_2428 ();
 sg13g2_decap_4 FILLER_37_2440 ();
 sg13g2_decap_8 FILLER_37_2457 ();
 sg13g2_fill_2 FILLER_37_2464 ();
 sg13g2_fill_1 FILLER_37_2466 ();
 sg13g2_decap_8 FILLER_37_2481 ();
 sg13g2_fill_2 FILLER_37_2488 ();
 sg13g2_fill_2 FILLER_37_2494 ();
 sg13g2_fill_1 FILLER_37_2496 ();
 sg13g2_fill_2 FILLER_37_2510 ();
 sg13g2_fill_1 FILLER_37_2512 ();
 sg13g2_fill_1 FILLER_37_2539 ();
 sg13g2_fill_1 FILLER_37_2545 ();
 sg13g2_fill_1 FILLER_37_2559 ();
 sg13g2_fill_1 FILLER_37_2574 ();
 sg13g2_fill_1 FILLER_37_2581 ();
 sg13g2_fill_2 FILLER_37_2607 ();
 sg13g2_fill_2 FILLER_37_2621 ();
 sg13g2_fill_2 FILLER_37_2635 ();
 sg13g2_fill_1 FILLER_37_2637 ();
 sg13g2_decap_4 FILLER_37_2664 ();
 sg13g2_fill_1 FILLER_37_2668 ();
 sg13g2_fill_2 FILLER_37_2690 ();
 sg13g2_fill_1 FILLER_37_2692 ();
 sg13g2_fill_2 FILLER_37_2702 ();
 sg13g2_fill_2 FILLER_37_2726 ();
 sg13g2_fill_1 FILLER_37_2728 ();
 sg13g2_fill_1 FILLER_37_2791 ();
 sg13g2_fill_2 FILLER_37_2818 ();
 sg13g2_fill_1 FILLER_37_2899 ();
 sg13g2_fill_2 FILLER_37_2964 ();
 sg13g2_fill_1 FILLER_37_2966 ();
 sg13g2_fill_1 FILLER_37_3004 ();
 sg13g2_fill_1 FILLER_37_3084 ();
 sg13g2_fill_2 FILLER_37_3090 ();
 sg13g2_fill_1 FILLER_37_3092 ();
 sg13g2_decap_4 FILLER_37_3124 ();
 sg13g2_fill_2 FILLER_37_3128 ();
 sg13g2_decap_8 FILLER_37_3143 ();
 sg13g2_decap_8 FILLER_37_3150 ();
 sg13g2_fill_1 FILLER_37_3157 ();
 sg13g2_decap_8 FILLER_37_3166 ();
 sg13g2_decap_8 FILLER_37_3173 ();
 sg13g2_fill_2 FILLER_37_3267 ();
 sg13g2_fill_2 FILLER_37_3325 ();
 sg13g2_fill_1 FILLER_37_3327 ();
 sg13g2_fill_2 FILLER_37_3356 ();
 sg13g2_fill_1 FILLER_37_3358 ();
 sg13g2_fill_2 FILLER_37_3368 ();
 sg13g2_decap_4 FILLER_37_3411 ();
 sg13g2_fill_1 FILLER_37_3415 ();
 sg13g2_decap_8 FILLER_37_3420 ();
 sg13g2_fill_2 FILLER_37_3427 ();
 sg13g2_fill_1 FILLER_37_3429 ();
 sg13g2_fill_2 FILLER_37_3443 ();
 sg13g2_fill_1 FILLER_37_3445 ();
 sg13g2_decap_4 FILLER_37_3465 ();
 sg13g2_fill_1 FILLER_37_3506 ();
 sg13g2_fill_1 FILLER_37_3541 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_44 ();
 sg13g2_fill_1 FILLER_38_46 ();
 sg13g2_fill_2 FILLER_38_68 ();
 sg13g2_fill_2 FILLER_38_85 ();
 sg13g2_fill_1 FILLER_38_87 ();
 sg13g2_fill_2 FILLER_38_100 ();
 sg13g2_fill_1 FILLER_38_102 ();
 sg13g2_fill_2 FILLER_38_244 ();
 sg13g2_fill_1 FILLER_38_246 ();
 sg13g2_fill_2 FILLER_38_257 ();
 sg13g2_fill_1 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_269 ();
 sg13g2_fill_2 FILLER_38_276 ();
 sg13g2_fill_1 FILLER_38_278 ();
 sg13g2_decap_4 FILLER_38_300 ();
 sg13g2_fill_1 FILLER_38_304 ();
 sg13g2_fill_1 FILLER_38_327 ();
 sg13g2_decap_4 FILLER_38_345 ();
 sg13g2_fill_1 FILLER_38_349 ();
 sg13g2_decap_8 FILLER_38_382 ();
 sg13g2_fill_2 FILLER_38_389 ();
 sg13g2_fill_1 FILLER_38_391 ();
 sg13g2_fill_2 FILLER_38_397 ();
 sg13g2_fill_1 FILLER_38_399 ();
 sg13g2_fill_1 FILLER_38_418 ();
 sg13g2_fill_2 FILLER_38_468 ();
 sg13g2_fill_1 FILLER_38_470 ();
 sg13g2_fill_1 FILLER_38_475 ();
 sg13g2_decap_4 FILLER_38_480 ();
 sg13g2_fill_1 FILLER_38_494 ();
 sg13g2_decap_8 FILLER_38_513 ();
 sg13g2_decap_4 FILLER_38_520 ();
 sg13g2_fill_1 FILLER_38_524 ();
 sg13g2_fill_1 FILLER_38_529 ();
 sg13g2_fill_1 FILLER_38_535 ();
 sg13g2_decap_4 FILLER_38_565 ();
 sg13g2_fill_1 FILLER_38_569 ();
 sg13g2_decap_8 FILLER_38_581 ();
 sg13g2_decap_8 FILLER_38_588 ();
 sg13g2_fill_2 FILLER_38_595 ();
 sg13g2_fill_1 FILLER_38_597 ();
 sg13g2_decap_4 FILLER_38_603 ();
 sg13g2_fill_1 FILLER_38_607 ();
 sg13g2_fill_1 FILLER_38_616 ();
 sg13g2_decap_8 FILLER_38_625 ();
 sg13g2_fill_2 FILLER_38_632 ();
 sg13g2_fill_1 FILLER_38_634 ();
 sg13g2_fill_2 FILLER_38_647 ();
 sg13g2_fill_1 FILLER_38_649 ();
 sg13g2_fill_1 FILLER_38_654 ();
 sg13g2_fill_2 FILLER_38_660 ();
 sg13g2_fill_1 FILLER_38_662 ();
 sg13g2_fill_2 FILLER_38_694 ();
 sg13g2_fill_1 FILLER_38_708 ();
 sg13g2_fill_1 FILLER_38_714 ();
 sg13g2_fill_2 FILLER_38_723 ();
 sg13g2_fill_2 FILLER_38_759 ();
 sg13g2_fill_1 FILLER_38_761 ();
 sg13g2_fill_2 FILLER_38_766 ();
 sg13g2_decap_8 FILLER_38_775 ();
 sg13g2_decap_4 FILLER_38_782 ();
 sg13g2_fill_2 FILLER_38_790 ();
 sg13g2_decap_8 FILLER_38_796 ();
 sg13g2_fill_2 FILLER_38_803 ();
 sg13g2_fill_1 FILLER_38_805 ();
 sg13g2_fill_1 FILLER_38_825 ();
 sg13g2_decap_8 FILLER_38_851 ();
 sg13g2_fill_1 FILLER_38_868 ();
 sg13g2_fill_2 FILLER_38_874 ();
 sg13g2_fill_2 FILLER_38_885 ();
 sg13g2_fill_1 FILLER_38_887 ();
 sg13g2_fill_1 FILLER_38_939 ();
 sg13g2_fill_2 FILLER_38_953 ();
 sg13g2_fill_1 FILLER_38_995 ();
 sg13g2_decap_4 FILLER_38_1005 ();
 sg13g2_fill_1 FILLER_38_1035 ();
 sg13g2_decap_4 FILLER_38_1040 ();
 sg13g2_fill_2 FILLER_38_1044 ();
 sg13g2_decap_8 FILLER_38_1051 ();
 sg13g2_fill_2 FILLER_38_1084 ();
 sg13g2_fill_2 FILLER_38_1108 ();
 sg13g2_fill_1 FILLER_38_1110 ();
 sg13g2_decap_8 FILLER_38_1132 ();
 sg13g2_fill_1 FILLER_38_1139 ();
 sg13g2_decap_4 FILLER_38_1159 ();
 sg13g2_fill_2 FILLER_38_1163 ();
 sg13g2_fill_1 FILLER_38_1191 ();
 sg13g2_fill_1 FILLER_38_1209 ();
 sg13g2_fill_2 FILLER_38_1220 ();
 sg13g2_fill_1 FILLER_38_1222 ();
 sg13g2_fill_2 FILLER_38_1305 ();
 sg13g2_fill_1 FILLER_38_1307 ();
 sg13g2_decap_4 FILLER_38_1350 ();
 sg13g2_fill_1 FILLER_38_1354 ();
 sg13g2_fill_2 FILLER_38_1359 ();
 sg13g2_decap_8 FILLER_38_1370 ();
 sg13g2_decap_4 FILLER_38_1377 ();
 sg13g2_fill_2 FILLER_38_1390 ();
 sg13g2_fill_1 FILLER_38_1401 ();
 sg13g2_decap_8 FILLER_38_1429 ();
 sg13g2_fill_1 FILLER_38_1436 ();
 sg13g2_decap_4 FILLER_38_1488 ();
 sg13g2_fill_2 FILLER_38_1492 ();
 sg13g2_fill_1 FILLER_38_1532 ();
 sg13g2_fill_1 FILLER_38_1542 ();
 sg13g2_decap_8 FILLER_38_1561 ();
 sg13g2_fill_2 FILLER_38_1580 ();
 sg13g2_fill_1 FILLER_38_1582 ();
 sg13g2_fill_1 FILLER_38_1601 ();
 sg13g2_fill_2 FILLER_38_1651 ();
 sg13g2_decap_8 FILLER_38_1683 ();
 sg13g2_decap_8 FILLER_38_1724 ();
 sg13g2_fill_1 FILLER_38_1731 ();
 sg13g2_fill_1 FILLER_38_1750 ();
 sg13g2_fill_1 FILLER_38_1754 ();
 sg13g2_fill_2 FILLER_38_1768 ();
 sg13g2_fill_1 FILLER_38_1770 ();
 sg13g2_decap_4 FILLER_38_1786 ();
 sg13g2_decap_4 FILLER_38_1823 ();
 sg13g2_decap_8 FILLER_38_1843 ();
 sg13g2_fill_2 FILLER_38_1850 ();
 sg13g2_fill_1 FILLER_38_1852 ();
 sg13g2_decap_4 FILLER_38_1866 ();
 sg13g2_fill_2 FILLER_38_1870 ();
 sg13g2_decap_8 FILLER_38_1892 ();
 sg13g2_decap_4 FILLER_38_1899 ();
 sg13g2_fill_2 FILLER_38_1916 ();
 sg13g2_fill_1 FILLER_38_1918 ();
 sg13g2_decap_4 FILLER_38_1928 ();
 sg13g2_fill_1 FILLER_38_1932 ();
 sg13g2_decap_8 FILLER_38_1937 ();
 sg13g2_decap_8 FILLER_38_1944 ();
 sg13g2_fill_2 FILLER_38_1951 ();
 sg13g2_fill_1 FILLER_38_1953 ();
 sg13g2_decap_4 FILLER_38_1978 ();
 sg13g2_fill_2 FILLER_38_1982 ();
 sg13g2_decap_4 FILLER_38_1987 ();
 sg13g2_fill_2 FILLER_38_1991 ();
 sg13g2_fill_2 FILLER_38_2011 ();
 sg13g2_decap_8 FILLER_38_2027 ();
 sg13g2_fill_2 FILLER_38_2065 ();
 sg13g2_fill_2 FILLER_38_2085 ();
 sg13g2_decap_8 FILLER_38_2138 ();
 sg13g2_fill_1 FILLER_38_2145 ();
 sg13g2_fill_2 FILLER_38_2150 ();
 sg13g2_fill_1 FILLER_38_2152 ();
 sg13g2_decap_8 FILLER_38_2157 ();
 sg13g2_fill_1 FILLER_38_2164 ();
 sg13g2_decap_8 FILLER_38_2175 ();
 sg13g2_fill_2 FILLER_38_2182 ();
 sg13g2_fill_1 FILLER_38_2184 ();
 sg13g2_fill_1 FILLER_38_2198 ();
 sg13g2_decap_8 FILLER_38_2202 ();
 sg13g2_decap_4 FILLER_38_2209 ();
 sg13g2_fill_1 FILLER_38_2213 ();
 sg13g2_fill_1 FILLER_38_2246 ();
 sg13g2_decap_4 FILLER_38_2260 ();
 sg13g2_fill_1 FILLER_38_2264 ();
 sg13g2_decap_4 FILLER_38_2295 ();
 sg13g2_fill_1 FILLER_38_2315 ();
 sg13g2_fill_1 FILLER_38_2326 ();
 sg13g2_fill_1 FILLER_38_2337 ();
 sg13g2_fill_1 FILLER_38_2356 ();
 sg13g2_fill_1 FILLER_38_2365 ();
 sg13g2_fill_2 FILLER_38_2374 ();
 sg13g2_fill_1 FILLER_38_2376 ();
 sg13g2_fill_1 FILLER_38_2425 ();
 sg13g2_fill_2 FILLER_38_2440 ();
 sg13g2_fill_1 FILLER_38_2454 ();
 sg13g2_fill_2 FILLER_38_2460 ();
 sg13g2_fill_1 FILLER_38_2462 ();
 sg13g2_decap_4 FILLER_38_2475 ();
 sg13g2_decap_4 FILLER_38_2484 ();
 sg13g2_decap_4 FILLER_38_2493 ();
 sg13g2_fill_1 FILLER_38_2497 ();
 sg13g2_fill_2 FILLER_38_2505 ();
 sg13g2_fill_2 FILLER_38_2524 ();
 sg13g2_fill_1 FILLER_38_2548 ();
 sg13g2_fill_1 FILLER_38_2565 ();
 sg13g2_fill_2 FILLER_38_2598 ();
 sg13g2_fill_2 FILLER_38_2617 ();
 sg13g2_fill_1 FILLER_38_2619 ();
 sg13g2_decap_8 FILLER_38_2625 ();
 sg13g2_decap_4 FILLER_38_2632 ();
 sg13g2_decap_4 FILLER_38_2659 ();
 sg13g2_fill_2 FILLER_38_2663 ();
 sg13g2_fill_2 FILLER_38_2682 ();
 sg13g2_fill_1 FILLER_38_2696 ();
 sg13g2_fill_1 FILLER_38_2710 ();
 sg13g2_fill_1 FILLER_38_2805 ();
 sg13g2_fill_2 FILLER_38_2814 ();
 sg13g2_fill_1 FILLER_38_2816 ();
 sg13g2_fill_2 FILLER_38_2891 ();
 sg13g2_fill_1 FILLER_38_2893 ();
 sg13g2_fill_2 FILLER_38_2917 ();
 sg13g2_fill_1 FILLER_38_2919 ();
 sg13g2_fill_2 FILLER_38_3002 ();
 sg13g2_fill_1 FILLER_38_3009 ();
 sg13g2_decap_8 FILLER_38_3038 ();
 sg13g2_fill_2 FILLER_38_3045 ();
 sg13g2_fill_1 FILLER_38_3084 ();
 sg13g2_fill_1 FILLER_38_3113 ();
 sg13g2_fill_1 FILLER_38_3193 ();
 sg13g2_decap_8 FILLER_38_3250 ();
 sg13g2_decap_8 FILLER_38_3257 ();
 sg13g2_decap_4 FILLER_38_3264 ();
 sg13g2_fill_2 FILLER_38_3277 ();
 sg13g2_fill_1 FILLER_38_3279 ();
 sg13g2_fill_2 FILLER_38_3308 ();
 sg13g2_fill_2 FILLER_38_3346 ();
 sg13g2_fill_2 FILLER_38_3376 ();
 sg13g2_fill_1 FILLER_38_3378 ();
 sg13g2_fill_2 FILLER_38_3480 ();
 sg13g2_fill_1 FILLER_38_3482 ();
 sg13g2_fill_2 FILLER_38_3510 ();
 sg13g2_fill_1 FILLER_38_3553 ();
 sg13g2_decap_4 FILLER_38_3576 ();
 sg13g2_decap_4 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_4 ();
 sg13g2_fill_1 FILLER_39_34 ();
 sg13g2_fill_1 FILLER_39_48 ();
 sg13g2_fill_2 FILLER_39_85 ();
 sg13g2_decap_8 FILLER_39_92 ();
 sg13g2_fill_1 FILLER_39_103 ();
 sg13g2_fill_1 FILLER_39_146 ();
 sg13g2_decap_8 FILLER_39_197 ();
 sg13g2_fill_1 FILLER_39_204 ();
 sg13g2_fill_2 FILLER_39_227 ();
 sg13g2_decap_4 FILLER_39_271 ();
 sg13g2_fill_2 FILLER_39_275 ();
 sg13g2_fill_1 FILLER_39_300 ();
 sg13g2_decap_8 FILLER_39_357 ();
 sg13g2_decap_4 FILLER_39_388 ();
 sg13g2_fill_1 FILLER_39_392 ();
 sg13g2_decap_8 FILLER_39_417 ();
 sg13g2_decap_8 FILLER_39_424 ();
 sg13g2_fill_2 FILLER_39_431 ();
 sg13g2_fill_1 FILLER_39_433 ();
 sg13g2_fill_1 FILLER_39_447 ();
 sg13g2_fill_2 FILLER_39_489 ();
 sg13g2_decap_8 FILLER_39_507 ();
 sg13g2_decap_4 FILLER_39_514 ();
 sg13g2_fill_1 FILLER_39_518 ();
 sg13g2_fill_2 FILLER_39_549 ();
 sg13g2_fill_1 FILLER_39_551 ();
 sg13g2_decap_4 FILLER_39_560 ();
 sg13g2_decap_4 FILLER_39_572 ();
 sg13g2_fill_1 FILLER_39_581 ();
 sg13g2_fill_2 FILLER_39_619 ();
 sg13g2_fill_1 FILLER_39_621 ();
 sg13g2_decap_8 FILLER_39_661 ();
 sg13g2_decap_4 FILLER_39_668 ();
 sg13g2_fill_1 FILLER_39_672 ();
 sg13g2_fill_2 FILLER_39_703 ();
 sg13g2_fill_1 FILLER_39_709 ();
 sg13g2_decap_8 FILLER_39_714 ();
 sg13g2_fill_2 FILLER_39_721 ();
 sg13g2_fill_1 FILLER_39_737 ();
 sg13g2_fill_1 FILLER_39_743 ();
 sg13g2_decap_8 FILLER_39_749 ();
 sg13g2_decap_4 FILLER_39_756 ();
 sg13g2_decap_4 FILLER_39_815 ();
 sg13g2_fill_2 FILLER_39_824 ();
 sg13g2_decap_4 FILLER_39_847 ();
 sg13g2_fill_1 FILLER_39_851 ();
 sg13g2_fill_1 FILLER_39_858 ();
 sg13g2_fill_2 FILLER_39_879 ();
 sg13g2_fill_1 FILLER_39_881 ();
 sg13g2_fill_1 FILLER_39_885 ();
 sg13g2_decap_8 FILLER_39_919 ();
 sg13g2_fill_2 FILLER_39_926 ();
 sg13g2_decap_8 FILLER_39_941 ();
 sg13g2_fill_2 FILLER_39_971 ();
 sg13g2_decap_8 FILLER_39_993 ();
 sg13g2_decap_4 FILLER_39_1000 ();
 sg13g2_fill_2 FILLER_39_1010 ();
 sg13g2_decap_8 FILLER_39_1025 ();
 sg13g2_decap_8 FILLER_39_1035 ();
 sg13g2_fill_1 FILLER_39_1042 ();
 sg13g2_decap_4 FILLER_39_1051 ();
 sg13g2_fill_2 FILLER_39_1083 ();
 sg13g2_fill_2 FILLER_39_1098 ();
 sg13g2_fill_2 FILLER_39_1131 ();
 sg13g2_fill_2 FILLER_39_1146 ();
 sg13g2_fill_1 FILLER_39_1148 ();
 sg13g2_fill_2 FILLER_39_1165 ();
 sg13g2_fill_1 FILLER_39_1190 ();
 sg13g2_decap_4 FILLER_39_1227 ();
 sg13g2_fill_2 FILLER_39_1231 ();
 sg13g2_fill_2 FILLER_39_1246 ();
 sg13g2_fill_1 FILLER_39_1248 ();
 sg13g2_fill_2 FILLER_39_1262 ();
 sg13g2_fill_1 FILLER_39_1264 ();
 sg13g2_decap_4 FILLER_39_1278 ();
 sg13g2_decap_8 FILLER_39_1286 ();
 sg13g2_decap_4 FILLER_39_1293 ();
 sg13g2_decap_4 FILLER_39_1301 ();
 sg13g2_fill_2 FILLER_39_1305 ();
 sg13g2_decap_4 FILLER_39_1313 ();
 sg13g2_fill_2 FILLER_39_1334 ();
 sg13g2_decap_8 FILLER_39_1346 ();
 sg13g2_fill_1 FILLER_39_1353 ();
 sg13g2_fill_2 FILLER_39_1387 ();
 sg13g2_fill_2 FILLER_39_1394 ();
 sg13g2_fill_1 FILLER_39_1396 ();
 sg13g2_decap_4 FILLER_39_1433 ();
 sg13g2_fill_1 FILLER_39_1437 ();
 sg13g2_fill_1 FILLER_39_1478 ();
 sg13g2_decap_8 FILLER_39_1483 ();
 sg13g2_fill_1 FILLER_39_1490 ();
 sg13g2_fill_2 FILLER_39_1508 ();
 sg13g2_fill_1 FILLER_39_1510 ();
 sg13g2_fill_1 FILLER_39_1516 ();
 sg13g2_fill_1 FILLER_39_1530 ();
 sg13g2_fill_2 FILLER_39_1556 ();
 sg13g2_decap_8 FILLER_39_1579 ();
 sg13g2_decap_4 FILLER_39_1586 ();
 sg13g2_fill_1 FILLER_39_1590 ();
 sg13g2_decap_8 FILLER_39_1630 ();
 sg13g2_decap_4 FILLER_39_1658 ();
 sg13g2_fill_1 FILLER_39_1662 ();
 sg13g2_fill_1 FILLER_39_1681 ();
 sg13g2_fill_2 FILLER_39_1690 ();
 sg13g2_fill_1 FILLER_39_1692 ();
 sg13g2_decap_8 FILLER_39_1731 ();
 sg13g2_fill_2 FILLER_39_1738 ();
 sg13g2_fill_1 FILLER_39_1740 ();
 sg13g2_fill_2 FILLER_39_1774 ();
 sg13g2_fill_1 FILLER_39_1776 ();
 sg13g2_fill_2 FILLER_39_1799 ();
 sg13g2_fill_2 FILLER_39_1809 ();
 sg13g2_decap_8 FILLER_39_1823 ();
 sg13g2_decap_4 FILLER_39_1830 ();
 sg13g2_fill_2 FILLER_39_1834 ();
 sg13g2_fill_2 FILLER_39_1873 ();
 sg13g2_fill_1 FILLER_39_1875 ();
 sg13g2_decap_8 FILLER_39_1892 ();
 sg13g2_fill_1 FILLER_39_1899 ();
 sg13g2_decap_4 FILLER_39_1932 ();
 sg13g2_fill_1 FILLER_39_1936 ();
 sg13g2_fill_2 FILLER_39_1977 ();
 sg13g2_decap_8 FILLER_39_1992 ();
 sg13g2_fill_1 FILLER_39_1999 ();
 sg13g2_fill_2 FILLER_39_2032 ();
 sg13g2_fill_1 FILLER_39_2034 ();
 sg13g2_fill_2 FILLER_39_2077 ();
 sg13g2_decap_4 FILLER_39_2085 ();
 sg13g2_fill_2 FILLER_39_2093 ();
 sg13g2_fill_1 FILLER_39_2099 ();
 sg13g2_decap_4 FILLER_39_2121 ();
 sg13g2_fill_1 FILLER_39_2148 ();
 sg13g2_decap_4 FILLER_39_2217 ();
 sg13g2_decap_8 FILLER_39_2229 ();
 sg13g2_decap_8 FILLER_39_2236 ();
 sg13g2_fill_2 FILLER_39_2243 ();
 sg13g2_fill_1 FILLER_39_2245 ();
 sg13g2_fill_2 FILLER_39_2251 ();
 sg13g2_decap_4 FILLER_39_2266 ();
 sg13g2_decap_8 FILLER_39_2295 ();
 sg13g2_decap_4 FILLER_39_2307 ();
 sg13g2_fill_2 FILLER_39_2311 ();
 sg13g2_fill_1 FILLER_39_2336 ();
 sg13g2_decap_8 FILLER_39_2352 ();
 sg13g2_fill_2 FILLER_39_2372 ();
 sg13g2_fill_2 FILLER_39_2403 ();
 sg13g2_fill_1 FILLER_39_2429 ();
 sg13g2_fill_1 FILLER_39_2443 ();
 sg13g2_fill_1 FILLER_39_2453 ();
 sg13g2_fill_2 FILLER_39_2459 ();
 sg13g2_decap_4 FILLER_39_2480 ();
 sg13g2_fill_2 FILLER_39_2484 ();
 sg13g2_fill_2 FILLER_39_2505 ();
 sg13g2_fill_1 FILLER_39_2507 ();
 sg13g2_decap_8 FILLER_39_2523 ();
 sg13g2_decap_4 FILLER_39_2548 ();
 sg13g2_fill_1 FILLER_39_2552 ();
 sg13g2_fill_2 FILLER_39_2557 ();
 sg13g2_fill_1 FILLER_39_2573 ();
 sg13g2_decap_4 FILLER_39_2587 ();
 sg13g2_fill_1 FILLER_39_2608 ();
 sg13g2_decap_8 FILLER_39_2617 ();
 sg13g2_decap_4 FILLER_39_2624 ();
 sg13g2_fill_2 FILLER_39_2628 ();
 sg13g2_decap_8 FILLER_39_2657 ();
 sg13g2_fill_2 FILLER_39_2664 ();
 sg13g2_fill_2 FILLER_39_2717 ();
 sg13g2_fill_1 FILLER_39_2755 ();
 sg13g2_fill_2 FILLER_39_2800 ();
 sg13g2_fill_2 FILLER_39_2819 ();
 sg13g2_fill_1 FILLER_39_2821 ();
 sg13g2_fill_2 FILLER_39_2856 ();
 sg13g2_fill_1 FILLER_39_2858 ();
 sg13g2_fill_1 FILLER_39_2885 ();
 sg13g2_fill_2 FILLER_39_2956 ();
 sg13g2_fill_1 FILLER_39_2958 ();
 sg13g2_fill_1 FILLER_39_2982 ();
 sg13g2_fill_1 FILLER_39_3015 ();
 sg13g2_fill_1 FILLER_39_3043 ();
 sg13g2_decap_8 FILLER_39_3070 ();
 sg13g2_decap_4 FILLER_39_3077 ();
 sg13g2_decap_8 FILLER_39_3086 ();
 sg13g2_fill_2 FILLER_39_3093 ();
 sg13g2_decap_4 FILLER_39_3099 ();
 sg13g2_fill_2 FILLER_39_3103 ();
 sg13g2_fill_2 FILLER_39_3195 ();
 sg13g2_fill_2 FILLER_39_3223 ();
 sg13g2_fill_2 FILLER_39_3244 ();
 sg13g2_decap_8 FILLER_39_3255 ();
 sg13g2_fill_1 FILLER_39_3262 ();
 sg13g2_fill_2 FILLER_39_3287 ();
 sg13g2_fill_2 FILLER_39_3293 ();
 sg13g2_fill_2 FILLER_39_3300 ();
 sg13g2_fill_2 FILLER_39_3307 ();
 sg13g2_fill_1 FILLER_39_3309 ();
 sg13g2_decap_4 FILLER_39_3378 ();
 sg13g2_decap_4 FILLER_39_3395 ();
 sg13g2_decap_8 FILLER_39_3420 ();
 sg13g2_fill_1 FILLER_39_3427 ();
 sg13g2_decap_8 FILLER_39_3445 ();
 sg13g2_fill_2 FILLER_39_3457 ();
 sg13g2_fill_1 FILLER_39_3459 ();
 sg13g2_fill_1 FILLER_39_3464 ();
 sg13g2_decap_8 FILLER_39_3474 ();
 sg13g2_fill_2 FILLER_39_3481 ();
 sg13g2_decap_4 FILLER_39_3487 ();
 sg13g2_fill_1 FILLER_39_3491 ();
 sg13g2_fill_1 FILLER_39_3542 ();
 sg13g2_fill_1 FILLER_39_3547 ();
 sg13g2_decap_4 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_36 ();
 sg13g2_fill_1 FILLER_40_55 ();
 sg13g2_fill_1 FILLER_40_98 ();
 sg13g2_decap_4 FILLER_40_115 ();
 sg13g2_fill_1 FILLER_40_170 ();
 sg13g2_fill_2 FILLER_40_180 ();
 sg13g2_fill_2 FILLER_40_196 ();
 sg13g2_fill_1 FILLER_40_198 ();
 sg13g2_fill_2 FILLER_40_204 ();
 sg13g2_fill_2 FILLER_40_220 ();
 sg13g2_fill_2 FILLER_40_261 ();
 sg13g2_fill_1 FILLER_40_303 ();
 sg13g2_fill_1 FILLER_40_317 ();
 sg13g2_fill_1 FILLER_40_340 ();
 sg13g2_fill_2 FILLER_40_381 ();
 sg13g2_fill_1 FILLER_40_383 ();
 sg13g2_fill_2 FILLER_40_399 ();
 sg13g2_decap_8 FILLER_40_417 ();
 sg13g2_decap_4 FILLER_40_424 ();
 sg13g2_fill_1 FILLER_40_428 ();
 sg13g2_fill_2 FILLER_40_433 ();
 sg13g2_fill_1 FILLER_40_452 ();
 sg13g2_fill_2 FILLER_40_517 ();
 sg13g2_fill_1 FILLER_40_519 ();
 sg13g2_decap_4 FILLER_40_524 ();
 sg13g2_fill_1 FILLER_40_528 ();
 sg13g2_fill_2 FILLER_40_534 ();
 sg13g2_fill_2 FILLER_40_541 ();
 sg13g2_decap_8 FILLER_40_547 ();
 sg13g2_decap_4 FILLER_40_554 ();
 sg13g2_fill_2 FILLER_40_558 ();
 sg13g2_fill_1 FILLER_40_565 ();
 sg13g2_fill_1 FILLER_40_589 ();
 sg13g2_fill_2 FILLER_40_613 ();
 sg13g2_fill_1 FILLER_40_615 ();
 sg13g2_fill_1 FILLER_40_640 ();
 sg13g2_fill_2 FILLER_40_651 ();
 sg13g2_decap_8 FILLER_40_662 ();
 sg13g2_fill_2 FILLER_40_669 ();
 sg13g2_fill_2 FILLER_40_676 ();
 sg13g2_fill_1 FILLER_40_694 ();
 sg13g2_fill_1 FILLER_40_713 ();
 sg13g2_fill_2 FILLER_40_727 ();
 sg13g2_fill_1 FILLER_40_750 ();
 sg13g2_fill_2 FILLER_40_764 ();
 sg13g2_fill_1 FILLER_40_766 ();
 sg13g2_fill_2 FILLER_40_783 ();
 sg13g2_fill_1 FILLER_40_785 ();
 sg13g2_fill_2 FILLER_40_790 ();
 sg13g2_fill_1 FILLER_40_792 ();
 sg13g2_decap_4 FILLER_40_797 ();
 sg13g2_decap_4 FILLER_40_820 ();
 sg13g2_decap_8 FILLER_40_831 ();
 sg13g2_decap_8 FILLER_40_854 ();
 sg13g2_decap_8 FILLER_40_861 ();
 sg13g2_fill_2 FILLER_40_868 ();
 sg13g2_fill_1 FILLER_40_870 ();
 sg13g2_fill_2 FILLER_40_874 ();
 sg13g2_decap_8 FILLER_40_892 ();
 sg13g2_fill_2 FILLER_40_899 ();
 sg13g2_decap_8 FILLER_40_909 ();
 sg13g2_decap_4 FILLER_40_916 ();
 sg13g2_fill_1 FILLER_40_920 ();
 sg13g2_decap_4 FILLER_40_924 ();
 sg13g2_decap_8 FILLER_40_979 ();
 sg13g2_fill_2 FILLER_40_998 ();
 sg13g2_fill_1 FILLER_40_1000 ();
 sg13g2_decap_4 FILLER_40_1009 ();
 sg13g2_fill_1 FILLER_40_1021 ();
 sg13g2_fill_1 FILLER_40_1028 ();
 sg13g2_decap_8 FILLER_40_1037 ();
 sg13g2_fill_1 FILLER_40_1044 ();
 sg13g2_fill_2 FILLER_40_1058 ();
 sg13g2_fill_1 FILLER_40_1064 ();
 sg13g2_decap_8 FILLER_40_1078 ();
 sg13g2_fill_2 FILLER_40_1118 ();
 sg13g2_fill_1 FILLER_40_1120 ();
 sg13g2_fill_2 FILLER_40_1139 ();
 sg13g2_fill_2 FILLER_40_1161 ();
 sg13g2_fill_1 FILLER_40_1163 ();
 sg13g2_fill_1 FILLER_40_1169 ();
 sg13g2_fill_2 FILLER_40_1190 ();
 sg13g2_fill_1 FILLER_40_1192 ();
 sg13g2_fill_1 FILLER_40_1249 ();
 sg13g2_decap_4 FILLER_40_1269 ();
 sg13g2_fill_1 FILLER_40_1273 ();
 sg13g2_decap_4 FILLER_40_1288 ();
 sg13g2_fill_2 FILLER_40_1323 ();
 sg13g2_fill_1 FILLER_40_1325 ();
 sg13g2_fill_2 FILLER_40_1335 ();
 sg13g2_decap_8 FILLER_40_1369 ();
 sg13g2_decap_4 FILLER_40_1376 ();
 sg13g2_fill_2 FILLER_40_1380 ();
 sg13g2_fill_2 FILLER_40_1399 ();
 sg13g2_fill_2 FILLER_40_1419 ();
 sg13g2_fill_2 FILLER_40_1430 ();
 sg13g2_fill_1 FILLER_40_1432 ();
 sg13g2_fill_2 FILLER_40_1475 ();
 sg13g2_decap_4 FILLER_40_1503 ();
 sg13g2_decap_8 FILLER_40_1557 ();
 sg13g2_fill_1 FILLER_40_1583 ();
 sg13g2_fill_2 FILLER_40_1601 ();
 sg13g2_decap_8 FILLER_40_1622 ();
 sg13g2_fill_2 FILLER_40_1629 ();
 sg13g2_decap_4 FILLER_40_1644 ();
 sg13g2_fill_2 FILLER_40_1648 ();
 sg13g2_decap_4 FILLER_40_1663 ();
 sg13g2_fill_2 FILLER_40_1680 ();
 sg13g2_fill_1 FILLER_40_1698 ();
 sg13g2_decap_8 FILLER_40_1736 ();
 sg13g2_fill_2 FILLER_40_1747 ();
 sg13g2_decap_8 FILLER_40_1758 ();
 sg13g2_fill_1 FILLER_40_1765 ();
 sg13g2_fill_2 FILLER_40_1794 ();
 sg13g2_fill_1 FILLER_40_1800 ();
 sg13g2_decap_4 FILLER_40_1817 ();
 sg13g2_decap_4 FILLER_40_1826 ();
 sg13g2_decap_8 FILLER_40_1843 ();
 sg13g2_fill_2 FILLER_40_1850 ();
 sg13g2_decap_8 FILLER_40_1864 ();
 sg13g2_fill_2 FILLER_40_1871 ();
 sg13g2_fill_1 FILLER_40_1873 ();
 sg13g2_fill_2 FILLER_40_1887 ();
 sg13g2_decap_4 FILLER_40_1909 ();
 sg13g2_fill_1 FILLER_40_1913 ();
 sg13g2_decap_4 FILLER_40_1936 ();
 sg13g2_fill_1 FILLER_40_1940 ();
 sg13g2_fill_1 FILLER_40_1949 ();
 sg13g2_fill_2 FILLER_40_2000 ();
 sg13g2_fill_1 FILLER_40_2002 ();
 sg13g2_fill_2 FILLER_40_2012 ();
 sg13g2_fill_1 FILLER_40_2014 ();
 sg13g2_fill_2 FILLER_40_2052 ();
 sg13g2_fill_1 FILLER_40_2054 ();
 sg13g2_decap_4 FILLER_40_2090 ();
 sg13g2_fill_2 FILLER_40_2099 ();
 sg13g2_decap_8 FILLER_40_2119 ();
 sg13g2_fill_1 FILLER_40_2126 ();
 sg13g2_fill_2 FILLER_40_2142 ();
 sg13g2_fill_1 FILLER_40_2144 ();
 sg13g2_decap_4 FILLER_40_2161 ();
 sg13g2_fill_1 FILLER_40_2165 ();
 sg13g2_fill_1 FILLER_40_2170 ();
 sg13g2_decap_4 FILLER_40_2183 ();
 sg13g2_fill_2 FILLER_40_2207 ();
 sg13g2_fill_1 FILLER_40_2209 ();
 sg13g2_fill_2 FILLER_40_2220 ();
 sg13g2_decap_8 FILLER_40_2255 ();
 sg13g2_fill_1 FILLER_40_2262 ();
 sg13g2_fill_1 FILLER_40_2276 ();
 sg13g2_decap_8 FILLER_40_2292 ();
 sg13g2_decap_4 FILLER_40_2299 ();
 sg13g2_fill_1 FILLER_40_2303 ();
 sg13g2_fill_1 FILLER_40_2317 ();
 sg13g2_decap_4 FILLER_40_2332 ();
 sg13g2_decap_8 FILLER_40_2351 ();
 sg13g2_fill_2 FILLER_40_2358 ();
 sg13g2_fill_1 FILLER_40_2360 ();
 sg13g2_decap_4 FILLER_40_2371 ();
 sg13g2_fill_2 FILLER_40_2384 ();
 sg13g2_fill_1 FILLER_40_2386 ();
 sg13g2_decap_8 FILLER_40_2399 ();
 sg13g2_fill_2 FILLER_40_2406 ();
 sg13g2_fill_1 FILLER_40_2408 ();
 sg13g2_fill_2 FILLER_40_2443 ();
 sg13g2_decap_8 FILLER_40_2476 ();
 sg13g2_fill_2 FILLER_40_2483 ();
 sg13g2_fill_1 FILLER_40_2485 ();
 sg13g2_fill_2 FILLER_40_2500 ();
 sg13g2_fill_1 FILLER_40_2502 ();
 sg13g2_decap_4 FILLER_40_2509 ();
 sg13g2_decap_4 FILLER_40_2518 ();
 sg13g2_fill_1 FILLER_40_2522 ();
 sg13g2_fill_1 FILLER_40_2529 ();
 sg13g2_decap_8 FILLER_40_2543 ();
 sg13g2_fill_2 FILLER_40_2550 ();
 sg13g2_fill_1 FILLER_40_2564 ();
 sg13g2_decap_8 FILLER_40_2593 ();
 sg13g2_fill_2 FILLER_40_2600 ();
 sg13g2_fill_1 FILLER_40_2602 ();
 sg13g2_decap_4 FILLER_40_2617 ();
 sg13g2_decap_4 FILLER_40_2693 ();
 sg13g2_fill_2 FILLER_40_2733 ();
 sg13g2_fill_2 FILLER_40_2750 ();
 sg13g2_fill_1 FILLER_40_2752 ();
 sg13g2_fill_1 FILLER_40_2848 ();
 sg13g2_fill_1 FILLER_40_2889 ();
 sg13g2_decap_4 FILLER_40_2916 ();
 sg13g2_fill_2 FILLER_40_2920 ();
 sg13g2_fill_1 FILLER_40_2971 ();
 sg13g2_fill_1 FILLER_40_2977 ();
 sg13g2_fill_2 FILLER_40_3028 ();
 sg13g2_fill_1 FILLER_40_3030 ();
 sg13g2_fill_2 FILLER_40_3047 ();
 sg13g2_fill_1 FILLER_40_3049 ();
 sg13g2_fill_1 FILLER_40_3058 ();
 sg13g2_fill_1 FILLER_40_3072 ();
 sg13g2_fill_1 FILLER_40_3086 ();
 sg13g2_decap_8 FILLER_40_3109 ();
 sg13g2_decap_8 FILLER_40_3116 ();
 sg13g2_fill_2 FILLER_40_3123 ();
 sg13g2_decap_8 FILLER_40_3138 ();
 sg13g2_fill_1 FILLER_40_3145 ();
 sg13g2_fill_1 FILLER_40_3169 ();
 sg13g2_fill_2 FILLER_40_3186 ();
 sg13g2_fill_1 FILLER_40_3209 ();
 sg13g2_fill_1 FILLER_40_3216 ();
 sg13g2_fill_2 FILLER_40_3222 ();
 sg13g2_fill_2 FILLER_40_3309 ();
 sg13g2_fill_2 FILLER_40_3319 ();
 sg13g2_decap_8 FILLER_40_3350 ();
 sg13g2_fill_2 FILLER_40_3357 ();
 sg13g2_fill_2 FILLER_40_3368 ();
 sg13g2_decap_4 FILLER_40_3428 ();
 sg13g2_fill_1 FILLER_40_3454 ();
 sg13g2_fill_2 FILLER_40_3561 ();
 sg13g2_fill_1 FILLER_40_3563 ();
 sg13g2_decap_8 FILLER_40_3573 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_7 ();
 sg13g2_fill_1 FILLER_41_39 ();
 sg13g2_fill_1 FILLER_41_62 ();
 sg13g2_fill_2 FILLER_41_71 ();
 sg13g2_fill_1 FILLER_41_82 ();
 sg13g2_decap_8 FILLER_41_93 ();
 sg13g2_decap_4 FILLER_41_100 ();
 sg13g2_fill_1 FILLER_41_104 ();
 sg13g2_fill_1 FILLER_41_109 ();
 sg13g2_decap_4 FILLER_41_120 ();
 sg13g2_fill_2 FILLER_41_124 ();
 sg13g2_fill_1 FILLER_41_154 ();
 sg13g2_fill_2 FILLER_41_177 ();
 sg13g2_fill_1 FILLER_41_221 ();
 sg13g2_fill_2 FILLER_41_241 ();
 sg13g2_fill_2 FILLER_41_248 ();
 sg13g2_fill_1 FILLER_41_250 ();
 sg13g2_decap_8 FILLER_41_257 ();
 sg13g2_fill_2 FILLER_41_277 ();
 sg13g2_fill_2 FILLER_41_371 ();
 sg13g2_fill_1 FILLER_41_373 ();
 sg13g2_decap_8 FILLER_41_388 ();
 sg13g2_fill_2 FILLER_41_395 ();
 sg13g2_fill_1 FILLER_41_397 ();
 sg13g2_fill_2 FILLER_41_416 ();
 sg13g2_fill_1 FILLER_41_418 ();
 sg13g2_fill_1 FILLER_41_438 ();
 sg13g2_decap_4 FILLER_41_449 ();
 sg13g2_fill_2 FILLER_41_472 ();
 sg13g2_fill_1 FILLER_41_496 ();
 sg13g2_fill_2 FILLER_41_525 ();
 sg13g2_fill_1 FILLER_41_527 ();
 sg13g2_fill_1 FILLER_41_545 ();
 sg13g2_decap_4 FILLER_41_551 ();
 sg13g2_fill_2 FILLER_41_555 ();
 sg13g2_decap_4 FILLER_41_573 ();
 sg13g2_fill_1 FILLER_41_577 ();
 sg13g2_fill_1 FILLER_41_583 ();
 sg13g2_fill_1 FILLER_41_602 ();
 sg13g2_fill_2 FILLER_41_647 ();
 sg13g2_fill_1 FILLER_41_649 ();
 sg13g2_decap_4 FILLER_41_684 ();
 sg13g2_fill_2 FILLER_41_688 ();
 sg13g2_fill_1 FILLER_41_704 ();
 sg13g2_decap_4 FILLER_41_718 ();
 sg13g2_fill_1 FILLER_41_733 ();
 sg13g2_fill_1 FILLER_41_739 ();
 sg13g2_decap_8 FILLER_41_749 ();
 sg13g2_decap_8 FILLER_41_756 ();
 sg13g2_fill_1 FILLER_41_773 ();
 sg13g2_fill_1 FILLER_41_821 ();
 sg13g2_fill_1 FILLER_41_827 ();
 sg13g2_fill_2 FILLER_41_858 ();
 sg13g2_fill_1 FILLER_41_860 ();
 sg13g2_decap_4 FILLER_41_869 ();
 sg13g2_fill_2 FILLER_41_873 ();
 sg13g2_fill_2 FILLER_41_893 ();
 sg13g2_fill_1 FILLER_41_895 ();
 sg13g2_fill_2 FILLER_41_909 ();
 sg13g2_fill_1 FILLER_41_911 ();
 sg13g2_fill_2 FILLER_41_941 ();
 sg13g2_fill_1 FILLER_41_943 ();
 sg13g2_fill_2 FILLER_41_960 ();
 sg13g2_fill_2 FILLER_41_987 ();
 sg13g2_decap_8 FILLER_41_1006 ();
 sg13g2_fill_2 FILLER_41_1013 ();
 sg13g2_fill_1 FILLER_41_1015 ();
 sg13g2_fill_2 FILLER_41_1028 ();
 sg13g2_fill_2 FILLER_41_1053 ();
 sg13g2_fill_1 FILLER_41_1062 ();
 sg13g2_fill_2 FILLER_41_1076 ();
 sg13g2_fill_1 FILLER_41_1078 ();
 sg13g2_decap_8 FILLER_41_1104 ();
 sg13g2_fill_1 FILLER_41_1111 ();
 sg13g2_fill_1 FILLER_41_1128 ();
 sg13g2_fill_2 FILLER_41_1142 ();
 sg13g2_fill_1 FILLER_41_1144 ();
 sg13g2_fill_2 FILLER_41_1162 ();
 sg13g2_decap_8 FILLER_41_1176 ();
 sg13g2_decap_8 FILLER_41_1213 ();
 sg13g2_decap_8 FILLER_41_1225 ();
 sg13g2_decap_4 FILLER_41_1232 ();
 sg13g2_fill_2 FILLER_41_1236 ();
 sg13g2_fill_1 FILLER_41_1266 ();
 sg13g2_decap_8 FILLER_41_1291 ();
 sg13g2_decap_4 FILLER_41_1298 ();
 sg13g2_fill_1 FILLER_41_1302 ();
 sg13g2_fill_1 FILLER_41_1308 ();
 sg13g2_decap_4 FILLER_41_1314 ();
 sg13g2_fill_1 FILLER_41_1318 ();
 sg13g2_fill_2 FILLER_41_1333 ();
 sg13g2_fill_1 FILLER_41_1335 ();
 sg13g2_decap_8 FILLER_41_1344 ();
 sg13g2_decap_8 FILLER_41_1351 ();
 sg13g2_fill_2 FILLER_41_1358 ();
 sg13g2_fill_1 FILLER_41_1360 ();
 sg13g2_fill_2 FILLER_41_1367 ();
 sg13g2_fill_1 FILLER_41_1369 ();
 sg13g2_fill_1 FILLER_41_1386 ();
 sg13g2_fill_1 FILLER_41_1396 ();
 sg13g2_fill_2 FILLER_41_1409 ();
 sg13g2_fill_1 FILLER_41_1411 ();
 sg13g2_fill_1 FILLER_41_1463 ();
 sg13g2_fill_2 FILLER_41_1480 ();
 sg13g2_fill_1 FILLER_41_1482 ();
 sg13g2_decap_4 FILLER_41_1495 ();
 sg13g2_fill_2 FILLER_41_1499 ();
 sg13g2_fill_1 FILLER_41_1518 ();
 sg13g2_decap_4 FILLER_41_1567 ();
 sg13g2_fill_2 FILLER_41_1571 ();
 sg13g2_fill_2 FILLER_41_1581 ();
 sg13g2_decap_8 FILLER_41_1593 ();
 sg13g2_fill_1 FILLER_41_1600 ();
 sg13g2_decap_8 FILLER_41_1609 ();
 sg13g2_fill_1 FILLER_41_1616 ();
 sg13g2_fill_2 FILLER_41_1632 ();
 sg13g2_fill_2 FILLER_41_1642 ();
 sg13g2_decap_4 FILLER_41_1648 ();
 sg13g2_fill_1 FILLER_41_1652 ();
 sg13g2_fill_1 FILLER_41_1679 ();
 sg13g2_decap_8 FILLER_41_1705 ();
 sg13g2_fill_1 FILLER_41_1712 ();
 sg13g2_fill_2 FILLER_41_1721 ();
 sg13g2_decap_4 FILLER_41_1744 ();
 sg13g2_fill_2 FILLER_41_1748 ();
 sg13g2_fill_2 FILLER_41_1760 ();
 sg13g2_fill_2 FILLER_41_1779 ();
 sg13g2_fill_1 FILLER_41_1830 ();
 sg13g2_fill_2 FILLER_41_1853 ();
 sg13g2_fill_1 FILLER_41_1869 ();
 sg13g2_decap_4 FILLER_41_1893 ();
 sg13g2_fill_2 FILLER_41_1897 ();
 sg13g2_decap_4 FILLER_41_1911 ();
 sg13g2_decap_8 FILLER_41_1925 ();
 sg13g2_fill_1 FILLER_41_1932 ();
 sg13g2_fill_2 FILLER_41_1946 ();
 sg13g2_decap_8 FILLER_41_1966 ();
 sg13g2_decap_8 FILLER_41_1973 ();
 sg13g2_decap_4 FILLER_41_1993 ();
 sg13g2_fill_2 FILLER_41_1997 ();
 sg13g2_fill_2 FILLER_41_2026 ();
 sg13g2_fill_1 FILLER_41_2028 ();
 sg13g2_fill_1 FILLER_41_2052 ();
 sg13g2_decap_8 FILLER_41_2081 ();
 sg13g2_decap_8 FILLER_41_2105 ();
 sg13g2_fill_2 FILLER_41_2112 ();
 sg13g2_fill_1 FILLER_41_2114 ();
 sg13g2_decap_8 FILLER_41_2126 ();
 sg13g2_fill_1 FILLER_41_2133 ();
 sg13g2_decap_8 FILLER_41_2138 ();
 sg13g2_decap_8 FILLER_41_2145 ();
 sg13g2_decap_8 FILLER_41_2152 ();
 sg13g2_fill_1 FILLER_41_2170 ();
 sg13g2_decap_8 FILLER_41_2175 ();
 sg13g2_decap_8 FILLER_41_2182 ();
 sg13g2_decap_8 FILLER_41_2189 ();
 sg13g2_fill_2 FILLER_41_2196 ();
 sg13g2_fill_1 FILLER_41_2198 ();
 sg13g2_fill_2 FILLER_41_2204 ();
 sg13g2_decap_8 FILLER_41_2210 ();
 sg13g2_decap_4 FILLER_41_2217 ();
 sg13g2_decap_4 FILLER_41_2231 ();
 sg13g2_fill_1 FILLER_41_2235 ();
 sg13g2_decap_4 FILLER_41_2240 ();
 sg13g2_fill_1 FILLER_41_2260 ();
 sg13g2_decap_8 FILLER_41_2265 ();
 sg13g2_fill_1 FILLER_41_2272 ();
 sg13g2_fill_2 FILLER_41_2286 ();
 sg13g2_fill_2 FILLER_41_2301 ();
 sg13g2_fill_2 FILLER_41_2334 ();
 sg13g2_decap_8 FILLER_41_2352 ();
 sg13g2_decap_4 FILLER_41_2359 ();
 sg13g2_fill_2 FILLER_41_2363 ();
 sg13g2_fill_1 FILLER_41_2370 ();
 sg13g2_decap_4 FILLER_41_2395 ();
 sg13g2_fill_2 FILLER_41_2399 ();
 sg13g2_fill_1 FILLER_41_2427 ();
 sg13g2_decap_4 FILLER_41_2433 ();
 sg13g2_fill_1 FILLER_41_2437 ();
 sg13g2_fill_2 FILLER_41_2446 ();
 sg13g2_fill_1 FILLER_41_2448 ();
 sg13g2_fill_1 FILLER_41_2454 ();
 sg13g2_decap_8 FILLER_41_2463 ();
 sg13g2_decap_4 FILLER_41_2470 ();
 sg13g2_fill_1 FILLER_41_2474 ();
 sg13g2_decap_8 FILLER_41_2521 ();
 sg13g2_fill_1 FILLER_41_2528 ();
 sg13g2_fill_2 FILLER_41_2553 ();
 sg13g2_fill_1 FILLER_41_2555 ();
 sg13g2_fill_1 FILLER_41_2566 ();
 sg13g2_decap_8 FILLER_41_2600 ();
 sg13g2_fill_2 FILLER_41_2607 ();
 sg13g2_fill_2 FILLER_41_2646 ();
 sg13g2_decap_8 FILLER_41_2678 ();
 sg13g2_fill_2 FILLER_41_2685 ();
 sg13g2_fill_1 FILLER_41_2715 ();
 sg13g2_fill_2 FILLER_41_2742 ();
 sg13g2_fill_1 FILLER_41_2744 ();
 sg13g2_fill_1 FILLER_41_2766 ();
 sg13g2_fill_1 FILLER_41_2776 ();
 sg13g2_fill_2 FILLER_41_2790 ();
 sg13g2_fill_1 FILLER_41_2820 ();
 sg13g2_fill_1 FILLER_41_2853 ();
 sg13g2_fill_1 FILLER_41_2859 ();
 sg13g2_fill_1 FILLER_41_2877 ();
 sg13g2_fill_2 FILLER_41_2964 ();
 sg13g2_fill_2 FILLER_41_3020 ();
 sg13g2_fill_2 FILLER_41_3035 ();
 sg13g2_fill_2 FILLER_41_3064 ();
 sg13g2_decap_8 FILLER_41_3075 ();
 sg13g2_decap_8 FILLER_41_3107 ();
 sg13g2_fill_2 FILLER_41_3114 ();
 sg13g2_decap_4 FILLER_41_3137 ();
 sg13g2_fill_2 FILLER_41_3141 ();
 sg13g2_fill_1 FILLER_41_3151 ();
 sg13g2_decap_8 FILLER_41_3165 ();
 sg13g2_fill_2 FILLER_41_3172 ();
 sg13g2_fill_1 FILLER_41_3212 ();
 sg13g2_fill_2 FILLER_41_3238 ();
 sg13g2_fill_2 FILLER_41_3245 ();
 sg13g2_decap_4 FILLER_41_3256 ();
 sg13g2_decap_4 FILLER_41_3264 ();
 sg13g2_decap_8 FILLER_41_3276 ();
 sg13g2_fill_2 FILLER_41_3283 ();
 sg13g2_fill_2 FILLER_41_3298 ();
 sg13g2_fill_1 FILLER_41_3300 ();
 sg13g2_fill_2 FILLER_41_3322 ();
 sg13g2_fill_1 FILLER_41_3324 ();
 sg13g2_fill_2 FILLER_41_3329 ();
 sg13g2_fill_2 FILLER_41_3339 ();
 sg13g2_fill_1 FILLER_41_3341 ();
 sg13g2_fill_2 FILLER_41_3370 ();
 sg13g2_fill_2 FILLER_41_3393 ();
 sg13g2_fill_2 FILLER_41_3417 ();
 sg13g2_decap_4 FILLER_41_3427 ();
 sg13g2_fill_2 FILLER_41_3468 ();
 sg13g2_fill_1 FILLER_41_3470 ();
 sg13g2_fill_2 FILLER_41_3493 ();
 sg13g2_fill_1 FILLER_41_3495 ();
 sg13g2_fill_1 FILLER_41_3505 ();
 sg13g2_fill_1 FILLER_41_3534 ();
 sg13g2_decap_4 FILLER_41_3544 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_39 ();
 sg13g2_fill_1 FILLER_42_62 ();
 sg13g2_decap_4 FILLER_42_86 ();
 sg13g2_fill_2 FILLER_42_114 ();
 sg13g2_fill_2 FILLER_42_256 ();
 sg13g2_fill_1 FILLER_42_258 ();
 sg13g2_fill_2 FILLER_42_302 ();
 sg13g2_fill_1 FILLER_42_304 ();
 sg13g2_fill_2 FILLER_42_318 ();
 sg13g2_fill_2 FILLER_42_329 ();
 sg13g2_decap_8 FILLER_42_384 ();
 sg13g2_fill_1 FILLER_42_391 ();
 sg13g2_fill_2 FILLER_42_423 ();
 sg13g2_decap_8 FILLER_42_452 ();
 sg13g2_decap_4 FILLER_42_459 ();
 sg13g2_fill_1 FILLER_42_463 ();
 sg13g2_decap_4 FILLER_42_478 ();
 sg13g2_fill_1 FILLER_42_508 ();
 sg13g2_fill_2 FILLER_42_518 ();
 sg13g2_fill_1 FILLER_42_520 ();
 sg13g2_fill_2 FILLER_42_525 ();
 sg13g2_fill_1 FILLER_42_535 ();
 sg13g2_fill_2 FILLER_42_541 ();
 sg13g2_decap_8 FILLER_42_546 ();
 sg13g2_fill_2 FILLER_42_553 ();
 sg13g2_fill_2 FILLER_42_571 ();
 sg13g2_fill_2 FILLER_42_594 ();
 sg13g2_fill_1 FILLER_42_596 ();
 sg13g2_fill_2 FILLER_42_614 ();
 sg13g2_fill_1 FILLER_42_616 ();
 sg13g2_fill_2 FILLER_42_625 ();
 sg13g2_fill_1 FILLER_42_627 ();
 sg13g2_decap_4 FILLER_42_655 ();
 sg13g2_fill_2 FILLER_42_659 ();
 sg13g2_decap_4 FILLER_42_679 ();
 sg13g2_fill_1 FILLER_42_688 ();
 sg13g2_decap_8 FILLER_42_694 ();
 sg13g2_fill_1 FILLER_42_705 ();
 sg13g2_fill_2 FILLER_42_729 ();
 sg13g2_fill_2 FILLER_42_777 ();
 sg13g2_fill_1 FILLER_42_779 ();
 sg13g2_fill_2 FILLER_42_796 ();
 sg13g2_fill_1 FILLER_42_810 ();
 sg13g2_fill_2 FILLER_42_827 ();
 sg13g2_fill_2 FILLER_42_835 ();
 sg13g2_fill_1 FILLER_42_837 ();
 sg13g2_fill_2 FILLER_42_855 ();
 sg13g2_fill_1 FILLER_42_857 ();
 sg13g2_fill_1 FILLER_42_907 ();
 sg13g2_decap_8 FILLER_42_921 ();
 sg13g2_fill_2 FILLER_42_928 ();
 sg13g2_decap_4 FILLER_42_935 ();
 sg13g2_fill_1 FILLER_42_939 ();
 sg13g2_decap_4 FILLER_42_1011 ();
 sg13g2_fill_1 FILLER_42_1051 ();
 sg13g2_decap_4 FILLER_42_1098 ();
 sg13g2_decap_4 FILLER_42_1147 ();
 sg13g2_fill_1 FILLER_42_1151 ();
 sg13g2_fill_1 FILLER_42_1156 ();
 sg13g2_decap_8 FILLER_42_1167 ();
 sg13g2_decap_4 FILLER_42_1174 ();
 sg13g2_fill_1 FILLER_42_1178 ();
 sg13g2_decap_4 FILLER_42_1215 ();
 sg13g2_fill_1 FILLER_42_1248 ();
 sg13g2_fill_2 FILLER_42_1254 ();
 sg13g2_fill_1 FILLER_42_1256 ();
 sg13g2_fill_2 FILLER_42_1263 ();
 sg13g2_fill_1 FILLER_42_1265 ();
 sg13g2_fill_2 FILLER_42_1274 ();
 sg13g2_fill_1 FILLER_42_1279 ();
 sg13g2_fill_2 FILLER_42_1290 ();
 sg13g2_decap_4 FILLER_42_1296 ();
 sg13g2_fill_2 FILLER_42_1339 ();
 sg13g2_decap_4 FILLER_42_1372 ();
 sg13g2_fill_1 FILLER_42_1376 ();
 sg13g2_fill_2 FILLER_42_1382 ();
 sg13g2_fill_2 FILLER_42_1399 ();
 sg13g2_fill_1 FILLER_42_1416 ();
 sg13g2_decap_4 FILLER_42_1458 ();
 sg13g2_fill_2 FILLER_42_1462 ();
 sg13g2_decap_8 FILLER_42_1480 ();
 sg13g2_decap_4 FILLER_42_1487 ();
 sg13g2_fill_2 FILLER_42_1532 ();
 sg13g2_fill_1 FILLER_42_1534 ();
 sg13g2_fill_2 FILLER_42_1552 ();
 sg13g2_fill_1 FILLER_42_1554 ();
 sg13g2_decap_4 FILLER_42_1565 ();
 sg13g2_fill_2 FILLER_42_1601 ();
 sg13g2_fill_1 FILLER_42_1603 ();
 sg13g2_decap_8 FILLER_42_1628 ();
 sg13g2_fill_2 FILLER_42_1635 ();
 sg13g2_decap_4 FILLER_42_1660 ();
 sg13g2_fill_1 FILLER_42_1664 ();
 sg13g2_fill_1 FILLER_42_1701 ();
 sg13g2_fill_1 FILLER_42_1706 ();
 sg13g2_fill_2 FILLER_42_1717 ();
 sg13g2_fill_2 FILLER_42_1732 ();
 sg13g2_fill_2 FILLER_42_1760 ();
 sg13g2_fill_1 FILLER_42_1762 ();
 sg13g2_decap_4 FILLER_42_1773 ();
 sg13g2_fill_1 FILLER_42_1777 ();
 sg13g2_fill_1 FILLER_42_1791 ();
 sg13g2_decap_8 FILLER_42_1807 ();
 sg13g2_decap_4 FILLER_42_1814 ();
 sg13g2_fill_1 FILLER_42_1818 ();
 sg13g2_decap_4 FILLER_42_1826 ();
 sg13g2_fill_1 FILLER_42_1830 ();
 sg13g2_decap_4 FILLER_42_1835 ();
 sg13g2_fill_2 FILLER_42_1848 ();
 sg13g2_fill_1 FILLER_42_1850 ();
 sg13g2_fill_2 FILLER_42_1862 ();
 sg13g2_fill_2 FILLER_42_1872 ();
 sg13g2_fill_1 FILLER_42_1874 ();
 sg13g2_decap_4 FILLER_42_1890 ();
 sg13g2_fill_2 FILLER_42_1894 ();
 sg13g2_fill_2 FILLER_42_1909 ();
 sg13g2_fill_1 FILLER_42_1911 ();
 sg13g2_fill_2 FILLER_42_1948 ();
 sg13g2_decap_8 FILLER_42_1955 ();
 sg13g2_decap_8 FILLER_42_1962 ();
 sg13g2_fill_1 FILLER_42_1969 ();
 sg13g2_fill_2 FILLER_42_1997 ();
 sg13g2_fill_2 FILLER_42_2032 ();
 sg13g2_fill_1 FILLER_42_2034 ();
 sg13g2_decap_8 FILLER_42_2062 ();
 sg13g2_fill_1 FILLER_42_2069 ();
 sg13g2_decap_4 FILLER_42_2076 ();
 sg13g2_fill_2 FILLER_42_2080 ();
 sg13g2_fill_1 FILLER_42_2092 ();
 sg13g2_fill_2 FILLER_42_2103 ();
 sg13g2_fill_2 FILLER_42_2149 ();
 sg13g2_fill_2 FILLER_42_2164 ();
 sg13g2_decap_4 FILLER_42_2194 ();
 sg13g2_decap_8 FILLER_42_2208 ();
 sg13g2_fill_2 FILLER_42_2221 ();
 sg13g2_fill_1 FILLER_42_2223 ();
 sg13g2_fill_2 FILLER_42_2230 ();
 sg13g2_decap_8 FILLER_42_2236 ();
 sg13g2_decap_8 FILLER_42_2243 ();
 sg13g2_decap_8 FILLER_42_2250 ();
 sg13g2_decap_8 FILLER_42_2283 ();
 sg13g2_fill_1 FILLER_42_2290 ();
 sg13g2_decap_8 FILLER_42_2312 ();
 sg13g2_fill_1 FILLER_42_2334 ();
 sg13g2_fill_1 FILLER_42_2344 ();
 sg13g2_fill_2 FILLER_42_2356 ();
 sg13g2_decap_4 FILLER_42_2371 ();
 sg13g2_fill_2 FILLER_42_2416 ();
 sg13g2_fill_1 FILLER_42_2418 ();
 sg13g2_decap_4 FILLER_42_2439 ();
 sg13g2_fill_2 FILLER_42_2443 ();
 sg13g2_fill_2 FILLER_42_2468 ();
 sg13g2_fill_2 FILLER_42_2474 ();
 sg13g2_fill_1 FILLER_42_2476 ();
 sg13g2_decap_4 FILLER_42_2490 ();
 sg13g2_fill_2 FILLER_42_2494 ();
 sg13g2_decap_8 FILLER_42_2518 ();
 sg13g2_decap_8 FILLER_42_2525 ();
 sg13g2_fill_2 FILLER_42_2540 ();
 sg13g2_fill_2 FILLER_42_2547 ();
 sg13g2_fill_2 FILLER_42_2557 ();
 sg13g2_fill_1 FILLER_42_2559 ();
 sg13g2_fill_2 FILLER_42_2573 ();
 sg13g2_fill_1 FILLER_42_2575 ();
 sg13g2_fill_2 FILLER_42_2597 ();
 sg13g2_fill_1 FILLER_42_2599 ();
 sg13g2_decap_4 FILLER_42_2610 ();
 sg13g2_decap_8 FILLER_42_2618 ();
 sg13g2_fill_2 FILLER_42_2668 ();
 sg13g2_decap_8 FILLER_42_2697 ();
 sg13g2_fill_1 FILLER_42_2704 ();
 sg13g2_decap_8 FILLER_42_2751 ();
 sg13g2_fill_1 FILLER_42_2795 ();
 sg13g2_fill_1 FILLER_42_2802 ();
 sg13g2_fill_2 FILLER_42_2809 ();
 sg13g2_fill_2 FILLER_42_2839 ();
 sg13g2_fill_2 FILLER_42_2849 ();
 sg13g2_decap_4 FILLER_42_2929 ();
 sg13g2_fill_2 FILLER_42_2933 ();
 sg13g2_fill_2 FILLER_42_2975 ();
 sg13g2_fill_1 FILLER_42_2977 ();
 sg13g2_decap_8 FILLER_42_3000 ();
 sg13g2_fill_1 FILLER_42_3007 ();
 sg13g2_fill_2 FILLER_42_3048 ();
 sg13g2_decap_8 FILLER_42_3055 ();
 sg13g2_decap_4 FILLER_42_3062 ();
 sg13g2_fill_1 FILLER_42_3066 ();
 sg13g2_decap_4 FILLER_42_3080 ();
 sg13g2_fill_1 FILLER_42_3084 ();
 sg13g2_fill_1 FILLER_42_3090 ();
 sg13g2_fill_2 FILLER_42_3099 ();
 sg13g2_fill_1 FILLER_42_3101 ();
 sg13g2_decap_8 FILLER_42_3107 ();
 sg13g2_decap_8 FILLER_42_3114 ();
 sg13g2_fill_2 FILLER_42_3121 ();
 sg13g2_fill_1 FILLER_42_3123 ();
 sg13g2_fill_2 FILLER_42_3144 ();
 sg13g2_decap_8 FILLER_42_3159 ();
 sg13g2_fill_1 FILLER_42_3166 ();
 sg13g2_fill_2 FILLER_42_3176 ();
 sg13g2_decap_8 FILLER_42_3182 ();
 sg13g2_fill_2 FILLER_42_3189 ();
 sg13g2_fill_1 FILLER_42_3191 ();
 sg13g2_decap_8 FILLER_42_3195 ();
 sg13g2_decap_4 FILLER_42_3202 ();
 sg13g2_fill_2 FILLER_42_3214 ();
 sg13g2_fill_1 FILLER_42_3216 ();
 sg13g2_fill_2 FILLER_42_3272 ();
 sg13g2_fill_1 FILLER_42_3274 ();
 sg13g2_decap_8 FILLER_42_3287 ();
 sg13g2_fill_2 FILLER_42_3294 ();
 sg13g2_fill_2 FILLER_42_3304 ();
 sg13g2_fill_2 FILLER_42_3318 ();
 sg13g2_fill_1 FILLER_42_3328 ();
 sg13g2_decap_4 FILLER_42_3341 ();
 sg13g2_fill_2 FILLER_42_3345 ();
 sg13g2_decap_8 FILLER_42_3351 ();
 sg13g2_decap_8 FILLER_42_3358 ();
 sg13g2_decap_4 FILLER_42_3365 ();
 sg13g2_fill_1 FILLER_42_3369 ();
 sg13g2_decap_4 FILLER_42_3387 ();
 sg13g2_fill_2 FILLER_42_3391 ();
 sg13g2_fill_1 FILLER_42_3400 ();
 sg13g2_fill_2 FILLER_42_3426 ();
 sg13g2_decap_8 FILLER_42_3458 ();
 sg13g2_fill_1 FILLER_42_3469 ();
 sg13g2_fill_2 FILLER_42_3490 ();
 sg13g2_fill_1 FILLER_42_3492 ();
 sg13g2_fill_1 FILLER_42_3514 ();
 sg13g2_decap_4 FILLER_42_3524 ();
 sg13g2_fill_1 FILLER_42_3528 ();
 sg13g2_fill_1 FILLER_42_3538 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_11 ();
 sg13g2_decap_8 FILLER_43_18 ();
 sg13g2_fill_2 FILLER_43_25 ();
 sg13g2_fill_1 FILLER_43_36 ();
 sg13g2_decap_8 FILLER_43_74 ();
 sg13g2_decap_4 FILLER_43_81 ();
 sg13g2_decap_4 FILLER_43_88 ();
 sg13g2_fill_2 FILLER_43_110 ();
 sg13g2_fill_1 FILLER_43_133 ();
 sg13g2_fill_2 FILLER_43_157 ();
 sg13g2_fill_1 FILLER_43_159 ();
 sg13g2_fill_2 FILLER_43_242 ();
 sg13g2_fill_2 FILLER_43_257 ();
 sg13g2_fill_1 FILLER_43_268 ();
 sg13g2_fill_2 FILLER_43_274 ();
 sg13g2_fill_1 FILLER_43_276 ();
 sg13g2_fill_2 FILLER_43_363 ();
 sg13g2_fill_1 FILLER_43_365 ();
 sg13g2_fill_1 FILLER_43_396 ();
 sg13g2_decap_4 FILLER_43_425 ();
 sg13g2_fill_1 FILLER_43_429 ();
 sg13g2_fill_1 FILLER_43_440 ();
 sg13g2_decap_8 FILLER_43_451 ();
 sg13g2_decap_4 FILLER_43_458 ();
 sg13g2_decap_8 FILLER_43_482 ();
 sg13g2_decap_8 FILLER_43_489 ();
 sg13g2_fill_2 FILLER_43_524 ();
 sg13g2_fill_1 FILLER_43_526 ();
 sg13g2_fill_2 FILLER_43_540 ();
 sg13g2_decap_8 FILLER_43_547 ();
 sg13g2_fill_1 FILLER_43_554 ();
 sg13g2_fill_1 FILLER_43_588 ();
 sg13g2_fill_2 FILLER_43_602 ();
 sg13g2_fill_2 FILLER_43_609 ();
 sg13g2_fill_1 FILLER_43_611 ();
 sg13g2_fill_2 FILLER_43_649 ();
 sg13g2_fill_1 FILLER_43_651 ();
 sg13g2_decap_8 FILLER_43_657 ();
 sg13g2_decap_4 FILLER_43_664 ();
 sg13g2_fill_2 FILLER_43_668 ();
 sg13g2_fill_2 FILLER_43_697 ();
 sg13g2_fill_2 FILLER_43_715 ();
 sg13g2_fill_1 FILLER_43_725 ();
 sg13g2_decap_4 FILLER_43_730 ();
 sg13g2_fill_2 FILLER_43_734 ();
 sg13g2_decap_8 FILLER_43_753 ();
 sg13g2_fill_2 FILLER_43_819 ();
 sg13g2_fill_2 FILLER_43_838 ();
 sg13g2_fill_2 FILLER_43_882 ();
 sg13g2_fill_1 FILLER_43_884 ();
 sg13g2_fill_2 FILLER_43_894 ();
 sg13g2_fill_2 FILLER_43_901 ();
 sg13g2_fill_1 FILLER_43_962 ();
 sg13g2_fill_2 FILLER_43_1019 ();
 sg13g2_fill_1 FILLER_43_1021 ();
 sg13g2_fill_2 FILLER_43_1050 ();
 sg13g2_fill_2 FILLER_43_1090 ();
 sg13g2_fill_1 FILLER_43_1092 ();
 sg13g2_fill_2 FILLER_43_1109 ();
 sg13g2_fill_1 FILLER_43_1111 ();
 sg13g2_fill_2 FILLER_43_1116 ();
 sg13g2_fill_1 FILLER_43_1118 ();
 sg13g2_decap_8 FILLER_43_1126 ();
 sg13g2_fill_2 FILLER_43_1133 ();
 sg13g2_fill_1 FILLER_43_1135 ();
 sg13g2_fill_2 FILLER_43_1139 ();
 sg13g2_fill_1 FILLER_43_1156 ();
 sg13g2_fill_2 FILLER_43_1170 ();
 sg13g2_fill_1 FILLER_43_1172 ();
 sg13g2_decap_4 FILLER_43_1185 ();
 sg13g2_decap_4 FILLER_43_1197 ();
 sg13g2_decap_8 FILLER_43_1206 ();
 sg13g2_fill_1 FILLER_43_1238 ();
 sg13g2_decap_8 FILLER_43_1302 ();
 sg13g2_fill_1 FILLER_43_1309 ();
 sg13g2_decap_8 FILLER_43_1318 ();
 sg13g2_fill_1 FILLER_43_1325 ();
 sg13g2_fill_2 FILLER_43_1330 ();
 sg13g2_fill_1 FILLER_43_1332 ();
 sg13g2_decap_4 FILLER_43_1343 ();
 sg13g2_fill_1 FILLER_43_1365 ();
 sg13g2_fill_2 FILLER_43_1378 ();
 sg13g2_decap_4 FILLER_43_1436 ();
 sg13g2_fill_1 FILLER_43_1440 ();
 sg13g2_decap_8 FILLER_43_1478 ();
 sg13g2_fill_1 FILLER_43_1517 ();
 sg13g2_fill_1 FILLER_43_1531 ();
 sg13g2_fill_1 FILLER_43_1548 ();
 sg13g2_fill_2 FILLER_43_1563 ();
 sg13g2_fill_1 FILLER_43_1565 ();
 sg13g2_decap_8 FILLER_43_1571 ();
 sg13g2_fill_1 FILLER_43_1578 ();
 sg13g2_decap_8 FILLER_43_1595 ();
 sg13g2_decap_4 FILLER_43_1602 ();
 sg13g2_fill_1 FILLER_43_1606 ();
 sg13g2_fill_2 FILLER_43_1612 ();
 sg13g2_fill_1 FILLER_43_1614 ();
 sg13g2_fill_1 FILLER_43_1628 ();
 sg13g2_fill_2 FILLER_43_1633 ();
 sg13g2_fill_1 FILLER_43_1635 ();
 sg13g2_decap_4 FILLER_43_1641 ();
 sg13g2_fill_2 FILLER_43_1645 ();
 sg13g2_decap_8 FILLER_43_1671 ();
 sg13g2_decap_4 FILLER_43_1678 ();
 sg13g2_fill_1 FILLER_43_1682 ();
 sg13g2_decap_8 FILLER_43_1713 ();
 sg13g2_decap_4 FILLER_43_1725 ();
 sg13g2_fill_1 FILLER_43_1729 ();
 sg13g2_fill_2 FILLER_43_1751 ();
 sg13g2_fill_1 FILLER_43_1753 ();
 sg13g2_fill_2 FILLER_43_1764 ();
 sg13g2_decap_8 FILLER_43_1778 ();
 sg13g2_decap_8 FILLER_43_1785 ();
 sg13g2_decap_8 FILLER_43_1792 ();
 sg13g2_fill_2 FILLER_43_1804 ();
 sg13g2_decap_4 FILLER_43_1822 ();
 sg13g2_fill_2 FILLER_43_1831 ();
 sg13g2_fill_1 FILLER_43_1833 ();
 sg13g2_fill_2 FILLER_43_1849 ();
 sg13g2_decap_4 FILLER_43_1867 ();
 sg13g2_fill_2 FILLER_43_1929 ();
 sg13g2_fill_1 FILLER_43_1931 ();
 sg13g2_fill_2 FILLER_43_1963 ();
 sg13g2_fill_1 FILLER_43_1965 ();
 sg13g2_decap_8 FILLER_43_1993 ();
 sg13g2_decap_8 FILLER_43_2000 ();
 sg13g2_fill_2 FILLER_43_2007 ();
 sg13g2_decap_4 FILLER_43_2025 ();
 sg13g2_fill_1 FILLER_43_2029 ();
 sg13g2_fill_2 FILLER_43_2057 ();
 sg13g2_fill_1 FILLER_43_2059 ();
 sg13g2_fill_2 FILLER_43_2081 ();
 sg13g2_decap_8 FILLER_43_2095 ();
 sg13g2_decap_8 FILLER_43_2102 ();
 sg13g2_fill_2 FILLER_43_2109 ();
 sg13g2_fill_1 FILLER_43_2117 ();
 sg13g2_fill_2 FILLER_43_2122 ();
 sg13g2_fill_1 FILLER_43_2124 ();
 sg13g2_decap_4 FILLER_43_2129 ();
 sg13g2_fill_2 FILLER_43_2133 ();
 sg13g2_fill_2 FILLER_43_2151 ();
 sg13g2_fill_1 FILLER_43_2153 ();
 sg13g2_fill_2 FILLER_43_2177 ();
 sg13g2_fill_1 FILLER_43_2179 ();
 sg13g2_fill_2 FILLER_43_2225 ();
 sg13g2_decap_4 FILLER_43_2260 ();
 sg13g2_fill_2 FILLER_43_2290 ();
 sg13g2_fill_1 FILLER_43_2292 ();
 sg13g2_decap_8 FILLER_43_2322 ();
 sg13g2_decap_4 FILLER_43_2329 ();
 sg13g2_fill_2 FILLER_43_2333 ();
 sg13g2_decap_8 FILLER_43_2385 ();
 sg13g2_decap_8 FILLER_43_2392 ();
 sg13g2_fill_1 FILLER_43_2399 ();
 sg13g2_decap_4 FILLER_43_2440 ();
 sg13g2_fill_2 FILLER_43_2444 ();
 sg13g2_fill_1 FILLER_43_2475 ();
 sg13g2_fill_1 FILLER_43_2486 ();
 sg13g2_fill_1 FILLER_43_2496 ();
 sg13g2_fill_2 FILLER_43_2502 ();
 sg13g2_fill_1 FILLER_43_2504 ();
 sg13g2_fill_1 FILLER_43_2512 ();
 sg13g2_decap_4 FILLER_43_2526 ();
 sg13g2_fill_1 FILLER_43_2530 ();
 sg13g2_fill_2 FILLER_43_2540 ();
 sg13g2_fill_1 FILLER_43_2542 ();
 sg13g2_fill_2 FILLER_43_2575 ();
 sg13g2_fill_2 FILLER_43_2581 ();
 sg13g2_fill_1 FILLER_43_2583 ();
 sg13g2_fill_2 FILLER_43_2598 ();
 sg13g2_fill_2 FILLER_43_2608 ();
 sg13g2_fill_1 FILLER_43_2610 ();
 sg13g2_fill_2 FILLER_43_2629 ();
 sg13g2_fill_1 FILLER_43_2631 ();
 sg13g2_fill_1 FILLER_43_2637 ();
 sg13g2_fill_2 FILLER_43_2659 ();
 sg13g2_decap_8 FILLER_43_2684 ();
 sg13g2_fill_2 FILLER_43_2691 ();
 sg13g2_fill_1 FILLER_43_2693 ();
 sg13g2_decap_8 FILLER_43_2749 ();
 sg13g2_fill_1 FILLER_43_2756 ();
 sg13g2_fill_1 FILLER_43_2782 ();
 sg13g2_decap_8 FILLER_43_2822 ();
 sg13g2_fill_2 FILLER_43_2829 ();
 sg13g2_fill_1 FILLER_43_2831 ();
 sg13g2_decap_8 FILLER_43_2840 ();
 sg13g2_fill_2 FILLER_43_2847 ();
 sg13g2_fill_1 FILLER_43_2849 ();
 sg13g2_fill_1 FILLER_43_2863 ();
 sg13g2_decap_4 FILLER_43_2877 ();
 sg13g2_fill_2 FILLER_43_2891 ();
 sg13g2_fill_1 FILLER_43_2893 ();
 sg13g2_fill_2 FILLER_43_2907 ();
 sg13g2_fill_1 FILLER_43_2955 ();
 sg13g2_fill_2 FILLER_43_2961 ();
 sg13g2_decap_4 FILLER_43_2976 ();
 sg13g2_fill_2 FILLER_43_2980 ();
 sg13g2_fill_1 FILLER_43_3030 ();
 sg13g2_decap_8 FILLER_43_3037 ();
 sg13g2_fill_1 FILLER_43_3044 ();
 sg13g2_fill_2 FILLER_43_3097 ();
 sg13g2_decap_8 FILLER_43_3148 ();
 sg13g2_fill_2 FILLER_43_3155 ();
 sg13g2_fill_1 FILLER_43_3276 ();
 sg13g2_fill_1 FILLER_43_3322 ();
 sg13g2_decap_8 FILLER_43_3358 ();
 sg13g2_decap_8 FILLER_43_3365 ();
 sg13g2_fill_2 FILLER_43_3372 ();
 sg13g2_fill_1 FILLER_43_3379 ();
 sg13g2_decap_4 FILLER_43_3389 ();
 sg13g2_fill_2 FILLER_43_3393 ();
 sg13g2_fill_2 FILLER_43_3404 ();
 sg13g2_decap_4 FILLER_43_3422 ();
 sg13g2_fill_1 FILLER_43_3439 ();
 sg13g2_fill_1 FILLER_43_3469 ();
 sg13g2_fill_1 FILLER_43_3479 ();
 sg13g2_fill_2 FILLER_43_3518 ();
 sg13g2_fill_1 FILLER_43_3520 ();
 sg13g2_fill_1 FILLER_43_3535 ();
 sg13g2_decap_8 FILLER_43_3568 ();
 sg13g2_decap_4 FILLER_43_3575 ();
 sg13g2_fill_1 FILLER_43_3579 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_2 ();
 sg13g2_fill_2 FILLER_44_31 ();
 sg13g2_fill_1 FILLER_44_33 ();
 sg13g2_fill_2 FILLER_44_47 ();
 sg13g2_decap_8 FILLER_44_59 ();
 sg13g2_decap_8 FILLER_44_76 ();
 sg13g2_decap_4 FILLER_44_83 ();
 sg13g2_fill_2 FILLER_44_87 ();
 sg13g2_decap_4 FILLER_44_141 ();
 sg13g2_fill_1 FILLER_44_169 ();
 sg13g2_decap_8 FILLER_44_184 ();
 sg13g2_fill_1 FILLER_44_191 ();
 sg13g2_fill_1 FILLER_44_227 ();
 sg13g2_fill_1 FILLER_44_246 ();
 sg13g2_fill_2 FILLER_44_278 ();
 sg13g2_fill_2 FILLER_44_321 ();
 sg13g2_fill_1 FILLER_44_323 ();
 sg13g2_fill_1 FILLER_44_353 ();
 sg13g2_decap_8 FILLER_44_382 ();
 sg13g2_decap_4 FILLER_44_389 ();
 sg13g2_decap_8 FILLER_44_424 ();
 sg13g2_fill_1 FILLER_44_431 ();
 sg13g2_fill_2 FILLER_44_478 ();
 sg13g2_fill_1 FILLER_44_480 ();
 sg13g2_decap_4 FILLER_44_490 ();
 sg13g2_fill_2 FILLER_44_494 ();
 sg13g2_decap_4 FILLER_44_516 ();
 sg13g2_fill_2 FILLER_44_520 ();
 sg13g2_decap_8 FILLER_44_548 ();
 sg13g2_fill_1 FILLER_44_555 ();
 sg13g2_decap_8 FILLER_44_575 ();
 sg13g2_decap_4 FILLER_44_582 ();
 sg13g2_fill_2 FILLER_44_586 ();
 sg13g2_decap_4 FILLER_44_610 ();
 sg13g2_fill_2 FILLER_44_614 ();
 sg13g2_fill_1 FILLER_44_624 ();
 sg13g2_decap_8 FILLER_44_635 ();
 sg13g2_fill_2 FILLER_44_642 ();
 sg13g2_fill_1 FILLER_44_644 ();
 sg13g2_decap_4 FILLER_44_665 ();
 sg13g2_fill_1 FILLER_44_669 ();
 sg13g2_decap_8 FILLER_44_692 ();
 sg13g2_fill_2 FILLER_44_703 ();
 sg13g2_fill_2 FILLER_44_719 ();
 sg13g2_decap_4 FILLER_44_757 ();
 sg13g2_fill_2 FILLER_44_765 ();
 sg13g2_fill_1 FILLER_44_767 ();
 sg13g2_fill_2 FILLER_44_781 ();
 sg13g2_fill_1 FILLER_44_783 ();
 sg13g2_decap_8 FILLER_44_852 ();
 sg13g2_decap_8 FILLER_44_859 ();
 sg13g2_fill_2 FILLER_44_866 ();
 sg13g2_decap_4 FILLER_44_872 ();
 sg13g2_fill_1 FILLER_44_876 ();
 sg13g2_decap_4 FILLER_44_909 ();
 sg13g2_fill_2 FILLER_44_927 ();
 sg13g2_fill_1 FILLER_44_929 ();
 sg13g2_decap_4 FILLER_44_936 ();
 sg13g2_fill_1 FILLER_44_940 ();
 sg13g2_decap_8 FILLER_44_960 ();
 sg13g2_decap_4 FILLER_44_967 ();
 sg13g2_fill_1 FILLER_44_975 ();
 sg13g2_fill_2 FILLER_44_1036 ();
 sg13g2_fill_1 FILLER_44_1087 ();
 sg13g2_fill_2 FILLER_44_1109 ();
 sg13g2_decap_4 FILLER_44_1139 ();
 sg13g2_fill_2 FILLER_44_1143 ();
 sg13g2_decap_4 FILLER_44_1153 ();
 sg13g2_decap_4 FILLER_44_1170 ();
 sg13g2_fill_1 FILLER_44_1174 ();
 sg13g2_fill_1 FILLER_44_1183 ();
 sg13g2_decap_4 FILLER_44_1200 ();
 sg13g2_decap_4 FILLER_44_1301 ();
 sg13g2_fill_1 FILLER_44_1305 ();
 sg13g2_decap_4 FILLER_44_1328 ();
 sg13g2_decap_4 FILLER_44_1337 ();
 sg13g2_decap_4 FILLER_44_1349 ();
 sg13g2_fill_2 FILLER_44_1353 ();
 sg13g2_decap_8 FILLER_44_1368 ();
 sg13g2_decap_4 FILLER_44_1375 ();
 sg13g2_fill_2 FILLER_44_1379 ();
 sg13g2_fill_2 FILLER_44_1394 ();
 sg13g2_fill_1 FILLER_44_1396 ();
 sg13g2_fill_1 FILLER_44_1406 ();
 sg13g2_decap_4 FILLER_44_1429 ();
 sg13g2_fill_2 FILLER_44_1433 ();
 sg13g2_fill_1 FILLER_44_1503 ();
 sg13g2_fill_2 FILLER_44_1518 ();
 sg13g2_fill_1 FILLER_44_1533 ();
 sg13g2_fill_1 FILLER_44_1573 ();
 sg13g2_fill_1 FILLER_44_1602 ();
 sg13g2_fill_2 FILLER_44_1631 ();
 sg13g2_fill_1 FILLER_44_1633 ();
 sg13g2_fill_2 FILLER_44_1651 ();
 sg13g2_fill_2 FILLER_44_1658 ();
 sg13g2_decap_8 FILLER_44_1673 ();
 sg13g2_fill_1 FILLER_44_1680 ();
 sg13g2_fill_2 FILLER_44_1687 ();
 sg13g2_fill_1 FILLER_44_1697 ();
 sg13g2_fill_2 FILLER_44_1707 ();
 sg13g2_fill_1 FILLER_44_1725 ();
 sg13g2_fill_2 FILLER_44_1764 ();
 sg13g2_fill_1 FILLER_44_1766 ();
 sg13g2_fill_2 FILLER_44_1789 ();
 sg13g2_fill_1 FILLER_44_1800 ();
 sg13g2_decap_4 FILLER_44_1822 ();
 sg13g2_fill_1 FILLER_44_1826 ();
 sg13g2_fill_2 FILLER_44_1886 ();
 sg13g2_fill_1 FILLER_44_1888 ();
 sg13g2_fill_1 FILLER_44_1894 ();
 sg13g2_decap_8 FILLER_44_1926 ();
 sg13g2_decap_4 FILLER_44_1933 ();
 sg13g2_fill_1 FILLER_44_1937 ();
 sg13g2_decap_4 FILLER_44_1981 ();
 sg13g2_fill_1 FILLER_44_1985 ();
 sg13g2_fill_1 FILLER_44_2025 ();
 sg13g2_fill_1 FILLER_44_2039 ();
 sg13g2_fill_2 FILLER_44_2044 ();
 sg13g2_fill_2 FILLER_44_2054 ();
 sg13g2_fill_1 FILLER_44_2084 ();
 sg13g2_decap_8 FILLER_44_2102 ();
 sg13g2_fill_2 FILLER_44_2109 ();
 sg13g2_fill_1 FILLER_44_2111 ();
 sg13g2_decap_4 FILLER_44_2125 ();
 sg13g2_fill_1 FILLER_44_2129 ();
 sg13g2_fill_1 FILLER_44_2147 ();
 sg13g2_fill_2 FILLER_44_2155 ();
 sg13g2_decap_4 FILLER_44_2162 ();
 sg13g2_fill_2 FILLER_44_2186 ();
 sg13g2_decap_8 FILLER_44_2213 ();
 sg13g2_fill_2 FILLER_44_2220 ();
 sg13g2_decap_4 FILLER_44_2263 ();
 sg13g2_fill_1 FILLER_44_2299 ();
 sg13g2_decap_4 FILLER_44_2316 ();
 sg13g2_decap_8 FILLER_44_2324 ();
 sg13g2_decap_8 FILLER_44_2331 ();
 sg13g2_fill_1 FILLER_44_2338 ();
 sg13g2_fill_1 FILLER_44_2349 ();
 sg13g2_decap_8 FILLER_44_2409 ();
 sg13g2_decap_4 FILLER_44_2416 ();
 sg13g2_fill_2 FILLER_44_2465 ();
 sg13g2_fill_1 FILLER_44_2467 ();
 sg13g2_fill_2 FILLER_44_2496 ();
 sg13g2_fill_1 FILLER_44_2498 ();
 sg13g2_fill_2 FILLER_44_2504 ();
 sg13g2_fill_1 FILLER_44_2521 ();
 sg13g2_fill_1 FILLER_44_2575 ();
 sg13g2_decap_4 FILLER_44_2579 ();
 sg13g2_fill_1 FILLER_44_2583 ();
 sg13g2_fill_1 FILLER_44_2721 ();
 sg13g2_fill_2 FILLER_44_2784 ();
 sg13g2_fill_1 FILLER_44_2799 ();
 sg13g2_decap_4 FILLER_44_2808 ();
 sg13g2_fill_2 FILLER_44_2829 ();
 sg13g2_decap_4 FILLER_44_2863 ();
 sg13g2_fill_2 FILLER_44_2880 ();
 sg13g2_fill_1 FILLER_44_2910 ();
 sg13g2_decap_8 FILLER_44_2947 ();
 sg13g2_fill_1 FILLER_44_2954 ();
 sg13g2_fill_1 FILLER_44_2958 ();
 sg13g2_fill_1 FILLER_44_3007 ();
 sg13g2_fill_2 FILLER_44_3012 ();
 sg13g2_fill_2 FILLER_44_3047 ();
 sg13g2_fill_2 FILLER_44_3087 ();
 sg13g2_fill_1 FILLER_44_3089 ();
 sg13g2_fill_1 FILLER_44_3110 ();
 sg13g2_fill_2 FILLER_44_3124 ();
 sg13g2_fill_1 FILLER_44_3126 ();
 sg13g2_fill_1 FILLER_44_3132 ();
 sg13g2_decap_8 FILLER_44_3161 ();
 sg13g2_fill_1 FILLER_44_3168 ();
 sg13g2_decap_8 FILLER_44_3173 ();
 sg13g2_fill_2 FILLER_44_3180 ();
 sg13g2_fill_1 FILLER_44_3182 ();
 sg13g2_fill_2 FILLER_44_3188 ();
 sg13g2_fill_1 FILLER_44_3227 ();
 sg13g2_decap_4 FILLER_44_3261 ();
 sg13g2_fill_1 FILLER_44_3265 ();
 sg13g2_decap_4 FILLER_44_3269 ();
 sg13g2_fill_1 FILLER_44_3278 ();
 sg13g2_decap_8 FILLER_44_3285 ();
 sg13g2_decap_4 FILLER_44_3292 ();
 sg13g2_fill_1 FILLER_44_3296 ();
 sg13g2_decap_4 FILLER_44_3305 ();
 sg13g2_decap_4 FILLER_44_3341 ();
 sg13g2_fill_1 FILLER_44_3345 ();
 sg13g2_fill_2 FILLER_44_3374 ();
 sg13g2_fill_1 FILLER_44_3376 ();
 sg13g2_fill_2 FILLER_44_3410 ();
 sg13g2_fill_1 FILLER_44_3412 ();
 sg13g2_fill_1 FILLER_44_3435 ();
 sg13g2_fill_2 FILLER_44_3444 ();
 sg13g2_fill_1 FILLER_44_3446 ();
 sg13g2_fill_2 FILLER_44_3452 ();
 sg13g2_fill_2 FILLER_44_3482 ();
 sg13g2_decap_8 FILLER_44_3488 ();
 sg13g2_fill_1 FILLER_44_3495 ();
 sg13g2_decap_8 FILLER_44_3514 ();
 sg13g2_fill_2 FILLER_44_3521 ();
 sg13g2_fill_2 FILLER_44_3533 ();
 sg13g2_fill_2 FILLER_44_3544 ();
 sg13g2_fill_1 FILLER_44_3546 ();
 sg13g2_fill_2 FILLER_44_3564 ();
 sg13g2_decap_8 FILLER_44_3571 ();
 sg13g2_fill_2 FILLER_44_3578 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_28 ();
 sg13g2_decap_4 FILLER_45_43 ();
 sg13g2_fill_2 FILLER_45_47 ();
 sg13g2_fill_1 FILLER_45_63 ();
 sg13g2_fill_2 FILLER_45_91 ();
 sg13g2_fill_2 FILLER_45_110 ();
 sg13g2_fill_1 FILLER_45_112 ();
 sg13g2_fill_1 FILLER_45_149 ();
 sg13g2_fill_2 FILLER_45_184 ();
 sg13g2_fill_1 FILLER_45_186 ();
 sg13g2_fill_2 FILLER_45_244 ();
 sg13g2_decap_4 FILLER_45_290 ();
 sg13g2_fill_1 FILLER_45_302 ();
 sg13g2_fill_2 FILLER_45_379 ();
 sg13g2_fill_1 FILLER_45_381 ();
 sg13g2_fill_2 FILLER_45_409 ();
 sg13g2_fill_2 FILLER_45_434 ();
 sg13g2_decap_4 FILLER_45_467 ();
 sg13g2_fill_1 FILLER_45_471 ();
 sg13g2_decap_8 FILLER_45_497 ();
 sg13g2_fill_2 FILLER_45_504 ();
 sg13g2_fill_1 FILLER_45_506 ();
 sg13g2_decap_4 FILLER_45_512 ();
 sg13g2_decap_8 FILLER_45_521 ();
 sg13g2_fill_2 FILLER_45_528 ();
 sg13g2_fill_1 FILLER_45_530 ();
 sg13g2_fill_1 FILLER_45_539 ();
 sg13g2_fill_1 FILLER_45_543 ();
 sg13g2_decap_4 FILLER_45_549 ();
 sg13g2_decap_4 FILLER_45_571 ();
 sg13g2_fill_1 FILLER_45_575 ();
 sg13g2_decap_4 FILLER_45_604 ();
 sg13g2_decap_4 FILLER_45_612 ();
 sg13g2_fill_1 FILLER_45_629 ();
 sg13g2_decap_4 FILLER_45_641 ();
 sg13g2_fill_2 FILLER_45_650 ();
 sg13g2_fill_1 FILLER_45_671 ();
 sg13g2_decap_8 FILLER_45_716 ();
 sg13g2_fill_2 FILLER_45_723 ();
 sg13g2_fill_1 FILLER_45_725 ();
 sg13g2_decap_8 FILLER_45_730 ();
 sg13g2_decap_4 FILLER_45_737 ();
 sg13g2_fill_2 FILLER_45_741 ();
 sg13g2_fill_2 FILLER_45_784 ();
 sg13g2_fill_1 FILLER_45_786 ();
 sg13g2_fill_2 FILLER_45_821 ();
 sg13g2_fill_1 FILLER_45_823 ();
 sg13g2_fill_2 FILLER_45_834 ();
 sg13g2_fill_1 FILLER_45_869 ();
 sg13g2_decap_8 FILLER_45_874 ();
 sg13g2_fill_2 FILLER_45_881 ();
 sg13g2_fill_2 FILLER_45_915 ();
 sg13g2_fill_1 FILLER_45_917 ();
 sg13g2_decap_8 FILLER_45_923 ();
 sg13g2_fill_1 FILLER_45_930 ();
 sg13g2_fill_1 FILLER_45_936 ();
 sg13g2_fill_1 FILLER_45_991 ();
 sg13g2_fill_1 FILLER_45_1025 ();
 sg13g2_fill_1 FILLER_45_1059 ();
 sg13g2_fill_2 FILLER_45_1077 ();
 sg13g2_fill_2 FILLER_45_1113 ();
 sg13g2_decap_8 FILLER_45_1122 ();
 sg13g2_fill_2 FILLER_45_1129 ();
 sg13g2_fill_1 FILLER_45_1131 ();
 sg13g2_decap_4 FILLER_45_1142 ();
 sg13g2_fill_1 FILLER_45_1154 ();
 sg13g2_fill_2 FILLER_45_1164 ();
 sg13g2_decap_4 FILLER_45_1170 ();
 sg13g2_decap_8 FILLER_45_1202 ();
 sg13g2_fill_2 FILLER_45_1274 ();
 sg13g2_fill_2 FILLER_45_1284 ();
 sg13g2_fill_1 FILLER_45_1286 ();
 sg13g2_fill_1 FILLER_45_1303 ();
 sg13g2_decap_8 FILLER_45_1309 ();
 sg13g2_decap_8 FILLER_45_1316 ();
 sg13g2_decap_8 FILLER_45_1323 ();
 sg13g2_fill_1 FILLER_45_1330 ();
 sg13g2_decap_8 FILLER_45_1340 ();
 sg13g2_fill_1 FILLER_45_1347 ();
 sg13g2_fill_2 FILLER_45_1354 ();
 sg13g2_decap_8 FILLER_45_1370 ();
 sg13g2_decap_8 FILLER_45_1377 ();
 sg13g2_fill_2 FILLER_45_1384 ();
 sg13g2_fill_2 FILLER_45_1389 ();
 sg13g2_fill_1 FILLER_45_1404 ();
 sg13g2_fill_1 FILLER_45_1437 ();
 sg13g2_decap_4 FILLER_45_1446 ();
 sg13g2_fill_2 FILLER_45_1513 ();
 sg13g2_fill_1 FILLER_45_1515 ();
 sg13g2_decap_4 FILLER_45_1549 ();
 sg13g2_fill_2 FILLER_45_1562 ();
 sg13g2_decap_8 FILLER_45_1570 ();
 sg13g2_fill_1 FILLER_45_1577 ();
 sg13g2_fill_1 FILLER_45_1604 ();
 sg13g2_fill_1 FILLER_45_1618 ();
 sg13g2_decap_8 FILLER_45_1636 ();
 sg13g2_decap_4 FILLER_45_1643 ();
 sg13g2_fill_2 FILLER_45_1660 ();
 sg13g2_fill_2 FILLER_45_1688 ();
 sg13g2_fill_1 FILLER_45_1690 ();
 sg13g2_fill_2 FILLER_45_1699 ();
 sg13g2_decap_4 FILLER_45_1726 ();
 sg13g2_fill_2 FILLER_45_1730 ();
 sg13g2_fill_2 FILLER_45_1749 ();
 sg13g2_fill_1 FILLER_45_1751 ();
 sg13g2_fill_2 FILLER_45_1776 ();
 sg13g2_fill_1 FILLER_45_1778 ();
 sg13g2_decap_4 FILLER_45_1797 ();
 sg13g2_decap_8 FILLER_45_1814 ();
 sg13g2_decap_8 FILLER_45_1821 ();
 sg13g2_fill_1 FILLER_45_1828 ();
 sg13g2_decap_8 FILLER_45_1833 ();
 sg13g2_decap_4 FILLER_45_1840 ();
 sg13g2_fill_1 FILLER_45_1844 ();
 sg13g2_fill_2 FILLER_45_1858 ();
 sg13g2_fill_2 FILLER_45_1869 ();
 sg13g2_fill_1 FILLER_45_1876 ();
 sg13g2_fill_2 FILLER_45_1903 ();
 sg13g2_fill_1 FILLER_45_1905 ();
 sg13g2_decap_4 FILLER_45_1933 ();
 sg13g2_fill_1 FILLER_45_1954 ();
 sg13g2_fill_2 FILLER_45_1965 ();
 sg13g2_fill_1 FILLER_45_1967 ();
 sg13g2_fill_2 FILLER_45_1996 ();
 sg13g2_fill_2 FILLER_45_2068 ();
 sg13g2_fill_1 FILLER_45_2084 ();
 sg13g2_fill_2 FILLER_45_2095 ();
 sg13g2_fill_1 FILLER_45_2097 ();
 sg13g2_fill_2 FILLER_45_2102 ();
 sg13g2_fill_1 FILLER_45_2104 ();
 sg13g2_decap_8 FILLER_45_2121 ();
 sg13g2_fill_2 FILLER_45_2128 ();
 sg13g2_fill_2 FILLER_45_2142 ();
 sg13g2_fill_1 FILLER_45_2144 ();
 sg13g2_decap_4 FILLER_45_2150 ();
 sg13g2_fill_2 FILLER_45_2154 ();
 sg13g2_fill_1 FILLER_45_2162 ();
 sg13g2_decap_4 FILLER_45_2168 ();
 sg13g2_fill_2 FILLER_45_2172 ();
 sg13g2_decap_8 FILLER_45_2186 ();
 sg13g2_fill_1 FILLER_45_2197 ();
 sg13g2_decap_8 FILLER_45_2206 ();
 sg13g2_fill_1 FILLER_45_2213 ();
 sg13g2_fill_2 FILLER_45_2250 ();
 sg13g2_fill_2 FILLER_45_2267 ();
 sg13g2_fill_1 FILLER_45_2274 ();
 sg13g2_decap_8 FILLER_45_2291 ();
 sg13g2_fill_2 FILLER_45_2316 ();
 sg13g2_fill_1 FILLER_45_2318 ();
 sg13g2_fill_1 FILLER_45_2330 ();
 sg13g2_fill_1 FILLER_45_2383 ();
 sg13g2_decap_8 FILLER_45_2388 ();
 sg13g2_fill_2 FILLER_45_2395 ();
 sg13g2_fill_1 FILLER_45_2397 ();
 sg13g2_decap_8 FILLER_45_2439 ();
 sg13g2_fill_2 FILLER_45_2446 ();
 sg13g2_fill_1 FILLER_45_2448 ();
 sg13g2_fill_2 FILLER_45_2454 ();
 sg13g2_fill_1 FILLER_45_2456 ();
 sg13g2_fill_2 FILLER_45_2470 ();
 sg13g2_fill_1 FILLER_45_2472 ();
 sg13g2_fill_2 FILLER_45_2494 ();
 sg13g2_decap_4 FILLER_45_2522 ();
 sg13g2_fill_1 FILLER_45_2563 ();
 sg13g2_fill_2 FILLER_45_2569 ();
 sg13g2_fill_2 FILLER_45_2600 ();
 sg13g2_fill_1 FILLER_45_2619 ();
 sg13g2_fill_2 FILLER_45_2659 ();
 sg13g2_fill_1 FILLER_45_2661 ();
 sg13g2_fill_2 FILLER_45_2705 ();
 sg13g2_fill_1 FILLER_45_2716 ();
 sg13g2_fill_1 FILLER_45_2736 ();
 sg13g2_fill_2 FILLER_45_2745 ();
 sg13g2_fill_1 FILLER_45_2747 ();
 sg13g2_decap_4 FILLER_45_2756 ();
 sg13g2_decap_4 FILLER_45_2781 ();
 sg13g2_fill_2 FILLER_45_2798 ();
 sg13g2_fill_1 FILLER_45_2800 ();
 sg13g2_fill_2 FILLER_45_2842 ();
 sg13g2_fill_2 FILLER_45_2853 ();
 sg13g2_decap_4 FILLER_45_2869 ();
 sg13g2_fill_2 FILLER_45_2873 ();
 sg13g2_fill_2 FILLER_45_2888 ();
 sg13g2_fill_2 FILLER_45_2894 ();
 sg13g2_fill_1 FILLER_45_2896 ();
 sg13g2_fill_2 FILLER_45_2910 ();
 sg13g2_fill_2 FILLER_45_2925 ();
 sg13g2_fill_1 FILLER_45_2927 ();
 sg13g2_fill_1 FILLER_45_2934 ();
 sg13g2_fill_1 FILLER_45_2956 ();
 sg13g2_decap_4 FILLER_45_2975 ();
 sg13g2_fill_2 FILLER_45_2982 ();
 sg13g2_fill_1 FILLER_45_2984 ();
 sg13g2_fill_2 FILLER_45_2994 ();
 sg13g2_fill_1 FILLER_45_3039 ();
 sg13g2_fill_1 FILLER_45_3147 ();
 sg13g2_decap_8 FILLER_45_3156 ();
 sg13g2_fill_1 FILLER_45_3163 ();
 sg13g2_fill_2 FILLER_45_3254 ();
 sg13g2_fill_1 FILLER_45_3256 ();
 sg13g2_fill_2 FILLER_45_3285 ();
 sg13g2_decap_8 FILLER_45_3328 ();
 sg13g2_fill_2 FILLER_45_3335 ();
 sg13g2_fill_1 FILLER_45_3337 ();
 sg13g2_fill_2 FILLER_45_3363 ();
 sg13g2_fill_2 FILLER_45_3375 ();
 sg13g2_fill_1 FILLER_45_3377 ();
 sg13g2_fill_2 FILLER_45_3392 ();
 sg13g2_fill_1 FILLER_45_3394 ();
 sg13g2_decap_8 FILLER_45_3404 ();
 sg13g2_decap_4 FILLER_45_3411 ();
 sg13g2_decap_4 FILLER_45_3443 ();
 sg13g2_fill_1 FILLER_45_3447 ();
 sg13g2_decap_4 FILLER_45_3460 ();
 sg13g2_fill_1 FILLER_45_3464 ();
 sg13g2_fill_2 FILLER_45_3473 ();
 sg13g2_fill_1 FILLER_45_3475 ();
 sg13g2_fill_2 FILLER_45_3493 ();
 sg13g2_fill_1 FILLER_45_3500 ();
 sg13g2_decap_4 FILLER_45_3517 ();
 sg13g2_fill_1 FILLER_45_3521 ();
 sg13g2_fill_2 FILLER_45_3547 ();
 sg13g2_decap_8 FILLER_45_3571 ();
 sg13g2_fill_2 FILLER_45_3578 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_2 ();
 sg13g2_fill_2 FILLER_46_40 ();
 sg13g2_fill_1 FILLER_46_42 ();
 sg13g2_fill_1 FILLER_46_61 ();
 sg13g2_decap_8 FILLER_46_67 ();
 sg13g2_fill_2 FILLER_46_78 ();
 sg13g2_decap_4 FILLER_46_93 ();
 sg13g2_fill_1 FILLER_46_97 ();
 sg13g2_fill_2 FILLER_46_114 ();
 sg13g2_fill_2 FILLER_46_143 ();
 sg13g2_fill_1 FILLER_46_145 ();
 sg13g2_fill_1 FILLER_46_156 ();
 sg13g2_fill_1 FILLER_46_178 ();
 sg13g2_decap_4 FILLER_46_195 ();
 sg13g2_fill_2 FILLER_46_215 ();
 sg13g2_fill_2 FILLER_46_226 ();
 sg13g2_fill_1 FILLER_46_228 ();
 sg13g2_fill_1 FILLER_46_238 ();
 sg13g2_fill_2 FILLER_46_264 ();
 sg13g2_fill_1 FILLER_46_302 ();
 sg13g2_fill_2 FILLER_46_336 ();
 sg13g2_decap_8 FILLER_46_387 ();
 sg13g2_fill_2 FILLER_46_407 ();
 sg13g2_fill_1 FILLER_46_409 ();
 sg13g2_fill_2 FILLER_46_426 ();
 sg13g2_fill_1 FILLER_46_465 ();
 sg13g2_fill_2 FILLER_46_474 ();
 sg13g2_fill_1 FILLER_46_476 ();
 sg13g2_decap_8 FILLER_46_487 ();
 sg13g2_decap_4 FILLER_46_494 ();
 sg13g2_fill_1 FILLER_46_521 ();
 sg13g2_fill_2 FILLER_46_551 ();
 sg13g2_fill_1 FILLER_46_566 ();
 sg13g2_fill_1 FILLER_46_573 ();
 sg13g2_fill_2 FILLER_46_579 ();
 sg13g2_fill_1 FILLER_46_581 ();
 sg13g2_decap_4 FILLER_46_599 ();
 sg13g2_fill_2 FILLER_46_603 ();
 sg13g2_decap_4 FILLER_46_618 ();
 sg13g2_fill_2 FILLER_46_622 ();
 sg13g2_fill_2 FILLER_46_634 ();
 sg13g2_fill_1 FILLER_46_636 ();
 sg13g2_fill_1 FILLER_46_651 ();
 sg13g2_decap_4 FILLER_46_692 ();
 sg13g2_decap_8 FILLER_46_741 ();
 sg13g2_decap_4 FILLER_46_761 ();
 sg13g2_fill_1 FILLER_46_770 ();
 sg13g2_fill_1 FILLER_46_812 ();
 sg13g2_fill_1 FILLER_46_850 ();
 sg13g2_fill_1 FILLER_46_864 ();
 sg13g2_fill_1 FILLER_46_893 ();
 sg13g2_fill_2 FILLER_46_938 ();
 sg13g2_fill_1 FILLER_46_940 ();
 sg13g2_fill_2 FILLER_46_946 ();
 sg13g2_fill_2 FILLER_46_957 ();
 sg13g2_fill_1 FILLER_46_959 ();
 sg13g2_decap_8 FILLER_46_969 ();
 sg13g2_fill_2 FILLER_46_976 ();
 sg13g2_fill_1 FILLER_46_978 ();
 sg13g2_decap_4 FILLER_46_1011 ();
 sg13g2_fill_2 FILLER_46_1044 ();
 sg13g2_fill_1 FILLER_46_1046 ();
 sg13g2_fill_1 FILLER_46_1051 ();
 sg13g2_fill_2 FILLER_46_1075 ();
 sg13g2_fill_1 FILLER_46_1077 ();
 sg13g2_decap_4 FILLER_46_1138 ();
 sg13g2_decap_4 FILLER_46_1150 ();
 sg13g2_decap_4 FILLER_46_1190 ();
 sg13g2_fill_2 FILLER_46_1194 ();
 sg13g2_fill_1 FILLER_46_1222 ();
 sg13g2_fill_2 FILLER_46_1249 ();
 sg13g2_fill_1 FILLER_46_1302 ();
 sg13g2_fill_1 FILLER_46_1311 ();
 sg13g2_fill_1 FILLER_46_1378 ();
 sg13g2_decap_4 FILLER_46_1406 ();
 sg13g2_fill_1 FILLER_46_1410 ();
 sg13g2_fill_2 FILLER_46_1423 ();
 sg13g2_fill_2 FILLER_46_1460 ();
 sg13g2_fill_2 FILLER_46_1489 ();
 sg13g2_fill_1 FILLER_46_1491 ();
 sg13g2_decap_8 FILLER_46_1548 ();
 sg13g2_decap_8 FILLER_46_1555 ();
 sg13g2_fill_2 FILLER_46_1570 ();
 sg13g2_fill_1 FILLER_46_1572 ();
 sg13g2_decap_8 FILLER_46_1581 ();
 sg13g2_decap_4 FILLER_46_1588 ();
 sg13g2_fill_2 FILLER_46_1592 ();
 sg13g2_fill_2 FILLER_46_1607 ();
 sg13g2_fill_1 FILLER_46_1622 ();
 sg13g2_fill_1 FILLER_46_1627 ();
 sg13g2_fill_2 FILLER_46_1649 ();
 sg13g2_fill_2 FILLER_46_1671 ();
 sg13g2_fill_1 FILLER_46_1673 ();
 sg13g2_decap_4 FILLER_46_1718 ();
 sg13g2_fill_1 FILLER_46_1722 ();
 sg13g2_fill_1 FILLER_46_1735 ();
 sg13g2_fill_1 FILLER_46_1740 ();
 sg13g2_fill_1 FILLER_46_1754 ();
 sg13g2_fill_2 FILLER_46_1761 ();
 sg13g2_decap_4 FILLER_46_1768 ();
 sg13g2_fill_1 FILLER_46_1794 ();
 sg13g2_fill_2 FILLER_46_1809 ();
 sg13g2_fill_1 FILLER_46_1811 ();
 sg13g2_fill_2 FILLER_46_1854 ();
 sg13g2_fill_1 FILLER_46_1856 ();
 sg13g2_fill_2 FILLER_46_2002 ();
 sg13g2_fill_1 FILLER_46_2004 ();
 sg13g2_fill_1 FILLER_46_2033 ();
 sg13g2_fill_2 FILLER_46_2047 ();
 sg13g2_fill_1 FILLER_46_2049 ();
 sg13g2_decap_4 FILLER_46_2060 ();
 sg13g2_fill_2 FILLER_46_2064 ();
 sg13g2_fill_2 FILLER_46_2088 ();
 sg13g2_fill_1 FILLER_46_2099 ();
 sg13g2_fill_2 FILLER_46_2116 ();
 sg13g2_fill_2 FILLER_46_2131 ();
 sg13g2_fill_1 FILLER_46_2133 ();
 sg13g2_fill_2 FILLER_46_2155 ();
 sg13g2_fill_1 FILLER_46_2157 ();
 sg13g2_decap_4 FILLER_46_2166 ();
 sg13g2_fill_1 FILLER_46_2181 ();
 sg13g2_decap_8 FILLER_46_2190 ();
 sg13g2_fill_2 FILLER_46_2197 ();
 sg13g2_decap_4 FILLER_46_2204 ();
 sg13g2_fill_1 FILLER_46_2208 ();
 sg13g2_fill_2 FILLER_46_2231 ();
 sg13g2_fill_2 FILLER_46_2245 ();
 sg13g2_fill_1 FILLER_46_2255 ();
 sg13g2_decap_8 FILLER_46_2264 ();
 sg13g2_decap_8 FILLER_46_2271 ();
 sg13g2_decap_8 FILLER_46_2278 ();
 sg13g2_fill_2 FILLER_46_2285 ();
 sg13g2_decap_4 FILLER_46_2300 ();
 sg13g2_decap_8 FILLER_46_2310 ();
 sg13g2_fill_2 FILLER_46_2317 ();
 sg13g2_fill_2 FILLER_46_2346 ();
 sg13g2_fill_1 FILLER_46_2348 ();
 sg13g2_decap_8 FILLER_46_2376 ();
 sg13g2_fill_2 FILLER_46_2383 ();
 sg13g2_fill_2 FILLER_46_2398 ();
 sg13g2_fill_1 FILLER_46_2400 ();
 sg13g2_fill_1 FILLER_46_2419 ();
 sg13g2_fill_2 FILLER_46_2428 ();
 sg13g2_decap_8 FILLER_46_2448 ();
 sg13g2_decap_4 FILLER_46_2455 ();
 sg13g2_fill_2 FILLER_46_2459 ();
 sg13g2_fill_1 FILLER_46_2487 ();
 sg13g2_decap_4 FILLER_46_2492 ();
 sg13g2_fill_2 FILLER_46_2496 ();
 sg13g2_decap_4 FILLER_46_2522 ();
 sg13g2_fill_2 FILLER_46_2526 ();
 sg13g2_fill_2 FILLER_46_2532 ();
 sg13g2_fill_2 FILLER_46_2542 ();
 sg13g2_fill_1 FILLER_46_2544 ();
 sg13g2_fill_2 FILLER_46_2553 ();
 sg13g2_fill_1 FILLER_46_2573 ();
 sg13g2_decap_8 FILLER_46_2588 ();
 sg13g2_fill_1 FILLER_46_2665 ();
 sg13g2_fill_2 FILLER_46_2675 ();
 sg13g2_fill_2 FILLER_46_2690 ();
 sg13g2_fill_2 FILLER_46_2727 ();
 sg13g2_fill_2 FILLER_46_2746 ();
 sg13g2_decap_4 FILLER_46_2764 ();
 sg13g2_decap_4 FILLER_46_2776 ();
 sg13g2_fill_2 FILLER_46_2780 ();
 sg13g2_fill_2 FILLER_46_2819 ();
 sg13g2_fill_1 FILLER_46_2834 ();
 sg13g2_fill_2 FILLER_46_2843 ();
 sg13g2_fill_1 FILLER_46_2923 ();
 sg13g2_fill_2 FILLER_46_3000 ();
 sg13g2_fill_1 FILLER_46_3002 ();
 sg13g2_fill_2 FILLER_46_3055 ();
 sg13g2_fill_1 FILLER_46_3085 ();
 sg13g2_fill_1 FILLER_46_3109 ();
 sg13g2_fill_1 FILLER_46_3120 ();
 sg13g2_decap_8 FILLER_46_3133 ();
 sg13g2_fill_2 FILLER_46_3140 ();
 sg13g2_fill_1 FILLER_46_3142 ();
 sg13g2_decap_8 FILLER_46_3168 ();
 sg13g2_decap_8 FILLER_46_3175 ();
 sg13g2_decap_4 FILLER_46_3182 ();
 sg13g2_fill_1 FILLER_46_3186 ();
 sg13g2_fill_2 FILLER_46_3197 ();
 sg13g2_fill_1 FILLER_46_3227 ();
 sg13g2_fill_2 FILLER_46_3233 ();
 sg13g2_decap_4 FILLER_46_3279 ();
 sg13g2_fill_2 FILLER_46_3283 ();
 sg13g2_fill_2 FILLER_46_3299 ();
 sg13g2_fill_1 FILLER_46_3301 ();
 sg13g2_fill_1 FILLER_46_3315 ();
 sg13g2_fill_2 FILLER_46_3336 ();
 sg13g2_fill_2 FILLER_46_3370 ();
 sg13g2_fill_2 FILLER_46_3388 ();
 sg13g2_fill_2 FILLER_46_3398 ();
 sg13g2_fill_1 FILLER_46_3400 ();
 sg13g2_decap_4 FILLER_46_3413 ();
 sg13g2_fill_2 FILLER_46_3417 ();
 sg13g2_fill_1 FILLER_46_3447 ();
 sg13g2_decap_4 FILLER_46_3457 ();
 sg13g2_fill_1 FILLER_46_3461 ();
 sg13g2_fill_2 FILLER_46_3470 ();
 sg13g2_fill_1 FILLER_46_3472 ();
 sg13g2_decap_8 FILLER_46_3483 ();
 sg13g2_fill_1 FILLER_46_3502 ();
 sg13g2_fill_2 FILLER_46_3512 ();
 sg13g2_fill_1 FILLER_46_3514 ();
 sg13g2_decap_8 FILLER_46_3519 ();
 sg13g2_decap_4 FILLER_46_3526 ();
 sg13g2_decap_4 FILLER_46_3540 ();
 sg13g2_fill_2 FILLER_46_3559 ();
 sg13g2_fill_2 FILLER_46_3577 ();
 sg13g2_fill_1 FILLER_46_3579 ();
 sg13g2_decap_4 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_4 ();
 sg13g2_fill_2 FILLER_47_33 ();
 sg13g2_fill_2 FILLER_47_47 ();
 sg13g2_decap_4 FILLER_47_68 ();
 sg13g2_decap_4 FILLER_47_88 ();
 sg13g2_fill_1 FILLER_47_131 ();
 sg13g2_fill_2 FILLER_47_168 ();
 sg13g2_fill_2 FILLER_47_232 ();
 sg13g2_fill_2 FILLER_47_319 ();
 sg13g2_fill_1 FILLER_47_334 ();
 sg13g2_fill_2 FILLER_47_370 ();
 sg13g2_fill_1 FILLER_47_424 ();
 sg13g2_fill_1 FILLER_47_432 ();
 sg13g2_decap_8 FILLER_47_456 ();
 sg13g2_fill_2 FILLER_47_463 ();
 sg13g2_fill_1 FILLER_47_465 ();
 sg13g2_fill_1 FILLER_47_478 ();
 sg13g2_fill_1 FILLER_47_489 ();
 sg13g2_decap_8 FILLER_47_510 ();
 sg13g2_fill_2 FILLER_47_517 ();
 sg13g2_fill_1 FILLER_47_519 ();
 sg13g2_fill_2 FILLER_47_537 ();
 sg13g2_fill_1 FILLER_47_539 ();
 sg13g2_decap_8 FILLER_47_567 ();
 sg13g2_decap_4 FILLER_47_574 ();
 sg13g2_fill_1 FILLER_47_623 ();
 sg13g2_fill_1 FILLER_47_678 ();
 sg13g2_fill_1 FILLER_47_716 ();
 sg13g2_fill_2 FILLER_47_750 ();
 sg13g2_fill_2 FILLER_47_765 ();
 sg13g2_fill_1 FILLER_47_767 ();
 sg13g2_fill_2 FILLER_47_794 ();
 sg13g2_fill_1 FILLER_47_796 ();
 sg13g2_decap_4 FILLER_47_838 ();
 sg13g2_fill_1 FILLER_47_875 ();
 sg13g2_decap_4 FILLER_47_942 ();
 sg13g2_fill_1 FILLER_47_946 ();
 sg13g2_decap_4 FILLER_47_974 ();
 sg13g2_decap_8 FILLER_47_1003 ();
 sg13g2_fill_2 FILLER_47_1010 ();
 sg13g2_fill_1 FILLER_47_1018 ();
 sg13g2_fill_2 FILLER_47_1040 ();
 sg13g2_decap_8 FILLER_47_1055 ();
 sg13g2_fill_2 FILLER_47_1062 ();
 sg13g2_fill_1 FILLER_47_1064 ();
 sg13g2_fill_1 FILLER_47_1104 ();
 sg13g2_fill_2 FILLER_47_1167 ();
 sg13g2_fill_1 FILLER_47_1169 ();
 sg13g2_fill_2 FILLER_47_1274 ();
 sg13g2_fill_2 FILLER_47_1284 ();
 sg13g2_fill_2 FILLER_47_1296 ();
 sg13g2_fill_2 FILLER_47_1308 ();
 sg13g2_fill_1 FILLER_47_1310 ();
 sg13g2_fill_2 FILLER_47_1324 ();
 sg13g2_fill_2 FILLER_47_1351 ();
 sg13g2_decap_4 FILLER_47_1372 ();
 sg13g2_fill_2 FILLER_47_1389 ();
 sg13g2_fill_1 FILLER_47_1417 ();
 sg13g2_fill_2 FILLER_47_1436 ();
 sg13g2_fill_1 FILLER_47_1438 ();
 sg13g2_fill_2 FILLER_47_1495 ();
 sg13g2_fill_1 FILLER_47_1497 ();
 sg13g2_fill_1 FILLER_47_1512 ();
 sg13g2_decap_4 FILLER_47_1531 ();
 sg13g2_fill_1 FILLER_47_1535 ();
 sg13g2_fill_1 FILLER_47_1576 ();
 sg13g2_fill_1 FILLER_47_1585 ();
 sg13g2_fill_1 FILLER_47_1655 ();
 sg13g2_fill_2 FILLER_47_1684 ();
 sg13g2_fill_1 FILLER_47_1686 ();
 sg13g2_fill_1 FILLER_47_1724 ();
 sg13g2_fill_1 FILLER_47_1748 ();
 sg13g2_fill_1 FILLER_47_1777 ();
 sg13g2_fill_2 FILLER_47_1818 ();
 sg13g2_fill_1 FILLER_47_1820 ();
 sg13g2_fill_1 FILLER_47_1826 ();
 sg13g2_fill_1 FILLER_47_1891 ();
 sg13g2_fill_2 FILLER_47_1929 ();
 sg13g2_fill_1 FILLER_47_1931 ();
 sg13g2_fill_2 FILLER_47_1964 ();
 sg13g2_fill_1 FILLER_47_1994 ();
 sg13g2_fill_1 FILLER_47_2036 ();
 sg13g2_fill_2 FILLER_47_2059 ();
 sg13g2_fill_2 FILLER_47_2104 ();
 sg13g2_fill_2 FILLER_47_2116 ();
 sg13g2_fill_2 FILLER_47_2123 ();
 sg13g2_fill_1 FILLER_47_2125 ();
 sg13g2_decap_8 FILLER_47_2139 ();
 sg13g2_decap_8 FILLER_47_2146 ();
 sg13g2_decap_8 FILLER_47_2153 ();
 sg13g2_decap_8 FILLER_47_2165 ();
 sg13g2_fill_2 FILLER_47_2172 ();
 sg13g2_fill_1 FILLER_47_2174 ();
 sg13g2_fill_1 FILLER_47_2179 ();
 sg13g2_fill_1 FILLER_47_2185 ();
 sg13g2_fill_2 FILLER_47_2219 ();
 sg13g2_fill_2 FILLER_47_2229 ();
 sg13g2_fill_1 FILLER_47_2231 ();
 sg13g2_fill_2 FILLER_47_2248 ();
 sg13g2_fill_1 FILLER_47_2250 ();
 sg13g2_fill_1 FILLER_47_2264 ();
 sg13g2_fill_2 FILLER_47_2285 ();
 sg13g2_decap_4 FILLER_47_2339 ();
 sg13g2_fill_1 FILLER_47_2343 ();
 sg13g2_decap_8 FILLER_47_2348 ();
 sg13g2_fill_1 FILLER_47_2355 ();
 sg13g2_decap_4 FILLER_47_2377 ();
 sg13g2_fill_1 FILLER_47_2416 ();
 sg13g2_fill_2 FILLER_47_2429 ();
 sg13g2_decap_8 FILLER_47_2457 ();
 sg13g2_fill_1 FILLER_47_2477 ();
 sg13g2_decap_8 FILLER_47_2515 ();
 sg13g2_fill_2 FILLER_47_2522 ();
 sg13g2_fill_2 FILLER_47_2545 ();
 sg13g2_fill_1 FILLER_47_2552 ();
 sg13g2_decap_8 FILLER_47_2584 ();
 sg13g2_decap_4 FILLER_47_2591 ();
 sg13g2_fill_1 FILLER_47_2595 ();
 sg13g2_fill_1 FILLER_47_2620 ();
 sg13g2_fill_2 FILLER_47_2625 ();
 sg13g2_fill_1 FILLER_47_2627 ();
 sg13g2_decap_4 FILLER_47_2660 ();
 sg13g2_decap_8 FILLER_47_2692 ();
 sg13g2_decap_4 FILLER_47_2699 ();
 sg13g2_fill_2 FILLER_47_2703 ();
 sg13g2_decap_4 FILLER_47_2779 ();
 sg13g2_fill_2 FILLER_47_2783 ();
 sg13g2_fill_2 FILLER_47_2812 ();
 sg13g2_fill_1 FILLER_47_2814 ();
 sg13g2_fill_1 FILLER_47_2867 ();
 sg13g2_fill_2 FILLER_47_2890 ();
 sg13g2_decap_8 FILLER_47_2906 ();
 sg13g2_fill_2 FILLER_47_2913 ();
 sg13g2_fill_2 FILLER_47_2924 ();
 sg13g2_fill_1 FILLER_47_2926 ();
 sg13g2_fill_2 FILLER_47_2939 ();
 sg13g2_fill_1 FILLER_47_2941 ();
 sg13g2_decap_4 FILLER_47_2958 ();
 sg13g2_decap_8 FILLER_47_2967 ();
 sg13g2_fill_1 FILLER_47_2974 ();
 sg13g2_decap_8 FILLER_47_2980 ();
 sg13g2_decap_4 FILLER_47_2987 ();
 sg13g2_fill_1 FILLER_47_2991 ();
 sg13g2_fill_2 FILLER_47_2997 ();
 sg13g2_fill_2 FILLER_47_3035 ();
 sg13g2_fill_1 FILLER_47_3046 ();
 sg13g2_fill_1 FILLER_47_3057 ();
 sg13g2_decap_4 FILLER_47_3067 ();
 sg13g2_decap_8 FILLER_47_3083 ();
 sg13g2_decap_8 FILLER_47_3090 ();
 sg13g2_fill_2 FILLER_47_3097 ();
 sg13g2_decap_8 FILLER_47_3137 ();
 sg13g2_decap_4 FILLER_47_3144 ();
 sg13g2_fill_1 FILLER_47_3148 ();
 sg13g2_fill_1 FILLER_47_3179 ();
 sg13g2_fill_2 FILLER_47_3196 ();
 sg13g2_fill_1 FILLER_47_3198 ();
 sg13g2_fill_1 FILLER_47_3202 ();
 sg13g2_fill_1 FILLER_47_3212 ();
 sg13g2_fill_1 FILLER_47_3226 ();
 sg13g2_decap_8 FILLER_47_3327 ();
 sg13g2_fill_1 FILLER_47_3334 ();
 sg13g2_decap_4 FILLER_47_3339 ();
 sg13g2_fill_1 FILLER_47_3369 ();
 sg13g2_decap_8 FILLER_47_3375 ();
 sg13g2_fill_1 FILLER_47_3387 ();
 sg13g2_decap_8 FILLER_47_3404 ();
 sg13g2_fill_1 FILLER_47_3411 ();
 sg13g2_decap_8 FILLER_47_3424 ();
 sg13g2_decap_8 FILLER_47_3431 ();
 sg13g2_fill_1 FILLER_47_3438 ();
 sg13g2_fill_2 FILLER_47_3459 ();
 sg13g2_fill_1 FILLER_47_3487 ();
 sg13g2_fill_1 FILLER_47_3501 ();
 sg13g2_fill_2 FILLER_47_3527 ();
 sg13g2_decap_8 FILLER_47_3542 ();
 sg13g2_fill_2 FILLER_47_3549 ();
 sg13g2_fill_1 FILLER_47_3579 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_7 ();
 sg13g2_fill_1 FILLER_48_9 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_fill_2 FILLER_48_21 ();
 sg13g2_fill_2 FILLER_48_35 ();
 sg13g2_decap_4 FILLER_48_70 ();
 sg13g2_fill_2 FILLER_48_94 ();
 sg13g2_fill_1 FILLER_48_96 ();
 sg13g2_fill_1 FILLER_48_136 ();
 sg13g2_fill_2 FILLER_48_157 ();
 sg13g2_fill_1 FILLER_48_174 ();
 sg13g2_fill_2 FILLER_48_203 ();
 sg13g2_fill_1 FILLER_48_205 ();
 sg13g2_decap_4 FILLER_48_215 ();
 sg13g2_fill_1 FILLER_48_228 ();
 sg13g2_fill_1 FILLER_48_239 ();
 sg13g2_decap_4 FILLER_48_255 ();
 sg13g2_fill_2 FILLER_48_259 ();
 sg13g2_fill_2 FILLER_48_280 ();
 sg13g2_fill_1 FILLER_48_310 ();
 sg13g2_fill_2 FILLER_48_348 ();
 sg13g2_fill_2 FILLER_48_390 ();
 sg13g2_fill_2 FILLER_48_409 ();
 sg13g2_fill_1 FILLER_48_411 ();
 sg13g2_fill_2 FILLER_48_427 ();
 sg13g2_fill_1 FILLER_48_429 ();
 sg13g2_fill_1 FILLER_48_435 ();
 sg13g2_fill_2 FILLER_48_452 ();
 sg13g2_fill_1 FILLER_48_454 ();
 sg13g2_fill_2 FILLER_48_472 ();
 sg13g2_fill_1 FILLER_48_474 ();
 sg13g2_decap_4 FILLER_48_489 ();
 sg13g2_fill_2 FILLER_48_493 ();
 sg13g2_fill_1 FILLER_48_504 ();
 sg13g2_decap_4 FILLER_48_514 ();
 sg13g2_decap_8 FILLER_48_541 ();
 sg13g2_fill_2 FILLER_48_548 ();
 sg13g2_fill_1 FILLER_48_550 ();
 sg13g2_decap_8 FILLER_48_572 ();
 sg13g2_fill_2 FILLER_48_579 ();
 sg13g2_fill_1 FILLER_48_594 ();
 sg13g2_fill_1 FILLER_48_619 ();
 sg13g2_decap_4 FILLER_48_650 ();
 sg13g2_fill_1 FILLER_48_680 ();
 sg13g2_decap_4 FILLER_48_743 ();
 sg13g2_fill_2 FILLER_48_747 ();
 sg13g2_fill_1 FILLER_48_762 ();
 sg13g2_fill_1 FILLER_48_786 ();
 sg13g2_decap_8 FILLER_48_795 ();
 sg13g2_decap_8 FILLER_48_807 ();
 sg13g2_fill_2 FILLER_48_837 ();
 sg13g2_fill_1 FILLER_48_839 ();
 sg13g2_fill_1 FILLER_48_854 ();
 sg13g2_fill_2 FILLER_48_901 ();
 sg13g2_fill_1 FILLER_48_911 ();
 sg13g2_decap_8 FILLER_48_947 ();
 sg13g2_fill_2 FILLER_48_954 ();
 sg13g2_fill_1 FILLER_48_956 ();
 sg13g2_decap_8 FILLER_48_969 ();
 sg13g2_decap_4 FILLER_48_976 ();
 sg13g2_fill_1 FILLER_48_980 ();
 sg13g2_decap_4 FILLER_48_1001 ();
 sg13g2_fill_1 FILLER_48_1005 ();
 sg13g2_fill_1 FILLER_48_1014 ();
 sg13g2_fill_2 FILLER_48_1035 ();
 sg13g2_fill_1 FILLER_48_1037 ();
 sg13g2_decap_4 FILLER_48_1050 ();
 sg13g2_fill_2 FILLER_48_1070 ();
 sg13g2_fill_2 FILLER_48_1184 ();
 sg13g2_fill_1 FILLER_48_1199 ();
 sg13g2_decap_4 FILLER_48_1222 ();
 sg13g2_fill_1 FILLER_48_1226 ();
 sg13g2_fill_1 FILLER_48_1248 ();
 sg13g2_fill_2 FILLER_48_1304 ();
 sg13g2_fill_1 FILLER_48_1306 ();
 sg13g2_fill_2 FILLER_48_1357 ();
 sg13g2_fill_1 FILLER_48_1359 ();
 sg13g2_fill_1 FILLER_48_1400 ();
 sg13g2_fill_2 FILLER_48_1414 ();
 sg13g2_decap_8 FILLER_48_1442 ();
 sg13g2_fill_2 FILLER_48_1463 ();
 sg13g2_fill_1 FILLER_48_1465 ();
 sg13g2_fill_2 FILLER_48_1479 ();
 sg13g2_fill_2 FILLER_48_1532 ();
 sg13g2_fill_1 FILLER_48_1534 ();
 sg13g2_decap_4 FILLER_48_1548 ();
 sg13g2_fill_1 FILLER_48_1552 ();
 sg13g2_fill_1 FILLER_48_1562 ();
 sg13g2_fill_1 FILLER_48_1568 ();
 sg13g2_decap_4 FILLER_48_1594 ();
 sg13g2_fill_2 FILLER_48_1632 ();
 sg13g2_fill_1 FILLER_48_1634 ();
 sg13g2_fill_1 FILLER_48_1663 ();
 sg13g2_fill_1 FILLER_48_1695 ();
 sg13g2_fill_2 FILLER_48_1733 ();
 sg13g2_decap_8 FILLER_48_1767 ();
 sg13g2_fill_2 FILLER_48_1774 ();
 sg13g2_fill_1 FILLER_48_1793 ();
 sg13g2_fill_2 FILLER_48_1849 ();
 sg13g2_fill_1 FILLER_48_1884 ();
 sg13g2_fill_2 FILLER_48_1896 ();
 sg13g2_fill_1 FILLER_48_1898 ();
 sg13g2_fill_2 FILLER_48_1953 ();
 sg13g2_fill_2 FILLER_48_2001 ();
 sg13g2_fill_2 FILLER_48_2074 ();
 sg13g2_fill_1 FILLER_48_2076 ();
 sg13g2_fill_1 FILLER_48_2146 ();
 sg13g2_decap_8 FILLER_48_2163 ();
 sg13g2_fill_2 FILLER_48_2170 ();
 sg13g2_fill_1 FILLER_48_2172 ();
 sg13g2_fill_2 FILLER_48_2198 ();
 sg13g2_fill_1 FILLER_48_2200 ();
 sg13g2_decap_4 FILLER_48_2206 ();
 sg13g2_fill_2 FILLER_48_2210 ();
 sg13g2_fill_2 FILLER_48_2234 ();
 sg13g2_fill_2 FILLER_48_2241 ();
 sg13g2_fill_1 FILLER_48_2243 ();
 sg13g2_decap_8 FILLER_48_2267 ();
 sg13g2_decap_8 FILLER_48_2274 ();
 sg13g2_fill_2 FILLER_48_2288 ();
 sg13g2_fill_1 FILLER_48_2290 ();
 sg13g2_decap_4 FILLER_48_2321 ();
 sg13g2_decap_4 FILLER_48_2333 ();
 sg13g2_fill_2 FILLER_48_2356 ();
 sg13g2_fill_2 FILLER_48_2380 ();
 sg13g2_fill_1 FILLER_48_2382 ();
 sg13g2_fill_2 FILLER_48_2391 ();
 sg13g2_fill_1 FILLER_48_2393 ();
 sg13g2_fill_2 FILLER_48_2418 ();
 sg13g2_fill_1 FILLER_48_2420 ();
 sg13g2_decap_4 FILLER_48_2432 ();
 sg13g2_decap_8 FILLER_48_2448 ();
 sg13g2_decap_8 FILLER_48_2455 ();
 sg13g2_fill_1 FILLER_48_2462 ();
 sg13g2_decap_8 FILLER_48_2480 ();
 sg13g2_decap_4 FILLER_48_2487 ();
 sg13g2_decap_4 FILLER_48_2495 ();
 sg13g2_fill_1 FILLER_48_2540 ();
 sg13g2_decap_8 FILLER_48_2563 ();
 sg13g2_fill_1 FILLER_48_2587 ();
 sg13g2_fill_1 FILLER_48_2601 ();
 sg13g2_decap_4 FILLER_48_2625 ();
 sg13g2_fill_2 FILLER_48_2629 ();
 sg13g2_fill_2 FILLER_48_2683 ();
 sg13g2_fill_1 FILLER_48_2685 ();
 sg13g2_fill_1 FILLER_48_2692 ();
 sg13g2_fill_2 FILLER_48_2715 ();
 sg13g2_fill_1 FILLER_48_2717 ();
 sg13g2_fill_2 FILLER_48_2727 ();
 sg13g2_decap_4 FILLER_48_2789 ();
 sg13g2_fill_1 FILLER_48_2793 ();
 sg13g2_fill_2 FILLER_48_2797 ();
 sg13g2_fill_2 FILLER_48_2804 ();
 sg13g2_fill_1 FILLER_48_2806 ();
 sg13g2_decap_4 FILLER_48_2816 ();
 sg13g2_fill_1 FILLER_48_2820 ();
 sg13g2_decap_8 FILLER_48_2834 ();
 sg13g2_fill_2 FILLER_48_2841 ();
 sg13g2_fill_1 FILLER_48_2843 ();
 sg13g2_fill_1 FILLER_48_2875 ();
 sg13g2_decap_4 FILLER_48_2909 ();
 sg13g2_fill_1 FILLER_48_2913 ();
 sg13g2_fill_2 FILLER_48_2999 ();
 sg13g2_fill_1 FILLER_48_3001 ();
 sg13g2_decap_4 FILLER_48_3011 ();
 sg13g2_fill_2 FILLER_48_3015 ();
 sg13g2_fill_1 FILLER_48_3022 ();
 sg13g2_fill_1 FILLER_48_3034 ();
 sg13g2_decap_8 FILLER_48_3039 ();
 sg13g2_decap_4 FILLER_48_3046 ();
 sg13g2_fill_1 FILLER_48_3050 ();
 sg13g2_fill_2 FILLER_48_3082 ();
 sg13g2_fill_2 FILLER_48_3104 ();
 sg13g2_fill_2 FILLER_48_3117 ();
 sg13g2_fill_2 FILLER_48_3145 ();
 sg13g2_fill_2 FILLER_48_3156 ();
 sg13g2_fill_1 FILLER_48_3158 ();
 sg13g2_decap_8 FILLER_48_3168 ();
 sg13g2_decap_4 FILLER_48_3175 ();
 sg13g2_fill_1 FILLER_48_3179 ();
 sg13g2_decap_8 FILLER_48_3193 ();
 sg13g2_decap_4 FILLER_48_3208 ();
 sg13g2_fill_2 FILLER_48_3212 ();
 sg13g2_decap_4 FILLER_48_3256 ();
 sg13g2_fill_2 FILLER_48_3260 ();
 sg13g2_fill_1 FILLER_48_3277 ();
 sg13g2_fill_2 FILLER_48_3282 ();
 sg13g2_fill_1 FILLER_48_3298 ();
 sg13g2_decap_8 FILLER_48_3312 ();
 sg13g2_decap_8 FILLER_48_3319 ();
 sg13g2_fill_2 FILLER_48_3326 ();
 sg13g2_fill_2 FILLER_48_3340 ();
 sg13g2_decap_4 FILLER_48_3347 ();
 sg13g2_fill_2 FILLER_48_3381 ();
 sg13g2_fill_1 FILLER_48_3383 ();
 sg13g2_fill_2 FILLER_48_3389 ();
 sg13g2_fill_2 FILLER_48_3412 ();
 sg13g2_decap_8 FILLER_48_3431 ();
 sg13g2_fill_2 FILLER_48_3438 ();
 sg13g2_fill_1 FILLER_48_3440 ();
 sg13g2_fill_1 FILLER_48_3458 ();
 sg13g2_fill_2 FILLER_48_3483 ();
 sg13g2_fill_1 FILLER_48_3485 ();
 sg13g2_decap_8 FILLER_48_3507 ();
 sg13g2_decap_8 FILLER_48_3526 ();
 sg13g2_decap_8 FILLER_48_3541 ();
 sg13g2_decap_4 FILLER_48_3575 ();
 sg13g2_fill_1 FILLER_48_3579 ();
 sg13g2_fill_1 FILLER_49_32 ();
 sg13g2_decap_8 FILLER_49_61 ();
 sg13g2_fill_2 FILLER_49_68 ();
 sg13g2_decap_8 FILLER_49_74 ();
 sg13g2_fill_1 FILLER_49_81 ();
 sg13g2_fill_2 FILLER_49_108 ();
 sg13g2_fill_1 FILLER_49_159 ();
 sg13g2_fill_2 FILLER_49_196 ();
 sg13g2_fill_1 FILLER_49_234 ();
 sg13g2_fill_2 FILLER_49_331 ();
 sg13g2_fill_1 FILLER_49_346 ();
 sg13g2_decap_4 FILLER_49_387 ();
 sg13g2_fill_1 FILLER_49_391 ();
 sg13g2_decap_4 FILLER_49_397 ();
 sg13g2_fill_2 FILLER_49_430 ();
 sg13g2_fill_1 FILLER_49_436 ();
 sg13g2_fill_2 FILLER_49_461 ();
 sg13g2_fill_1 FILLER_49_463 ();
 sg13g2_fill_1 FILLER_49_468 ();
 sg13g2_fill_2 FILLER_49_484 ();
 sg13g2_fill_1 FILLER_49_491 ();
 sg13g2_decap_8 FILLER_49_507 ();
 sg13g2_fill_1 FILLER_49_514 ();
 sg13g2_fill_1 FILLER_49_533 ();
 sg13g2_fill_1 FILLER_49_539 ();
 sg13g2_decap_4 FILLER_49_552 ();
 sg13g2_decap_8 FILLER_49_560 ();
 sg13g2_decap_8 FILLER_49_567 ();
 sg13g2_fill_2 FILLER_49_574 ();
 sg13g2_fill_2 FILLER_49_604 ();
 sg13g2_fill_1 FILLER_49_606 ();
 sg13g2_decap_4 FILLER_49_624 ();
 sg13g2_fill_2 FILLER_49_656 ();
 sg13g2_fill_2 FILLER_49_677 ();
 sg13g2_fill_1 FILLER_49_679 ();
 sg13g2_fill_2 FILLER_49_690 ();
 sg13g2_fill_2 FILLER_49_698 ();
 sg13g2_decap_4 FILLER_49_704 ();
 sg13g2_decap_8 FILLER_49_712 ();
 sg13g2_decap_8 FILLER_49_719 ();
 sg13g2_fill_2 FILLER_49_726 ();
 sg13g2_fill_1 FILLER_49_728 ();
 sg13g2_fill_1 FILLER_49_737 ();
 sg13g2_decap_4 FILLER_49_750 ();
 sg13g2_fill_2 FILLER_49_767 ();
 sg13g2_decap_8 FILLER_49_789 ();
 sg13g2_fill_2 FILLER_49_796 ();
 sg13g2_fill_2 FILLER_49_810 ();
 sg13g2_decap_4 FILLER_49_816 ();
 sg13g2_decap_4 FILLER_49_831 ();
 sg13g2_fill_1 FILLER_49_839 ();
 sg13g2_decap_8 FILLER_49_844 ();
 sg13g2_decap_4 FILLER_49_851 ();
 sg13g2_fill_1 FILLER_49_855 ();
 sg13g2_fill_2 FILLER_49_869 ();
 sg13g2_fill_1 FILLER_49_871 ();
 sg13g2_fill_2 FILLER_49_908 ();
 sg13g2_fill_1 FILLER_49_922 ();
 sg13g2_decap_8 FILLER_49_942 ();
 sg13g2_fill_2 FILLER_49_949 ();
 sg13g2_fill_1 FILLER_49_951 ();
 sg13g2_decap_4 FILLER_49_969 ();
 sg13g2_decap_8 FILLER_49_978 ();
 sg13g2_decap_8 FILLER_49_999 ();
 sg13g2_decap_8 FILLER_49_1022 ();
 sg13g2_decap_8 FILLER_49_1029 ();
 sg13g2_fill_1 FILLER_49_1045 ();
 sg13g2_fill_2 FILLER_49_1053 ();
 sg13g2_fill_1 FILLER_49_1055 ();
 sg13g2_fill_2 FILLER_49_1061 ();
 sg13g2_fill_2 FILLER_49_1072 ();
 sg13g2_fill_2 FILLER_49_1093 ();
 sg13g2_fill_1 FILLER_49_1109 ();
 sg13g2_decap_8 FILLER_49_1143 ();
 sg13g2_decap_4 FILLER_49_1150 ();
 sg13g2_fill_2 FILLER_49_1154 ();
 sg13g2_fill_2 FILLER_49_1192 ();
 sg13g2_decap_4 FILLER_49_1222 ();
 sg13g2_fill_2 FILLER_49_1226 ();
 sg13g2_fill_1 FILLER_49_1275 ();
 sg13g2_fill_2 FILLER_49_1284 ();
 sg13g2_fill_1 FILLER_49_1286 ();
 sg13g2_decap_8 FILLER_49_1292 ();
 sg13g2_decap_4 FILLER_49_1299 ();
 sg13g2_fill_1 FILLER_49_1307 ();
 sg13g2_fill_2 FILLER_49_1342 ();
 sg13g2_fill_1 FILLER_49_1344 ();
 sg13g2_fill_1 FILLER_49_1371 ();
 sg13g2_fill_2 FILLER_49_1413 ();
 sg13g2_decap_4 FILLER_49_1420 ();
 sg13g2_decap_8 FILLER_49_1437 ();
 sg13g2_fill_2 FILLER_49_1466 ();
 sg13g2_decap_4 FILLER_49_1474 ();
 sg13g2_fill_2 FILLER_49_1478 ();
 sg13g2_fill_2 FILLER_49_1591 ();
 sg13g2_fill_2 FILLER_49_1661 ();
 sg13g2_decap_8 FILLER_49_1703 ();
 sg13g2_fill_2 FILLER_49_1710 ();
 sg13g2_fill_2 FILLER_49_1753 ();
 sg13g2_fill_2 FILLER_49_1763 ();
 sg13g2_fill_1 FILLER_49_1773 ();
 sg13g2_decap_8 FILLER_49_1778 ();
 sg13g2_fill_1 FILLER_49_1785 ();
 sg13g2_fill_1 FILLER_49_1832 ();
 sg13g2_decap_8 FILLER_49_1842 ();
 sg13g2_decap_4 FILLER_49_1849 ();
 sg13g2_fill_2 FILLER_49_1966 ();
 sg13g2_fill_1 FILLER_49_1990 ();
 sg13g2_fill_2 FILLER_49_2056 ();
 sg13g2_fill_1 FILLER_49_2095 ();
 sg13g2_decap_4 FILLER_49_2109 ();
 sg13g2_decap_4 FILLER_49_2131 ();
 sg13g2_fill_2 FILLER_49_2180 ();
 sg13g2_fill_1 FILLER_49_2182 ();
 sg13g2_decap_8 FILLER_49_2193 ();
 sg13g2_fill_2 FILLER_49_2200 ();
 sg13g2_fill_1 FILLER_49_2202 ();
 sg13g2_fill_2 FILLER_49_2209 ();
 sg13g2_fill_1 FILLER_49_2211 ();
 sg13g2_fill_2 FILLER_49_2218 ();
 sg13g2_fill_2 FILLER_49_2252 ();
 sg13g2_fill_2 FILLER_49_2263 ();
 sg13g2_fill_1 FILLER_49_2265 ();
 sg13g2_fill_1 FILLER_49_2282 ();
 sg13g2_fill_1 FILLER_49_2291 ();
 sg13g2_fill_1 FILLER_49_2298 ();
 sg13g2_decap_8 FILLER_49_2307 ();
 sg13g2_decap_8 FILLER_49_2314 ();
 sg13g2_fill_2 FILLER_49_2321 ();
 sg13g2_decap_8 FILLER_49_2353 ();
 sg13g2_decap_4 FILLER_49_2360 ();
 sg13g2_fill_1 FILLER_49_2383 ();
 sg13g2_decap_4 FILLER_49_2409 ();
 sg13g2_fill_2 FILLER_49_2416 ();
 sg13g2_fill_1 FILLER_49_2435 ();
 sg13g2_fill_2 FILLER_49_2485 ();
 sg13g2_decap_4 FILLER_49_2499 ();
 sg13g2_decap_4 FILLER_49_2529 ();
 sg13g2_fill_1 FILLER_49_2533 ();
 sg13g2_decap_8 FILLER_49_2547 ();
 sg13g2_fill_2 FILLER_49_2565 ();
 sg13g2_fill_1 FILLER_49_2567 ();
 sg13g2_decap_4 FILLER_49_2583 ();
 sg13g2_fill_2 FILLER_49_2605 ();
 sg13g2_fill_1 FILLER_49_2607 ();
 sg13g2_fill_1 FILLER_49_2632 ();
 sg13g2_fill_2 FILLER_49_2646 ();
 sg13g2_fill_1 FILLER_49_2686 ();
 sg13g2_decap_4 FILLER_49_2711 ();
 sg13g2_fill_2 FILLER_49_2731 ();
 sg13g2_fill_1 FILLER_49_2733 ();
 sg13g2_fill_1 FILLER_49_2739 ();
 sg13g2_decap_4 FILLER_49_2790 ();
 sg13g2_fill_2 FILLER_49_2794 ();
 sg13g2_fill_1 FILLER_49_2813 ();
 sg13g2_decap_8 FILLER_49_2842 ();
 sg13g2_fill_2 FILLER_49_2849 ();
 sg13g2_fill_1 FILLER_49_2877 ();
 sg13g2_decap_4 FILLER_49_2891 ();
 sg13g2_fill_2 FILLER_49_2895 ();
 sg13g2_fill_2 FILLER_49_2910 ();
 sg13g2_fill_1 FILLER_49_2912 ();
 sg13g2_fill_1 FILLER_49_2926 ();
 sg13g2_decap_8 FILLER_49_2937 ();
 sg13g2_decap_4 FILLER_49_2965 ();
 sg13g2_fill_2 FILLER_49_2969 ();
 sg13g2_fill_2 FILLER_49_2980 ();
 sg13g2_decap_4 FILLER_49_3012 ();
 sg13g2_fill_1 FILLER_49_3039 ();
 sg13g2_fill_1 FILLER_49_3048 ();
 sg13g2_decap_8 FILLER_49_3066 ();
 sg13g2_fill_1 FILLER_49_3094 ();
 sg13g2_decap_8 FILLER_49_3116 ();
 sg13g2_decap_8 FILLER_49_3137 ();
 sg13g2_decap_8 FILLER_49_3144 ();
 sg13g2_fill_2 FILLER_49_3151 ();
 sg13g2_fill_2 FILLER_49_3186 ();
 sg13g2_fill_1 FILLER_49_3188 ();
 sg13g2_fill_1 FILLER_49_3220 ();
 sg13g2_fill_2 FILLER_49_3226 ();
 sg13g2_fill_1 FILLER_49_3228 ();
 sg13g2_fill_1 FILLER_49_3266 ();
 sg13g2_fill_1 FILLER_49_3275 ();
 sg13g2_fill_2 FILLER_49_3289 ();
 sg13g2_fill_1 FILLER_49_3291 ();
 sg13g2_fill_1 FILLER_49_3305 ();
 sg13g2_fill_2 FILLER_49_3311 ();
 sg13g2_fill_2 FILLER_49_3323 ();
 sg13g2_fill_1 FILLER_49_3325 ();
 sg13g2_fill_1 FILLER_49_3385 ();
 sg13g2_fill_2 FILLER_49_3438 ();
 sg13g2_fill_1 FILLER_49_3440 ();
 sg13g2_fill_2 FILLER_49_3445 ();
 sg13g2_fill_2 FILLER_49_3452 ();
 sg13g2_fill_1 FILLER_49_3463 ();
 sg13g2_fill_2 FILLER_49_3476 ();
 sg13g2_fill_1 FILLER_49_3478 ();
 sg13g2_decap_4 FILLER_49_3492 ();
 sg13g2_decap_4 FILLER_49_3500 ();
 sg13g2_fill_2 FILLER_49_3504 ();
 sg13g2_fill_1 FILLER_49_3514 ();
 sg13g2_fill_2 FILLER_49_3523 ();
 sg13g2_fill_1 FILLER_49_3525 ();
 sg13g2_fill_2 FILLER_49_3531 ();
 sg13g2_decap_4 FILLER_49_3537 ();
 sg13g2_fill_2 FILLER_49_3577 ();
 sg13g2_fill_1 FILLER_49_3579 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_fill_1 FILLER_50_30 ();
 sg13g2_fill_2 FILLER_50_44 ();
 sg13g2_fill_1 FILLER_50_46 ();
 sg13g2_fill_2 FILLER_50_52 ();
 sg13g2_fill_1 FILLER_50_54 ();
 sg13g2_decap_8 FILLER_50_94 ();
 sg13g2_fill_1 FILLER_50_101 ();
 sg13g2_fill_2 FILLER_50_109 ();
 sg13g2_fill_1 FILLER_50_111 ();
 sg13g2_fill_2 FILLER_50_148 ();
 sg13g2_fill_1 FILLER_50_150 ();
 sg13g2_fill_1 FILLER_50_164 ();
 sg13g2_fill_2 FILLER_50_197 ();
 sg13g2_fill_1 FILLER_50_199 ();
 sg13g2_fill_2 FILLER_50_220 ();
 sg13g2_fill_1 FILLER_50_277 ();
 sg13g2_fill_2 FILLER_50_292 ();
 sg13g2_fill_2 FILLER_50_429 ();
 sg13g2_fill_1 FILLER_50_461 ();
 sg13g2_decap_4 FILLER_50_482 ();
 sg13g2_fill_1 FILLER_50_505 ();
 sg13g2_decap_4 FILLER_50_519 ();
 sg13g2_fill_2 FILLER_50_523 ();
 sg13g2_fill_2 FILLER_50_533 ();
 sg13g2_fill_1 FILLER_50_548 ();
 sg13g2_fill_2 FILLER_50_557 ();
 sg13g2_fill_1 FILLER_50_559 ();
 sg13g2_decap_4 FILLER_50_569 ();
 sg13g2_fill_2 FILLER_50_573 ();
 sg13g2_fill_1 FILLER_50_585 ();
 sg13g2_fill_1 FILLER_50_603 ();
 sg13g2_decap_4 FILLER_50_629 ();
 sg13g2_fill_2 FILLER_50_637 ();
 sg13g2_fill_1 FILLER_50_639 ();
 sg13g2_fill_1 FILLER_50_680 ();
 sg13g2_fill_2 FILLER_50_690 ();
 sg13g2_decap_4 FILLER_50_733 ();
 sg13g2_fill_2 FILLER_50_754 ();
 sg13g2_fill_1 FILLER_50_756 ();
 sg13g2_fill_1 FILLER_50_762 ();
 sg13g2_fill_2 FILLER_50_794 ();
 sg13g2_fill_1 FILLER_50_810 ();
 sg13g2_decap_8 FILLER_50_866 ();
 sg13g2_decap_4 FILLER_50_873 ();
 sg13g2_fill_2 FILLER_50_877 ();
 sg13g2_fill_1 FILLER_50_892 ();
 sg13g2_fill_2 FILLER_50_904 ();
 sg13g2_decap_4 FILLER_50_947 ();
 sg13g2_fill_1 FILLER_50_951 ();
 sg13g2_fill_1 FILLER_50_963 ();
 sg13g2_decap_8 FILLER_50_976 ();
 sg13g2_fill_1 FILLER_50_992 ();
 sg13g2_fill_2 FILLER_50_1024 ();
 sg13g2_fill_1 FILLER_50_1026 ();
 sg13g2_fill_2 FILLER_50_1066 ();
 sg13g2_fill_2 FILLER_50_1111 ();
 sg13g2_fill_2 FILLER_50_1122 ();
 sg13g2_fill_1 FILLER_50_1124 ();
 sg13g2_fill_2 FILLER_50_1137 ();
 sg13g2_fill_1 FILLER_50_1139 ();
 sg13g2_decap_4 FILLER_50_1156 ();
 sg13g2_fill_2 FILLER_50_1165 ();
 sg13g2_fill_2 FILLER_50_1188 ();
 sg13g2_fill_1 FILLER_50_1198 ();
 sg13g2_decap_4 FILLER_50_1203 ();
 sg13g2_fill_2 FILLER_50_1207 ();
 sg13g2_fill_2 FILLER_50_1242 ();
 sg13g2_fill_1 FILLER_50_1244 ();
 sg13g2_decap_4 FILLER_50_1252 ();
 sg13g2_fill_1 FILLER_50_1260 ();
 sg13g2_fill_1 FILLER_50_1324 ();
 sg13g2_fill_1 FILLER_50_1356 ();
 sg13g2_fill_2 FILLER_50_1365 ();
 sg13g2_fill_1 FILLER_50_1367 ();
 sg13g2_fill_1 FILLER_50_1393 ();
 sg13g2_fill_2 FILLER_50_1421 ();
 sg13g2_fill_1 FILLER_50_1423 ();
 sg13g2_fill_1 FILLER_50_1450 ();
 sg13g2_fill_1 FILLER_50_1455 ();
 sg13g2_decap_4 FILLER_50_1469 ();
 sg13g2_fill_1 FILLER_50_1522 ();
 sg13g2_fill_1 FILLER_50_1529 ();
 sg13g2_fill_1 FILLER_50_1548 ();
 sg13g2_fill_2 FILLER_50_1567 ();
 sg13g2_fill_1 FILLER_50_1569 ();
 sg13g2_fill_1 FILLER_50_1579 ();
 sg13g2_fill_2 FILLER_50_1590 ();
 sg13g2_decap_4 FILLER_50_1611 ();
 sg13g2_fill_1 FILLER_50_1615 ();
 sg13g2_decap_8 FILLER_50_1702 ();
 sg13g2_decap_4 FILLER_50_1709 ();
 sg13g2_fill_1 FILLER_50_1713 ();
 sg13g2_decap_4 FILLER_50_1742 ();
 sg13g2_fill_1 FILLER_50_1746 ();
 sg13g2_fill_1 FILLER_50_1755 ();
 sg13g2_decap_8 FILLER_50_1783 ();
 sg13g2_decap_8 FILLER_50_1790 ();
 sg13g2_decap_4 FILLER_50_1815 ();
 sg13g2_decap_4 FILLER_50_1875 ();
 sg13g2_fill_2 FILLER_50_1879 ();
 sg13g2_fill_2 FILLER_50_1890 ();
 sg13g2_fill_1 FILLER_50_1892 ();
 sg13g2_fill_2 FILLER_50_1905 ();
 sg13g2_fill_2 FILLER_50_1992 ();
 sg13g2_decap_4 FILLER_50_2135 ();
 sg13g2_fill_1 FILLER_50_2139 ();
 sg13g2_fill_1 FILLER_50_2155 ();
 sg13g2_fill_2 FILLER_50_2169 ();
 sg13g2_fill_1 FILLER_50_2171 ();
 sg13g2_fill_1 FILLER_50_2180 ();
 sg13g2_decap_4 FILLER_50_2200 ();
 sg13g2_decap_4 FILLER_50_2213 ();
 sg13g2_fill_1 FILLER_50_2217 ();
 sg13g2_decap_4 FILLER_50_2241 ();
 sg13g2_decap_4 FILLER_50_2250 ();
 sg13g2_decap_4 FILLER_50_2292 ();
 sg13g2_fill_2 FILLER_50_2314 ();
 sg13g2_fill_1 FILLER_50_2316 ();
 sg13g2_fill_2 FILLER_50_2321 ();
 sg13g2_fill_1 FILLER_50_2323 ();
 sg13g2_decap_4 FILLER_50_2333 ();
 sg13g2_fill_2 FILLER_50_2337 ();
 sg13g2_fill_1 FILLER_50_2344 ();
 sg13g2_decap_8 FILLER_50_2358 ();
 sg13g2_decap_8 FILLER_50_2423 ();
 sg13g2_fill_2 FILLER_50_2430 ();
 sg13g2_fill_2 FILLER_50_2460 ();
 sg13g2_fill_1 FILLER_50_2462 ();
 sg13g2_fill_2 FILLER_50_2497 ();
 sg13g2_decap_8 FILLER_50_2509 ();
 sg13g2_decap_4 FILLER_50_2516 ();
 sg13g2_decap_4 FILLER_50_2529 ();
 sg13g2_fill_1 FILLER_50_2533 ();
 sg13g2_decap_4 FILLER_50_2539 ();
 sg13g2_fill_2 FILLER_50_2579 ();
 sg13g2_fill_1 FILLER_50_2581 ();
 sg13g2_fill_2 FILLER_50_2592 ();
 sg13g2_fill_1 FILLER_50_2594 ();
 sg13g2_fill_1 FILLER_50_2608 ();
 sg13g2_decap_8 FILLER_50_2614 ();
 sg13g2_decap_8 FILLER_50_2621 ();
 sg13g2_decap_8 FILLER_50_2628 ();
 sg13g2_decap_8 FILLER_50_2635 ();
 sg13g2_fill_2 FILLER_50_2642 ();
 sg13g2_decap_8 FILLER_50_2681 ();
 sg13g2_decap_4 FILLER_50_2688 ();
 sg13g2_fill_1 FILLER_50_2692 ();
 sg13g2_fill_1 FILLER_50_2766 ();
 sg13g2_fill_2 FILLER_50_2820 ();
 sg13g2_decap_4 FILLER_50_2844 ();
 sg13g2_fill_1 FILLER_50_2874 ();
 sg13g2_fill_2 FILLER_50_2891 ();
 sg13g2_decap_8 FILLER_50_2932 ();
 sg13g2_fill_2 FILLER_50_2939 ();
 sg13g2_decap_4 FILLER_50_2964 ();
 sg13g2_fill_2 FILLER_50_2993 ();
 sg13g2_fill_1 FILLER_50_2995 ();
 sg13g2_decap_8 FILLER_50_3005 ();
 sg13g2_decap_8 FILLER_50_3042 ();
 sg13g2_decap_4 FILLER_50_3049 ();
 sg13g2_fill_2 FILLER_50_3053 ();
 sg13g2_decap_8 FILLER_50_3068 ();
 sg13g2_fill_2 FILLER_50_3075 ();
 sg13g2_fill_1 FILLER_50_3077 ();
 sg13g2_fill_2 FILLER_50_3100 ();
 sg13g2_fill_1 FILLER_50_3102 ();
 sg13g2_fill_2 FILLER_50_3132 ();
 sg13g2_fill_1 FILLER_50_3134 ();
 sg13g2_decap_8 FILLER_50_3142 ();
 sg13g2_fill_2 FILLER_50_3149 ();
 sg13g2_fill_1 FILLER_50_3151 ();
 sg13g2_fill_2 FILLER_50_3170 ();
 sg13g2_fill_2 FILLER_50_3190 ();
 sg13g2_fill_2 FILLER_50_3197 ();
 sg13g2_fill_1 FILLER_50_3199 ();
 sg13g2_fill_1 FILLER_50_3209 ();
 sg13g2_fill_2 FILLER_50_3229 ();
 sg13g2_fill_1 FILLER_50_3235 ();
 sg13g2_decap_8 FILLER_50_3248 ();
 sg13g2_fill_2 FILLER_50_3255 ();
 sg13g2_fill_1 FILLER_50_3257 ();
 sg13g2_decap_8 FILLER_50_3279 ();
 sg13g2_decap_4 FILLER_50_3286 ();
 sg13g2_fill_1 FILLER_50_3290 ();
 sg13g2_fill_2 FILLER_50_3324 ();
 sg13g2_decap_8 FILLER_50_3349 ();
 sg13g2_fill_2 FILLER_50_3356 ();
 sg13g2_decap_4 FILLER_50_3363 ();
 sg13g2_decap_4 FILLER_50_3393 ();
 sg13g2_fill_2 FILLER_50_3397 ();
 sg13g2_decap_8 FILLER_50_3407 ();
 sg13g2_decap_4 FILLER_50_3431 ();
 sg13g2_fill_1 FILLER_50_3435 ();
 sg13g2_fill_1 FILLER_50_3464 ();
 sg13g2_fill_2 FILLER_50_3477 ();
 sg13g2_decap_8 FILLER_50_3492 ();
 sg13g2_fill_2 FILLER_50_3499 ();
 sg13g2_fill_1 FILLER_50_3501 ();
 sg13g2_decap_4 FILLER_50_3523 ();
 sg13g2_decap_4 FILLER_50_3575 ();
 sg13g2_fill_1 FILLER_50_3579 ();
 sg13g2_fill_1 FILLER_51_31 ();
 sg13g2_fill_1 FILLER_51_37 ();
 sg13g2_decap_4 FILLER_51_69 ();
 sg13g2_fill_2 FILLER_51_73 ();
 sg13g2_decap_8 FILLER_51_89 ();
 sg13g2_decap_4 FILLER_51_96 ();
 sg13g2_fill_1 FILLER_51_113 ();
 sg13g2_fill_2 FILLER_51_138 ();
 sg13g2_fill_1 FILLER_51_140 ();
 sg13g2_fill_2 FILLER_51_149 ();
 sg13g2_decap_4 FILLER_51_164 ();
 sg13g2_fill_2 FILLER_51_186 ();
 sg13g2_fill_1 FILLER_51_188 ();
 sg13g2_fill_1 FILLER_51_220 ();
 sg13g2_fill_2 FILLER_51_257 ();
 sg13g2_fill_1 FILLER_51_309 ();
 sg13g2_decap_4 FILLER_51_350 ();
 sg13g2_fill_2 FILLER_51_367 ();
 sg13g2_fill_1 FILLER_51_369 ();
 sg13g2_fill_2 FILLER_51_400 ();
 sg13g2_fill_1 FILLER_51_402 ();
 sg13g2_fill_2 FILLER_51_417 ();
 sg13g2_decap_4 FILLER_51_451 ();
 sg13g2_decap_8 FILLER_51_460 ();
 sg13g2_fill_2 FILLER_51_467 ();
 sg13g2_fill_1 FILLER_51_469 ();
 sg13g2_decap_8 FILLER_51_484 ();
 sg13g2_fill_2 FILLER_51_500 ();
 sg13g2_decap_8 FILLER_51_507 ();
 sg13g2_fill_1 FILLER_51_514 ();
 sg13g2_fill_2 FILLER_51_543 ();
 sg13g2_decap_8 FILLER_51_549 ();
 sg13g2_fill_2 FILLER_51_556 ();
 sg13g2_fill_2 FILLER_51_562 ();
 sg13g2_fill_1 FILLER_51_564 ();
 sg13g2_decap_4 FILLER_51_593 ();
 sg13g2_fill_1 FILLER_51_597 ();
 sg13g2_fill_2 FILLER_51_619 ();
 sg13g2_fill_1 FILLER_51_621 ();
 sg13g2_decap_8 FILLER_51_632 ();
 sg13g2_fill_2 FILLER_51_639 ();
 sg13g2_fill_1 FILLER_51_641 ();
 sg13g2_fill_1 FILLER_51_667 ();
 sg13g2_fill_2 FILLER_51_675 ();
 sg13g2_fill_1 FILLER_51_677 ();
 sg13g2_decap_4 FILLER_51_689 ();
 sg13g2_fill_2 FILLER_51_693 ();
 sg13g2_decap_8 FILLER_51_700 ();
 sg13g2_fill_1 FILLER_51_707 ();
 sg13g2_decap_8 FILLER_51_726 ();
 sg13g2_decap_8 FILLER_51_753 ();
 sg13g2_fill_2 FILLER_51_760 ();
 sg13g2_fill_1 FILLER_51_762 ();
 sg13g2_decap_4 FILLER_51_793 ();
 sg13g2_fill_1 FILLER_51_797 ();
 sg13g2_fill_1 FILLER_51_810 ();
 sg13g2_decap_8 FILLER_51_815 ();
 sg13g2_decap_8 FILLER_51_830 ();
 sg13g2_decap_4 FILLER_51_837 ();
 sg13g2_fill_1 FILLER_51_841 ();
 sg13g2_fill_2 FILLER_51_848 ();
 sg13g2_fill_2 FILLER_51_858 ();
 sg13g2_decap_8 FILLER_51_872 ();
 sg13g2_fill_1 FILLER_51_879 ();
 sg13g2_fill_2 FILLER_51_902 ();
 sg13g2_fill_2 FILLER_51_909 ();
 sg13g2_decap_8 FILLER_51_915 ();
 sg13g2_decap_8 FILLER_51_945 ();
 sg13g2_fill_1 FILLER_51_952 ();
 sg13g2_decap_8 FILLER_51_969 ();
 sg13g2_fill_1 FILLER_51_976 ();
 sg13g2_fill_2 FILLER_51_995 ();
 sg13g2_fill_2 FILLER_51_1012 ();
 sg13g2_fill_1 FILLER_51_1014 ();
 sg13g2_fill_1 FILLER_51_1060 ();
 sg13g2_decap_8 FILLER_51_1069 ();
 sg13g2_decap_4 FILLER_51_1076 ();
 sg13g2_fill_2 FILLER_51_1080 ();
 sg13g2_fill_2 FILLER_51_1086 ();
 sg13g2_fill_1 FILLER_51_1088 ();
 sg13g2_decap_8 FILLER_51_1097 ();
 sg13g2_fill_2 FILLER_51_1104 ();
 sg13g2_fill_1 FILLER_51_1124 ();
 sg13g2_decap_8 FILLER_51_1133 ();
 sg13g2_fill_1 FILLER_51_1140 ();
 sg13g2_fill_2 FILLER_51_1154 ();
 sg13g2_fill_1 FILLER_51_1172 ();
 sg13g2_fill_1 FILLER_51_1183 ();
 sg13g2_decap_8 FILLER_51_1200 ();
 sg13g2_decap_4 FILLER_51_1229 ();
 sg13g2_fill_1 FILLER_51_1233 ();
 sg13g2_fill_2 FILLER_51_1271 ();
 sg13g2_fill_2 FILLER_51_1278 ();
 sg13g2_fill_1 FILLER_51_1308 ();
 sg13g2_fill_1 FILLER_51_1354 ();
 sg13g2_fill_2 FILLER_51_1400 ();
 sg13g2_fill_1 FILLER_51_1402 ();
 sg13g2_fill_1 FILLER_51_1419 ();
 sg13g2_decap_4 FILLER_51_1460 ();
 sg13g2_fill_2 FILLER_51_1464 ();
 sg13g2_decap_4 FILLER_51_1474 ();
 sg13g2_fill_1 FILLER_51_1478 ();
 sg13g2_fill_2 FILLER_51_1487 ();
 sg13g2_fill_2 FILLER_51_1497 ();
 sg13g2_fill_2 FILLER_51_1504 ();
 sg13g2_fill_1 FILLER_51_1506 ();
 sg13g2_decap_4 FILLER_51_1532 ();
 sg13g2_fill_2 FILLER_51_1536 ();
 sg13g2_fill_2 FILLER_51_1579 ();
 sg13g2_fill_2 FILLER_51_1589 ();
 sg13g2_fill_2 FILLER_51_1605 ();
 sg13g2_fill_2 FILLER_51_1638 ();
 sg13g2_fill_2 FILLER_51_1653 ();
 sg13g2_fill_1 FILLER_51_1655 ();
 sg13g2_fill_2 FILLER_51_1673 ();
 sg13g2_fill_1 FILLER_51_1675 ();
 sg13g2_fill_2 FILLER_51_1712 ();
 sg13g2_fill_1 FILLER_51_1768 ();
 sg13g2_decap_4 FILLER_51_1819 ();
 sg13g2_fill_2 FILLER_51_1862 ();
 sg13g2_decap_8 FILLER_51_1872 ();
 sg13g2_fill_2 FILLER_51_1879 ();
 sg13g2_fill_1 FILLER_51_1881 ();
 sg13g2_fill_1 FILLER_51_1915 ();
 sg13g2_fill_1 FILLER_51_1935 ();
 sg13g2_fill_2 FILLER_51_2053 ();
 sg13g2_decap_8 FILLER_51_2108 ();
 sg13g2_fill_1 FILLER_51_2131 ();
 sg13g2_fill_1 FILLER_51_2150 ();
 sg13g2_decap_4 FILLER_51_2160 ();
 sg13g2_decap_8 FILLER_51_2180 ();
 sg13g2_fill_2 FILLER_51_2187 ();
 sg13g2_fill_2 FILLER_51_2217 ();
 sg13g2_fill_1 FILLER_51_2219 ();
 sg13g2_fill_2 FILLER_51_2287 ();
 sg13g2_fill_1 FILLER_51_2289 ();
 sg13g2_fill_1 FILLER_51_2315 ();
 sg13g2_fill_1 FILLER_51_2349 ();
 sg13g2_fill_2 FILLER_51_2356 ();
 sg13g2_decap_8 FILLER_51_2371 ();
 sg13g2_decap_8 FILLER_51_2378 ();
 sg13g2_decap_4 FILLER_51_2385 ();
 sg13g2_fill_2 FILLER_51_2389 ();
 sg13g2_fill_2 FILLER_51_2404 ();
 sg13g2_fill_1 FILLER_51_2406 ();
 sg13g2_decap_8 FILLER_51_2431 ();
 sg13g2_decap_4 FILLER_51_2438 ();
 sg13g2_fill_2 FILLER_51_2442 ();
 sg13g2_decap_4 FILLER_51_2457 ();
 sg13g2_fill_1 FILLER_51_2461 ();
 sg13g2_decap_4 FILLER_51_2469 ();
 sg13g2_decap_8 FILLER_51_2501 ();
 sg13g2_fill_2 FILLER_51_2508 ();
 sg13g2_fill_1 FILLER_51_2510 ();
 sg13g2_fill_2 FILLER_51_2540 ();
 sg13g2_fill_1 FILLER_51_2542 ();
 sg13g2_fill_2 FILLER_51_2556 ();
 sg13g2_fill_1 FILLER_51_2558 ();
 sg13g2_fill_1 FILLER_51_2564 ();
 sg13g2_fill_2 FILLER_51_2593 ();
 sg13g2_fill_1 FILLER_51_2612 ();
 sg13g2_fill_2 FILLER_51_2627 ();
 sg13g2_fill_1 FILLER_51_2629 ();
 sg13g2_fill_1 FILLER_51_2643 ();
 sg13g2_fill_2 FILLER_51_2657 ();
 sg13g2_fill_2 FILLER_51_2705 ();
 sg13g2_fill_1 FILLER_51_2707 ();
 sg13g2_decap_4 FILLER_51_2730 ();
 sg13g2_fill_2 FILLER_51_2808 ();
 sg13g2_fill_1 FILLER_51_2810 ();
 sg13g2_fill_2 FILLER_51_2815 ();
 sg13g2_fill_2 FILLER_51_2822 ();
 sg13g2_fill_1 FILLER_51_2875 ();
 sg13g2_fill_2 FILLER_51_2890 ();
 sg13g2_fill_1 FILLER_51_2892 ();
 sg13g2_fill_1 FILLER_51_2902 ();
 sg13g2_fill_2 FILLER_51_2909 ();
 sg13g2_fill_2 FILLER_51_2917 ();
 sg13g2_decap_4 FILLER_51_2933 ();
 sg13g2_decap_4 FILLER_51_2970 ();
 sg13g2_fill_2 FILLER_51_2992 ();
 sg13g2_fill_2 FILLER_51_3016 ();
 sg13g2_fill_1 FILLER_51_3018 ();
 sg13g2_fill_1 FILLER_51_3043 ();
 sg13g2_decap_4 FILLER_51_3060 ();
 sg13g2_fill_1 FILLER_51_3073 ();
 sg13g2_fill_2 FILLER_51_3122 ();
 sg13g2_decap_4 FILLER_51_3137 ();
 sg13g2_fill_1 FILLER_51_3141 ();
 sg13g2_decap_4 FILLER_51_3222 ();
 sg13g2_fill_2 FILLER_51_3226 ();
 sg13g2_decap_4 FILLER_51_3254 ();
 sg13g2_fill_2 FILLER_51_3263 ();
 sg13g2_fill_1 FILLER_51_3265 ();
 sg13g2_decap_4 FILLER_51_3281 ();
 sg13g2_fill_1 FILLER_51_3285 ();
 sg13g2_decap_4 FILLER_51_3313 ();
 sg13g2_fill_1 FILLER_51_3362 ();
 sg13g2_decap_8 FILLER_51_3385 ();
 sg13g2_decap_4 FILLER_51_3392 ();
 sg13g2_fill_2 FILLER_51_3435 ();
 sg13g2_decap_8 FILLER_51_3470 ();
 sg13g2_decap_4 FILLER_51_3477 ();
 sg13g2_fill_1 FILLER_51_3481 ();
 sg13g2_decap_8 FILLER_51_3500 ();
 sg13g2_decap_4 FILLER_51_3521 ();
 sg13g2_fill_1 FILLER_51_3525 ();
 sg13g2_fill_1 FILLER_51_3544 ();
 sg13g2_fill_2 FILLER_51_3550 ();
 sg13g2_fill_2 FILLER_52_51 ();
 sg13g2_fill_1 FILLER_52_53 ();
 sg13g2_fill_2 FILLER_52_64 ();
 sg13g2_fill_1 FILLER_52_66 ();
 sg13g2_fill_2 FILLER_52_79 ();
 sg13g2_fill_1 FILLER_52_81 ();
 sg13g2_decap_8 FILLER_52_90 ();
 sg13g2_fill_2 FILLER_52_97 ();
 sg13g2_fill_2 FILLER_52_115 ();
 sg13g2_fill_2 FILLER_52_122 ();
 sg13g2_fill_1 FILLER_52_132 ();
 sg13g2_fill_1 FILLER_52_254 ();
 sg13g2_fill_2 FILLER_52_442 ();
 sg13g2_decap_4 FILLER_52_456 ();
 sg13g2_fill_2 FILLER_52_460 ();
 sg13g2_decap_4 FILLER_52_483 ();
 sg13g2_fill_1 FILLER_52_515 ();
 sg13g2_decap_4 FILLER_52_533 ();
 sg13g2_fill_1 FILLER_52_537 ();
 sg13g2_fill_2 FILLER_52_547 ();
 sg13g2_fill_1 FILLER_52_549 ();
 sg13g2_fill_1 FILLER_52_563 ();
 sg13g2_fill_1 FILLER_52_569 ();
 sg13g2_fill_1 FILLER_52_597 ();
 sg13g2_fill_1 FILLER_52_620 ();
 sg13g2_decap_8 FILLER_52_631 ();
 sg13g2_fill_1 FILLER_52_638 ();
 sg13g2_fill_2 FILLER_52_657 ();
 sg13g2_fill_2 FILLER_52_671 ();
 sg13g2_fill_1 FILLER_52_673 ();
 sg13g2_fill_2 FILLER_52_696 ();
 sg13g2_fill_2 FILLER_52_713 ();
 sg13g2_fill_2 FILLER_52_723 ();
 sg13g2_decap_8 FILLER_52_749 ();
 sg13g2_decap_8 FILLER_52_756 ();
 sg13g2_decap_4 FILLER_52_763 ();
 sg13g2_decap_4 FILLER_52_785 ();
 sg13g2_fill_1 FILLER_52_797 ();
 sg13g2_fill_2 FILLER_52_806 ();
 sg13g2_fill_1 FILLER_52_808 ();
 sg13g2_fill_2 FILLER_52_814 ();
 sg13g2_fill_1 FILLER_52_816 ();
 sg13g2_decap_8 FILLER_52_833 ();
 sg13g2_fill_2 FILLER_52_850 ();
 sg13g2_decap_4 FILLER_52_873 ();
 sg13g2_fill_2 FILLER_52_877 ();
 sg13g2_fill_2 FILLER_52_896 ();
 sg13g2_fill_1 FILLER_52_898 ();
 sg13g2_decap_4 FILLER_52_904 ();
 sg13g2_fill_1 FILLER_52_908 ();
 sg13g2_fill_2 FILLER_52_923 ();
 sg13g2_fill_1 FILLER_52_925 ();
 sg13g2_fill_2 FILLER_52_931 ();
 sg13g2_fill_1 FILLER_52_938 ();
 sg13g2_fill_2 FILLER_52_952 ();
 sg13g2_decap_4 FILLER_52_1007 ();
 sg13g2_decap_4 FILLER_52_1024 ();
 sg13g2_fill_2 FILLER_52_1028 ();
 sg13g2_fill_2 FILLER_52_1039 ();
 sg13g2_fill_2 FILLER_52_1050 ();
 sg13g2_fill_2 FILLER_52_1057 ();
 sg13g2_decap_8 FILLER_52_1073 ();
 sg13g2_fill_2 FILLER_52_1080 ();
 sg13g2_fill_1 FILLER_52_1082 ();
 sg13g2_fill_2 FILLER_52_1091 ();
 sg13g2_decap_8 FILLER_52_1102 ();
 sg13g2_fill_1 FILLER_52_1109 ();
 sg13g2_decap_4 FILLER_52_1128 ();
 sg13g2_fill_2 FILLER_52_1132 ();
 sg13g2_fill_2 FILLER_52_1141 ();
 sg13g2_fill_1 FILLER_52_1143 ();
 sg13g2_fill_2 FILLER_52_1157 ();
 sg13g2_fill_1 FILLER_52_1159 ();
 sg13g2_decap_4 FILLER_52_1165 ();
 sg13g2_fill_2 FILLER_52_1169 ();
 sg13g2_fill_1 FILLER_52_1182 ();
 sg13g2_decap_4 FILLER_52_1204 ();
 sg13g2_fill_2 FILLER_52_1236 ();
 sg13g2_decap_4 FILLER_52_1259 ();
 sg13g2_fill_1 FILLER_52_1263 ();
 sg13g2_decap_8 FILLER_52_1295 ();
 sg13g2_fill_2 FILLER_52_1325 ();
 sg13g2_fill_1 FILLER_52_1327 ();
 sg13g2_fill_2 FILLER_52_1373 ();
 sg13g2_fill_1 FILLER_52_1391 ();
 sg13g2_decap_8 FILLER_52_1443 ();
 sg13g2_decap_8 FILLER_52_1478 ();
 sg13g2_decap_4 FILLER_52_1485 ();
 sg13g2_fill_2 FILLER_52_1517 ();
 sg13g2_fill_1 FILLER_52_1519 ();
 sg13g2_fill_2 FILLER_52_1533 ();
 sg13g2_fill_1 FILLER_52_1535 ();
 sg13g2_decap_8 FILLER_52_1544 ();
 sg13g2_decap_8 FILLER_52_1551 ();
 sg13g2_decap_8 FILLER_52_1558 ();
 sg13g2_decap_8 FILLER_52_1565 ();
 sg13g2_decap_4 FILLER_52_1572 ();
 sg13g2_fill_1 FILLER_52_1576 ();
 sg13g2_decap_8 FILLER_52_1590 ();
 sg13g2_fill_2 FILLER_52_1597 ();
 sg13g2_fill_1 FILLER_52_1599 ();
 sg13g2_fill_2 FILLER_52_1614 ();
 sg13g2_fill_1 FILLER_52_1616 ();
 sg13g2_decap_4 FILLER_52_1620 ();
 sg13g2_fill_1 FILLER_52_1624 ();
 sg13g2_fill_2 FILLER_52_1638 ();
 sg13g2_fill_1 FILLER_52_1640 ();
 sg13g2_fill_2 FILLER_52_1658 ();
 sg13g2_decap_8 FILLER_52_1666 ();
 sg13g2_decap_8 FILLER_52_1673 ();
 sg13g2_fill_1 FILLER_52_1742 ();
 sg13g2_fill_1 FILLER_52_1751 ();
 sg13g2_fill_2 FILLER_52_1789 ();
 sg13g2_fill_1 FILLER_52_1791 ();
 sg13g2_fill_1 FILLER_52_1855 ();
 sg13g2_fill_2 FILLER_52_1884 ();
 sg13g2_fill_1 FILLER_52_1891 ();
 sg13g2_fill_1 FILLER_52_1916 ();
 sg13g2_fill_2 FILLER_52_1954 ();
 sg13g2_fill_1 FILLER_52_1956 ();
 sg13g2_fill_2 FILLER_52_1985 ();
 sg13g2_fill_1 FILLER_52_2028 ();
 sg13g2_fill_1 FILLER_52_2064 ();
 sg13g2_fill_2 FILLER_52_2074 ();
 sg13g2_fill_1 FILLER_52_2076 ();
 sg13g2_fill_2 FILLER_52_2098 ();
 sg13g2_decap_4 FILLER_52_2113 ();
 sg13g2_fill_2 FILLER_52_2142 ();
 sg13g2_fill_2 FILLER_52_2170 ();
 sg13g2_fill_2 FILLER_52_2181 ();
 sg13g2_decap_8 FILLER_52_2193 ();
 sg13g2_fill_2 FILLER_52_2233 ();
 sg13g2_decap_4 FILLER_52_2257 ();
 sg13g2_fill_2 FILLER_52_2269 ();
 sg13g2_fill_1 FILLER_52_2271 ();
 sg13g2_decap_4 FILLER_52_2277 ();
 sg13g2_decap_4 FILLER_52_2305 ();
 sg13g2_fill_1 FILLER_52_2309 ();
 sg13g2_fill_1 FILLER_52_2330 ();
 sg13g2_fill_1 FILLER_52_2344 ();
 sg13g2_fill_1 FILLER_52_2431 ();
 sg13g2_fill_2 FILLER_52_2454 ();
 sg13g2_fill_1 FILLER_52_2456 ();
 sg13g2_fill_2 FILLER_52_2477 ();
 sg13g2_fill_1 FILLER_52_2491 ();
 sg13g2_fill_2 FILLER_52_2532 ();
 sg13g2_fill_1 FILLER_52_2534 ();
 sg13g2_fill_1 FILLER_52_2557 ();
 sg13g2_decap_4 FILLER_52_2586 ();
 sg13g2_fill_2 FILLER_52_2590 ();
 sg13g2_decap_4 FILLER_52_2618 ();
 sg13g2_fill_2 FILLER_52_2622 ();
 sg13g2_fill_1 FILLER_52_2652 ();
 sg13g2_decap_4 FILLER_52_2690 ();
 sg13g2_fill_2 FILLER_52_2720 ();
 sg13g2_fill_1 FILLER_52_2722 ();
 sg13g2_fill_1 FILLER_52_2759 ();
 sg13g2_fill_2 FILLER_52_2769 ();
 sg13g2_fill_1 FILLER_52_2785 ();
 sg13g2_fill_1 FILLER_52_2795 ();
 sg13g2_fill_2 FILLER_52_2846 ();
 sg13g2_fill_1 FILLER_52_2848 ();
 sg13g2_fill_2 FILLER_52_2867 ();
 sg13g2_fill_1 FILLER_52_2877 ();
 sg13g2_decap_8 FILLER_52_2894 ();
 sg13g2_fill_2 FILLER_52_2915 ();
 sg13g2_decap_8 FILLER_52_2934 ();
 sg13g2_fill_2 FILLER_52_2941 ();
 sg13g2_fill_1 FILLER_52_2943 ();
 sg13g2_fill_1 FILLER_52_2997 ();
 sg13g2_decap_4 FILLER_52_3005 ();
 sg13g2_fill_1 FILLER_52_3009 ();
 sg13g2_fill_1 FILLER_52_3042 ();
 sg13g2_fill_2 FILLER_52_3095 ();
 sg13g2_decap_4 FILLER_52_3103 ();
 sg13g2_fill_2 FILLER_52_3107 ();
 sg13g2_fill_2 FILLER_52_3127 ();
 sg13g2_decap_8 FILLER_52_3138 ();
 sg13g2_decap_4 FILLER_52_3145 ();
 sg13g2_fill_1 FILLER_52_3178 ();
 sg13g2_fill_1 FILLER_52_3185 ();
 sg13g2_fill_2 FILLER_52_3195 ();
 sg13g2_fill_1 FILLER_52_3207 ();
 sg13g2_fill_2 FILLER_52_3241 ();
 sg13g2_fill_2 FILLER_52_3259 ();
 sg13g2_fill_1 FILLER_52_3261 ();
 sg13g2_decap_4 FILLER_52_3283 ();
 sg13g2_fill_2 FILLER_52_3287 ();
 sg13g2_fill_1 FILLER_52_3300 ();
 sg13g2_decap_4 FILLER_52_3308 ();
 sg13g2_fill_1 FILLER_52_3312 ();
 sg13g2_decap_4 FILLER_52_3318 ();
 sg13g2_fill_1 FILLER_52_3322 ();
 sg13g2_fill_2 FILLER_52_3335 ();
 sg13g2_decap_8 FILLER_52_3348 ();
 sg13g2_decap_4 FILLER_52_3355 ();
 sg13g2_fill_1 FILLER_52_3359 ();
 sg13g2_decap_8 FILLER_52_3379 ();
 sg13g2_fill_2 FILLER_52_3386 ();
 sg13g2_decap_8 FILLER_52_3392 ();
 sg13g2_fill_2 FILLER_52_3399 ();
 sg13g2_decap_4 FILLER_52_3415 ();
 sg13g2_fill_2 FILLER_52_3428 ();
 sg13g2_fill_1 FILLER_52_3430 ();
 sg13g2_fill_1 FILLER_52_3444 ();
 sg13g2_fill_2 FILLER_52_3449 ();
 sg13g2_fill_2 FILLER_52_3475 ();
 sg13g2_decap_8 FILLER_52_3502 ();
 sg13g2_fill_2 FILLER_52_3509 ();
 sg13g2_decap_4 FILLER_52_3542 ();
 sg13g2_fill_1 FILLER_52_3546 ();
 sg13g2_decap_8 FILLER_52_3572 ();
 sg13g2_fill_1 FILLER_52_3579 ();
 sg13g2_decap_4 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_4 ();
 sg13g2_fill_1 FILLER_53_38 ();
 sg13g2_fill_1 FILLER_53_43 ();
 sg13g2_fill_2 FILLER_53_57 ();
 sg13g2_decap_4 FILLER_53_83 ();
 sg13g2_fill_1 FILLER_53_87 ();
 sg13g2_fill_1 FILLER_53_129 ();
 sg13g2_fill_1 FILLER_53_148 ();
 sg13g2_fill_2 FILLER_53_158 ();
 sg13g2_fill_1 FILLER_53_160 ();
 sg13g2_fill_1 FILLER_53_174 ();
 sg13g2_fill_2 FILLER_53_189 ();
 sg13g2_fill_1 FILLER_53_219 ();
 sg13g2_fill_1 FILLER_53_273 ();
 sg13g2_fill_1 FILLER_53_290 ();
 sg13g2_decap_4 FILLER_53_342 ();
 sg13g2_fill_1 FILLER_53_390 ();
 sg13g2_fill_2 FILLER_53_399 ();
 sg13g2_decap_8 FILLER_53_415 ();
 sg13g2_decap_8 FILLER_53_422 ();
 sg13g2_fill_2 FILLER_53_429 ();
 sg13g2_fill_1 FILLER_53_431 ();
 sg13g2_fill_2 FILLER_53_452 ();
 sg13g2_fill_1 FILLER_53_454 ();
 sg13g2_fill_2 FILLER_53_462 ();
 sg13g2_fill_1 FILLER_53_464 ();
 sg13g2_fill_2 FILLER_53_480 ();
 sg13g2_fill_1 FILLER_53_491 ();
 sg13g2_decap_8 FILLER_53_503 ();
 sg13g2_decap_4 FILLER_53_510 ();
 sg13g2_fill_1 FILLER_53_514 ();
 sg13g2_decap_8 FILLER_53_519 ();
 sg13g2_fill_2 FILLER_53_526 ();
 sg13g2_fill_1 FILLER_53_528 ();
 sg13g2_fill_2 FILLER_53_571 ();
 sg13g2_fill_1 FILLER_53_573 ();
 sg13g2_fill_2 FILLER_53_583 ();
 sg13g2_fill_1 FILLER_53_585 ();
 sg13g2_decap_8 FILLER_53_591 ();
 sg13g2_fill_2 FILLER_53_598 ();
 sg13g2_decap_8 FILLER_53_627 ();
 sg13g2_fill_1 FILLER_53_647 ();
 sg13g2_fill_2 FILLER_53_655 ();
 sg13g2_fill_2 FILLER_53_667 ();
 sg13g2_fill_2 FILLER_53_679 ();
 sg13g2_decap_8 FILLER_53_691 ();
 sg13g2_decap_4 FILLER_53_731 ();
 sg13g2_fill_1 FILLER_53_735 ();
 sg13g2_fill_1 FILLER_53_751 ();
 sg13g2_fill_2 FILLER_53_790 ();
 sg13g2_fill_2 FILLER_53_802 ();
 sg13g2_decap_4 FILLER_53_835 ();
 sg13g2_fill_2 FILLER_53_839 ();
 sg13g2_decap_4 FILLER_53_875 ();
 sg13g2_fill_1 FILLER_53_879 ();
 sg13g2_decap_4 FILLER_53_902 ();
 sg13g2_fill_2 FILLER_53_906 ();
 sg13g2_decap_8 FILLER_53_920 ();
 sg13g2_decap_8 FILLER_53_944 ();
 sg13g2_decap_8 FILLER_53_951 ();
 sg13g2_fill_1 FILLER_53_958 ();
 sg13g2_decap_8 FILLER_53_972 ();
 sg13g2_decap_8 FILLER_53_979 ();
 sg13g2_decap_4 FILLER_53_1024 ();
 sg13g2_decap_4 FILLER_53_1054 ();
 sg13g2_fill_1 FILLER_53_1058 ();
 sg13g2_fill_2 FILLER_53_1063 ();
 sg13g2_decap_4 FILLER_53_1070 ();
 sg13g2_fill_1 FILLER_53_1074 ();
 sg13g2_fill_1 FILLER_53_1088 ();
 sg13g2_fill_2 FILLER_53_1130 ();
 sg13g2_fill_2 FILLER_53_1144 ();
 sg13g2_decap_8 FILLER_53_1204 ();
 sg13g2_decap_8 FILLER_53_1235 ();
 sg13g2_decap_8 FILLER_53_1251 ();
 sg13g2_decap_4 FILLER_53_1258 ();
 sg13g2_fill_1 FILLER_53_1262 ();
 sg13g2_decap_4 FILLER_53_1295 ();
 sg13g2_fill_2 FILLER_53_1299 ();
 sg13g2_fill_1 FILLER_53_1342 ();
 sg13g2_fill_2 FILLER_53_1370 ();
 sg13g2_fill_1 FILLER_53_1400 ();
 sg13g2_fill_1 FILLER_53_1412 ();
 sg13g2_fill_1 FILLER_53_1434 ();
 sg13g2_fill_2 FILLER_53_1440 ();
 sg13g2_fill_1 FILLER_53_1442 ();
 sg13g2_fill_1 FILLER_53_1446 ();
 sg13g2_fill_2 FILLER_53_1461 ();
 sg13g2_decap_8 FILLER_53_1477 ();
 sg13g2_fill_1 FILLER_53_1492 ();
 sg13g2_fill_2 FILLER_53_1517 ();
 sg13g2_decap_8 FILLER_53_1544 ();
 sg13g2_fill_2 FILLER_53_1551 ();
 sg13g2_decap_8 FILLER_53_1585 ();
 sg13g2_fill_2 FILLER_53_1592 ();
 sg13g2_fill_2 FILLER_53_1620 ();
 sg13g2_fill_1 FILLER_53_1622 ();
 sg13g2_decap_4 FILLER_53_1629 ();
 sg13g2_fill_2 FILLER_53_1659 ();
 sg13g2_fill_1 FILLER_53_1661 ();
 sg13g2_fill_1 FILLER_53_1688 ();
 sg13g2_fill_2 FILLER_53_1711 ();
 sg13g2_fill_1 FILLER_53_1713 ();
 sg13g2_fill_2 FILLER_53_1731 ();
 sg13g2_fill_1 FILLER_53_1733 ();
 sg13g2_fill_2 FILLER_53_1744 ();
 sg13g2_fill_1 FILLER_53_1746 ();
 sg13g2_decap_8 FILLER_53_1750 ();
 sg13g2_fill_2 FILLER_53_1767 ();
 sg13g2_fill_1 FILLER_53_1797 ();
 sg13g2_fill_2 FILLER_53_1835 ();
 sg13g2_fill_1 FILLER_53_1837 ();
 sg13g2_fill_1 FILLER_53_1912 ();
 sg13g2_fill_2 FILLER_53_1990 ();
 sg13g2_fill_2 FILLER_53_2038 ();
 sg13g2_fill_1 FILLER_53_2080 ();
 sg13g2_fill_2 FILLER_53_2146 ();
 sg13g2_fill_2 FILLER_53_2174 ();
 sg13g2_fill_1 FILLER_53_2176 ();
 sg13g2_decap_4 FILLER_53_2202 ();
 sg13g2_fill_2 FILLER_53_2266 ();
 sg13g2_decap_4 FILLER_53_2293 ();
 sg13g2_fill_2 FILLER_53_2297 ();
 sg13g2_fill_2 FILLER_53_2312 ();
 sg13g2_fill_1 FILLER_53_2314 ();
 sg13g2_decap_8 FILLER_53_2389 ();
 sg13g2_fill_1 FILLER_53_2396 ();
 sg13g2_fill_2 FILLER_53_2425 ();
 sg13g2_fill_2 FILLER_53_2455 ();
 sg13g2_fill_1 FILLER_53_2457 ();
 sg13g2_fill_1 FILLER_53_2473 ();
 sg13g2_fill_2 FILLER_53_2499 ();
 sg13g2_fill_2 FILLER_53_2537 ();
 sg13g2_fill_1 FILLER_53_2546 ();
 sg13g2_fill_2 FILLER_53_2585 ();
 sg13g2_fill_2 FILLER_53_2645 ();
 sg13g2_fill_2 FILLER_53_2697 ();
 sg13g2_fill_1 FILLER_53_2699 ();
 sg13g2_fill_2 FILLER_53_2705 ();
 sg13g2_fill_2 FILLER_53_2712 ();
 sg13g2_fill_1 FILLER_53_2714 ();
 sg13g2_fill_2 FILLER_53_2734 ();
 sg13g2_fill_1 FILLER_53_2736 ();
 sg13g2_decap_8 FILLER_53_2779 ();
 sg13g2_fill_1 FILLER_53_2786 ();
 sg13g2_fill_1 FILLER_53_2814 ();
 sg13g2_decap_4 FILLER_53_2828 ();
 sg13g2_fill_2 FILLER_53_2832 ();
 sg13g2_decap_4 FILLER_53_2847 ();
 sg13g2_fill_2 FILLER_53_2865 ();
 sg13g2_fill_1 FILLER_53_2867 ();
 sg13g2_fill_2 FILLER_53_2875 ();
 sg13g2_fill_1 FILLER_53_2877 ();
 sg13g2_fill_2 FILLER_53_2892 ();
 sg13g2_fill_1 FILLER_53_2894 ();
 sg13g2_fill_2 FILLER_53_2910 ();
 sg13g2_fill_1 FILLER_53_2912 ();
 sg13g2_fill_2 FILLER_53_2932 ();
 sg13g2_decap_8 FILLER_53_2938 ();
 sg13g2_fill_2 FILLER_53_2945 ();
 sg13g2_fill_2 FILLER_53_2973 ();
 sg13g2_fill_1 FILLER_53_2975 ();
 sg13g2_decap_4 FILLER_53_3010 ();
 sg13g2_fill_1 FILLER_53_3014 ();
 sg13g2_decap_4 FILLER_53_3028 ();
 sg13g2_fill_2 FILLER_53_3073 ();
 sg13g2_fill_1 FILLER_53_3075 ();
 sg13g2_decap_4 FILLER_53_3105 ();
 sg13g2_fill_2 FILLER_53_3109 ();
 sg13g2_decap_8 FILLER_53_3138 ();
 sg13g2_decap_4 FILLER_53_3145 ();
 sg13g2_fill_1 FILLER_53_3175 ();
 sg13g2_decap_8 FILLER_53_3208 ();
 sg13g2_fill_1 FILLER_53_3215 ();
 sg13g2_decap_4 FILLER_53_3225 ();
 sg13g2_fill_2 FILLER_53_3229 ();
 sg13g2_decap_4 FILLER_53_3254 ();
 sg13g2_fill_1 FILLER_53_3258 ();
 sg13g2_fill_1 FILLER_53_3263 ();
 sg13g2_fill_1 FILLER_53_3272 ();
 sg13g2_fill_2 FILLER_53_3314 ();
 sg13g2_fill_1 FILLER_53_3316 ();
 sg13g2_decap_4 FILLER_53_3333 ();
 sg13g2_fill_2 FILLER_53_3358 ();
 sg13g2_fill_1 FILLER_53_3395 ();
 sg13g2_fill_2 FILLER_53_3416 ();
 sg13g2_fill_1 FILLER_53_3418 ();
 sg13g2_decap_4 FILLER_53_3446 ();
 sg13g2_decap_8 FILLER_53_3498 ();
 sg13g2_decap_8 FILLER_53_3535 ();
 sg13g2_fill_1 FILLER_53_3579 ();
 sg13g2_decap_4 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_30 ();
 sg13g2_fill_1 FILLER_54_32 ();
 sg13g2_fill_2 FILLER_54_41 ();
 sg13g2_fill_2 FILLER_54_68 ();
 sg13g2_fill_2 FILLER_54_75 ();
 sg13g2_fill_1 FILLER_54_129 ();
 sg13g2_fill_1 FILLER_54_160 ();
 sg13g2_fill_1 FILLER_54_169 ();
 sg13g2_fill_1 FILLER_54_189 ();
 sg13g2_fill_2 FILLER_54_205 ();
 sg13g2_fill_2 FILLER_54_227 ();
 sg13g2_fill_2 FILLER_54_297 ();
 sg13g2_decap_4 FILLER_54_349 ();
 sg13g2_fill_1 FILLER_54_353 ();
 sg13g2_fill_1 FILLER_54_362 ();
 sg13g2_fill_2 FILLER_54_380 ();
 sg13g2_fill_1 FILLER_54_390 ();
 sg13g2_decap_4 FILLER_54_408 ();
 sg13g2_decap_8 FILLER_54_417 ();
 sg13g2_decap_4 FILLER_54_424 ();
 sg13g2_fill_1 FILLER_54_428 ();
 sg13g2_fill_1 FILLER_54_442 ();
 sg13g2_fill_1 FILLER_54_459 ();
 sg13g2_fill_2 FILLER_54_484 ();
 sg13g2_fill_1 FILLER_54_486 ();
 sg13g2_decap_8 FILLER_54_501 ();
 sg13g2_fill_1 FILLER_54_508 ();
 sg13g2_decap_4 FILLER_54_543 ();
 sg13g2_fill_1 FILLER_54_555 ();
 sg13g2_decap_4 FILLER_54_573 ();
 sg13g2_fill_1 FILLER_54_577 ();
 sg13g2_decap_4 FILLER_54_595 ();
 sg13g2_fill_1 FILLER_54_599 ();
 sg13g2_fill_1 FILLER_54_612 ();
 sg13g2_decap_8 FILLER_54_623 ();
 sg13g2_fill_2 FILLER_54_630 ();
 sg13g2_fill_1 FILLER_54_632 ();
 sg13g2_fill_2 FILLER_54_646 ();
 sg13g2_fill_2 FILLER_54_664 ();
 sg13g2_decap_8 FILLER_54_694 ();
 sg13g2_fill_1 FILLER_54_701 ();
 sg13g2_fill_1 FILLER_54_715 ();
 sg13g2_fill_1 FILLER_54_726 ();
 sg13g2_fill_2 FILLER_54_747 ();
 sg13g2_fill_1 FILLER_54_749 ();
 sg13g2_decap_8 FILLER_54_785 ();
 sg13g2_fill_1 FILLER_54_792 ();
 sg13g2_fill_2 FILLER_54_805 ();
 sg13g2_decap_8 FILLER_54_812 ();
 sg13g2_fill_2 FILLER_54_843 ();
 sg13g2_decap_8 FILLER_54_878 ();
 sg13g2_decap_4 FILLER_54_885 ();
 sg13g2_fill_1 FILLER_54_894 ();
 sg13g2_decap_8 FILLER_54_900 ();
 sg13g2_decap_4 FILLER_54_918 ();
 sg13g2_fill_2 FILLER_54_946 ();
 sg13g2_fill_1 FILLER_54_948 ();
 sg13g2_fill_2 FILLER_54_977 ();
 sg13g2_fill_1 FILLER_54_979 ();
 sg13g2_fill_2 FILLER_54_996 ();
 sg13g2_decap_4 FILLER_54_1016 ();
 sg13g2_fill_1 FILLER_54_1033 ();
 sg13g2_fill_2 FILLER_54_1081 ();
 sg13g2_fill_1 FILLER_54_1083 ();
 sg13g2_decap_4 FILLER_54_1103 ();
 sg13g2_decap_8 FILLER_54_1112 ();
 sg13g2_decap_8 FILLER_54_1132 ();
 sg13g2_decap_4 FILLER_54_1139 ();
 sg13g2_fill_2 FILLER_54_1167 ();
 sg13g2_fill_1 FILLER_54_1169 ();
 sg13g2_fill_1 FILLER_54_1193 ();
 sg13g2_decap_4 FILLER_54_1199 ();
 sg13g2_decap_8 FILLER_54_1262 ();
 sg13g2_fill_2 FILLER_54_1269 ();
 sg13g2_fill_1 FILLER_54_1271 ();
 sg13g2_fill_1 FILLER_54_1282 ();
 sg13g2_fill_2 FILLER_54_1291 ();
 sg13g2_fill_2 FILLER_54_1297 ();
 sg13g2_fill_1 FILLER_54_1299 ();
 sg13g2_fill_1 FILLER_54_1332 ();
 sg13g2_fill_1 FILLER_54_1340 ();
 sg13g2_fill_2 FILLER_54_1364 ();
 sg13g2_fill_1 FILLER_54_1366 ();
 sg13g2_fill_1 FILLER_54_1457 ();
 sg13g2_fill_2 FILLER_54_1496 ();
 sg13g2_fill_1 FILLER_54_1498 ();
 sg13g2_fill_2 FILLER_54_1520 ();
 sg13g2_fill_1 FILLER_54_1522 ();
 sg13g2_fill_2 FILLER_54_1563 ();
 sg13g2_fill_1 FILLER_54_1565 ();
 sg13g2_fill_2 FILLER_54_1574 ();
 sg13g2_fill_2 FILLER_54_1609 ();
 sg13g2_fill_1 FILLER_54_1611 ();
 sg13g2_fill_1 FILLER_54_1620 ();
 sg13g2_fill_1 FILLER_54_1631 ();
 sg13g2_decap_8 FILLER_54_1637 ();
 sg13g2_decap_4 FILLER_54_1654 ();
 sg13g2_fill_2 FILLER_54_1658 ();
 sg13g2_fill_1 FILLER_54_1692 ();
 sg13g2_decap_8 FILLER_54_1748 ();
 sg13g2_fill_2 FILLER_54_1755 ();
 sg13g2_decap_8 FILLER_54_1766 ();
 sg13g2_fill_1 FILLER_54_1778 ();
 sg13g2_decap_8 FILLER_54_1788 ();
 sg13g2_decap_8 FILLER_54_1795 ();
 sg13g2_decap_8 FILLER_54_1809 ();
 sg13g2_fill_2 FILLER_54_1825 ();
 sg13g2_fill_1 FILLER_54_1827 ();
 sg13g2_fill_1 FILLER_54_1836 ();
 sg13g2_fill_1 FILLER_54_1864 ();
 sg13g2_decap_4 FILLER_54_1883 ();
 sg13g2_fill_1 FILLER_54_1887 ();
 sg13g2_decap_4 FILLER_54_1898 ();
 sg13g2_fill_2 FILLER_54_1902 ();
 sg13g2_fill_1 FILLER_54_1913 ();
 sg13g2_fill_2 FILLER_54_1976 ();
 sg13g2_fill_1 FILLER_54_1978 ();
 sg13g2_fill_2 FILLER_54_2050 ();
 sg13g2_fill_1 FILLER_54_2052 ();
 sg13g2_fill_2 FILLER_54_2066 ();
 sg13g2_fill_1 FILLER_54_2082 ();
 sg13g2_fill_1 FILLER_54_2128 ();
 sg13g2_fill_2 FILLER_54_2133 ();
 sg13g2_fill_1 FILLER_54_2135 ();
 sg13g2_decap_4 FILLER_54_2149 ();
 sg13g2_decap_8 FILLER_54_2178 ();
 sg13g2_fill_1 FILLER_54_2185 ();
 sg13g2_fill_1 FILLER_54_2195 ();
 sg13g2_fill_1 FILLER_54_2200 ();
 sg13g2_decap_8 FILLER_54_2241 ();
 sg13g2_fill_2 FILLER_54_2248 ();
 sg13g2_fill_1 FILLER_54_2250 ();
 sg13g2_fill_2 FILLER_54_2283 ();
 sg13g2_fill_1 FILLER_54_2285 ();
 sg13g2_decap_8 FILLER_54_2307 ();
 sg13g2_decap_4 FILLER_54_2342 ();
 sg13g2_decap_4 FILLER_54_2359 ();
 sg13g2_fill_2 FILLER_54_2363 ();
 sg13g2_fill_2 FILLER_54_2390 ();
 sg13g2_fill_1 FILLER_54_2392 ();
 sg13g2_decap_4 FILLER_54_2411 ();
 sg13g2_fill_1 FILLER_54_2415 ();
 sg13g2_fill_2 FILLER_54_2425 ();
 sg13g2_decap_8 FILLER_54_2453 ();
 sg13g2_fill_1 FILLER_54_2460 ();
 sg13g2_decap_4 FILLER_54_2503 ();
 sg13g2_fill_2 FILLER_54_2507 ();
 sg13g2_fill_1 FILLER_54_2530 ();
 sg13g2_fill_2 FILLER_54_2536 ();
 sg13g2_fill_1 FILLER_54_2538 ();
 sg13g2_fill_1 FILLER_54_2557 ();
 sg13g2_fill_2 FILLER_54_2607 ();
 sg13g2_fill_1 FILLER_54_2609 ();
 sg13g2_fill_2 FILLER_54_2629 ();
 sg13g2_fill_2 FILLER_54_2693 ();
 sg13g2_fill_2 FILLER_54_2751 ();
 sg13g2_fill_1 FILLER_54_2753 ();
 sg13g2_fill_2 FILLER_54_2789 ();
 sg13g2_fill_1 FILLER_54_2791 ();
 sg13g2_fill_2 FILLER_54_2807 ();
 sg13g2_fill_2 FILLER_54_2817 ();
 sg13g2_fill_1 FILLER_54_2819 ();
 sg13g2_fill_2 FILLER_54_2841 ();
 sg13g2_fill_2 FILLER_54_2857 ();
 sg13g2_fill_2 FILLER_54_2872 ();
 sg13g2_fill_1 FILLER_54_2907 ();
 sg13g2_fill_2 FILLER_54_2944 ();
 sg13g2_fill_1 FILLER_54_2946 ();
 sg13g2_fill_1 FILLER_54_2964 ();
 sg13g2_fill_2 FILLER_54_2981 ();
 sg13g2_fill_1 FILLER_54_2983 ();
 sg13g2_decap_4 FILLER_54_2992 ();
 sg13g2_decap_8 FILLER_54_3006 ();
 sg13g2_decap_8 FILLER_54_3013 ();
 sg13g2_decap_8 FILLER_54_3036 ();
 sg13g2_fill_2 FILLER_54_3043 ();
 sg13g2_fill_1 FILLER_54_3045 ();
 sg13g2_decap_8 FILLER_54_3057 ();
 sg13g2_decap_8 FILLER_54_3064 ();
 sg13g2_decap_8 FILLER_54_3071 ();
 sg13g2_fill_2 FILLER_54_3102 ();
 sg13g2_decap_8 FILLER_54_3113 ();
 sg13g2_fill_2 FILLER_54_3120 ();
 sg13g2_decap_8 FILLER_54_3152 ();
 sg13g2_fill_1 FILLER_54_3159 ();
 sg13g2_decap_8 FILLER_54_3173 ();
 sg13g2_fill_2 FILLER_54_3180 ();
 sg13g2_fill_2 FILLER_54_3199 ();
 sg13g2_fill_2 FILLER_54_3250 ();
 sg13g2_fill_1 FILLER_54_3252 ();
 sg13g2_fill_1 FILLER_54_3276 ();
 sg13g2_fill_2 FILLER_54_3290 ();
 sg13g2_decap_4 FILLER_54_3304 ();
 sg13g2_fill_2 FILLER_54_3308 ();
 sg13g2_fill_1 FILLER_54_3326 ();
 sg13g2_decap_8 FILLER_54_3337 ();
 sg13g2_decap_4 FILLER_54_3344 ();
 sg13g2_decap_8 FILLER_54_3357 ();
 sg13g2_fill_2 FILLER_54_3381 ();
 sg13g2_fill_1 FILLER_54_3383 ();
 sg13g2_fill_2 FILLER_54_3396 ();
 sg13g2_fill_1 FILLER_54_3398 ();
 sg13g2_fill_1 FILLER_54_3420 ();
 sg13g2_decap_8 FILLER_54_3444 ();
 sg13g2_fill_2 FILLER_54_3496 ();
 sg13g2_fill_1 FILLER_54_3498 ();
 sg13g2_fill_1 FILLER_54_3507 ();
 sg13g2_fill_2 FILLER_54_3520 ();
 sg13g2_fill_1 FILLER_54_3527 ();
 sg13g2_fill_2 FILLER_54_3540 ();
 sg13g2_decap_4 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_4 ();
 sg13g2_fill_2 FILLER_55_46 ();
 sg13g2_decap_4 FILLER_55_85 ();
 sg13g2_fill_1 FILLER_55_89 ();
 sg13g2_fill_2 FILLER_55_129 ();
 sg13g2_fill_2 FILLER_55_136 ();
 sg13g2_fill_1 FILLER_55_138 ();
 sg13g2_fill_2 FILLER_55_158 ();
 sg13g2_fill_1 FILLER_55_160 ();
 sg13g2_fill_2 FILLER_55_174 ();
 sg13g2_fill_2 FILLER_55_189 ();
 sg13g2_fill_2 FILLER_55_205 ();
 sg13g2_fill_2 FILLER_55_212 ();
 sg13g2_fill_1 FILLER_55_259 ();
 sg13g2_fill_2 FILLER_55_370 ();
 sg13g2_fill_1 FILLER_55_443 ();
 sg13g2_decap_8 FILLER_55_470 ();
 sg13g2_decap_8 FILLER_55_477 ();
 sg13g2_fill_1 FILLER_55_484 ();
 sg13g2_fill_2 FILLER_55_492 ();
 sg13g2_fill_1 FILLER_55_494 ();
 sg13g2_fill_2 FILLER_55_500 ();
 sg13g2_fill_1 FILLER_55_502 ();
 sg13g2_fill_2 FILLER_55_533 ();
 sg13g2_fill_1 FILLER_55_535 ();
 sg13g2_fill_1 FILLER_55_551 ();
 sg13g2_fill_2 FILLER_55_570 ();
 sg13g2_decap_4 FILLER_55_580 ();
 sg13g2_fill_2 FILLER_55_584 ();
 sg13g2_decap_8 FILLER_55_595 ();
 sg13g2_fill_2 FILLER_55_602 ();
 sg13g2_decap_4 FILLER_55_629 ();
 sg13g2_fill_2 FILLER_55_633 ();
 sg13g2_fill_2 FILLER_55_641 ();
 sg13g2_fill_1 FILLER_55_643 ();
 sg13g2_fill_1 FILLER_55_661 ();
 sg13g2_fill_1 FILLER_55_705 ();
 sg13g2_fill_2 FILLER_55_727 ();
 sg13g2_fill_1 FILLER_55_729 ();
 sg13g2_fill_1 FILLER_55_735 ();
 sg13g2_decap_8 FILLER_55_749 ();
 sg13g2_decap_4 FILLER_55_756 ();
 sg13g2_fill_1 FILLER_55_760 ();
 sg13g2_decap_4 FILLER_55_780 ();
 sg13g2_decap_8 FILLER_55_789 ();
 sg13g2_fill_1 FILLER_55_809 ();
 sg13g2_fill_2 FILLER_55_815 ();
 sg13g2_fill_1 FILLER_55_817 ();
 sg13g2_decap_8 FILLER_55_850 ();
 sg13g2_fill_1 FILLER_55_857 ();
 sg13g2_fill_2 FILLER_55_908 ();
 sg13g2_fill_2 FILLER_55_920 ();
 sg13g2_fill_1 FILLER_55_931 ();
 sg13g2_fill_2 FILLER_55_962 ();
 sg13g2_fill_1 FILLER_55_964 ();
 sg13g2_decap_4 FILLER_55_973 ();
 sg13g2_fill_1 FILLER_55_977 ();
 sg13g2_fill_1 FILLER_55_991 ();
 sg13g2_fill_1 FILLER_55_1027 ();
 sg13g2_decap_4 FILLER_55_1041 ();
 sg13g2_fill_1 FILLER_55_1045 ();
 sg13g2_fill_1 FILLER_55_1064 ();
 sg13g2_fill_2 FILLER_55_1119 ();
 sg13g2_fill_1 FILLER_55_1121 ();
 sg13g2_decap_4 FILLER_55_1140 ();
 sg13g2_fill_1 FILLER_55_1144 ();
 sg13g2_fill_1 FILLER_55_1156 ();
 sg13g2_decap_4 FILLER_55_1166 ();
 sg13g2_fill_1 FILLER_55_1170 ();
 sg13g2_decap_8 FILLER_55_1194 ();
 sg13g2_decap_4 FILLER_55_1201 ();
 sg13g2_fill_2 FILLER_55_1222 ();
 sg13g2_fill_2 FILLER_55_1237 ();
 sg13g2_decap_4 FILLER_55_1243 ();
 sg13g2_fill_1 FILLER_55_1263 ();
 sg13g2_fill_2 FILLER_55_1293 ();
 sg13g2_fill_1 FILLER_55_1295 ();
 sg13g2_fill_2 FILLER_55_1328 ();
 sg13g2_fill_2 FILLER_55_1381 ();
 sg13g2_fill_1 FILLER_55_1383 ();
 sg13g2_decap_4 FILLER_55_1398 ();
 sg13g2_decap_8 FILLER_55_1433 ();
 sg13g2_fill_2 FILLER_55_1440 ();
 sg13g2_fill_1 FILLER_55_1442 ();
 sg13g2_decap_4 FILLER_55_1456 ();
 sg13g2_decap_8 FILLER_55_1473 ();
 sg13g2_decap_8 FILLER_55_1480 ();
 sg13g2_fill_1 FILLER_55_1497 ();
 sg13g2_fill_1 FILLER_55_1526 ();
 sg13g2_fill_2 FILLER_55_1532 ();
 sg13g2_decap_4 FILLER_55_1564 ();
 sg13g2_fill_2 FILLER_55_1568 ();
 sg13g2_decap_8 FILLER_55_1603 ();
 sg13g2_decap_4 FILLER_55_1623 ();
 sg13g2_fill_2 FILLER_55_1627 ();
 sg13g2_fill_2 FILLER_55_1634 ();
 sg13g2_fill_1 FILLER_55_1636 ();
 sg13g2_fill_2 FILLER_55_1665 ();
 sg13g2_decap_4 FILLER_55_1693 ();
 sg13g2_fill_1 FILLER_55_1714 ();
 sg13g2_fill_2 FILLER_55_1727 ();
 sg13g2_fill_2 FILLER_55_1749 ();
 sg13g2_fill_1 FILLER_55_1751 ();
 sg13g2_fill_1 FILLER_55_1778 ();
 sg13g2_decap_4 FILLER_55_1794 ();
 sg13g2_fill_1 FILLER_55_1816 ();
 sg13g2_fill_2 FILLER_55_1855 ();
 sg13g2_fill_1 FILLER_55_1870 ();
 sg13g2_fill_1 FILLER_55_1875 ();
 sg13g2_fill_2 FILLER_55_1907 ();
 sg13g2_fill_1 FILLER_55_1919 ();
 sg13g2_fill_2 FILLER_55_1933 ();
 sg13g2_fill_1 FILLER_55_1958 ();
 sg13g2_fill_2 FILLER_55_1977 ();
 sg13g2_fill_2 FILLER_55_1992 ();
 sg13g2_fill_1 FILLER_55_2034 ();
 sg13g2_decap_4 FILLER_55_2056 ();
 sg13g2_fill_1 FILLER_55_2073 ();
 sg13g2_fill_1 FILLER_55_2102 ();
 sg13g2_decap_4 FILLER_55_2153 ();
 sg13g2_fill_2 FILLER_55_2157 ();
 sg13g2_decap_4 FILLER_55_2177 ();
 sg13g2_fill_2 FILLER_55_2181 ();
 sg13g2_fill_2 FILLER_55_2204 ();
 sg13g2_fill_2 FILLER_55_2232 ();
 sg13g2_fill_1 FILLER_55_2234 ();
 sg13g2_fill_1 FILLER_55_2244 ();
 sg13g2_fill_2 FILLER_55_2253 ();
 sg13g2_decap_4 FILLER_55_2260 ();
 sg13g2_fill_2 FILLER_55_2264 ();
 sg13g2_fill_2 FILLER_55_2271 ();
 sg13g2_fill_1 FILLER_55_2277 ();
 sg13g2_fill_2 FILLER_55_2281 ();
 sg13g2_fill_1 FILLER_55_2283 ();
 sg13g2_fill_2 FILLER_55_2289 ();
 sg13g2_decap_4 FILLER_55_2338 ();
 sg13g2_fill_2 FILLER_55_2342 ();
 sg13g2_decap_8 FILLER_55_2357 ();
 sg13g2_fill_2 FILLER_55_2364 ();
 sg13g2_fill_1 FILLER_55_2366 ();
 sg13g2_fill_1 FILLER_55_2376 ();
 sg13g2_decap_4 FILLER_55_2393 ();
 sg13g2_fill_1 FILLER_55_2397 ();
 sg13g2_fill_1 FILLER_55_2406 ();
 sg13g2_decap_8 FILLER_55_2442 ();
 sg13g2_decap_4 FILLER_55_2481 ();
 sg13g2_fill_2 FILLER_55_2485 ();
 sg13g2_fill_2 FILLER_55_2500 ();
 sg13g2_fill_1 FILLER_55_2514 ();
 sg13g2_fill_2 FILLER_55_2527 ();
 sg13g2_fill_1 FILLER_55_2529 ();
 sg13g2_fill_2 FILLER_55_2555 ();
 sg13g2_fill_1 FILLER_55_2557 ();
 sg13g2_fill_1 FILLER_55_2567 ();
 sg13g2_fill_2 FILLER_55_2577 ();
 sg13g2_fill_1 FILLER_55_2579 ();
 sg13g2_fill_2 FILLER_55_2593 ();
 sg13g2_fill_1 FILLER_55_2595 ();
 sg13g2_fill_2 FILLER_55_2625 ();
 sg13g2_fill_1 FILLER_55_2627 ();
 sg13g2_fill_2 FILLER_55_2649 ();
 sg13g2_fill_2 FILLER_55_2677 ();
 sg13g2_decap_4 FILLER_55_2692 ();
 sg13g2_fill_2 FILLER_55_2696 ();
 sg13g2_fill_1 FILLER_55_2706 ();
 sg13g2_decap_8 FILLER_55_2720 ();
 sg13g2_fill_2 FILLER_55_2727 ();
 sg13g2_fill_2 FILLER_55_2772 ();
 sg13g2_fill_1 FILLER_55_2787 ();
 sg13g2_decap_8 FILLER_55_2812 ();
 sg13g2_fill_2 FILLER_55_2819 ();
 sg13g2_fill_1 FILLER_55_2825 ();
 sg13g2_decap_4 FILLER_55_2845 ();
 sg13g2_decap_4 FILLER_55_2888 ();
 sg13g2_fill_1 FILLER_55_2892 ();
 sg13g2_decap_4 FILLER_55_2906 ();
 sg13g2_fill_1 FILLER_55_2931 ();
 sg13g2_fill_2 FILLER_55_2937 ();
 sg13g2_fill_2 FILLER_55_2949 ();
 sg13g2_fill_2 FILLER_55_2974 ();
 sg13g2_fill_1 FILLER_55_2976 ();
 sg13g2_decap_8 FILLER_55_2985 ();
 sg13g2_fill_1 FILLER_55_2992 ();
 sg13g2_fill_1 FILLER_55_3004 ();
 sg13g2_fill_1 FILLER_55_3048 ();
 sg13g2_fill_1 FILLER_55_3053 ();
 sg13g2_decap_4 FILLER_55_3082 ();
 sg13g2_fill_2 FILLER_55_3086 ();
 sg13g2_fill_1 FILLER_55_3121 ();
 sg13g2_decap_8 FILLER_55_3143 ();
 sg13g2_decap_4 FILLER_55_3150 ();
 sg13g2_fill_2 FILLER_55_3167 ();
 sg13g2_fill_1 FILLER_55_3181 ();
 sg13g2_fill_2 FILLER_55_3208 ();
 sg13g2_decap_8 FILLER_55_3223 ();
 sg13g2_decap_4 FILLER_55_3230 ();
 sg13g2_fill_2 FILLER_55_3234 ();
 sg13g2_fill_2 FILLER_55_3253 ();
 sg13g2_fill_1 FILLER_55_3255 ();
 sg13g2_fill_2 FILLER_55_3292 ();
 sg13g2_fill_1 FILLER_55_3294 ();
 sg13g2_fill_1 FILLER_55_3310 ();
 sg13g2_fill_1 FILLER_55_3318 ();
 sg13g2_decap_8 FILLER_55_3327 ();
 sg13g2_decap_8 FILLER_55_3334 ();
 sg13g2_decap_4 FILLER_55_3368 ();
 sg13g2_decap_4 FILLER_55_3377 ();
 sg13g2_fill_1 FILLER_55_3381 ();
 sg13g2_decap_8 FILLER_55_3397 ();
 sg13g2_decap_4 FILLER_55_3404 ();
 sg13g2_fill_2 FILLER_55_3408 ();
 sg13g2_decap_8 FILLER_55_3450 ();
 sg13g2_fill_1 FILLER_55_3478 ();
 sg13g2_decap_4 FILLER_55_3497 ();
 sg13g2_fill_1 FILLER_55_3501 ();
 sg13g2_decap_8 FILLER_55_3514 ();
 sg13g2_decap_8 FILLER_55_3521 ();
 sg13g2_fill_2 FILLER_55_3528 ();
 sg13g2_decap_4 FILLER_55_3547 ();
 sg13g2_fill_1 FILLER_55_3579 ();
 sg13g2_fill_1 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_27 ();
 sg13g2_fill_1 FILLER_56_29 ();
 sg13g2_decap_4 FILLER_56_47 ();
 sg13g2_fill_2 FILLER_56_51 ();
 sg13g2_fill_2 FILLER_56_75 ();
 sg13g2_fill_1 FILLER_56_77 ();
 sg13g2_fill_2 FILLER_56_83 ();
 sg13g2_fill_1 FILLER_56_85 ();
 sg13g2_decap_4 FILLER_56_100 ();
 sg13g2_fill_2 FILLER_56_104 ();
 sg13g2_fill_1 FILLER_56_125 ();
 sg13g2_fill_2 FILLER_56_153 ();
 sg13g2_fill_1 FILLER_56_155 ();
 sg13g2_fill_2 FILLER_56_169 ();
 sg13g2_fill_2 FILLER_56_179 ();
 sg13g2_fill_2 FILLER_56_213 ();
 sg13g2_fill_2 FILLER_56_336 ();
 sg13g2_fill_1 FILLER_56_366 ();
 sg13g2_fill_2 FILLER_56_384 ();
 sg13g2_fill_2 FILLER_56_413 ();
 sg13g2_decap_8 FILLER_56_423 ();
 sg13g2_decap_4 FILLER_56_430 ();
 sg13g2_fill_2 FILLER_56_434 ();
 sg13g2_decap_8 FILLER_56_502 ();
 sg13g2_fill_2 FILLER_56_509 ();
 sg13g2_fill_1 FILLER_56_511 ();
 sg13g2_decap_8 FILLER_56_516 ();
 sg13g2_fill_2 FILLER_56_523 ();
 sg13g2_decap_4 FILLER_56_540 ();
 sg13g2_fill_2 FILLER_56_544 ();
 sg13g2_fill_2 FILLER_56_558 ();
 sg13g2_fill_1 FILLER_56_560 ();
 sg13g2_fill_2 FILLER_56_569 ();
 sg13g2_fill_1 FILLER_56_571 ();
 sg13g2_fill_2 FILLER_56_581 ();
 sg13g2_fill_1 FILLER_56_583 ();
 sg13g2_fill_2 FILLER_56_590 ();
 sg13g2_decap_8 FILLER_56_605 ();
 sg13g2_fill_1 FILLER_56_612 ();
 sg13g2_fill_1 FILLER_56_624 ();
 sg13g2_decap_4 FILLER_56_638 ();
 sg13g2_fill_2 FILLER_56_672 ();
 sg13g2_fill_2 FILLER_56_694 ();
 sg13g2_decap_4 FILLER_56_702 ();
 sg13g2_decap_8 FILLER_56_719 ();
 sg13g2_decap_8 FILLER_56_758 ();
 sg13g2_fill_1 FILLER_56_765 ();
 sg13g2_decap_4 FILLER_56_789 ();
 sg13g2_fill_1 FILLER_56_793 ();
 sg13g2_fill_1 FILLER_56_804 ();
 sg13g2_decap_4 FILLER_56_826 ();
 sg13g2_fill_2 FILLER_56_866 ();
 sg13g2_fill_1 FILLER_56_882 ();
 sg13g2_fill_2 FILLER_56_897 ();
 sg13g2_fill_1 FILLER_56_899 ();
 sg13g2_fill_1 FILLER_56_928 ();
 sg13g2_fill_2 FILLER_56_941 ();
 sg13g2_fill_1 FILLER_56_948 ();
 sg13g2_fill_2 FILLER_56_966 ();
 sg13g2_fill_1 FILLER_56_968 ();
 sg13g2_decap_4 FILLER_56_995 ();
 sg13g2_fill_2 FILLER_56_1014 ();
 sg13g2_fill_2 FILLER_56_1036 ();
 sg13g2_fill_1 FILLER_56_1038 ();
 sg13g2_fill_1 FILLER_56_1057 ();
 sg13g2_decap_4 FILLER_56_1085 ();
 sg13g2_fill_1 FILLER_56_1105 ();
 sg13g2_decap_4 FILLER_56_1115 ();
 sg13g2_fill_1 FILLER_56_1119 ();
 sg13g2_fill_2 FILLER_56_1145 ();
 sg13g2_fill_1 FILLER_56_1147 ();
 sg13g2_fill_1 FILLER_56_1158 ();
 sg13g2_decap_8 FILLER_56_1170 ();
 sg13g2_fill_1 FILLER_56_1177 ();
 sg13g2_fill_2 FILLER_56_1198 ();
 sg13g2_fill_1 FILLER_56_1200 ();
 sg13g2_fill_2 FILLER_56_1224 ();
 sg13g2_fill_1 FILLER_56_1226 ();
 sg13g2_decap_4 FILLER_56_1235 ();
 sg13g2_fill_1 FILLER_56_1239 ();
 sg13g2_decap_8 FILLER_56_1294 ();
 sg13g2_decap_4 FILLER_56_1301 ();
 sg13g2_fill_2 FILLER_56_1305 ();
 sg13g2_fill_2 FILLER_56_1325 ();
 sg13g2_fill_2 FILLER_56_1370 ();
 sg13g2_fill_1 FILLER_56_1372 ();
 sg13g2_fill_2 FILLER_56_1386 ();
 sg13g2_fill_2 FILLER_56_1396 ();
 sg13g2_fill_2 FILLER_56_1403 ();
 sg13g2_fill_1 FILLER_56_1405 ();
 sg13g2_fill_2 FILLER_56_1436 ();
 sg13g2_fill_2 FILLER_56_1453 ();
 sg13g2_fill_2 FILLER_56_1459 ();
 sg13g2_decap_8 FILLER_56_1477 ();
 sg13g2_decap_4 FILLER_56_1484 ();
 sg13g2_fill_1 FILLER_56_1496 ();
 sg13g2_fill_1 FILLER_56_1579 ();
 sg13g2_decap_4 FILLER_56_1621 ();
 sg13g2_fill_2 FILLER_56_1657 ();
 sg13g2_fill_1 FILLER_56_1659 ();
 sg13g2_fill_2 FILLER_56_1683 ();
 sg13g2_decap_4 FILLER_56_1717 ();
 sg13g2_fill_1 FILLER_56_1721 ();
 sg13g2_fill_2 FILLER_56_1735 ();
 sg13g2_decap_8 FILLER_56_1760 ();
 sg13g2_fill_2 FILLER_56_1767 ();
 sg13g2_fill_2 FILLER_56_1777 ();
 sg13g2_fill_2 FILLER_56_1803 ();
 sg13g2_decap_8 FILLER_56_1812 ();
 sg13g2_decap_8 FILLER_56_1819 ();
 sg13g2_fill_2 FILLER_56_1826 ();
 sg13g2_fill_1 FILLER_56_1836 ();
 sg13g2_fill_1 FILLER_56_1842 ();
 sg13g2_decap_4 FILLER_56_1859 ();
 sg13g2_fill_1 FILLER_56_1863 ();
 sg13g2_fill_2 FILLER_56_1881 ();
 sg13g2_fill_2 FILLER_56_1888 ();
 sg13g2_decap_8 FILLER_56_1902 ();
 sg13g2_fill_2 FILLER_56_1909 ();
 sg13g2_fill_2 FILLER_56_1952 ();
 sg13g2_fill_1 FILLER_56_1954 ();
 sg13g2_fill_2 FILLER_56_1971 ();
 sg13g2_fill_1 FILLER_56_1973 ();
 sg13g2_fill_1 FILLER_56_2012 ();
 sg13g2_fill_2 FILLER_56_2033 ();
 sg13g2_fill_1 FILLER_56_2035 ();
 sg13g2_fill_1 FILLER_56_2073 ();
 sg13g2_fill_2 FILLER_56_2082 ();
 sg13g2_fill_1 FILLER_56_2084 ();
 sg13g2_decap_4 FILLER_56_2099 ();
 sg13g2_fill_2 FILLER_56_2121 ();
 sg13g2_fill_1 FILLER_56_2123 ();
 sg13g2_fill_2 FILLER_56_2154 ();
 sg13g2_decap_4 FILLER_56_2182 ();
 sg13g2_fill_2 FILLER_56_2186 ();
 sg13g2_fill_1 FILLER_56_2219 ();
 sg13g2_decap_4 FILLER_56_2258 ();
 sg13g2_fill_2 FILLER_56_2267 ();
 sg13g2_fill_1 FILLER_56_2280 ();
 sg13g2_fill_2 FILLER_56_2327 ();
 sg13g2_fill_1 FILLER_56_2342 ();
 sg13g2_decap_4 FILLER_56_2352 ();
 sg13g2_fill_1 FILLER_56_2356 ();
 sg13g2_fill_1 FILLER_56_2369 ();
 sg13g2_fill_2 FILLER_56_2399 ();
 sg13g2_fill_1 FILLER_56_2401 ();
 sg13g2_fill_1 FILLER_56_2407 ();
 sg13g2_decap_4 FILLER_56_2416 ();
 sg13g2_fill_1 FILLER_56_2420 ();
 sg13g2_decap_4 FILLER_56_2460 ();
 sg13g2_decap_8 FILLER_56_2490 ();
 sg13g2_fill_1 FILLER_56_2497 ();
 sg13g2_fill_2 FILLER_56_2502 ();
 sg13g2_fill_1 FILLER_56_2535 ();
 sg13g2_fill_2 FILLER_56_2563 ();
 sg13g2_fill_1 FILLER_56_2565 ();
 sg13g2_fill_1 FILLER_56_2577 ();
 sg13g2_fill_2 FILLER_56_2599 ();
 sg13g2_fill_1 FILLER_56_2601 ();
 sg13g2_fill_2 FILLER_56_2607 ();
 sg13g2_fill_1 FILLER_56_2609 ();
 sg13g2_decap_8 FILLER_56_2672 ();
 sg13g2_fill_2 FILLER_56_2679 ();
 sg13g2_decap_4 FILLER_56_2725 ();
 sg13g2_decap_4 FILLER_56_2735 ();
 sg13g2_fill_2 FILLER_56_2739 ();
 sg13g2_fill_2 FILLER_56_2753 ();
 sg13g2_fill_1 FILLER_56_2755 ();
 sg13g2_decap_8 FILLER_56_2816 ();
 sg13g2_fill_1 FILLER_56_2823 ();
 sg13g2_fill_1 FILLER_56_2850 ();
 sg13g2_fill_2 FILLER_56_2856 ();
 sg13g2_fill_1 FILLER_56_2891 ();
 sg13g2_decap_8 FILLER_56_2912 ();
 sg13g2_fill_1 FILLER_56_2919 ();
 sg13g2_fill_2 FILLER_56_2957 ();
 sg13g2_fill_1 FILLER_56_2959 ();
 sg13g2_decap_8 FILLER_56_2977 ();
 sg13g2_fill_2 FILLER_56_2984 ();
 sg13g2_fill_2 FILLER_56_3011 ();
 sg13g2_fill_1 FILLER_56_3013 ();
 sg13g2_fill_2 FILLER_56_3022 ();
 sg13g2_fill_2 FILLER_56_3038 ();
 sg13g2_decap_8 FILLER_56_3065 ();
 sg13g2_fill_1 FILLER_56_3072 ();
 sg13g2_fill_1 FILLER_56_3080 ();
 sg13g2_fill_2 FILLER_56_3097 ();
 sg13g2_fill_1 FILLER_56_3104 ();
 sg13g2_decap_4 FILLER_56_3115 ();
 sg13g2_fill_1 FILLER_56_3129 ();
 sg13g2_decap_8 FILLER_56_3143 ();
 sg13g2_fill_2 FILLER_56_3150 ();
 sg13g2_fill_1 FILLER_56_3152 ();
 sg13g2_fill_2 FILLER_56_3178 ();
 sg13g2_fill_1 FILLER_56_3180 ();
 sg13g2_fill_2 FILLER_56_3226 ();
 sg13g2_fill_1 FILLER_56_3228 ();
 sg13g2_fill_2 FILLER_56_3255 ();
 sg13g2_fill_1 FILLER_56_3257 ();
 sg13g2_fill_2 FILLER_56_3294 ();
 sg13g2_fill_1 FILLER_56_3296 ();
 sg13g2_fill_2 FILLER_56_3309 ();
 sg13g2_fill_1 FILLER_56_3339 ();
 sg13g2_decap_4 FILLER_56_3386 ();
 sg13g2_decap_8 FILLER_56_3446 ();
 sg13g2_decap_8 FILLER_56_3470 ();
 sg13g2_fill_1 FILLER_56_3497 ();
 sg13g2_fill_1 FILLER_56_3525 ();
 sg13g2_fill_1 FILLER_56_3554 ();
 sg13g2_decap_8 FILLER_56_3564 ();
 sg13g2_decap_8 FILLER_56_3571 ();
 sg13g2_fill_2 FILLER_56_3578 ();
 sg13g2_fill_1 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_38 ();
 sg13g2_fill_1 FILLER_57_60 ();
 sg13g2_fill_1 FILLER_57_69 ();
 sg13g2_fill_2 FILLER_57_82 ();
 sg13g2_fill_1 FILLER_57_84 ();
 sg13g2_fill_1 FILLER_57_93 ();
 sg13g2_fill_2 FILLER_57_102 ();
 sg13g2_fill_2 FILLER_57_118 ();
 sg13g2_fill_1 FILLER_57_120 ();
 sg13g2_decap_4 FILLER_57_125 ();
 sg13g2_fill_1 FILLER_57_129 ();
 sg13g2_fill_2 FILLER_57_147 ();
 sg13g2_fill_1 FILLER_57_149 ();
 sg13g2_fill_2 FILLER_57_155 ();
 sg13g2_fill_2 FILLER_57_192 ();
 sg13g2_fill_1 FILLER_57_262 ();
 sg13g2_fill_1 FILLER_57_331 ();
 sg13g2_fill_2 FILLER_57_364 ();
 sg13g2_fill_1 FILLER_57_472 ();
 sg13g2_fill_1 FILLER_57_478 ();
 sg13g2_fill_2 FILLER_57_488 ();
 sg13g2_fill_1 FILLER_57_490 ();
 sg13g2_decap_8 FILLER_57_496 ();
 sg13g2_fill_1 FILLER_57_503 ();
 sg13g2_fill_2 FILLER_57_541 ();
 sg13g2_fill_1 FILLER_57_543 ();
 sg13g2_decap_4 FILLER_57_547 ();
 sg13g2_fill_2 FILLER_57_551 ();
 sg13g2_fill_1 FILLER_57_581 ();
 sg13g2_decap_4 FILLER_57_595 ();
 sg13g2_decap_8 FILLER_57_615 ();
 sg13g2_decap_4 FILLER_57_622 ();
 sg13g2_fill_1 FILLER_57_648 ();
 sg13g2_fill_1 FILLER_57_662 ();
 sg13g2_fill_1 FILLER_57_685 ();
 sg13g2_decap_4 FILLER_57_703 ();
 sg13g2_fill_1 FILLER_57_730 ();
 sg13g2_fill_2 FILLER_57_785 ();
 sg13g2_fill_2 FILLER_57_802 ();
 sg13g2_fill_1 FILLER_57_804 ();
 sg13g2_fill_1 FILLER_57_818 ();
 sg13g2_fill_2 FILLER_57_824 ();
 sg13g2_fill_1 FILLER_57_826 ();
 sg13g2_fill_2 FILLER_57_836 ();
 sg13g2_fill_1 FILLER_57_838 ();
 sg13g2_fill_1 FILLER_57_865 ();
 sg13g2_decap_8 FILLER_57_898 ();
 sg13g2_fill_2 FILLER_57_905 ();
 sg13g2_fill_1 FILLER_57_912 ();
 sg13g2_fill_2 FILLER_57_923 ();
 sg13g2_fill_2 FILLER_57_939 ();
 sg13g2_fill_2 FILLER_57_945 ();
 sg13g2_fill_1 FILLER_57_1006 ();
 sg13g2_decap_8 FILLER_57_1020 ();
 sg13g2_fill_2 FILLER_57_1027 ();
 sg13g2_fill_1 FILLER_57_1029 ();
 sg13g2_decap_8 FILLER_57_1034 ();
 sg13g2_decap_4 FILLER_57_1065 ();
 sg13g2_fill_1 FILLER_57_1069 ();
 sg13g2_fill_2 FILLER_57_1078 ();
 sg13g2_fill_1 FILLER_57_1080 ();
 sg13g2_fill_1 FILLER_57_1101 ();
 sg13g2_decap_8 FILLER_57_1107 ();
 sg13g2_decap_4 FILLER_57_1114 ();
 sg13g2_decap_8 FILLER_57_1137 ();
 sg13g2_decap_4 FILLER_57_1144 ();
 sg13g2_fill_2 FILLER_57_1148 ();
 sg13g2_fill_2 FILLER_57_1176 ();
 sg13g2_decap_4 FILLER_57_1186 ();
 sg13g2_fill_2 FILLER_57_1190 ();
 sg13g2_decap_4 FILLER_57_1200 ();
 sg13g2_fill_2 FILLER_57_1231 ();
 sg13g2_decap_4 FILLER_57_1241 ();
 sg13g2_decap_4 FILLER_57_1296 ();
 sg13g2_fill_1 FILLER_57_1300 ();
 sg13g2_fill_2 FILLER_57_1331 ();
 sg13g2_decap_8 FILLER_57_1336 ();
 sg13g2_fill_1 FILLER_57_1343 ();
 sg13g2_fill_1 FILLER_57_1378 ();
 sg13g2_fill_1 FILLER_57_1393 ();
 sg13g2_fill_1 FILLER_57_1402 ();
 sg13g2_fill_2 FILLER_57_1414 ();
 sg13g2_decap_4 FILLER_57_1426 ();
 sg13g2_fill_2 FILLER_57_1430 ();
 sg13g2_decap_4 FILLER_57_1437 ();
 sg13g2_fill_1 FILLER_57_1441 ();
 sg13g2_fill_1 FILLER_57_1447 ();
 sg13g2_fill_2 FILLER_57_1453 ();
 sg13g2_fill_1 FILLER_57_1455 ();
 sg13g2_fill_1 FILLER_57_1461 ();
 sg13g2_decap_8 FILLER_57_1475 ();
 sg13g2_fill_2 FILLER_57_1482 ();
 sg13g2_fill_1 FILLER_57_1504 ();
 sg13g2_fill_1 FILLER_57_1510 ();
 sg13g2_decap_4 FILLER_57_1527 ();
 sg13g2_decap_8 FILLER_57_1535 ();
 sg13g2_fill_1 FILLER_57_1542 ();
 sg13g2_fill_2 FILLER_57_1571 ();
 sg13g2_fill_2 FILLER_57_1606 ();
 sg13g2_fill_1 FILLER_57_1616 ();
 sg13g2_fill_1 FILLER_57_1624 ();
 sg13g2_fill_2 FILLER_57_1653 ();
 sg13g2_fill_1 FILLER_57_1655 ();
 sg13g2_fill_2 FILLER_57_1660 ();
 sg13g2_fill_1 FILLER_57_1662 ();
 sg13g2_fill_1 FILLER_57_1671 ();
 sg13g2_fill_2 FILLER_57_1685 ();
 sg13g2_fill_1 FILLER_57_1687 ();
 sg13g2_fill_1 FILLER_57_1712 ();
 sg13g2_decap_4 FILLER_57_1737 ();
 sg13g2_fill_1 FILLER_57_1741 ();
 sg13g2_decap_8 FILLER_57_1758 ();
 sg13g2_fill_2 FILLER_57_1765 ();
 sg13g2_fill_1 FILLER_57_1767 ();
 sg13g2_decap_8 FILLER_57_1783 ();
 sg13g2_fill_2 FILLER_57_1790 ();
 sg13g2_fill_1 FILLER_57_1792 ();
 sg13g2_decap_4 FILLER_57_1823 ();
 sg13g2_fill_1 FILLER_57_1827 ();
 sg13g2_decap_4 FILLER_57_1847 ();
 sg13g2_fill_1 FILLER_57_1851 ();
 sg13g2_fill_1 FILLER_57_1884 ();
 sg13g2_decap_8 FILLER_57_1908 ();
 sg13g2_decap_4 FILLER_57_1915 ();
 sg13g2_fill_1 FILLER_57_1933 ();
 sg13g2_decap_4 FILLER_57_1938 ();
 sg13g2_fill_2 FILLER_57_1942 ();
 sg13g2_fill_1 FILLER_57_1970 ();
 sg13g2_fill_2 FILLER_57_1984 ();
 sg13g2_decap_4 FILLER_57_2015 ();
 sg13g2_fill_1 FILLER_57_2019 ();
 sg13g2_decap_8 FILLER_57_2037 ();
 sg13g2_fill_1 FILLER_57_2044 ();
 sg13g2_fill_2 FILLER_57_2053 ();
 sg13g2_fill_2 FILLER_57_2063 ();
 sg13g2_fill_2 FILLER_57_2078 ();
 sg13g2_fill_2 FILLER_57_2100 ();
 sg13g2_fill_1 FILLER_57_2119 ();
 sg13g2_fill_2 FILLER_57_2133 ();
 sg13g2_fill_1 FILLER_57_2135 ();
 sg13g2_fill_2 FILLER_57_2162 ();
 sg13g2_fill_1 FILLER_57_2164 ();
 sg13g2_fill_2 FILLER_57_2192 ();
 sg13g2_decap_4 FILLER_57_2199 ();
 sg13g2_fill_2 FILLER_57_2203 ();
 sg13g2_decap_4 FILLER_57_2229 ();
 sg13g2_fill_2 FILLER_57_2242 ();
 sg13g2_decap_4 FILLER_57_2257 ();
 sg13g2_decap_8 FILLER_57_2275 ();
 sg13g2_decap_4 FILLER_57_2330 ();
 sg13g2_fill_1 FILLER_57_2334 ();
 sg13g2_decap_4 FILLER_57_2359 ();
 sg13g2_fill_1 FILLER_57_2363 ();
 sg13g2_decap_8 FILLER_57_2390 ();
 sg13g2_fill_1 FILLER_57_2421 ();
 sg13g2_fill_1 FILLER_57_2449 ();
 sg13g2_fill_2 FILLER_57_2459 ();
 sg13g2_fill_1 FILLER_57_2461 ();
 sg13g2_decap_4 FILLER_57_2473 ();
 sg13g2_fill_1 FILLER_57_2477 ();
 sg13g2_fill_2 FILLER_57_2515 ();
 sg13g2_fill_1 FILLER_57_2517 ();
 sg13g2_decap_4 FILLER_57_2526 ();
 sg13g2_fill_1 FILLER_57_2530 ();
 sg13g2_fill_2 FILLER_57_2535 ();
 sg13g2_fill_1 FILLER_57_2537 ();
 sg13g2_fill_2 FILLER_57_2571 ();
 sg13g2_fill_2 FILLER_57_2601 ();
 sg13g2_fill_1 FILLER_57_2644 ();
 sg13g2_fill_1 FILLER_57_2653 ();
 sg13g2_fill_2 FILLER_57_2670 ();
 sg13g2_fill_1 FILLER_57_2672 ();
 sg13g2_fill_1 FILLER_57_2699 ();
 sg13g2_fill_2 FILLER_57_2719 ();
 sg13g2_fill_1 FILLER_57_2721 ();
 sg13g2_fill_2 FILLER_57_2796 ();
 sg13g2_fill_1 FILLER_57_2815 ();
 sg13g2_decap_4 FILLER_57_2821 ();
 sg13g2_fill_2 FILLER_57_2825 ();
 sg13g2_fill_1 FILLER_57_2835 ();
 sg13g2_fill_2 FILLER_57_2868 ();
 sg13g2_fill_2 FILLER_57_2887 ();
 sg13g2_decap_8 FILLER_57_2902 ();
 sg13g2_fill_2 FILLER_57_2909 ();
 sg13g2_fill_1 FILLER_57_2911 ();
 sg13g2_decap_8 FILLER_57_2916 ();
 sg13g2_fill_2 FILLER_57_2923 ();
 sg13g2_decap_4 FILLER_57_2960 ();
 sg13g2_fill_1 FILLER_57_2964 ();
 sg13g2_decap_8 FILLER_57_2975 ();
 sg13g2_decap_8 FILLER_57_2982 ();
 sg13g2_fill_1 FILLER_57_3006 ();
 sg13g2_fill_2 FILLER_57_3012 ();
 sg13g2_fill_1 FILLER_57_3014 ();
 sg13g2_fill_2 FILLER_57_3028 ();
 sg13g2_decap_8 FILLER_57_3048 ();
 sg13g2_decap_8 FILLER_57_3055 ();
 sg13g2_fill_2 FILLER_57_3075 ();
 sg13g2_fill_1 FILLER_57_3077 ();
 sg13g2_fill_2 FILLER_57_3091 ();
 sg13g2_fill_2 FILLER_57_3098 ();
 sg13g2_decap_4 FILLER_57_3113 ();
 sg13g2_fill_1 FILLER_57_3133 ();
 sg13g2_fill_2 FILLER_57_3148 ();
 sg13g2_fill_1 FILLER_57_3150 ();
 sg13g2_fill_1 FILLER_57_3164 ();
 sg13g2_fill_2 FILLER_57_3174 ();
 sg13g2_fill_1 FILLER_57_3176 ();
 sg13g2_fill_2 FILLER_57_3182 ();
 sg13g2_fill_1 FILLER_57_3205 ();
 sg13g2_fill_2 FILLER_57_3211 ();
 sg13g2_fill_1 FILLER_57_3213 ();
 sg13g2_fill_2 FILLER_57_3227 ();
 sg13g2_fill_2 FILLER_57_3232 ();
 sg13g2_fill_1 FILLER_57_3234 ();
 sg13g2_fill_2 FILLER_57_3271 ();
 sg13g2_fill_1 FILLER_57_3278 ();
 sg13g2_fill_1 FILLER_57_3284 ();
 sg13g2_fill_1 FILLER_57_3295 ();
 sg13g2_fill_2 FILLER_57_3301 ();
 sg13g2_fill_1 FILLER_57_3303 ();
 sg13g2_decap_4 FILLER_57_3312 ();
 sg13g2_decap_8 FILLER_57_3320 ();
 sg13g2_decap_4 FILLER_57_3327 ();
 sg13g2_fill_1 FILLER_57_3331 ();
 sg13g2_decap_4 FILLER_57_3335 ();
 sg13g2_decap_8 FILLER_57_3344 ();
 sg13g2_fill_2 FILLER_57_3351 ();
 sg13g2_fill_1 FILLER_57_3353 ();
 sg13g2_decap_8 FILLER_57_3364 ();
 sg13g2_fill_2 FILLER_57_3371 ();
 sg13g2_decap_4 FILLER_57_3380 ();
 sg13g2_fill_1 FILLER_57_3384 ();
 sg13g2_decap_4 FILLER_57_3390 ();
 sg13g2_fill_1 FILLER_57_3394 ();
 sg13g2_decap_8 FILLER_57_3399 ();
 sg13g2_decap_4 FILLER_57_3406 ();
 sg13g2_fill_2 FILLER_57_3410 ();
 sg13g2_fill_2 FILLER_57_3425 ();
 sg13g2_fill_1 FILLER_57_3427 ();
 sg13g2_fill_1 FILLER_57_3441 ();
 sg13g2_fill_2 FILLER_57_3447 ();
 sg13g2_decap_4 FILLER_57_3473 ();
 sg13g2_decap_4 FILLER_57_3503 ();
 sg13g2_fill_2 FILLER_57_3507 ();
 sg13g2_fill_1 FILLER_57_3526 ();
 sg13g2_decap_8 FILLER_57_3536 ();
 sg13g2_decap_8 FILLER_57_3543 ();
 sg13g2_decap_4 FILLER_57_3550 ();
 sg13g2_fill_2 FILLER_57_3554 ();
 sg13g2_decap_8 FILLER_57_3564 ();
 sg13g2_decap_8 FILLER_57_3571 ();
 sg13g2_fill_2 FILLER_57_3578 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_fill_1 FILLER_58_14 ();
 sg13g2_fill_2 FILLER_58_61 ();
 sg13g2_fill_1 FILLER_58_63 ();
 sg13g2_fill_2 FILLER_58_67 ();
 sg13g2_fill_1 FILLER_58_69 ();
 sg13g2_decap_8 FILLER_58_75 ();
 sg13g2_fill_1 FILLER_58_82 ();
 sg13g2_fill_2 FILLER_58_99 ();
 sg13g2_fill_1 FILLER_58_107 ();
 sg13g2_fill_2 FILLER_58_120 ();
 sg13g2_fill_1 FILLER_58_122 ();
 sg13g2_fill_2 FILLER_58_132 ();
 sg13g2_fill_2 FILLER_58_145 ();
 sg13g2_fill_1 FILLER_58_147 ();
 sg13g2_fill_1 FILLER_58_173 ();
 sg13g2_fill_1 FILLER_58_307 ();
 sg13g2_fill_1 FILLER_58_316 ();
 sg13g2_fill_1 FILLER_58_332 ();
 sg13g2_fill_1 FILLER_58_353 ();
 sg13g2_fill_2 FILLER_58_371 ();
 sg13g2_fill_2 FILLER_58_382 ();
 sg13g2_decap_4 FILLER_58_397 ();
 sg13g2_fill_1 FILLER_58_427 ();
 sg13g2_fill_2 FILLER_58_436 ();
 sg13g2_fill_1 FILLER_58_438 ();
 sg13g2_decap_8 FILLER_58_471 ();
 sg13g2_fill_1 FILLER_58_478 ();
 sg13g2_fill_1 FILLER_58_507 ();
 sg13g2_decap_8 FILLER_58_512 ();
 sg13g2_decap_8 FILLER_58_519 ();
 sg13g2_fill_2 FILLER_58_533 ();
 sg13g2_fill_1 FILLER_58_535 ();
 sg13g2_fill_2 FILLER_58_549 ();
 sg13g2_fill_2 FILLER_58_555 ();
 sg13g2_decap_8 FILLER_58_561 ();
 sg13g2_fill_1 FILLER_58_572 ();
 sg13g2_fill_1 FILLER_58_579 ();
 sg13g2_decap_4 FILLER_58_626 ();
 sg13g2_fill_1 FILLER_58_635 ();
 sg13g2_decap_8 FILLER_58_640 ();
 sg13g2_decap_4 FILLER_58_647 ();
 sg13g2_fill_2 FILLER_58_651 ();
 sg13g2_fill_2 FILLER_58_727 ();
 sg13g2_fill_1 FILLER_58_729 ();
 sg13g2_decap_8 FILLER_58_757 ();
 sg13g2_decap_4 FILLER_58_764 ();
 sg13g2_fill_2 FILLER_58_768 ();
 sg13g2_fill_2 FILLER_58_799 ();
 sg13g2_fill_1 FILLER_58_801 ();
 sg13g2_fill_1 FILLER_58_846 ();
 sg13g2_fill_2 FILLER_58_874 ();
 sg13g2_fill_2 FILLER_58_927 ();
 sg13g2_decap_8 FILLER_58_941 ();
 sg13g2_fill_1 FILLER_58_948 ();
 sg13g2_fill_2 FILLER_58_975 ();
 sg13g2_decap_4 FILLER_58_987 ();
 sg13g2_decap_8 FILLER_58_996 ();
 sg13g2_decap_4 FILLER_58_1003 ();
 sg13g2_decap_8 FILLER_58_1039 ();
 sg13g2_fill_2 FILLER_58_1090 ();
 sg13g2_fill_1 FILLER_58_1092 ();
 sg13g2_fill_1 FILLER_58_1119 ();
 sg13g2_decap_4 FILLER_58_1144 ();
 sg13g2_decap_8 FILLER_58_1188 ();
 sg13g2_fill_1 FILLER_58_1211 ();
 sg13g2_decap_4 FILLER_58_1232 ();
 sg13g2_fill_1 FILLER_58_1236 ();
 sg13g2_fill_1 FILLER_58_1242 ();
 sg13g2_decap_8 FILLER_58_1258 ();
 sg13g2_decap_8 FILLER_58_1265 ();
 sg13g2_fill_2 FILLER_58_1272 ();
 sg13g2_fill_1 FILLER_58_1277 ();
 sg13g2_decap_8 FILLER_58_1298 ();
 sg13g2_decap_4 FILLER_58_1337 ();
 sg13g2_fill_1 FILLER_58_1341 ();
 sg13g2_fill_1 FILLER_58_1362 ();
 sg13g2_fill_2 FILLER_58_1377 ();
 sg13g2_decap_4 FILLER_58_1396 ();
 sg13g2_fill_2 FILLER_58_1409 ();
 sg13g2_fill_1 FILLER_58_1411 ();
 sg13g2_decap_8 FILLER_58_1430 ();
 sg13g2_decap_8 FILLER_58_1437 ();
 sg13g2_fill_2 FILLER_58_1444 ();
 sg13g2_fill_1 FILLER_58_1446 ();
 sg13g2_fill_2 FILLER_58_1472 ();
 sg13g2_fill_2 FILLER_58_1483 ();
 sg13g2_fill_2 FILLER_58_1503 ();
 sg13g2_fill_2 FILLER_58_1510 ();
 sg13g2_fill_2 FILLER_58_1527 ();
 sg13g2_decap_8 FILLER_58_1542 ();
 sg13g2_fill_2 FILLER_58_1549 ();
 sg13g2_decap_8 FILLER_58_1561 ();
 sg13g2_fill_1 FILLER_58_1568 ();
 sg13g2_fill_2 FILLER_58_1607 ();
 sg13g2_fill_1 FILLER_58_1609 ();
 sg13g2_fill_2 FILLER_58_1632 ();
 sg13g2_fill_1 FILLER_58_1634 ();
 sg13g2_fill_1 FILLER_58_1699 ();
 sg13g2_decap_4 FILLER_58_1754 ();
 sg13g2_fill_2 FILLER_58_1758 ();
 sg13g2_decap_8 FILLER_58_1791 ();
 sg13g2_decap_4 FILLER_58_1798 ();
 sg13g2_fill_1 FILLER_58_1802 ();
 sg13g2_fill_2 FILLER_58_1831 ();
 sg13g2_fill_1 FILLER_58_1841 ();
 sg13g2_decap_8 FILLER_58_1852 ();
 sg13g2_decap_8 FILLER_58_1868 ();
 sg13g2_decap_4 FILLER_58_1875 ();
 sg13g2_fill_2 FILLER_58_1908 ();
 sg13g2_fill_1 FILLER_58_1938 ();
 sg13g2_fill_2 FILLER_58_1952 ();
 sg13g2_decap_4 FILLER_58_1968 ();
 sg13g2_fill_1 FILLER_58_1972 ();
 sg13g2_fill_2 FILLER_58_1976 ();
 sg13g2_fill_1 FILLER_58_1978 ();
 sg13g2_fill_2 FILLER_58_1997 ();
 sg13g2_decap_8 FILLER_58_2007 ();
 sg13g2_decap_8 FILLER_58_2046 ();
 sg13g2_fill_2 FILLER_58_2053 ();
 sg13g2_fill_1 FILLER_58_2055 ();
 sg13g2_decap_8 FILLER_58_2078 ();
 sg13g2_fill_2 FILLER_58_2098 ();
 sg13g2_fill_1 FILLER_58_2100 ();
 sg13g2_fill_1 FILLER_58_2105 ();
 sg13g2_decap_4 FILLER_58_2134 ();
 sg13g2_fill_1 FILLER_58_2151 ();
 sg13g2_fill_2 FILLER_58_2187 ();
 sg13g2_decap_4 FILLER_58_2197 ();
 sg13g2_fill_2 FILLER_58_2201 ();
 sg13g2_fill_2 FILLER_58_2258 ();
 sg13g2_fill_1 FILLER_58_2268 ();
 sg13g2_fill_1 FILLER_58_2355 ();
 sg13g2_decap_8 FILLER_58_2393 ();
 sg13g2_fill_2 FILLER_58_2400 ();
 sg13g2_fill_1 FILLER_58_2402 ();
 sg13g2_fill_2 FILLER_58_2420 ();
 sg13g2_fill_1 FILLER_58_2422 ();
 sg13g2_decap_4 FILLER_58_2443 ();
 sg13g2_fill_2 FILLER_58_2447 ();
 sg13g2_fill_2 FILLER_58_2469 ();
 sg13g2_fill_1 FILLER_58_2471 ();
 sg13g2_fill_1 FILLER_58_2478 ();
 sg13g2_decap_4 FILLER_58_2584 ();
 sg13g2_fill_2 FILLER_58_2588 ();
 sg13g2_fill_1 FILLER_58_2607 ();
 sg13g2_fill_1 FILLER_58_2679 ();
 sg13g2_decap_4 FILLER_58_2684 ();
 sg13g2_fill_1 FILLER_58_2688 ();
 sg13g2_fill_2 FILLER_58_2724 ();
 sg13g2_fill_1 FILLER_58_2744 ();
 sg13g2_fill_2 FILLER_58_2776 ();
 sg13g2_fill_1 FILLER_58_2778 ();
 sg13g2_fill_1 FILLER_58_2791 ();
 sg13g2_fill_1 FILLER_58_2814 ();
 sg13g2_fill_2 FILLER_58_2845 ();
 sg13g2_fill_1 FILLER_58_2851 ();
 sg13g2_fill_2 FILLER_58_2861 ();
 sg13g2_fill_1 FILLER_58_2863 ();
 sg13g2_fill_2 FILLER_58_2872 ();
 sg13g2_fill_2 FILLER_58_2916 ();
 sg13g2_fill_1 FILLER_58_2931 ();
 sg13g2_fill_2 FILLER_58_2969 ();
 sg13g2_decap_8 FILLER_58_2979 ();
 sg13g2_decap_8 FILLER_58_3012 ();
 sg13g2_fill_1 FILLER_58_3019 ();
 sg13g2_fill_1 FILLER_58_3024 ();
 sg13g2_decap_4 FILLER_58_3049 ();
 sg13g2_fill_2 FILLER_58_3053 ();
 sg13g2_fill_2 FILLER_58_3090 ();
 sg13g2_decap_8 FILLER_58_3105 ();
 sg13g2_fill_1 FILLER_58_3112 ();
 sg13g2_decap_4 FILLER_58_3116 ();
 sg13g2_decap_8 FILLER_58_3141 ();
 sg13g2_fill_1 FILLER_58_3148 ();
 sg13g2_fill_2 FILLER_58_3162 ();
 sg13g2_fill_1 FILLER_58_3164 ();
 sg13g2_fill_1 FILLER_58_3178 ();
 sg13g2_fill_1 FILLER_58_3189 ();
 sg13g2_fill_2 FILLER_58_3203 ();
 sg13g2_fill_2 FILLER_58_3209 ();
 sg13g2_fill_1 FILLER_58_3211 ();
 sg13g2_decap_4 FILLER_58_3219 ();
 sg13g2_decap_8 FILLER_58_3244 ();
 sg13g2_decap_8 FILLER_58_3251 ();
 sg13g2_fill_1 FILLER_58_3267 ();
 sg13g2_fill_1 FILLER_58_3273 ();
 sg13g2_fill_2 FILLER_58_3291 ();
 sg13g2_fill_2 FILLER_58_3298 ();
 sg13g2_fill_1 FILLER_58_3300 ();
 sg13g2_fill_2 FILLER_58_3311 ();
 sg13g2_decap_8 FILLER_58_3318 ();
 sg13g2_fill_1 FILLER_58_3343 ();
 sg13g2_fill_2 FILLER_58_3356 ();
 sg13g2_fill_1 FILLER_58_3364 ();
 sg13g2_fill_1 FILLER_58_3372 ();
 sg13g2_fill_1 FILLER_58_3393 ();
 sg13g2_fill_1 FILLER_58_3427 ();
 sg13g2_fill_2 FILLER_58_3448 ();
 sg13g2_fill_1 FILLER_58_3450 ();
 sg13g2_fill_1 FILLER_58_3480 ();
 sg13g2_fill_2 FILLER_58_3507 ();
 sg13g2_fill_1 FILLER_58_3509 ();
 sg13g2_fill_2 FILLER_58_3527 ();
 sg13g2_fill_2 FILLER_58_3543 ();
 sg13g2_fill_1 FILLER_58_3545 ();
 sg13g2_fill_2 FILLER_58_3549 ();
 sg13g2_fill_1 FILLER_58_3551 ();
 sg13g2_fill_1 FILLER_59_0 ();
 sg13g2_fill_2 FILLER_59_41 ();
 sg13g2_fill_1 FILLER_59_43 ();
 sg13g2_fill_2 FILLER_59_68 ();
 sg13g2_fill_1 FILLER_59_70 ();
 sg13g2_decap_4 FILLER_59_104 ();
 sg13g2_fill_1 FILLER_59_108 ();
 sg13g2_fill_1 FILLER_59_114 ();
 sg13g2_fill_1 FILLER_59_131 ();
 sg13g2_fill_2 FILLER_59_155 ();
 sg13g2_fill_2 FILLER_59_167 ();
 sg13g2_fill_1 FILLER_59_169 ();
 sg13g2_fill_1 FILLER_59_179 ();
 sg13g2_fill_2 FILLER_59_190 ();
 sg13g2_fill_2 FILLER_59_265 ();
 sg13g2_fill_2 FILLER_59_280 ();
 sg13g2_fill_1 FILLER_59_336 ();
 sg13g2_fill_2 FILLER_59_373 ();
 sg13g2_fill_1 FILLER_59_375 ();
 sg13g2_fill_2 FILLER_59_403 ();
 sg13g2_fill_1 FILLER_59_410 ();
 sg13g2_fill_2 FILLER_59_443 ();
 sg13g2_fill_1 FILLER_59_445 ();
 sg13g2_fill_1 FILLER_59_475 ();
 sg13g2_fill_2 FILLER_59_480 ();
 sg13g2_decap_8 FILLER_59_493 ();
 sg13g2_fill_2 FILLER_59_500 ();
 sg13g2_fill_1 FILLER_59_502 ();
 sg13g2_fill_1 FILLER_59_531 ();
 sg13g2_fill_1 FILLER_59_554 ();
 sg13g2_fill_2 FILLER_59_563 ();
 sg13g2_fill_1 FILLER_59_565 ();
 sg13g2_fill_2 FILLER_59_581 ();
 sg13g2_fill_1 FILLER_59_583 ();
 sg13g2_decap_4 FILLER_59_592 ();
 sg13g2_fill_2 FILLER_59_596 ();
 sg13g2_fill_2 FILLER_59_609 ();
 sg13g2_fill_2 FILLER_59_616 ();
 sg13g2_decap_8 FILLER_59_622 ();
 sg13g2_fill_2 FILLER_59_629 ();
 sg13g2_fill_2 FILLER_59_659 ();
 sg13g2_fill_1 FILLER_59_682 ();
 sg13g2_decap_8 FILLER_59_692 ();
 sg13g2_fill_1 FILLER_59_699 ();
 sg13g2_fill_1 FILLER_59_727 ();
 sg13g2_fill_1 FILLER_59_736 ();
 sg13g2_fill_2 FILLER_59_749 ();
 sg13g2_fill_1 FILLER_59_751 ();
 sg13g2_fill_1 FILLER_59_780 ();
 sg13g2_fill_1 FILLER_59_789 ();
 sg13g2_decap_8 FILLER_59_816 ();
 sg13g2_fill_2 FILLER_59_823 ();
 sg13g2_fill_1 FILLER_59_825 ();
 sg13g2_fill_2 FILLER_59_862 ();
 sg13g2_fill_1 FILLER_59_890 ();
 sg13g2_decap_4 FILLER_59_902 ();
 sg13g2_fill_1 FILLER_59_906 ();
 sg13g2_decap_4 FILLER_59_939 ();
 sg13g2_fill_2 FILLER_59_943 ();
 sg13g2_fill_2 FILLER_59_975 ();
 sg13g2_fill_2 FILLER_59_980 ();
 sg13g2_fill_1 FILLER_59_982 ();
 sg13g2_decap_8 FILLER_59_1004 ();
 sg13g2_fill_1 FILLER_59_1011 ();
 sg13g2_fill_1 FILLER_59_1066 ();
 sg13g2_decap_4 FILLER_59_1071 ();
 sg13g2_fill_2 FILLER_59_1075 ();
 sg13g2_fill_1 FILLER_59_1082 ();
 sg13g2_decap_8 FILLER_59_1090 ();
 sg13g2_decap_4 FILLER_59_1097 ();
 sg13g2_fill_1 FILLER_59_1101 ();
 sg13g2_decap_8 FILLER_59_1106 ();
 sg13g2_fill_1 FILLER_59_1113 ();
 sg13g2_decap_8 FILLER_59_1139 ();
 sg13g2_decap_8 FILLER_59_1146 ();
 sg13g2_fill_2 FILLER_59_1153 ();
 sg13g2_decap_8 FILLER_59_1168 ();
 sg13g2_fill_2 FILLER_59_1207 ();
 sg13g2_fill_1 FILLER_59_1209 ();
 sg13g2_decap_8 FILLER_59_1233 ();
 sg13g2_fill_1 FILLER_59_1240 ();
 sg13g2_decap_8 FILLER_59_1269 ();
 sg13g2_decap_8 FILLER_59_1291 ();
 sg13g2_decap_4 FILLER_59_1298 ();
 sg13g2_fill_2 FILLER_59_1302 ();
 sg13g2_fill_2 FILLER_59_1321 ();
 sg13g2_fill_1 FILLER_59_1323 ();
 sg13g2_decap_8 FILLER_59_1337 ();
 sg13g2_fill_2 FILLER_59_1344 ();
 sg13g2_fill_1 FILLER_59_1346 ();
 sg13g2_fill_1 FILLER_59_1405 ();
 sg13g2_fill_1 FILLER_59_1424 ();
 sg13g2_fill_1 FILLER_59_1451 ();
 sg13g2_fill_2 FILLER_59_1473 ();
 sg13g2_fill_1 FILLER_59_1475 ();
 sg13g2_fill_2 FILLER_59_1483 ();
 sg13g2_fill_1 FILLER_59_1485 ();
 sg13g2_fill_2 FILLER_59_1506 ();
 sg13g2_decap_8 FILLER_59_1533 ();
 sg13g2_decap_8 FILLER_59_1540 ();
 sg13g2_fill_1 FILLER_59_1547 ();
 sg13g2_fill_1 FILLER_59_1569 ();
 sg13g2_decap_4 FILLER_59_1584 ();
 sg13g2_fill_1 FILLER_59_1639 ();
 sg13g2_decap_4 FILLER_59_1661 ();
 sg13g2_fill_2 FILLER_59_1665 ();
 sg13g2_decap_8 FILLER_59_1675 ();
 sg13g2_fill_2 FILLER_59_1709 ();
 sg13g2_fill_1 FILLER_59_1720 ();
 sg13g2_fill_1 FILLER_59_1775 ();
 sg13g2_decap_8 FILLER_59_1789 ();
 sg13g2_fill_1 FILLER_59_1823 ();
 sg13g2_fill_2 FILLER_59_1851 ();
 sg13g2_decap_8 FILLER_59_1881 ();
 sg13g2_fill_2 FILLER_59_1888 ();
 sg13g2_fill_1 FILLER_59_1939 ();
 sg13g2_fill_2 FILLER_59_2001 ();
 sg13g2_fill_2 FILLER_59_2034 ();
 sg13g2_fill_1 FILLER_59_2036 ();
 sg13g2_fill_1 FILLER_59_2074 ();
 sg13g2_fill_2 FILLER_59_2103 ();
 sg13g2_fill_1 FILLER_59_2152 ();
 sg13g2_fill_2 FILLER_59_2181 ();
 sg13g2_fill_2 FILLER_59_2188 ();
 sg13g2_fill_1 FILLER_59_2190 ();
 sg13g2_fill_2 FILLER_59_2228 ();
 sg13g2_fill_1 FILLER_59_2230 ();
 sg13g2_decap_8 FILLER_59_2249 ();
 sg13g2_decap_8 FILLER_59_2282 ();
 sg13g2_decap_8 FILLER_59_2289 ();
 sg13g2_fill_2 FILLER_59_2296 ();
 sg13g2_fill_2 FILLER_59_2311 ();
 sg13g2_fill_1 FILLER_59_2313 ();
 sg13g2_fill_2 FILLER_59_2331 ();
 sg13g2_fill_1 FILLER_59_2333 ();
 sg13g2_decap_8 FILLER_59_2390 ();
 sg13g2_decap_4 FILLER_59_2397 ();
 sg13g2_fill_1 FILLER_59_2401 ();
 sg13g2_decap_8 FILLER_59_2419 ();
 sg13g2_decap_8 FILLER_59_2446 ();
 sg13g2_fill_2 FILLER_59_2453 ();
 sg13g2_fill_1 FILLER_59_2455 ();
 sg13g2_decap_4 FILLER_59_2460 ();
 sg13g2_fill_2 FILLER_59_2475 ();
 sg13g2_decap_4 FILLER_59_2488 ();
 sg13g2_fill_2 FILLER_59_2492 ();
 sg13g2_decap_4 FILLER_59_2503 ();
 sg13g2_fill_1 FILLER_59_2526 ();
 sg13g2_fill_1 FILLER_59_2531 ();
 sg13g2_fill_2 FILLER_59_2606 ();
 sg13g2_fill_1 FILLER_59_2608 ();
 sg13g2_fill_1 FILLER_59_2659 ();
 sg13g2_fill_1 FILLER_59_2697 ();
 sg13g2_fill_2 FILLER_59_2703 ();
 sg13g2_fill_1 FILLER_59_2705 ();
 sg13g2_decap_8 FILLER_59_2747 ();
 sg13g2_decap_4 FILLER_59_2758 ();
 sg13g2_fill_1 FILLER_59_2762 ();
 sg13g2_fill_2 FILLER_59_2772 ();
 sg13g2_fill_1 FILLER_59_2774 ();
 sg13g2_fill_1 FILLER_59_2785 ();
 sg13g2_fill_1 FILLER_59_2790 ();
 sg13g2_fill_1 FILLER_59_2800 ();
 sg13g2_fill_2 FILLER_59_2842 ();
 sg13g2_fill_2 FILLER_59_2857 ();
 sg13g2_fill_2 FILLER_59_2881 ();
 sg13g2_fill_2 FILLER_59_2901 ();
 sg13g2_fill_1 FILLER_59_2903 ();
 sg13g2_fill_1 FILLER_59_2917 ();
 sg13g2_fill_2 FILLER_59_2949 ();
 sg13g2_fill_1 FILLER_59_2951 ();
 sg13g2_decap_8 FILLER_59_2967 ();
 sg13g2_fill_1 FILLER_59_2974 ();
 sg13g2_decap_4 FILLER_59_2988 ();
 sg13g2_fill_1 FILLER_59_2992 ();
 sg13g2_decap_4 FILLER_59_3014 ();
 sg13g2_fill_2 FILLER_59_3018 ();
 sg13g2_decap_8 FILLER_59_3040 ();
 sg13g2_fill_2 FILLER_59_3047 ();
 sg13g2_fill_1 FILLER_59_3049 ();
 sg13g2_decap_8 FILLER_59_3075 ();
 sg13g2_fill_2 FILLER_59_3114 ();
 sg13g2_decap_8 FILLER_59_3144 ();
 sg13g2_fill_2 FILLER_59_3151 ();
 sg13g2_fill_1 FILLER_59_3153 ();
 sg13g2_fill_1 FILLER_59_3201 ();
 sg13g2_fill_2 FILLER_59_3228 ();
 sg13g2_decap_4 FILLER_59_3248 ();
 sg13g2_fill_1 FILLER_59_3268 ();
 sg13g2_fill_1 FILLER_59_3305 ();
 sg13g2_fill_2 FILLER_59_3321 ();
 sg13g2_fill_1 FILLER_59_3323 ();
 sg13g2_fill_1 FILLER_59_3336 ();
 sg13g2_decap_4 FILLER_59_3364 ();
 sg13g2_fill_2 FILLER_59_3368 ();
 sg13g2_fill_2 FILLER_59_3378 ();
 sg13g2_decap_4 FILLER_59_3396 ();
 sg13g2_fill_2 FILLER_59_3400 ();
 sg13g2_decap_8 FILLER_59_3410 ();
 sg13g2_decap_4 FILLER_59_3417 ();
 sg13g2_fill_2 FILLER_59_3425 ();
 sg13g2_decap_4 FILLER_59_3441 ();
 sg13g2_fill_1 FILLER_59_3445 ();
 sg13g2_fill_2 FILLER_59_3451 ();
 sg13g2_fill_1 FILLER_59_3453 ();
 sg13g2_decap_8 FILLER_59_3477 ();
 sg13g2_decap_8 FILLER_59_3510 ();
 sg13g2_decap_4 FILLER_59_3517 ();
 sg13g2_fill_1 FILLER_59_3521 ();
 sg13g2_decap_4 FILLER_59_3575 ();
 sg13g2_fill_1 FILLER_59_3579 ();
 sg13g2_decap_4 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_4 ();
 sg13g2_fill_1 FILLER_60_36 ();
 sg13g2_fill_1 FILLER_60_46 ();
 sg13g2_decap_4 FILLER_60_57 ();
 sg13g2_fill_2 FILLER_60_61 ();
 sg13g2_fill_1 FILLER_60_67 ();
 sg13g2_decap_8 FILLER_60_76 ();
 sg13g2_decap_8 FILLER_60_83 ();
 sg13g2_fill_2 FILLER_60_90 ();
 sg13g2_fill_1 FILLER_60_92 ();
 sg13g2_fill_2 FILLER_60_98 ();
 sg13g2_fill_2 FILLER_60_107 ();
 sg13g2_fill_1 FILLER_60_109 ();
 sg13g2_fill_2 FILLER_60_116 ();
 sg13g2_fill_1 FILLER_60_118 ();
 sg13g2_fill_2 FILLER_60_137 ();
 sg13g2_fill_1 FILLER_60_139 ();
 sg13g2_fill_1 FILLER_60_179 ();
 sg13g2_fill_2 FILLER_60_212 ();
 sg13g2_fill_1 FILLER_60_214 ();
 sg13g2_fill_2 FILLER_60_246 ();
 sg13g2_fill_1 FILLER_60_262 ();
 sg13g2_fill_2 FILLER_60_325 ();
 sg13g2_decap_8 FILLER_60_347 ();
 sg13g2_fill_2 FILLER_60_358 ();
 sg13g2_fill_1 FILLER_60_365 ();
 sg13g2_fill_2 FILLER_60_426 ();
 sg13g2_fill_1 FILLER_60_428 ();
 sg13g2_fill_2 FILLER_60_446 ();
 sg13g2_fill_2 FILLER_60_465 ();
 sg13g2_fill_1 FILLER_60_467 ();
 sg13g2_decap_8 FILLER_60_489 ();
 sg13g2_decap_4 FILLER_60_496 ();
 sg13g2_decap_8 FILLER_60_519 ();
 sg13g2_fill_1 FILLER_60_526 ();
 sg13g2_decap_8 FILLER_60_563 ();
 sg13g2_fill_1 FILLER_60_570 ();
 sg13g2_fill_2 FILLER_60_591 ();
 sg13g2_fill_1 FILLER_60_593 ();
 sg13g2_fill_2 FILLER_60_607 ();
 sg13g2_decap_8 FILLER_60_639 ();
 sg13g2_decap_4 FILLER_60_646 ();
 sg13g2_fill_2 FILLER_60_666 ();
 sg13g2_fill_2 FILLER_60_698 ();
 sg13g2_fill_1 FILLER_60_700 ();
 sg13g2_fill_1 FILLER_60_723 ();
 sg13g2_fill_1 FILLER_60_744 ();
 sg13g2_decap_8 FILLER_60_749 ();
 sg13g2_fill_2 FILLER_60_756 ();
 sg13g2_fill_1 FILLER_60_758 ();
 sg13g2_fill_2 FILLER_60_790 ();
 sg13g2_fill_1 FILLER_60_792 ();
 sg13g2_decap_4 FILLER_60_818 ();
 sg13g2_decap_8 FILLER_60_844 ();
 sg13g2_fill_2 FILLER_60_851 ();
 sg13g2_decap_8 FILLER_60_865 ();
 sg13g2_decap_4 FILLER_60_872 ();
 sg13g2_fill_1 FILLER_60_876 ();
 sg13g2_fill_1 FILLER_60_898 ();
 sg13g2_fill_2 FILLER_60_911 ();
 sg13g2_decap_8 FILLER_60_939 ();
 sg13g2_fill_2 FILLER_60_946 ();
 sg13g2_fill_1 FILLER_60_956 ();
 sg13g2_fill_2 FILLER_60_983 ();
 sg13g2_fill_1 FILLER_60_985 ();
 sg13g2_decap_8 FILLER_60_1013 ();
 sg13g2_fill_2 FILLER_60_1020 ();
 sg13g2_fill_1 FILLER_60_1022 ();
 sg13g2_fill_2 FILLER_60_1039 ();
 sg13g2_fill_1 FILLER_60_1041 ();
 sg13g2_decap_4 FILLER_60_1046 ();
 sg13g2_decap_8 FILLER_60_1069 ();
 sg13g2_fill_1 FILLER_60_1076 ();
 sg13g2_fill_2 FILLER_60_1108 ();
 sg13g2_decap_4 FILLER_60_1140 ();
 sg13g2_fill_1 FILLER_60_1144 ();
 sg13g2_fill_1 FILLER_60_1162 ();
 sg13g2_fill_1 FILLER_60_1175 ();
 sg13g2_fill_1 FILLER_60_1180 ();
 sg13g2_decap_8 FILLER_60_1185 ();
 sg13g2_decap_8 FILLER_60_1199 ();
 sg13g2_fill_1 FILLER_60_1206 ();
 sg13g2_fill_2 FILLER_60_1226 ();
 sg13g2_fill_1 FILLER_60_1228 ();
 sg13g2_fill_1 FILLER_60_1266 ();
 sg13g2_fill_2 FILLER_60_1272 ();
 sg13g2_decap_4 FILLER_60_1300 ();
 sg13g2_fill_1 FILLER_60_1314 ();
 sg13g2_fill_2 FILLER_60_1320 ();
 sg13g2_fill_1 FILLER_60_1322 ();
 sg13g2_fill_1 FILLER_60_1335 ();
 sg13g2_fill_2 FILLER_60_1371 ();
 sg13g2_decap_4 FILLER_60_1399 ();
 sg13g2_decap_4 FILLER_60_1437 ();
 sg13g2_fill_2 FILLER_60_1441 ();
 sg13g2_fill_2 FILLER_60_1451 ();
 sg13g2_fill_1 FILLER_60_1453 ();
 sg13g2_decap_4 FILLER_60_1464 ();
 sg13g2_fill_1 FILLER_60_1484 ();
 sg13g2_fill_2 FILLER_60_1509 ();
 sg13g2_fill_1 FILLER_60_1528 ();
 sg13g2_fill_1 FILLER_60_1551 ();
 sg13g2_fill_2 FILLER_60_1569 ();
 sg13g2_fill_2 FILLER_60_1588 ();
 sg13g2_fill_2 FILLER_60_1595 ();
 sg13g2_fill_2 FILLER_60_1607 ();
 sg13g2_fill_2 FILLER_60_1718 ();
 sg13g2_decap_4 FILLER_60_1753 ();
 sg13g2_fill_1 FILLER_60_1836 ();
 sg13g2_fill_1 FILLER_60_1870 ();
 sg13g2_fill_2 FILLER_60_1874 ();
 sg13g2_fill_1 FILLER_60_1876 ();
 sg13g2_decap_8 FILLER_60_1882 ();
 sg13g2_decap_4 FILLER_60_1906 ();
 sg13g2_fill_2 FILLER_60_1933 ();
 sg13g2_decap_4 FILLER_60_1962 ();
 sg13g2_fill_2 FILLER_60_1966 ();
 sg13g2_decap_4 FILLER_60_1972 ();
 sg13g2_fill_2 FILLER_60_2011 ();
 sg13g2_fill_1 FILLER_60_2049 ();
 sg13g2_fill_2 FILLER_60_2059 ();
 sg13g2_fill_1 FILLER_60_2071 ();
 sg13g2_fill_2 FILLER_60_2090 ();
 sg13g2_fill_2 FILLER_60_2145 ();
 sg13g2_fill_2 FILLER_60_2175 ();
 sg13g2_fill_1 FILLER_60_2177 ();
 sg13g2_decap_8 FILLER_60_2215 ();
 sg13g2_fill_1 FILLER_60_2222 ();
 sg13g2_fill_1 FILLER_60_2259 ();
 sg13g2_decap_4 FILLER_60_2342 ();
 sg13g2_fill_2 FILLER_60_2346 ();
 sg13g2_decap_4 FILLER_60_2356 ();
 sg13g2_fill_2 FILLER_60_2372 ();
 sg13g2_fill_1 FILLER_60_2374 ();
 sg13g2_fill_1 FILLER_60_2425 ();
 sg13g2_fill_1 FILLER_60_2454 ();
 sg13g2_fill_2 FILLER_60_2478 ();
 sg13g2_fill_1 FILLER_60_2480 ();
 sg13g2_decap_8 FILLER_60_2518 ();
 sg13g2_decap_4 FILLER_60_2525 ();
 sg13g2_fill_1 FILLER_60_2558 ();
 sg13g2_decap_8 FILLER_60_2581 ();
 sg13g2_decap_4 FILLER_60_2588 ();
 sg13g2_fill_1 FILLER_60_2592 ();
 sg13g2_fill_2 FILLER_60_2632 ();
 sg13g2_fill_1 FILLER_60_2659 ();
 sg13g2_fill_2 FILLER_60_2674 ();
 sg13g2_decap_4 FILLER_60_2684 ();
 sg13g2_fill_1 FILLER_60_2697 ();
 sg13g2_fill_1 FILLER_60_2772 ();
 sg13g2_fill_1 FILLER_60_2810 ();
 sg13g2_decap_8 FILLER_60_2816 ();
 sg13g2_fill_1 FILLER_60_2823 ();
 sg13g2_fill_2 FILLER_60_2831 ();
 sg13g2_fill_1 FILLER_60_2833 ();
 sg13g2_fill_2 FILLER_60_2852 ();
 sg13g2_fill_2 FILLER_60_2887 ();
 sg13g2_fill_1 FILLER_60_2926 ();
 sg13g2_fill_2 FILLER_60_2945 ();
 sg13g2_fill_2 FILLER_60_2967 ();
 sg13g2_fill_1 FILLER_60_2969 ();
 sg13g2_fill_1 FILLER_60_2991 ();
 sg13g2_fill_2 FILLER_60_3021 ();
 sg13g2_decap_4 FILLER_60_3048 ();
 sg13g2_fill_2 FILLER_60_3052 ();
 sg13g2_decap_4 FILLER_60_3071 ();
 sg13g2_fill_2 FILLER_60_3080 ();
 sg13g2_fill_1 FILLER_60_3082 ();
 sg13g2_fill_2 FILLER_60_3088 ();
 sg13g2_fill_1 FILLER_60_3090 ();
 sg13g2_decap_4 FILLER_60_3095 ();
 sg13g2_fill_2 FILLER_60_3108 ();
 sg13g2_fill_2 FILLER_60_3116 ();
 sg13g2_fill_1 FILLER_60_3118 ();
 sg13g2_decap_8 FILLER_60_3124 ();
 sg13g2_decap_8 FILLER_60_3131 ();
 sg13g2_fill_2 FILLER_60_3167 ();
 sg13g2_decap_8 FILLER_60_3191 ();
 sg13g2_fill_1 FILLER_60_3211 ();
 sg13g2_fill_1 FILLER_60_3225 ();
 sg13g2_fill_1 FILLER_60_3244 ();
 sg13g2_fill_1 FILLER_60_3265 ();
 sg13g2_fill_2 FILLER_60_3276 ();
 sg13g2_decap_4 FILLER_60_3288 ();
 sg13g2_fill_1 FILLER_60_3305 ();
 sg13g2_decap_8 FILLER_60_3311 ();
 sg13g2_fill_1 FILLER_60_3318 ();
 sg13g2_decap_4 FILLER_60_3337 ();
 sg13g2_fill_2 FILLER_60_3341 ();
 sg13g2_decap_8 FILLER_60_3359 ();
 sg13g2_decap_8 FILLER_60_3366 ();
 sg13g2_decap_4 FILLER_60_3373 ();
 sg13g2_fill_1 FILLER_60_3377 ();
 sg13g2_fill_2 FILLER_60_3403 ();
 sg13g2_fill_1 FILLER_60_3405 ();
 sg13g2_fill_1 FILLER_60_3411 ();
 sg13g2_fill_1 FILLER_60_3438 ();
 sg13g2_fill_2 FILLER_60_3484 ();
 sg13g2_fill_2 FILLER_60_3495 ();
 sg13g2_fill_1 FILLER_60_3497 ();
 sg13g2_decap_8 FILLER_60_3508 ();
 sg13g2_fill_1 FILLER_60_3515 ();
 sg13g2_fill_2 FILLER_60_3548 ();
 sg13g2_fill_1 FILLER_60_3550 ();
 sg13g2_fill_1 FILLER_60_3579 ();
 sg13g2_fill_1 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_65 ();
 sg13g2_fill_1 FILLER_61_86 ();
 sg13g2_fill_1 FILLER_61_92 ();
 sg13g2_decap_4 FILLER_61_102 ();
 sg13g2_fill_2 FILLER_61_106 ();
 sg13g2_fill_2 FILLER_61_121 ();
 sg13g2_fill_1 FILLER_61_123 ();
 sg13g2_fill_2 FILLER_61_132 ();
 sg13g2_fill_2 FILLER_61_152 ();
 sg13g2_fill_1 FILLER_61_154 ();
 sg13g2_fill_2 FILLER_61_164 ();
 sg13g2_fill_1 FILLER_61_166 ();
 sg13g2_fill_2 FILLER_61_181 ();
 sg13g2_fill_1 FILLER_61_219 ();
 sg13g2_fill_2 FILLER_61_291 ();
 sg13g2_fill_2 FILLER_61_305 ();
 sg13g2_decap_4 FILLER_61_319 ();
 sg13g2_decap_4 FILLER_61_334 ();
 sg13g2_fill_2 FILLER_61_338 ();
 sg13g2_decap_8 FILLER_61_359 ();
 sg13g2_fill_1 FILLER_61_366 ();
 sg13g2_decap_8 FILLER_61_387 ();
 sg13g2_fill_1 FILLER_61_394 ();
 sg13g2_decap_4 FILLER_61_414 ();
 sg13g2_fill_2 FILLER_61_418 ();
 sg13g2_decap_8 FILLER_61_433 ();
 sg13g2_decap_8 FILLER_61_440 ();
 sg13g2_decap_8 FILLER_61_447 ();
 sg13g2_fill_2 FILLER_61_466 ();
 sg13g2_fill_2 FILLER_61_507 ();
 sg13g2_decap_4 FILLER_61_522 ();
 sg13g2_decap_8 FILLER_61_562 ();
 sg13g2_fill_1 FILLER_61_569 ();
 sg13g2_fill_2 FILLER_61_579 ();
 sg13g2_fill_2 FILLER_61_594 ();
 sg13g2_decap_8 FILLER_61_625 ();
 sg13g2_fill_1 FILLER_61_650 ();
 sg13g2_fill_1 FILLER_61_667 ();
 sg13g2_decap_8 FILLER_61_674 ();
 sg13g2_fill_2 FILLER_61_690 ();
 sg13g2_fill_2 FILLER_61_704 ();
 sg13g2_fill_2 FILLER_61_731 ();
 sg13g2_decap_4 FILLER_61_757 ();
 sg13g2_fill_2 FILLER_61_761 ();
 sg13g2_decap_4 FILLER_61_789 ();
 sg13g2_fill_1 FILLER_61_793 ();
 sg13g2_decap_8 FILLER_61_815 ();
 sg13g2_decap_4 FILLER_61_822 ();
 sg13g2_fill_2 FILLER_61_844 ();
 sg13g2_fill_1 FILLER_61_846 ();
 sg13g2_fill_1 FILLER_61_868 ();
 sg13g2_decap_8 FILLER_61_877 ();
 sg13g2_fill_1 FILLER_61_884 ();
 sg13g2_decap_8 FILLER_61_910 ();
 sg13g2_decap_4 FILLER_61_939 ();
 sg13g2_fill_1 FILLER_61_943 ();
 sg13g2_decap_8 FILLER_61_966 ();
 sg13g2_decap_8 FILLER_61_973 ();
 sg13g2_fill_1 FILLER_61_980 ();
 sg13g2_fill_2 FILLER_61_996 ();
 sg13g2_decap_8 FILLER_61_1016 ();
 sg13g2_fill_2 FILLER_61_1023 ();
 sg13g2_fill_1 FILLER_61_1025 ();
 sg13g2_fill_2 FILLER_61_1080 ();
 sg13g2_fill_1 FILLER_61_1082 ();
 sg13g2_decap_4 FILLER_61_1146 ();
 sg13g2_fill_1 FILLER_61_1150 ();
 sg13g2_fill_1 FILLER_61_1182 ();
 sg13g2_fill_2 FILLER_61_1194 ();
 sg13g2_fill_1 FILLER_61_1196 ();
 sg13g2_decap_8 FILLER_61_1202 ();
 sg13g2_fill_1 FILLER_61_1209 ();
 sg13g2_fill_2 FILLER_61_1232 ();
 sg13g2_fill_1 FILLER_61_1243 ();
 sg13g2_fill_2 FILLER_61_1267 ();
 sg13g2_decap_8 FILLER_61_1291 ();
 sg13g2_fill_1 FILLER_61_1298 ();
 sg13g2_decap_8 FILLER_61_1302 ();
 sg13g2_fill_2 FILLER_61_1309 ();
 sg13g2_fill_2 FILLER_61_1355 ();
 sg13g2_fill_1 FILLER_61_1390 ();
 sg13g2_fill_1 FILLER_61_1443 ();
 sg13g2_decap_4 FILLER_61_1474 ();
 sg13g2_fill_2 FILLER_61_1491 ();
 sg13g2_fill_1 FILLER_61_1493 ();
 sg13g2_decap_8 FILLER_61_1517 ();
 sg13g2_decap_8 FILLER_61_1546 ();
 sg13g2_decap_4 FILLER_61_1553 ();
 sg13g2_fill_2 FILLER_61_1564 ();
 sg13g2_fill_2 FILLER_61_1575 ();
 sg13g2_decap_8 FILLER_61_1587 ();
 sg13g2_decap_4 FILLER_61_1623 ();
 sg13g2_decap_4 FILLER_61_1635 ();
 sg13g2_fill_2 FILLER_61_1639 ();
 sg13g2_fill_2 FILLER_61_1651 ();
 sg13g2_fill_1 FILLER_61_1653 ();
 sg13g2_fill_1 FILLER_61_1659 ();
 sg13g2_decap_4 FILLER_61_1664 ();
 sg13g2_decap_8 FILLER_61_1672 ();
 sg13g2_fill_1 FILLER_61_1679 ();
 sg13g2_fill_2 FILLER_61_1684 ();
 sg13g2_fill_1 FILLER_61_1686 ();
 sg13g2_fill_1 FILLER_61_1695 ();
 sg13g2_fill_2 FILLER_61_1704 ();
 sg13g2_decap_8 FILLER_61_1710 ();
 sg13g2_fill_2 FILLER_61_1725 ();
 sg13g2_fill_1 FILLER_61_1731 ();
 sg13g2_decap_8 FILLER_61_1736 ();
 sg13g2_fill_2 FILLER_61_1743 ();
 sg13g2_fill_2 FILLER_61_1763 ();
 sg13g2_fill_1 FILLER_61_1765 ();
 sg13g2_decap_8 FILLER_61_1779 ();
 sg13g2_decap_8 FILLER_61_1786 ();
 sg13g2_decap_8 FILLER_61_1802 ();
 sg13g2_decap_4 FILLER_61_1809 ();
 sg13g2_fill_1 FILLER_61_1813 ();
 sg13g2_fill_1 FILLER_61_1823 ();
 sg13g2_decap_4 FILLER_61_1829 ();
 sg13g2_fill_1 FILLER_61_1833 ();
 sg13g2_fill_2 FILLER_61_1837 ();
 sg13g2_fill_1 FILLER_61_1839 ();
 sg13g2_fill_2 FILLER_61_1847 ();
 sg13g2_fill_1 FILLER_61_1849 ();
 sg13g2_fill_2 FILLER_61_1863 ();
 sg13g2_decap_8 FILLER_61_1902 ();
 sg13g2_decap_8 FILLER_61_1953 ();
 sg13g2_decap_4 FILLER_61_1960 ();
 sg13g2_fill_1 FILLER_61_2070 ();
 sg13g2_fill_1 FILLER_61_2076 ();
 sg13g2_fill_1 FILLER_61_2099 ();
 sg13g2_fill_1 FILLER_61_2115 ();
 sg13g2_decap_8 FILLER_61_2144 ();
 sg13g2_fill_1 FILLER_61_2151 ();
 sg13g2_fill_2 FILLER_61_2156 ();
 sg13g2_decap_8 FILLER_61_2162 ();
 sg13g2_decap_8 FILLER_61_2169 ();
 sg13g2_decap_4 FILLER_61_2200 ();
 sg13g2_fill_1 FILLER_61_2204 ();
 sg13g2_fill_1 FILLER_61_2209 ();
 sg13g2_decap_8 FILLER_61_2231 ();
 sg13g2_decap_8 FILLER_61_2238 ();
 sg13g2_decap_4 FILLER_61_2245 ();
 sg13g2_fill_2 FILLER_61_2253 ();
 sg13g2_fill_1 FILLER_61_2255 ();
 sg13g2_decap_4 FILLER_61_2273 ();
 sg13g2_fill_2 FILLER_61_2277 ();
 sg13g2_decap_8 FILLER_61_2291 ();
 sg13g2_decap_8 FILLER_61_2298 ();
 sg13g2_fill_2 FILLER_61_2305 ();
 sg13g2_fill_1 FILLER_61_2307 ();
 sg13g2_fill_2 FILLER_61_2331 ();
 sg13g2_decap_8 FILLER_61_2346 ();
 sg13g2_fill_2 FILLER_61_2369 ();
 sg13g2_fill_1 FILLER_61_2371 ();
 sg13g2_fill_2 FILLER_61_2393 ();
 sg13g2_decap_4 FILLER_61_2418 ();
 sg13g2_fill_2 FILLER_61_2430 ();
 sg13g2_fill_2 FILLER_61_2438 ();
 sg13g2_fill_1 FILLER_61_2440 ();
 sg13g2_fill_2 FILLER_61_2446 ();
 sg13g2_fill_1 FILLER_61_2448 ();
 sg13g2_fill_2 FILLER_61_2457 ();
 sg13g2_fill_1 FILLER_61_2459 ();
 sg13g2_fill_1 FILLER_61_2470 ();
 sg13g2_fill_2 FILLER_61_2476 ();
 sg13g2_fill_1 FILLER_61_2478 ();
 sg13g2_decap_4 FILLER_61_2482 ();
 sg13g2_decap_8 FILLER_61_2490 ();
 sg13g2_fill_1 FILLER_61_2497 ();
 sg13g2_fill_2 FILLER_61_2515 ();
 sg13g2_fill_1 FILLER_61_2517 ();
 sg13g2_fill_2 FILLER_61_2551 ();
 sg13g2_fill_1 FILLER_61_2553 ();
 sg13g2_fill_2 FILLER_61_2559 ();
 sg13g2_fill_2 FILLER_61_2569 ();
 sg13g2_fill_1 FILLER_61_2571 ();
 sg13g2_fill_2 FILLER_61_2580 ();
 sg13g2_fill_2 FILLER_61_2595 ();
 sg13g2_decap_8 FILLER_61_2625 ();
 sg13g2_decap_8 FILLER_61_2632 ();
 sg13g2_fill_2 FILLER_61_2662 ();
 sg13g2_fill_1 FILLER_61_2664 ();
 sg13g2_fill_2 FILLER_61_2686 ();
 sg13g2_decap_8 FILLER_61_2734 ();
 sg13g2_decap_4 FILLER_61_2741 ();
 sg13g2_fill_2 FILLER_61_2745 ();
 sg13g2_decap_4 FILLER_61_2751 ();
 sg13g2_fill_1 FILLER_61_2755 ();
 sg13g2_fill_2 FILLER_61_2773 ();
 sg13g2_fill_1 FILLER_61_2775 ();
 sg13g2_fill_2 FILLER_61_2790 ();
 sg13g2_fill_2 FILLER_61_2801 ();
 sg13g2_decap_8 FILLER_61_2821 ();
 sg13g2_decap_8 FILLER_61_2828 ();
 sg13g2_fill_2 FILLER_61_2843 ();
 sg13g2_decap_8 FILLER_61_2849 ();
 sg13g2_decap_4 FILLER_61_2856 ();
 sg13g2_fill_2 FILLER_61_2860 ();
 sg13g2_fill_1 FILLER_61_2871 ();
 sg13g2_fill_1 FILLER_61_2882 ();
 sg13g2_decap_8 FILLER_61_2908 ();
 sg13g2_fill_2 FILLER_61_2915 ();
 sg13g2_decap_4 FILLER_61_2925 ();
 sg13g2_fill_2 FILLER_61_2996 ();
 sg13g2_fill_1 FILLER_61_2998 ();
 sg13g2_fill_2 FILLER_61_3012 ();
 sg13g2_fill_1 FILLER_61_3014 ();
 sg13g2_decap_8 FILLER_61_3047 ();
 sg13g2_decap_4 FILLER_61_3054 ();
 sg13g2_fill_1 FILLER_61_3058 ();
 sg13g2_decap_4 FILLER_61_3085 ();
 sg13g2_fill_1 FILLER_61_3089 ();
 sg13g2_decap_4 FILLER_61_3103 ();
 sg13g2_fill_1 FILLER_61_3107 ();
 sg13g2_fill_2 FILLER_61_3113 ();
 sg13g2_decap_8 FILLER_61_3133 ();
 sg13g2_fill_1 FILLER_61_3155 ();
 sg13g2_decap_4 FILLER_61_3185 ();
 sg13g2_decap_4 FILLER_61_3193 ();
 sg13g2_fill_1 FILLER_61_3197 ();
 sg13g2_fill_2 FILLER_61_3224 ();
 sg13g2_decap_8 FILLER_61_3245 ();
 sg13g2_fill_2 FILLER_61_3263 ();
 sg13g2_fill_1 FILLER_61_3265 ();
 sg13g2_fill_1 FILLER_61_3305 ();
 sg13g2_fill_2 FILLER_61_3314 ();
 sg13g2_fill_1 FILLER_61_3316 ();
 sg13g2_decap_4 FILLER_61_3321 ();
 sg13g2_fill_1 FILLER_61_3331 ();
 sg13g2_decap_8 FILLER_61_3385 ();
 sg13g2_decap_8 FILLER_61_3396 ();
 sg13g2_decap_4 FILLER_61_3403 ();
 sg13g2_fill_2 FILLER_61_3407 ();
 sg13g2_fill_1 FILLER_61_3437 ();
 sg13g2_decap_8 FILLER_61_3454 ();
 sg13g2_decap_4 FILLER_61_3461 ();
 sg13g2_decap_8 FILLER_61_3478 ();
 sg13g2_fill_1 FILLER_61_3489 ();
 sg13g2_fill_1 FILLER_61_3517 ();
 sg13g2_decap_8 FILLER_61_3529 ();
 sg13g2_fill_2 FILLER_61_3536 ();
 sg13g2_decap_8 FILLER_61_3546 ();
 sg13g2_decap_4 FILLER_61_3553 ();
 sg13g2_fill_1 FILLER_61_3557 ();
 sg13g2_decap_8 FILLER_61_3573 ();
 sg13g2_decap_4 FILLER_62_0 ();
 sg13g2_fill_2 FILLER_62_4 ();
 sg13g2_fill_2 FILLER_62_10 ();
 sg13g2_decap_4 FILLER_62_54 ();
 sg13g2_fill_2 FILLER_62_58 ();
 sg13g2_fill_2 FILLER_62_68 ();
 sg13g2_fill_2 FILLER_62_75 ();
 sg13g2_decap_8 FILLER_62_103 ();
 sg13g2_fill_2 FILLER_62_128 ();
 sg13g2_fill_1 FILLER_62_130 ();
 sg13g2_fill_2 FILLER_62_220 ();
 sg13g2_fill_2 FILLER_62_239 ();
 sg13g2_fill_2 FILLER_62_311 ();
 sg13g2_fill_2 FILLER_62_328 ();
 sg13g2_fill_2 FILLER_62_354 ();
 sg13g2_decap_8 FILLER_62_377 ();
 sg13g2_fill_1 FILLER_62_384 ();
 sg13g2_fill_2 FILLER_62_390 ();
 sg13g2_fill_2 FILLER_62_409 ();
 sg13g2_fill_1 FILLER_62_411 ();
 sg13g2_fill_1 FILLER_62_428 ();
 sg13g2_fill_2 FILLER_62_475 ();
 sg13g2_fill_2 FILLER_62_481 ();
 sg13g2_fill_1 FILLER_62_483 ();
 sg13g2_fill_1 FILLER_62_501 ();
 sg13g2_fill_2 FILLER_62_535 ();
 sg13g2_fill_1 FILLER_62_550 ();
 sg13g2_fill_2 FILLER_62_571 ();
 sg13g2_fill_2 FILLER_62_581 ();
 sg13g2_decap_8 FILLER_62_592 ();
 sg13g2_decap_4 FILLER_62_599 ();
 sg13g2_fill_1 FILLER_62_603 ();
 sg13g2_decap_8 FILLER_62_618 ();
 sg13g2_decap_8 FILLER_62_625 ();
 sg13g2_fill_2 FILLER_62_632 ();
 sg13g2_fill_2 FILLER_62_664 ();
 sg13g2_fill_2 FILLER_62_698 ();
 sg13g2_decap_4 FILLER_62_729 ();
 sg13g2_fill_1 FILLER_62_733 ();
 sg13g2_decap_8 FILLER_62_750 ();
 sg13g2_fill_2 FILLER_62_757 ();
 sg13g2_fill_1 FILLER_62_759 ();
 sg13g2_fill_1 FILLER_62_797 ();
 sg13g2_decap_4 FILLER_62_822 ();
 sg13g2_fill_2 FILLER_62_826 ();
 sg13g2_decap_4 FILLER_62_849 ();
 sg13g2_fill_2 FILLER_62_853 ();
 sg13g2_fill_2 FILLER_62_860 ();
 sg13g2_decap_4 FILLER_62_884 ();
 sg13g2_fill_2 FILLER_62_893 ();
 sg13g2_fill_1 FILLER_62_895 ();
 sg13g2_fill_2 FILLER_62_904 ();
 sg13g2_fill_1 FILLER_62_980 ();
 sg13g2_fill_2 FILLER_62_1006 ();
 sg13g2_fill_1 FILLER_62_1008 ();
 sg13g2_fill_1 FILLER_62_1026 ();
 sg13g2_fill_2 FILLER_62_1040 ();
 sg13g2_decap_4 FILLER_62_1072 ();
 sg13g2_fill_2 FILLER_62_1076 ();
 sg13g2_fill_2 FILLER_62_1086 ();
 sg13g2_fill_1 FILLER_62_1088 ();
 sg13g2_fill_1 FILLER_62_1093 ();
 sg13g2_fill_2 FILLER_62_1104 ();
 sg13g2_fill_2 FILLER_62_1120 ();
 sg13g2_fill_1 FILLER_62_1122 ();
 sg13g2_fill_1 FILLER_62_1129 ();
 sg13g2_decap_8 FILLER_62_1143 ();
 sg13g2_decap_8 FILLER_62_1150 ();
 sg13g2_decap_4 FILLER_62_1157 ();
 sg13g2_fill_2 FILLER_62_1161 ();
 sg13g2_fill_1 FILLER_62_1174 ();
 sg13g2_decap_8 FILLER_62_1200 ();
 sg13g2_decap_4 FILLER_62_1207 ();
 sg13g2_decap_4 FILLER_62_1241 ();
 sg13g2_fill_2 FILLER_62_1245 ();
 sg13g2_decap_4 FILLER_62_1251 ();
 sg13g2_decap_4 FILLER_62_1259 ();
 sg13g2_fill_2 FILLER_62_1263 ();
 sg13g2_fill_2 FILLER_62_1293 ();
 sg13g2_fill_2 FILLER_62_1336 ();
 sg13g2_fill_1 FILLER_62_1338 ();
 sg13g2_fill_2 FILLER_62_1347 ();
 sg13g2_decap_4 FILLER_62_1373 ();
 sg13g2_fill_2 FILLER_62_1377 ();
 sg13g2_decap_4 FILLER_62_1393 ();
 sg13g2_fill_2 FILLER_62_1397 ();
 sg13g2_fill_2 FILLER_62_1406 ();
 sg13g2_fill_1 FILLER_62_1440 ();
 sg13g2_fill_2 FILLER_62_1456 ();
 sg13g2_decap_8 FILLER_62_1472 ();
 sg13g2_fill_1 FILLER_62_1479 ();
 sg13g2_fill_2 FILLER_62_1497 ();
 sg13g2_decap_8 FILLER_62_1509 ();
 sg13g2_fill_2 FILLER_62_1516 ();
 sg13g2_fill_1 FILLER_62_1518 ();
 sg13g2_fill_2 FILLER_62_1532 ();
 sg13g2_decap_8 FILLER_62_1542 ();
 sg13g2_fill_1 FILLER_62_1563 ();
 sg13g2_decap_8 FILLER_62_1586 ();
 sg13g2_fill_1 FILLER_62_1593 ();
 sg13g2_fill_1 FILLER_62_1607 ();
 sg13g2_fill_2 FILLER_62_1618 ();
 sg13g2_fill_1 FILLER_62_1620 ();
 sg13g2_decap_8 FILLER_62_1625 ();
 sg13g2_fill_2 FILLER_62_1665 ();
 sg13g2_fill_1 FILLER_62_1667 ();
 sg13g2_fill_2 FILLER_62_1681 ();
 sg13g2_decap_8 FILLER_62_1688 ();
 sg13g2_fill_2 FILLER_62_1695 ();
 sg13g2_fill_1 FILLER_62_1697 ();
 sg13g2_fill_2 FILLER_62_1713 ();
 sg13g2_fill_2 FILLER_62_1748 ();
 sg13g2_fill_1 FILLER_62_1750 ();
 sg13g2_fill_2 FILLER_62_1765 ();
 sg13g2_decap_4 FILLER_62_1787 ();
 sg13g2_fill_1 FILLER_62_1791 ();
 sg13g2_fill_1 FILLER_62_1797 ();
 sg13g2_decap_8 FILLER_62_1806 ();
 sg13g2_fill_2 FILLER_62_1821 ();
 sg13g2_decap_4 FILLER_62_1857 ();
 sg13g2_fill_2 FILLER_62_1877 ();
 sg13g2_decap_8 FILLER_62_1883 ();
 sg13g2_fill_2 FILLER_62_1890 ();
 sg13g2_fill_1 FILLER_62_1905 ();
 sg13g2_fill_2 FILLER_62_1917 ();
 sg13g2_decap_4 FILLER_62_1937 ();
 sg13g2_fill_2 FILLER_62_1945 ();
 sg13g2_fill_1 FILLER_62_1947 ();
 sg13g2_fill_2 FILLER_62_1961 ();
 sg13g2_fill_1 FILLER_62_2017 ();
 sg13g2_decap_4 FILLER_62_2043 ();
 sg13g2_fill_1 FILLER_62_2047 ();
 sg13g2_decap_4 FILLER_62_2053 ();
 sg13g2_fill_2 FILLER_62_2062 ();
 sg13g2_fill_1 FILLER_62_2124 ();
 sg13g2_fill_2 FILLER_62_2133 ();
 sg13g2_decap_4 FILLER_62_2143 ();
 sg13g2_decap_4 FILLER_62_2159 ();
 sg13g2_fill_1 FILLER_62_2163 ();
 sg13g2_fill_2 FILLER_62_2168 ();
 sg13g2_fill_1 FILLER_62_2194 ();
 sg13g2_decap_8 FILLER_62_2210 ();
 sg13g2_fill_1 FILLER_62_2232 ();
 sg13g2_fill_2 FILLER_62_2253 ();
 sg13g2_fill_1 FILLER_62_2255 ();
 sg13g2_decap_8 FILLER_62_2334 ();
 sg13g2_decap_4 FILLER_62_2345 ();
 sg13g2_fill_2 FILLER_62_2349 ();
 sg13g2_decap_4 FILLER_62_2398 ();
 sg13g2_fill_2 FILLER_62_2402 ();
 sg13g2_decap_8 FILLER_62_2431 ();
 sg13g2_fill_1 FILLER_62_2438 ();
 sg13g2_fill_2 FILLER_62_2464 ();
 sg13g2_fill_1 FILLER_62_2466 ();
 sg13g2_fill_1 FILLER_62_2487 ();
 sg13g2_fill_1 FILLER_62_2497 ();
 sg13g2_decap_8 FILLER_62_2501 ();
 sg13g2_decap_4 FILLER_62_2511 ();
 sg13g2_decap_4 FILLER_62_2536 ();
 sg13g2_fill_1 FILLER_62_2540 ();
 sg13g2_decap_8 FILLER_62_2553 ();
 sg13g2_fill_2 FILLER_62_2560 ();
 sg13g2_fill_2 FILLER_62_2565 ();
 sg13g2_fill_2 FILLER_62_2609 ();
 sg13g2_decap_8 FILLER_62_2634 ();
 sg13g2_decap_8 FILLER_62_2662 ();
 sg13g2_decap_8 FILLER_62_2669 ();
 sg13g2_fill_1 FILLER_62_2676 ();
 sg13g2_decap_4 FILLER_62_2687 ();
 sg13g2_fill_1 FILLER_62_2699 ();
 sg13g2_fill_2 FILLER_62_2705 ();
 sg13g2_fill_1 FILLER_62_2715 ();
 sg13g2_fill_2 FILLER_62_2770 ();
 sg13g2_fill_1 FILLER_62_2772 ();
 sg13g2_decap_4 FILLER_62_2785 ();
 sg13g2_fill_2 FILLER_62_2789 ();
 sg13g2_fill_2 FILLER_62_2803 ();
 sg13g2_fill_1 FILLER_62_2805 ();
 sg13g2_decap_4 FILLER_62_2821 ();
 sg13g2_fill_2 FILLER_62_2825 ();
 sg13g2_fill_1 FILLER_62_2868 ();
 sg13g2_decap_4 FILLER_62_2899 ();
 sg13g2_fill_2 FILLER_62_2903 ();
 sg13g2_fill_2 FILLER_62_2937 ();
 sg13g2_fill_1 FILLER_62_2939 ();
 sg13g2_decap_4 FILLER_62_2945 ();
 sg13g2_fill_2 FILLER_62_2949 ();
 sg13g2_decap_8 FILLER_62_2968 ();
 sg13g2_decap_4 FILLER_62_2975 ();
 sg13g2_decap_4 FILLER_62_2992 ();
 sg13g2_fill_2 FILLER_62_2996 ();
 sg13g2_decap_4 FILLER_62_3026 ();
 sg13g2_fill_2 FILLER_62_3030 ();
 sg13g2_decap_4 FILLER_62_3037 ();
 sg13g2_fill_1 FILLER_62_3041 ();
 sg13g2_fill_2 FILLER_62_3068 ();
 sg13g2_fill_1 FILLER_62_3070 ();
 sg13g2_fill_2 FILLER_62_3081 ();
 sg13g2_fill_1 FILLER_62_3083 ();
 sg13g2_decap_4 FILLER_62_3088 ();
 sg13g2_decap_4 FILLER_62_3102 ();
 sg13g2_fill_1 FILLER_62_3132 ();
 sg13g2_fill_2 FILLER_62_3155 ();
 sg13g2_fill_1 FILLER_62_3161 ();
 sg13g2_fill_2 FILLER_62_3183 ();
 sg13g2_fill_2 FILLER_62_3201 ();
 sg13g2_decap_4 FILLER_62_3239 ();
 sg13g2_fill_1 FILLER_62_3243 ();
 sg13g2_fill_1 FILLER_62_3262 ();
 sg13g2_decap_4 FILLER_62_3267 ();
 sg13g2_fill_1 FILLER_62_3274 ();
 sg13g2_fill_1 FILLER_62_3288 ();
 sg13g2_decap_4 FILLER_62_3294 ();
 sg13g2_decap_8 FILLER_62_3333 ();
 sg13g2_fill_1 FILLER_62_3340 ();
 sg13g2_fill_2 FILLER_62_3356 ();
 sg13g2_fill_1 FILLER_62_3376 ();
 sg13g2_fill_2 FILLER_62_3404 ();
 sg13g2_fill_2 FILLER_62_3437 ();
 sg13g2_decap_4 FILLER_62_3448 ();
 sg13g2_fill_1 FILLER_62_3452 ();
 sg13g2_decap_8 FILLER_62_3467 ();
 sg13g2_fill_2 FILLER_62_3474 ();
 sg13g2_fill_2 FILLER_62_3502 ();
 sg13g2_decap_4 FILLER_62_3509 ();
 sg13g2_fill_2 FILLER_62_3513 ();
 sg13g2_fill_2 FILLER_62_3549 ();
 sg13g2_decap_4 FILLER_62_3574 ();
 sg13g2_fill_2 FILLER_62_3578 ();
 sg13g2_decap_4 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_32 ();
 sg13g2_fill_2 FILLER_63_51 ();
 sg13g2_decap_4 FILLER_63_71 ();
 sg13g2_fill_1 FILLER_63_75 ();
 sg13g2_decap_4 FILLER_63_96 ();
 sg13g2_fill_1 FILLER_63_100 ();
 sg13g2_fill_1 FILLER_63_171 ();
 sg13g2_fill_2 FILLER_63_216 ();
 sg13g2_fill_1 FILLER_63_218 ();
 sg13g2_fill_1 FILLER_63_245 ();
 sg13g2_fill_1 FILLER_63_271 ();
 sg13g2_fill_1 FILLER_63_277 ();
 sg13g2_fill_2 FILLER_63_333 ();
 sg13g2_fill_1 FILLER_63_340 ();
 sg13g2_fill_1 FILLER_63_346 ();
 sg13g2_decap_8 FILLER_63_352 ();
 sg13g2_decap_8 FILLER_63_359 ();
 sg13g2_fill_2 FILLER_63_366 ();
 sg13g2_decap_8 FILLER_63_378 ();
 sg13g2_fill_2 FILLER_63_385 ();
 sg13g2_decap_4 FILLER_63_412 ();
 sg13g2_fill_1 FILLER_63_416 ();
 sg13g2_fill_2 FILLER_63_435 ();
 sg13g2_decap_8 FILLER_63_446 ();
 sg13g2_fill_2 FILLER_63_453 ();
 sg13g2_decap_4 FILLER_63_462 ();
 sg13g2_decap_8 FILLER_63_479 ();
 sg13g2_fill_2 FILLER_63_486 ();
 sg13g2_fill_1 FILLER_63_488 ();
 sg13g2_fill_1 FILLER_63_507 ();
 sg13g2_decap_4 FILLER_63_549 ();
 sg13g2_fill_2 FILLER_63_553 ();
 sg13g2_decap_8 FILLER_63_568 ();
 sg13g2_fill_2 FILLER_63_575 ();
 sg13g2_fill_1 FILLER_63_577 ();
 sg13g2_decap_4 FILLER_63_589 ();
 sg13g2_decap_4 FILLER_63_598 ();
 sg13g2_fill_1 FILLER_63_602 ();
 sg13g2_decap_8 FILLER_63_620 ();
 sg13g2_fill_2 FILLER_63_627 ();
 sg13g2_fill_1 FILLER_63_629 ();
 sg13g2_decap_4 FILLER_63_668 ();
 sg13g2_fill_2 FILLER_63_676 ();
 sg13g2_fill_1 FILLER_63_678 ();
 sg13g2_decap_8 FILLER_63_696 ();
 sg13g2_fill_2 FILLER_63_703 ();
 sg13g2_decap_8 FILLER_63_717 ();
 sg13g2_decap_8 FILLER_63_724 ();
 sg13g2_decap_4 FILLER_63_731 ();
 sg13g2_fill_1 FILLER_63_735 ();
 sg13g2_fill_2 FILLER_63_761 ();
 sg13g2_fill_1 FILLER_63_763 ();
 sg13g2_decap_4 FILLER_63_874 ();
 sg13g2_fill_2 FILLER_63_878 ();
 sg13g2_fill_2 FILLER_63_893 ();
 sg13g2_fill_1 FILLER_63_895 ();
 sg13g2_fill_2 FILLER_63_913 ();
 sg13g2_decap_4 FILLER_63_932 ();
 sg13g2_fill_2 FILLER_63_993 ();
 sg13g2_fill_2 FILLER_63_1003 ();
 sg13g2_fill_2 FILLER_63_1021 ();
 sg13g2_fill_1 FILLER_63_1044 ();
 sg13g2_decap_4 FILLER_63_1066 ();
 sg13g2_fill_1 FILLER_63_1070 ();
 sg13g2_fill_2 FILLER_63_1092 ();
 sg13g2_fill_1 FILLER_63_1094 ();
 sg13g2_fill_1 FILLER_63_1121 ();
 sg13g2_fill_2 FILLER_63_1146 ();
 sg13g2_fill_2 FILLER_63_1180 ();
 sg13g2_fill_1 FILLER_63_1182 ();
 sg13g2_fill_2 FILLER_63_1192 ();
 sg13g2_fill_1 FILLER_63_1194 ();
 sg13g2_fill_2 FILLER_63_1200 ();
 sg13g2_fill_2 FILLER_63_1215 ();
 sg13g2_fill_2 FILLER_63_1234 ();
 sg13g2_decap_8 FILLER_63_1256 ();
 sg13g2_decap_4 FILLER_63_1263 ();
 sg13g2_fill_2 FILLER_63_1302 ();
 sg13g2_fill_2 FILLER_63_1309 ();
 sg13g2_fill_1 FILLER_63_1311 ();
 sg13g2_fill_1 FILLER_63_1347 ();
 sg13g2_fill_1 FILLER_63_1357 ();
 sg13g2_fill_1 FILLER_63_1399 ();
 sg13g2_fill_2 FILLER_63_1428 ();
 sg13g2_decap_4 FILLER_63_1438 ();
 sg13g2_decap_4 FILLER_63_1478 ();
 sg13g2_decap_4 FILLER_63_1508 ();
 sg13g2_decap_8 FILLER_63_1531 ();
 sg13g2_decap_4 FILLER_63_1538 ();
 sg13g2_fill_2 FILLER_63_1542 ();
 sg13g2_fill_1 FILLER_63_1557 ();
 sg13g2_decap_8 FILLER_63_1612 ();
 sg13g2_fill_1 FILLER_63_1619 ();
 sg13g2_fill_1 FILLER_63_1633 ();
 sg13g2_fill_2 FILLER_63_1647 ();
 sg13g2_decap_4 FILLER_63_1659 ();
 sg13g2_fill_1 FILLER_63_1663 ();
 sg13g2_fill_1 FILLER_63_1692 ();
 sg13g2_decap_8 FILLER_63_1707 ();
 sg13g2_decap_8 FILLER_63_1714 ();
 sg13g2_fill_1 FILLER_63_1721 ();
 sg13g2_decap_8 FILLER_63_1735 ();
 sg13g2_decap_4 FILLER_63_1747 ();
 sg13g2_fill_1 FILLER_63_1751 ();
 sg13g2_decap_4 FILLER_63_1757 ();
 sg13g2_fill_2 FILLER_63_1761 ();
 sg13g2_fill_2 FILLER_63_1772 ();
 sg13g2_fill_1 FILLER_63_1774 ();
 sg13g2_fill_1 FILLER_63_1789 ();
 sg13g2_decap_8 FILLER_63_1810 ();
 sg13g2_decap_4 FILLER_63_1817 ();
 sg13g2_fill_1 FILLER_63_1821 ();
 sg13g2_decap_4 FILLER_63_1829 ();
 sg13g2_fill_2 FILLER_63_1833 ();
 sg13g2_fill_1 FILLER_63_1840 ();
 sg13g2_fill_2 FILLER_63_1846 ();
 sg13g2_fill_1 FILLER_63_1848 ();
 sg13g2_fill_2 FILLER_63_1859 ();
 sg13g2_fill_1 FILLER_63_1861 ();
 sg13g2_fill_1 FILLER_63_1890 ();
 sg13g2_fill_2 FILLER_63_1910 ();
 sg13g2_fill_2 FILLER_63_1924 ();
 sg13g2_fill_1 FILLER_63_1926 ();
 sg13g2_decap_8 FILLER_63_1967 ();
 sg13g2_decap_8 FILLER_63_1974 ();
 sg13g2_decap_8 FILLER_63_1981 ();
 sg13g2_fill_1 FILLER_63_1988 ();
 sg13g2_fill_2 FILLER_63_2007 ();
 sg13g2_fill_1 FILLER_63_2013 ();
 sg13g2_fill_1 FILLER_63_2018 ();
 sg13g2_decap_4 FILLER_63_2038 ();
 sg13g2_fill_1 FILLER_63_2081 ();
 sg13g2_fill_2 FILLER_63_2092 ();
 sg13g2_fill_1 FILLER_63_2094 ();
 sg13g2_fill_2 FILLER_63_2118 ();
 sg13g2_fill_1 FILLER_63_2130 ();
 sg13g2_fill_2 FILLER_63_2157 ();
 sg13g2_fill_2 FILLER_63_2183 ();
 sg13g2_fill_1 FILLER_63_2185 ();
 sg13g2_decap_4 FILLER_63_2191 ();
 sg13g2_decap_8 FILLER_63_2208 ();
 sg13g2_fill_2 FILLER_63_2215 ();
 sg13g2_fill_1 FILLER_63_2217 ();
 sg13g2_decap_4 FILLER_63_2231 ();
 sg13g2_fill_1 FILLER_63_2235 ();
 sg13g2_decap_8 FILLER_63_2252 ();
 sg13g2_decap_8 FILLER_63_2273 ();
 sg13g2_decap_8 FILLER_63_2284 ();
 sg13g2_decap_4 FILLER_63_2291 ();
 sg13g2_fill_1 FILLER_63_2308 ();
 sg13g2_fill_2 FILLER_63_2321 ();
 sg13g2_fill_1 FILLER_63_2356 ();
 sg13g2_fill_2 FILLER_63_2369 ();
 sg13g2_fill_1 FILLER_63_2384 ();
 sg13g2_decap_8 FILLER_63_2397 ();
 sg13g2_decap_8 FILLER_63_2404 ();
 sg13g2_decap_4 FILLER_63_2411 ();
 sg13g2_fill_2 FILLER_63_2420 ();
 sg13g2_decap_8 FILLER_63_2435 ();
 sg13g2_decap_4 FILLER_63_2442 ();
 sg13g2_fill_1 FILLER_63_2446 ();
 sg13g2_fill_1 FILLER_63_2466 ();
 sg13g2_fill_2 FILLER_63_2476 ();
 sg13g2_fill_1 FILLER_63_2478 ();
 sg13g2_fill_2 FILLER_63_2497 ();
 sg13g2_fill_1 FILLER_63_2499 ();
 sg13g2_fill_2 FILLER_63_2520 ();
 sg13g2_fill_1 FILLER_63_2522 ();
 sg13g2_fill_2 FILLER_63_2546 ();
 sg13g2_fill_1 FILLER_63_2548 ();
 sg13g2_fill_1 FILLER_63_2554 ();
 sg13g2_fill_1 FILLER_63_2561 ();
 sg13g2_decap_8 FILLER_63_2575 ();
 sg13g2_fill_2 FILLER_63_2647 ();
 sg13g2_fill_1 FILLER_63_2649 ();
 sg13g2_decap_8 FILLER_63_2667 ();
 sg13g2_fill_2 FILLER_63_2674 ();
 sg13g2_fill_1 FILLER_63_2676 ();
 sg13g2_fill_2 FILLER_63_2681 ();
 sg13g2_fill_2 FILLER_63_2697 ();
 sg13g2_fill_1 FILLER_63_2699 ();
 sg13g2_fill_2 FILLER_63_2716 ();
 sg13g2_fill_2 FILLER_63_2731 ();
 sg13g2_decap_8 FILLER_63_2746 ();
 sg13g2_decap_8 FILLER_63_2753 ();
 sg13g2_fill_2 FILLER_63_2760 ();
 sg13g2_decap_4 FILLER_63_2792 ();
 sg13g2_fill_2 FILLER_63_2796 ();
 sg13g2_decap_8 FILLER_63_2807 ();
 sg13g2_fill_2 FILLER_63_2814 ();
 sg13g2_fill_1 FILLER_63_2816 ();
 sg13g2_decap_4 FILLER_63_2831 ();
 sg13g2_fill_2 FILLER_63_2849 ();
 sg13g2_fill_1 FILLER_63_2856 ();
 sg13g2_fill_1 FILLER_63_2956 ();
 sg13g2_fill_2 FILLER_63_2967 ();
 sg13g2_fill_1 FILLER_63_2969 ();
 sg13g2_fill_2 FILLER_63_2980 ();
 sg13g2_decap_8 FILLER_63_2992 ();
 sg13g2_decap_8 FILLER_63_3014 ();
 sg13g2_fill_2 FILLER_63_3029 ();
 sg13g2_fill_1 FILLER_63_3059 ();
 sg13g2_fill_2 FILLER_63_3070 ();
 sg13g2_fill_1 FILLER_63_3072 ();
 sg13g2_fill_2 FILLER_63_3086 ();
 sg13g2_decap_8 FILLER_63_3096 ();
 sg13g2_fill_2 FILLER_63_3103 ();
 sg13g2_fill_1 FILLER_63_3105 ();
 sg13g2_decap_4 FILLER_63_3128 ();
 sg13g2_fill_2 FILLER_63_3132 ();
 sg13g2_fill_2 FILLER_63_3156 ();
 sg13g2_fill_1 FILLER_63_3158 ();
 sg13g2_decap_8 FILLER_63_3176 ();
 sg13g2_decap_8 FILLER_63_3183 ();
 sg13g2_fill_1 FILLER_63_3190 ();
 sg13g2_fill_2 FILLER_63_3200 ();
 sg13g2_decap_8 FILLER_63_3211 ();
 sg13g2_fill_1 FILLER_63_3218 ();
 sg13g2_fill_1 FILLER_63_3223 ();
 sg13g2_fill_2 FILLER_63_3241 ();
 sg13g2_fill_1 FILLER_63_3243 ();
 sg13g2_fill_2 FILLER_63_3261 ();
 sg13g2_fill_1 FILLER_63_3288 ();
 sg13g2_fill_2 FILLER_63_3315 ();
 sg13g2_fill_2 FILLER_63_3325 ();
 sg13g2_fill_2 FILLER_63_3370 ();
 sg13g2_decap_8 FILLER_63_3400 ();
 sg13g2_decap_4 FILLER_63_3407 ();
 sg13g2_fill_2 FILLER_63_3424 ();
 sg13g2_fill_1 FILLER_63_3426 ();
 sg13g2_fill_2 FILLER_63_3435 ();
 sg13g2_fill_1 FILLER_63_3445 ();
 sg13g2_fill_1 FILLER_63_3467 ();
 sg13g2_fill_2 FILLER_63_3482 ();
 sg13g2_fill_1 FILLER_63_3484 ();
 sg13g2_fill_1 FILLER_63_3514 ();
 sg13g2_fill_1 FILLER_63_3562 ();
 sg13g2_fill_2 FILLER_63_3577 ();
 sg13g2_fill_1 FILLER_63_3579 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_7 ();
 sg13g2_fill_1 FILLER_64_48 ();
 sg13g2_decap_4 FILLER_64_69 ();
 sg13g2_fill_2 FILLER_64_73 ();
 sg13g2_fill_2 FILLER_64_96 ();
 sg13g2_fill_1 FILLER_64_98 ();
 sg13g2_fill_1 FILLER_64_116 ();
 sg13g2_fill_2 FILLER_64_130 ();
 sg13g2_fill_1 FILLER_64_150 ();
 sg13g2_fill_1 FILLER_64_184 ();
 sg13g2_fill_1 FILLER_64_267 ();
 sg13g2_decap_8 FILLER_64_301 ();
 sg13g2_fill_2 FILLER_64_308 ();
 sg13g2_decap_8 FILLER_64_315 ();
 sg13g2_fill_2 FILLER_64_322 ();
 sg13g2_fill_1 FILLER_64_324 ();
 sg13g2_fill_2 FILLER_64_359 ();
 sg13g2_decap_4 FILLER_64_377 ();
 sg13g2_fill_2 FILLER_64_381 ();
 sg13g2_fill_1 FILLER_64_394 ();
 sg13g2_decap_4 FILLER_64_418 ();
 sg13g2_fill_1 FILLER_64_422 ();
 sg13g2_fill_2 FILLER_64_439 ();
 sg13g2_decap_8 FILLER_64_451 ();
 sg13g2_fill_2 FILLER_64_458 ();
 sg13g2_fill_2 FILLER_64_483 ();
 sg13g2_fill_1 FILLER_64_485 ();
 sg13g2_fill_2 FILLER_64_494 ();
 sg13g2_fill_1 FILLER_64_507 ();
 sg13g2_fill_1 FILLER_64_517 ();
 sg13g2_fill_2 FILLER_64_527 ();
 sg13g2_fill_2 FILLER_64_546 ();
 sg13g2_fill_2 FILLER_64_565 ();
 sg13g2_fill_2 FILLER_64_576 ();
 sg13g2_fill_1 FILLER_64_578 ();
 sg13g2_decap_4 FILLER_64_612 ();
 sg13g2_decap_4 FILLER_64_629 ();
 sg13g2_fill_2 FILLER_64_646 ();
 sg13g2_fill_1 FILLER_64_648 ();
 sg13g2_decap_4 FILLER_64_654 ();
 sg13g2_decap_8 FILLER_64_666 ();
 sg13g2_decap_8 FILLER_64_673 ();
 sg13g2_fill_1 FILLER_64_680 ();
 sg13g2_decap_8 FILLER_64_685 ();
 sg13g2_decap_8 FILLER_64_692 ();
 sg13g2_decap_4 FILLER_64_699 ();
 sg13g2_decap_4 FILLER_64_742 ();
 sg13g2_fill_1 FILLER_64_746 ();
 sg13g2_decap_8 FILLER_64_752 ();
 sg13g2_fill_2 FILLER_64_759 ();
 sg13g2_decap_4 FILLER_64_787 ();
 sg13g2_fill_1 FILLER_64_791 ();
 sg13g2_decap_8 FILLER_64_809 ();
 sg13g2_decap_8 FILLER_64_816 ();
 sg13g2_fill_1 FILLER_64_823 ();
 sg13g2_decap_4 FILLER_64_828 ();
 sg13g2_fill_1 FILLER_64_832 ();
 sg13g2_decap_8 FILLER_64_841 ();
 sg13g2_decap_8 FILLER_64_848 ();
 sg13g2_fill_2 FILLER_64_855 ();
 sg13g2_decap_4 FILLER_64_883 ();
 sg13g2_fill_1 FILLER_64_887 ();
 sg13g2_fill_2 FILLER_64_918 ();
 sg13g2_fill_1 FILLER_64_920 ();
 sg13g2_fill_2 FILLER_64_975 ();
 sg13g2_decap_8 FILLER_64_998 ();
 sg13g2_fill_1 FILLER_64_1031 ();
 sg13g2_decap_4 FILLER_64_1043 ();
 sg13g2_fill_2 FILLER_64_1047 ();
 sg13g2_decap_4 FILLER_64_1052 ();
 sg13g2_fill_2 FILLER_64_1056 ();
 sg13g2_decap_8 FILLER_64_1069 ();
 sg13g2_fill_2 FILLER_64_1076 ();
 sg13g2_decap_8 FILLER_64_1086 ();
 sg13g2_decap_4 FILLER_64_1093 ();
 sg13g2_fill_1 FILLER_64_1097 ();
 sg13g2_fill_1 FILLER_64_1124 ();
 sg13g2_fill_1 FILLER_64_1138 ();
 sg13g2_decap_4 FILLER_64_1145 ();
 sg13g2_fill_2 FILLER_64_1149 ();
 sg13g2_decap_8 FILLER_64_1171 ();
 sg13g2_fill_1 FILLER_64_1178 ();
 sg13g2_decap_4 FILLER_64_1205 ();
 sg13g2_fill_2 FILLER_64_1209 ();
 sg13g2_fill_2 FILLER_64_1233 ();
 sg13g2_fill_2 FILLER_64_1267 ();
 sg13g2_fill_2 FILLER_64_1290 ();
 sg13g2_fill_1 FILLER_64_1292 ();
 sg13g2_fill_2 FILLER_64_1298 ();
 sg13g2_fill_2 FILLER_64_1312 ();
 sg13g2_fill_1 FILLER_64_1314 ();
 sg13g2_fill_2 FILLER_64_1336 ();
 sg13g2_fill_1 FILLER_64_1338 ();
 sg13g2_decap_8 FILLER_64_1389 ();
 sg13g2_decap_4 FILLER_64_1401 ();
 sg13g2_decap_8 FILLER_64_1409 ();
 sg13g2_decap_8 FILLER_64_1416 ();
 sg13g2_fill_1 FILLER_64_1423 ();
 sg13g2_decap_8 FILLER_64_1428 ();
 sg13g2_fill_2 FILLER_64_1435 ();
 sg13g2_fill_1 FILLER_64_1437 ();
 sg13g2_decap_8 FILLER_64_1451 ();
 sg13g2_decap_4 FILLER_64_1458 ();
 sg13g2_fill_1 FILLER_64_1471 ();
 sg13g2_decap_4 FILLER_64_1485 ();
 sg13g2_fill_2 FILLER_64_1499 ();
 sg13g2_fill_1 FILLER_64_1501 ();
 sg13g2_decap_4 FILLER_64_1530 ();
 sg13g2_fill_1 FILLER_64_1534 ();
 sg13g2_fill_2 FILLER_64_1576 ();
 sg13g2_fill_1 FILLER_64_1578 ();
 sg13g2_fill_2 FILLER_64_1588 ();
 sg13g2_fill_1 FILLER_64_1590 ();
 sg13g2_decap_4 FILLER_64_1613 ();
 sg13g2_fill_1 FILLER_64_1617 ();
 sg13g2_fill_2 FILLER_64_1662 ();
 sg13g2_fill_1 FILLER_64_1678 ();
 sg13g2_fill_2 FILLER_64_1694 ();
 sg13g2_fill_1 FILLER_64_1696 ();
 sg13g2_decap_4 FILLER_64_1710 ();
 sg13g2_fill_1 FILLER_64_1714 ();
 sg13g2_fill_2 FILLER_64_1724 ();
 sg13g2_fill_1 FILLER_64_1726 ();
 sg13g2_fill_2 FILLER_64_1735 ();
 sg13g2_decap_8 FILLER_64_1752 ();
 sg13g2_decap_4 FILLER_64_1759 ();
 sg13g2_fill_1 FILLER_64_1763 ();
 sg13g2_fill_1 FILLER_64_1769 ();
 sg13g2_decap_8 FILLER_64_1775 ();
 sg13g2_fill_2 FILLER_64_1782 ();
 sg13g2_fill_1 FILLER_64_1784 ();
 sg13g2_fill_2 FILLER_64_1794 ();
 sg13g2_decap_8 FILLER_64_1802 ();
 sg13g2_decap_4 FILLER_64_1809 ();
 sg13g2_fill_2 FILLER_64_1813 ();
 sg13g2_fill_2 FILLER_64_1846 ();
 sg13g2_decap_4 FILLER_64_1853 ();
 sg13g2_fill_1 FILLER_64_1887 ();
 sg13g2_fill_1 FILLER_64_1897 ();
 sg13g2_fill_1 FILLER_64_1906 ();
 sg13g2_fill_1 FILLER_64_1912 ();
 sg13g2_fill_1 FILLER_64_1928 ();
 sg13g2_fill_1 FILLER_64_1944 ();
 sg13g2_fill_2 FILLER_64_1950 ();
 sg13g2_decap_8 FILLER_64_1973 ();
 sg13g2_fill_1 FILLER_64_1980 ();
 sg13g2_decap_4 FILLER_64_1985 ();
 sg13g2_fill_2 FILLER_64_1989 ();
 sg13g2_fill_2 FILLER_64_2014 ();
 sg13g2_fill_1 FILLER_64_2016 ();
 sg13g2_fill_1 FILLER_64_2022 ();
 sg13g2_decap_4 FILLER_64_2033 ();
 sg13g2_decap_8 FILLER_64_2047 ();
 sg13g2_fill_1 FILLER_64_2054 ();
 sg13g2_fill_2 FILLER_64_2067 ();
 sg13g2_fill_1 FILLER_64_2069 ();
 sg13g2_fill_2 FILLER_64_2074 ();
 sg13g2_decap_8 FILLER_64_2089 ();
 sg13g2_fill_2 FILLER_64_2096 ();
 sg13g2_fill_1 FILLER_64_2098 ();
 sg13g2_fill_2 FILLER_64_2120 ();
 sg13g2_fill_2 FILLER_64_2135 ();
 sg13g2_fill_1 FILLER_64_2185 ();
 sg13g2_fill_2 FILLER_64_2237 ();
 sg13g2_fill_1 FILLER_64_2239 ();
 sg13g2_decap_4 FILLER_64_2256 ();
 sg13g2_decap_8 FILLER_64_2276 ();
 sg13g2_decap_8 FILLER_64_2304 ();
 sg13g2_fill_1 FILLER_64_2311 ();
 sg13g2_fill_2 FILLER_64_2321 ();
 sg13g2_decap_8 FILLER_64_2341 ();
 sg13g2_fill_2 FILLER_64_2348 ();
 sg13g2_fill_1 FILLER_64_2350 ();
 sg13g2_fill_2 FILLER_64_2382 ();
 sg13g2_fill_2 FILLER_64_2409 ();
 sg13g2_fill_1 FILLER_64_2411 ();
 sg13g2_decap_8 FILLER_64_2437 ();
 sg13g2_fill_2 FILLER_64_2444 ();
 sg13g2_decap_8 FILLER_64_2467 ();
 sg13g2_fill_2 FILLER_64_2474 ();
 sg13g2_decap_8 FILLER_64_2492 ();
 sg13g2_decap_8 FILLER_64_2499 ();
 sg13g2_fill_2 FILLER_64_2506 ();
 sg13g2_decap_8 FILLER_64_2513 ();
 sg13g2_fill_2 FILLER_64_2537 ();
 sg13g2_fill_1 FILLER_64_2539 ();
 sg13g2_decap_8 FILLER_64_2558 ();
 sg13g2_fill_1 FILLER_64_2565 ();
 sg13g2_decap_4 FILLER_64_2637 ();
 sg13g2_fill_1 FILLER_64_2641 ();
 sg13g2_fill_2 FILLER_64_2661 ();
 sg13g2_fill_1 FILLER_64_2663 ();
 sg13g2_fill_1 FILLER_64_2673 ();
 sg13g2_fill_1 FILLER_64_2719 ();
 sg13g2_decap_8 FILLER_64_2732 ();
 sg13g2_decap_4 FILLER_64_2739 ();
 sg13g2_fill_1 FILLER_64_2743 ();
 sg13g2_fill_1 FILLER_64_2763 ();
 sg13g2_fill_1 FILLER_64_2840 ();
 sg13g2_fill_1 FILLER_64_2861 ();
 sg13g2_decap_8 FILLER_64_2893 ();
 sg13g2_decap_8 FILLER_64_2908 ();
 sg13g2_decap_8 FILLER_64_2920 ();
 sg13g2_fill_1 FILLER_64_2940 ();
 sg13g2_fill_1 FILLER_64_2946 ();
 sg13g2_fill_1 FILLER_64_2953 ();
 sg13g2_fill_2 FILLER_64_2962 ();
 sg13g2_decap_4 FILLER_64_2984 ();
 sg13g2_fill_1 FILLER_64_2988 ();
 sg13g2_decap_4 FILLER_64_3012 ();
 sg13g2_fill_1 FILLER_64_3016 ();
 sg13g2_fill_2 FILLER_64_3030 ();
 sg13g2_fill_1 FILLER_64_3032 ();
 sg13g2_fill_1 FILLER_64_3057 ();
 sg13g2_fill_2 FILLER_64_3083 ();
 sg13g2_fill_1 FILLER_64_3085 ();
 sg13g2_fill_2 FILLER_64_3096 ();
 sg13g2_fill_2 FILLER_64_3112 ();
 sg13g2_fill_2 FILLER_64_3122 ();
 sg13g2_fill_1 FILLER_64_3124 ();
 sg13g2_fill_2 FILLER_64_3158 ();
 sg13g2_fill_2 FILLER_64_3186 ();
 sg13g2_decap_8 FILLER_64_3204 ();
 sg13g2_decap_4 FILLER_64_3211 ();
 sg13g2_decap_8 FILLER_64_3236 ();
 sg13g2_decap_8 FILLER_64_3263 ();
 sg13g2_fill_2 FILLER_64_3270 ();
 sg13g2_fill_1 FILLER_64_3272 ();
 sg13g2_decap_8 FILLER_64_3284 ();
 sg13g2_decap_4 FILLER_64_3291 ();
 sg13g2_fill_2 FILLER_64_3295 ();
 sg13g2_decap_4 FILLER_64_3310 ();
 sg13g2_decap_4 FILLER_64_3319 ();
 sg13g2_fill_1 FILLER_64_3323 ();
 sg13g2_decap_8 FILLER_64_3331 ();
 sg13g2_decap_4 FILLER_64_3338 ();
 sg13g2_fill_1 FILLER_64_3342 ();
 sg13g2_decap_4 FILLER_64_3350 ();
 sg13g2_fill_2 FILLER_64_3361 ();
 sg13g2_fill_2 FILLER_64_3372 ();
 sg13g2_decap_8 FILLER_64_3391 ();
 sg13g2_decap_4 FILLER_64_3398 ();
 sg13g2_fill_2 FILLER_64_3420 ();
 sg13g2_decap_4 FILLER_64_3447 ();
 sg13g2_fill_1 FILLER_64_3451 ();
 sg13g2_fill_1 FILLER_64_3510 ();
 sg13g2_fill_2 FILLER_64_3532 ();
 sg13g2_fill_2 FILLER_64_3543 ();
 sg13g2_fill_2 FILLER_64_3561 ();
 sg13g2_fill_1 FILLER_64_3563 ();
 sg13g2_fill_2 FILLER_64_3577 ();
 sg13g2_fill_1 FILLER_64_3579 ();
 sg13g2_decap_4 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_4 ();
 sg13g2_decap_8 FILLER_65_65 ();
 sg13g2_fill_2 FILLER_65_72 ();
 sg13g2_fill_1 FILLER_65_74 ();
 sg13g2_fill_2 FILLER_65_87 ();
 sg13g2_fill_2 FILLER_65_144 ();
 sg13g2_fill_2 FILLER_65_228 ();
 sg13g2_fill_1 FILLER_65_230 ();
 sg13g2_fill_2 FILLER_65_308 ();
 sg13g2_fill_1 FILLER_65_315 ();
 sg13g2_fill_1 FILLER_65_344 ();
 sg13g2_decap_8 FILLER_65_380 ();
 sg13g2_decap_4 FILLER_65_387 ();
 sg13g2_fill_2 FILLER_65_391 ();
 sg13g2_fill_2 FILLER_65_405 ();
 sg13g2_fill_1 FILLER_65_407 ();
 sg13g2_decap_8 FILLER_65_445 ();
 sg13g2_decap_4 FILLER_65_452 ();
 sg13g2_fill_2 FILLER_65_493 ();
 sg13g2_fill_1 FILLER_65_495 ();
 sg13g2_decap_4 FILLER_65_520 ();
 sg13g2_fill_1 FILLER_65_524 ();
 sg13g2_fill_2 FILLER_65_529 ();
 sg13g2_fill_1 FILLER_65_531 ();
 sg13g2_decap_4 FILLER_65_549 ();
 sg13g2_fill_2 FILLER_65_575 ();
 sg13g2_fill_1 FILLER_65_605 ();
 sg13g2_decap_8 FILLER_65_620 ();
 sg13g2_fill_2 FILLER_65_632 ();
 sg13g2_fill_2 FILLER_65_661 ();
 sg13g2_decap_8 FILLER_65_704 ();
 sg13g2_decap_8 FILLER_65_711 ();
 sg13g2_fill_1 FILLER_65_718 ();
 sg13g2_decap_4 FILLER_65_723 ();
 sg13g2_decap_8 FILLER_65_736 ();
 sg13g2_fill_1 FILLER_65_743 ();
 sg13g2_decap_8 FILLER_65_748 ();
 sg13g2_fill_2 FILLER_65_755 ();
 sg13g2_fill_2 FILLER_65_823 ();
 sg13g2_decap_8 FILLER_65_853 ();
 sg13g2_decap_4 FILLER_65_860 ();
 sg13g2_fill_1 FILLER_65_864 ();
 sg13g2_fill_2 FILLER_65_933 ();
 sg13g2_decap_4 FILLER_65_963 ();
 sg13g2_fill_1 FILLER_65_967 ();
 sg13g2_decap_4 FILLER_65_1000 ();
 sg13g2_fill_2 FILLER_65_1009 ();
 sg13g2_decap_4 FILLER_65_1016 ();
 sg13g2_fill_2 FILLER_65_1020 ();
 sg13g2_decap_4 FILLER_65_1050 ();
 sg13g2_fill_2 FILLER_65_1054 ();
 sg13g2_decap_4 FILLER_65_1084 ();
 sg13g2_decap_8 FILLER_65_1144 ();
 sg13g2_fill_2 FILLER_65_1160 ();
 sg13g2_fill_1 FILLER_65_1166 ();
 sg13g2_fill_2 FILLER_65_1171 ();
 sg13g2_fill_2 FILLER_65_1186 ();
 sg13g2_decap_4 FILLER_65_1214 ();
 sg13g2_fill_2 FILLER_65_1218 ();
 sg13g2_fill_2 FILLER_65_1228 ();
 sg13g2_fill_2 FILLER_65_1294 ();
 sg13g2_fill_2 FILLER_65_1304 ();
 sg13g2_fill_2 FILLER_65_1311 ();
 sg13g2_fill_2 FILLER_65_1317 ();
 sg13g2_decap_8 FILLER_65_1337 ();
 sg13g2_fill_1 FILLER_65_1356 ();
 sg13g2_fill_2 FILLER_65_1363 ();
 sg13g2_fill_1 FILLER_65_1365 ();
 sg13g2_fill_2 FILLER_65_1374 ();
 sg13g2_fill_1 FILLER_65_1386 ();
 sg13g2_fill_2 FILLER_65_1400 ();
 sg13g2_decap_8 FILLER_65_1407 ();
 sg13g2_decap_4 FILLER_65_1414 ();
 sg13g2_decap_4 FILLER_65_1434 ();
 sg13g2_decap_4 FILLER_65_1455 ();
 sg13g2_fill_1 FILLER_65_1459 ();
 sg13g2_fill_2 FILLER_65_1493 ();
 sg13g2_decap_4 FILLER_65_1503 ();
 sg13g2_fill_1 FILLER_65_1516 ();
 sg13g2_decap_4 FILLER_65_1521 ();
 sg13g2_fill_2 FILLER_65_1525 ();
 sg13g2_fill_2 FILLER_65_1547 ();
 sg13g2_fill_1 FILLER_65_1549 ();
 sg13g2_fill_2 FILLER_65_1564 ();
 sg13g2_fill_2 FILLER_65_1576 ();
 sg13g2_fill_1 FILLER_65_1583 ();
 sg13g2_fill_2 FILLER_65_1597 ();
 sg13g2_fill_2 FILLER_65_1647 ();
 sg13g2_fill_2 FILLER_65_1666 ();
 sg13g2_fill_1 FILLER_65_1668 ();
 sg13g2_fill_2 FILLER_65_1692 ();
 sg13g2_fill_1 FILLER_65_1694 ();
 sg13g2_fill_2 FILLER_65_1713 ();
 sg13g2_fill_1 FILLER_65_1742 ();
 sg13g2_decap_4 FILLER_65_1755 ();
 sg13g2_fill_1 FILLER_65_1759 ();
 sg13g2_decap_4 FILLER_65_1775 ();
 sg13g2_fill_1 FILLER_65_1779 ();
 sg13g2_fill_2 FILLER_65_1790 ();
 sg13g2_fill_1 FILLER_65_1792 ();
 sg13g2_decap_8 FILLER_65_1798 ();
 sg13g2_fill_2 FILLER_65_1805 ();
 sg13g2_fill_1 FILLER_65_1835 ();
 sg13g2_fill_2 FILLER_65_1853 ();
 sg13g2_fill_1 FILLER_65_1855 ();
 sg13g2_fill_2 FILLER_65_1869 ();
 sg13g2_fill_1 FILLER_65_1871 ();
 sg13g2_decap_8 FILLER_65_1891 ();
 sg13g2_decap_4 FILLER_65_1898 ();
 sg13g2_fill_1 FILLER_65_1902 ();
 sg13g2_fill_2 FILLER_65_1908 ();
 sg13g2_fill_1 FILLER_65_1934 ();
 sg13g2_fill_2 FILLER_65_1975 ();
 sg13g2_fill_1 FILLER_65_1990 ();
 sg13g2_decap_8 FILLER_65_2010 ();
 sg13g2_fill_2 FILLER_65_2017 ();
 sg13g2_fill_2 FILLER_65_2040 ();
 sg13g2_fill_1 FILLER_65_2042 ();
 sg13g2_decap_4 FILLER_65_2093 ();
 sg13g2_fill_2 FILLER_65_2097 ();
 sg13g2_decap_4 FILLER_65_2107 ();
 sg13g2_fill_2 FILLER_65_2128 ();
 sg13g2_fill_1 FILLER_65_2135 ();
 sg13g2_fill_2 FILLER_65_2154 ();
 sg13g2_fill_1 FILLER_65_2156 ();
 sg13g2_fill_1 FILLER_65_2170 ();
 sg13g2_fill_1 FILLER_65_2183 ();
 sg13g2_fill_1 FILLER_65_2198 ();
 sg13g2_decap_4 FILLER_65_2214 ();
 sg13g2_fill_2 FILLER_65_2233 ();
 sg13g2_decap_8 FILLER_65_2253 ();
 sg13g2_fill_1 FILLER_65_2260 ();
 sg13g2_decap_8 FILLER_65_2307 ();
 sg13g2_fill_2 FILLER_65_2325 ();
 sg13g2_decap_4 FILLER_65_2340 ();
 sg13g2_decap_4 FILLER_65_2374 ();
 sg13g2_fill_2 FILLER_65_2386 ();
 sg13g2_fill_1 FILLER_65_2388 ();
 sg13g2_decap_8 FILLER_65_2404 ();
 sg13g2_fill_1 FILLER_65_2411 ();
 sg13g2_decap_8 FILLER_65_2437 ();
 sg13g2_decap_4 FILLER_65_2444 ();
 sg13g2_fill_2 FILLER_65_2448 ();
 sg13g2_decap_8 FILLER_65_2463 ();
 sg13g2_decap_4 FILLER_65_2470 ();
 sg13g2_decap_8 FILLER_65_2499 ();
 sg13g2_fill_2 FILLER_65_2506 ();
 sg13g2_decap_4 FILLER_65_2526 ();
 sg13g2_fill_2 FILLER_65_2534 ();
 sg13g2_decap_8 FILLER_65_2550 ();
 sg13g2_fill_1 FILLER_65_2589 ();
 sg13g2_fill_2 FILLER_65_2627 ();
 sg13g2_fill_1 FILLER_65_2629 ();
 sg13g2_decap_4 FILLER_65_2638 ();
 sg13g2_decap_8 FILLER_65_2664 ();
 sg13g2_fill_2 FILLER_65_2671 ();
 sg13g2_decap_4 FILLER_65_2696 ();
 sg13g2_fill_1 FILLER_65_2705 ();
 sg13g2_decap_4 FILLER_65_2711 ();
 sg13g2_fill_1 FILLER_65_2724 ();
 sg13g2_decap_8 FILLER_65_2737 ();
 sg13g2_fill_1 FILLER_65_2744 ();
 sg13g2_fill_1 FILLER_65_2812 ();
 sg13g2_decap_8 FILLER_65_2818 ();
 sg13g2_fill_1 FILLER_65_2825 ();
 sg13g2_fill_2 FILLER_65_2843 ();
 sg13g2_fill_1 FILLER_65_2845 ();
 sg13g2_fill_2 FILLER_65_2866 ();
 sg13g2_fill_2 FILLER_65_2873 ();
 sg13g2_fill_1 FILLER_65_2875 ();
 sg13g2_fill_2 FILLER_65_2882 ();
 sg13g2_decap_8 FILLER_65_2917 ();
 sg13g2_fill_2 FILLER_65_2935 ();
 sg13g2_fill_1 FILLER_65_2937 ();
 sg13g2_fill_2 FILLER_65_2946 ();
 sg13g2_fill_1 FILLER_65_2948 ();
 sg13g2_decap_8 FILLER_65_3016 ();
 sg13g2_fill_2 FILLER_65_3023 ();
 sg13g2_fill_1 FILLER_65_3025 ();
 sg13g2_decap_8 FILLER_65_3053 ();
 sg13g2_fill_2 FILLER_65_3060 ();
 sg13g2_fill_1 FILLER_65_3080 ();
 sg13g2_decap_8 FILLER_65_3095 ();
 sg13g2_decap_4 FILLER_65_3102 ();
 sg13g2_fill_1 FILLER_65_3106 ();
 sg13g2_decap_8 FILLER_65_3122 ();
 sg13g2_fill_2 FILLER_65_3129 ();
 sg13g2_fill_1 FILLER_65_3156 ();
 sg13g2_decap_8 FILLER_65_3181 ();
 sg13g2_decap_4 FILLER_65_3188 ();
 sg13g2_fill_1 FILLER_65_3192 ();
 sg13g2_decap_8 FILLER_65_3214 ();
 sg13g2_decap_4 FILLER_65_3221 ();
 sg13g2_fill_1 FILLER_65_3225 ();
 sg13g2_fill_1 FILLER_65_3239 ();
 sg13g2_fill_1 FILLER_65_3265 ();
 sg13g2_decap_8 FILLER_65_3295 ();
 sg13g2_fill_1 FILLER_65_3302 ();
 sg13g2_decap_8 FILLER_65_3313 ();
 sg13g2_decap_4 FILLER_65_3320 ();
 sg13g2_decap_8 FILLER_65_3341 ();
 sg13g2_decap_8 FILLER_65_3348 ();
 sg13g2_decap_4 FILLER_65_3358 ();
 sg13g2_fill_2 FILLER_65_3362 ();
 sg13g2_decap_4 FILLER_65_3368 ();
 sg13g2_fill_1 FILLER_65_3372 ();
 sg13g2_decap_8 FILLER_65_3419 ();
 sg13g2_fill_2 FILLER_65_3426 ();
 sg13g2_decap_4 FILLER_65_3445 ();
 sg13g2_fill_1 FILLER_65_3449 ();
 sg13g2_decap_4 FILLER_65_3480 ();
 sg13g2_fill_1 FILLER_65_3484 ();
 sg13g2_decap_4 FILLER_65_3495 ();
 sg13g2_fill_1 FILLER_65_3499 ();
 sg13g2_decap_4 FILLER_65_3509 ();
 sg13g2_fill_2 FILLER_65_3513 ();
 sg13g2_decap_8 FILLER_65_3545 ();
 sg13g2_fill_1 FILLER_65_3552 ();
 sg13g2_fill_2 FILLER_65_3558 ();
 sg13g2_fill_1 FILLER_65_3560 ();
 sg13g2_decap_4 FILLER_65_3574 ();
 sg13g2_fill_2 FILLER_65_3578 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_7 ();
 sg13g2_fill_1 FILLER_66_9 ();
 sg13g2_decap_4 FILLER_66_14 ();
 sg13g2_fill_1 FILLER_66_18 ();
 sg13g2_fill_1 FILLER_66_105 ();
 sg13g2_fill_2 FILLER_66_173 ();
 sg13g2_fill_1 FILLER_66_175 ();
 sg13g2_fill_2 FILLER_66_203 ();
 sg13g2_fill_2 FILLER_66_228 ();
 sg13g2_fill_2 FILLER_66_277 ();
 sg13g2_fill_1 FILLER_66_279 ();
 sg13g2_fill_1 FILLER_66_291 ();
 sg13g2_fill_2 FILLER_66_321 ();
 sg13g2_fill_1 FILLER_66_327 ();
 sg13g2_fill_2 FILLER_66_345 ();
 sg13g2_fill_1 FILLER_66_347 ();
 sg13g2_decap_4 FILLER_66_361 ();
 sg13g2_fill_2 FILLER_66_375 ();
 sg13g2_decap_4 FILLER_66_385 ();
 sg13g2_fill_2 FILLER_66_389 ();
 sg13g2_decap_4 FILLER_66_416 ();
 sg13g2_decap_8 FILLER_66_440 ();
 sg13g2_decap_4 FILLER_66_447 ();
 sg13g2_fill_2 FILLER_66_479 ();
 sg13g2_decap_8 FILLER_66_492 ();
 sg13g2_fill_2 FILLER_66_499 ();
 sg13g2_fill_1 FILLER_66_501 ();
 sg13g2_decap_8 FILLER_66_520 ();
 sg13g2_fill_1 FILLER_66_527 ();
 sg13g2_decap_8 FILLER_66_550 ();
 sg13g2_fill_2 FILLER_66_557 ();
 sg13g2_fill_2 FILLER_66_582 ();
 sg13g2_fill_1 FILLER_66_595 ();
 sg13g2_decap_8 FILLER_66_615 ();
 sg13g2_fill_2 FILLER_66_622 ();
 sg13g2_fill_1 FILLER_66_624 ();
 sg13g2_fill_2 FILLER_66_666 ();
 sg13g2_fill_1 FILLER_66_668 ();
 sg13g2_decap_8 FILLER_66_683 ();
 sg13g2_fill_2 FILLER_66_690 ();
 sg13g2_fill_1 FILLER_66_692 ();
 sg13g2_decap_8 FILLER_66_707 ();
 sg13g2_fill_1 FILLER_66_714 ();
 sg13g2_fill_2 FILLER_66_752 ();
 sg13g2_fill_1 FILLER_66_758 ();
 sg13g2_decap_4 FILLER_66_809 ();
 sg13g2_fill_2 FILLER_66_823 ();
 sg13g2_fill_1 FILLER_66_825 ();
 sg13g2_fill_2 FILLER_66_831 ();
 sg13g2_fill_1 FILLER_66_833 ();
 sg13g2_decap_8 FILLER_66_884 ();
 sg13g2_decap_4 FILLER_66_891 ();
 sg13g2_decap_4 FILLER_66_909 ();
 sg13g2_fill_1 FILLER_66_940 ();
 sg13g2_decap_8 FILLER_66_961 ();
 sg13g2_decap_8 FILLER_66_1019 ();
 sg13g2_fill_1 FILLER_66_1026 ();
 sg13g2_fill_1 FILLER_66_1031 ();
 sg13g2_decap_8 FILLER_66_1035 ();
 sg13g2_decap_4 FILLER_66_1042 ();
 sg13g2_decap_4 FILLER_66_1067 ();
 sg13g2_fill_1 FILLER_66_1071 ();
 sg13g2_decap_8 FILLER_66_1107 ();
 sg13g2_decap_8 FILLER_66_1114 ();
 sg13g2_decap_8 FILLER_66_1121 ();
 sg13g2_fill_1 FILLER_66_1128 ();
 sg13g2_fill_1 FILLER_66_1195 ();
 sg13g2_fill_2 FILLER_66_1201 ();
 sg13g2_fill_1 FILLER_66_1203 ();
 sg13g2_decap_8 FILLER_66_1232 ();
 sg13g2_fill_2 FILLER_66_1239 ();
 sg13g2_fill_1 FILLER_66_1262 ();
 sg13g2_decap_8 FILLER_66_1269 ();
 sg13g2_fill_1 FILLER_66_1303 ();
 sg13g2_fill_2 FILLER_66_1333 ();
 sg13g2_fill_1 FILLER_66_1364 ();
 sg13g2_fill_2 FILLER_66_1386 ();
 sg13g2_fill_2 FILLER_66_1408 ();
 sg13g2_fill_1 FILLER_66_1410 ();
 sg13g2_fill_1 FILLER_66_1432 ();
 sg13g2_fill_2 FILLER_66_1448 ();
 sg13g2_fill_2 FILLER_66_1475 ();
 sg13g2_fill_1 FILLER_66_1486 ();
 sg13g2_decap_4 FILLER_66_1508 ();
 sg13g2_fill_1 FILLER_66_1512 ();
 sg13g2_fill_1 FILLER_66_1518 ();
 sg13g2_fill_2 FILLER_66_1544 ();
 sg13g2_fill_2 FILLER_66_1567 ();
 sg13g2_fill_1 FILLER_66_1569 ();
 sg13g2_decap_4 FILLER_66_1610 ();
 sg13g2_fill_2 FILLER_66_1651 ();
 sg13g2_decap_8 FILLER_66_1658 ();
 sg13g2_decap_4 FILLER_66_1665 ();
 sg13g2_decap_4 FILLER_66_1673 ();
 sg13g2_fill_1 FILLER_66_1677 ();
 sg13g2_fill_2 FILLER_66_1688 ();
 sg13g2_fill_1 FILLER_66_1699 ();
 sg13g2_fill_2 FILLER_66_1705 ();
 sg13g2_fill_1 FILLER_66_1707 ();
 sg13g2_decap_8 FILLER_66_1713 ();
 sg13g2_fill_2 FILLER_66_1720 ();
 sg13g2_decap_4 FILLER_66_1739 ();
 sg13g2_fill_1 FILLER_66_1754 ();
 sg13g2_decap_8 FILLER_66_1798 ();
 sg13g2_fill_1 FILLER_66_1822 ();
 sg13g2_fill_2 FILLER_66_1831 ();
 sg13g2_fill_1 FILLER_66_1833 ();
 sg13g2_decap_8 FILLER_66_1855 ();
 sg13g2_fill_2 FILLER_66_1897 ();
 sg13g2_fill_1 FILLER_66_1899 ();
 sg13g2_fill_1 FILLER_66_1905 ();
 sg13g2_decap_4 FILLER_66_1917 ();
 sg13g2_fill_2 FILLER_66_1927 ();
 sg13g2_decap_4 FILLER_66_1944 ();
 sg13g2_fill_2 FILLER_66_1989 ();
 sg13g2_fill_1 FILLER_66_1991 ();
 sg13g2_fill_1 FILLER_66_2020 ();
 sg13g2_fill_1 FILLER_66_2043 ();
 sg13g2_decap_4 FILLER_66_2066 ();
 sg13g2_fill_2 FILLER_66_2070 ();
 sg13g2_decap_4 FILLER_66_2096 ();
 sg13g2_decap_8 FILLER_66_2115 ();
 sg13g2_fill_2 FILLER_66_2147 ();
 sg13g2_decap_8 FILLER_66_2195 ();
 sg13g2_fill_1 FILLER_66_2202 ();
 sg13g2_decap_4 FILLER_66_2208 ();
 sg13g2_fill_1 FILLER_66_2212 ();
 sg13g2_fill_1 FILLER_66_2241 ();
 sg13g2_decap_8 FILLER_66_2255 ();
 sg13g2_fill_1 FILLER_66_2262 ();
 sg13g2_fill_2 FILLER_66_2298 ();
 sg13g2_fill_2 FILLER_66_2344 ();
 sg13g2_fill_1 FILLER_66_2346 ();
 sg13g2_decap_8 FILLER_66_2400 ();
 sg13g2_fill_1 FILLER_66_2407 ();
 sg13g2_fill_1 FILLER_66_2413 ();
 sg13g2_decap_8 FILLER_66_2433 ();
 sg13g2_fill_1 FILLER_66_2440 ();
 sg13g2_fill_1 FILLER_66_2472 ();
 sg13g2_fill_2 FILLER_66_2485 ();
 sg13g2_fill_2 FILLER_66_2493 ();
 sg13g2_decap_8 FILLER_66_2521 ();
 sg13g2_fill_1 FILLER_66_2528 ();
 sg13g2_fill_2 FILLER_66_2534 ();
 sg13g2_fill_1 FILLER_66_2536 ();
 sg13g2_fill_1 FILLER_66_2562 ();
 sg13g2_fill_1 FILLER_66_2604 ();
 sg13g2_fill_1 FILLER_66_2646 ();
 sg13g2_decap_8 FILLER_66_2663 ();
 sg13g2_decap_8 FILLER_66_2670 ();
 sg13g2_decap_4 FILLER_66_2690 ();
 sg13g2_fill_2 FILLER_66_2718 ();
 sg13g2_fill_1 FILLER_66_2720 ();
 sg13g2_fill_1 FILLER_66_2740 ();
 sg13g2_decap_8 FILLER_66_2745 ();
 sg13g2_fill_2 FILLER_66_2752 ();
 sg13g2_fill_1 FILLER_66_2754 ();
 sg13g2_decap_4 FILLER_66_2790 ();
 sg13g2_decap_8 FILLER_66_2809 ();
 sg13g2_decap_4 FILLER_66_2816 ();
 sg13g2_fill_2 FILLER_66_2820 ();
 sg13g2_fill_1 FILLER_66_2840 ();
 sg13g2_fill_2 FILLER_66_2870 ();
 sg13g2_fill_1 FILLER_66_2872 ();
 sg13g2_decap_8 FILLER_66_2904 ();
 sg13g2_decap_8 FILLER_66_2911 ();
 sg13g2_fill_2 FILLER_66_2927 ();
 sg13g2_fill_1 FILLER_66_2929 ();
 sg13g2_decap_8 FILLER_66_2956 ();
 sg13g2_decap_4 FILLER_66_2966 ();
 sg13g2_fill_2 FILLER_66_2975 ();
 sg13g2_fill_1 FILLER_66_2982 ();
 sg13g2_decap_8 FILLER_66_3007 ();
 sg13g2_fill_2 FILLER_66_3014 ();
 sg13g2_fill_1 FILLER_66_3016 ();
 sg13g2_fill_2 FILLER_66_3041 ();
 sg13g2_fill_1 FILLER_66_3059 ();
 sg13g2_fill_1 FILLER_66_3072 ();
 sg13g2_decap_4 FILLER_66_3095 ();
 sg13g2_fill_1 FILLER_66_3099 ();
 sg13g2_decap_8 FILLER_66_3128 ();
 sg13g2_fill_2 FILLER_66_3135 ();
 sg13g2_fill_1 FILLER_66_3137 ();
 sg13g2_decap_4 FILLER_66_3151 ();
 sg13g2_fill_1 FILLER_66_3155 ();
 sg13g2_fill_2 FILLER_66_3169 ();
 sg13g2_fill_1 FILLER_66_3171 ();
 sg13g2_decap_8 FILLER_66_3185 ();
 sg13g2_decap_4 FILLER_66_3195 ();
 sg13g2_fill_2 FILLER_66_3244 ();
 sg13g2_fill_1 FILLER_66_3246 ();
 sg13g2_decap_4 FILLER_66_3271 ();
 sg13g2_fill_2 FILLER_66_3275 ();
 sg13g2_decap_8 FILLER_66_3285 ();
 sg13g2_fill_2 FILLER_66_3292 ();
 sg13g2_fill_1 FILLER_66_3294 ();
 sg13g2_fill_2 FILLER_66_3323 ();
 sg13g2_fill_1 FILLER_66_3325 ();
 sg13g2_fill_1 FILLER_66_3354 ();
 sg13g2_decap_8 FILLER_66_3387 ();
 sg13g2_decap_4 FILLER_66_3394 ();
 sg13g2_fill_1 FILLER_66_3398 ();
 sg13g2_decap_4 FILLER_66_3422 ();
 sg13g2_decap_8 FILLER_66_3434 ();
 sg13g2_decap_8 FILLER_66_3441 ();
 sg13g2_decap_4 FILLER_66_3448 ();
 sg13g2_fill_1 FILLER_66_3452 ();
 sg13g2_decap_8 FILLER_66_3457 ();
 sg13g2_decap_4 FILLER_66_3464 ();
 sg13g2_fill_1 FILLER_66_3468 ();
 sg13g2_decap_8 FILLER_66_3472 ();
 sg13g2_fill_2 FILLER_66_3479 ();
 sg13g2_fill_1 FILLER_66_3481 ();
 sg13g2_decap_8 FILLER_66_3500 ();
 sg13g2_decap_8 FILLER_66_3507 ();
 sg13g2_decap_8 FILLER_66_3514 ();
 sg13g2_decap_4 FILLER_66_3521 ();
 sg13g2_fill_1 FILLER_66_3529 ();
 sg13g2_fill_1 FILLER_66_3543 ();
 sg13g2_fill_2 FILLER_66_3550 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_4 FILLER_67_7 ();
 sg13g2_fill_2 FILLER_67_11 ();
 sg13g2_fill_2 FILLER_67_41 ();
 sg13g2_fill_1 FILLER_67_43 ();
 sg13g2_fill_2 FILLER_67_84 ();
 sg13g2_fill_1 FILLER_67_86 ();
 sg13g2_fill_2 FILLER_67_155 ();
 sg13g2_fill_1 FILLER_67_157 ();
 sg13g2_fill_2 FILLER_67_176 ();
 sg13g2_fill_1 FILLER_67_178 ();
 sg13g2_fill_2 FILLER_67_193 ();
 sg13g2_fill_2 FILLER_67_228 ();
 sg13g2_fill_2 FILLER_67_274 ();
 sg13g2_fill_1 FILLER_67_276 ();
 sg13g2_decap_8 FILLER_67_293 ();
 sg13g2_decap_4 FILLER_67_300 ();
 sg13g2_fill_1 FILLER_67_304 ();
 sg13g2_fill_2 FILLER_67_313 ();
 sg13g2_fill_1 FILLER_67_315 ();
 sg13g2_fill_1 FILLER_67_320 ();
 sg13g2_fill_2 FILLER_67_326 ();
 sg13g2_fill_2 FILLER_67_348 ();
 sg13g2_fill_1 FILLER_67_350 ();
 sg13g2_fill_1 FILLER_67_364 ();
 sg13g2_fill_1 FILLER_67_395 ();
 sg13g2_decap_4 FILLER_67_417 ();
 sg13g2_decap_8 FILLER_67_445 ();
 sg13g2_fill_1 FILLER_67_452 ();
 sg13g2_decap_8 FILLER_67_464 ();
 sg13g2_decap_8 FILLER_67_471 ();
 sg13g2_decap_8 FILLER_67_484 ();
 sg13g2_fill_2 FILLER_67_504 ();
 sg13g2_decap_8 FILLER_67_526 ();
 sg13g2_fill_2 FILLER_67_542 ();
 sg13g2_decap_4 FILLER_67_548 ();
 sg13g2_fill_2 FILLER_67_552 ();
 sg13g2_decap_4 FILLER_67_577 ();
 sg13g2_fill_2 FILLER_67_581 ();
 sg13g2_fill_1 FILLER_67_604 ();
 sg13g2_decap_8 FILLER_67_609 ();
 sg13g2_decap_8 FILLER_67_616 ();
 sg13g2_decap_4 FILLER_67_623 ();
 sg13g2_fill_2 FILLER_67_657 ();
 sg13g2_fill_1 FILLER_67_659 ();
 sg13g2_fill_2 FILLER_67_720 ();
 sg13g2_fill_2 FILLER_67_731 ();
 sg13g2_fill_1 FILLER_67_746 ();
 sg13g2_fill_1 FILLER_67_762 ();
 sg13g2_fill_2 FILLER_67_791 ();
 sg13g2_decap_4 FILLER_67_872 ();
 sg13g2_fill_1 FILLER_67_876 ();
 sg13g2_decap_4 FILLER_67_881 ();
 sg13g2_fill_2 FILLER_67_885 ();
 sg13g2_fill_2 FILLER_67_896 ();
 sg13g2_fill_1 FILLER_67_898 ();
 sg13g2_fill_2 FILLER_67_931 ();
 sg13g2_decap_4 FILLER_67_1000 ();
 sg13g2_decap_8 FILLER_67_1018 ();
 sg13g2_fill_2 FILLER_67_1025 ();
 sg13g2_fill_1 FILLER_67_1027 ();
 sg13g2_fill_2 FILLER_67_1033 ();
 sg13g2_fill_2 FILLER_67_1040 ();
 sg13g2_fill_1 FILLER_67_1042 ();
 sg13g2_fill_1 FILLER_67_1096 ();
 sg13g2_fill_2 FILLER_67_1116 ();
 sg13g2_fill_1 FILLER_67_1133 ();
 sg13g2_decap_8 FILLER_67_1138 ();
 sg13g2_decap_4 FILLER_67_1145 ();
 sg13g2_fill_1 FILLER_67_1149 ();
 sg13g2_decap_4 FILLER_67_1164 ();
 sg13g2_fill_1 FILLER_67_1168 ();
 sg13g2_fill_1 FILLER_67_1205 ();
 sg13g2_fill_1 FILLER_67_1216 ();
 sg13g2_fill_1 FILLER_67_1221 ();
 sg13g2_decap_8 FILLER_67_1231 ();
 sg13g2_fill_1 FILLER_67_1238 ();
 sg13g2_decap_4 FILLER_67_1252 ();
 sg13g2_fill_1 FILLER_67_1256 ();
 sg13g2_fill_2 FILLER_67_1261 ();
 sg13g2_fill_1 FILLER_67_1263 ();
 sg13g2_fill_2 FILLER_67_1277 ();
 sg13g2_fill_2 FILLER_67_1300 ();
 sg13g2_fill_1 FILLER_67_1302 ();
 sg13g2_fill_2 FILLER_67_1307 ();
 sg13g2_decap_8 FILLER_67_1334 ();
 sg13g2_fill_2 FILLER_67_1341 ();
 sg13g2_fill_1 FILLER_67_1356 ();
 sg13g2_fill_1 FILLER_67_1402 ();
 sg13g2_decap_8 FILLER_67_1412 ();
 sg13g2_fill_2 FILLER_67_1441 ();
 sg13g2_decap_8 FILLER_67_1479 ();
 sg13g2_fill_2 FILLER_67_1486 ();
 sg13g2_fill_1 FILLER_67_1488 ();
 sg13g2_fill_2 FILLER_67_1545 ();
 sg13g2_fill_2 FILLER_67_1552 ();
 sg13g2_fill_1 FILLER_67_1572 ();
 sg13g2_fill_2 FILLER_67_1578 ();
 sg13g2_fill_2 FILLER_67_1620 ();
 sg13g2_fill_2 FILLER_67_1644 ();
 sg13g2_fill_2 FILLER_67_1672 ();
 sg13g2_fill_1 FILLER_67_1674 ();
 sg13g2_decap_4 FILLER_67_1699 ();
 sg13g2_fill_2 FILLER_67_1703 ();
 sg13g2_decap_8 FILLER_67_1720 ();
 sg13g2_decap_8 FILLER_67_1727 ();
 sg13g2_fill_2 FILLER_67_1734 ();
 sg13g2_decap_4 FILLER_67_1756 ();
 sg13g2_fill_2 FILLER_67_1760 ();
 sg13g2_decap_8 FILLER_67_1802 ();
 sg13g2_decap_8 FILLER_67_1809 ();
 sg13g2_decap_4 FILLER_67_1816 ();
 sg13g2_fill_1 FILLER_67_1820 ();
 sg13g2_decap_4 FILLER_67_1848 ();
 sg13g2_decap_8 FILLER_67_1857 ();
 sg13g2_fill_1 FILLER_67_1864 ();
 sg13g2_decap_8 FILLER_67_1881 ();
 sg13g2_fill_1 FILLER_67_1888 ();
 sg13g2_fill_2 FILLER_67_1894 ();
 sg13g2_fill_1 FILLER_67_1896 ();
 sg13g2_fill_1 FILLER_67_1946 ();
 sg13g2_decap_8 FILLER_67_1966 ();
 sg13g2_fill_1 FILLER_67_1973 ();
 sg13g2_fill_2 FILLER_67_1991 ();
 sg13g2_decap_8 FILLER_67_2013 ();
 sg13g2_fill_1 FILLER_67_2020 ();
 sg13g2_fill_2 FILLER_67_2029 ();
 sg13g2_fill_2 FILLER_67_2040 ();
 sg13g2_decap_8 FILLER_67_2054 ();
 sg13g2_decap_4 FILLER_67_2061 ();
 sg13g2_decap_8 FILLER_67_2070 ();
 sg13g2_decap_4 FILLER_67_2077 ();
 sg13g2_fill_1 FILLER_67_2081 ();
 sg13g2_decap_8 FILLER_67_2087 ();
 sg13g2_decap_8 FILLER_67_2094 ();
 sg13g2_fill_1 FILLER_67_2114 ();
 sg13g2_decap_8 FILLER_67_2123 ();
 sg13g2_fill_2 FILLER_67_2130 ();
 sg13g2_fill_1 FILLER_67_2132 ();
 sg13g2_fill_1 FILLER_67_2171 ();
 sg13g2_decap_8 FILLER_67_2184 ();
 sg13g2_fill_2 FILLER_67_2191 ();
 sg13g2_fill_1 FILLER_67_2200 ();
 sg13g2_decap_8 FILLER_67_2209 ();
 sg13g2_decap_4 FILLER_67_2216 ();
 sg13g2_fill_1 FILLER_67_2234 ();
 sg13g2_fill_2 FILLER_67_2240 ();
 sg13g2_fill_2 FILLER_67_2255 ();
 sg13g2_fill_1 FILLER_67_2257 ();
 sg13g2_decap_4 FILLER_67_2284 ();
 sg13g2_fill_1 FILLER_67_2288 ();
 sg13g2_fill_1 FILLER_67_2297 ();
 sg13g2_fill_1 FILLER_67_2311 ();
 sg13g2_decap_4 FILLER_67_2347 ();
 sg13g2_fill_2 FILLER_67_2351 ();
 sg13g2_fill_2 FILLER_67_2366 ();
 sg13g2_fill_1 FILLER_67_2381 ();
 sg13g2_fill_1 FILLER_67_2402 ();
 sg13g2_fill_2 FILLER_67_2421 ();
 sg13g2_decap_8 FILLER_67_2440 ();
 sg13g2_decap_4 FILLER_67_2447 ();
 sg13g2_decap_8 FILLER_67_2459 ();
 sg13g2_fill_1 FILLER_67_2466 ();
 sg13g2_fill_2 FILLER_67_2476 ();
 sg13g2_fill_2 FILLER_67_2497 ();
 sg13g2_decap_8 FILLER_67_2504 ();
 sg13g2_fill_2 FILLER_67_2511 ();
 sg13g2_decap_4 FILLER_67_2529 ();
 sg13g2_fill_1 FILLER_67_2533 ();
 sg13g2_decap_8 FILLER_67_2554 ();
 sg13g2_fill_2 FILLER_67_2587 ();
 sg13g2_fill_2 FILLER_67_2593 ();
 sg13g2_decap_8 FILLER_67_2610 ();
 sg13g2_decap_4 FILLER_67_2617 ();
 sg13g2_fill_2 FILLER_67_2621 ();
 sg13g2_fill_1 FILLER_67_2640 ();
 sg13g2_decap_8 FILLER_67_2663 ();
 sg13g2_fill_2 FILLER_67_2670 ();
 sg13g2_fill_2 FILLER_67_2695 ();
 sg13g2_fill_1 FILLER_67_2697 ();
 sg13g2_decap_8 FILLER_67_2710 ();
 sg13g2_fill_2 FILLER_67_2721 ();
 sg13g2_fill_2 FILLER_67_2733 ();
 sg13g2_fill_1 FILLER_67_2735 ();
 sg13g2_fill_1 FILLER_67_2776 ();
 sg13g2_decap_8 FILLER_67_2785 ();
 sg13g2_fill_2 FILLER_67_2792 ();
 sg13g2_fill_1 FILLER_67_2794 ();
 sg13g2_fill_2 FILLER_67_2817 ();
 sg13g2_fill_1 FILLER_67_2819 ();
 sg13g2_fill_1 FILLER_67_2856 ();
 sg13g2_fill_2 FILLER_67_2870 ();
 sg13g2_fill_1 FILLER_67_2872 ();
 sg13g2_decap_8 FILLER_67_2899 ();
 sg13g2_fill_2 FILLER_67_2906 ();
 sg13g2_fill_1 FILLER_67_2908 ();
 sg13g2_fill_2 FILLER_67_2931 ();
 sg13g2_fill_1 FILLER_67_2933 ();
 sg13g2_fill_1 FILLER_67_2947 ();
 sg13g2_decap_4 FILLER_67_2951 ();
 sg13g2_decap_8 FILLER_67_2967 ();
 sg13g2_decap_8 FILLER_67_2989 ();
 sg13g2_decap_4 FILLER_67_2996 ();
 sg13g2_fill_1 FILLER_67_3009 ();
 sg13g2_decap_4 FILLER_67_3029 ();
 sg13g2_decap_4 FILLER_67_3057 ();
 sg13g2_fill_2 FILLER_67_3061 ();
 sg13g2_decap_8 FILLER_67_3076 ();
 sg13g2_decap_8 FILLER_67_3083 ();
 sg13g2_fill_2 FILLER_67_3100 ();
 sg13g2_decap_8 FILLER_67_3118 ();
 sg13g2_decap_4 FILLER_67_3125 ();
 sg13g2_fill_2 FILLER_67_3129 ();
 sg13g2_fill_2 FILLER_67_3135 ();
 sg13g2_fill_1 FILLER_67_3137 ();
 sg13g2_fill_1 FILLER_67_3151 ();
 sg13g2_decap_4 FILLER_67_3202 ();
 sg13g2_fill_2 FILLER_67_3206 ();
 sg13g2_fill_1 FILLER_67_3221 ();
 sg13g2_fill_1 FILLER_67_3267 ();
 sg13g2_decap_8 FILLER_67_3296 ();
 sg13g2_fill_1 FILLER_67_3303 ();
 sg13g2_fill_1 FILLER_67_3308 ();
 sg13g2_fill_2 FILLER_67_3326 ();
 sg13g2_fill_1 FILLER_67_3328 ();
 sg13g2_fill_2 FILLER_67_3333 ();
 sg13g2_fill_1 FILLER_67_3335 ();
 sg13g2_fill_1 FILLER_67_3354 ();
 sg13g2_fill_1 FILLER_67_3369 ();
 sg13g2_decap_4 FILLER_67_3392 ();
 sg13g2_fill_2 FILLER_67_3396 ();
 sg13g2_fill_1 FILLER_67_3402 ();
 sg13g2_fill_2 FILLER_67_3542 ();
 sg13g2_fill_1 FILLER_67_3549 ();
 sg13g2_fill_2 FILLER_67_3563 ();
 sg13g2_decap_8 FILLER_67_3569 ();
 sg13g2_decap_4 FILLER_67_3576 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_4 FILLER_68_21 ();
 sg13g2_fill_2 FILLER_68_34 ();
 sg13g2_fill_2 FILLER_68_100 ();
 sg13g2_fill_2 FILLER_68_133 ();
 sg13g2_fill_1 FILLER_68_135 ();
 sg13g2_fill_1 FILLER_68_149 ();
 sg13g2_fill_2 FILLER_68_243 ();
 sg13g2_fill_2 FILLER_68_266 ();
 sg13g2_fill_2 FILLER_68_295 ();
 sg13g2_fill_1 FILLER_68_297 ();
 sg13g2_fill_1 FILLER_68_314 ();
 sg13g2_fill_1 FILLER_68_323 ();
 sg13g2_fill_2 FILLER_68_332 ();
 sg13g2_fill_1 FILLER_68_339 ();
 sg13g2_decap_4 FILLER_68_350 ();
 sg13g2_fill_1 FILLER_68_354 ();
 sg13g2_decap_8 FILLER_68_383 ();
 sg13g2_fill_1 FILLER_68_390 ();
 sg13g2_decap_4 FILLER_68_417 ();
 sg13g2_fill_2 FILLER_68_421 ();
 sg13g2_fill_2 FILLER_68_479 ();
 sg13g2_fill_1 FILLER_68_494 ();
 sg13g2_fill_1 FILLER_68_520 ();
 sg13g2_fill_1 FILLER_68_526 ();
 sg13g2_fill_1 FILLER_68_544 ();
 sg13g2_decap_8 FILLER_68_551 ();
 sg13g2_fill_2 FILLER_68_575 ();
 sg13g2_decap_8 FILLER_68_585 ();
 sg13g2_decap_4 FILLER_68_592 ();
 sg13g2_fill_2 FILLER_68_605 ();
 sg13g2_fill_2 FILLER_68_628 ();
 sg13g2_fill_2 FILLER_68_643 ();
 sg13g2_decap_8 FILLER_68_672 ();
 sg13g2_fill_2 FILLER_68_679 ();
 sg13g2_fill_1 FILLER_68_681 ();
 sg13g2_decap_8 FILLER_68_708 ();
 sg13g2_fill_1 FILLER_68_715 ();
 sg13g2_fill_2 FILLER_68_727 ();
 sg13g2_fill_1 FILLER_68_729 ();
 sg13g2_decap_4 FILLER_68_739 ();
 sg13g2_fill_2 FILLER_68_743 ();
 sg13g2_decap_4 FILLER_68_764 ();
 sg13g2_fill_2 FILLER_68_772 ();
 sg13g2_decap_8 FILLER_68_778 ();
 sg13g2_decap_8 FILLER_68_785 ();
 sg13g2_decap_4 FILLER_68_792 ();
 sg13g2_fill_1 FILLER_68_796 ();
 sg13g2_fill_2 FILLER_68_801 ();
 sg13g2_decap_4 FILLER_68_807 ();
 sg13g2_fill_1 FILLER_68_811 ();
 sg13g2_decap_4 FILLER_68_825 ();
 sg13g2_fill_2 FILLER_68_829 ();
 sg13g2_fill_2 FILLER_68_849 ();
 sg13g2_fill_1 FILLER_68_864 ();
 sg13g2_decap_8 FILLER_68_898 ();
 sg13g2_fill_2 FILLER_68_905 ();
 sg13g2_fill_1 FILLER_68_907 ();
 sg13g2_fill_1 FILLER_68_949 ();
 sg13g2_decap_8 FILLER_68_960 ();
 sg13g2_decap_8 FILLER_68_967 ();
 sg13g2_fill_1 FILLER_68_974 ();
 sg13g2_fill_2 FILLER_68_992 ();
 sg13g2_fill_1 FILLER_68_994 ();
 sg13g2_decap_4 FILLER_68_1011 ();
 sg13g2_fill_1 FILLER_68_1015 ();
 sg13g2_fill_2 FILLER_68_1044 ();
 sg13g2_fill_2 FILLER_68_1055 ();
 sg13g2_fill_1 FILLER_68_1057 ();
 sg13g2_decap_8 FILLER_68_1066 ();
 sg13g2_decap_4 FILLER_68_1073 ();
 sg13g2_fill_2 FILLER_68_1107 ();
 sg13g2_fill_1 FILLER_68_1109 ();
 sg13g2_decap_8 FILLER_68_1128 ();
 sg13g2_fill_2 FILLER_68_1135 ();
 sg13g2_fill_1 FILLER_68_1137 ();
 sg13g2_decap_4 FILLER_68_1141 ();
 sg13g2_fill_2 FILLER_68_1167 ();
 sg13g2_fill_1 FILLER_68_1169 ();
 sg13g2_fill_1 FILLER_68_1201 ();
 sg13g2_decap_8 FILLER_68_1239 ();
 sg13g2_fill_2 FILLER_68_1246 ();
 sg13g2_fill_1 FILLER_68_1248 ();
 sg13g2_decap_4 FILLER_68_1277 ();
 sg13g2_fill_1 FILLER_68_1281 ();
 sg13g2_fill_2 FILLER_68_1295 ();
 sg13g2_decap_4 FILLER_68_1307 ();
 sg13g2_fill_2 FILLER_68_1311 ();
 sg13g2_fill_2 FILLER_68_1334 ();
 sg13g2_fill_2 FILLER_68_1377 ();
 sg13g2_fill_1 FILLER_68_1379 ();
 sg13g2_decap_8 FILLER_68_1410 ();
 sg13g2_decap_4 FILLER_68_1446 ();
 sg13g2_fill_2 FILLER_68_1450 ();
 sg13g2_fill_2 FILLER_68_1464 ();
 sg13g2_decap_4 FILLER_68_1470 ();
 sg13g2_fill_1 FILLER_68_1474 ();
 sg13g2_fill_1 FILLER_68_1488 ();
 sg13g2_decap_4 FILLER_68_1514 ();
 sg13g2_fill_1 FILLER_68_1518 ();
 sg13g2_fill_1 FILLER_68_1532 ();
 sg13g2_fill_1 FILLER_68_1549 ();
 sg13g2_fill_1 FILLER_68_1576 ();
 sg13g2_decap_8 FILLER_68_1589 ();
 sg13g2_fill_2 FILLER_68_1596 ();
 sg13g2_fill_1 FILLER_68_1598 ();
 sg13g2_decap_8 FILLER_68_1620 ();
 sg13g2_fill_1 FILLER_68_1627 ();
 sg13g2_fill_2 FILLER_68_1672 ();
 sg13g2_fill_1 FILLER_68_1674 ();
 sg13g2_decap_4 FILLER_68_1701 ();
 sg13g2_fill_1 FILLER_68_1705 ();
 sg13g2_fill_1 FILLER_68_1750 ();
 sg13g2_fill_2 FILLER_68_1766 ();
 sg13g2_fill_2 FILLER_68_1773 ();
 sg13g2_fill_1 FILLER_68_1775 ();
 sg13g2_decap_4 FILLER_68_1797 ();
 sg13g2_fill_1 FILLER_68_1801 ();
 sg13g2_decap_8 FILLER_68_1817 ();
 sg13g2_fill_1 FILLER_68_1824 ();
 sg13g2_fill_2 FILLER_68_1838 ();
 sg13g2_fill_1 FILLER_68_1840 ();
 sg13g2_fill_2 FILLER_68_1862 ();
 sg13g2_decap_8 FILLER_68_1893 ();
 sg13g2_fill_2 FILLER_68_1900 ();
 sg13g2_fill_1 FILLER_68_1902 ();
 sg13g2_fill_2 FILLER_68_1941 ();
 sg13g2_fill_1 FILLER_68_1943 ();
 sg13g2_decap_4 FILLER_68_1965 ();
 sg13g2_decap_8 FILLER_68_2004 ();
 sg13g2_fill_2 FILLER_68_2024 ();
 sg13g2_fill_1 FILLER_68_2026 ();
 sg13g2_fill_2 FILLER_68_2053 ();
 sg13g2_fill_1 FILLER_68_2107 ();
 sg13g2_decap_4 FILLER_68_2127 ();
 sg13g2_fill_1 FILLER_68_2131 ();
 sg13g2_fill_1 FILLER_68_2169 ();
 sg13g2_decap_4 FILLER_68_2179 ();
 sg13g2_fill_2 FILLER_68_2217 ();
 sg13g2_fill_2 FILLER_68_2244 ();
 sg13g2_decap_8 FILLER_68_2254 ();
 sg13g2_decap_8 FILLER_68_2261 ();
 sg13g2_decap_4 FILLER_68_2268 ();
 sg13g2_fill_2 FILLER_68_2272 ();
 sg13g2_fill_1 FILLER_68_2287 ();
 sg13g2_fill_1 FILLER_68_2301 ();
 sg13g2_fill_1 FILLER_68_2353 ();
 sg13g2_decap_8 FILLER_68_2366 ();
 sg13g2_decap_8 FILLER_68_2373 ();
 sg13g2_decap_8 FILLER_68_2380 ();
 sg13g2_fill_2 FILLER_68_2387 ();
 sg13g2_decap_8 FILLER_68_2394 ();
 sg13g2_decap_8 FILLER_68_2401 ();
 sg13g2_fill_2 FILLER_68_2428 ();
 sg13g2_decap_8 FILLER_68_2435 ();
 sg13g2_fill_2 FILLER_68_2442 ();
 sg13g2_fill_1 FILLER_68_2444 ();
 sg13g2_fill_1 FILLER_68_2470 ();
 sg13g2_fill_2 FILLER_68_2527 ();
 sg13g2_decap_8 FILLER_68_2545 ();
 sg13g2_decap_4 FILLER_68_2552 ();
 sg13g2_fill_1 FILLER_68_2556 ();
 sg13g2_fill_2 FILLER_68_2585 ();
 sg13g2_fill_2 FILLER_68_2591 ();
 sg13g2_fill_1 FILLER_68_2593 ();
 sg13g2_decap_8 FILLER_68_2622 ();
 sg13g2_decap_8 FILLER_68_2629 ();
 sg13g2_decap_4 FILLER_68_2636 ();
 sg13g2_fill_1 FILLER_68_2640 ();
 sg13g2_fill_2 FILLER_68_2660 ();
 sg13g2_decap_4 FILLER_68_2675 ();
 sg13g2_fill_2 FILLER_68_2679 ();
 sg13g2_decap_8 FILLER_68_2692 ();
 sg13g2_decap_4 FILLER_68_2699 ();
 sg13g2_fill_2 FILLER_68_2703 ();
 sg13g2_fill_1 FILLER_68_2709 ();
 sg13g2_decap_4 FILLER_68_2718 ();
 sg13g2_fill_1 FILLER_68_2722 ();
 sg13g2_decap_4 FILLER_68_2727 ();
 sg13g2_fill_2 FILLER_68_2731 ();
 sg13g2_fill_1 FILLER_68_2738 ();
 sg13g2_decap_8 FILLER_68_2743 ();
 sg13g2_decap_8 FILLER_68_2750 ();
 sg13g2_fill_2 FILLER_68_2757 ();
 sg13g2_fill_1 FILLER_68_2771 ();
 sg13g2_fill_2 FILLER_68_2777 ();
 sg13g2_fill_2 FILLER_68_2792 ();
 sg13g2_fill_1 FILLER_68_2794 ();
 sg13g2_decap_8 FILLER_68_2823 ();
 sg13g2_decap_8 FILLER_68_2830 ();
 sg13g2_fill_2 FILLER_68_2837 ();
 sg13g2_fill_2 FILLER_68_2862 ();
 sg13g2_fill_1 FILLER_68_2886 ();
 sg13g2_fill_1 FILLER_68_2899 ();
 sg13g2_decap_4 FILLER_68_2941 ();
 sg13g2_fill_2 FILLER_68_2945 ();
 sg13g2_fill_2 FILLER_68_2955 ();
 sg13g2_fill_2 FILLER_68_2989 ();
 sg13g2_fill_1 FILLER_68_2991 ();
 sg13g2_fill_1 FILLER_68_3013 ();
 sg13g2_fill_2 FILLER_68_3042 ();
 sg13g2_decap_8 FILLER_68_3051 ();
 sg13g2_decap_4 FILLER_68_3058 ();
 sg13g2_fill_2 FILLER_68_3067 ();
 sg13g2_fill_1 FILLER_68_3069 ();
 sg13g2_decap_8 FILLER_68_3074 ();
 sg13g2_decap_4 FILLER_68_3081 ();
 sg13g2_decap_4 FILLER_68_3099 ();
 sg13g2_decap_8 FILLER_68_3108 ();
 sg13g2_decap_8 FILLER_68_3115 ();
 sg13g2_decap_8 FILLER_68_3122 ();
 sg13g2_decap_4 FILLER_68_3129 ();
 sg13g2_decap_8 FILLER_68_3139 ();
 sg13g2_decap_4 FILLER_68_3146 ();
 sg13g2_fill_2 FILLER_68_3154 ();
 sg13g2_decap_4 FILLER_68_3179 ();
 sg13g2_fill_1 FILLER_68_3183 ();
 sg13g2_fill_2 FILLER_68_3194 ();
 sg13g2_fill_1 FILLER_68_3196 ();
 sg13g2_fill_2 FILLER_68_3228 ();
 sg13g2_fill_2 FILLER_68_3239 ();
 sg13g2_fill_2 FILLER_68_3246 ();
 sg13g2_fill_2 FILLER_68_3266 ();
 sg13g2_fill_2 FILLER_68_3287 ();
 sg13g2_fill_2 FILLER_68_3331 ();
 sg13g2_fill_1 FILLER_68_3359 ();
 sg13g2_fill_2 FILLER_68_3411 ();
 sg13g2_fill_1 FILLER_68_3413 ();
 sg13g2_fill_2 FILLER_68_3428 ();
 sg13g2_fill_1 FILLER_68_3430 ();
 sg13g2_decap_8 FILLER_68_3456 ();
 sg13g2_fill_2 FILLER_68_3475 ();
 sg13g2_decap_4 FILLER_68_3495 ();
 sg13g2_fill_1 FILLER_68_3499 ();
 sg13g2_fill_2 FILLER_68_3508 ();
 sg13g2_fill_1 FILLER_68_3518 ();
 sg13g2_decap_8 FILLER_68_3523 ();
 sg13g2_fill_1 FILLER_68_3530 ();
 sg13g2_fill_2 FILLER_68_3541 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_4 FILLER_69_35 ();
 sg13g2_fill_2 FILLER_69_39 ();
 sg13g2_fill_2 FILLER_69_45 ();
 sg13g2_fill_1 FILLER_69_47 ();
 sg13g2_fill_2 FILLER_69_57 ();
 sg13g2_fill_1 FILLER_69_59 ();
 sg13g2_fill_2 FILLER_69_181 ();
 sg13g2_fill_1 FILLER_69_201 ();
 sg13g2_fill_2 FILLER_69_254 ();
 sg13g2_decap_8 FILLER_69_296 ();
 sg13g2_decap_8 FILLER_69_303 ();
 sg13g2_decap_4 FILLER_69_310 ();
 sg13g2_fill_2 FILLER_69_314 ();
 sg13g2_fill_2 FILLER_69_337 ();
 sg13g2_fill_1 FILLER_69_365 ();
 sg13g2_decap_4 FILLER_69_395 ();
 sg13g2_fill_1 FILLER_69_444 ();
 sg13g2_fill_2 FILLER_69_453 ();
 sg13g2_fill_1 FILLER_69_455 ();
 sg13g2_decap_4 FILLER_69_465 ();
 sg13g2_fill_1 FILLER_69_469 ();
 sg13g2_fill_1 FILLER_69_478 ();
 sg13g2_decap_8 FILLER_69_487 ();
 sg13g2_decap_8 FILLER_69_494 ();
 sg13g2_fill_2 FILLER_69_514 ();
 sg13g2_fill_1 FILLER_69_516 ();
 sg13g2_decap_4 FILLER_69_539 ();
 sg13g2_fill_2 FILLER_69_543 ();
 sg13g2_decap_4 FILLER_69_554 ();
 sg13g2_fill_2 FILLER_69_558 ();
 sg13g2_fill_1 FILLER_69_563 ();
 sg13g2_decap_8 FILLER_69_577 ();
 sg13g2_decap_8 FILLER_69_611 ();
 sg13g2_decap_8 FILLER_69_618 ();
 sg13g2_fill_1 FILLER_69_638 ();
 sg13g2_fill_2 FILLER_69_652 ();
 sg13g2_fill_1 FILLER_69_654 ();
 sg13g2_fill_2 FILLER_69_665 ();
 sg13g2_fill_1 FILLER_69_667 ();
 sg13g2_decap_8 FILLER_69_680 ();
 sg13g2_fill_1 FILLER_69_687 ();
 sg13g2_fill_2 FILLER_69_714 ();
 sg13g2_fill_1 FILLER_69_731 ();
 sg13g2_fill_2 FILLER_69_745 ();
 sg13g2_fill_1 FILLER_69_747 ();
 sg13g2_decap_8 FILLER_69_769 ();
 sg13g2_fill_1 FILLER_69_776 ();
 sg13g2_fill_1 FILLER_69_811 ();
 sg13g2_fill_1 FILLER_69_841 ();
 sg13g2_decap_4 FILLER_69_859 ();
 sg13g2_decap_4 FILLER_69_880 ();
 sg13g2_fill_1 FILLER_69_884 ();
 sg13g2_fill_2 FILLER_69_893 ();
 sg13g2_fill_2 FILLER_69_912 ();
 sg13g2_fill_2 FILLER_69_933 ();
 sg13g2_fill_1 FILLER_69_935 ();
 sg13g2_decap_8 FILLER_69_965 ();
 sg13g2_fill_2 FILLER_69_990 ();
 sg13g2_fill_1 FILLER_69_992 ();
 sg13g2_decap_8 FILLER_69_1016 ();
 sg13g2_fill_2 FILLER_69_1023 ();
 sg13g2_fill_2 FILLER_69_1043 ();
 sg13g2_fill_1 FILLER_69_1045 ();
 sg13g2_fill_1 FILLER_69_1066 ();
 sg13g2_decap_8 FILLER_69_1071 ();
 sg13g2_decap_8 FILLER_69_1078 ();
 sg13g2_fill_2 FILLER_69_1101 ();
 sg13g2_decap_8 FILLER_69_1132 ();
 sg13g2_decap_4 FILLER_69_1139 ();
 sg13g2_fill_1 FILLER_69_1143 ();
 sg13g2_decap_8 FILLER_69_1165 ();
 sg13g2_fill_2 FILLER_69_1172 ();
 sg13g2_fill_1 FILLER_69_1174 ();
 sg13g2_fill_2 FILLER_69_1201 ();
 sg13g2_decap_8 FILLER_69_1220 ();
 sg13g2_decap_4 FILLER_69_1227 ();
 sg13g2_fill_2 FILLER_69_1249 ();
 sg13g2_fill_1 FILLER_69_1265 ();
 sg13g2_decap_8 FILLER_69_1279 ();
 sg13g2_decap_8 FILLER_69_1286 ();
 sg13g2_fill_1 FILLER_69_1293 ();
 sg13g2_decap_8 FILLER_69_1325 ();
 sg13g2_fill_1 FILLER_69_1332 ();
 sg13g2_fill_2 FILLER_69_1355 ();
 sg13g2_decap_8 FILLER_69_1381 ();
 sg13g2_fill_2 FILLER_69_1388 ();
 sg13g2_fill_1 FILLER_69_1390 ();
 sg13g2_fill_1 FILLER_69_1403 ();
 sg13g2_decap_8 FILLER_69_1409 ();
 sg13g2_decap_8 FILLER_69_1416 ();
 sg13g2_decap_8 FILLER_69_1423 ();
 sg13g2_decap_8 FILLER_69_1447 ();
 sg13g2_fill_2 FILLER_69_1454 ();
 sg13g2_decap_8 FILLER_69_1464 ();
 sg13g2_fill_2 FILLER_69_1471 ();
 sg13g2_fill_1 FILLER_69_1473 ();
 sg13g2_decap_4 FILLER_69_1478 ();
 sg13g2_decap_8 FILLER_69_1486 ();
 sg13g2_decap_4 FILLER_69_1505 ();
 sg13g2_fill_1 FILLER_69_1509 ();
 sg13g2_decap_8 FILLER_69_1530 ();
 sg13g2_fill_1 FILLER_69_1537 ();
 sg13g2_decap_8 FILLER_69_1543 ();
 sg13g2_fill_1 FILLER_69_1550 ();
 sg13g2_decap_8 FILLER_69_1583 ();
 sg13g2_decap_8 FILLER_69_1590 ();
 sg13g2_fill_2 FILLER_69_1597 ();
 sg13g2_decap_8 FILLER_69_1627 ();
 sg13g2_fill_1 FILLER_69_1634 ();
 sg13g2_fill_1 FILLER_69_1648 ();
 sg13g2_decap_8 FILLER_69_1668 ();
 sg13g2_decap_8 FILLER_69_1695 ();
 sg13g2_fill_2 FILLER_69_1702 ();
 sg13g2_decap_4 FILLER_69_1732 ();
 sg13g2_fill_2 FILLER_69_1736 ();
 sg13g2_decap_4 FILLER_69_1754 ();
 sg13g2_fill_1 FILLER_69_1808 ();
 sg13g2_fill_2 FILLER_69_1814 ();
 sg13g2_fill_1 FILLER_69_1854 ();
 sg13g2_fill_2 FILLER_69_1860 ();
 sg13g2_fill_1 FILLER_69_1876 ();
 sg13g2_fill_2 FILLER_69_1916 ();
 sg13g2_fill_1 FILLER_69_1918 ();
 sg13g2_fill_2 FILLER_69_1927 ();
 sg13g2_fill_2 FILLER_69_1936 ();
 sg13g2_fill_2 FILLER_69_1942 ();
 sg13g2_fill_1 FILLER_69_1944 ();
 sg13g2_fill_1 FILLER_69_1949 ();
 sg13g2_decap_8 FILLER_69_1966 ();
 sg13g2_decap_4 FILLER_69_1973 ();
 sg13g2_fill_2 FILLER_69_1977 ();
 sg13g2_decap_4 FILLER_69_2005 ();
 sg13g2_fill_1 FILLER_69_2022 ();
 sg13g2_decap_8 FILLER_69_2053 ();
 sg13g2_fill_1 FILLER_69_2060 ();
 sg13g2_fill_1 FILLER_69_2077 ();
 sg13g2_decap_8 FILLER_69_2089 ();
 sg13g2_fill_1 FILLER_69_2118 ();
 sg13g2_fill_1 FILLER_69_2127 ();
 sg13g2_fill_1 FILLER_69_2136 ();
 sg13g2_fill_2 FILLER_69_2141 ();
 sg13g2_fill_2 FILLER_69_2148 ();
 sg13g2_fill_1 FILLER_69_2176 ();
 sg13g2_fill_2 FILLER_69_2190 ();
 sg13g2_fill_1 FILLER_69_2192 ();
 sg13g2_decap_4 FILLER_69_2222 ();
 sg13g2_fill_1 FILLER_69_2226 ();
 sg13g2_fill_2 FILLER_69_2244 ();
 sg13g2_fill_2 FILLER_69_2272 ();
 sg13g2_fill_2 FILLER_69_2279 ();
 sg13g2_fill_1 FILLER_69_2281 ();
 sg13g2_fill_2 FILLER_69_2309 ();
 sg13g2_fill_2 FILLER_69_2324 ();
 sg13g2_decap_4 FILLER_69_2343 ();
 sg13g2_fill_2 FILLER_69_2347 ();
 sg13g2_decap_4 FILLER_69_2403 ();
 sg13g2_decap_4 FILLER_69_2436 ();
 sg13g2_fill_1 FILLER_69_2440 ();
 sg13g2_fill_2 FILLER_69_2506 ();
 sg13g2_fill_1 FILLER_69_2516 ();
 sg13g2_fill_1 FILLER_69_2529 ();
 sg13g2_decap_4 FILLER_69_2551 ();
 sg13g2_fill_1 FILLER_69_2555 ();
 sg13g2_fill_2 FILLER_69_2582 ();
 sg13g2_fill_1 FILLER_69_2584 ();
 sg13g2_fill_2 FILLER_69_2619 ();
 sg13g2_fill_2 FILLER_69_2638 ();
 sg13g2_fill_1 FILLER_69_2640 ();
 sg13g2_decap_8 FILLER_69_2663 ();
 sg13g2_fill_2 FILLER_69_2670 ();
 sg13g2_fill_1 FILLER_69_2672 ();
 sg13g2_decap_8 FILLER_69_2696 ();
 sg13g2_fill_2 FILLER_69_2703 ();
 sg13g2_fill_1 FILLER_69_2705 ();
 sg13g2_fill_2 FILLER_69_2710 ();
 sg13g2_fill_1 FILLER_69_2712 ();
 sg13g2_fill_2 FILLER_69_2789 ();
 sg13g2_fill_1 FILLER_69_2806 ();
 sg13g2_decap_4 FILLER_69_2826 ();
 sg13g2_fill_2 FILLER_69_2830 ();
 sg13g2_fill_1 FILLER_69_2850 ();
 sg13g2_fill_1 FILLER_69_2886 ();
 sg13g2_fill_1 FILLER_69_2942 ();
 sg13g2_fill_2 FILLER_69_2951 ();
 sg13g2_fill_1 FILLER_69_2953 ();
 sg13g2_decap_4 FILLER_69_2969 ();
 sg13g2_fill_1 FILLER_69_2973 ();
 sg13g2_fill_2 FILLER_69_2984 ();
 sg13g2_fill_1 FILLER_69_2986 ();
 sg13g2_decap_8 FILLER_69_2994 ();
 sg13g2_fill_1 FILLER_69_3001 ();
 sg13g2_decap_8 FILLER_69_3007 ();
 sg13g2_decap_4 FILLER_69_3014 ();
 sg13g2_fill_1 FILLER_69_3018 ();
 sg13g2_decap_8 FILLER_69_3023 ();
 sg13g2_decap_8 FILLER_69_3030 ();
 sg13g2_fill_2 FILLER_69_3037 ();
 sg13g2_fill_2 FILLER_69_3057 ();
 sg13g2_decap_4 FILLER_69_3080 ();
 sg13g2_fill_2 FILLER_69_3084 ();
 sg13g2_decap_4 FILLER_69_3115 ();
 sg13g2_fill_1 FILLER_69_3119 ();
 sg13g2_fill_1 FILLER_69_3163 ();
 sg13g2_fill_2 FILLER_69_3178 ();
 sg13g2_fill_1 FILLER_69_3180 ();
 sg13g2_fill_1 FILLER_69_3192 ();
 sg13g2_fill_2 FILLER_69_3256 ();
 sg13g2_decap_4 FILLER_69_3283 ();
 sg13g2_fill_2 FILLER_69_3287 ();
 sg13g2_fill_2 FILLER_69_3307 ();
 sg13g2_fill_1 FILLER_69_3309 ();
 sg13g2_fill_1 FILLER_69_3365 ();
 sg13g2_fill_1 FILLER_69_3430 ();
 sg13g2_fill_1 FILLER_69_3439 ();
 sg13g2_fill_2 FILLER_69_3460 ();
 sg13g2_fill_1 FILLER_69_3470 ();
 sg13g2_fill_2 FILLER_69_3481 ();
 sg13g2_fill_1 FILLER_69_3483 ();
 sg13g2_decap_8 FILLER_69_3503 ();
 sg13g2_fill_1 FILLER_69_3510 ();
 sg13g2_fill_1 FILLER_69_3579 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_fill_1 FILLER_70_49 ();
 sg13g2_fill_1 FILLER_70_54 ();
 sg13g2_fill_2 FILLER_70_68 ();
 sg13g2_decap_4 FILLER_70_108 ();
 sg13g2_fill_2 FILLER_70_112 ();
 sg13g2_fill_1 FILLER_70_195 ();
 sg13g2_decap_4 FILLER_70_250 ();
 sg13g2_fill_2 FILLER_70_278 ();
 sg13g2_fill_2 FILLER_70_313 ();
 sg13g2_fill_1 FILLER_70_320 ();
 sg13g2_decap_8 FILLER_70_326 ();
 sg13g2_decap_8 FILLER_70_333 ();
 sg13g2_fill_1 FILLER_70_340 ();
 sg13g2_fill_1 FILLER_70_346 ();
 sg13g2_decap_8 FILLER_70_360 ();
 sg13g2_fill_2 FILLER_70_367 ();
 sg13g2_decap_8 FILLER_70_382 ();
 sg13g2_fill_2 FILLER_70_389 ();
 sg13g2_decap_8 FILLER_70_408 ();
 sg13g2_fill_1 FILLER_70_415 ();
 sg13g2_fill_2 FILLER_70_421 ();
 sg13g2_fill_1 FILLER_70_423 ();
 sg13g2_fill_2 FILLER_70_442 ();
 sg13g2_fill_1 FILLER_70_460 ();
 sg13g2_fill_2 FILLER_70_475 ();
 sg13g2_fill_1 FILLER_70_482 ();
 sg13g2_decap_4 FILLER_70_493 ();
 sg13g2_fill_1 FILLER_70_497 ();
 sg13g2_fill_1 FILLER_70_513 ();
 sg13g2_decap_8 FILLER_70_525 ();
 sg13g2_decap_4 FILLER_70_532 ();
 sg13g2_fill_1 FILLER_70_536 ();
 sg13g2_fill_1 FILLER_70_558 ();
 sg13g2_decap_8 FILLER_70_586 ();
 sg13g2_fill_2 FILLER_70_593 ();
 sg13g2_fill_2 FILLER_70_608 ();
 sg13g2_fill_2 FILLER_70_658 ();
 sg13g2_decap_8 FILLER_70_732 ();
 sg13g2_decap_4 FILLER_70_739 ();
 sg13g2_fill_1 FILLER_70_743 ();
 sg13g2_fill_1 FILLER_70_779 ();
 sg13g2_decap_4 FILLER_70_795 ();
 sg13g2_fill_1 FILLER_70_812 ();
 sg13g2_fill_1 FILLER_70_821 ();
 sg13g2_decap_8 FILLER_70_843 ();
 sg13g2_decap_8 FILLER_70_850 ();
 sg13g2_fill_1 FILLER_70_857 ();
 sg13g2_fill_2 FILLER_70_874 ();
 sg13g2_fill_1 FILLER_70_876 ();
 sg13g2_fill_2 FILLER_70_908 ();
 sg13g2_fill_2 FILLER_70_917 ();
 sg13g2_decap_8 FILLER_70_943 ();
 sg13g2_fill_2 FILLER_70_950 ();
 sg13g2_fill_1 FILLER_70_952 ();
 sg13g2_decap_8 FILLER_70_959 ();
 sg13g2_decap_4 FILLER_70_966 ();
 sg13g2_fill_1 FILLER_70_970 ();
 sg13g2_fill_2 FILLER_70_993 ();
 sg13g2_fill_2 FILLER_70_1025 ();
 sg13g2_fill_1 FILLER_70_1031 ();
 sg13g2_fill_2 FILLER_70_1036 ();
 sg13g2_fill_2 FILLER_70_1052 ();
 sg13g2_fill_1 FILLER_70_1054 ();
 sg13g2_fill_1 FILLER_70_1080 ();
 sg13g2_decap_4 FILLER_70_1106 ();
 sg13g2_fill_2 FILLER_70_1110 ();
 sg13g2_fill_2 FILLER_70_1122 ();
 sg13g2_decap_8 FILLER_70_1132 ();
 sg13g2_fill_1 FILLER_70_1139 ();
 sg13g2_fill_2 FILLER_70_1163 ();
 sg13g2_fill_1 FILLER_70_1182 ();
 sg13g2_fill_2 FILLER_70_1196 ();
 sg13g2_fill_1 FILLER_70_1198 ();
 sg13g2_fill_1 FILLER_70_1215 ();
 sg13g2_decap_4 FILLER_70_1241 ();
 sg13g2_fill_2 FILLER_70_1245 ();
 sg13g2_decap_4 FILLER_70_1252 ();
 sg13g2_fill_2 FILLER_70_1256 ();
 sg13g2_decap_4 FILLER_70_1296 ();
 sg13g2_fill_1 FILLER_70_1300 ();
 sg13g2_fill_2 FILLER_70_1310 ();
 sg13g2_fill_1 FILLER_70_1325 ();
 sg13g2_fill_2 FILLER_70_1356 ();
 sg13g2_fill_1 FILLER_70_1358 ();
 sg13g2_decap_8 FILLER_70_1387 ();
 sg13g2_decap_4 FILLER_70_1394 ();
 sg13g2_fill_1 FILLER_70_1398 ();
 sg13g2_fill_2 FILLER_70_1427 ();
 sg13g2_fill_1 FILLER_70_1429 ();
 sg13g2_fill_1 FILLER_70_1497 ();
 sg13g2_fill_2 FILLER_70_1511 ();
 sg13g2_fill_2 FILLER_70_1518 ();
 sg13g2_fill_2 FILLER_70_1555 ();
 sg13g2_decap_8 FILLER_70_1571 ();
 sg13g2_decap_4 FILLER_70_1587 ();
 sg13g2_fill_1 FILLER_70_1596 ();
 sg13g2_fill_1 FILLER_70_1604 ();
 sg13g2_decap_8 FILLER_70_1609 ();
 sg13g2_decap_8 FILLER_70_1616 ();
 sg13g2_fill_1 FILLER_70_1623 ();
 sg13g2_decap_8 FILLER_70_1637 ();
 sg13g2_decap_8 FILLER_70_1644 ();
 sg13g2_fill_2 FILLER_70_1695 ();
 sg13g2_fill_2 FILLER_70_1706 ();
 sg13g2_fill_2 FILLER_70_1720 ();
 sg13g2_decap_8 FILLER_70_1730 ();
 sg13g2_decap_4 FILLER_70_1737 ();
 sg13g2_fill_1 FILLER_70_1741 ();
 sg13g2_fill_2 FILLER_70_1777 ();
 sg13g2_fill_1 FILLER_70_1795 ();
 sg13g2_fill_1 FILLER_70_1809 ();
 sg13g2_decap_8 FILLER_70_1815 ();
 sg13g2_fill_2 FILLER_70_1822 ();
 sg13g2_decap_8 FILLER_70_1848 ();
 sg13g2_fill_2 FILLER_70_1855 ();
 sg13g2_fill_1 FILLER_70_1857 ();
 sg13g2_decap_4 FILLER_70_1883 ();
 sg13g2_decap_8 FILLER_70_1891 ();
 sg13g2_fill_2 FILLER_70_1898 ();
 sg13g2_fill_2 FILLER_70_1939 ();
 sg13g2_fill_1 FILLER_70_1941 ();
 sg13g2_fill_2 FILLER_70_1950 ();
 sg13g2_decap_4 FILLER_70_1968 ();
 sg13g2_fill_1 FILLER_70_1972 ();
 sg13g2_fill_2 FILLER_70_1999 ();
 sg13g2_fill_1 FILLER_70_2001 ();
 sg13g2_fill_2 FILLER_70_2015 ();
 sg13g2_fill_1 FILLER_70_2021 ();
 sg13g2_fill_1 FILLER_70_2035 ();
 sg13g2_decap_4 FILLER_70_2046 ();
 sg13g2_fill_1 FILLER_70_2050 ();
 sg13g2_fill_1 FILLER_70_2073 ();
 sg13g2_decap_8 FILLER_70_2089 ();
 sg13g2_decap_4 FILLER_70_2096 ();
 sg13g2_fill_1 FILLER_70_2100 ();
 sg13g2_decap_8 FILLER_70_2118 ();
 sg13g2_fill_2 FILLER_70_2125 ();
 sg13g2_fill_1 FILLER_70_2127 ();
 sg13g2_decap_8 FILLER_70_2132 ();
 sg13g2_decap_4 FILLER_70_2139 ();
 sg13g2_decap_8 FILLER_70_2149 ();
 sg13g2_fill_1 FILLER_70_2156 ();
 sg13g2_fill_2 FILLER_70_2183 ();
 sg13g2_fill_1 FILLER_70_2232 ();
 sg13g2_decap_4 FILLER_70_2241 ();
 sg13g2_fill_2 FILLER_70_2260 ();
 sg13g2_fill_1 FILLER_70_2262 ();
 sg13g2_decap_8 FILLER_70_2290 ();
 sg13g2_fill_2 FILLER_70_2297 ();
 sg13g2_fill_1 FILLER_70_2299 ();
 sg13g2_fill_1 FILLER_70_2346 ();
 sg13g2_fill_2 FILLER_70_2351 ();
 sg13g2_decap_8 FILLER_70_2366 ();
 sg13g2_fill_2 FILLER_70_2373 ();
 sg13g2_decap_4 FILLER_70_2388 ();
 sg13g2_decap_8 FILLER_70_2410 ();
 sg13g2_fill_1 FILLER_70_2424 ();
 sg13g2_fill_2 FILLER_70_2438 ();
 sg13g2_fill_1 FILLER_70_2440 ();
 sg13g2_decap_4 FILLER_70_2462 ();
 sg13g2_fill_1 FILLER_70_2484 ();
 sg13g2_fill_1 FILLER_70_2498 ();
 sg13g2_fill_1 FILLER_70_2514 ();
 sg13g2_fill_2 FILLER_70_2525 ();
 sg13g2_fill_1 FILLER_70_2527 ();
 sg13g2_decap_4 FILLER_70_2564 ();
 sg13g2_fill_1 FILLER_70_2568 ();
 sg13g2_fill_1 FILLER_70_2577 ();
 sg13g2_fill_2 FILLER_70_2614 ();
 sg13g2_fill_2 FILLER_70_2629 ();
 sg13g2_fill_1 FILLER_70_2644 ();
 sg13g2_fill_2 FILLER_70_2666 ();
 sg13g2_fill_2 FILLER_70_2702 ();
 sg13g2_fill_2 FILLER_70_2721 ();
 sg13g2_decap_8 FILLER_70_2727 ();
 sg13g2_fill_1 FILLER_70_2734 ();
 sg13g2_decap_8 FILLER_70_2744 ();
 sg13g2_decap_4 FILLER_70_2751 ();
 sg13g2_fill_2 FILLER_70_2755 ();
 sg13g2_fill_1 FILLER_70_2782 ();
 sg13g2_decap_8 FILLER_70_2795 ();
 sg13g2_fill_1 FILLER_70_2802 ();
 sg13g2_decap_8 FILLER_70_2844 ();
 sg13g2_decap_8 FILLER_70_2851 ();
 sg13g2_decap_4 FILLER_70_2858 ();
 sg13g2_fill_2 FILLER_70_2867 ();
 sg13g2_fill_1 FILLER_70_2869 ();
 sg13g2_decap_8 FILLER_70_2883 ();
 sg13g2_fill_1 FILLER_70_2959 ();
 sg13g2_decap_8 FILLER_70_2967 ();
 sg13g2_fill_1 FILLER_70_2995 ();
 sg13g2_decap_8 FILLER_70_3008 ();
 sg13g2_fill_2 FILLER_70_3015 ();
 sg13g2_fill_1 FILLER_70_3021 ();
 sg13g2_fill_1 FILLER_70_3067 ();
 sg13g2_fill_2 FILLER_70_3076 ();
 sg13g2_fill_1 FILLER_70_3078 ();
 sg13g2_fill_2 FILLER_70_3093 ();
 sg13g2_fill_1 FILLER_70_3095 ();
 sg13g2_fill_2 FILLER_70_3114 ();
 sg13g2_fill_1 FILLER_70_3116 ();
 sg13g2_fill_2 FILLER_70_3127 ();
 sg13g2_decap_8 FILLER_70_3137 ();
 sg13g2_fill_2 FILLER_70_3158 ();
 sg13g2_decap_8 FILLER_70_3178 ();
 sg13g2_decap_4 FILLER_70_3185 ();
 sg13g2_fill_2 FILLER_70_3189 ();
 sg13g2_decap_8 FILLER_70_3278 ();
 sg13g2_fill_2 FILLER_70_3285 ();
 sg13g2_fill_1 FILLER_70_3287 ();
 sg13g2_decap_4 FILLER_70_3313 ();
 sg13g2_fill_1 FILLER_70_3325 ();
 sg13g2_fill_2 FILLER_70_3392 ();
 sg13g2_fill_1 FILLER_70_3410 ();
 sg13g2_decap_4 FILLER_70_3446 ();
 sg13g2_fill_1 FILLER_70_3450 ();
 sg13g2_decap_8 FILLER_70_3467 ();
 sg13g2_decap_4 FILLER_70_3474 ();
 sg13g2_fill_1 FILLER_70_3478 ();
 sg13g2_decap_4 FILLER_70_3497 ();
 sg13g2_fill_1 FILLER_70_3501 ();
 sg13g2_fill_1 FILLER_70_3538 ();
 sg13g2_fill_2 FILLER_70_3561 ();
 sg13g2_fill_1 FILLER_70_3563 ();
 sg13g2_decap_8 FILLER_70_3573 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_4 FILLER_71_42 ();
 sg13g2_decap_4 FILLER_71_83 ();
 sg13g2_fill_2 FILLER_71_152 ();
 sg13g2_fill_2 FILLER_71_232 ();
 sg13g2_fill_1 FILLER_71_234 ();
 sg13g2_fill_2 FILLER_71_278 ();
 sg13g2_fill_2 FILLER_71_288 ();
 sg13g2_decap_4 FILLER_71_298 ();
 sg13g2_fill_2 FILLER_71_302 ();
 sg13g2_decap_8 FILLER_71_356 ();
 sg13g2_decap_8 FILLER_71_388 ();
 sg13g2_fill_2 FILLER_71_395 ();
 sg13g2_decap_8 FILLER_71_442 ();
 sg13g2_fill_2 FILLER_71_449 ();
 sg13g2_fill_2 FILLER_71_465 ();
 sg13g2_fill_1 FILLER_71_467 ();
 sg13g2_decap_8 FILLER_71_483 ();
 sg13g2_decap_8 FILLER_71_490 ();
 sg13g2_decap_4 FILLER_71_497 ();
 sg13g2_fill_1 FILLER_71_501 ();
 sg13g2_fill_1 FILLER_71_509 ();
 sg13g2_fill_2 FILLER_71_518 ();
 sg13g2_fill_1 FILLER_71_520 ();
 sg13g2_fill_1 FILLER_71_547 ();
 sg13g2_fill_1 FILLER_71_553 ();
 sg13g2_fill_1 FILLER_71_562 ();
 sg13g2_fill_1 FILLER_71_568 ();
 sg13g2_fill_1 FILLER_71_579 ();
 sg13g2_fill_1 FILLER_71_601 ();
 sg13g2_decap_8 FILLER_71_611 ();
 sg13g2_decap_8 FILLER_71_618 ();
 sg13g2_fill_1 FILLER_71_625 ();
 sg13g2_fill_2 FILLER_71_647 ();
 sg13g2_fill_1 FILLER_71_649 ();
 sg13g2_fill_1 FILLER_71_666 ();
 sg13g2_fill_1 FILLER_71_672 ();
 sg13g2_fill_1 FILLER_71_682 ();
 sg13g2_fill_1 FILLER_71_716 ();
 sg13g2_decap_4 FILLER_71_723 ();
 sg13g2_fill_1 FILLER_71_727 ();
 sg13g2_fill_1 FILLER_71_736 ();
 sg13g2_decap_8 FILLER_71_747 ();
 sg13g2_fill_2 FILLER_71_754 ();
 sg13g2_decap_8 FILLER_71_769 ();
 sg13g2_decap_4 FILLER_71_776 ();
 sg13g2_decap_8 FILLER_71_797 ();
 sg13g2_fill_2 FILLER_71_804 ();
 sg13g2_fill_1 FILLER_71_806 ();
 sg13g2_fill_1 FILLER_71_819 ();
 sg13g2_decap_8 FILLER_71_836 ();
 sg13g2_decap_8 FILLER_71_843 ();
 sg13g2_decap_4 FILLER_71_850 ();
 sg13g2_fill_1 FILLER_71_854 ();
 sg13g2_decap_4 FILLER_71_879 ();
 sg13g2_fill_1 FILLER_71_900 ();
 sg13g2_fill_2 FILLER_71_906 ();
 sg13g2_decap_8 FILLER_71_915 ();
 sg13g2_fill_2 FILLER_71_922 ();
 sg13g2_decap_4 FILLER_71_927 ();
 sg13g2_fill_1 FILLER_71_931 ();
 sg13g2_fill_2 FILLER_71_941 ();
 sg13g2_fill_1 FILLER_71_943 ();
 sg13g2_fill_2 FILLER_71_947 ();
 sg13g2_fill_1 FILLER_71_949 ();
 sg13g2_decap_8 FILLER_71_965 ();
 sg13g2_decap_4 FILLER_71_972 ();
 sg13g2_decap_8 FILLER_71_992 ();
 sg13g2_fill_2 FILLER_71_999 ();
 sg13g2_fill_1 FILLER_71_1006 ();
 sg13g2_decap_8 FILLER_71_1020 ();
 sg13g2_decap_4 FILLER_71_1027 ();
 sg13g2_fill_2 FILLER_71_1031 ();
 sg13g2_decap_4 FILLER_71_1046 ();
 sg13g2_fill_1 FILLER_71_1055 ();
 sg13g2_fill_2 FILLER_71_1082 ();
 sg13g2_fill_1 FILLER_71_1100 ();
 sg13g2_decap_8 FILLER_71_1111 ();
 sg13g2_fill_1 FILLER_71_1133 ();
 sg13g2_fill_2 FILLER_71_1144 ();
 sg13g2_fill_2 FILLER_71_1196 ();
 sg13g2_decap_4 FILLER_71_1219 ();
 sg13g2_fill_2 FILLER_71_1238 ();
 sg13g2_fill_2 FILLER_71_1260 ();
 sg13g2_fill_2 FILLER_71_1269 ();
 sg13g2_decap_8 FILLER_71_1279 ();
 sg13g2_fill_2 FILLER_71_1286 ();
 sg13g2_fill_1 FILLER_71_1288 ();
 sg13g2_decap_4 FILLER_71_1297 ();
 sg13g2_fill_1 FILLER_71_1301 ();
 sg13g2_decap_4 FILLER_71_1333 ();
 sg13g2_fill_1 FILLER_71_1342 ();
 sg13g2_decap_8 FILLER_71_1356 ();
 sg13g2_decap_8 FILLER_71_1363 ();
 sg13g2_fill_2 FILLER_71_1370 ();
 sg13g2_decap_4 FILLER_71_1375 ();
 sg13g2_fill_1 FILLER_71_1389 ();
 sg13g2_fill_1 FILLER_71_1405 ();
 sg13g2_fill_2 FILLER_71_1414 ();
 sg13g2_decap_4 FILLER_71_1425 ();
 sg13g2_decap_8 FILLER_71_1466 ();
 sg13g2_fill_2 FILLER_71_1473 ();
 sg13g2_fill_2 FILLER_71_1531 ();
 sg13g2_fill_1 FILLER_71_1537 ();
 sg13g2_decap_8 FILLER_71_1606 ();
 sg13g2_fill_2 FILLER_71_1651 ();
 sg13g2_fill_1 FILLER_71_1653 ();
 sg13g2_fill_2 FILLER_71_1676 ();
 sg13g2_decap_8 FILLER_71_1695 ();
 sg13g2_decap_8 FILLER_71_1702 ();
 sg13g2_decap_8 FILLER_71_1709 ();
 sg13g2_fill_2 FILLER_71_1716 ();
 sg13g2_fill_2 FILLER_71_1722 ();
 sg13g2_fill_1 FILLER_71_1724 ();
 sg13g2_decap_8 FILLER_71_1734 ();
 sg13g2_fill_2 FILLER_71_1759 ();
 sg13g2_fill_1 FILLER_71_1761 ();
 sg13g2_decap_8 FILLER_71_1775 ();
 sg13g2_fill_1 FILLER_71_1794 ();
 sg13g2_fill_1 FILLER_71_1816 ();
 sg13g2_decap_4 FILLER_71_1821 ();
 sg13g2_fill_1 FILLER_71_1825 ();
 sg13g2_decap_4 FILLER_71_1840 ();
 sg13g2_fill_1 FILLER_71_1844 ();
 sg13g2_decap_8 FILLER_71_1861 ();
 sg13g2_fill_2 FILLER_71_1868 ();
 sg13g2_fill_1 FILLER_71_1879 ();
 sg13g2_decap_8 FILLER_71_1893 ();
 sg13g2_fill_2 FILLER_71_1900 ();
 sg13g2_fill_1 FILLER_71_1902 ();
 sg13g2_fill_1 FILLER_71_1915 ();
 sg13g2_decap_4 FILLER_71_1925 ();
 sg13g2_fill_1 FILLER_71_1929 ();
 sg13g2_fill_2 FILLER_71_1935 ();
 sg13g2_fill_2 FILLER_71_1954 ();
 sg13g2_fill_1 FILLER_71_1956 ();
 sg13g2_decap_4 FILLER_71_1966 ();
 sg13g2_fill_1 FILLER_71_1970 ();
 sg13g2_fill_2 FILLER_71_1978 ();
 sg13g2_decap_8 FILLER_71_2053 ();
 sg13g2_fill_2 FILLER_71_2060 ();
 sg13g2_fill_1 FILLER_71_2062 ();
 sg13g2_decap_8 FILLER_71_2085 ();
 sg13g2_decap_8 FILLER_71_2157 ();
 sg13g2_fill_2 FILLER_71_2164 ();
 sg13g2_decap_4 FILLER_71_2197 ();
 sg13g2_fill_2 FILLER_71_2244 ();
 sg13g2_decap_8 FILLER_71_2311 ();
 sg13g2_decap_8 FILLER_71_2318 ();
 sg13g2_fill_1 FILLER_71_2338 ();
 sg13g2_fill_1 FILLER_71_2370 ();
 sg13g2_decap_8 FILLER_71_2444 ();
 sg13g2_fill_2 FILLER_71_2503 ();
 sg13g2_fill_1 FILLER_71_2505 ();
 sg13g2_fill_2 FILLER_71_2523 ();
 sg13g2_fill_1 FILLER_71_2525 ();
 sg13g2_decap_4 FILLER_71_2552 ();
 sg13g2_fill_1 FILLER_71_2556 ();
 sg13g2_decap_8 FILLER_71_2580 ();
 sg13g2_decap_8 FILLER_71_2600 ();
 sg13g2_decap_4 FILLER_71_2607 ();
 sg13g2_fill_2 FILLER_71_2616 ();
 sg13g2_decap_8 FILLER_71_2623 ();
 sg13g2_fill_1 FILLER_71_2648 ();
 sg13g2_decap_4 FILLER_71_2665 ();
 sg13g2_fill_2 FILLER_71_2669 ();
 sg13g2_fill_1 FILLER_71_2709 ();
 sg13g2_fill_2 FILLER_71_2728 ();
 sg13g2_decap_4 FILLER_71_2748 ();
 sg13g2_fill_2 FILLER_71_2782 ();
 sg13g2_fill_1 FILLER_71_2804 ();
 sg13g2_decap_4 FILLER_71_2809 ();
 sg13g2_fill_2 FILLER_71_2813 ();
 sg13g2_decap_8 FILLER_71_2822 ();
 sg13g2_fill_2 FILLER_71_2829 ();
 sg13g2_fill_1 FILLER_71_2831 ();
 sg13g2_fill_2 FILLER_71_2836 ();
 sg13g2_fill_2 FILLER_71_2843 ();
 sg13g2_fill_1 FILLER_71_2845 ();
 sg13g2_fill_1 FILLER_71_2885 ();
 sg13g2_fill_1 FILLER_71_2925 ();
 sg13g2_fill_2 FILLER_71_2934 ();
 sg13g2_decap_4 FILLER_71_2952 ();
 sg13g2_fill_1 FILLER_71_2956 ();
 sg13g2_fill_1 FILLER_71_2965 ();
 sg13g2_fill_2 FILLER_71_2982 ();
 sg13g2_decap_4 FILLER_71_2994 ();
 sg13g2_decap_4 FILLER_71_3005 ();
 sg13g2_fill_1 FILLER_71_3009 ();
 sg13g2_fill_1 FILLER_71_3035 ();
 sg13g2_decap_8 FILLER_71_3053 ();
 sg13g2_decap_4 FILLER_71_3060 ();
 sg13g2_fill_2 FILLER_71_3064 ();
 sg13g2_fill_2 FILLER_71_3077 ();
 sg13g2_fill_2 FILLER_71_3089 ();
 sg13g2_fill_1 FILLER_71_3108 ();
 sg13g2_decap_4 FILLER_71_3142 ();
 sg13g2_fill_1 FILLER_71_3146 ();
 sg13g2_fill_2 FILLER_71_3157 ();
 sg13g2_decap_8 FILLER_71_3169 ();
 sg13g2_fill_2 FILLER_71_3176 ();
 sg13g2_fill_1 FILLER_71_3178 ();
 sg13g2_fill_1 FILLER_71_3183 ();
 sg13g2_decap_8 FILLER_71_3248 ();
 sg13g2_decap_4 FILLER_71_3342 ();
 sg13g2_fill_2 FILLER_71_3346 ();
 sg13g2_fill_1 FILLER_71_3361 ();
 sg13g2_fill_2 FILLER_71_3366 ();
 sg13g2_fill_1 FILLER_71_3377 ();
 sg13g2_fill_2 FILLER_71_3399 ();
 sg13g2_fill_2 FILLER_71_3414 ();
 sg13g2_fill_1 FILLER_71_3416 ();
 sg13g2_fill_2 FILLER_71_3429 ();
 sg13g2_fill_2 FILLER_71_3436 ();
 sg13g2_fill_1 FILLER_71_3438 ();
 sg13g2_decap_8 FILLER_71_3470 ();
 sg13g2_fill_2 FILLER_71_3477 ();
 sg13g2_decap_8 FILLER_71_3484 ();
 sg13g2_fill_2 FILLER_71_3491 ();
 sg13g2_fill_1 FILLER_71_3493 ();
 sg13g2_decap_4 FILLER_71_3505 ();
 sg13g2_decap_4 FILLER_71_3514 ();
 sg13g2_fill_1 FILLER_71_3518 ();
 sg13g2_decap_8 FILLER_71_3537 ();
 sg13g2_fill_2 FILLER_71_3564 ();
 sg13g2_fill_2 FILLER_71_3578 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_fill_1 FILLER_72_86 ();
 sg13g2_fill_2 FILLER_72_152 ();
 sg13g2_fill_1 FILLER_72_198 ();
 sg13g2_fill_2 FILLER_72_204 ();
 sg13g2_fill_2 FILLER_72_219 ();
 sg13g2_fill_1 FILLER_72_221 ();
 sg13g2_fill_2 FILLER_72_230 ();
 sg13g2_fill_1 FILLER_72_232 ();
 sg13g2_fill_1 FILLER_72_274 ();
 sg13g2_fill_1 FILLER_72_284 ();
 sg13g2_fill_1 FILLER_72_304 ();
 sg13g2_decap_8 FILLER_72_327 ();
 sg13g2_decap_4 FILLER_72_334 ();
 sg13g2_decap_8 FILLER_72_346 ();
 sg13g2_decap_8 FILLER_72_353 ();
 sg13g2_decap_8 FILLER_72_389 ();
 sg13g2_fill_2 FILLER_72_403 ();
 sg13g2_decap_8 FILLER_72_410 ();
 sg13g2_decap_8 FILLER_72_431 ();
 sg13g2_decap_8 FILLER_72_438 ();
 sg13g2_fill_1 FILLER_72_445 ();
 sg13g2_fill_1 FILLER_72_471 ();
 sg13g2_decap_8 FILLER_72_492 ();
 sg13g2_decap_8 FILLER_72_526 ();
 sg13g2_decap_4 FILLER_72_546 ();
 sg13g2_fill_2 FILLER_72_558 ();
 sg13g2_decap_8 FILLER_72_585 ();
 sg13g2_decap_8 FILLER_72_592 ();
 sg13g2_fill_1 FILLER_72_599 ();
 sg13g2_fill_2 FILLER_72_616 ();
 sg13g2_decap_4 FILLER_72_650 ();
 sg13g2_fill_2 FILLER_72_654 ();
 sg13g2_decap_8 FILLER_72_691 ();
 sg13g2_fill_2 FILLER_72_711 ();
 sg13g2_fill_1 FILLER_72_721 ();
 sg13g2_fill_1 FILLER_72_739 ();
 sg13g2_fill_1 FILLER_72_750 ();
 sg13g2_fill_2 FILLER_72_778 ();
 sg13g2_fill_1 FILLER_72_780 ();
 sg13g2_decap_4 FILLER_72_802 ();
 sg13g2_fill_2 FILLER_72_806 ();
 sg13g2_fill_2 FILLER_72_833 ();
 sg13g2_fill_2 FILLER_72_839 ();
 sg13g2_fill_1 FILLER_72_841 ();
 sg13g2_decap_8 FILLER_72_850 ();
 sg13g2_fill_2 FILLER_72_857 ();
 sg13g2_fill_1 FILLER_72_859 ();
 sg13g2_fill_2 FILLER_72_877 ();
 sg13g2_fill_1 FILLER_72_879 ();
 sg13g2_decap_8 FILLER_72_905 ();
 sg13g2_decap_4 FILLER_72_912 ();
 sg13g2_fill_1 FILLER_72_922 ();
 sg13g2_fill_1 FILLER_72_948 ();
 sg13g2_fill_2 FILLER_72_974 ();
 sg13g2_fill_1 FILLER_72_976 ();
 sg13g2_fill_1 FILLER_72_981 ();
 sg13g2_fill_2 FILLER_72_987 ();
 sg13g2_fill_1 FILLER_72_1002 ();
 sg13g2_decap_4 FILLER_72_1019 ();
 sg13g2_fill_1 FILLER_72_1031 ();
 sg13g2_fill_1 FILLER_72_1039 ();
 sg13g2_decap_8 FILLER_72_1049 ();
 sg13g2_decap_4 FILLER_72_1077 ();
 sg13g2_fill_1 FILLER_72_1081 ();
 sg13g2_decap_8 FILLER_72_1107 ();
 sg13g2_fill_2 FILLER_72_1114 ();
 sg13g2_fill_1 FILLER_72_1116 ();
 sg13g2_decap_4 FILLER_72_1121 ();
 sg13g2_decap_8 FILLER_72_1146 ();
 sg13g2_decap_8 FILLER_72_1153 ();
 sg13g2_decap_4 FILLER_72_1160 ();
 sg13g2_fill_2 FILLER_72_1164 ();
 sg13g2_fill_2 FILLER_72_1204 ();
 sg13g2_fill_1 FILLER_72_1206 ();
 sg13g2_fill_2 FILLER_72_1211 ();
 sg13g2_fill_2 FILLER_72_1221 ();
 sg13g2_fill_1 FILLER_72_1223 ();
 sg13g2_decap_4 FILLER_72_1228 ();
 sg13g2_fill_1 FILLER_72_1243 ();
 sg13g2_decap_4 FILLER_72_1256 ();
 sg13g2_fill_1 FILLER_72_1260 ();
 sg13g2_decap_4 FILLER_72_1274 ();
 sg13g2_fill_2 FILLER_72_1278 ();
 sg13g2_fill_2 FILLER_72_1298 ();
 sg13g2_decap_8 FILLER_72_1323 ();
 sg13g2_fill_1 FILLER_72_1330 ();
 sg13g2_fill_1 FILLER_72_1336 ();
 sg13g2_fill_2 FILLER_72_1350 ();
 sg13g2_fill_1 FILLER_72_1352 ();
 sg13g2_decap_4 FILLER_72_1357 ();
 sg13g2_fill_2 FILLER_72_1366 ();
 sg13g2_decap_4 FILLER_72_1388 ();
 sg13g2_decap_4 FILLER_72_1402 ();
 sg13g2_fill_2 FILLER_72_1410 ();
 sg13g2_fill_1 FILLER_72_1412 ();
 sg13g2_fill_2 FILLER_72_1421 ();
 sg13g2_fill_1 FILLER_72_1423 ();
 sg13g2_decap_4 FILLER_72_1437 ();
 sg13g2_fill_2 FILLER_72_1441 ();
 sg13g2_fill_1 FILLER_72_1447 ();
 sg13g2_decap_8 FILLER_72_1458 ();
 sg13g2_fill_2 FILLER_72_1481 ();
 sg13g2_fill_1 FILLER_72_1497 ();
 sg13g2_decap_4 FILLER_72_1507 ();
 sg13g2_fill_2 FILLER_72_1511 ();
 sg13g2_fill_2 FILLER_72_1518 ();
 sg13g2_fill_1 FILLER_72_1520 ();
 sg13g2_decap_8 FILLER_72_1531 ();
 sg13g2_fill_2 FILLER_72_1538 ();
 sg13g2_fill_1 FILLER_72_1540 ();
 sg13g2_decap_4 FILLER_72_1551 ();
 sg13g2_fill_2 FILLER_72_1555 ();
 sg13g2_decap_8 FILLER_72_1570 ();
 sg13g2_fill_2 FILLER_72_1577 ();
 sg13g2_fill_1 FILLER_72_1579 ();
 sg13g2_fill_1 FILLER_72_1624 ();
 sg13g2_fill_1 FILLER_72_1659 ();
 sg13g2_fill_1 FILLER_72_1677 ();
 sg13g2_fill_1 FILLER_72_1719 ();
 sg13g2_decap_8 FILLER_72_1753 ();
 sg13g2_fill_1 FILLER_72_1760 ();
 sg13g2_decap_8 FILLER_72_1789 ();
 sg13g2_decap_4 FILLER_72_1796 ();
 sg13g2_fill_1 FILLER_72_1800 ();
 sg13g2_decap_8 FILLER_72_1805 ();
 sg13g2_fill_2 FILLER_72_1817 ();
 sg13g2_fill_1 FILLER_72_1819 ();
 sg13g2_fill_2 FILLER_72_1833 ();
 sg13g2_decap_4 FILLER_72_1843 ();
 sg13g2_decap_4 FILLER_72_1856 ();
 sg13g2_decap_8 FILLER_72_1867 ();
 sg13g2_fill_2 FILLER_72_1874 ();
 sg13g2_fill_2 FILLER_72_1928 ();
 sg13g2_fill_1 FILLER_72_1930 ();
 sg13g2_fill_1 FILLER_72_1997 ();
 sg13g2_fill_2 FILLER_72_2002 ();
 sg13g2_fill_2 FILLER_72_2018 ();
 sg13g2_fill_2 FILLER_72_2029 ();
 sg13g2_fill_2 FILLER_72_2059 ();
 sg13g2_fill_1 FILLER_72_2061 ();
 sg13g2_decap_8 FILLER_72_2118 ();
 sg13g2_decap_4 FILLER_72_2125 ();
 sg13g2_fill_2 FILLER_72_2129 ();
 sg13g2_decap_4 FILLER_72_2134 ();
 sg13g2_fill_2 FILLER_72_2149 ();
 sg13g2_fill_2 FILLER_72_2179 ();
 sg13g2_fill_1 FILLER_72_2226 ();
 sg13g2_fill_1 FILLER_72_2264 ();
 sg13g2_decap_8 FILLER_72_2270 ();
 sg13g2_fill_1 FILLER_72_2277 ();
 sg13g2_decap_8 FILLER_72_2291 ();
 sg13g2_fill_2 FILLER_72_2298 ();
 sg13g2_fill_1 FILLER_72_2300 ();
 sg13g2_fill_1 FILLER_72_2329 ();
 sg13g2_decap_8 FILLER_72_2358 ();
 sg13g2_fill_2 FILLER_72_2365 ();
 sg13g2_fill_1 FILLER_72_2367 ();
 sg13g2_fill_2 FILLER_72_2381 ();
 sg13g2_fill_1 FILLER_72_2383 ();
 sg13g2_fill_2 FILLER_72_2415 ();
 sg13g2_decap_8 FILLER_72_2435 ();
 sg13g2_decap_4 FILLER_72_2442 ();
 sg13g2_fill_1 FILLER_72_2446 ();
 sg13g2_decap_4 FILLER_72_2465 ();
 sg13g2_decap_8 FILLER_72_2473 ();
 sg13g2_fill_2 FILLER_72_2480 ();
 sg13g2_fill_2 FILLER_72_2489 ();
 sg13g2_fill_2 FILLER_72_2496 ();
 sg13g2_decap_8 FILLER_72_2516 ();
 sg13g2_fill_2 FILLER_72_2553 ();
 sg13g2_decap_8 FILLER_72_2592 ();
 sg13g2_fill_2 FILLER_72_2599 ();
 sg13g2_fill_2 FILLER_72_2645 ();
 sg13g2_fill_1 FILLER_72_2647 ();
 sg13g2_decap_4 FILLER_72_2704 ();
 sg13g2_fill_2 FILLER_72_2708 ();
 sg13g2_decap_8 FILLER_72_2722 ();
 sg13g2_decap_4 FILLER_72_2729 ();
 sg13g2_decap_8 FILLER_72_2751 ();
 sg13g2_fill_1 FILLER_72_2758 ();
 sg13g2_decap_8 FILLER_72_2776 ();
 sg13g2_fill_2 FILLER_72_2783 ();
 sg13g2_fill_1 FILLER_72_2794 ();
 sg13g2_fill_2 FILLER_72_2803 ();
 sg13g2_fill_1 FILLER_72_2810 ();
 sg13g2_fill_2 FILLER_72_2821 ();
 sg13g2_fill_1 FILLER_72_2843 ();
 sg13g2_fill_2 FILLER_72_2876 ();
 sg13g2_fill_2 FILLER_72_2919 ();
 sg13g2_fill_2 FILLER_72_2929 ();
 sg13g2_fill_1 FILLER_72_2931 ();
 sg13g2_decap_4 FILLER_72_2947 ();
 sg13g2_fill_2 FILLER_72_2964 ();
 sg13g2_fill_1 FILLER_72_2971 ();
 sg13g2_fill_2 FILLER_72_2976 ();
 sg13g2_fill_2 FILLER_72_2991 ();
 sg13g2_decap_4 FILLER_72_3016 ();
 sg13g2_fill_2 FILLER_72_3020 ();
 sg13g2_fill_2 FILLER_72_3067 ();
 sg13g2_fill_1 FILLER_72_3090 ();
 sg13g2_fill_2 FILLER_72_3100 ();
 sg13g2_decap_8 FILLER_72_3107 ();
 sg13g2_decap_4 FILLER_72_3114 ();
 sg13g2_fill_1 FILLER_72_3118 ();
 sg13g2_fill_2 FILLER_72_3126 ();
 sg13g2_fill_2 FILLER_72_3133 ();
 sg13g2_fill_1 FILLER_72_3135 ();
 sg13g2_fill_1 FILLER_72_3146 ();
 sg13g2_fill_2 FILLER_72_3160 ();
 sg13g2_decap_8 FILLER_72_3167 ();
 sg13g2_fill_2 FILLER_72_3202 ();
 sg13g2_fill_1 FILLER_72_3204 ();
 sg13g2_decap_4 FILLER_72_3224 ();
 sg13g2_fill_1 FILLER_72_3228 ();
 sg13g2_decap_8 FILLER_72_3244 ();
 sg13g2_decap_8 FILLER_72_3251 ();
 sg13g2_fill_1 FILLER_72_3262 ();
 sg13g2_decap_8 FILLER_72_3278 ();
 sg13g2_decap_8 FILLER_72_3285 ();
 sg13g2_fill_2 FILLER_72_3318 ();
 sg13g2_fill_1 FILLER_72_3320 ();
 sg13g2_decap_8 FILLER_72_3334 ();
 sg13g2_decap_8 FILLER_72_3345 ();
 sg13g2_decap_4 FILLER_72_3352 ();
 sg13g2_fill_1 FILLER_72_3393 ();
 sg13g2_fill_1 FILLER_72_3403 ();
 sg13g2_decap_4 FILLER_72_3428 ();
 sg13g2_fill_2 FILLER_72_3432 ();
 sg13g2_fill_2 FILLER_72_3438 ();
 sg13g2_decap_8 FILLER_72_3444 ();
 sg13g2_decap_4 FILLER_72_3451 ();
 sg13g2_fill_2 FILLER_72_3508 ();
 sg13g2_decap_8 FILLER_72_3519 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_fill_1 FILLER_73_49 ();
 sg13g2_fill_2 FILLER_73_87 ();
 sg13g2_fill_2 FILLER_73_131 ();
 sg13g2_fill_2 FILLER_73_183 ();
 sg13g2_fill_2 FILLER_73_205 ();
 sg13g2_fill_2 FILLER_73_262 ();
 sg13g2_fill_2 FILLER_73_277 ();
 sg13g2_decap_8 FILLER_73_295 ();
 sg13g2_decap_4 FILLER_73_302 ();
 sg13g2_decap_4 FILLER_73_326 ();
 sg13g2_fill_2 FILLER_73_335 ();
 sg13g2_fill_1 FILLER_73_337 ();
 sg13g2_decap_8 FILLER_73_352 ();
 sg13g2_decap_8 FILLER_73_359 ();
 sg13g2_fill_2 FILLER_73_366 ();
 sg13g2_fill_2 FILLER_73_389 ();
 sg13g2_decap_8 FILLER_73_408 ();
 sg13g2_fill_1 FILLER_73_415 ();
 sg13g2_fill_2 FILLER_73_424 ();
 sg13g2_fill_1 FILLER_73_426 ();
 sg13g2_decap_4 FILLER_73_440 ();
 sg13g2_fill_1 FILLER_73_462 ();
 sg13g2_fill_1 FILLER_73_470 ();
 sg13g2_fill_2 FILLER_73_482 ();
 sg13g2_decap_8 FILLER_73_510 ();
 sg13g2_decap_4 FILLER_73_517 ();
 sg13g2_decap_8 FILLER_73_544 ();
 sg13g2_fill_2 FILLER_73_560 ();
 sg13g2_fill_1 FILLER_73_562 ();
 sg13g2_decap_4 FILLER_73_577 ();
 sg13g2_decap_4 FILLER_73_586 ();
 sg13g2_fill_1 FILLER_73_590 ();
 sg13g2_fill_2 FILLER_73_623 ();
 sg13g2_fill_1 FILLER_73_625 ();
 sg13g2_decap_4 FILLER_73_645 ();
 sg13g2_fill_2 FILLER_73_649 ();
 sg13g2_decap_4 FILLER_73_655 ();
 sg13g2_fill_1 FILLER_73_678 ();
 sg13g2_decap_8 FILLER_73_692 ();
 sg13g2_decap_8 FILLER_73_699 ();
 sg13g2_decap_8 FILLER_73_727 ();
 sg13g2_decap_4 FILLER_73_734 ();
 sg13g2_fill_1 FILLER_73_738 ();
 sg13g2_decap_8 FILLER_73_747 ();
 sg13g2_decap_8 FILLER_73_754 ();
 sg13g2_decap_4 FILLER_73_761 ();
 sg13g2_fill_2 FILLER_73_776 ();
 sg13g2_decap_8 FILLER_73_802 ();
 sg13g2_decap_8 FILLER_73_834 ();
 sg13g2_fill_2 FILLER_73_856 ();
 sg13g2_fill_1 FILLER_73_858 ();
 sg13g2_decap_8 FILLER_73_871 ();
 sg13g2_decap_4 FILLER_73_878 ();
 sg13g2_fill_1 FILLER_73_890 ();
 sg13g2_fill_1 FILLER_73_905 ();
 sg13g2_decap_4 FILLER_73_911 ();
 sg13g2_fill_1 FILLER_73_933 ();
 sg13g2_fill_2 FILLER_73_942 ();
 sg13g2_decap_4 FILLER_73_947 ();
 sg13g2_fill_2 FILLER_73_966 ();
 sg13g2_fill_2 FILLER_73_982 ();
 sg13g2_decap_8 FILLER_73_1000 ();
 sg13g2_decap_4 FILLER_73_1007 ();
 sg13g2_fill_2 FILLER_73_1011 ();
 sg13g2_decap_8 FILLER_73_1026 ();
 sg13g2_decap_4 FILLER_73_1050 ();
 sg13g2_fill_1 FILLER_73_1054 ();
 sg13g2_decap_4 FILLER_73_1059 ();
 sg13g2_fill_2 FILLER_73_1063 ();
 sg13g2_fill_1 FILLER_73_1070 ();
 sg13g2_fill_2 FILLER_73_1090 ();
 sg13g2_fill_1 FILLER_73_1092 ();
 sg13g2_decap_4 FILLER_73_1114 ();
 sg13g2_fill_1 FILLER_73_1118 ();
 sg13g2_decap_4 FILLER_73_1147 ();
 sg13g2_fill_1 FILLER_73_1151 ();
 sg13g2_decap_8 FILLER_73_1164 ();
 sg13g2_fill_1 FILLER_73_1171 ();
 sg13g2_fill_1 FILLER_73_1210 ();
 sg13g2_decap_4 FILLER_73_1215 ();
 sg13g2_fill_2 FILLER_73_1224 ();
 sg13g2_fill_1 FILLER_73_1226 ();
 sg13g2_decap_8 FILLER_73_1232 ();
 sg13g2_fill_2 FILLER_73_1239 ();
 sg13g2_decap_8 FILLER_73_1251 ();
 sg13g2_fill_2 FILLER_73_1265 ();
 sg13g2_decap_4 FILLER_73_1284 ();
 sg13g2_fill_2 FILLER_73_1288 ();
 sg13g2_fill_1 FILLER_73_1298 ();
 sg13g2_fill_2 FILLER_73_1305 ();
 sg13g2_fill_2 FILLER_73_1317 ();
 sg13g2_decap_4 FILLER_73_1327 ();
 sg13g2_fill_2 FILLER_73_1347 ();
 sg13g2_fill_2 FILLER_73_1367 ();
 sg13g2_fill_1 FILLER_73_1369 ();
 sg13g2_fill_2 FILLER_73_1383 ();
 sg13g2_fill_1 FILLER_73_1397 ();
 sg13g2_decap_4 FILLER_73_1406 ();
 sg13g2_fill_1 FILLER_73_1410 ();
 sg13g2_fill_2 FILLER_73_1421 ();
 sg13g2_fill_2 FILLER_73_1429 ();
 sg13g2_fill_2 FILLER_73_1443 ();
 sg13g2_decap_8 FILLER_73_1461 ();
 sg13g2_decap_4 FILLER_73_1501 ();
 sg13g2_fill_1 FILLER_73_1505 ();
 sg13g2_fill_2 FILLER_73_1515 ();
 sg13g2_fill_1 FILLER_73_1525 ();
 sg13g2_fill_2 FILLER_73_1571 ();
 sg13g2_fill_1 FILLER_73_1573 ();
 sg13g2_fill_1 FILLER_73_1600 ();
 sg13g2_decap_8 FILLER_73_1605 ();
 sg13g2_fill_2 FILLER_73_1617 ();
 sg13g2_fill_1 FILLER_73_1619 ();
 sg13g2_fill_2 FILLER_73_1633 ();
 sg13g2_fill_1 FILLER_73_1635 ();
 sg13g2_fill_2 FILLER_73_1645 ();
 sg13g2_fill_1 FILLER_73_1647 ();
 sg13g2_decap_8 FILLER_73_1656 ();
 sg13g2_fill_1 FILLER_73_1663 ();
 sg13g2_fill_1 FILLER_73_1668 ();
 sg13g2_decap_8 FILLER_73_1682 ();
 sg13g2_fill_1 FILLER_73_1695 ();
 sg13g2_decap_8 FILLER_73_1700 ();
 sg13g2_decap_8 FILLER_73_1707 ();
 sg13g2_fill_2 FILLER_73_1714 ();
 sg13g2_fill_1 FILLER_73_1716 ();
 sg13g2_decap_8 FILLER_73_1721 ();
 sg13g2_decap_4 FILLER_73_1728 ();
 sg13g2_fill_2 FILLER_73_1732 ();
 sg13g2_decap_8 FILLER_73_1747 ();
 sg13g2_decap_4 FILLER_73_1754 ();
 sg13g2_fill_1 FILLER_73_1758 ();
 sg13g2_decap_8 FILLER_73_1770 ();
 sg13g2_decap_4 FILLER_73_1777 ();
 sg13g2_fill_2 FILLER_73_1781 ();
 sg13g2_fill_2 FILLER_73_1824 ();
 sg13g2_decap_4 FILLER_73_1898 ();
 sg13g2_fill_1 FILLER_73_1902 ();
 sg13g2_fill_2 FILLER_73_1912 ();
 sg13g2_fill_1 FILLER_73_1919 ();
 sg13g2_decap_8 FILLER_73_1924 ();
 sg13g2_decap_4 FILLER_73_1931 ();
 sg13g2_fill_1 FILLER_73_1935 ();
 sg13g2_decap_8 FILLER_73_1951 ();
 sg13g2_decap_8 FILLER_73_1958 ();
 sg13g2_decap_4 FILLER_73_1965 ();
 sg13g2_fill_1 FILLER_73_1969 ();
 sg13g2_fill_1 FILLER_73_1974 ();
 sg13g2_decap_4 FILLER_73_1985 ();
 sg13g2_fill_1 FILLER_73_1989 ();
 sg13g2_fill_1 FILLER_73_2018 ();
 sg13g2_fill_2 FILLER_73_2062 ();
 sg13g2_fill_2 FILLER_73_2072 ();
 sg13g2_decap_8 FILLER_73_2085 ();
 sg13g2_decap_8 FILLER_73_2092 ();
 sg13g2_fill_1 FILLER_73_2104 ();
 sg13g2_fill_1 FILLER_73_2110 ();
 sg13g2_decap_8 FILLER_73_2119 ();
 sg13g2_fill_2 FILLER_73_2126 ();
 sg13g2_fill_1 FILLER_73_2128 ();
 sg13g2_fill_1 FILLER_73_2155 ();
 sg13g2_fill_2 FILLER_73_2160 ();
 sg13g2_fill_1 FILLER_73_2162 ();
 sg13g2_fill_1 FILLER_73_2167 ();
 sg13g2_decap_8 FILLER_73_2172 ();
 sg13g2_fill_1 FILLER_73_2179 ();
 sg13g2_decap_8 FILLER_73_2210 ();
 sg13g2_decap_8 FILLER_73_2217 ();
 sg13g2_decap_8 FILLER_73_2224 ();
 sg13g2_decap_4 FILLER_73_2231 ();
 sg13g2_fill_2 FILLER_73_2235 ();
 sg13g2_decap_4 FILLER_73_2244 ();
 sg13g2_fill_2 FILLER_73_2352 ();
 sg13g2_fill_1 FILLER_73_2364 ();
 sg13g2_fill_1 FILLER_73_2391 ();
 sg13g2_decap_4 FILLER_73_2396 ();
 sg13g2_fill_2 FILLER_73_2405 ();
 sg13g2_fill_1 FILLER_73_2422 ();
 sg13g2_fill_1 FILLER_73_2431 ();
 sg13g2_fill_1 FILLER_73_2443 ();
 sg13g2_fill_1 FILLER_73_2449 ();
 sg13g2_fill_2 FILLER_73_2491 ();
 sg13g2_fill_1 FILLER_73_2493 ();
 sg13g2_decap_4 FILLER_73_2548 ();
 sg13g2_decap_4 FILLER_73_2578 ();
 sg13g2_fill_2 FILLER_73_2582 ();
 sg13g2_fill_1 FILLER_73_2588 ();
 sg13g2_decap_4 FILLER_73_2599 ();
 sg13g2_fill_2 FILLER_73_2603 ();
 sg13g2_decap_8 FILLER_73_2619 ();
 sg13g2_fill_1 FILLER_73_2626 ();
 sg13g2_fill_2 FILLER_73_2632 ();
 sg13g2_fill_1 FILLER_73_2652 ();
 sg13g2_decap_8 FILLER_73_2657 ();
 sg13g2_decap_8 FILLER_73_2664 ();
 sg13g2_fill_2 FILLER_73_2671 ();
 sg13g2_fill_1 FILLER_73_2673 ();
 sg13g2_fill_2 FILLER_73_2679 ();
 sg13g2_fill_2 FILLER_73_2685 ();
 sg13g2_fill_2 FILLER_73_2698 ();
 sg13g2_fill_1 FILLER_73_2700 ();
 sg13g2_decap_8 FILLER_73_2705 ();
 sg13g2_decap_8 FILLER_73_2712 ();
 sg13g2_fill_2 FILLER_73_2719 ();
 sg13g2_fill_1 FILLER_73_2721 ();
 sg13g2_decap_4 FILLER_73_2732 ();
 sg13g2_decap_4 FILLER_73_2749 ();
 sg13g2_fill_2 FILLER_73_2753 ();
 sg13g2_decap_8 FILLER_73_2778 ();
 sg13g2_fill_2 FILLER_73_2785 ();
 sg13g2_fill_1 FILLER_73_2787 ();
 sg13g2_fill_2 FILLER_73_2812 ();
 sg13g2_decap_8 FILLER_73_2820 ();
 sg13g2_decap_4 FILLER_73_2827 ();
 sg13g2_fill_1 FILLER_73_2831 ();
 sg13g2_fill_1 FILLER_73_2863 ();
 sg13g2_fill_1 FILLER_73_2873 ();
 sg13g2_fill_2 FILLER_73_2883 ();
 sg13g2_fill_2 FILLER_73_2898 ();
 sg13g2_fill_1 FILLER_73_2900 ();
 sg13g2_fill_1 FILLER_73_2909 ();
 sg13g2_fill_2 FILLER_73_2928 ();
 sg13g2_fill_1 FILLER_73_2930 ();
 sg13g2_fill_2 FILLER_73_2945 ();
 sg13g2_fill_2 FILLER_73_2951 ();
 sg13g2_fill_1 FILLER_73_2953 ();
 sg13g2_fill_1 FILLER_73_2967 ();
 sg13g2_decap_4 FILLER_73_2972 ();
 sg13g2_fill_1 FILLER_73_2976 ();
 sg13g2_fill_2 FILLER_73_2991 ();
 sg13g2_fill_2 FILLER_73_2999 ();
 sg13g2_fill_1 FILLER_73_3057 ();
 sg13g2_fill_2 FILLER_73_3121 ();
 sg13g2_fill_1 FILLER_73_3123 ();
 sg13g2_decap_4 FILLER_73_3128 ();
 sg13g2_fill_2 FILLER_73_3141 ();
 sg13g2_fill_1 FILLER_73_3143 ();
 sg13g2_decap_4 FILLER_73_3158 ();
 sg13g2_fill_2 FILLER_73_3162 ();
 sg13g2_decap_8 FILLER_73_3177 ();
 sg13g2_decap_4 FILLER_73_3197 ();
 sg13g2_fill_2 FILLER_73_3201 ();
 sg13g2_fill_2 FILLER_73_3208 ();
 sg13g2_fill_2 FILLER_73_3223 ();
 sg13g2_fill_1 FILLER_73_3225 ();
 sg13g2_fill_1 FILLER_73_3253 ();
 sg13g2_decap_8 FILLER_73_3270 ();
 sg13g2_decap_8 FILLER_73_3303 ();
 sg13g2_fill_1 FILLER_73_3364 ();
 sg13g2_fill_1 FILLER_73_3382 ();
 sg13g2_fill_1 FILLER_73_3411 ();
 sg13g2_fill_2 FILLER_73_3442 ();
 sg13g2_fill_2 FILLER_73_3466 ();
 sg13g2_decap_8 FILLER_73_3472 ();
 sg13g2_decap_8 FILLER_73_3479 ();
 sg13g2_decap_4 FILLER_73_3486 ();
 sg13g2_fill_1 FILLER_73_3490 ();
 sg13g2_fill_1 FILLER_73_3504 ();
 sg13g2_fill_2 FILLER_73_3525 ();
 sg13g2_fill_1 FILLER_73_3527 ();
 sg13g2_fill_2 FILLER_73_3554 ();
 sg13g2_fill_1 FILLER_73_3556 ();
 sg13g2_decap_8 FILLER_73_3565 ();
 sg13g2_decap_8 FILLER_73_3572 ();
 sg13g2_fill_1 FILLER_73_3579 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_fill_2 FILLER_74_42 ();
 sg13g2_fill_1 FILLER_74_128 ();
 sg13g2_fill_1 FILLER_74_173 ();
 sg13g2_fill_1 FILLER_74_239 ();
 sg13g2_fill_2 FILLER_74_290 ();
 sg13g2_decap_4 FILLER_74_300 ();
 sg13g2_decap_4 FILLER_74_320 ();
 sg13g2_decap_4 FILLER_74_356 ();
 sg13g2_fill_1 FILLER_74_360 ();
 sg13g2_fill_2 FILLER_74_383 ();
 sg13g2_fill_1 FILLER_74_385 ();
 sg13g2_fill_2 FILLER_74_412 ();
 sg13g2_fill_2 FILLER_74_430 ();
 sg13g2_fill_1 FILLER_74_472 ();
 sg13g2_decap_4 FILLER_74_487 ();
 sg13g2_decap_8 FILLER_74_504 ();
 sg13g2_decap_4 FILLER_74_511 ();
 sg13g2_fill_1 FILLER_74_515 ();
 sg13g2_decap_4 FILLER_74_525 ();
 sg13g2_fill_1 FILLER_74_537 ();
 sg13g2_fill_1 FILLER_74_551 ();
 sg13g2_decap_8 FILLER_74_593 ();
 sg13g2_decap_4 FILLER_74_600 ();
 sg13g2_fill_2 FILLER_74_608 ();
 sg13g2_fill_1 FILLER_74_610 ();
 sg13g2_decap_4 FILLER_74_621 ();
 sg13g2_fill_1 FILLER_74_629 ();
 sg13g2_fill_2 FILLER_74_657 ();
 sg13g2_fill_1 FILLER_74_659 ();
 sg13g2_decap_4 FILLER_74_669 ();
 sg13g2_fill_1 FILLER_74_673 ();
 sg13g2_fill_2 FILLER_74_687 ();
 sg13g2_fill_2 FILLER_74_693 ();
 sg13g2_fill_1 FILLER_74_695 ();
 sg13g2_decap_4 FILLER_74_706 ();
 sg13g2_fill_1 FILLER_74_710 ();
 sg13g2_fill_2 FILLER_74_717 ();
 sg13g2_decap_8 FILLER_74_723 ();
 sg13g2_decap_4 FILLER_74_730 ();
 sg13g2_fill_1 FILLER_74_734 ();
 sg13g2_decap_4 FILLER_74_739 ();
 sg13g2_fill_1 FILLER_74_743 ();
 sg13g2_decap_8 FILLER_74_763 ();
 sg13g2_decap_8 FILLER_74_774 ();
 sg13g2_decap_4 FILLER_74_781 ();
 sg13g2_decap_8 FILLER_74_804 ();
 sg13g2_fill_2 FILLER_74_811 ();
 sg13g2_fill_1 FILLER_74_813 ();
 sg13g2_fill_1 FILLER_74_832 ();
 sg13g2_fill_2 FILLER_74_841 ();
 sg13g2_fill_2 FILLER_74_856 ();
 sg13g2_decap_4 FILLER_74_877 ();
 sg13g2_decap_8 FILLER_74_901 ();
 sg13g2_fill_2 FILLER_74_918 ();
 sg13g2_fill_1 FILLER_74_920 ();
 sg13g2_decap_4 FILLER_74_949 ();
 sg13g2_fill_2 FILLER_74_953 ();
 sg13g2_decap_4 FILLER_74_963 ();
 sg13g2_fill_1 FILLER_74_967 ();
 sg13g2_fill_1 FILLER_74_978 ();
 sg13g2_decap_8 FILLER_74_994 ();
 sg13g2_decap_4 FILLER_74_1064 ();
 sg13g2_fill_1 FILLER_74_1068 ();
 sg13g2_fill_1 FILLER_74_1073 ();
 sg13g2_fill_2 FILLER_74_1087 ();
 sg13g2_fill_1 FILLER_74_1089 ();
 sg13g2_fill_1 FILLER_74_1131 ();
 sg13g2_decap_8 FILLER_74_1137 ();
 sg13g2_fill_2 FILLER_74_1144 ();
 sg13g2_decap_8 FILLER_74_1182 ();
 sg13g2_fill_2 FILLER_74_1189 ();
 sg13g2_fill_1 FILLER_74_1191 ();
 sg13g2_decap_4 FILLER_74_1226 ();
 sg13g2_fill_1 FILLER_74_1230 ();
 sg13g2_fill_2 FILLER_74_1239 ();
 sg13g2_fill_1 FILLER_74_1241 ();
 sg13g2_fill_2 FILLER_74_1277 ();
 sg13g2_fill_1 FILLER_74_1279 ();
 sg13g2_decap_8 FILLER_74_1307 ();
 sg13g2_fill_1 FILLER_74_1314 ();
 sg13g2_decap_8 FILLER_74_1327 ();
 sg13g2_fill_1 FILLER_74_1334 ();
 sg13g2_decap_4 FILLER_74_1355 ();
 sg13g2_fill_2 FILLER_74_1359 ();
 sg13g2_decap_8 FILLER_74_1365 ();
 sg13g2_fill_2 FILLER_74_1385 ();
 sg13g2_fill_2 FILLER_74_1392 ();
 sg13g2_fill_1 FILLER_74_1394 ();
 sg13g2_fill_2 FILLER_74_1400 ();
 sg13g2_fill_1 FILLER_74_1402 ();
 sg13g2_fill_2 FILLER_74_1411 ();
 sg13g2_fill_2 FILLER_74_1445 ();
 sg13g2_fill_2 FILLER_74_1450 ();
 sg13g2_fill_1 FILLER_74_1452 ();
 sg13g2_decap_8 FILLER_74_1465 ();
 sg13g2_decap_4 FILLER_74_1472 ();
 sg13g2_fill_1 FILLER_74_1476 ();
 sg13g2_decap_8 FILLER_74_1482 ();
 sg13g2_fill_1 FILLER_74_1494 ();
 sg13g2_fill_2 FILLER_74_1499 ();
 sg13g2_fill_1 FILLER_74_1510 ();
 sg13g2_decap_8 FILLER_74_1539 ();
 sg13g2_decap_4 FILLER_74_1554 ();
 sg13g2_fill_1 FILLER_74_1607 ();
 sg13g2_fill_1 FILLER_74_1629 ();
 sg13g2_decap_4 FILLER_74_1660 ();
 sg13g2_fill_1 FILLER_74_1679 ();
 sg13g2_fill_1 FILLER_74_1691 ();
 sg13g2_fill_2 FILLER_74_1709 ();
 sg13g2_fill_1 FILLER_74_1711 ();
 sg13g2_decap_4 FILLER_74_1748 ();
 sg13g2_fill_1 FILLER_74_1752 ();
 sg13g2_decap_8 FILLER_74_1772 ();
 sg13g2_decap_4 FILLER_74_1779 ();
 sg13g2_decap_4 FILLER_74_1796 ();
 sg13g2_fill_1 FILLER_74_1805 ();
 sg13g2_fill_1 FILLER_74_1828 ();
 sg13g2_fill_2 FILLER_74_1843 ();
 sg13g2_fill_1 FILLER_74_1845 ();
 sg13g2_decap_4 FILLER_74_1851 ();
 sg13g2_fill_2 FILLER_74_1874 ();
 sg13g2_decap_4 FILLER_74_1888 ();
 sg13g2_fill_1 FILLER_74_1892 ();
 sg13g2_decap_4 FILLER_74_1896 ();
 sg13g2_fill_2 FILLER_74_1900 ();
 sg13g2_decap_8 FILLER_74_1907 ();
 sg13g2_fill_2 FILLER_74_1942 ();
 sg13g2_fill_1 FILLER_74_1944 ();
 sg13g2_fill_2 FILLER_74_1962 ();
 sg13g2_fill_1 FILLER_74_1981 ();
 sg13g2_fill_1 FILLER_74_1985 ();
 sg13g2_fill_2 FILLER_74_1990 ();
 sg13g2_fill_2 FILLER_74_2032 ();
 sg13g2_fill_1 FILLER_74_2042 ();
 sg13g2_fill_1 FILLER_74_2055 ();
 sg13g2_decap_8 FILLER_74_2080 ();
 sg13g2_decap_8 FILLER_74_2087 ();
 sg13g2_fill_1 FILLER_74_2094 ();
 sg13g2_fill_2 FILLER_74_2116 ();
 sg13g2_fill_1 FILLER_74_2118 ();
 sg13g2_fill_2 FILLER_74_2151 ();
 sg13g2_fill_1 FILLER_74_2153 ();
 sg13g2_decap_8 FILLER_74_2175 ();
 sg13g2_decap_8 FILLER_74_2182 ();
 sg13g2_decap_4 FILLER_74_2189 ();
 sg13g2_fill_1 FILLER_74_2193 ();
 sg13g2_fill_2 FILLER_74_2215 ();
 sg13g2_fill_1 FILLER_74_2217 ();
 sg13g2_decap_4 FILLER_74_2227 ();
 sg13g2_fill_2 FILLER_74_2231 ();
 sg13g2_fill_1 FILLER_74_2254 ();
 sg13g2_fill_1 FILLER_74_2276 ();
 sg13g2_fill_1 FILLER_74_2281 ();
 sg13g2_fill_2 FILLER_74_2287 ();
 sg13g2_fill_1 FILLER_74_2289 ();
 sg13g2_fill_2 FILLER_74_2311 ();
 sg13g2_decap_8 FILLER_74_2319 ();
 sg13g2_fill_2 FILLER_74_2326 ();
 sg13g2_fill_1 FILLER_74_2328 ();
 sg13g2_decap_8 FILLER_74_2356 ();
 sg13g2_fill_2 FILLER_74_2363 ();
 sg13g2_fill_1 FILLER_74_2391 ();
 sg13g2_fill_1 FILLER_74_2431 ();
 sg13g2_fill_1 FILLER_74_2476 ();
 sg13g2_decap_8 FILLER_74_2490 ();
 sg13g2_decap_4 FILLER_74_2505 ();
 sg13g2_fill_1 FILLER_74_2509 ();
 sg13g2_fill_1 FILLER_74_2519 ();
 sg13g2_fill_2 FILLER_74_2554 ();
 sg13g2_fill_1 FILLER_74_2556 ();
 sg13g2_decap_8 FILLER_74_2571 ();
 sg13g2_decap_8 FILLER_74_2578 ();
 sg13g2_decap_4 FILLER_74_2585 ();
 sg13g2_fill_1 FILLER_74_2589 ();
 sg13g2_decap_4 FILLER_74_2600 ();
 sg13g2_fill_2 FILLER_74_2604 ();
 sg13g2_fill_1 FILLER_74_2611 ();
 sg13g2_decap_8 FILLER_74_2627 ();
 sg13g2_decap_4 FILLER_74_2634 ();
 sg13g2_fill_1 FILLER_74_2638 ();
 sg13g2_decap_8 FILLER_74_2657 ();
 sg13g2_fill_2 FILLER_74_2677 ();
 sg13g2_decap_4 FILLER_74_2692 ();
 sg13g2_decap_8 FILLER_74_2724 ();
 sg13g2_fill_2 FILLER_74_2783 ();
 sg13g2_fill_1 FILLER_74_2785 ();
 sg13g2_fill_1 FILLER_74_2798 ();
 sg13g2_decap_4 FILLER_74_2817 ();
 sg13g2_fill_1 FILLER_74_2821 ();
 sg13g2_fill_2 FILLER_74_2840 ();
 sg13g2_decap_4 FILLER_74_2873 ();
 sg13g2_decap_8 FILLER_74_2889 ();
 sg13g2_fill_1 FILLER_74_2896 ();
 sg13g2_fill_2 FILLER_74_2905 ();
 sg13g2_fill_1 FILLER_74_2907 ();
 sg13g2_fill_2 FILLER_74_2924 ();
 sg13g2_fill_2 FILLER_74_2947 ();
 sg13g2_fill_2 FILLER_74_2969 ();
 sg13g2_fill_1 FILLER_74_2971 ();
 sg13g2_decap_8 FILLER_74_2988 ();
 sg13g2_decap_4 FILLER_74_2995 ();
 sg13g2_fill_2 FILLER_74_2999 ();
 sg13g2_fill_2 FILLER_74_3018 ();
 sg13g2_fill_1 FILLER_74_3033 ();
 sg13g2_fill_1 FILLER_74_3062 ();
 sg13g2_decap_4 FILLER_74_3081 ();
 sg13g2_decap_8 FILLER_74_3108 ();
 sg13g2_decap_4 FILLER_74_3115 ();
 sg13g2_fill_1 FILLER_74_3119 ();
 sg13g2_decap_4 FILLER_74_3160 ();
 sg13g2_fill_1 FILLER_74_3164 ();
 sg13g2_decap_8 FILLER_74_3173 ();
 sg13g2_fill_1 FILLER_74_3180 ();
 sg13g2_fill_1 FILLER_74_3202 ();
 sg13g2_decap_8 FILLER_74_3216 ();
 sg13g2_decap_4 FILLER_74_3223 ();
 sg13g2_fill_1 FILLER_74_3227 ();
 sg13g2_fill_2 FILLER_74_3256 ();
 sg13g2_fill_2 FILLER_74_3266 ();
 sg13g2_decap_4 FILLER_74_3281 ();
 sg13g2_fill_1 FILLER_74_3285 ();
 sg13g2_decap_4 FILLER_74_3314 ();
 sg13g2_fill_1 FILLER_74_3318 ();
 sg13g2_decap_4 FILLER_74_3366 ();
 sg13g2_fill_1 FILLER_74_3370 ();
 sg13g2_decap_4 FILLER_74_3392 ();
 sg13g2_fill_1 FILLER_74_3396 ();
 sg13g2_decap_4 FILLER_74_3410 ();
 sg13g2_decap_4 FILLER_74_3429 ();
 sg13g2_decap_4 FILLER_74_3449 ();
 sg13g2_fill_2 FILLER_74_3478 ();
 sg13g2_fill_1 FILLER_74_3480 ();
 sg13g2_decap_8 FILLER_74_3494 ();
 sg13g2_fill_1 FILLER_74_3501 ();
 sg13g2_fill_1 FILLER_74_3511 ();
 sg13g2_decap_8 FILLER_74_3517 ();
 sg13g2_decap_4 FILLER_74_3524 ();
 sg13g2_fill_2 FILLER_74_3528 ();
 sg13g2_decap_4 FILLER_74_3549 ();
 sg13g2_fill_2 FILLER_74_3577 ();
 sg13g2_fill_1 FILLER_74_3579 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_4 FILLER_75_28 ();
 sg13g2_fill_2 FILLER_75_32 ();
 sg13g2_fill_2 FILLER_75_78 ();
 sg13g2_fill_1 FILLER_75_89 ();
 sg13g2_fill_1 FILLER_75_162 ();
 sg13g2_fill_2 FILLER_75_210 ();
 sg13g2_fill_1 FILLER_75_212 ();
 sg13g2_fill_1 FILLER_75_221 ();
 sg13g2_fill_1 FILLER_75_257 ();
 sg13g2_decap_8 FILLER_75_271 ();
 sg13g2_decap_8 FILLER_75_278 ();
 sg13g2_decap_8 FILLER_75_299 ();
 sg13g2_decap_4 FILLER_75_306 ();
 sg13g2_fill_2 FILLER_75_310 ();
 sg13g2_fill_1 FILLER_75_322 ();
 sg13g2_fill_2 FILLER_75_327 ();
 sg13g2_fill_1 FILLER_75_329 ();
 sg13g2_fill_2 FILLER_75_335 ();
 sg13g2_fill_1 FILLER_75_342 ();
 sg13g2_fill_2 FILLER_75_348 ();
 sg13g2_decap_8 FILLER_75_356 ();
 sg13g2_fill_1 FILLER_75_363 ();
 sg13g2_fill_1 FILLER_75_372 ();
 sg13g2_fill_2 FILLER_75_382 ();
 sg13g2_fill_2 FILLER_75_407 ();
 sg13g2_fill_1 FILLER_75_409 ();
 sg13g2_decap_8 FILLER_75_432 ();
 sg13g2_fill_2 FILLER_75_439 ();
 sg13g2_fill_1 FILLER_75_441 ();
 sg13g2_decap_8 FILLER_75_468 ();
 sg13g2_decap_4 FILLER_75_475 ();
 sg13g2_fill_2 FILLER_75_479 ();
 sg13g2_fill_1 FILLER_75_491 ();
 sg13g2_fill_2 FILLER_75_497 ();
 sg13g2_fill_2 FILLER_75_543 ();
 sg13g2_fill_1 FILLER_75_545 ();
 sg13g2_fill_2 FILLER_75_588 ();
 sg13g2_fill_2 FILLER_75_600 ();
 sg13g2_fill_2 FILLER_75_618 ();
 sg13g2_fill_1 FILLER_75_637 ();
 sg13g2_fill_2 FILLER_75_651 ();
 sg13g2_fill_1 FILLER_75_653 ();
 sg13g2_fill_2 FILLER_75_660 ();
 sg13g2_fill_1 FILLER_75_662 ();
 sg13g2_decap_8 FILLER_75_678 ();
 sg13g2_fill_2 FILLER_75_685 ();
 sg13g2_decap_4 FILLER_75_696 ();
 sg13g2_fill_1 FILLER_75_700 ();
 sg13g2_fill_2 FILLER_75_710 ();
 sg13g2_fill_1 FILLER_75_712 ();
 sg13g2_decap_4 FILLER_75_723 ();
 sg13g2_fill_2 FILLER_75_727 ();
 sg13g2_fill_2 FILLER_75_756 ();
 sg13g2_fill_2 FILLER_75_763 ();
 sg13g2_fill_1 FILLER_75_765 ();
 sg13g2_fill_2 FILLER_75_771 ();
 sg13g2_fill_1 FILLER_75_778 ();
 sg13g2_decap_4 FILLER_75_796 ();
 sg13g2_fill_2 FILLER_75_800 ();
 sg13g2_decap_4 FILLER_75_828 ();
 sg13g2_fill_2 FILLER_75_832 ();
 sg13g2_decap_8 FILLER_75_845 ();
 sg13g2_decap_8 FILLER_75_852 ();
 sg13g2_fill_2 FILLER_75_859 ();
 sg13g2_fill_1 FILLER_75_861 ();
 sg13g2_decap_8 FILLER_75_877 ();
 sg13g2_fill_1 FILLER_75_884 ();
 sg13g2_fill_2 FILLER_75_901 ();
 sg13g2_fill_1 FILLER_75_903 ();
 sg13g2_decap_4 FILLER_75_915 ();
 sg13g2_fill_1 FILLER_75_937 ();
 sg13g2_fill_1 FILLER_75_981 ();
 sg13g2_fill_2 FILLER_75_1004 ();
 sg13g2_fill_2 FILLER_75_1011 ();
 sg13g2_fill_1 FILLER_75_1017 ();
 sg13g2_decap_4 FILLER_75_1027 ();
 sg13g2_fill_2 FILLER_75_1031 ();
 sg13g2_fill_2 FILLER_75_1063 ();
 sg13g2_fill_2 FILLER_75_1070 ();
 sg13g2_fill_1 FILLER_75_1072 ();
 sg13g2_fill_2 FILLER_75_1096 ();
 sg13g2_fill_1 FILLER_75_1098 ();
 sg13g2_fill_2 FILLER_75_1106 ();
 sg13g2_fill_1 FILLER_75_1108 ();
 sg13g2_decap_4 FILLER_75_1119 ();
 sg13g2_fill_1 FILLER_75_1140 ();
 sg13g2_fill_1 FILLER_75_1154 ();
 sg13g2_decap_4 FILLER_75_1170 ();
 sg13g2_fill_2 FILLER_75_1174 ();
 sg13g2_fill_2 FILLER_75_1201 ();
 sg13g2_decap_8 FILLER_75_1207 ();
 sg13g2_decap_8 FILLER_75_1214 ();
 sg13g2_fill_2 FILLER_75_1221 ();
 sg13g2_fill_1 FILLER_75_1233 ();
 sg13g2_decap_4 FILLER_75_1242 ();
 sg13g2_decap_8 FILLER_75_1264 ();
 sg13g2_fill_1 FILLER_75_1271 ();
 sg13g2_fill_2 FILLER_75_1284 ();
 sg13g2_fill_1 FILLER_75_1286 ();
 sg13g2_fill_2 FILLER_75_1296 ();
 sg13g2_decap_8 FILLER_75_1315 ();
 sg13g2_decap_4 FILLER_75_1365 ();
 sg13g2_fill_1 FILLER_75_1369 ();
 sg13g2_fill_1 FILLER_75_1387 ();
 sg13g2_fill_2 FILLER_75_1396 ();
 sg13g2_fill_1 FILLER_75_1445 ();
 sg13g2_decap_8 FILLER_75_1450 ();
 sg13g2_fill_2 FILLER_75_1457 ();
 sg13g2_decap_8 FILLER_75_1464 ();
 sg13g2_decap_8 FILLER_75_1471 ();
 sg13g2_fill_1 FILLER_75_1492 ();
 sg13g2_decap_8 FILLER_75_1509 ();
 sg13g2_fill_2 FILLER_75_1516 ();
 sg13g2_fill_1 FILLER_75_1518 ();
 sg13g2_decap_4 FILLER_75_1528 ();
 sg13g2_fill_1 FILLER_75_1532 ();
 sg13g2_fill_2 FILLER_75_1546 ();
 sg13g2_fill_1 FILLER_75_1552 ();
 sg13g2_decap_4 FILLER_75_1565 ();
 sg13g2_decap_4 FILLER_75_1577 ();
 sg13g2_fill_1 FILLER_75_1581 ();
 sg13g2_decap_4 FILLER_75_1609 ();
 sg13g2_fill_2 FILLER_75_1613 ();
 sg13g2_decap_8 FILLER_75_1624 ();
 sg13g2_decap_4 FILLER_75_1631 ();
 sg13g2_fill_2 FILLER_75_1635 ();
 sg13g2_fill_2 FILLER_75_1646 ();
 sg13g2_decap_4 FILLER_75_1653 ();
 sg13g2_fill_2 FILLER_75_1657 ();
 sg13g2_fill_2 FILLER_75_1668 ();
 sg13g2_fill_1 FILLER_75_1670 ();
 sg13g2_fill_2 FILLER_75_1713 ();
 sg13g2_fill_1 FILLER_75_1725 ();
 sg13g2_fill_1 FILLER_75_1731 ();
 sg13g2_fill_2 FILLER_75_1742 ();
 sg13g2_fill_1 FILLER_75_1744 ();
 sg13g2_fill_2 FILLER_75_1754 ();
 sg13g2_fill_1 FILLER_75_1756 ();
 sg13g2_fill_2 FILLER_75_1794 ();
 sg13g2_decap_8 FILLER_75_1808 ();
 sg13g2_fill_2 FILLER_75_1815 ();
 sg13g2_decap_8 FILLER_75_1829 ();
 sg13g2_fill_2 FILLER_75_1836 ();
 sg13g2_decap_4 FILLER_75_1843 ();
 sg13g2_decap_4 FILLER_75_1875 ();
 sg13g2_decap_4 FILLER_75_1914 ();
 sg13g2_fill_1 FILLER_75_1918 ();
 sg13g2_fill_1 FILLER_75_1923 ();
 sg13g2_fill_2 FILLER_75_1932 ();
 sg13g2_fill_1 FILLER_75_1934 ();
 sg13g2_decap_4 FILLER_75_1948 ();
 sg13g2_fill_2 FILLER_75_2018 ();
 sg13g2_fill_1 FILLER_75_2020 ();
 sg13g2_fill_2 FILLER_75_2030 ();
 sg13g2_decap_4 FILLER_75_2050 ();
 sg13g2_fill_1 FILLER_75_2060 ();
 sg13g2_decap_4 FILLER_75_2073 ();
 sg13g2_fill_2 FILLER_75_2077 ();
 sg13g2_fill_1 FILLER_75_2083 ();
 sg13g2_decap_4 FILLER_75_2092 ();
 sg13g2_fill_2 FILLER_75_2096 ();
 sg13g2_fill_2 FILLER_75_2101 ();
 sg13g2_fill_2 FILLER_75_2116 ();
 sg13g2_decap_4 FILLER_75_2121 ();
 sg13g2_fill_1 FILLER_75_2137 ();
 sg13g2_fill_1 FILLER_75_2145 ();
 sg13g2_fill_2 FILLER_75_2151 ();
 sg13g2_fill_2 FILLER_75_2158 ();
 sg13g2_fill_1 FILLER_75_2160 ();
 sg13g2_decap_8 FILLER_75_2177 ();
 sg13g2_fill_2 FILLER_75_2184 ();
 sg13g2_fill_1 FILLER_75_2205 ();
 sg13g2_fill_2 FILLER_75_2217 ();
 sg13g2_decap_4 FILLER_75_2248 ();
 sg13g2_fill_2 FILLER_75_2252 ();
 sg13g2_decap_8 FILLER_75_2263 ();
 sg13g2_decap_4 FILLER_75_2270 ();
 sg13g2_fill_1 FILLER_75_2274 ();
 sg13g2_fill_2 FILLER_75_2303 ();
 sg13g2_fill_1 FILLER_75_2305 ();
 sg13g2_decap_4 FILLER_75_2338 ();
 sg13g2_decap_8 FILLER_75_2375 ();
 sg13g2_fill_1 FILLER_75_2382 ();
 sg13g2_decap_8 FILLER_75_2402 ();
 sg13g2_decap_4 FILLER_75_2409 ();
 sg13g2_fill_1 FILLER_75_2413 ();
 sg13g2_fill_1 FILLER_75_2426 ();
 sg13g2_fill_2 FILLER_75_2435 ();
 sg13g2_fill_1 FILLER_75_2437 ();
 sg13g2_fill_1 FILLER_75_2443 ();
 sg13g2_fill_2 FILLER_75_2461 ();
 sg13g2_fill_1 FILLER_75_2517 ();
 sg13g2_decap_4 FILLER_75_2526 ();
 sg13g2_fill_2 FILLER_75_2530 ();
 sg13g2_fill_2 FILLER_75_2540 ();
 sg13g2_fill_1 FILLER_75_2542 ();
 sg13g2_decap_4 FILLER_75_2547 ();
 sg13g2_fill_2 FILLER_75_2551 ();
 sg13g2_decap_8 FILLER_75_2568 ();
 sg13g2_fill_2 FILLER_75_2580 ();
 sg13g2_fill_2 FILLER_75_2611 ();
 sg13g2_decap_4 FILLER_75_2621 ();
 sg13g2_fill_1 FILLER_75_2625 ();
 sg13g2_fill_2 FILLER_75_2644 ();
 sg13g2_fill_1 FILLER_75_2659 ();
 sg13g2_fill_2 FILLER_75_2679 ();
 sg13g2_fill_2 FILLER_75_2687 ();
 sg13g2_decap_4 FILLER_75_2694 ();
 sg13g2_fill_1 FILLER_75_2702 ();
 sg13g2_fill_1 FILLER_75_2707 ();
 sg13g2_decap_8 FILLER_75_2723 ();
 sg13g2_fill_2 FILLER_75_2730 ();
 sg13g2_fill_2 FILLER_75_2754 ();
 sg13g2_fill_1 FILLER_75_2756 ();
 sg13g2_decap_4 FILLER_75_2787 ();
 sg13g2_fill_1 FILLER_75_2791 ();
 sg13g2_fill_1 FILLER_75_2804 ();
 sg13g2_decap_8 FILLER_75_2832 ();
 sg13g2_fill_2 FILLER_75_2839 ();
 sg13g2_fill_1 FILLER_75_2841 ();
 sg13g2_fill_2 FILLER_75_2854 ();
 sg13g2_decap_4 FILLER_75_2861 ();
 sg13g2_fill_1 FILLER_75_2865 ();
 sg13g2_decap_4 FILLER_75_2877 ();
 sg13g2_fill_2 FILLER_75_2881 ();
 sg13g2_fill_2 FILLER_75_2891 ();
 sg13g2_fill_1 FILLER_75_2893 ();
 sg13g2_fill_2 FILLER_75_2923 ();
 sg13g2_fill_1 FILLER_75_2925 ();
 sg13g2_fill_2 FILLER_75_2954 ();
 sg13g2_fill_2 FILLER_75_2965 ();
 sg13g2_fill_1 FILLER_75_2967 ();
 sg13g2_fill_2 FILLER_75_2990 ();
 sg13g2_fill_1 FILLER_75_2992 ();
 sg13g2_decap_8 FILLER_75_2998 ();
 sg13g2_fill_2 FILLER_75_3005 ();
 sg13g2_decap_4 FILLER_75_3033 ();
 sg13g2_fill_2 FILLER_75_3037 ();
 sg13g2_decap_8 FILLER_75_3043 ();
 sg13g2_fill_2 FILLER_75_3050 ();
 sg13g2_fill_1 FILLER_75_3052 ();
 sg13g2_decap_4 FILLER_75_3060 ();
 sg13g2_fill_1 FILLER_75_3098 ();
 sg13g2_decap_8 FILLER_75_3105 ();
 sg13g2_fill_2 FILLER_75_3112 ();
 sg13g2_fill_1 FILLER_75_3114 ();
 sg13g2_fill_2 FILLER_75_3127 ();
 sg13g2_fill_1 FILLER_75_3129 ();
 sg13g2_fill_1 FILLER_75_3133 ();
 sg13g2_fill_2 FILLER_75_3157 ();
 sg13g2_fill_1 FILLER_75_3159 ();
 sg13g2_decap_4 FILLER_75_3199 ();
 sg13g2_decap_8 FILLER_75_3219 ();
 sg13g2_fill_1 FILLER_75_3226 ();
 sg13g2_decap_8 FILLER_75_3233 ();
 sg13g2_fill_2 FILLER_75_3250 ();
 sg13g2_decap_4 FILLER_75_3266 ();
 sg13g2_fill_1 FILLER_75_3270 ();
 sg13g2_decap_4 FILLER_75_3276 ();
 sg13g2_fill_2 FILLER_75_3280 ();
 sg13g2_fill_2 FILLER_75_3304 ();
 sg13g2_fill_1 FILLER_75_3306 ();
 sg13g2_fill_2 FILLER_75_3316 ();
 sg13g2_fill_1 FILLER_75_3346 ();
 sg13g2_decap_4 FILLER_75_3361 ();
 sg13g2_decap_8 FILLER_75_3386 ();
 sg13g2_decap_8 FILLER_75_3393 ();
 sg13g2_fill_1 FILLER_75_3400 ();
 sg13g2_fill_2 FILLER_75_3418 ();
 sg13g2_fill_1 FILLER_75_3420 ();
 sg13g2_decap_8 FILLER_75_3431 ();
 sg13g2_fill_2 FILLER_75_3438 ();
 sg13g2_fill_1 FILLER_75_3440 ();
 sg13g2_decap_4 FILLER_75_3454 ();
 sg13g2_fill_1 FILLER_75_3473 ();
 sg13g2_fill_1 FILLER_75_3479 ();
 sg13g2_fill_2 FILLER_75_3485 ();
 sg13g2_decap_4 FILLER_75_3498 ();
 sg13g2_decap_8 FILLER_75_3538 ();
 sg13g2_fill_2 FILLER_75_3545 ();
 sg13g2_decap_8 FILLER_75_3571 ();
 sg13g2_fill_2 FILLER_75_3578 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_fill_2 FILLER_76_42 ();
 sg13g2_fill_1 FILLER_76_224 ();
 sg13g2_fill_2 FILLER_76_229 ();
 sg13g2_fill_1 FILLER_76_258 ();
 sg13g2_fill_2 FILLER_76_276 ();
 sg13g2_decap_4 FILLER_76_313 ();
 sg13g2_fill_2 FILLER_76_327 ();
 sg13g2_fill_1 FILLER_76_340 ();
 sg13g2_decap_4 FILLER_76_354 ();
 sg13g2_fill_1 FILLER_76_358 ();
 sg13g2_fill_2 FILLER_76_384 ();
 sg13g2_fill_1 FILLER_76_386 ();
 sg13g2_decap_8 FILLER_76_403 ();
 sg13g2_decap_8 FILLER_76_438 ();
 sg13g2_fill_2 FILLER_76_445 ();
 sg13g2_fill_1 FILLER_76_447 ();
 sg13g2_decap_8 FILLER_76_466 ();
 sg13g2_decap_4 FILLER_76_501 ();
 sg13g2_fill_2 FILLER_76_513 ();
 sg13g2_fill_1 FILLER_76_515 ();
 sg13g2_fill_1 FILLER_76_529 ();
 sg13g2_decap_8 FILLER_76_536 ();
 sg13g2_fill_1 FILLER_76_566 ();
 sg13g2_fill_2 FILLER_76_572 ();
 sg13g2_fill_1 FILLER_76_574 ();
 sg13g2_fill_2 FILLER_76_591 ();
 sg13g2_fill_1 FILLER_76_593 ();
 sg13g2_decap_4 FILLER_76_599 ();
 sg13g2_fill_1 FILLER_76_646 ();
 sg13g2_decap_8 FILLER_76_666 ();
 sg13g2_fill_1 FILLER_76_673 ();
 sg13g2_fill_2 FILLER_76_697 ();
 sg13g2_fill_2 FILLER_76_714 ();
 sg13g2_decap_8 FILLER_76_734 ();
 sg13g2_fill_1 FILLER_76_741 ();
 sg13g2_fill_1 FILLER_76_769 ();
 sg13g2_decap_4 FILLER_76_778 ();
 sg13g2_fill_1 FILLER_76_798 ();
 sg13g2_fill_2 FILLER_76_827 ();
 sg13g2_fill_2 FILLER_76_834 ();
 sg13g2_fill_1 FILLER_76_836 ();
 sg13g2_fill_2 FILLER_76_851 ();
 sg13g2_fill_1 FILLER_76_853 ();
 sg13g2_decap_4 FILLER_76_857 ();
 sg13g2_fill_1 FILLER_76_861 ();
 sg13g2_fill_1 FILLER_76_876 ();
 sg13g2_fill_1 FILLER_76_885 ();
 sg13g2_fill_2 FILLER_76_901 ();
 sg13g2_fill_1 FILLER_76_903 ();
 sg13g2_decap_8 FILLER_76_913 ();
 sg13g2_fill_2 FILLER_76_920 ();
 sg13g2_fill_1 FILLER_76_922 ();
 sg13g2_fill_2 FILLER_76_941 ();
 sg13g2_fill_1 FILLER_76_943 ();
 sg13g2_decap_8 FILLER_76_948 ();
 sg13g2_fill_2 FILLER_76_955 ();
 sg13g2_fill_1 FILLER_76_957 ();
 sg13g2_decap_8 FILLER_76_966 ();
 sg13g2_decap_8 FILLER_76_978 ();
 sg13g2_fill_1 FILLER_76_985 ();
 sg13g2_fill_1 FILLER_76_993 ();
 sg13g2_fill_2 FILLER_76_1002 ();
 sg13g2_fill_1 FILLER_76_1004 ();
 sg13g2_decap_8 FILLER_76_1022 ();
 sg13g2_decap_4 FILLER_76_1029 ();
 sg13g2_fill_2 FILLER_76_1038 ();
 sg13g2_fill_1 FILLER_76_1045 ();
 sg13g2_fill_1 FILLER_76_1058 ();
 sg13g2_decap_8 FILLER_76_1064 ();
 sg13g2_decap_8 FILLER_76_1071 ();
 sg13g2_decap_4 FILLER_76_1078 ();
 sg13g2_decap_8 FILLER_76_1090 ();
 sg13g2_fill_2 FILLER_76_1097 ();
 sg13g2_fill_2 FILLER_76_1104 ();
 sg13g2_fill_1 FILLER_76_1166 ();
 sg13g2_fill_2 FILLER_76_1178 ();
 sg13g2_fill_1 FILLER_76_1180 ();
 sg13g2_fill_2 FILLER_76_1202 ();
 sg13g2_fill_1 FILLER_76_1204 ();
 sg13g2_fill_2 FILLER_76_1213 ();
 sg13g2_decap_8 FILLER_76_1238 ();
 sg13g2_decap_4 FILLER_76_1245 ();
 sg13g2_decap_8 FILLER_76_1287 ();
 sg13g2_decap_4 FILLER_76_1294 ();
 sg13g2_fill_1 FILLER_76_1309 ();
 sg13g2_fill_2 FILLER_76_1323 ();
 sg13g2_fill_1 FILLER_76_1349 ();
 sg13g2_fill_2 FILLER_76_1354 ();
 sg13g2_decap_4 FILLER_76_1385 ();
 sg13g2_fill_1 FILLER_76_1401 ();
 sg13g2_decap_8 FILLER_76_1412 ();
 sg13g2_decap_4 FILLER_76_1419 ();
 sg13g2_fill_1 FILLER_76_1423 ();
 sg13g2_decap_4 FILLER_76_1435 ();
 sg13g2_fill_1 FILLER_76_1439 ();
 sg13g2_fill_2 FILLER_76_1457 ();
 sg13g2_fill_2 FILLER_76_1463 ();
 sg13g2_decap_4 FILLER_76_1473 ();
 sg13g2_decap_4 FILLER_76_1491 ();
 sg13g2_fill_1 FILLER_76_1495 ();
 sg13g2_decap_4 FILLER_76_1565 ();
 sg13g2_fill_1 FILLER_76_1573 ();
 sg13g2_fill_2 FILLER_76_1579 ();
 sg13g2_fill_2 FILLER_76_1585 ();
 sg13g2_fill_1 FILLER_76_1587 ();
 sg13g2_fill_1 FILLER_76_1607 ();
 sg13g2_decap_8 FILLER_76_1636 ();
 sg13g2_decap_4 FILLER_76_1647 ();
 sg13g2_fill_1 FILLER_76_1651 ();
 sg13g2_fill_2 FILLER_76_1674 ();
 sg13g2_fill_1 FILLER_76_1676 ();
 sg13g2_decap_4 FILLER_76_1681 ();
 sg13g2_fill_2 FILLER_76_1685 ();
 sg13g2_fill_2 FILLER_76_1693 ();
 sg13g2_fill_2 FILLER_76_1705 ();
 sg13g2_fill_2 FILLER_76_1720 ();
 sg13g2_fill_1 FILLER_76_1726 ();
 sg13g2_decap_8 FILLER_76_1744 ();
 sg13g2_decap_8 FILLER_76_1751 ();
 sg13g2_fill_1 FILLER_76_1758 ();
 sg13g2_fill_2 FILLER_76_1777 ();
 sg13g2_decap_8 FILLER_76_1803 ();
 sg13g2_fill_2 FILLER_76_1810 ();
 sg13g2_fill_2 FILLER_76_1838 ();
 sg13g2_decap_8 FILLER_76_1848 ();
 sg13g2_decap_4 FILLER_76_1878 ();
 sg13g2_fill_1 FILLER_76_1882 ();
 sg13g2_decap_4 FILLER_76_1893 ();
 sg13g2_fill_1 FILLER_76_1902 ();
 sg13g2_decap_4 FILLER_76_1907 ();
 sg13g2_fill_2 FILLER_76_1911 ();
 sg13g2_fill_1 FILLER_76_1937 ();
 sg13g2_fill_1 FILLER_76_1964 ();
 sg13g2_decap_8 FILLER_76_1976 ();
 sg13g2_fill_2 FILLER_76_1983 ();
 sg13g2_fill_1 FILLER_76_1985 ();
 sg13g2_fill_2 FILLER_76_1989 ();
 sg13g2_fill_1 FILLER_76_1991 ();
 sg13g2_fill_2 FILLER_76_2009 ();
 sg13g2_fill_1 FILLER_76_2011 ();
 sg13g2_fill_2 FILLER_76_2027 ();
 sg13g2_fill_1 FILLER_76_2029 ();
 sg13g2_fill_2 FILLER_76_2054 ();
 sg13g2_fill_1 FILLER_76_2056 ();
 sg13g2_fill_2 FILLER_76_2070 ();
 sg13g2_fill_1 FILLER_76_2072 ();
 sg13g2_fill_1 FILLER_76_2079 ();
 sg13g2_decap_4 FILLER_76_2088 ();
 sg13g2_fill_1 FILLER_76_2092 ();
 sg13g2_fill_2 FILLER_76_2131 ();
 sg13g2_fill_1 FILLER_76_2138 ();
 sg13g2_fill_2 FILLER_76_2151 ();
 sg13g2_fill_2 FILLER_76_2161 ();
 sg13g2_fill_1 FILLER_76_2171 ();
 sg13g2_fill_2 FILLER_76_2188 ();
 sg13g2_fill_1 FILLER_76_2190 ();
 sg13g2_fill_2 FILLER_76_2200 ();
 sg13g2_fill_1 FILLER_76_2202 ();
 sg13g2_fill_1 FILLER_76_2220 ();
 sg13g2_fill_1 FILLER_76_2229 ();
 sg13g2_fill_1 FILLER_76_2243 ();
 sg13g2_fill_2 FILLER_76_2264 ();
 sg13g2_fill_1 FILLER_76_2266 ();
 sg13g2_decap_8 FILLER_76_2272 ();
 sg13g2_fill_2 FILLER_76_2279 ();
 sg13g2_fill_1 FILLER_76_2281 ();
 sg13g2_fill_2 FILLER_76_2307 ();
 sg13g2_fill_2 FILLER_76_2325 ();
 sg13g2_fill_1 FILLER_76_2327 ();
 sg13g2_fill_2 FILLER_76_2343 ();
 sg13g2_fill_1 FILLER_76_2354 ();
 sg13g2_fill_2 FILLER_76_2381 ();
 sg13g2_fill_1 FILLER_76_2401 ();
 sg13g2_decap_8 FILLER_76_2414 ();
 sg13g2_fill_1 FILLER_76_2426 ();
 sg13g2_decap_8 FILLER_76_2452 ();
 sg13g2_fill_2 FILLER_76_2459 ();
 sg13g2_fill_1 FILLER_76_2461 ();
 sg13g2_fill_2 FILLER_76_2555 ();
 sg13g2_fill_1 FILLER_76_2557 ();
 sg13g2_decap_8 FILLER_76_2593 ();
 sg13g2_fill_2 FILLER_76_2600 ();
 sg13g2_fill_1 FILLER_76_2602 ();
 sg13g2_fill_1 FILLER_76_2612 ();
 sg13g2_fill_2 FILLER_76_2623 ();
 sg13g2_fill_1 FILLER_76_2625 ();
 sg13g2_decap_4 FILLER_76_2630 ();
 sg13g2_fill_1 FILLER_76_2634 ();
 sg13g2_fill_2 FILLER_76_2640 ();
 sg13g2_decap_8 FILLER_76_2674 ();
 sg13g2_fill_2 FILLER_76_2681 ();
 sg13g2_fill_1 FILLER_76_2683 ();
 sg13g2_fill_2 FILLER_76_2687 ();
 sg13g2_fill_2 FILLER_76_2697 ();
 sg13g2_decap_4 FILLER_76_2729 ();
 sg13g2_fill_1 FILLER_76_2733 ();
 sg13g2_fill_2 FILLER_76_2739 ();
 sg13g2_fill_1 FILLER_76_2746 ();
 sg13g2_decap_4 FILLER_76_2763 ();
 sg13g2_decap_8 FILLER_76_2785 ();
 sg13g2_fill_2 FILLER_76_2805 ();
 sg13g2_fill_1 FILLER_76_2807 ();
 sg13g2_fill_1 FILLER_76_2816 ();
 sg13g2_fill_2 FILLER_76_2852 ();
 sg13g2_decap_4 FILLER_76_2873 ();
 sg13g2_fill_1 FILLER_76_2877 ();
 sg13g2_decap_8 FILLER_76_2887 ();
 sg13g2_decap_4 FILLER_76_2894 ();
 sg13g2_fill_2 FILLER_76_2928 ();
 sg13g2_fill_1 FILLER_76_2930 ();
 sg13g2_fill_2 FILLER_76_2943 ();
 sg13g2_fill_1 FILLER_76_2945 ();
 sg13g2_decap_4 FILLER_76_2989 ();
 sg13g2_fill_1 FILLER_76_2993 ();
 sg13g2_decap_8 FILLER_76_3004 ();
 sg13g2_fill_1 FILLER_76_3020 ();
 sg13g2_fill_1 FILLER_76_3049 ();
 sg13g2_decap_4 FILLER_76_3090 ();
 sg13g2_decap_4 FILLER_76_3120 ();
 sg13g2_decap_4 FILLER_76_3137 ();
 sg13g2_decap_8 FILLER_76_3154 ();
 sg13g2_fill_1 FILLER_76_3161 ();
 sg13g2_decap_8 FILLER_76_3186 ();
 sg13g2_decap_4 FILLER_76_3193 ();
 sg13g2_fill_2 FILLER_76_3225 ();
 sg13g2_fill_1 FILLER_76_3227 ();
 sg13g2_fill_2 FILLER_76_3233 ();
 sg13g2_fill_1 FILLER_76_3235 ();
 sg13g2_fill_2 FILLER_76_3242 ();
 sg13g2_fill_2 FILLER_76_3273 ();
 sg13g2_decap_8 FILLER_76_3283 ();
 sg13g2_decap_8 FILLER_76_3303 ();
 sg13g2_decap_4 FILLER_76_3310 ();
 sg13g2_fill_2 FILLER_76_3314 ();
 sg13g2_fill_1 FILLER_76_3337 ();
 sg13g2_fill_2 FILLER_76_3355 ();
 sg13g2_fill_1 FILLER_76_3367 ();
 sg13g2_fill_2 FILLER_76_3375 ();
 sg13g2_decap_8 FILLER_76_3385 ();
 sg13g2_decap_4 FILLER_76_3392 ();
 sg13g2_fill_1 FILLER_76_3409 ();
 sg13g2_fill_2 FILLER_76_3415 ();
 sg13g2_fill_1 FILLER_76_3417 ();
 sg13g2_fill_2 FILLER_76_3426 ();
 sg13g2_decap_8 FILLER_76_3438 ();
 sg13g2_decap_4 FILLER_76_3445 ();
 sg13g2_fill_2 FILLER_76_3449 ();
 sg13g2_decap_4 FILLER_76_3472 ();
 sg13g2_fill_1 FILLER_76_3476 ();
 sg13g2_fill_2 FILLER_76_3516 ();
 sg13g2_fill_1 FILLER_76_3518 ();
 sg13g2_decap_4 FILLER_76_3524 ();
 sg13g2_fill_1 FILLER_76_3528 ();
 sg13g2_fill_1 FILLER_76_3546 ();
 sg13g2_decap_4 FILLER_76_3576 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_fill_2 FILLER_77_35 ();
 sg13g2_fill_1 FILLER_77_129 ();
 sg13g2_fill_2 FILLER_77_151 ();
 sg13g2_fill_1 FILLER_77_267 ();
 sg13g2_fill_1 FILLER_77_273 ();
 sg13g2_fill_2 FILLER_77_283 ();
 sg13g2_fill_1 FILLER_77_285 ();
 sg13g2_decap_8 FILLER_77_299 ();
 sg13g2_fill_1 FILLER_77_306 ();
 sg13g2_decap_8 FILLER_77_321 ();
 sg13g2_fill_1 FILLER_77_328 ();
 sg13g2_fill_2 FILLER_77_339 ();
 sg13g2_fill_1 FILLER_77_341 ();
 sg13g2_decap_4 FILLER_77_352 ();
 sg13g2_decap_4 FILLER_77_387 ();
 sg13g2_fill_2 FILLER_77_391 ();
 sg13g2_decap_8 FILLER_77_406 ();
 sg13g2_fill_2 FILLER_77_413 ();
 sg13g2_fill_1 FILLER_77_415 ();
 sg13g2_fill_1 FILLER_77_420 ();
 sg13g2_decap_4 FILLER_77_436 ();
 sg13g2_fill_2 FILLER_77_440 ();
 sg13g2_fill_2 FILLER_77_460 ();
 sg13g2_fill_1 FILLER_77_474 ();
 sg13g2_fill_2 FILLER_77_484 ();
 sg13g2_decap_4 FILLER_77_489 ();
 sg13g2_fill_2 FILLER_77_493 ();
 sg13g2_decap_8 FILLER_77_499 ();
 sg13g2_decap_4 FILLER_77_506 ();
 sg13g2_decap_4 FILLER_77_519 ();
 sg13g2_fill_2 FILLER_77_523 ();
 sg13g2_decap_4 FILLER_77_545 ();
 sg13g2_decap_8 FILLER_77_571 ();
 sg13g2_decap_4 FILLER_77_578 ();
 sg13g2_decap_4 FILLER_77_604 ();
 sg13g2_fill_2 FILLER_77_608 ();
 sg13g2_decap_8 FILLER_77_615 ();
 sg13g2_decap_4 FILLER_77_622 ();
 sg13g2_fill_2 FILLER_77_634 ();
 sg13g2_fill_1 FILLER_77_636 ();
 sg13g2_decap_8 FILLER_77_663 ();
 sg13g2_decap_8 FILLER_77_670 ();
 sg13g2_fill_1 FILLER_77_677 ();
 sg13g2_fill_2 FILLER_77_700 ();
 sg13g2_fill_1 FILLER_77_702 ();
 sg13g2_decap_8 FILLER_77_732 ();
 sg13g2_fill_2 FILLER_77_739 ();
 sg13g2_fill_1 FILLER_77_741 ();
 sg13g2_fill_2 FILLER_77_763 ();
 sg13g2_fill_1 FILLER_77_770 ();
 sg13g2_decap_8 FILLER_77_792 ();
 sg13g2_fill_2 FILLER_77_799 ();
 sg13g2_fill_2 FILLER_77_809 ();
 sg13g2_fill_1 FILLER_77_819 ();
 sg13g2_decap_4 FILLER_77_838 ();
 sg13g2_fill_2 FILLER_77_842 ();
 sg13g2_fill_1 FILLER_77_852 ();
 sg13g2_fill_1 FILLER_77_872 ();
 sg13g2_fill_2 FILLER_77_878 ();
 sg13g2_decap_8 FILLER_77_889 ();
 sg13g2_decap_8 FILLER_77_912 ();
 sg13g2_fill_1 FILLER_77_919 ();
 sg13g2_decap_4 FILLER_77_954 ();
 sg13g2_fill_1 FILLER_77_971 ();
 sg13g2_fill_1 FILLER_77_988 ();
 sg13g2_fill_2 FILLER_77_999 ();
 sg13g2_fill_1 FILLER_77_1009 ();
 sg13g2_fill_2 FILLER_77_1014 ();
 sg13g2_fill_1 FILLER_77_1016 ();
 sg13g2_fill_2 FILLER_77_1022 ();
 sg13g2_fill_1 FILLER_77_1024 ();
 sg13g2_fill_2 FILLER_77_1049 ();
 sg13g2_decap_4 FILLER_77_1067 ();
 sg13g2_fill_1 FILLER_77_1071 ();
 sg13g2_fill_2 FILLER_77_1093 ();
 sg13g2_fill_1 FILLER_77_1095 ();
 sg13g2_fill_1 FILLER_77_1108 ();
 sg13g2_decap_8 FILLER_77_1114 ();
 sg13g2_decap_4 FILLER_77_1121 ();
 sg13g2_fill_2 FILLER_77_1125 ();
 sg13g2_decap_8 FILLER_77_1132 ();
 sg13g2_decap_8 FILLER_77_1139 ();
 sg13g2_decap_8 FILLER_77_1146 ();
 sg13g2_fill_1 FILLER_77_1153 ();
 sg13g2_fill_2 FILLER_77_1172 ();
 sg13g2_decap_8 FILLER_77_1186 ();
 sg13g2_fill_2 FILLER_77_1211 ();
 sg13g2_decap_8 FILLER_77_1239 ();
 sg13g2_decap_4 FILLER_77_1246 ();
 sg13g2_fill_1 FILLER_77_1250 ();
 sg13g2_fill_2 FILLER_77_1264 ();
 sg13g2_fill_1 FILLER_77_1286 ();
 sg13g2_decap_8 FILLER_77_1316 ();
 sg13g2_decap_8 FILLER_77_1323 ();
 sg13g2_decap_8 FILLER_77_1348 ();
 sg13g2_decap_8 FILLER_77_1355 ();
 sg13g2_fill_2 FILLER_77_1366 ();
 sg13g2_decap_4 FILLER_77_1376 ();
 sg13g2_fill_2 FILLER_77_1385 ();
 sg13g2_decap_8 FILLER_77_1396 ();
 sg13g2_decap_8 FILLER_77_1403 ();
 sg13g2_fill_1 FILLER_77_1410 ();
 sg13g2_fill_1 FILLER_77_1415 ();
 sg13g2_fill_2 FILLER_77_1434 ();
 sg13g2_fill_1 FILLER_77_1436 ();
 sg13g2_fill_2 FILLER_77_1460 ();
 sg13g2_fill_1 FILLER_77_1462 ();
 sg13g2_fill_2 FILLER_77_1498 ();
 sg13g2_fill_2 FILLER_77_1505 ();
 sg13g2_fill_1 FILLER_77_1507 ();
 sg13g2_decap_8 FILLER_77_1513 ();
 sg13g2_fill_1 FILLER_77_1520 ();
 sg13g2_decap_8 FILLER_77_1536 ();
 sg13g2_fill_2 FILLER_77_1543 ();
 sg13g2_fill_1 FILLER_77_1545 ();
 sg13g2_fill_1 FILLER_77_1555 ();
 sg13g2_fill_1 FILLER_77_1561 ();
 sg13g2_fill_1 FILLER_77_1579 ();
 sg13g2_decap_4 FILLER_77_1612 ();
 sg13g2_fill_2 FILLER_77_1616 ();
 sg13g2_fill_2 FILLER_77_1624 ();
 sg13g2_fill_1 FILLER_77_1638 ();
 sg13g2_decap_8 FILLER_77_1648 ();
 sg13g2_fill_2 FILLER_77_1655 ();
 sg13g2_decap_8 FILLER_77_1669 ();
 sg13g2_fill_2 FILLER_77_1676 ();
 sg13g2_fill_1 FILLER_77_1696 ();
 sg13g2_decap_8 FILLER_77_1705 ();
 sg13g2_fill_2 FILLER_77_1712 ();
 sg13g2_fill_2 FILLER_77_1719 ();
 sg13g2_fill_1 FILLER_77_1726 ();
 sg13g2_fill_2 FILLER_77_1749 ();
 sg13g2_fill_1 FILLER_77_1751 ();
 sg13g2_decap_4 FILLER_77_1778 ();
 sg13g2_fill_1 FILLER_77_1782 ();
 sg13g2_decap_8 FILLER_77_1799 ();
 sg13g2_decap_8 FILLER_77_1806 ();
 sg13g2_decap_4 FILLER_77_1813 ();
 sg13g2_fill_1 FILLER_77_1835 ();
 sg13g2_decap_4 FILLER_77_1841 ();
 sg13g2_decap_4 FILLER_77_1849 ();
 sg13g2_fill_2 FILLER_77_1870 ();
 sg13g2_fill_1 FILLER_77_1872 ();
 sg13g2_decap_8 FILLER_77_1878 ();
 sg13g2_fill_2 FILLER_77_1896 ();
 sg13g2_decap_8 FILLER_77_1906 ();
 sg13g2_fill_1 FILLER_77_1913 ();
 sg13g2_decap_8 FILLER_77_1931 ();
 sg13g2_fill_2 FILLER_77_1938 ();
 sg13g2_fill_1 FILLER_77_1940 ();
 sg13g2_fill_1 FILLER_77_1961 ();
 sg13g2_fill_2 FILLER_77_1988 ();
 sg13g2_fill_1 FILLER_77_1990 ();
 sg13g2_decap_8 FILLER_77_2006 ();
 sg13g2_decap_8 FILLER_77_2052 ();
 sg13g2_fill_2 FILLER_77_2059 ();
 sg13g2_fill_1 FILLER_77_2061 ();
 sg13g2_decap_8 FILLER_77_2079 ();
 sg13g2_fill_1 FILLER_77_2086 ();
 sg13g2_decap_4 FILLER_77_2100 ();
 sg13g2_fill_2 FILLER_77_2104 ();
 sg13g2_decap_8 FILLER_77_2119 ();
 sg13g2_decap_4 FILLER_77_2126 ();
 sg13g2_fill_2 FILLER_77_2134 ();
 sg13g2_fill_1 FILLER_77_2136 ();
 sg13g2_fill_2 FILLER_77_2156 ();
 sg13g2_decap_8 FILLER_77_2167 ();
 sg13g2_decap_4 FILLER_77_2174 ();
 sg13g2_fill_1 FILLER_77_2178 ();
 sg13g2_fill_1 FILLER_77_2187 ();
 sg13g2_decap_8 FILLER_77_2206 ();
 sg13g2_fill_2 FILLER_77_2213 ();
 sg13g2_fill_2 FILLER_77_2248 ();
 sg13g2_decap_4 FILLER_77_2255 ();
 sg13g2_fill_1 FILLER_77_2269 ();
 sg13g2_fill_2 FILLER_77_2274 ();
 sg13g2_decap_8 FILLER_77_2282 ();
 sg13g2_fill_2 FILLER_77_2289 ();
 sg13g2_fill_1 FILLER_77_2291 ();
 sg13g2_decap_4 FILLER_77_2295 ();
 sg13g2_fill_2 FILLER_77_2299 ();
 sg13g2_fill_2 FILLER_77_2306 ();
 sg13g2_fill_1 FILLER_77_2308 ();
 sg13g2_fill_2 FILLER_77_2314 ();
 sg13g2_decap_8 FILLER_77_2329 ();
 sg13g2_fill_2 FILLER_77_2336 ();
 sg13g2_fill_1 FILLER_77_2338 ();
 sg13g2_decap_8 FILLER_77_2349 ();
 sg13g2_decap_4 FILLER_77_2356 ();
 sg13g2_fill_2 FILLER_77_2385 ();
 sg13g2_fill_1 FILLER_77_2387 ();
 sg13g2_fill_2 FILLER_77_2409 ();
 sg13g2_decap_8 FILLER_77_2423 ();
 sg13g2_fill_2 FILLER_77_2430 ();
 sg13g2_fill_1 FILLER_77_2432 ();
 sg13g2_decap_4 FILLER_77_2451 ();
 sg13g2_fill_1 FILLER_77_2455 ();
 sg13g2_fill_2 FILLER_77_2479 ();
 sg13g2_decap_8 FILLER_77_2489 ();
 sg13g2_decap_4 FILLER_77_2496 ();
 sg13g2_fill_2 FILLER_77_2513 ();
 sg13g2_fill_1 FILLER_77_2528 ();
 sg13g2_fill_2 FILLER_77_2542 ();
 sg13g2_fill_1 FILLER_77_2544 ();
 sg13g2_fill_1 FILLER_77_2563 ();
 sg13g2_decap_8 FILLER_77_2584 ();
 sg13g2_decap_4 FILLER_77_2591 ();
 sg13g2_fill_1 FILLER_77_2595 ();
 sg13g2_decap_4 FILLER_77_2634 ();
 sg13g2_fill_2 FILLER_77_2658 ();
 sg13g2_fill_1 FILLER_77_2660 ();
 sg13g2_decap_4 FILLER_77_2677 ();
 sg13g2_fill_1 FILLER_77_2681 ();
 sg13g2_fill_2 FILLER_77_2690 ();
 sg13g2_fill_1 FILLER_77_2714 ();
 sg13g2_decap_8 FILLER_77_2723 ();
 sg13g2_decap_4 FILLER_77_2730 ();
 sg13g2_fill_2 FILLER_77_2743 ();
 sg13g2_fill_1 FILLER_77_2745 ();
 sg13g2_decap_4 FILLER_77_2770 ();
 sg13g2_decap_8 FILLER_77_2779 ();
 sg13g2_decap_8 FILLER_77_2786 ();
 sg13g2_fill_2 FILLER_77_2819 ();
 sg13g2_fill_1 FILLER_77_2821 ();
 sg13g2_fill_2 FILLER_77_2830 ();
 sg13g2_decap_4 FILLER_77_2840 ();
 sg13g2_decap_4 FILLER_77_2861 ();
 sg13g2_fill_2 FILLER_77_2865 ();
 sg13g2_fill_1 FILLER_77_2872 ();
 sg13g2_decap_8 FILLER_77_2889 ();
 sg13g2_fill_2 FILLER_77_2906 ();
 sg13g2_fill_1 FILLER_77_2908 ();
 sg13g2_fill_2 FILLER_77_2930 ();
 sg13g2_fill_1 FILLER_77_2932 ();
 sg13g2_fill_2 FILLER_77_2968 ();
 sg13g2_fill_1 FILLER_77_2970 ();
 sg13g2_fill_1 FILLER_77_2998 ();
 sg13g2_decap_4 FILLER_77_3004 ();
 sg13g2_fill_2 FILLER_77_3008 ();
 sg13g2_decap_4 FILLER_77_3020 ();
 sg13g2_fill_1 FILLER_77_3065 ();
 sg13g2_fill_1 FILLER_77_3071 ();
 sg13g2_decap_4 FILLER_77_3088 ();
 sg13g2_fill_1 FILLER_77_3092 ();
 sg13g2_fill_2 FILLER_77_3103 ();
 sg13g2_fill_1 FILLER_77_3105 ();
 sg13g2_fill_2 FILLER_77_3111 ();
 sg13g2_fill_1 FILLER_77_3113 ();
 sg13g2_fill_1 FILLER_77_3140 ();
 sg13g2_fill_2 FILLER_77_3166 ();
 sg13g2_decap_4 FILLER_77_3185 ();
 sg13g2_decap_4 FILLER_77_3198 ();
 sg13g2_fill_2 FILLER_77_3202 ();
 sg13g2_decap_8 FILLER_77_3208 ();
 sg13g2_decap_8 FILLER_77_3232 ();
 sg13g2_fill_2 FILLER_77_3239 ();
 sg13g2_fill_2 FILLER_77_3246 ();
 sg13g2_fill_1 FILLER_77_3252 ();
 sg13g2_fill_2 FILLER_77_3262 ();
 sg13g2_fill_1 FILLER_77_3288 ();
 sg13g2_decap_4 FILLER_77_3309 ();
 sg13g2_decap_4 FILLER_77_3323 ();
 sg13g2_fill_2 FILLER_77_3327 ();
 sg13g2_fill_1 FILLER_77_3341 ();
 sg13g2_fill_2 FILLER_77_3360 ();
 sg13g2_decap_8 FILLER_77_3395 ();
 sg13g2_fill_2 FILLER_77_3425 ();
 sg13g2_decap_8 FILLER_77_3447 ();
 sg13g2_fill_2 FILLER_77_3454 ();
 sg13g2_fill_1 FILLER_77_3456 ();
 sg13g2_decap_8 FILLER_77_3470 ();
 sg13g2_fill_2 FILLER_77_3509 ();
 sg13g2_fill_1 FILLER_77_3511 ();
 sg13g2_fill_1 FILLER_77_3529 ();
 sg13g2_decap_8 FILLER_77_3543 ();
 sg13g2_fill_1 FILLER_77_3550 ();
 sg13g2_decap_4 FILLER_77_3576 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_4 FILLER_78_35 ();
 sg13g2_fill_1 FILLER_78_39 ();
 sg13g2_fill_2 FILLER_78_105 ();
 sg13g2_fill_2 FILLER_78_133 ();
 sg13g2_fill_2 FILLER_78_240 ();
 sg13g2_fill_1 FILLER_78_251 ();
 sg13g2_decap_4 FILLER_78_334 ();
 sg13g2_fill_1 FILLER_78_338 ();
 sg13g2_fill_1 FILLER_78_343 ();
 sg13g2_decap_8 FILLER_78_348 ();
 sg13g2_decap_4 FILLER_78_355 ();
 sg13g2_fill_2 FILLER_78_359 ();
 sg13g2_fill_2 FILLER_78_383 ();
 sg13g2_fill_2 FILLER_78_396 ();
 sg13g2_decap_8 FILLER_78_410 ();
 sg13g2_fill_2 FILLER_78_474 ();
 sg13g2_decap_8 FILLER_78_484 ();
 sg13g2_decap_4 FILLER_78_523 ();
 sg13g2_fill_1 FILLER_78_527 ();
 sg13g2_fill_1 FILLER_78_539 ();
 sg13g2_fill_2 FILLER_78_545 ();
 sg13g2_fill_2 FILLER_78_568 ();
 sg13g2_decap_8 FILLER_78_575 ();
 sg13g2_fill_1 FILLER_78_582 ();
 sg13g2_fill_2 FILLER_78_595 ();
 sg13g2_decap_4 FILLER_78_609 ();
 sg13g2_fill_1 FILLER_78_613 ();
 sg13g2_fill_2 FILLER_78_627 ();
 sg13g2_decap_4 FILLER_78_648 ();
 sg13g2_fill_1 FILLER_78_663 ();
 sg13g2_fill_1 FILLER_78_672 ();
 sg13g2_fill_1 FILLER_78_687 ();
 sg13g2_decap_8 FILLER_78_695 ();
 sg13g2_decap_4 FILLER_78_702 ();
 sg13g2_fill_1 FILLER_78_719 ();
 sg13g2_decap_8 FILLER_78_733 ();
 sg13g2_decap_4 FILLER_78_740 ();
 sg13g2_decap_8 FILLER_78_780 ();
 sg13g2_decap_4 FILLER_78_787 ();
 sg13g2_fill_2 FILLER_78_791 ();
 sg13g2_decap_8 FILLER_78_840 ();
 sg13g2_decap_8 FILLER_78_847 ();
 sg13g2_decap_4 FILLER_78_854 ();
 sg13g2_fill_2 FILLER_78_858 ();
 sg13g2_fill_2 FILLER_78_888 ();
 sg13g2_fill_2 FILLER_78_903 ();
 sg13g2_decap_8 FILLER_78_918 ();
 sg13g2_fill_2 FILLER_78_925 ();
 sg13g2_fill_1 FILLER_78_927 ();
 sg13g2_fill_2 FILLER_78_946 ();
 sg13g2_fill_1 FILLER_78_948 ();
 sg13g2_decap_4 FILLER_78_965 ();
 sg13g2_fill_1 FILLER_78_981 ();
 sg13g2_fill_2 FILLER_78_997 ();
 sg13g2_decap_4 FILLER_78_1028 ();
 sg13g2_fill_2 FILLER_78_1032 ();
 sg13g2_decap_8 FILLER_78_1065 ();
 sg13g2_fill_1 FILLER_78_1072 ();
 sg13g2_fill_1 FILLER_78_1090 ();
 sg13g2_fill_1 FILLER_78_1124 ();
 sg13g2_fill_1 FILLER_78_1145 ();
 sg13g2_fill_2 FILLER_78_1169 ();
 sg13g2_fill_1 FILLER_78_1171 ();
 sg13g2_decap_8 FILLER_78_1178 ();
 sg13g2_fill_1 FILLER_78_1189 ();
 sg13g2_fill_1 FILLER_78_1195 ();
 sg13g2_fill_2 FILLER_78_1201 ();
 sg13g2_fill_1 FILLER_78_1203 ();
 sg13g2_fill_1 FILLER_78_1217 ();
 sg13g2_fill_2 FILLER_78_1227 ();
 sg13g2_decap_8 FILLER_78_1239 ();
 sg13g2_decap_4 FILLER_78_1246 ();
 sg13g2_fill_1 FILLER_78_1258 ();
 sg13g2_fill_1 FILLER_78_1287 ();
 sg13g2_decap_8 FILLER_78_1305 ();
 sg13g2_decap_8 FILLER_78_1312 ();
 sg13g2_fill_1 FILLER_78_1319 ();
 sg13g2_fill_1 FILLER_78_1349 ();
 sg13g2_fill_1 FILLER_78_1393 ();
 sg13g2_fill_2 FILLER_78_1398 ();
 sg13g2_fill_1 FILLER_78_1400 ();
 sg13g2_fill_1 FILLER_78_1409 ();
 sg13g2_fill_1 FILLER_78_1423 ();
 sg13g2_fill_1 FILLER_78_1428 ();
 sg13g2_decap_4 FILLER_78_1434 ();
 sg13g2_fill_2 FILLER_78_1446 ();
 sg13g2_fill_1 FILLER_78_1448 ();
 sg13g2_decap_8 FILLER_78_1454 ();
 sg13g2_decap_8 FILLER_78_1461 ();
 sg13g2_decap_8 FILLER_78_1468 ();
 sg13g2_fill_1 FILLER_78_1503 ();
 sg13g2_decap_8 FILLER_78_1509 ();
 sg13g2_decap_8 FILLER_78_1528 ();
 sg13g2_decap_8 FILLER_78_1535 ();
 sg13g2_fill_2 FILLER_78_1542 ();
 sg13g2_fill_1 FILLER_78_1544 ();
 sg13g2_fill_2 FILLER_78_1555 ();
 sg13g2_decap_4 FILLER_78_1565 ();
 sg13g2_fill_2 FILLER_78_1582 ();
 sg13g2_fill_1 FILLER_78_1592 ();
 sg13g2_decap_4 FILLER_78_1605 ();
 sg13g2_fill_1 FILLER_78_1609 ();
 sg13g2_fill_1 FILLER_78_1614 ();
 sg13g2_decap_4 FILLER_78_1620 ();
 sg13g2_fill_1 FILLER_78_1644 ();
 sg13g2_decap_4 FILLER_78_1672 ();
 sg13g2_fill_1 FILLER_78_1676 ();
 sg13g2_decap_8 FILLER_78_1694 ();
 sg13g2_decap_8 FILLER_78_1701 ();
 sg13g2_decap_8 FILLER_78_1708 ();
 sg13g2_decap_8 FILLER_78_1715 ();
 sg13g2_fill_2 FILLER_78_1722 ();
 sg13g2_fill_1 FILLER_78_1724 ();
 sg13g2_decap_8 FILLER_78_1745 ();
 sg13g2_fill_2 FILLER_78_1762 ();
 sg13g2_fill_1 FILLER_78_1764 ();
 sg13g2_decap_4 FILLER_78_1775 ();
 sg13g2_fill_2 FILLER_78_1789 ();
 sg13g2_decap_8 FILLER_78_1837 ();
 sg13g2_decap_4 FILLER_78_1844 ();
 sg13g2_fill_2 FILLER_78_1848 ();
 sg13g2_decap_8 FILLER_78_1869 ();
 sg13g2_fill_2 FILLER_78_1876 ();
 sg13g2_decap_4 FILLER_78_1888 ();
 sg13g2_fill_1 FILLER_78_1896 ();
 sg13g2_decap_8 FILLER_78_1902 ();
 sg13g2_fill_1 FILLER_78_1909 ();
 sg13g2_fill_2 FILLER_78_1916 ();
 sg13g2_fill_1 FILLER_78_1918 ();
 sg13g2_fill_1 FILLER_78_1924 ();
 sg13g2_decap_4 FILLER_78_1930 ();
 sg13g2_decap_8 FILLER_78_1953 ();
 sg13g2_decap_4 FILLER_78_1960 ();
 sg13g2_fill_1 FILLER_78_1974 ();
 sg13g2_decap_8 FILLER_78_1980 ();
 sg13g2_fill_1 FILLER_78_1987 ();
 sg13g2_fill_2 FILLER_78_1997 ();
 sg13g2_decap_4 FILLER_78_2008 ();
 sg13g2_fill_2 FILLER_78_2012 ();
 sg13g2_fill_1 FILLER_78_2024 ();
 sg13g2_fill_1 FILLER_78_2052 ();
 sg13g2_fill_1 FILLER_78_2067 ();
 sg13g2_fill_1 FILLER_78_2073 ();
 sg13g2_decap_8 FILLER_78_2085 ();
 sg13g2_decap_4 FILLER_78_2092 ();
 sg13g2_decap_8 FILLER_78_2099 ();
 sg13g2_decap_4 FILLER_78_2106 ();
 sg13g2_decap_4 FILLER_78_2120 ();
 sg13g2_decap_4 FILLER_78_2145 ();
 sg13g2_fill_1 FILLER_78_2149 ();
 sg13g2_fill_1 FILLER_78_2155 ();
 sg13g2_decap_4 FILLER_78_2166 ();
 sg13g2_fill_2 FILLER_78_2170 ();
 sg13g2_fill_2 FILLER_78_2189 ();
 sg13g2_fill_1 FILLER_78_2191 ();
 sg13g2_decap_8 FILLER_78_2210 ();
 sg13g2_fill_2 FILLER_78_2217 ();
 sg13g2_fill_2 FILLER_78_2227 ();
 sg13g2_fill_1 FILLER_78_2229 ();
 sg13g2_decap_8 FILLER_78_2241 ();
 sg13g2_decap_4 FILLER_78_2252 ();
 sg13g2_fill_1 FILLER_78_2256 ();
 sg13g2_decap_4 FILLER_78_2270 ();
 sg13g2_fill_1 FILLER_78_2274 ();
 sg13g2_fill_2 FILLER_78_2280 ();
 sg13g2_fill_1 FILLER_78_2282 ();
 sg13g2_fill_1 FILLER_78_2303 ();
 sg13g2_decap_4 FILLER_78_2312 ();
 sg13g2_fill_2 FILLER_78_2334 ();
 sg13g2_decap_8 FILLER_78_2354 ();
 sg13g2_fill_2 FILLER_78_2361 ();
 sg13g2_decap_8 FILLER_78_2433 ();
 sg13g2_decap_4 FILLER_78_2440 ();
 sg13g2_fill_1 FILLER_78_2444 ();
 sg13g2_decap_8 FILLER_78_2459 ();
 sg13g2_fill_2 FILLER_78_2478 ();
 sg13g2_fill_1 FILLER_78_2496 ();
 sg13g2_fill_2 FILLER_78_2506 ();
 sg13g2_fill_1 FILLER_78_2539 ();
 sg13g2_fill_2 FILLER_78_2549 ();
 sg13g2_decap_4 FILLER_78_2563 ();
 sg13g2_fill_2 FILLER_78_2567 ();
 sg13g2_decap_8 FILLER_78_2579 ();
 sg13g2_decap_4 FILLER_78_2586 ();
 sg13g2_fill_1 FILLER_78_2590 ();
 sg13g2_fill_1 FILLER_78_2609 ();
 sg13g2_decap_8 FILLER_78_2625 ();
 sg13g2_decap_8 FILLER_78_2632 ();
 sg13g2_fill_1 FILLER_78_2639 ();
 sg13g2_decap_4 FILLER_78_2662 ();
 sg13g2_fill_1 FILLER_78_2666 ();
 sg13g2_fill_2 FILLER_78_2675 ();
 sg13g2_decap_4 FILLER_78_2685 ();
 sg13g2_fill_2 FILLER_78_2689 ();
 sg13g2_fill_2 FILLER_78_2704 ();
 sg13g2_decap_4 FILLER_78_2732 ();
 sg13g2_fill_2 FILLER_78_2748 ();
 sg13g2_fill_1 FILLER_78_2764 ();
 sg13g2_fill_1 FILLER_78_2770 ();
 sg13g2_decap_8 FILLER_78_2776 ();
 sg13g2_fill_2 FILLER_78_2783 ();
 sg13g2_fill_1 FILLER_78_2785 ();
 sg13g2_decap_4 FILLER_78_2806 ();
 sg13g2_fill_2 FILLER_78_2810 ();
 sg13g2_fill_2 FILLER_78_2825 ();
 sg13g2_fill_2 FILLER_78_2836 ();
 sg13g2_decap_4 FILLER_78_2842 ();
 sg13g2_fill_2 FILLER_78_2846 ();
 sg13g2_decap_4 FILLER_78_2890 ();
 sg13g2_fill_2 FILLER_78_2894 ();
 sg13g2_decap_8 FILLER_78_2907 ();
 sg13g2_fill_1 FILLER_78_2914 ();
 sg13g2_decap_8 FILLER_78_2930 ();
 sg13g2_fill_2 FILLER_78_2937 ();
 sg13g2_fill_1 FILLER_78_2939 ();
 sg13g2_fill_2 FILLER_78_2948 ();
 sg13g2_fill_1 FILLER_78_2950 ();
 sg13g2_fill_2 FILLER_78_2964 ();
 sg13g2_fill_1 FILLER_78_2971 ();
 sg13g2_fill_1 FILLER_78_2985 ();
 sg13g2_fill_2 FILLER_78_2995 ();
 sg13g2_fill_1 FILLER_78_2997 ();
 sg13g2_fill_2 FILLER_78_3027 ();
 sg13g2_fill_1 FILLER_78_3029 ();
 sg13g2_fill_1 FILLER_78_3040 ();
 sg13g2_fill_1 FILLER_78_3051 ();
 sg13g2_fill_2 FILLER_78_3058 ();
 sg13g2_fill_1 FILLER_78_3060 ();
 sg13g2_fill_2 FILLER_78_3084 ();
 sg13g2_fill_1 FILLER_78_3086 ();
 sg13g2_decap_8 FILLER_78_3090 ();
 sg13g2_fill_1 FILLER_78_3137 ();
 sg13g2_fill_2 FILLER_78_3143 ();
 sg13g2_decap_8 FILLER_78_3174 ();
 sg13g2_fill_2 FILLER_78_3181 ();
 sg13g2_fill_1 FILLER_78_3183 ();
 sg13g2_fill_2 FILLER_78_3224 ();
 sg13g2_fill_2 FILLER_78_3239 ();
 sg13g2_fill_1 FILLER_78_3241 ();
 sg13g2_decap_4 FILLER_78_3246 ();
 sg13g2_fill_1 FILLER_78_3250 ();
 sg13g2_fill_2 FILLER_78_3257 ();
 sg13g2_fill_2 FILLER_78_3272 ();
 sg13g2_fill_1 FILLER_78_3274 ();
 sg13g2_fill_2 FILLER_78_3279 ();
 sg13g2_fill_2 FILLER_78_3296 ();
 sg13g2_fill_2 FILLER_78_3306 ();
 sg13g2_decap_8 FILLER_78_3320 ();
 sg13g2_decap_4 FILLER_78_3327 ();
 sg13g2_fill_1 FILLER_78_3331 ();
 sg13g2_fill_1 FILLER_78_3369 ();
 sg13g2_fill_1 FILLER_78_3374 ();
 sg13g2_decap_8 FILLER_78_3396 ();
 sg13g2_decap_4 FILLER_78_3403 ();
 sg13g2_fill_2 FILLER_78_3415 ();
 sg13g2_fill_1 FILLER_78_3417 ();
 sg13g2_decap_4 FILLER_78_3423 ();
 sg13g2_fill_2 FILLER_78_3427 ();
 sg13g2_fill_2 FILLER_78_3453 ();
 sg13g2_fill_1 FILLER_78_3455 ();
 sg13g2_fill_1 FILLER_78_3461 ();
 sg13g2_fill_1 FILLER_78_3467 ();
 sg13g2_decap_8 FILLER_78_3479 ();
 sg13g2_fill_2 FILLER_78_3490 ();
 sg13g2_fill_1 FILLER_78_3499 ();
 sg13g2_decap_8 FILLER_78_3509 ();
 sg13g2_decap_4 FILLER_78_3516 ();
 sg13g2_fill_2 FILLER_78_3520 ();
 sg13g2_fill_2 FILLER_78_3527 ();
 sg13g2_fill_2 FILLER_78_3534 ();
 sg13g2_fill_1 FILLER_78_3536 ();
 sg13g2_fill_1 FILLER_78_3555 ();
 sg13g2_decap_4 FILLER_78_3576 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_fill_2 FILLER_79_35 ();
 sg13g2_fill_1 FILLER_79_107 ();
 sg13g2_fill_2 FILLER_79_136 ();
 sg13g2_fill_1 FILLER_79_190 ();
 sg13g2_fill_1 FILLER_79_200 ();
 sg13g2_fill_2 FILLER_79_228 ();
 sg13g2_fill_2 FILLER_79_257 ();
 sg13g2_fill_1 FILLER_79_269 ();
 sg13g2_fill_2 FILLER_79_274 ();
 sg13g2_fill_2 FILLER_79_296 ();
 sg13g2_fill_1 FILLER_79_340 ();
 sg13g2_fill_2 FILLER_79_357 ();
 sg13g2_fill_1 FILLER_79_359 ();
 sg13g2_fill_2 FILLER_79_364 ();
 sg13g2_decap_4 FILLER_79_384 ();
 sg13g2_fill_2 FILLER_79_396 ();
 sg13g2_fill_2 FILLER_79_410 ();
 sg13g2_fill_2 FILLER_79_421 ();
 sg13g2_fill_1 FILLER_79_423 ();
 sg13g2_fill_2 FILLER_79_469 ();
 sg13g2_fill_1 FILLER_79_471 ();
 sg13g2_fill_2 FILLER_79_483 ();
 sg13g2_fill_1 FILLER_79_494 ();
 sg13g2_decap_4 FILLER_79_499 ();
 sg13g2_decap_4 FILLER_79_512 ();
 sg13g2_decap_8 FILLER_79_525 ();
 sg13g2_fill_1 FILLER_79_532 ();
 sg13g2_fill_1 FILLER_79_537 ();
 sg13g2_decap_8 FILLER_79_542 ();
 sg13g2_fill_2 FILLER_79_549 ();
 sg13g2_fill_1 FILLER_79_556 ();
 sg13g2_fill_1 FILLER_79_573 ();
 sg13g2_decap_8 FILLER_79_606 ();
 sg13g2_decap_4 FILLER_79_613 ();
 sg13g2_decap_8 FILLER_79_630 ();
 sg13g2_fill_1 FILLER_79_641 ();
 sg13g2_decap_4 FILLER_79_667 ();
 sg13g2_fill_2 FILLER_79_671 ();
 sg13g2_decap_8 FILLER_79_685 ();
 sg13g2_decap_8 FILLER_79_692 ();
 sg13g2_fill_2 FILLER_79_699 ();
 sg13g2_fill_1 FILLER_79_701 ();
 sg13g2_decap_4 FILLER_79_734 ();
 sg13g2_fill_2 FILLER_79_774 ();
 sg13g2_fill_1 FILLER_79_776 ();
 sg13g2_decap_4 FILLER_79_781 ();
 sg13g2_fill_2 FILLER_79_808 ();
 sg13g2_decap_4 FILLER_79_835 ();
 sg13g2_decap_8 FILLER_79_859 ();
 sg13g2_fill_2 FILLER_79_866 ();
 sg13g2_decap_8 FILLER_79_880 ();
 sg13g2_decap_8 FILLER_79_887 ();
 sg13g2_decap_4 FILLER_79_894 ();
 sg13g2_decap_8 FILLER_79_910 ();
 sg13g2_fill_2 FILLER_79_917 ();
 sg13g2_fill_1 FILLER_79_919 ();
 sg13g2_decap_8 FILLER_79_969 ();
 sg13g2_fill_2 FILLER_79_994 ();
 sg13g2_fill_2 FILLER_79_1004 ();
 sg13g2_fill_1 FILLER_79_1006 ();
 sg13g2_fill_1 FILLER_79_1020 ();
 sg13g2_fill_1 FILLER_79_1045 ();
 sg13g2_decap_4 FILLER_79_1087 ();
 sg13g2_fill_2 FILLER_79_1095 ();
 sg13g2_decap_8 FILLER_79_1116 ();
 sg13g2_fill_1 FILLER_79_1123 ();
 sg13g2_fill_1 FILLER_79_1138 ();
 sg13g2_fill_1 FILLER_79_1201 ();
 sg13g2_fill_2 FILLER_79_1207 ();
 sg13g2_fill_1 FILLER_79_1209 ();
 sg13g2_fill_2 FILLER_79_1218 ();
 sg13g2_fill_1 FILLER_79_1220 ();
 sg13g2_fill_2 FILLER_79_1226 ();
 sg13g2_fill_2 FILLER_79_1241 ();
 sg13g2_fill_2 FILLER_79_1258 ();
 sg13g2_fill_1 FILLER_79_1260 ();
 sg13g2_fill_1 FILLER_79_1266 ();
 sg13g2_fill_1 FILLER_79_1280 ();
 sg13g2_fill_2 FILLER_79_1311 ();
 sg13g2_fill_1 FILLER_79_1313 ();
 sg13g2_fill_1 FILLER_79_1327 ();
 sg13g2_fill_2 FILLER_79_1357 ();
 sg13g2_fill_1 FILLER_79_1359 ();
 sg13g2_decap_4 FILLER_79_1364 ();
 sg13g2_decap_8 FILLER_79_1372 ();
 sg13g2_fill_2 FILLER_79_1379 ();
 sg13g2_fill_1 FILLER_79_1381 ();
 sg13g2_fill_1 FILLER_79_1386 ();
 sg13g2_fill_1 FILLER_79_1426 ();
 sg13g2_decap_8 FILLER_79_1456 ();
 sg13g2_fill_1 FILLER_79_1463 ();
 sg13g2_fill_2 FILLER_79_1502 ();
 sg13g2_fill_1 FILLER_79_1504 ();
 sg13g2_fill_1 FILLER_79_1539 ();
 sg13g2_fill_1 FILLER_79_1560 ();
 sg13g2_decap_4 FILLER_79_1582 ();
 sg13g2_fill_2 FILLER_79_1591 ();
 sg13g2_fill_1 FILLER_79_1593 ();
 sg13g2_fill_1 FILLER_79_1615 ();
 sg13g2_fill_2 FILLER_79_1670 ();
 sg13g2_fill_1 FILLER_79_1672 ();
 sg13g2_fill_1 FILLER_79_1692 ();
 sg13g2_fill_2 FILLER_79_1704 ();
 sg13g2_fill_1 FILLER_79_1706 ();
 sg13g2_fill_2 FILLER_79_1728 ();
 sg13g2_fill_2 FILLER_79_1738 ();
 sg13g2_fill_2 FILLER_79_1755 ();
 sg13g2_fill_2 FILLER_79_1822 ();
 sg13g2_fill_2 FILLER_79_1864 ();
 sg13g2_fill_1 FILLER_79_1866 ();
 sg13g2_decap_4 FILLER_79_1875 ();
 sg13g2_decap_8 FILLER_79_1900 ();
 sg13g2_fill_2 FILLER_79_1907 ();
 sg13g2_fill_1 FILLER_79_1938 ();
 sg13g2_fill_2 FILLER_79_1952 ();
 sg13g2_fill_2 FILLER_79_1966 ();
 sg13g2_fill_2 FILLER_79_1984 ();
 sg13g2_fill_1 FILLER_79_1999 ();
 sg13g2_fill_2 FILLER_79_2008 ();
 sg13g2_fill_1 FILLER_79_2010 ();
 sg13g2_decap_4 FILLER_79_2019 ();
 sg13g2_fill_1 FILLER_79_2038 ();
 sg13g2_fill_2 FILLER_79_2047 ();
 sg13g2_fill_2 FILLER_79_2057 ();
 sg13g2_fill_2 FILLER_79_2083 ();
 sg13g2_decap_8 FILLER_79_2185 ();
 sg13g2_fill_2 FILLER_79_2192 ();
 sg13g2_fill_1 FILLER_79_2215 ();
 sg13g2_fill_1 FILLER_79_2252 ();
 sg13g2_fill_2 FILLER_79_2290 ();
 sg13g2_fill_1 FILLER_79_2292 ();
 sg13g2_fill_2 FILLER_79_2305 ();
 sg13g2_fill_1 FILLER_79_2307 ();
 sg13g2_fill_1 FILLER_79_2322 ();
 sg13g2_decap_8 FILLER_79_2356 ();
 sg13g2_fill_2 FILLER_79_2363 ();
 sg13g2_fill_2 FILLER_79_2373 ();
 sg13g2_fill_1 FILLER_79_2375 ();
 sg13g2_fill_2 FILLER_79_2385 ();
 sg13g2_fill_1 FILLER_79_2399 ();
 sg13g2_decap_4 FILLER_79_2410 ();
 sg13g2_decap_4 FILLER_79_2436 ();
 sg13g2_fill_1 FILLER_79_2440 ();
 sg13g2_fill_2 FILLER_79_2463 ();
 sg13g2_fill_2 FILLER_79_2474 ();
 sg13g2_decap_8 FILLER_79_2492 ();
 sg13g2_fill_2 FILLER_79_2508 ();
 sg13g2_fill_1 FILLER_79_2549 ();
 sg13g2_decap_4 FILLER_79_2564 ();
 sg13g2_fill_2 FILLER_79_2584 ();
 sg13g2_fill_2 FILLER_79_2598 ();
 sg13g2_fill_1 FILLER_79_2600 ();
 sg13g2_fill_1 FILLER_79_2631 ();
 sg13g2_fill_1 FILLER_79_2662 ();
 sg13g2_decap_8 FILLER_79_2685 ();
 sg13g2_fill_2 FILLER_79_2697 ();
 sg13g2_fill_1 FILLER_79_2699 ();
 sg13g2_fill_2 FILLER_79_2705 ();
 sg13g2_fill_1 FILLER_79_2707 ();
 sg13g2_fill_1 FILLER_79_2724 ();
 sg13g2_decap_8 FILLER_79_2738 ();
 sg13g2_fill_1 FILLER_79_2759 ();
 sg13g2_fill_2 FILLER_79_2823 ();
 sg13g2_fill_2 FILLER_79_2833 ();
 sg13g2_fill_1 FILLER_79_2835 ();
 sg13g2_fill_2 FILLER_79_2847 ();
 sg13g2_fill_2 FILLER_79_2912 ();
 sg13g2_fill_1 FILLER_79_2914 ();
 sg13g2_fill_1 FILLER_79_2936 ();
 sg13g2_fill_2 FILLER_79_2971 ();
 sg13g2_fill_2 FILLER_79_3008 ();
 sg13g2_fill_1 FILLER_79_3010 ();
 sg13g2_fill_2 FILLER_79_3108 ();
 sg13g2_fill_2 FILLER_79_3123 ();
 sg13g2_decap_4 FILLER_79_3146 ();
 sg13g2_decap_4 FILLER_79_3222 ();
 sg13g2_fill_1 FILLER_79_3242 ();
 sg13g2_decap_4 FILLER_79_3256 ();
 sg13g2_fill_1 FILLER_79_3260 ();
 sg13g2_fill_1 FILLER_79_3269 ();
 sg13g2_fill_2 FILLER_79_3274 ();
 sg13g2_fill_2 FILLER_79_3292 ();
 sg13g2_fill_1 FILLER_79_3294 ();
 sg13g2_decap_8 FILLER_79_3320 ();
 sg13g2_decap_4 FILLER_79_3327 ();
 sg13g2_decap_4 FILLER_79_3342 ();
 sg13g2_fill_1 FILLER_79_3374 ();
 sg13g2_fill_1 FILLER_79_3394 ();
 sg13g2_fill_1 FILLER_79_3399 ();
 sg13g2_fill_2 FILLER_79_3432 ();
 sg13g2_decap_4 FILLER_79_3450 ();
 sg13g2_fill_2 FILLER_79_3454 ();
 sg13g2_fill_1 FILLER_79_3489 ();
 sg13g2_fill_2 FILLER_79_3511 ();
 sg13g2_fill_2 FILLER_79_3545 ();
 sg13g2_fill_2 FILLER_79_3577 ();
 sg13g2_fill_1 FILLER_79_3579 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_fill_2 FILLER_80_28 ();
 sg13g2_fill_1 FILLER_80_67 ();
 sg13g2_fill_1 FILLER_80_81 ();
 sg13g2_fill_1 FILLER_80_144 ();
 sg13g2_fill_2 FILLER_80_176 ();
 sg13g2_fill_2 FILLER_80_261 ();
 sg13g2_fill_1 FILLER_80_279 ();
 sg13g2_fill_1 FILLER_80_296 ();
 sg13g2_fill_2 FILLER_80_331 ();
 sg13g2_decap_4 FILLER_80_373 ();
 sg13g2_fill_2 FILLER_80_382 ();
 sg13g2_decap_8 FILLER_80_405 ();
 sg13g2_decap_4 FILLER_80_444 ();
 sg13g2_decap_8 FILLER_80_453 ();
 sg13g2_decap_4 FILLER_80_460 ();
 sg13g2_fill_2 FILLER_80_472 ();
 sg13g2_fill_1 FILLER_80_474 ();
 sg13g2_decap_8 FILLER_80_488 ();
 sg13g2_fill_1 FILLER_80_495 ();
 sg13g2_decap_8 FILLER_80_556 ();
 sg13g2_fill_2 FILLER_80_563 ();
 sg13g2_fill_2 FILLER_80_573 ();
 sg13g2_fill_2 FILLER_80_579 ();
 sg13g2_decap_8 FILLER_80_600 ();
 sg13g2_decap_4 FILLER_80_607 ();
 sg13g2_fill_2 FILLER_80_642 ();
 sg13g2_fill_1 FILLER_80_644 ();
 sg13g2_decap_8 FILLER_80_661 ();
 sg13g2_decap_8 FILLER_80_700 ();
 sg13g2_decap_4 FILLER_80_725 ();
 sg13g2_fill_2 FILLER_80_729 ();
 sg13g2_decap_8 FILLER_80_734 ();
 sg13g2_decap_4 FILLER_80_741 ();
 sg13g2_decap_4 FILLER_80_754 ();
 sg13g2_decap_8 FILLER_80_763 ();
 sg13g2_fill_1 FILLER_80_770 ();
 sg13g2_fill_2 FILLER_80_799 ();
 sg13g2_fill_1 FILLER_80_801 ();
 sg13g2_fill_2 FILLER_80_824 ();
 sg13g2_fill_1 FILLER_80_826 ();
 sg13g2_decap_8 FILLER_80_831 ();
 sg13g2_decap_4 FILLER_80_866 ();
 sg13g2_fill_1 FILLER_80_870 ();
 sg13g2_fill_2 FILLER_80_899 ();
 sg13g2_decap_8 FILLER_80_937 ();
 sg13g2_decap_4 FILLER_80_944 ();
 sg13g2_fill_1 FILLER_80_948 ();
 sg13g2_fill_2 FILLER_80_954 ();
 sg13g2_fill_1 FILLER_80_956 ();
 sg13g2_decap_8 FILLER_80_962 ();
 sg13g2_decap_8 FILLER_80_969 ();
 sg13g2_decap_8 FILLER_80_976 ();
 sg13g2_fill_2 FILLER_80_983 ();
 sg13g2_fill_2 FILLER_80_990 ();
 sg13g2_fill_1 FILLER_80_992 ();
 sg13g2_fill_1 FILLER_80_1001 ();
 sg13g2_decap_4 FILLER_80_1028 ();
 sg13g2_fill_1 FILLER_80_1032 ();
 sg13g2_fill_2 FILLER_80_1046 ();
 sg13g2_fill_1 FILLER_80_1048 ();
 sg13g2_fill_1 FILLER_80_1055 ();
 sg13g2_decap_8 FILLER_80_1064 ();
 sg13g2_fill_2 FILLER_80_1071 ();
 sg13g2_fill_2 FILLER_80_1083 ();
 sg13g2_fill_1 FILLER_80_1085 ();
 sg13g2_decap_4 FILLER_80_1114 ();
 sg13g2_decap_8 FILLER_80_1134 ();
 sg13g2_decap_4 FILLER_80_1141 ();
 sg13g2_decap_8 FILLER_80_1162 ();
 sg13g2_decap_8 FILLER_80_1169 ();
 sg13g2_decap_8 FILLER_80_1176 ();
 sg13g2_decap_4 FILLER_80_1183 ();
 sg13g2_fill_1 FILLER_80_1187 ();
 sg13g2_fill_1 FILLER_80_1201 ();
 sg13g2_fill_1 FILLER_80_1215 ();
 sg13g2_decap_8 FILLER_80_1232 ();
 sg13g2_fill_1 FILLER_80_1239 ();
 sg13g2_decap_8 FILLER_80_1258 ();
 sg13g2_decap_8 FILLER_80_1265 ();
 sg13g2_fill_2 FILLER_80_1272 ();
 sg13g2_decap_8 FILLER_80_1278 ();
 sg13g2_decap_4 FILLER_80_1285 ();
 sg13g2_fill_2 FILLER_80_1289 ();
 sg13g2_decap_8 FILLER_80_1308 ();
 sg13g2_decap_4 FILLER_80_1315 ();
 sg13g2_fill_1 FILLER_80_1332 ();
 sg13g2_fill_2 FILLER_80_1355 ();
 sg13g2_fill_1 FILLER_80_1357 ();
 sg13g2_decap_4 FILLER_80_1368 ();
 sg13g2_fill_1 FILLER_80_1372 ();
 sg13g2_decap_4 FILLER_80_1386 ();
 sg13g2_fill_1 FILLER_80_1393 ();
 sg13g2_decap_8 FILLER_80_1403 ();
 sg13g2_decap_8 FILLER_80_1422 ();
 sg13g2_decap_8 FILLER_80_1429 ();
 sg13g2_fill_1 FILLER_80_1446 ();
 sg13g2_fill_2 FILLER_80_1452 ();
 sg13g2_fill_1 FILLER_80_1454 ();
 sg13g2_decap_8 FILLER_80_1460 ();
 sg13g2_decap_4 FILLER_80_1467 ();
 sg13g2_fill_2 FILLER_80_1484 ();
 sg13g2_decap_8 FILLER_80_1509 ();
 sg13g2_fill_1 FILLER_80_1516 ();
 sg13g2_fill_1 FILLER_80_1527 ();
 sg13g2_decap_8 FILLER_80_1533 ();
 sg13g2_decap_8 FILLER_80_1540 ();
 sg13g2_decap_4 FILLER_80_1557 ();
 sg13g2_decap_4 FILLER_80_1565 ();
 sg13g2_decap_4 FILLER_80_1572 ();
 sg13g2_fill_1 FILLER_80_1576 ();
 sg13g2_decap_4 FILLER_80_1581 ();
 sg13g2_fill_1 FILLER_80_1594 ();
 sg13g2_decap_8 FILLER_80_1599 ();
 sg13g2_decap_8 FILLER_80_1606 ();
 sg13g2_decap_8 FILLER_80_1613 ();
 sg13g2_fill_2 FILLER_80_1620 ();
 sg13g2_fill_1 FILLER_80_1622 ();
 sg13g2_decap_8 FILLER_80_1644 ();
 sg13g2_decap_4 FILLER_80_1651 ();
 sg13g2_fill_1 FILLER_80_1655 ();
 sg13g2_fill_2 FILLER_80_1664 ();
 sg13g2_decap_4 FILLER_80_1670 ();
 sg13g2_fill_2 FILLER_80_1686 ();
 sg13g2_decap_8 FILLER_80_1694 ();
 sg13g2_fill_2 FILLER_80_1701 ();
 sg13g2_decap_4 FILLER_80_1720 ();
 sg13g2_fill_1 FILLER_80_1724 ();
 sg13g2_decap_8 FILLER_80_1744 ();
 sg13g2_decap_4 FILLER_80_1751 ();
 sg13g2_decap_8 FILLER_80_1774 ();
 sg13g2_decap_8 FILLER_80_1786 ();
 sg13g2_decap_8 FILLER_80_1793 ();
 sg13g2_fill_1 FILLER_80_1826 ();
 sg13g2_fill_2 FILLER_80_1831 ();
 sg13g2_fill_2 FILLER_80_1850 ();
 sg13g2_fill_1 FILLER_80_1860 ();
 sg13g2_decap_8 FILLER_80_1870 ();
 sg13g2_decap_4 FILLER_80_1877 ();
 sg13g2_fill_1 FILLER_80_1881 ();
 sg13g2_fill_1 FILLER_80_1887 ();
 sg13g2_fill_2 FILLER_80_1898 ();
 sg13g2_decap_8 FILLER_80_1911 ();
 sg13g2_fill_2 FILLER_80_1918 ();
 sg13g2_decap_8 FILLER_80_1938 ();
 sg13g2_decap_8 FILLER_80_1945 ();
 sg13g2_decap_4 FILLER_80_1952 ();
 sg13g2_fill_1 FILLER_80_1956 ();
 sg13g2_fill_1 FILLER_80_1967 ();
 sg13g2_decap_8 FILLER_80_1973 ();
 sg13g2_decap_4 FILLER_80_1980 ();
 sg13g2_decap_8 FILLER_80_1996 ();
 sg13g2_decap_8 FILLER_80_2003 ();
 sg13g2_decap_4 FILLER_80_2010 ();
 sg13g2_decap_8 FILLER_80_2035 ();
 sg13g2_fill_1 FILLER_80_2042 ();
 sg13g2_decap_8 FILLER_80_2048 ();
 sg13g2_decap_4 FILLER_80_2055 ();
 sg13g2_fill_2 FILLER_80_2059 ();
 sg13g2_decap_8 FILLER_80_2075 ();
 sg13g2_decap_4 FILLER_80_2082 ();
 sg13g2_fill_1 FILLER_80_2086 ();
 sg13g2_decap_8 FILLER_80_2107 ();
 sg13g2_decap_4 FILLER_80_2114 ();
 sg13g2_fill_1 FILLER_80_2118 ();
 sg13g2_decap_8 FILLER_80_2141 ();
 sg13g2_fill_2 FILLER_80_2148 ();
 sg13g2_decap_4 FILLER_80_2168 ();
 sg13g2_fill_2 FILLER_80_2172 ();
 sg13g2_fill_2 FILLER_80_2187 ();
 sg13g2_fill_1 FILLER_80_2189 ();
 sg13g2_decap_8 FILLER_80_2214 ();
 sg13g2_fill_2 FILLER_80_2221 ();
 sg13g2_decap_8 FILLER_80_2237 ();
 sg13g2_decap_8 FILLER_80_2244 ();
 sg13g2_fill_2 FILLER_80_2251 ();
 sg13g2_fill_1 FILLER_80_2253 ();
 sg13g2_decap_8 FILLER_80_2271 ();
 sg13g2_fill_1 FILLER_80_2278 ();
 sg13g2_decap_4 FILLER_80_2283 ();
 sg13g2_fill_2 FILLER_80_2287 ();
 sg13g2_decap_8 FILLER_80_2312 ();
 sg13g2_decap_8 FILLER_80_2319 ();
 sg13g2_fill_2 FILLER_80_2326 ();
 sg13g2_fill_1 FILLER_80_2328 ();
 sg13g2_fill_2 FILLER_80_2349 ();
 sg13g2_fill_2 FILLER_80_2391 ();
 sg13g2_fill_1 FILLER_80_2393 ();
 sg13g2_fill_1 FILLER_80_2478 ();
 sg13g2_fill_1 FILLER_80_2511 ();
 sg13g2_decap_8 FILLER_80_2540 ();
 sg13g2_fill_2 FILLER_80_2551 ();
 sg13g2_fill_1 FILLER_80_2553 ();
 sg13g2_decap_8 FILLER_80_2559 ();
 sg13g2_decap_4 FILLER_80_2566 ();
 sg13g2_decap_8 FILLER_80_2587 ();
 sg13g2_decap_4 FILLER_80_2594 ();
 sg13g2_fill_1 FILLER_80_2598 ();
 sg13g2_decap_4 FILLER_80_2603 ();
 sg13g2_decap_8 FILLER_80_2624 ();
 sg13g2_decap_8 FILLER_80_2631 ();
 sg13g2_decap_4 FILLER_80_2638 ();
 sg13g2_fill_1 FILLER_80_2642 ();
 sg13g2_decap_8 FILLER_80_2659 ();
 sg13g2_decap_4 FILLER_80_2666 ();
 sg13g2_fill_2 FILLER_80_2679 ();
 sg13g2_fill_1 FILLER_80_2681 ();
 sg13g2_decap_8 FILLER_80_2695 ();
 sg13g2_decap_4 FILLER_80_2702 ();
 sg13g2_fill_2 FILLER_80_2706 ();
 sg13g2_fill_1 FILLER_80_2730 ();
 sg13g2_decap_8 FILLER_80_2739 ();
 sg13g2_decap_8 FILLER_80_2746 ();
 sg13g2_fill_2 FILLER_80_2753 ();
 sg13g2_fill_1 FILLER_80_2755 ();
 sg13g2_fill_2 FILLER_80_2761 ();
 sg13g2_decap_8 FILLER_80_2776 ();
 sg13g2_decap_8 FILLER_80_2783 ();
 sg13g2_fill_1 FILLER_80_2790 ();
 sg13g2_decap_8 FILLER_80_2806 ();
 sg13g2_decap_4 FILLER_80_2831 ();
 sg13g2_fill_2 FILLER_80_2835 ();
 sg13g2_decap_8 FILLER_80_2845 ();
 sg13g2_decap_8 FILLER_80_2856 ();
 sg13g2_decap_8 FILLER_80_2863 ();
 sg13g2_fill_2 FILLER_80_2870 ();
 sg13g2_fill_1 FILLER_80_2872 ();
 sg13g2_decap_8 FILLER_80_2888 ();
 sg13g2_fill_2 FILLER_80_2895 ();
 sg13g2_fill_1 FILLER_80_2897 ();
 sg13g2_decap_8 FILLER_80_2906 ();
 sg13g2_decap_4 FILLER_80_2913 ();
 sg13g2_decap_8 FILLER_80_2931 ();
 sg13g2_decap_8 FILLER_80_2938 ();
 sg13g2_decap_8 FILLER_80_2945 ();
 sg13g2_decap_4 FILLER_80_2952 ();
 sg13g2_decap_4 FILLER_80_2961 ();
 sg13g2_fill_1 FILLER_80_2965 ();
 sg13g2_decap_4 FILLER_80_2993 ();
 sg13g2_fill_2 FILLER_80_2997 ();
 sg13g2_decap_8 FILLER_80_3027 ();
 sg13g2_decap_8 FILLER_80_3034 ();
 sg13g2_decap_8 FILLER_80_3041 ();
 sg13g2_decap_8 FILLER_80_3048 ();
 sg13g2_fill_1 FILLER_80_3055 ();
 sg13g2_fill_2 FILLER_80_3060 ();
 sg13g2_fill_1 FILLER_80_3062 ();
 sg13g2_decap_4 FILLER_80_3067 ();
 sg13g2_fill_2 FILLER_80_3071 ();
 sg13g2_decap_8 FILLER_80_3082 ();
 sg13g2_decap_8 FILLER_80_3089 ();
 sg13g2_fill_2 FILLER_80_3096 ();
 sg13g2_fill_1 FILLER_80_3098 ();
 sg13g2_fill_1 FILLER_80_3104 ();
 sg13g2_decap_8 FILLER_80_3115 ();
 sg13g2_fill_1 FILLER_80_3126 ();
 sg13g2_decap_8 FILLER_80_3139 ();
 sg13g2_decap_8 FILLER_80_3146 ();
 sg13g2_fill_2 FILLER_80_3153 ();
 sg13g2_decap_8 FILLER_80_3169 ();
 sg13g2_decap_8 FILLER_80_3176 ();
 sg13g2_decap_4 FILLER_80_3183 ();
 sg13g2_fill_2 FILLER_80_3187 ();
 sg13g2_decap_4 FILLER_80_3207 ();
 sg13g2_fill_1 FILLER_80_3211 ();
 sg13g2_fill_2 FILLER_80_3222 ();
 sg13g2_fill_1 FILLER_80_3224 ();
 sg13g2_decap_8 FILLER_80_3237 ();
 sg13g2_decap_4 FILLER_80_3244 ();
 sg13g2_decap_8 FILLER_80_3253 ();
 sg13g2_decap_4 FILLER_80_3273 ();
 sg13g2_decap_8 FILLER_80_3292 ();
 sg13g2_fill_1 FILLER_80_3299 ();
 sg13g2_decap_8 FILLER_80_3312 ();
 sg13g2_fill_2 FILLER_80_3319 ();
 sg13g2_fill_1 FILLER_80_3321 ();
 sg13g2_decap_8 FILLER_80_3343 ();
 sg13g2_fill_2 FILLER_80_3350 ();
 sg13g2_fill_1 FILLER_80_3352 ();
 sg13g2_decap_8 FILLER_80_3365 ();
 sg13g2_decap_8 FILLER_80_3372 ();
 sg13g2_decap_8 FILLER_80_3398 ();
 sg13g2_fill_1 FILLER_80_3405 ();
 sg13g2_fill_1 FILLER_80_3414 ();
 sg13g2_fill_1 FILLER_80_3424 ();
 sg13g2_decap_4 FILLER_80_3435 ();
 sg13g2_fill_2 FILLER_80_3439 ();
 sg13g2_decap_4 FILLER_80_3454 ();
 sg13g2_fill_2 FILLER_80_3458 ();
 sg13g2_decap_8 FILLER_80_3477 ();
 sg13g2_decap_4 FILLER_80_3484 ();
 sg13g2_decap_8 FILLER_80_3506 ();
 sg13g2_decap_8 FILLER_80_3513 ();
 sg13g2_fill_2 FILLER_80_3520 ();
 sg13g2_fill_1 FILLER_80_3526 ();
 sg13g2_decap_8 FILLER_80_3532 ();
 sg13g2_decap_8 FILLER_80_3539 ();
 sg13g2_fill_2 FILLER_80_3546 ();
 sg13g2_fill_1 FILLER_80_3548 ();
 sg13g2_decap_4 FILLER_80_3558 ();
 sg13g2_decap_4 FILLER_80_3575 ();
 sg13g2_fill_1 FILLER_80_3579 ();
 assign uio_oe[0] = net1059;
 assign uio_oe[1] = net1060;
 assign uio_oe[2] = net14;
 assign uio_oe[3] = net15;
 assign uio_oe[4] = net1061;
 assign uio_oe[5] = net1062;
 assign uio_oe[6] = net1063;
 assign uio_oe[7] = net16;
 assign uio_out[2] = net17;
 assign uio_out[3] = net18;
 assign uio_out[5] = net19;
 assign uio_out[7] = net20;
endmodule
