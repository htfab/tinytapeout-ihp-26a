module tt_um_snake_game (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire audio;
 wire eat;
 wire failure;
 wire \game_inst.apple_inst.apple_x[0] ;
 wire \game_inst.apple_inst.apple_x[1] ;
 wire \game_inst.apple_inst.apple_x[2] ;
 wire \game_inst.apple_inst.apple_x[3] ;
 wire \game_inst.apple_inst.apple_x[4] ;
 wire \game_inst.apple_inst.apple_y[0] ;
 wire \game_inst.apple_inst.apple_y[1] ;
 wire \game_inst.apple_inst.apple_y[2] ;
 wire \game_inst.apple_inst.apple_y[3] ;
 wire \game_inst.apple_inst.i_snake_valid ;
 wire \game_inst.apple_inst.i_snake_x[0] ;
 wire \game_inst.apple_inst.i_snake_x[1] ;
 wire \game_inst.apple_inst.i_snake_x[2] ;
 wire \game_inst.apple_inst.i_snake_x[3] ;
 wire \game_inst.apple_inst.i_snake_x[4] ;
 wire \game_inst.apple_inst.i_snake_y[0] ;
 wire \game_inst.apple_inst.i_snake_y[1] ;
 wire \game_inst.apple_inst.i_snake_y[2] ;
 wire \game_inst.apple_inst.i_snake_y[3] ;
 wire \game_inst.apple_inst.o_ready ;
 wire \game_inst.apple_inst.random_inst.lfsr4[0] ;
 wire \game_inst.apple_inst.random_inst.lfsr4[1] ;
 wire \game_inst.apple_inst.random_inst.lfsr4[2] ;
 wire \game_inst.apple_inst.random_inst.lfsr4[3] ;
 wire \game_inst.apple_inst.random_inst.lfsr5[0] ;
 wire \game_inst.apple_inst.random_inst.lfsr5[1] ;
 wire \game_inst.apple_inst.random_inst.lfsr5[2] ;
 wire \game_inst.apple_inst.random_inst.lfsr5[3] ;
 wire \game_inst.apple_inst.random_inst.lfsr5[4] ;
 wire \game_inst.apple_inst.test ;
 wire \game_inst.control_inst.backwards[1] ;
 wire \game_inst.control_inst.dir[0] ;
 wire \game_inst.control_inst.dir[1] ;
 wire \game_inst.control_inst.i_head_dir[0] ;
 wire \game_inst.control_inst.o_start ;
 wire \game_inst.head_x[0] ;
 wire \game_inst.head_x[1] ;
 wire \game_inst.head_x[2] ;
 wire \game_inst.head_x[3] ;
 wire \game_inst.head_x[4] ;
 wire \game_inst.head_y[0] ;
 wire \game_inst.head_y[1] ;
 wire \game_inst.head_y[2] ;
 wire \game_inst.head_y[3] ;
 wire \game_inst.o_success ;
 wire \game_inst.o_tick ;
 wire \game_inst.o_vga_hsync ;
 wire \game_inst.o_vga_vsync ;
 wire \game_inst.pwm_base ;
 wire \game_inst.snake_inst.length[0] ;
 wire \game_inst.snake_inst.length[1] ;
 wire \game_inst.snake_inst.length[2] ;
 wire \game_inst.snake_inst.length[3] ;
 wire \game_inst.snake_inst.length[4] ;
 wire \game_inst.snake_inst.length[5] ;
 wire \game_inst.snake_inst.length[6] ;
 wire \game_inst.snake_inst.length[7] ;
 wire \game_inst.snake_inst.pos[0] ;
 wire \game_inst.snake_inst.pos[1] ;
 wire \game_inst.snake_inst.pos[2] ;
 wire \game_inst.snake_inst.pos[3] ;
 wire \game_inst.snake_inst.pos[4] ;
 wire \game_inst.snake_inst.pos[5] ;
 wire \game_inst.snake_inst.pos[6] ;
 wire \game_inst.snake_inst.pos[7] ;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire clknet_leaf_0_clk;
 wire \game_inst.sound_inst.counter[0] ;
 wire \game_inst.sound_inst.counter[1] ;
 wire \game_inst.sound_inst.counter[2] ;
 wire \game_inst.sound_inst.counter[3] ;
 wire \game_inst.sound_inst.max_counter[0] ;
 wire \game_inst.sound_inst.max_counter[1] ;
 wire \game_inst.sound_inst.max_counter[2] ;
 wire \game_inst.sound_inst.max_counter[3] ;
 wire \game_inst.sound_inst.mode[0] ;
 wire \game_inst.sound_inst.mode[1] ;
 wire \game_inst.sound_inst.phase[0] ;
 wire \game_inst.sound_inst.phase[1] ;
 wire \game_inst.sound_inst.phase[2] ;
 wire \game_inst.sound_inst.phase[3] ;
 wire \game_inst.sound_inst.phase[4] ;
 wire \game_inst.sound_inst.prev_pwm_base ;
 wire \game_inst.sound_inst.prev_vsync ;
 wire \game_inst.sound_inst.vsync_pulse ;
 wire \game_inst.tick ;
 wire \game_inst.tickgen_inst.counter[0] ;
 wire \game_inst.tickgen_inst.counter[1] ;
 wire \game_inst.tickgen_inst.counter[2] ;
 wire \game_inst.tickgen_inst.counter[3] ;
 wire \game_inst.tickgen_inst.counter_max[1] ;
 wire \game_inst.tickgen_inst.counter_max[2] ;
 wire \game_inst.tickgen_inst.counter_max[3] ;
 wire \game_inst.tickgen_inst.prev_user_input ;
 wire \game_inst.vga_inst.color[1] ;
 wire \game_inst.vga_inst.color[2] ;
 wire \game_inst.vga_inst.color[3] ;
 wire \game_inst.vga_inst.prev_dir[0] ;
 wire \game_inst.vga_inst.prev_dir[1] ;
 wire \game_inst.vga_inst.px[0] ;
 wire \game_inst.vga_inst.px[1] ;
 wire \game_inst.vga_inst.px[2] ;
 wire \game_inst.vga_inst.px[3] ;
 wire \game_inst.vga_inst.px[4] ;
 wire \game_inst.vga_inst.px[5] ;
 wire \game_inst.vga_inst.px[6] ;
 wire \game_inst.vga_inst.px[7] ;
 wire \game_inst.vga_inst.px[8] ;
 wire \game_inst.vga_inst.px[9] ;
 wire \game_inst.vga_inst.py[0] ;
 wire \game_inst.vga_inst.py[1] ;
 wire \game_inst.vga_inst.py[2] ;
 wire \game_inst.vga_inst.py[4] ;
 wire \game_inst.vga_inst.py[5] ;
 wire \game_inst.vga_inst.py[6] ;
 wire \game_inst.vga_inst.py[7] ;
 wire \game_inst.vga_inst.py[8] ;
 wire \game_inst.vga_inst.py[9] ;
 wire \game_inst.vga_inst.row_buffer[0][0] ;
 wire \game_inst.vga_inst.row_buffer[0][1] ;
 wire \game_inst.vga_inst.row_buffer[0][2] ;
 wire \game_inst.vga_inst.row_buffer[0][3] ;
 wire \game_inst.vga_inst.row_buffer[1][0] ;
 wire \game_inst.vga_inst.row_buffer[1][1] ;
 wire \game_inst.vga_inst.row_buffer[1][2] ;
 wire \game_inst.vga_inst.row_buffer[1][3] ;
 wire \game_inst.vga_inst.row_buffer[2][0] ;
 wire \game_inst.vga_inst.row_buffer[2][1] ;
 wire \game_inst.vga_inst.row_buffer[2][2] ;
 wire \game_inst.vga_inst.row_buffer[2][3] ;
 wire \game_inst.vga_inst.row_buffer[3][0] ;
 wire \game_inst.vga_inst.row_buffer[3][1] ;
 wire \game_inst.vga_inst.row_buffer[3][2] ;
 wire \game_inst.vga_inst.row_buffer[3][3] ;
 wire \game_inst.vga_inst.row_buffer[4][0] ;
 wire \game_inst.vga_inst.row_buffer[4][1] ;
 wire \game_inst.vga_inst.row_buffer[4][2] ;
 wire \game_inst.vga_inst.row_buffer[4][3] ;
 wire \game_inst.vga_inst.row_buffer[5][0] ;
 wire \game_inst.vga_inst.row_buffer[5][1] ;
 wire \game_inst.vga_inst.row_buffer[5][2] ;
 wire \game_inst.vga_inst.row_buffer[5][3] ;
 wire \game_inst.vga_inst.row_buffer[6][0] ;
 wire \game_inst.vga_inst.row_buffer[6][1] ;
 wire \game_inst.vga_inst.row_buffer[6][2] ;
 wire \game_inst.vga_inst.row_buffer[6][3] ;
 wire \game_inst.vga_inst.row_buffer[7][0] ;
 wire \game_inst.vga_inst.row_buffer[7][1] ;
 wire \game_inst.vga_inst.row_buffer[7][2] ;
 wire \game_inst.vga_inst.row_buffer[7][3] ;
 wire \game_inst.vga_inst.row_buffer[8][0] ;
 wire \game_inst.vga_inst.row_buffer[8][1] ;
 wire \game_inst.vga_inst.row_buffer[8][2] ;
 wire \game_inst.vga_inst.row_buffer[8][3] ;
 wire \game_inst.vga_inst.s_hsync ;
 wire \game_inst.vga_inst.s_vsync ;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net8;
 wire net9;
 wire net10;
 wire net222;
 wire net11;
 wire net12;
 wire net13;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[0] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[100] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[101] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[102] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[103] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[104] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[105] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[106] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[107] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[108] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[109] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[10] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[110] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[111] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[112] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[113] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[114] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[115] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[116] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[117] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[118] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[119] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[11] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[120] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[121] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[122] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[123] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[124] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[125] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[126] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[127] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[128] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[129] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[12] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[130] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[131] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[132] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[133] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[134] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[135] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[136] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[137] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[138] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[139] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[13] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[140] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[141] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[142] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[143] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[144] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[145] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[146] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[147] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[148] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[149] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[14] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[150] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[151] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[152] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[153] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[154] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[155] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[156] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[157] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[158] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[159] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[15] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[160] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[161] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[162] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[163] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[164] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[165] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[166] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[167] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[168] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[169] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[16] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[170] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[171] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[172] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[173] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[174] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[175] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[176] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[177] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[178] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[179] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[17] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[180] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[181] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[182] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[183] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[184] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[185] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[186] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[187] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[188] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[189] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[18] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[190] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[191] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[192] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[193] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[194] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[195] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[196] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[197] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[198] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[199] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[19] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[1] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[200] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[201] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[202] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[203] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[204] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[205] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[206] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[207] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[208] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[209] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[20] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[210] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[211] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[212] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[213] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[214] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[215] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[216] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[217] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[218] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[219] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[21] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[220] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[221] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[222] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[223] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[224] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[225] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[226] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[227] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[228] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[229] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[22] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[230] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[231] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[232] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[233] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[23] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[24] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[25] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[26] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[27] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[28] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[29] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[2] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[30] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[31] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[32] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[33] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[34] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[35] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[36] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[37] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[38] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[39] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[3] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[40] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[41] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[42] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[43] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[44] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[45] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[46] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[47] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[48] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[49] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[4] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[50] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[51] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[52] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[53] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[54] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[55] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[56] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[57] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[58] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[59] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[5] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[60] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[61] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[62] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[63] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[64] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[65] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[66] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[67] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[68] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[69] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[6] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[70] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[71] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[72] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[73] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[74] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[75] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[76] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[77] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[78] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[79] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[7] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[80] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[81] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[82] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[83] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[84] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[85] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[86] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[87] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[88] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[89] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[8] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[90] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[91] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[92] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[93] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[94] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[95] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[96] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[97] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[98] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[99] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[9] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[0] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[100] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[101] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[102] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[103] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[104] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[105] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[106] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[107] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[108] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[109] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[10] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[110] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[111] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[112] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[113] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[114] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[115] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[116] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[117] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[118] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[119] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[11] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[120] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[121] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[122] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[123] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[124] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[125] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[126] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[127] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[128] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[129] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[12] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[130] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[131] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[132] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[133] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[134] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[135] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[136] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[137] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[138] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[139] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[13] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[140] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[141] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[142] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[143] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[144] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[145] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[146] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[147] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[148] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[149] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[14] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[150] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[151] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[152] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[153] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[154] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[155] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[156] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[157] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[158] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[159] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[15] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[160] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[161] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[162] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[163] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[164] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[165] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[166] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[167] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[168] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[169] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[16] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[170] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[171] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[172] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[173] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[174] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[175] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[176] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[177] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[178] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[179] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[17] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[180] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[181] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[182] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[183] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[184] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[185] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[186] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[187] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[188] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[189] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[18] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[190] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[191] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[192] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[193] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[194] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[195] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[196] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[197] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[198] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[199] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[19] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[1] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[200] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[201] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[202] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[203] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[204] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[205] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[206] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[207] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[208] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[209] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[20] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[210] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[211] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[212] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[213] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[214] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[215] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[216] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[217] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[218] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[219] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[21] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[220] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[221] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[222] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[223] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[224] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[225] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[226] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[227] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[228] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[229] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[22] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[230] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[231] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[232] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[233] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[23] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[24] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[25] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[26] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[27] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[28] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[29] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[2] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[30] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[31] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[32] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[33] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[34] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[35] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[36] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[37] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[38] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[39] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[3] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[40] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[41] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[42] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[43] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[44] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[45] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[46] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[47] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[48] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[49] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[4] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[50] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[51] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[52] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[53] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[54] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[55] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[56] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[57] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[58] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[59] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[5] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[60] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[61] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[62] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[63] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[64] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[65] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[66] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[67] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[68] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[69] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[6] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[70] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[71] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[72] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[73] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[74] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[75] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[76] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[77] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[78] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[79] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[7] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[80] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[81] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[82] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[83] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[84] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[85] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[86] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[87] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[88] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[89] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[8] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[90] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[91] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[92] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[93] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[94] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[95] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[96] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[97] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[98] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[99] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[9] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[0] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[100] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[101] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[102] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[103] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[104] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[105] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[106] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[107] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[108] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[109] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[10] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[110] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[111] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[112] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[113] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[114] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[115] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[116] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[117] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[118] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[119] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[11] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[120] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[121] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[122] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[123] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[124] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[125] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[126] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[127] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[128] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[129] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[12] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[130] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[131] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[132] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[133] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[134] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[135] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[136] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[137] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[138] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[139] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[13] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[140] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[141] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[142] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[143] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[144] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[145] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[146] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[147] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[148] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[149] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[14] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[150] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[151] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[152] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[153] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[154] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[155] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[156] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[157] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[158] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[159] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[15] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[160] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[161] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[162] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[163] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[164] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[165] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[166] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[167] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[168] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[169] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[16] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[170] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[171] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[172] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[173] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[174] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[175] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[176] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[177] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[178] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[179] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[17] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[180] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[181] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[182] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[183] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[184] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[185] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[186] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[187] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[188] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[189] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[18] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[190] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[191] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[192] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[193] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[194] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[195] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[196] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[197] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[198] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[199] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[19] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[1] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[200] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[201] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[202] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[203] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[204] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[205] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[206] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[207] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[208] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[209] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[20] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[210] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[211] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[212] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[213] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[214] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[215] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[216] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[217] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[218] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[219] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[21] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[220] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[221] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[222] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[223] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[224] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[225] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[226] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[227] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[228] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[229] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[22] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[230] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[231] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[232] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[233] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[23] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[24] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[25] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[26] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[27] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[28] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[29] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[2] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[30] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[31] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[32] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[33] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[34] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[35] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[36] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[37] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[38] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[39] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[3] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[40] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[41] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[42] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[43] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[44] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[45] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[46] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[47] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[48] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[49] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[4] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[50] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[51] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[52] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[53] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[54] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[55] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[56] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[57] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[58] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[59] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[5] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[60] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[61] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[62] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[63] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[64] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[65] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[66] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[67] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[68] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[69] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[6] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[70] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[71] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[72] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[73] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[74] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[75] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[76] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[77] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[78] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[79] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[7] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[80] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[81] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[82] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[83] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[84] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[85] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[86] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[87] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[88] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[89] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[8] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[90] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[91] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[92] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[93] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[94] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[95] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[96] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[97] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[98] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[99] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[9] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[0] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[100] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[101] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[102] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[103] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[104] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[105] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[106] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[107] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[108] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[109] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[10] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[110] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[111] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[112] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[113] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[114] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[115] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[116] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[117] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[118] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[119] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[11] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[120] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[121] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[122] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[123] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[124] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[125] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[126] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[127] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[128] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[129] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[12] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[130] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[131] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[132] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[133] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[134] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[135] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[136] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[137] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[138] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[139] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[13] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[140] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[141] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[142] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[143] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[144] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[145] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[146] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[147] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[148] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[149] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[14] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[150] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[151] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[152] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[153] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[154] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[155] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[156] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[157] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[158] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[159] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[15] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[160] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[161] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[162] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[163] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[164] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[165] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[166] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[167] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[168] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[169] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[16] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[170] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[171] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[172] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[173] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[174] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[175] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[176] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[177] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[178] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[179] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[17] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[180] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[181] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[182] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[183] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[184] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[185] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[186] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[187] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[188] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[189] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[18] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[190] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[191] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[192] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[193] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[194] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[195] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[196] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[197] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[198] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[199] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[19] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[1] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[200] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[201] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[202] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[203] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[204] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[205] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[206] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[207] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[208] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[209] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[20] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[210] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[211] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[212] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[213] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[214] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[215] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[216] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[217] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[218] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[219] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[21] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[220] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[221] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[222] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[223] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[224] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[225] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[226] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[227] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[228] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[229] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[22] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[230] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[231] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[232] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[233] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[23] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[24] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[25] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[26] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[27] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[28] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[29] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[2] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[30] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[31] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[32] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[33] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[34] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[35] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[36] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[37] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[38] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[39] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[3] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[40] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[41] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[42] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[43] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[44] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[45] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[46] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[47] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[48] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[49] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[4] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[50] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[51] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[52] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[53] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[54] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[55] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[56] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[57] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[58] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[59] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[5] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[60] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[61] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[62] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[63] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[64] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[65] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[66] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[67] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[68] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[69] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[6] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[70] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[71] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[72] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[73] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[74] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[75] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[76] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[77] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[78] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[79] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[7] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[80] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[81] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[82] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[83] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[84] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[85] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[86] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[87] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[88] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[89] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[8] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[90] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[91] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[92] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[93] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[94] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[95] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[96] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[97] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[98] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[99] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[9] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[0] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[100] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[101] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[102] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[103] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[104] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[105] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[106] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[107] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[108] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[109] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[10] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[110] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[111] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[112] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[113] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[114] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[115] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[116] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[11] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[12] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[13] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[14] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[15] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[16] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[17] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[18] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[19] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[1] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[20] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[21] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[22] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[23] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[24] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[25] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[26] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[27] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[28] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[29] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[2] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[30] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[31] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[32] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[33] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[34] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[35] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[36] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[37] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[38] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[39] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[3] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[40] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[41] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[42] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[43] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[44] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[45] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[46] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[47] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[48] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[49] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[4] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[50] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[51] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[52] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[53] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[54] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[55] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[56] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[57] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[58] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[59] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[5] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[60] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[61] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[62] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[63] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[64] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[65] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[66] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[67] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[68] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[69] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[6] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[70] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[71] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[72] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[73] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[74] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[75] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[76] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[77] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[78] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[79] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[7] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[80] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[81] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[82] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[83] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[84] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[85] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[86] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[87] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[88] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[89] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[8] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[90] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[91] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[92] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[93] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[94] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[95] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[96] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[97] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[98] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[99] ;
 wire [0:0] \game_inst.snake_inst.shiftreg_inst.high[9] ;

 sg13g2_nand2_1 _0938_ (.Y(_0713_),
    .A(net531),
    .B(net119));
 sg13g2_nand3_1 _0939_ (.B(_0712_),
    .C(_0713_),
    .A(net131),
    .Y(_0105_));
 sg13g2_nand2_1 _0940_ (.Y(_0714_),
    .A(net503),
    .B(net119));
 sg13g2_and2_1 _0941_ (.A(\game_inst.head_x[2] ),
    .B(_0708_),
    .X(_0715_));
 sg13g2_xor2_1 _0942_ (.B(_0708_),
    .A(\game_inst.head_x[2] ),
    .X(_0716_));
 sg13g2_a21o_1 _0943_ (.A2(_0710_),
    .A1(\game_inst.head_x[0] ),
    .B1(_0709_),
    .X(_0717_));
 sg13g2_xor2_1 _0944_ (.B(_0717_),
    .A(_0716_),
    .X(_0718_));
 sg13g2_a22oi_1 _0945_ (.Y(_0719_),
    .B1(_0718_),
    .B2(_0495_),
    .A2(_0704_),
    .A1(net503));
 sg13g2_a21oi_1 _0946_ (.A1(_0714_),
    .A2(_0719_),
    .Y(_0106_),
    .B1(net151));
 sg13g2_a21oi_1 _0947_ (.A1(_0716_),
    .A2(_0717_),
    .Y(_0720_),
    .B1(_0715_));
 sg13g2_xnor2_1 _0948_ (.Y(_0721_),
    .A(\game_inst.head_x[3] ),
    .B(_0720_));
 sg13g2_xnor2_1 _0949_ (.Y(_0722_),
    .A(\game_inst.control_inst.dir[0] ),
    .B(_0721_));
 sg13g2_a22oi_1 _0950_ (.Y(_0723_),
    .B1(_0722_),
    .B2(_0495_),
    .A2(_0704_),
    .A1(net529));
 sg13g2_nand2_1 _0951_ (.Y(_0724_),
    .A(net529),
    .B(net119));
 sg13g2_nand3_1 _0952_ (.B(_0723_),
    .C(_0724_),
    .A(net131),
    .Y(_0107_));
 sg13g2_nand2_1 _0953_ (.Y(_0725_),
    .A(net497),
    .B(net119));
 sg13g2_and4_1 _0954_ (.A(_0237_),
    .B(net141),
    .C(_0240_),
    .D(_0720_),
    .X(_0726_));
 sg13g2_nor3_1 _0955_ (.A(_0237_),
    .B(_0708_),
    .C(_0720_),
    .Y(_0727_));
 sg13g2_o21ai_1 _0956_ (.B1(net497),
    .Y(_0728_),
    .A1(_0726_),
    .A2(_0727_));
 sg13g2_nor3_1 _0957_ (.A(net497),
    .B(_0726_),
    .C(_0727_),
    .Y(_0729_));
 sg13g2_nor2_1 _0958_ (.A(net119),
    .B(_0729_),
    .Y(_0730_));
 sg13g2_nand2_1 _0959_ (.Y(_0731_),
    .A(_0728_),
    .B(_0730_));
 sg13g2_a21oi_1 _0960_ (.A1(_0725_),
    .A2(_0731_),
    .Y(_0108_),
    .B1(net151));
 sg13g2_xnor2_1 _0961_ (.Y(_0732_),
    .A(net505),
    .B(net141));
 sg13g2_nand2_1 _0962_ (.Y(_0733_),
    .A(net505),
    .B(net121));
 sg13g2_a21oi_1 _0963_ (.A1(_0493_),
    .A2(_0732_),
    .Y(_0734_),
    .B1(net151));
 sg13g2_nand2_1 _0964_ (.Y(_0109_),
    .A(_0733_),
    .B(_0734_));
 sg13g2_nand2_1 _0965_ (.Y(_0735_),
    .A(_0239_),
    .B(\game_inst.control_inst.dir[0] ));
 sg13g2_and2_1 _0966_ (.A(\game_inst.head_y[1] ),
    .B(_0735_),
    .X(_0736_));
 sg13g2_xor2_1 _0967_ (.B(_0735_),
    .A(\game_inst.head_y[1] ),
    .X(_0737_));
 sg13g2_xor2_1 _0968_ (.B(_0737_),
    .A(net505),
    .X(_0738_));
 sg13g2_a22oi_1 _0969_ (.Y(_0739_),
    .B1(_0704_),
    .B2(_0738_),
    .A2(_0495_),
    .A1(net533));
 sg13g2_nand2_1 _0970_ (.Y(_0740_),
    .A(net533),
    .B(net121));
 sg13g2_nand3_1 _0971_ (.B(_0739_),
    .C(_0740_),
    .A(net131),
    .Y(_0110_));
 sg13g2_a21oi_1 _0972_ (.A1(\game_inst.head_y[0] ),
    .A2(_0737_),
    .Y(_0741_),
    .B1(_0736_));
 sg13g2_xnor2_1 _0973_ (.Y(_0742_),
    .A(\game_inst.head_y[2] ),
    .B(_0735_));
 sg13g2_xor2_1 _0974_ (.B(_0742_),
    .A(_0741_),
    .X(_0743_));
 sg13g2_a22oi_1 _0975_ (.Y(_0744_),
    .B1(_0704_),
    .B2(_0743_),
    .A2(_0495_),
    .A1(net528));
 sg13g2_nand2_1 _0976_ (.Y(_0745_),
    .A(net528),
    .B(net121));
 sg13g2_nand3_1 _0977_ (.B(_0744_),
    .C(_0745_),
    .A(net132),
    .Y(_0111_));
 sg13g2_nand2b_1 _0978_ (.Y(_0746_),
    .B(\game_inst.control_inst.dir[0] ),
    .A_N(\game_inst.head_y[0] ));
 sg13g2_a21oi_1 _0979_ (.A1(\game_inst.head_y[0] ),
    .A2(_0240_),
    .Y(_0747_),
    .B1(net141));
 sg13g2_nand3_1 _0980_ (.B(_0746_),
    .C(_0747_),
    .A(_0737_),
    .Y(_0748_));
 sg13g2_nor2_1 _0981_ (.A(_0742_),
    .B(_0748_),
    .Y(_0749_));
 sg13g2_o21ai_1 _0982_ (.B1(_0493_),
    .Y(_0750_),
    .A1(net567),
    .A2(_0749_));
 sg13g2_a21oi_1 _0983_ (.A1(net567),
    .A2(_0749_),
    .Y(_0751_),
    .B1(_0750_));
 sg13g2_nand2_1 _0984_ (.Y(_0752_),
    .A(net567),
    .B(net121));
 sg13g2_nor2b_1 _0985_ (.A(_0751_),
    .B_N(_0752_),
    .Y(_0753_));
 sg13g2_nor2_1 _0986_ (.A(net151),
    .B(_0753_),
    .Y(_0112_));
 sg13g2_nor2_1 _0987_ (.A(net153),
    .B(_0682_),
    .Y(_0113_));
 sg13g2_nand2_1 _0988_ (.Y(_0114_),
    .A(net133),
    .B(_0686_));
 sg13g2_nand2_2 _0989_ (.Y(_0754_),
    .A(_0270_),
    .B(_0499_));
 sg13g2_a22oi_1 _0990_ (.Y(_0755_),
    .B1(net117),
    .B2(_0703_),
    .A2(net118),
    .A1(net140));
 sg13g2_nor3_1 _0991_ (.A(_0705_),
    .B(_0706_),
    .C(_0755_),
    .Y(_0756_));
 sg13g2_xor2_1 _0992_ (.B(_0756_),
    .A(_0754_),
    .X(_0115_));
 sg13g2_nor2_1 _0993_ (.A(net138),
    .B(_0754_),
    .Y(_0757_));
 sg13g2_nand2_2 _0994_ (.Y(_0758_),
    .A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[0] [0]),
    .B(net134));
 sg13g2_nand3_1 _0995_ (.B(net138),
    .C(net134),
    .A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[0] [0]),
    .Y(_0759_));
 sg13g2_a21o_1 _0996_ (.A2(net134),
    .A1(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[0] [0]),
    .B1(net138),
    .X(_0760_));
 sg13g2_nand3_1 _0997_ (.B(_0759_),
    .C(_0760_),
    .A(net139),
    .Y(_0761_));
 sg13g2_a21o_1 _0998_ (.A2(_0760_),
    .A1(_0759_),
    .B1(net139),
    .X(_0762_));
 sg13g2_nand2_1 _0999_ (.Y(_0763_),
    .A(_0761_),
    .B(_0762_));
 sg13g2_a21oi_1 _1000_ (.A1(net134),
    .A2(_0763_),
    .Y(_0764_),
    .B1(net117));
 sg13g2_o21ai_1 _1001_ (.B1(_0712_),
    .Y(_0765_),
    .A1(net118),
    .A2(_0713_));
 sg13g2_nor2_1 _1002_ (.A(_0764_),
    .B(_0765_),
    .Y(_0766_));
 sg13g2_nor2_1 _1003_ (.A(_0757_),
    .B(_0766_),
    .Y(_0116_));
 sg13g2_and3_1 _1004_ (.X(_0767_),
    .A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[0] [0]),
    .B(net137),
    .C(net135));
 sg13g2_xor2_1 _1005_ (.B(_0758_),
    .A(net137),
    .X(_0768_));
 sg13g2_nand2_1 _1006_ (.Y(_0769_),
    .A(_0759_),
    .B(_0761_));
 sg13g2_a21oi_1 _1007_ (.A1(_0759_),
    .A2(_0761_),
    .Y(_0770_),
    .B1(_0768_));
 sg13g2_xor2_1 _1008_ (.B(_0769_),
    .A(_0768_),
    .X(_0771_));
 sg13g2_a22oi_1 _1009_ (.Y(_0772_),
    .B1(_0771_),
    .B2(net118),
    .A2(_0714_),
    .A1(net117));
 sg13g2_nand2b_1 _1010_ (.Y(_0773_),
    .B(_0719_),
    .A_N(_0772_));
 sg13g2_mux2_1 _1011_ (.A0(net137),
    .A1(_0773_),
    .S(_0754_),
    .X(_0117_));
 sg13g2_nor2_1 _1012_ (.A(net136),
    .B(_0754_),
    .Y(_0774_));
 sg13g2_o21ai_1 _1013_ (.B1(net136),
    .Y(_0775_),
    .A1(_0767_),
    .A2(_0770_));
 sg13g2_or3_1 _1014_ (.A(net136),
    .B(_0767_),
    .C(_0770_),
    .X(_0776_));
 sg13g2_nand2_1 _1015_ (.Y(_0777_),
    .A(_0775_),
    .B(_0776_));
 sg13g2_xnor2_1 _1016_ (.Y(_0778_),
    .A(_0758_),
    .B(_0777_));
 sg13g2_a22oi_1 _1017_ (.Y(_0779_),
    .B1(_0778_),
    .B2(net118),
    .A2(_0724_),
    .A1(net117));
 sg13g2_nor2b_1 _1018_ (.A(_0779_),
    .B_N(_0723_),
    .Y(_0780_));
 sg13g2_a21oi_1 _1019_ (.A1(_0754_),
    .A2(_0780_),
    .Y(_0118_),
    .B1(_0774_));
 sg13g2_mux2_1 _1020_ (.A0(_0776_),
    .A1(_0775_),
    .S(_0758_),
    .X(_0781_));
 sg13g2_xor2_1 _1021_ (.B(_0781_),
    .A(net516),
    .X(_0782_));
 sg13g2_a22oi_1 _1022_ (.Y(_0783_),
    .B1(_0782_),
    .B2(net118),
    .A2(_0725_),
    .A1(net117));
 sg13g2_a21oi_1 _1023_ (.A1(_0728_),
    .A2(_0730_),
    .Y(_0149_),
    .B1(_0783_));
 sg13g2_nor2_1 _1024_ (.A(net516),
    .B(_0754_),
    .Y(_0150_));
 sg13g2_a21oi_1 _1025_ (.A1(_0754_),
    .A2(_0149_),
    .Y(_0119_),
    .B1(_0150_));
 sg13g2_nand2_1 _1026_ (.Y(_0151_),
    .A(net435),
    .B(_0335_));
 sg13g2_a21oi_1 _1027_ (.A1(_0499_),
    .A2(_0151_),
    .Y(_0120_),
    .B1(net151));
 sg13g2_nand2_2 _1028_ (.Y(_0152_),
    .A(net134),
    .B(_0499_));
 sg13g2_inv_2 _1029_ (.Y(_0153_),
    .A(_0152_));
 sg13g2_a22oi_1 _1030_ (.Y(_0154_),
    .B1(_0500_),
    .B2(_0733_),
    .A2(_0498_),
    .A1(net578));
 sg13g2_a21oi_1 _1031_ (.A1(_0493_),
    .A2(_0732_),
    .Y(_0155_),
    .B1(_0154_));
 sg13g2_xnor2_1 _1032_ (.Y(_0121_),
    .A(_0153_),
    .B(_0155_));
 sg13g2_nor2_1 _1033_ (.A(net118),
    .B(_0740_),
    .Y(_0156_));
 sg13g2_nor2_2 _1034_ (.A(_0038_),
    .B(net134),
    .Y(_0157_));
 sg13g2_and2_1 _1035_ (.A(\game_inst.apple_inst.i_snake_y[1] ),
    .B(_0157_),
    .X(_0158_));
 sg13g2_xnor2_1 _1036_ (.Y(_0159_),
    .A(_0266_),
    .B(_0157_));
 sg13g2_xor2_1 _1037_ (.B(_0159_),
    .A(\game_inst.apple_inst.i_snake_y[0] ),
    .X(_0160_));
 sg13g2_a21oi_1 _1038_ (.A1(_0499_),
    .A2(_0160_),
    .Y(_0161_),
    .B1(_0156_));
 sg13g2_nand3_1 _1039_ (.B(_0152_),
    .C(_0161_),
    .A(_0739_),
    .Y(_0162_));
 sg13g2_o21ai_1 _1040_ (.B1(_0162_),
    .Y(_0163_),
    .A1(net521),
    .A2(_0152_));
 sg13g2_inv_1 _1041_ (.Y(_0122_),
    .A(net522));
 sg13g2_nand2_1 _1042_ (.Y(_0164_),
    .A(\game_inst.apple_inst.i_snake_y[2] ),
    .B(_0157_));
 sg13g2_xnor2_1 _1043_ (.Y(_0165_),
    .A(\game_inst.apple_inst.i_snake_y[2] ),
    .B(_0157_));
 sg13g2_a21oi_1 _1044_ (.A1(\game_inst.apple_inst.i_snake_y[0] ),
    .A2(_0159_),
    .Y(_0166_),
    .B1(_0158_));
 sg13g2_xnor2_1 _1045_ (.Y(_0167_),
    .A(_0165_),
    .B(_0166_));
 sg13g2_a22oi_1 _1046_ (.Y(_0168_),
    .B1(_0167_),
    .B2(net118),
    .A2(_0745_),
    .A1(net117));
 sg13g2_nand2b_1 _1047_ (.Y(_0169_),
    .B(_0744_),
    .A_N(_0168_));
 sg13g2_mux2_1 _1048_ (.A0(net526),
    .A1(_0169_),
    .S(_0152_),
    .X(_0123_));
 sg13g2_o21ai_1 _1049_ (.B1(_0164_),
    .Y(_0170_),
    .A1(_0165_),
    .A2(_0166_));
 sg13g2_xnor2_1 _1050_ (.Y(_0171_),
    .A(_0268_),
    .B(_0157_));
 sg13g2_xnor2_1 _1051_ (.Y(_0172_),
    .A(_0170_),
    .B(_0171_));
 sg13g2_a22oi_1 _1052_ (.Y(_0173_),
    .B1(_0172_),
    .B2(net118),
    .A2(_0752_),
    .A1(net117));
 sg13g2_nor3_1 _1053_ (.A(_0751_),
    .B(_0153_),
    .C(_0173_),
    .Y(_0174_));
 sg13g2_a21oi_1 _1054_ (.A1(_0268_),
    .A2(_0153_),
    .Y(_0124_),
    .B1(_0174_));
 sg13g2_nor2_1 _1055_ (.A(net518),
    .B(_0582_),
    .Y(_0175_));
 sg13g2_and4_1 _1056_ (.A(net419),
    .B(net518),
    .C(_0340_),
    .D(_0580_),
    .X(_0176_));
 sg13g2_o21ai_1 _1057_ (.B1(net132),
    .Y(_0125_),
    .A1(_0175_),
    .A2(_0176_));
 sg13g2_nor2_1 _1058_ (.A(net480),
    .B(_0176_),
    .Y(_0177_));
 sg13g2_and2_1 _1059_ (.A(net480),
    .B(_0176_),
    .X(_0178_));
 sg13g2_nor3_1 _1060_ (.A(net150),
    .B(net481),
    .C(_0178_),
    .Y(_0126_));
 sg13g2_nor2_1 _1061_ (.A(net495),
    .B(_0178_),
    .Y(_0179_));
 sg13g2_and4_1 _1062_ (.A(\game_inst.snake_inst.length[0] ),
    .B(net480),
    .C(net495),
    .D(_0582_),
    .X(_0180_));
 sg13g2_nand3_1 _1063_ (.B(\game_inst.snake_inst.length[2] ),
    .C(_0176_),
    .A(\game_inst.snake_inst.length[1] ),
    .Y(_0181_));
 sg13g2_nor3_1 _1064_ (.A(net150),
    .B(_0179_),
    .C(_0180_),
    .Y(_0127_));
 sg13g2_nor2_1 _1065_ (.A(net465),
    .B(_0180_),
    .Y(_0182_));
 sg13g2_nor2_1 _1066_ (.A(_0254_),
    .B(_0181_),
    .Y(_0183_));
 sg13g2_nor3_1 _1067_ (.A(net151),
    .B(net466),
    .C(_0183_),
    .Y(_0128_));
 sg13g2_nor2_1 _1068_ (.A(net450),
    .B(_0183_),
    .Y(_0184_));
 sg13g2_and3_2 _1069_ (.X(_0185_),
    .A(net465),
    .B(net450),
    .C(_0180_));
 sg13g2_nor3_1 _1070_ (.A(net150),
    .B(net451),
    .C(_0185_),
    .Y(_0129_));
 sg13g2_xnor2_1 _1071_ (.Y(_0186_),
    .A(net498),
    .B(_0185_));
 sg13g2_nor2_1 _1072_ (.A(net150),
    .B(_0186_),
    .Y(_0130_));
 sg13g2_a21oi_1 _1073_ (.A1(\game_inst.snake_inst.length[5] ),
    .A2(_0185_),
    .Y(_0187_),
    .B1(net410));
 sg13g2_and3_1 _1074_ (.X(_0188_),
    .A(\game_inst.snake_inst.length[5] ),
    .B(net410),
    .C(_0185_));
 sg13g2_nor3_1 _1075_ (.A(net150),
    .B(net411),
    .C(_0188_),
    .Y(_0131_));
 sg13g2_o21ai_1 _1076_ (.B1(net132),
    .Y(_0189_),
    .A1(net349),
    .A2(_0188_));
 sg13g2_a21oi_1 _1077_ (.A1(net349),
    .A2(_0188_),
    .Y(_0132_),
    .B1(_0189_));
 sg13g2_nand2_1 _1078_ (.Y(_0190_),
    .A(net131),
    .B(_0499_));
 sg13g2_nor3_1 _1079_ (.A(_0338_),
    .B(_0501_),
    .C(_0190_),
    .Y(_0133_));
 sg13g2_nor2_1 _1080_ (.A(net460),
    .B(_0501_),
    .Y(_0191_));
 sg13g2_nor3_1 _1081_ (.A(_0502_),
    .B(_0190_),
    .C(net461),
    .Y(_0134_));
 sg13g2_a21oi_1 _1082_ (.A1(\game_inst.snake_inst.pos[3] ),
    .A2(_0502_),
    .Y(_0192_),
    .B1(net393));
 sg13g2_nor3_1 _1083_ (.A(_0504_),
    .B(_0190_),
    .C(net394),
    .Y(_0135_));
 sg13g2_nand2_1 _1084_ (.Y(_0193_),
    .A(net378),
    .B(_0662_));
 sg13g2_o21ai_1 _1085_ (.B1(net379),
    .Y(_0136_),
    .A1(_0243_),
    .A2(net112));
 sg13g2_nor2_1 _1086_ (.A(net388),
    .B(net112),
    .Y(_0194_));
 sg13g2_a21oi_1 _1087_ (.A1(_0267_),
    .A2(net110),
    .Y(_0137_),
    .B1(_0194_));
 sg13g2_mux2_1 _1088_ (.A0(net415),
    .A1(net457),
    .S(_0662_),
    .X(_0138_));
 sg13g2_nand2_1 _1089_ (.Y(_0195_),
    .A(net408),
    .B(net110));
 sg13g2_o21ai_1 _1090_ (.B1(_0195_),
    .Y(_0139_),
    .A1(_0241_),
    .A2(net112));
 sg13g2_nor3_1 _1091_ (.A(_0239_),
    .B(\game_inst.control_inst.dir[0] ),
    .C(net463),
    .Y(_0196_));
 sg13g2_nor2_1 _1092_ (.A(net152),
    .B(net464),
    .Y(_0140_));
 sg13g2_nand3b_1 _1093_ (.B(_0003_),
    .C(net153),
    .Y(_0197_),
    .A_N(\game_inst.tickgen_inst.prev_user_input ));
 sg13g2_a21oi_1 _1094_ (.A1(net399),
    .A2(_0197_),
    .Y(_0198_),
    .B1(net154));
 sg13g2_o21ai_1 _1095_ (.B1(_0198_),
    .Y(_0141_),
    .A1(net399),
    .A2(_0197_));
 sg13g2_nor2b_1 _1096_ (.A(net1),
    .B_N(net487),
    .Y(_0199_));
 sg13g2_xnor2_1 _1097_ (.Y(_0200_),
    .A(net487),
    .B(net1));
 sg13g2_a21oi_1 _1098_ (.A1(net399),
    .A2(_0200_),
    .Y(_0201_),
    .B1(_0197_));
 sg13g2_o21ai_1 _1099_ (.B1(_0201_),
    .Y(_0202_),
    .A1(net399),
    .A2(_0200_));
 sg13g2_a21oi_1 _1100_ (.A1(net487),
    .A2(_0197_),
    .Y(_0203_),
    .B1(net155));
 sg13g2_nand2_1 _1101_ (.Y(_0142_),
    .A(_0202_),
    .B(net488));
 sg13g2_a21oi_1 _1102_ (.A1(net399),
    .A2(_0200_),
    .Y(_0204_),
    .B1(_0199_));
 sg13g2_xor2_1 _1103_ (.B(net1),
    .A(net511),
    .X(_0205_));
 sg13g2_a21oi_1 _1104_ (.A1(_0204_),
    .A2(_0205_),
    .Y(_0206_),
    .B1(_0197_));
 sg13g2_o21ai_1 _1105_ (.B1(_0206_),
    .Y(_0207_),
    .A1(_0204_),
    .A2(_0205_));
 sg13g2_a21oi_1 _1106_ (.A1(net511),
    .A2(_0197_),
    .Y(_0208_),
    .B1(net155));
 sg13g2_nand2_1 _1107_ (.Y(_0143_),
    .A(_0207_),
    .B(net512));
 sg13g2_nor2_1 _1108_ (.A(net5),
    .B(net346),
    .Y(_0209_));
 sg13g2_nand3_1 _1109_ (.B(\game_inst.sound_inst.vsync_pulse ),
    .C(_0209_),
    .A(net463),
    .Y(_0210_));
 sg13g2_nor2_1 _1110_ (.A(\game_inst.o_success ),
    .B(_0210_),
    .Y(_0211_));
 sg13g2_or2_1 _1111_ (.X(_0212_),
    .B(_0210_),
    .A(\game_inst.o_success ));
 sg13g2_a21oi_1 _1112_ (.A1(_0231_),
    .A2(\game_inst.tickgen_inst.counter_max[3] ),
    .Y(_0213_),
    .B1(net357));
 sg13g2_xnor2_1 _1113_ (.Y(_0214_),
    .A(net386),
    .B(\game_inst.tickgen_inst.counter_max[2] ));
 sg13g2_nand2b_1 _1114_ (.Y(_0215_),
    .B(net399),
    .A_N(\game_inst.tickgen_inst.counter[1] ));
 sg13g2_a22oi_1 _1115_ (.Y(_0216_),
    .B1(_0233_),
    .B2(\game_inst.tickgen_inst.counter[1] ),
    .A2(_0232_),
    .A1(net344));
 sg13g2_nand4_1 _1116_ (.B(_0214_),
    .C(_0215_),
    .A(_0213_),
    .Y(_0217_),
    .D(_0216_));
 sg13g2_or2_1 _1117_ (.X(_0218_),
    .B(_0217_),
    .A(_0212_));
 sg13g2_o21ai_1 _1118_ (.B1(net401),
    .Y(_0219_),
    .A1(_0540_),
    .A2(_0211_));
 sg13g2_a21oi_1 _1119_ (.A1(_0218_),
    .A2(net402),
    .Y(_0144_),
    .B1(net153));
 sg13g2_and2_1 _1120_ (.A(_0211_),
    .B(_0217_),
    .X(_0220_));
 sg13g2_o21ai_1 _1121_ (.B1(net133),
    .Y(_0221_),
    .A1(net357),
    .A2(_0220_));
 sg13g2_a21oi_1 _1122_ (.A1(net357),
    .A2(_0211_),
    .Y(_0145_),
    .B1(_0221_));
 sg13g2_and2_1 _1123_ (.A(\game_inst.tickgen_inst.counter[1] ),
    .B(net357),
    .X(_0222_));
 sg13g2_nand2_1 _1124_ (.Y(_0223_),
    .A(net499),
    .B(net357));
 sg13g2_a22oi_1 _1125_ (.Y(_0224_),
    .B1(_0220_),
    .B2(_0223_),
    .A2(_0212_),
    .A1(net499));
 sg13g2_o21ai_1 _1126_ (.B1(net133),
    .Y(_0225_),
    .A1(net499),
    .A2(net357));
 sg13g2_nor2_1 _1127_ (.A(_0224_),
    .B(_0225_),
    .Y(_0146_));
 sg13g2_a21oi_1 _1128_ (.A1(_0220_),
    .A2(_0222_),
    .Y(_0226_),
    .B1(net386));
 sg13g2_nand2_1 _1129_ (.Y(_0227_),
    .A(net386),
    .B(_0222_));
 sg13g2_a21oi_1 _1130_ (.A1(_0217_),
    .A2(_0227_),
    .Y(_0228_),
    .B1(_0212_));
 sg13g2_nor3_1 _1131_ (.A(net152),
    .B(net387),
    .C(_0228_),
    .Y(_0147_));
 sg13g2_o21ai_1 _1132_ (.B1(_0231_),
    .Y(_0229_),
    .A1(_0212_),
    .A2(_0227_));
 sg13g2_nand2_1 _1133_ (.Y(_0230_),
    .A(net133),
    .B(_0229_));
 sg13g2_a21oi_1 _1134_ (.A1(net344),
    .A2(_0228_),
    .Y(_0148_),
    .B1(_0230_));
 sg13g2_buf_1 _1135_ (.A(\game_inst.vga_inst.color[3] ),
    .X(uo_out[6]));
 sg13g2_inv_1 _1136_ (.Y(_0231_),
    .A(net344));
 sg13g2_inv_1 _1137_ (.Y(_0232_),
    .A(\game_inst.tickgen_inst.counter_max[3] ));
 sg13g2_inv_1 _1138_ (.Y(_0233_),
    .A(net399));
 sg13g2_inv_1 _1139_ (.Y(_0234_),
    .A(\game_inst.apple_inst.i_snake_valid ));
 sg13g2_inv_1 _1140_ (.Y(_0235_),
    .A(\game_inst.head_y[2] ));
 sg13g2_inv_1 _1141_ (.Y(_0236_),
    .A(\game_inst.head_y[0] ));
 sg13g2_inv_1 _1142_ (.Y(_0237_),
    .A(\game_inst.head_x[3] ));
 sg13g2_inv_2 _1143_ (.Y(_0238_),
    .A(net500));
 sg13g2_inv_2 _1144_ (.Y(_0239_),
    .A(net581));
 sg13g2_inv_4 _1145_ (.A(\game_inst.control_inst.dir[0] ),
    .Y(_0240_));
 sg13g2_inv_1 _1146_ (.Y(_0241_),
    .A(net458));
 sg13g2_inv_1 _1147_ (.Y(_0242_),
    .A(net388));
 sg13g2_inv_1 _1148_ (.Y(_0243_),
    .A(net375));
 sg13g2_inv_1 _1149_ (.Y(_0244_),
    .A(net397));
 sg13g2_inv_1 _1150_ (.Y(_0245_),
    .A(net417));
 sg13g2_inv_1 _1151_ (.Y(_0246_),
    .A(net416));
 sg13g2_inv_1 _1152_ (.Y(_0247_),
    .A(net406));
 sg13g2_inv_1 _1153_ (.Y(_0248_),
    .A(\game_inst.vga_inst.py[7] ));
 sg13g2_inv_1 _1154_ (.Y(_0249_),
    .A(\game_inst.sound_inst.phase[0] ));
 sg13g2_inv_1 _1155_ (.Y(_0250_),
    .A(\game_inst.sound_inst.max_counter[0] ));
 sg13g2_inv_1 _1156_ (.Y(_0251_),
    .A(\game_inst.sound_inst.counter[1] ));
 sg13g2_inv_1 _1157_ (.Y(_0252_),
    .A(\game_inst.sound_inst.max_counter[2] ));
 sg13g2_inv_1 _1158_ (.Y(_0038_),
    .A(net459));
 sg13g2_inv_1 _1159_ (.Y(_0253_),
    .A(net346));
 sg13g2_inv_1 _1160_ (.Y(_0254_),
    .A(net465));
 sg13g2_inv_1 _1161_ (.Y(_0255_),
    .A(\game_inst.snake_inst.length[4] ));
 sg13g2_inv_1 _1162_ (.Y(_0256_),
    .A(\game_inst.o_tick ));
 sg13g2_inv_1 _1163_ (.Y(_0257_),
    .A(\game_inst.snake_inst.pos[0] ));
 sg13g2_inv_1 _1164_ (.Y(_0258_),
    .A(\game_inst.snake_inst.pos[4] ));
 sg13g2_inv_1 _1165_ (.Y(_0259_),
    .A(\game_inst.apple_inst.apple_x[0] ));
 sg13g2_inv_1 _1166_ (.Y(_0260_),
    .A(net140));
 sg13g2_inv_1 _1167_ (.Y(_0261_),
    .A(net138));
 sg13g2_inv_1 _1168_ (.Y(_0262_),
    .A(\game_inst.apple_inst.apple_x[1] ));
 sg13g2_inv_1 _1169_ (.Y(_0263_),
    .A(\game_inst.apple_inst.i_snake_x[4] ));
 sg13g2_inv_2 _1170_ (.Y(_0264_),
    .A(\game_inst.apple_inst.apple_x[4] ));
 sg13g2_inv_1 _1171_ (.Y(_0265_),
    .A(\game_inst.apple_inst.apple_y[0] ));
 sg13g2_inv_1 _1172_ (.Y(_0266_),
    .A(\game_inst.apple_inst.i_snake_y[1] ));
 sg13g2_inv_1 _1173_ (.Y(_0267_),
    .A(\game_inst.apple_inst.apple_y[1] ));
 sg13g2_inv_1 _1174_ (.Y(_0268_),
    .A(net514));
 sg13g2_inv_1 _1175_ (.Y(_0269_),
    .A(net156));
 sg13g2_inv_2 _1176_ (.Y(_0270_),
    .A(net134));
 sg13g2_inv_1 _1177_ (.Y(_0271_),
    .A(net145));
 sg13g2_inv_2 _1178_ (.Y(_0272_),
    .A(net147));
 sg13g2_nor2b_2 _1179_ (.A(net342),
    .B_N(net340),
    .Y(\game_inst.sound_inst.vsync_pulse ));
 sg13g2_nand4_1 _1180_ (.B(\game_inst.snake_inst.length[5] ),
    .C(\game_inst.snake_inst.length[6] ),
    .A(_0255_),
    .Y(_0273_),
    .D(\game_inst.snake_inst.length[7] ));
 sg13g2_nand2b_1 _1181_ (.Y(_0274_),
    .B(\game_inst.snake_inst.length[0] ),
    .A_N(\game_inst.snake_inst.length[1] ));
 sg13g2_nor4_2 _1182_ (.A(\game_inst.snake_inst.length[2] ),
    .B(_0254_),
    .C(_0273_),
    .Y(\game_inst.o_success ),
    .D(_0274_));
 sg13g2_or2_1 _1183_ (.X(_0003_),
    .B(net1),
    .A(net2));
 sg13g2_or3_1 _1184_ (.A(\game_inst.vga_inst.py[8] ),
    .B(\game_inst.vga_inst.py[7] ),
    .C(net142),
    .X(_0275_));
 sg13g2_nand3_1 _1185_ (.B(\game_inst.vga_inst.py[7] ),
    .C(net142),
    .A(\game_inst.vga_inst.py[8] ),
    .Y(_0276_));
 sg13g2_a21oi_1 _1186_ (.A1(_0275_),
    .A2(_0276_),
    .Y(_0277_),
    .B1(net484));
 sg13g2_nor2_1 _1187_ (.A(net148),
    .B(\game_inst.vga_inst.px[6] ),
    .Y(_0278_));
 sg13g2_or2_1 _1188_ (.X(_0279_),
    .B(\game_inst.vga_inst.px[6] ),
    .A(net148));
 sg13g2_nor2_1 _1189_ (.A(net146),
    .B(net147),
    .Y(_0280_));
 sg13g2_nand2_2 _1190_ (.Y(_0281_),
    .A(net148),
    .B(net475));
 sg13g2_o21ai_1 _1191_ (.B1(_0280_),
    .Y(_0282_),
    .A1(net144),
    .A2(_0278_));
 sg13g2_a21oi_1 _1192_ (.A1(net144),
    .A2(_0281_),
    .Y(_0283_),
    .B1(_0282_));
 sg13g2_nor2_1 _1193_ (.A(_0277_),
    .B(_0283_),
    .Y(_0284_));
 sg13g2_nand4_1 _1194_ (.B(\game_inst.vga_inst.py[7] ),
    .C(net142),
    .A(\game_inst.vga_inst.py[8] ),
    .Y(_0285_),
    .D(\game_inst.vga_inst.py[5] ));
 sg13g2_o21ai_1 _1195_ (.B1(net144),
    .Y(_0286_),
    .A1(net146),
    .A2(net147));
 sg13g2_nand3b_1 _1196_ (.B(_0285_),
    .C(_0286_),
    .Y(_0287_),
    .A_N(net353));
 sg13g2_or3_1 _1197_ (.A(_0253_),
    .B(_0284_),
    .C(_0287_),
    .X(_0288_));
 sg13g2_or3_1 _1198_ (.A(_0277_),
    .B(_0283_),
    .C(_0287_),
    .X(_0289_));
 sg13g2_nand3_1 _1199_ (.B(net143),
    .C(net453),
    .A(net351),
    .Y(_0290_));
 sg13g2_or2_1 _1200_ (.X(_0291_),
    .B(\game_inst.vga_inst.py[2] ),
    .A(net351));
 sg13g2_o21ai_1 _1201_ (.B1(_0290_),
    .Y(_0292_),
    .A1(net143),
    .A2(_0291_));
 sg13g2_and2_1 _1202_ (.A(net149),
    .B(net548),
    .X(_0293_));
 sg13g2_nor3_1 _1203_ (.A(net149),
    .B(net517),
    .C(net383),
    .Y(_0294_));
 sg13g2_a21oi_1 _1204_ (.A1(net383),
    .A2(_0293_),
    .Y(_0295_),
    .B1(_0294_));
 sg13g2_nand2b_1 _1205_ (.Y(_0296_),
    .B(net569),
    .A_N(net142));
 sg13g2_a22oi_1 _1206_ (.Y(_0297_),
    .B1(_0267_),
    .B2(net142),
    .A2(_0265_),
    .A1(\game_inst.vga_inst.py[5] ));
 sg13g2_xnor2_1 _1207_ (.Y(_0298_),
    .A(net446),
    .B(net145));
 sg13g2_nand2b_1 _1208_ (.Y(_0299_),
    .B(\game_inst.vga_inst.py[7] ),
    .A_N(net457));
 sg13g2_xnor2_1 _1209_ (.Y(_0300_),
    .A(net437),
    .B(net475));
 sg13g2_xnor2_1 _1210_ (.Y(_0301_),
    .A(\game_inst.apple_inst.apple_x[0] ),
    .B(net148));
 sg13g2_nor4_1 _1211_ (.A(net455),
    .B(net439),
    .C(net444),
    .D(net447),
    .Y(_0302_));
 sg13g2_nand2b_1 _1212_ (.Y(_0303_),
    .B(net378),
    .A_N(net484));
 sg13g2_xnor2_1 _1213_ (.Y(_0304_),
    .A(\game_inst.vga_inst.py[8] ),
    .B(net408));
 sg13g2_nand4_1 _1214_ (.B(_0299_),
    .C(_0301_),
    .A(net419),
    .Y(_0305_),
    .D(_0304_));
 sg13g2_nand2b_1 _1215_ (.Y(_0306_),
    .B(net147),
    .A_N(\game_inst.apple_inst.apple_x[2] ));
 sg13g2_nand3_1 _1216_ (.B(_0297_),
    .C(_0306_),
    .A(_0296_),
    .Y(_0307_));
 sg13g2_a22oi_1 _1217_ (.Y(_0308_),
    .B1(_0272_),
    .B2(net425),
    .A2(net457),
    .A1(_0248_));
 sg13g2_xnor2_1 _1218_ (.Y(_0309_),
    .A(\game_inst.apple_inst.apple_x[4] ),
    .B(net144));
 sg13g2_nand4_1 _1219_ (.B(_0302_),
    .C(_0308_),
    .A(_0298_),
    .Y(_0310_),
    .D(_0309_));
 sg13g2_nor4_1 _1220_ (.A(_0292_),
    .B(_0305_),
    .C(net570),
    .D(_0310_),
    .Y(_0311_));
 sg13g2_nand4_1 _1221_ (.B(_0300_),
    .C(_0303_),
    .A(_0295_),
    .Y(_0312_),
    .D(net571));
 sg13g2_o21ai_1 _1222_ (.B1(_0288_),
    .Y(_0000_),
    .A1(_0289_),
    .A2(_0312_));
 sg13g2_nor3_1 _1223_ (.A(net346),
    .B(_0284_),
    .C(_0287_),
    .Y(_0002_));
 sg13g2_mux2_1 _1224_ (.A0(net447),
    .A1(net444),
    .S(net149),
    .X(_0313_));
 sg13g2_nand2b_1 _1225_ (.Y(_0314_),
    .B(_0313_),
    .A_N(_0292_));
 sg13g2_nor3_1 _1226_ (.A(net143),
    .B(net439),
    .C(_0291_),
    .Y(_0315_));
 sg13g2_o21ai_1 _1227_ (.B1(_0290_),
    .Y(_0316_),
    .A1(_0302_),
    .A2(_0315_));
 sg13g2_o21ai_1 _1228_ (.B1(_0295_),
    .Y(_0317_),
    .A1(net455),
    .A2(_0290_));
 sg13g2_nand2b_1 _1229_ (.Y(_0318_),
    .B(_0316_),
    .A_N(_0317_));
 sg13g2_a21oi_1 _1230_ (.A1(_0314_),
    .A2(_0318_),
    .Y(_0001_),
    .B1(_0289_));
 sg13g2_nand2_1 _1231_ (.Y(_0319_),
    .A(net143),
    .B(\game_inst.vga_inst.py[1] ));
 sg13g2_nor4_1 _1232_ (.A(net353),
    .B(_0285_),
    .C(_0291_),
    .D(_0319_),
    .Y(_0037_));
 sg13g2_mux2_1 _1233_ (.A0(_0279_),
    .A1(_0281_),
    .S(net149),
    .X(_0320_));
 sg13g2_and4_1 _1234_ (.A(net144),
    .B(_0271_),
    .C(net473),
    .D(_0320_),
    .X(_0036_));
 sg13g2_nor2b_1 _1235_ (.A(\game_inst.apple_inst.o_ready ),
    .B_N(\game_inst.control_inst.o_start ),
    .Y(eat));
 sg13g2_and3_2 _1236_ (.X(_0321_),
    .A(net343),
    .B(net436),
    .C(net383));
 sg13g2_and2_1 _1237_ (.A(net517),
    .B(_0321_),
    .X(_0322_));
 sg13g2_and2_1 _1238_ (.A(_0293_),
    .B(_0321_),
    .X(_0323_));
 sg13g2_nand2_2 _1239_ (.Y(_0324_),
    .A(_0293_),
    .B(_0321_));
 sg13g2_xor2_1 _1240_ (.B(\game_inst.snake_inst.pos[7] ),
    .A(\game_inst.snake_inst.length[7] ),
    .X(_0325_));
 sg13g2_xor2_1 _1241_ (.B(\game_inst.snake_inst.pos[1] ),
    .A(\game_inst.snake_inst.length[1] ),
    .X(_0326_));
 sg13g2_xor2_1 _1242_ (.B(\game_inst.snake_inst.pos[0] ),
    .A(\game_inst.snake_inst.length[0] ),
    .X(_0327_));
 sg13g2_xor2_1 _1243_ (.B(\game_inst.snake_inst.pos[5] ),
    .A(\game_inst.snake_inst.length[5] ),
    .X(_0328_));
 sg13g2_xor2_1 _1244_ (.B(\game_inst.snake_inst.pos[4] ),
    .A(\game_inst.snake_inst.length[4] ),
    .X(_0329_));
 sg13g2_xor2_1 _1245_ (.B(\game_inst.snake_inst.pos[6] ),
    .A(\game_inst.snake_inst.length[6] ),
    .X(_0330_));
 sg13g2_xnor2_1 _1246_ (.Y(_0331_),
    .A(\game_inst.snake_inst.length[3] ),
    .B(\game_inst.snake_inst.pos[3] ));
 sg13g2_xor2_1 _1247_ (.B(\game_inst.snake_inst.pos[2] ),
    .A(\game_inst.snake_inst.length[2] ),
    .X(_0332_));
 sg13g2_nor3_1 _1248_ (.A(_0325_),
    .B(_0327_),
    .C(_0329_),
    .Y(_0333_));
 sg13g2_nor4_1 _1249_ (.A(_0326_),
    .B(_0328_),
    .C(_0330_),
    .D(_0332_),
    .Y(_0334_));
 sg13g2_nand3_1 _1250_ (.B(_0333_),
    .C(_0334_),
    .A(_0331_),
    .Y(_0335_));
 sg13g2_nand2_1 _1251_ (.Y(_0336_),
    .A(_0038_),
    .B(_0335_));
 sg13g2_nor4_1 _1252_ (.A(\game_inst.snake_inst.pos[2] ),
    .B(\game_inst.snake_inst.pos[5] ),
    .C(net393),
    .D(\game_inst.snake_inst.pos[6] ),
    .Y(_0337_));
 sg13g2_nor2_1 _1253_ (.A(net534),
    .B(net359),
    .Y(_0338_));
 sg13g2_nor2_1 _1254_ (.A(net428),
    .B(\game_inst.snake_inst.pos[3] ),
    .Y(_0339_));
 sg13g2_and3_2 _1255_ (.X(_0340_),
    .A(_0337_),
    .B(_0338_),
    .C(_0339_));
 sg13g2_nand3_1 _1256_ (.B(_0338_),
    .C(_0339_),
    .A(_0337_),
    .Y(_0341_));
 sg13g2_nor2_1 _1257_ (.A(\game_inst.vga_inst.prev_dir[0] ),
    .B(_0340_),
    .Y(_0342_));
 sg13g2_nand2b_1 _1258_ (.Y(_0343_),
    .B(_0342_),
    .A_N(\game_inst.vga_inst.prev_dir[1] ));
 sg13g2_o21ai_1 _1259_ (.B1(_0343_),
    .Y(_0344_),
    .A1(net135),
    .A2(_0336_));
 sg13g2_nor2b_1 _1260_ (.A(net147),
    .B_N(net137),
    .Y(_0345_));
 sg13g2_nor2b_1 _1261_ (.A(\game_inst.vga_inst.px[6] ),
    .B_N(net138),
    .Y(_0346_));
 sg13g2_nand2b_2 _1262_ (.Y(_0347_),
    .B(net148),
    .A_N(net139));
 sg13g2_nand2b_2 _1263_ (.Y(_0348_),
    .B(\game_inst.vga_inst.px[6] ),
    .A_N(net138));
 sg13g2_nor2b_2 _1264_ (.A(_0346_),
    .B_N(_0348_),
    .Y(_0349_));
 sg13g2_a21o_2 _1265_ (.A2(_0348_),
    .A1(_0347_),
    .B1(_0346_),
    .X(_0350_));
 sg13g2_xnor2_1 _1266_ (.Y(_0351_),
    .A(net137),
    .B(net147));
 sg13g2_a21oi_2 _1267_ (.B1(_0345_),
    .Y(_0352_),
    .A2(_0351_),
    .A1(_0350_));
 sg13g2_nor2b_1 _1268_ (.A(net145),
    .B_N(net136),
    .Y(_0353_));
 sg13g2_xnor2_1 _1269_ (.Y(_0354_),
    .A(net136),
    .B(net145));
 sg13g2_inv_1 _1270_ (.Y(_0355_),
    .A(_0354_));
 sg13g2_xnor2_1 _1271_ (.Y(_0356_),
    .A(_0352_),
    .B(_0354_));
 sg13g2_xnor2_1 _1272_ (.Y(_0357_),
    .A(_0352_),
    .B(_0355_));
 sg13g2_nand2_2 _1273_ (.Y(_0358_),
    .A(net420),
    .B(net377));
 sg13g2_nand3_1 _1274_ (.B(net420),
    .C(net377),
    .A(net453),
    .Y(_0359_));
 sg13g2_and4_1 _1275_ (.A(net143),
    .B(\game_inst.vga_inst.py[2] ),
    .C(\game_inst.vga_inst.py[1] ),
    .D(\game_inst.vga_inst.py[0] ),
    .X(_0360_));
 sg13g2_and2_1 _1276_ (.A(\game_inst.vga_inst.py[5] ),
    .B(\game_inst.vga_inst.py[4] ),
    .X(_0361_));
 sg13g2_and4_1 _1277_ (.A(\game_inst.vga_inst.py[7] ),
    .B(net142),
    .C(_0360_),
    .D(_0361_),
    .X(_0362_));
 sg13g2_xnor2_1 _1278_ (.Y(_0363_),
    .A(\game_inst.vga_inst.py[8] ),
    .B(\game_inst.apple_inst.i_snake_y[3] ));
 sg13g2_xnor2_1 _1279_ (.Y(_0364_),
    .A(_0362_),
    .B(_0363_));
 sg13g2_xnor2_1 _1280_ (.Y(_0365_),
    .A(net142),
    .B(\game_inst.apple_inst.i_snake_y[1] ));
 sg13g2_xnor2_1 _1281_ (.Y(_0366_),
    .A(\game_inst.vga_inst.py[7] ),
    .B(\game_inst.apple_inst.i_snake_y[2] ));
 sg13g2_nor2_1 _1282_ (.A(_0290_),
    .B(_0358_),
    .Y(_0367_));
 sg13g2_xnor2_1 _1283_ (.Y(_0368_),
    .A(\game_inst.vga_inst.py[5] ),
    .B(\game_inst.apple_inst.i_snake_y[0] ));
 sg13g2_xnor2_1 _1284_ (.Y(_0369_),
    .A(_0367_),
    .B(_0368_));
 sg13g2_nand2b_1 _1285_ (.Y(_0370_),
    .B(net144),
    .A_N(\game_inst.apple_inst.i_snake_x[4] ));
 sg13g2_nor2_1 _1286_ (.A(_0353_),
    .B(_0370_),
    .Y(_0371_));
 sg13g2_nand3_1 _1287_ (.B(_0360_),
    .C(_0361_),
    .A(net142),
    .Y(_0372_));
 sg13g2_xor2_1 _1288_ (.B(_0372_),
    .A(_0366_),
    .X(_0373_));
 sg13g2_nand3_1 _1289_ (.B(_0361_),
    .C(_0365_),
    .A(_0360_),
    .Y(_0374_));
 sg13g2_a21oi_1 _1290_ (.A1(_0360_),
    .A2(_0361_),
    .Y(_0375_),
    .B1(_0365_));
 sg13g2_nand3b_1 _1291_ (.B(_0371_),
    .C(_0374_),
    .Y(_0376_),
    .A_N(_0375_));
 sg13g2_nor4_2 _1292_ (.A(_0364_),
    .B(_0369_),
    .C(_0373_),
    .Y(_0377_),
    .D(_0376_));
 sg13g2_and2_1 _1293_ (.A(_0356_),
    .B(_0377_),
    .X(_0378_));
 sg13g2_nand3_1 _1294_ (.B(_0356_),
    .C(_0377_),
    .A(\game_inst.apple_inst.i_snake_valid ),
    .Y(_0379_));
 sg13g2_nor2b_1 _1295_ (.A(\game_inst.vga_inst.px[9] ),
    .B_N(\game_inst.apple_inst.i_snake_x[4] ),
    .Y(_0380_));
 sg13g2_nor2_1 _1296_ (.A(_0353_),
    .B(_0380_),
    .Y(_0381_));
 sg13g2_o21ai_1 _1297_ (.B1(_0381_),
    .Y(_0382_),
    .A1(_0352_),
    .A2(_0355_));
 sg13g2_nor2b_1 _1298_ (.A(_0380_),
    .B_N(_0349_),
    .Y(_0383_));
 sg13g2_nor2b_2 _1299_ (.A(\game_inst.vga_inst.px[5] ),
    .B_N(net139),
    .Y(_0384_));
 sg13g2_xnor2_1 _1300_ (.Y(_0385_),
    .A(net139),
    .B(net148));
 sg13g2_nand4_1 _1301_ (.B(_0354_),
    .C(_0383_),
    .A(_0351_),
    .Y(_0386_),
    .D(_0385_));
 sg13g2_nand3_1 _1302_ (.B(_0366_),
    .C(_0368_),
    .A(_0363_),
    .Y(_0387_));
 sg13g2_nor2_2 _1303_ (.A(_0272_),
    .B(_0281_),
    .Y(_0388_));
 sg13g2_nor4_1 _1304_ (.A(_0263_),
    .B(\game_inst.vga_inst.px[9] ),
    .C(net145),
    .D(_0388_),
    .Y(_0389_));
 sg13g2_nand3_1 _1305_ (.B(_0365_),
    .C(_0370_),
    .A(\game_inst.apple_inst.i_snake_valid ),
    .Y(_0390_));
 sg13g2_nor3_1 _1306_ (.A(_0387_),
    .B(_0389_),
    .C(_0390_),
    .Y(_0391_));
 sg13g2_nand2_1 _1307_ (.Y(_0392_),
    .A(_0281_),
    .B(_0351_));
 sg13g2_a21oi_1 _1308_ (.A1(_0348_),
    .A2(_0384_),
    .Y(_0393_),
    .B1(_0346_));
 sg13g2_nor2_1 _1309_ (.A(_0392_),
    .B(_0393_),
    .Y(_0394_));
 sg13g2_a21oi_1 _1310_ (.A1(net136),
    .A2(net145),
    .Y(_0395_),
    .B1(_0345_));
 sg13g2_nand2b_1 _1311_ (.Y(_0396_),
    .B(_0395_),
    .A_N(_0388_));
 sg13g2_o21ai_1 _1312_ (.B1(_0380_),
    .Y(_0397_),
    .A1(\game_inst.apple_inst.i_snake_x[3] ),
    .A2(_0271_));
 sg13g2_o21ai_1 _1313_ (.B1(_0397_),
    .Y(_0398_),
    .A1(_0381_),
    .A2(_0388_));
 sg13g2_o21ai_1 _1314_ (.B1(_0398_),
    .Y(_0399_),
    .A1(_0394_),
    .A2(_0396_));
 sg13g2_nand4_1 _1315_ (.B(_0386_),
    .C(_0391_),
    .A(_0382_),
    .Y(_0400_),
    .D(_0399_));
 sg13g2_nand2_1 _1316_ (.Y(_0401_),
    .A(net139),
    .B(net138));
 sg13g2_nand3_1 _1317_ (.B(\game_inst.apple_inst.i_snake_x[1] ),
    .C(net137),
    .A(net139),
    .Y(_0402_));
 sg13g2_a21o_1 _1318_ (.A2(\game_inst.apple_inst.i_snake_x[1] ),
    .A1(net139),
    .B1(\game_inst.apple_inst.i_snake_x[2] ),
    .X(_0403_));
 sg13g2_and3_1 _1319_ (.X(_0404_),
    .A(_0272_),
    .B(_0402_),
    .C(_0403_));
 sg13g2_o21ai_1 _1320_ (.B1(_0401_),
    .Y(_0405_),
    .A1(_0348_),
    .A2(_0384_));
 sg13g2_nand2_1 _1321_ (.Y(_0406_),
    .A(_0279_),
    .B(_0405_));
 sg13g2_nand3_1 _1322_ (.B(_0402_),
    .C(_0403_),
    .A(net147),
    .Y(_0407_));
 sg13g2_a21o_1 _1323_ (.A2(_0403_),
    .A1(_0402_),
    .B1(net147),
    .X(_0408_));
 sg13g2_nand2_1 _1324_ (.Y(_0409_),
    .A(_0407_),
    .B(_0408_));
 sg13g2_a22oi_1 _1325_ (.Y(_0410_),
    .B1(_0407_),
    .B2(_0408_),
    .A2(_0405_),
    .A1(_0279_));
 sg13g2_xnor2_1 _1326_ (.Y(_0411_),
    .A(_0354_),
    .B(_0402_));
 sg13g2_or3_1 _1327_ (.A(_0404_),
    .B(_0410_),
    .C(_0411_),
    .X(_0412_));
 sg13g2_o21ai_1 _1328_ (.B1(_0411_),
    .Y(_0413_),
    .A1(_0404_),
    .A2(_0410_));
 sg13g2_and2_1 _1329_ (.A(_0412_),
    .B(_0413_),
    .X(_0414_));
 sg13g2_nand4_1 _1330_ (.B(_0377_),
    .C(_0412_),
    .A(_0356_),
    .Y(_0415_),
    .D(_0413_));
 sg13g2_a221oi_1 _1331_ (.B2(_0378_),
    .C1(_0357_),
    .B1(_0414_),
    .A1(_0379_),
    .Y(_0416_),
    .A2(_0400_));
 sg13g2_a21oi_1 _1332_ (.A1(net116),
    .A2(_0416_),
    .Y(_0417_),
    .B1(net352));
 sg13g2_nor2_1 _1333_ (.A(net127),
    .B(_0417_),
    .Y(_0032_));
 sg13g2_nand3b_1 _1334_ (.B(_0341_),
    .C(\game_inst.vga_inst.prev_dir[0] ),
    .Y(_0418_),
    .A_N(\game_inst.vga_inst.prev_dir[1] ));
 sg13g2_nand2_1 _1335_ (.Y(_0419_),
    .A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[0] [0]),
    .B(_0335_));
 sg13g2_o21ai_1 _1336_ (.B1(_0418_),
    .Y(_0420_),
    .A1(net134),
    .A2(_0419_));
 sg13g2_a21oi_1 _1337_ (.A1(_0416_),
    .A2(net115),
    .Y(_0421_),
    .B1(net356));
 sg13g2_nor2_1 _1338_ (.A(net127),
    .B(_0421_),
    .Y(_0033_));
 sg13g2_nand2_1 _1339_ (.Y(_0422_),
    .A(\game_inst.vga_inst.prev_dir[1] ),
    .B(_0342_));
 sg13g2_o21ai_1 _1340_ (.B1(_0422_),
    .Y(_0423_),
    .A1(_0270_),
    .A2(_0336_));
 sg13g2_a21oi_1 _1341_ (.A1(_0416_),
    .A2(net114),
    .Y(_0424_),
    .B1(net348));
 sg13g2_nor2_1 _1342_ (.A(net128),
    .B(_0424_),
    .Y(_0034_));
 sg13g2_nand3_1 _1343_ (.B(\game_inst.vga_inst.prev_dir[1] ),
    .C(_0341_),
    .A(\game_inst.vga_inst.prev_dir[0] ),
    .Y(_0425_));
 sg13g2_o21ai_1 _1344_ (.B1(_0425_),
    .Y(_0426_),
    .A1(_0270_),
    .A2(_0419_));
 sg13g2_a21oi_1 _1345_ (.A1(_0416_),
    .A2(net113),
    .Y(_0427_),
    .B1(net355));
 sg13g2_nor2_1 _1346_ (.A(net128),
    .B(_0427_),
    .Y(_0035_));
 sg13g2_o21ai_1 _1347_ (.B1(_0356_),
    .Y(_0428_),
    .A1(_0234_),
    .A2(_0415_));
 sg13g2_xnor2_1 _1348_ (.Y(_0429_),
    .A(_0406_),
    .B(_0409_));
 sg13g2_xor2_1 _1349_ (.B(_0351_),
    .A(_0350_),
    .X(_0430_));
 sg13g2_a21oi_1 _1350_ (.A1(_0356_),
    .A2(_0377_),
    .Y(_0431_),
    .B1(_0430_));
 sg13g2_a21o_1 _1351_ (.A2(_0429_),
    .A1(_0378_),
    .B1(_0431_),
    .X(_0432_));
 sg13g2_a21oi_1 _1352_ (.A1(_0378_),
    .A2(_0429_),
    .Y(_0433_),
    .B1(_0431_));
 sg13g2_xor2_1 _1353_ (.B(_0349_),
    .A(_0347_),
    .X(_0434_));
 sg13g2_xnor2_1 _1354_ (.Y(_0435_),
    .A(_0347_),
    .B(_0349_));
 sg13g2_a21oi_1 _1355_ (.A1(_0356_),
    .A2(_0377_),
    .Y(_0436_),
    .B1(_0434_));
 sg13g2_xnor2_1 _1356_ (.Y(_0437_),
    .A(_0349_),
    .B(_0384_));
 sg13g2_xor2_1 _1357_ (.B(_0384_),
    .A(_0349_),
    .X(_0438_));
 sg13g2_a21oi_1 _1358_ (.A1(_0356_),
    .A2(_0377_),
    .Y(_0439_),
    .B1(_0435_));
 sg13g2_a221oi_1 _1359_ (.B2(_0378_),
    .C1(_0436_),
    .B1(_0438_),
    .A1(_0379_),
    .Y(_0440_),
    .A2(_0400_));
 sg13g2_xnor2_1 _1360_ (.Y(_0441_),
    .A(_0379_),
    .B(_0385_));
 sg13g2_xor2_1 _1361_ (.B(_0385_),
    .A(_0379_),
    .X(_0442_));
 sg13g2_and4_1 _1362_ (.A(_0428_),
    .B(_0433_),
    .C(_0440_),
    .D(_0442_),
    .X(_0443_));
 sg13g2_a21oi_1 _1363_ (.A1(net116),
    .A2(_0443_),
    .Y(_0444_),
    .B1(net443));
 sg13g2_and2_1 _1364_ (.A(net127),
    .B(_0417_),
    .X(_0445_));
 sg13g2_a21oi_1 _1365_ (.A1(net124),
    .A2(_0444_),
    .Y(_0028_),
    .B1(_0445_));
 sg13g2_a21oi_1 _1366_ (.A1(net115),
    .A2(_0443_),
    .Y(_0446_),
    .B1(net449));
 sg13g2_and2_1 _1367_ (.A(net127),
    .B(_0421_),
    .X(_0447_));
 sg13g2_a21oi_1 _1368_ (.A1(net124),
    .A2(_0446_),
    .Y(_0029_),
    .B1(_0447_));
 sg13g2_a21oi_1 _1369_ (.A1(net114),
    .A2(_0443_),
    .Y(_0448_),
    .B1(net413));
 sg13g2_and2_1 _1370_ (.A(net127),
    .B(_0424_),
    .X(_0449_));
 sg13g2_a21oi_1 _1371_ (.A1(net124),
    .A2(_0448_),
    .Y(_0030_),
    .B1(_0449_));
 sg13g2_a21oi_1 _1372_ (.A1(net113),
    .A2(_0443_),
    .Y(_0450_),
    .B1(net438));
 sg13g2_and2_1 _1373_ (.A(net128),
    .B(_0427_),
    .X(_0451_));
 sg13g2_a21oi_1 _1374_ (.A1(net124),
    .A2(_0450_),
    .Y(_0031_),
    .B1(_0451_));
 sg13g2_and4_1 _1375_ (.A(_0428_),
    .B(_0433_),
    .C(_0440_),
    .D(_0441_),
    .X(_0452_));
 sg13g2_a21o_1 _1376_ (.A2(_0452_),
    .A1(net116),
    .B1(net369),
    .X(_0453_));
 sg13g2_a221oi_1 _1377_ (.B2(_0452_),
    .C1(net369),
    .B1(net116),
    .A1(net149),
    .Y(_0454_),
    .A2(_0322_));
 sg13g2_a21oi_1 _1378_ (.A1(net127),
    .A2(_0444_),
    .Y(_0024_),
    .B1(net370));
 sg13g2_a21o_1 _1379_ (.A2(_0452_),
    .A1(net115),
    .B1(net372),
    .X(_0455_));
 sg13g2_a221oi_1 _1380_ (.B2(_0452_),
    .C1(net372),
    .B1(net115),
    .A1(net149),
    .Y(_0456_),
    .A2(_0322_));
 sg13g2_a21oi_1 _1381_ (.A1(net127),
    .A2(_0446_),
    .Y(_0025_),
    .B1(net373));
 sg13g2_a21o_1 _1382_ (.A2(_0452_),
    .A1(net114),
    .B1(net360),
    .X(_0457_));
 sg13g2_a221oi_1 _1383_ (.B2(_0452_),
    .C1(net360),
    .B1(net114),
    .A1(net149),
    .Y(_0458_),
    .A2(_0322_));
 sg13g2_a21oi_1 _1384_ (.A1(net127),
    .A2(_0448_),
    .Y(_0026_),
    .B1(net361));
 sg13g2_a21o_1 _1385_ (.A2(_0452_),
    .A1(net113),
    .B1(net366),
    .X(_0459_));
 sg13g2_a221oi_1 _1386_ (.B2(_0452_),
    .C1(net366),
    .B1(net113),
    .A1(net149),
    .Y(_0460_),
    .A2(_0322_));
 sg13g2_a21oi_1 _1387_ (.A1(net130),
    .A2(_0450_),
    .Y(_0027_),
    .B1(net367));
 sg13g2_a221oi_1 _1388_ (.B2(_0378_),
    .C1(_0439_),
    .B1(_0437_),
    .A1(_0379_),
    .Y(_0461_),
    .A2(_0400_));
 sg13g2_and4_1 _1389_ (.A(_0428_),
    .B(_0433_),
    .C(_0442_),
    .D(_0461_),
    .X(_0462_));
 sg13g2_a21o_1 _1390_ (.A2(_0462_),
    .A1(net116),
    .B1(net539),
    .X(_0463_));
 sg13g2_mux2_1 _1391_ (.A0(_0453_),
    .A1(_0463_),
    .S(net123),
    .X(_0020_));
 sg13g2_a21o_1 _1392_ (.A2(_0462_),
    .A1(net115),
    .B1(net538),
    .X(_0464_));
 sg13g2_mux2_1 _1393_ (.A0(_0455_),
    .A1(_0464_),
    .S(net123),
    .X(_0021_));
 sg13g2_a21o_1 _1394_ (.A2(_0462_),
    .A1(net114),
    .B1(net547),
    .X(_0465_));
 sg13g2_mux2_1 _1395_ (.A0(_0457_),
    .A1(_0465_),
    .S(net123),
    .X(_0022_));
 sg13g2_a21o_1 _1396_ (.A2(_0462_),
    .A1(net113),
    .B1(net549),
    .X(_0466_));
 sg13g2_mux2_1 _1397_ (.A0(_0459_),
    .A1(_0466_),
    .S(net123),
    .X(_0023_));
 sg13g2_and4_1 _1398_ (.A(_0428_),
    .B(_0433_),
    .C(_0441_),
    .D(_0461_),
    .X(_0467_));
 sg13g2_a21o_1 _1399_ (.A2(_0467_),
    .A1(net116),
    .B1(net550),
    .X(_0468_));
 sg13g2_mux2_1 _1400_ (.A0(_0463_),
    .A1(_0468_),
    .S(net123),
    .X(_0016_));
 sg13g2_a21o_1 _1401_ (.A2(_0467_),
    .A1(net115),
    .B1(net536),
    .X(_0469_));
 sg13g2_mux2_1 _1402_ (.A0(_0464_),
    .A1(_0469_),
    .S(net123),
    .X(_0017_));
 sg13g2_a21o_1 _1403_ (.A2(_0467_),
    .A1(net114),
    .B1(net543),
    .X(_0470_));
 sg13g2_mux2_1 _1404_ (.A0(_0465_),
    .A1(_0470_),
    .S(net124),
    .X(_0018_));
 sg13g2_a21o_1 _1405_ (.A2(_0467_),
    .A1(net113),
    .B1(net554),
    .X(_0471_));
 sg13g2_mux2_1 _1406_ (.A0(_0466_),
    .A1(_0471_),
    .S(net125),
    .X(_0019_));
 sg13g2_and4_1 _1407_ (.A(_0428_),
    .B(_0432_),
    .C(_0440_),
    .D(_0442_),
    .X(_0472_));
 sg13g2_a21o_1 _1408_ (.A2(_0472_),
    .A1(net116),
    .B1(net553),
    .X(_0473_));
 sg13g2_mux2_1 _1409_ (.A0(_0468_),
    .A1(_0473_),
    .S(net123),
    .X(_0012_));
 sg13g2_a21o_1 _1410_ (.A2(_0472_),
    .A1(net115),
    .B1(net555),
    .X(_0474_));
 sg13g2_mux2_1 _1411_ (.A0(_0469_),
    .A1(_0474_),
    .S(net123),
    .X(_0013_));
 sg13g2_a21o_1 _1412_ (.A2(_0472_),
    .A1(net114),
    .B1(net558),
    .X(_0475_));
 sg13g2_mux2_1 _1413_ (.A0(_0470_),
    .A1(_0475_),
    .S(net125),
    .X(_0014_));
 sg13g2_a21o_1 _1414_ (.A2(_0472_),
    .A1(net113),
    .B1(net551),
    .X(_0476_));
 sg13g2_mux2_1 _1415_ (.A0(_0471_),
    .A1(_0476_),
    .S(net125),
    .X(_0015_));
 sg13g2_and4_1 _1416_ (.A(_0428_),
    .B(_0432_),
    .C(_0440_),
    .D(_0441_),
    .X(_0477_));
 sg13g2_a21o_1 _1417_ (.A2(_0477_),
    .A1(net116),
    .B1(net540),
    .X(_0478_));
 sg13g2_mux2_1 _1418_ (.A0(_0473_),
    .A1(_0478_),
    .S(net125),
    .X(_0008_));
 sg13g2_a21o_1 _1419_ (.A2(_0477_),
    .A1(net115),
    .B1(net545),
    .X(_0479_));
 sg13g2_mux2_1 _1420_ (.A0(_0474_),
    .A1(_0479_),
    .S(net125),
    .X(_0009_));
 sg13g2_a21o_1 _1421_ (.A2(_0477_),
    .A1(net114),
    .B1(\game_inst.vga_inst.row_buffer[2][2] ),
    .X(_0480_));
 sg13g2_mux2_1 _1422_ (.A0(_0475_),
    .A1(_0480_),
    .S(net126),
    .X(_0010_));
 sg13g2_a21o_1 _1423_ (.A2(_0477_),
    .A1(net113),
    .B1(net560),
    .X(_0481_));
 sg13g2_mux2_1 _1424_ (.A0(_0476_),
    .A1(_0481_),
    .S(net126),
    .X(_0011_));
 sg13g2_and4_1 _1425_ (.A(_0428_),
    .B(_0432_),
    .C(_0442_),
    .D(_0461_),
    .X(_0482_));
 sg13g2_a21o_1 _1426_ (.A2(_0482_),
    .A1(_0344_),
    .B1(net542),
    .X(_0483_));
 sg13g2_mux2_1 _1427_ (.A0(_0478_),
    .A1(_0483_),
    .S(net125),
    .X(_0004_));
 sg13g2_a21o_1 _1428_ (.A2(_0482_),
    .A1(_0420_),
    .B1(\game_inst.vga_inst.row_buffer[1][1] ),
    .X(_0484_));
 sg13g2_mux2_1 _1429_ (.A0(_0479_),
    .A1(_0484_),
    .S(net125),
    .X(_0005_));
 sg13g2_a21o_1 _1430_ (.A2(_0482_),
    .A1(_0423_),
    .B1(net562),
    .X(_0485_));
 sg13g2_mux2_1 _1431_ (.A0(_0480_),
    .A1(_0485_),
    .S(net125),
    .X(_0006_));
 sg13g2_a21o_1 _1432_ (.A2(_0482_),
    .A1(_0426_),
    .B1(\game_inst.vga_inst.row_buffer[1][3] ),
    .X(_0486_));
 sg13g2_mux2_1 _1433_ (.A0(_0481_),
    .A1(_0486_),
    .S(net126),
    .X(_0007_));
 sg13g2_nor2_1 _1434_ (.A(net155),
    .B(net6),
    .Y(_0487_));
 sg13g2_nand2b_1 _1435_ (.Y(_0488_),
    .B(net157),
    .A_N(net6));
 sg13g2_nand4_1 _1436_ (.B(\game_inst.snake_inst.pos[5] ),
    .C(_0258_),
    .A(\game_inst.snake_inst.pos[7] ),
    .Y(_0489_),
    .D(\game_inst.snake_inst.pos[6] ));
 sg13g2_nand2b_1 _1437_ (.Y(_0490_),
    .B(\game_inst.snake_inst.pos[3] ),
    .A_N(\game_inst.snake_inst.pos[2] ));
 sg13g2_nand3_1 _1438_ (.B(\game_inst.apple_inst.o_ready ),
    .C(_0338_),
    .A(\game_inst.tick ),
    .Y(_0491_));
 sg13g2_or3_1 _1439_ (.A(_0489_),
    .B(_0490_),
    .C(_0491_),
    .X(_0492_));
 sg13g2_inv_2 _1440_ (.Y(_0493_),
    .A(net121));
 sg13g2_o21ai_1 _1441_ (.B1(net132),
    .Y(_0494_),
    .A1(_0240_),
    .A2(net122));
 sg13g2_a21o_2 _1442_ (.A2(net120),
    .A1(net482),
    .B1(_0494_),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[0] [0]));
 sg13g2_nor2_2 _1443_ (.A(_0239_),
    .B(net121),
    .Y(_0495_));
 sg13g2_nand2_1 _1444_ (.Y(_0496_),
    .A(net141),
    .B(_0493_));
 sg13g2_nand2_1 _1445_ (.Y(_0497_),
    .A(net131),
    .B(_0496_));
 sg13g2_a21o_2 _1446_ (.A2(net120),
    .A1(net478),
    .B1(_0497_),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[0] [0]));
 sg13g2_or2_1 _1447_ (.X(uo_out[5]),
    .B(\game_inst.vga_inst.color[2] ),
    .A(\game_inst.vga_inst.color[3] ));
 sg13g2_or2_1 _1448_ (.X(uo_out[4]),
    .B(\game_inst.vga_inst.color[3] ),
    .A(\game_inst.vga_inst.color[1] ));
 sg13g2_o21ai_1 _1449_ (.B1(net131),
    .Y(_0039_),
    .A1(net359),
    .A2(_0493_));
 sg13g2_or4_1 _1450_ (.A(\game_inst.snake_inst.pos[1] ),
    .B(_0257_),
    .C(_0489_),
    .D(_0490_),
    .X(_0498_));
 sg13g2_and2_1 _1451_ (.A(net120),
    .B(_0498_),
    .X(_0499_));
 sg13g2_nand2_2 _1452_ (.Y(_0500_),
    .A(net120),
    .B(_0498_));
 sg13g2_and2_1 _1453_ (.A(net534),
    .B(net359),
    .X(_0501_));
 sg13g2_and2_1 _1454_ (.A(net460),
    .B(_0501_),
    .X(_0502_));
 sg13g2_xnor2_1 _1455_ (.Y(_0503_),
    .A(net535),
    .B(_0502_));
 sg13g2_o21ai_1 _1456_ (.B1(net131),
    .Y(_0040_),
    .A1(_0500_),
    .A2(_0503_));
 sg13g2_and3_2 _1457_ (.X(_0504_),
    .A(net535),
    .B(net393),
    .C(_0502_));
 sg13g2_a21oi_1 _1458_ (.A1(net564),
    .A2(_0504_),
    .Y(_0505_),
    .B1(net117));
 sg13g2_o21ai_1 _1459_ (.B1(_0505_),
    .Y(_0506_),
    .A1(net564),
    .A2(_0504_));
 sg13g2_nand2_1 _1460_ (.Y(_0041_),
    .A(net132),
    .B(_0506_));
 sg13g2_a21oi_1 _1461_ (.A1(\game_inst.snake_inst.pos[5] ),
    .A2(_0504_),
    .Y(_0507_),
    .B1(net508));
 sg13g2_nand3_1 _1462_ (.B(net508),
    .C(_0504_),
    .A(net564),
    .Y(_0508_));
 sg13g2_nand2_1 _1463_ (.Y(_0509_),
    .A(_0499_),
    .B(_0508_));
 sg13g2_o21ai_1 _1464_ (.B1(net132),
    .Y(_0042_),
    .A1(net509),
    .A2(_0509_));
 sg13g2_xor2_1 _1465_ (.B(_0508_),
    .A(net404),
    .X(_0510_));
 sg13g2_o21ai_1 _1466_ (.B1(net131),
    .Y(_0043_),
    .A1(_0500_),
    .A2(_0510_));
 sg13g2_nor2b_1 _1467_ (.A(\game_inst.vga_inst.px[7] ),
    .B_N(net144),
    .Y(_0511_));
 sg13g2_and4_1 _1468_ (.A(net146),
    .B(_0278_),
    .C(net129),
    .D(_0511_),
    .X(_0512_));
 sg13g2_nand4_1 _1469_ (.B(_0278_),
    .C(net129),
    .A(net146),
    .Y(_0513_),
    .D(_0511_));
 sg13g2_nor2_2 _1470_ (.A(net154),
    .B(_0512_),
    .Y(_0514_));
 sg13g2_nand2_2 _1471_ (.Y(_0515_),
    .A(net156),
    .B(_0513_));
 sg13g2_nor2_1 _1472_ (.A(net343),
    .B(net154),
    .Y(_0044_));
 sg13g2_xnor2_1 _1473_ (.Y(_0516_),
    .A(net343),
    .B(net436));
 sg13g2_nor2_1 _1474_ (.A(_0515_),
    .B(_0516_),
    .Y(_0045_));
 sg13g2_a21oi_1 _1475_ (.A1(net343),
    .A2(\game_inst.vga_inst.px[1] ),
    .Y(_0517_),
    .B1(net383));
 sg13g2_nor3_1 _1476_ (.A(net154),
    .B(_0321_),
    .C(net384),
    .Y(_0046_));
 sg13g2_o21ai_1 _1477_ (.B1(net156),
    .Y(_0518_),
    .A1(net517),
    .A2(_0321_));
 sg13g2_nor2_1 _1478_ (.A(_0322_),
    .B(_0518_),
    .Y(_0047_));
 sg13g2_o21ai_1 _1479_ (.B1(net156),
    .Y(_0519_),
    .A1(net493),
    .A2(_0322_));
 sg13g2_nor2_1 _1480_ (.A(net129),
    .B(net494),
    .Y(_0048_));
 sg13g2_xnor2_1 _1481_ (.Y(_0520_),
    .A(net148),
    .B(net129));
 sg13g2_nor2_1 _1482_ (.A(_0515_),
    .B(_0520_),
    .Y(_0049_));
 sg13g2_a21oi_1 _1483_ (.A1(net148),
    .A2(net129),
    .Y(_0521_),
    .B1(net475));
 sg13g2_nor2_1 _1484_ (.A(net476),
    .B(net126),
    .Y(_0522_));
 sg13g2_nor3_1 _1485_ (.A(_0515_),
    .B(_0521_),
    .C(_0522_),
    .Y(_0050_));
 sg13g2_and2_1 _1486_ (.A(net129),
    .B(_0388_),
    .X(_0523_));
 sg13g2_nor2_1 _1487_ (.A(net473),
    .B(_0522_),
    .Y(_0524_));
 sg13g2_nor3_1 _1488_ (.A(_0515_),
    .B(_0523_),
    .C(_0524_),
    .Y(_0051_));
 sg13g2_or2_1 _1489_ (.X(_0525_),
    .B(_0523_),
    .A(net145));
 sg13g2_nand2_1 _1490_ (.Y(_0526_),
    .A(net145),
    .B(_0523_));
 sg13g2_and3_1 _1491_ (.X(_0052_),
    .A(_0514_),
    .B(_0525_),
    .C(_0526_));
 sg13g2_xor2_1 _1492_ (.B(_0526_),
    .A(net144),
    .X(_0527_));
 sg13g2_nor2_1 _1493_ (.A(_0515_),
    .B(net574),
    .Y(_0053_));
 sg13g2_a21oi_2 _1494_ (.B1(\game_inst.sound_inst.phase[4] ),
    .Y(_0528_),
    .A2(\game_inst.sound_inst.phase[2] ),
    .A1(\game_inst.sound_inst.phase[3] ));
 sg13g2_xnor2_1 _1495_ (.Y(_0529_),
    .A(\game_inst.sound_inst.max_counter[2] ),
    .B(_0528_));
 sg13g2_nand2b_1 _1496_ (.Y(_0530_),
    .B(\game_inst.sound_inst.max_counter[1] ),
    .A_N(_0528_));
 sg13g2_xor2_1 _1497_ (.B(_0528_),
    .A(\game_inst.sound_inst.max_counter[1] ),
    .X(_0531_));
 sg13g2_o21ai_1 _1498_ (.B1(_0530_),
    .Y(_0532_),
    .A1(_0250_),
    .A2(_0531_));
 sg13g2_nand2_1 _1499_ (.Y(_0533_),
    .A(_0529_),
    .B(_0532_));
 sg13g2_nor2b_1 _1500_ (.A(\game_inst.sound_inst.prev_vsync ),
    .B_N(\game_inst.sound_inst.vsync_pulse ),
    .Y(_0534_));
 sg13g2_nand2_1 _1501_ (.Y(_0535_),
    .A(net430),
    .B(_0534_));
 sg13g2_nor2_2 _1502_ (.A(net432),
    .B(_0535_),
    .Y(_0536_));
 sg13g2_inv_1 _1503_ (.Y(_0537_),
    .A(_0536_));
 sg13g2_o21ai_1 _1504_ (.B1(_0536_),
    .Y(_0538_),
    .A1(_0529_),
    .A2(_0532_));
 sg13g2_inv_1 _1505_ (.Y(_0539_),
    .A(_0538_));
 sg13g2_nand2_1 _1506_ (.Y(_0540_),
    .A(\game_inst.o_tick ),
    .B(net404));
 sg13g2_nor2_1 _1507_ (.A(net430),
    .B(net432),
    .Y(_0541_));
 sg13g2_nor2b_2 _1508_ (.A(_0540_),
    .B_N(_0541_),
    .Y(_0542_));
 sg13g2_inv_1 _1509_ (.Y(_0543_),
    .A(_0542_));
 sg13g2_a221oi_1 _1510_ (.B2(_0533_),
    .C1(_0542_),
    .B1(_0539_),
    .A1(net556),
    .Y(_0544_),
    .A2(_0537_));
 sg13g2_xor2_1 _1511_ (.B(net136),
    .A(\game_inst.head_x[3] ),
    .X(_0545_));
 sg13g2_xor2_1 _1512_ (.B(\game_inst.apple_inst.i_snake_y[3] ),
    .A(\game_inst.head_y[3] ),
    .X(_0546_));
 sg13g2_xor2_1 _1513_ (.B(net137),
    .A(\game_inst.head_x[2] ),
    .X(_0547_));
 sg13g2_nor2b_1 _1514_ (.A(\game_inst.apple_inst.i_snake_y[2] ),
    .B_N(\game_inst.head_y[2] ),
    .Y(_0548_));
 sg13g2_xor2_1 _1515_ (.B(\game_inst.apple_inst.i_snake_y[1] ),
    .A(\game_inst.head_y[1] ),
    .X(_0549_));
 sg13g2_xor2_1 _1516_ (.B(net138),
    .A(\game_inst.head_x[1] ),
    .X(_0550_));
 sg13g2_nor2b_1 _1517_ (.A(\game_inst.apple_inst.i_snake_y[0] ),
    .B_N(\game_inst.head_y[0] ),
    .Y(_0551_));
 sg13g2_xor2_1 _1518_ (.B(\game_inst.apple_inst.i_snake_x[4] ),
    .A(\game_inst.head_x[4] ),
    .X(_0552_));
 sg13g2_nor3_1 _1519_ (.A(_0545_),
    .B(_0546_),
    .C(_0549_),
    .Y(_0553_));
 sg13g2_a221oi_1 _1520_ (.B2(_0236_),
    .C1(_0547_),
    .B1(\game_inst.apple_inst.i_snake_y[0] ),
    .A1(\game_inst.head_x[0] ),
    .Y(_0554_),
    .A2(_0260_));
 sg13g2_a22oi_1 _1521_ (.Y(_0555_),
    .B1(\game_inst.apple_inst.i_snake_y[2] ),
    .B2(_0235_),
    .A2(net140),
    .A1(_0238_));
 sg13g2_nor4_1 _1522_ (.A(_0548_),
    .B(_0550_),
    .C(_0551_),
    .D(_0552_),
    .Y(_0556_));
 sg13g2_nand4_1 _1523_ (.B(_0554_),
    .C(_0555_),
    .A(_0553_),
    .Y(_0557_),
    .D(_0556_));
 sg13g2_nand2_1 _1524_ (.Y(_0558_),
    .A(\game_inst.head_x[4] ),
    .B(\game_inst.head_x[1] ));
 sg13g2_o21ai_1 _1525_ (.B1(_0238_),
    .Y(_0559_),
    .A1(\game_inst.head_x[4] ),
    .A2(\game_inst.head_x[1] ));
 sg13g2_a21oi_1 _1526_ (.A1(\game_inst.head_x[0] ),
    .A2(_0558_),
    .Y(_0560_),
    .B1(\game_inst.head_x[3] ));
 sg13g2_nand3b_1 _1527_ (.B(_0559_),
    .C(_0560_),
    .Y(_0561_),
    .A_N(\game_inst.head_x[2] ));
 sg13g2_and3_1 _1528_ (.X(_0562_),
    .A(\game_inst.head_y[3] ),
    .B(\game_inst.head_y[2] ),
    .C(\game_inst.head_y[1] ));
 sg13g2_nor3_1 _1529_ (.A(\game_inst.head_y[3] ),
    .B(\game_inst.head_y[2] ),
    .C(\game_inst.head_y[1] ),
    .Y(_0563_));
 sg13g2_o21ai_1 _1530_ (.B1(_0236_),
    .Y(_0564_),
    .A1(_0562_),
    .A2(_0563_));
 sg13g2_nand3_1 _1531_ (.B(_0561_),
    .C(_0564_),
    .A(_0557_),
    .Y(_0565_));
 sg13g2_nand3_1 _1532_ (.B(_0341_),
    .C(_0565_),
    .A(net435),
    .Y(_0566_));
 sg13g2_and4_1 _1533_ (.A(net435),
    .B(\game_inst.o_tick ),
    .C(_0341_),
    .D(_0565_),
    .X(_0567_));
 sg13g2_and2_1 _1534_ (.A(\game_inst.o_tick ),
    .B(\game_inst.o_success ),
    .X(_0568_));
 sg13g2_xnor2_1 _1535_ (.Y(_0569_),
    .A(\game_inst.apple_inst.i_snake_y[3] ),
    .B(\game_inst.apple_inst.apple_y[3] ));
 sg13g2_xnor2_1 _1536_ (.Y(_0570_),
    .A(net137),
    .B(\game_inst.apple_inst.apple_x[2] ));
 sg13g2_a22oi_1 _1537_ (.Y(_0571_),
    .B1(\game_inst.apple_inst.i_snake_y[1] ),
    .B2(_0267_),
    .A2(_0260_),
    .A1(\game_inst.apple_inst.apple_x[0] ));
 sg13g2_xnor2_1 _1538_ (.Y(_0572_),
    .A(net136),
    .B(\game_inst.apple_inst.apple_x[3] ));
 sg13g2_a22oi_1 _1539_ (.Y(_0573_),
    .B1(_0266_),
    .B2(\game_inst.apple_inst.apple_y[1] ),
    .A2(net140),
    .A1(_0259_));
 sg13g2_a22oi_1 _1540_ (.Y(_0574_),
    .B1(_0263_),
    .B2(\game_inst.apple_inst.apple_x[4] ),
    .A2(_0262_),
    .A1(\game_inst.apple_inst.i_snake_x[1] ));
 sg13g2_nand4_1 _1541_ (.B(_0572_),
    .C(_0573_),
    .A(_0571_),
    .Y(_0575_),
    .D(_0574_));
 sg13g2_xor2_1 _1542_ (.B(\game_inst.apple_inst.i_snake_y[0] ),
    .A(\game_inst.apple_inst.apple_y[0] ),
    .X(_0576_));
 sg13g2_a221oi_1 _1543_ (.B2(_0264_),
    .C1(_0576_),
    .B1(\game_inst.apple_inst.i_snake_x[4] ),
    .A1(_0261_),
    .Y(_0577_),
    .A2(\game_inst.apple_inst.apple_x[1] ));
 sg13g2_xnor2_1 _1544_ (.Y(_0578_),
    .A(\game_inst.apple_inst.i_snake_y[2] ),
    .B(\game_inst.apple_inst.apple_y[2] ));
 sg13g2_nand4_1 _1545_ (.B(_0570_),
    .C(_0577_),
    .A(_0569_),
    .Y(_0579_),
    .D(_0578_));
 sg13g2_nor2_1 _1546_ (.A(_0575_),
    .B(_0579_),
    .Y(_0580_));
 sg13g2_nand2_1 _1547_ (.Y(_0581_),
    .A(net419),
    .B(_0340_));
 sg13g2_nor3_2 _1548_ (.A(_0575_),
    .B(_0579_),
    .C(_0581_),
    .Y(_0582_));
 sg13g2_or2_1 _1549_ (.X(_0583_),
    .B(_0582_),
    .A(_0568_));
 sg13g2_or2_1 _1550_ (.X(_0584_),
    .B(_0583_),
    .A(_0567_));
 sg13g2_nor3_1 _1551_ (.A(net152),
    .B(net557),
    .C(_0584_),
    .Y(_0054_));
 sg13g2_xnor2_1 _1552_ (.Y(_0585_),
    .A(net519),
    .B(_0531_));
 sg13g2_nor2b_1 _1553_ (.A(_0536_),
    .B_N(net575),
    .Y(_0586_));
 sg13g2_a221oi_1 _1554_ (.B2(_0543_),
    .C1(_0583_),
    .B1(_0586_),
    .A1(_0536_),
    .Y(_0587_),
    .A2(_0585_));
 sg13g2_nor3_1 _1555_ (.A(net150),
    .B(_0567_),
    .C(net576),
    .Y(_0055_));
 sg13g2_nor2b_2 _1556_ (.A(\game_inst.sound_inst.prev_pwm_base ),
    .B_N(net341),
    .Y(_0588_));
 sg13g2_o21ai_1 _1557_ (.B1(_0588_),
    .Y(_0589_),
    .A1(_0251_),
    .A2(\game_inst.sound_inst.max_counter[1] ));
 sg13g2_a21oi_1 _1558_ (.A1(_0251_),
    .A2(\game_inst.sound_inst.max_counter[1] ),
    .Y(_0590_),
    .B1(_0589_));
 sg13g2_xnor2_1 _1559_ (.Y(_0591_),
    .A(\game_inst.sound_inst.max_counter[3] ),
    .B(\game_inst.sound_inst.counter[3] ));
 sg13g2_xnor2_1 _1560_ (.Y(_0592_),
    .A(\game_inst.sound_inst.counter[2] ),
    .B(\game_inst.sound_inst.max_counter[2] ));
 sg13g2_xnor2_1 _1561_ (.Y(_0593_),
    .A(\game_inst.sound_inst.max_counter[0] ),
    .B(\game_inst.sound_inst.counter[0] ));
 sg13g2_nand4_1 _1562_ (.B(_0591_),
    .C(_0592_),
    .A(_0590_),
    .Y(_0594_),
    .D(_0593_));
 sg13g2_and3_1 _1563_ (.X(_0595_),
    .A(\game_inst.sound_inst.phase[2] ),
    .B(\game_inst.sound_inst.mode[1] ),
    .C(\game_inst.sound_inst.mode[0] ));
 sg13g2_nand2_2 _1564_ (.Y(_0596_),
    .A(net132),
    .B(_0594_));
 sg13g2_nand2_1 _1565_ (.Y(_0597_),
    .A(net363),
    .B(_0594_));
 sg13g2_or4_1 _1566_ (.A(net363),
    .B(_0541_),
    .C(_0594_),
    .D(_0595_),
    .X(_0598_));
 sg13g2_a21oi_1 _1567_ (.A1(net364),
    .A2(_0598_),
    .Y(_0056_),
    .B1(net152));
 sg13g2_nor3_1 _1568_ (.A(_0542_),
    .B(_0567_),
    .C(_0568_),
    .Y(_0599_));
 sg13g2_nor2_1 _1569_ (.A(_0542_),
    .B(_0583_),
    .Y(_0600_));
 sg13g2_nor3_1 _1570_ (.A(_0542_),
    .B(_0567_),
    .C(_0583_),
    .Y(_0601_));
 sg13g2_or3_1 _1571_ (.A(_0542_),
    .B(_0567_),
    .C(_0583_),
    .X(_0602_));
 sg13g2_nor3_1 _1572_ (.A(\game_inst.sound_inst.phase[4] ),
    .B(\game_inst.sound_inst.phase[3] ),
    .C(\game_inst.sound_inst.mode[1] ),
    .Y(_0603_));
 sg13g2_a21oi_1 _1573_ (.A1(\game_inst.sound_inst.mode[0] ),
    .A2(_0603_),
    .Y(_0604_),
    .B1(_0249_));
 sg13g2_a21oi_1 _1574_ (.A1(\game_inst.sound_inst.phase[4] ),
    .A2(\game_inst.sound_inst.phase[3] ),
    .Y(_0605_),
    .B1(\game_inst.sound_inst.phase[0] ));
 sg13g2_nor4_1 _1575_ (.A(\game_inst.sound_inst.phase[2] ),
    .B(net390),
    .C(_0604_),
    .D(_0605_),
    .Y(_0606_));
 sg13g2_nor2_1 _1576_ (.A(_0602_),
    .B(_0606_),
    .Y(_0607_));
 sg13g2_nand2_1 _1577_ (.Y(_0608_),
    .A(net432),
    .B(_0607_));
 sg13g2_a21oi_1 _1578_ (.A1(_0599_),
    .A2(net433),
    .Y(_0057_),
    .B1(net152));
 sg13g2_a21oi_1 _1579_ (.A1(net430),
    .A2(_0607_),
    .Y(_0609_),
    .B1(_0584_));
 sg13g2_nor2_1 _1580_ (.A(net152),
    .B(net431),
    .Y(_0058_));
 sg13g2_and2_1 _1581_ (.A(net422),
    .B(_0588_),
    .X(_0610_));
 sg13g2_nor2_1 _1582_ (.A(net422),
    .B(_0588_),
    .Y(_0611_));
 sg13g2_nor3_1 _1583_ (.A(_0596_),
    .B(_0610_),
    .C(net423),
    .Y(_0059_));
 sg13g2_and2_1 _1584_ (.A(net441),
    .B(_0610_),
    .X(_0612_));
 sg13g2_nor2_1 _1585_ (.A(net441),
    .B(_0610_),
    .Y(_0613_));
 sg13g2_nor3_1 _1586_ (.A(_0596_),
    .B(_0612_),
    .C(net442),
    .Y(_0060_));
 sg13g2_nand2_1 _1587_ (.Y(_0614_),
    .A(net454),
    .B(_0612_));
 sg13g2_xnor2_1 _1588_ (.Y(_0615_),
    .A(net454),
    .B(_0612_));
 sg13g2_nor2_1 _1589_ (.A(_0596_),
    .B(_0615_),
    .Y(_0061_));
 sg13g2_xor2_1 _1590_ (.B(_0614_),
    .A(net479),
    .X(_0616_));
 sg13g2_nor2_1 _1591_ (.A(_0596_),
    .B(_0616_),
    .Y(_0062_));
 sg13g2_xnor2_1 _1592_ (.Y(_0617_),
    .A(net519),
    .B(_0536_));
 sg13g2_a21oi_1 _1593_ (.A1(_0601_),
    .A2(net520),
    .Y(_0063_),
    .B1(net150));
 sg13g2_o21ai_1 _1594_ (.B1(_0533_),
    .Y(_0618_),
    .A1(_0252_),
    .A2(_0528_));
 sg13g2_xor2_1 _1595_ (.B(_0528_),
    .A(net523),
    .X(_0619_));
 sg13g2_a21oi_1 _1596_ (.A1(_0618_),
    .A2(_0619_),
    .Y(_0620_),
    .B1(_0537_));
 sg13g2_o21ai_1 _1597_ (.B1(_0620_),
    .Y(_0621_),
    .A1(_0618_),
    .A2(_0619_));
 sg13g2_a21oi_1 _1598_ (.A1(_0600_),
    .A2(_0621_),
    .Y(_0622_),
    .B1(_0567_));
 sg13g2_nor3_1 _1599_ (.A(net523),
    .B(_0536_),
    .C(_0602_),
    .Y(_0623_));
 sg13g2_nor3_1 _1600_ (.A(net150),
    .B(_0622_),
    .C(net524),
    .Y(_0064_));
 sg13g2_nand2_2 _1601_ (.Y(_0624_),
    .A(net133),
    .B(_0601_));
 sg13g2_and2_1 _1602_ (.A(net470),
    .B(_0534_),
    .X(_0625_));
 sg13g2_nor2_1 _1603_ (.A(net470),
    .B(_0534_),
    .Y(_0626_));
 sg13g2_nor3_1 _1604_ (.A(_0624_),
    .B(_0625_),
    .C(net471),
    .Y(_0065_));
 sg13g2_and2_1 _1605_ (.A(net390),
    .B(_0625_),
    .X(_0627_));
 sg13g2_nor2_1 _1606_ (.A(net390),
    .B(_0625_),
    .Y(_0628_));
 sg13g2_nor3_1 _1607_ (.A(_0624_),
    .B(_0627_),
    .C(net391),
    .Y(_0066_));
 sg13g2_and2_1 _1608_ (.A(net490),
    .B(_0627_),
    .X(_0629_));
 sg13g2_nor2_1 _1609_ (.A(net490),
    .B(_0627_),
    .Y(_0630_));
 sg13g2_nor3_1 _1610_ (.A(_0624_),
    .B(_0629_),
    .C(_0630_),
    .Y(_0067_));
 sg13g2_nand2_1 _1611_ (.Y(_0631_),
    .A(net491),
    .B(_0629_));
 sg13g2_xnor2_1 _1612_ (.Y(_0632_),
    .A(net491),
    .B(_0629_));
 sg13g2_nor2_1 _1613_ (.A(_0624_),
    .B(_0632_),
    .Y(_0068_));
 sg13g2_xor2_1 _1614_ (.B(_0631_),
    .A(net502),
    .X(_0633_));
 sg13g2_nor2_1 _1615_ (.A(_0624_),
    .B(_0633_),
    .Y(_0069_));
 sg13g2_o21ai_1 _1616_ (.B1(net121),
    .Y(_0070_),
    .A1(_0256_),
    .A2(net404));
 sg13g2_mux2_1 _1617_ (.A0(net455),
    .A1(_0483_),
    .S(net129),
    .X(_0071_));
 sg13g2_mux2_1 _1618_ (.A0(net439),
    .A1(_0484_),
    .S(net129),
    .X(_0072_));
 sg13g2_mux2_1 _1619_ (.A0(net444),
    .A1(_0485_),
    .S(net130),
    .X(_0073_));
 sg13g2_mux2_1 _1620_ (.A0(net447),
    .A1(_0486_),
    .S(net130),
    .X(_0074_));
 sg13g2_or3_1 _1621_ (.A(\game_inst.vga_inst.py[4] ),
    .B(\game_inst.vga_inst.py[1] ),
    .C(\game_inst.vga_inst.py[0] ),
    .X(_0634_));
 sg13g2_nand3_1 _1622_ (.B(net143),
    .C(\game_inst.vga_inst.py[2] ),
    .A(net353),
    .Y(_0635_));
 sg13g2_nor4_1 _1623_ (.A(\game_inst.vga_inst.py[5] ),
    .B(_0275_),
    .C(_0634_),
    .D(_0635_),
    .Y(_0636_));
 sg13g2_nor2_1 _1624_ (.A(_0513_),
    .B(_0636_),
    .Y(_0637_));
 sg13g2_o21ai_1 _1625_ (.B1(net156),
    .Y(_0638_),
    .A1(net377),
    .A2(net565));
 sg13g2_a21oi_1 _1626_ (.A1(net377),
    .A2(_0512_),
    .Y(_0075_),
    .B1(_0638_));
 sg13g2_a21oi_1 _1627_ (.A1(net377),
    .A2(_0512_),
    .Y(_0639_),
    .B1(net420));
 sg13g2_o21ai_1 _1628_ (.B1(net156),
    .Y(_0640_),
    .A1(_0358_),
    .A2(_0513_));
 sg13g2_nor2_1 _1629_ (.A(_0639_),
    .B(_0640_),
    .Y(_0076_));
 sg13g2_nand2_1 _1630_ (.Y(_0641_),
    .A(net453),
    .B(_0514_));
 sg13g2_nand2_1 _1631_ (.Y(_0642_),
    .A(net156),
    .B(_0637_));
 sg13g2_xor2_1 _1632_ (.B(_0358_),
    .A(net453),
    .X(_0643_));
 sg13g2_o21ai_1 _1633_ (.B1(_0641_),
    .Y(_0077_),
    .A1(_0642_),
    .A2(_0643_));
 sg13g2_nand2_1 _1634_ (.Y(_0644_),
    .A(net143),
    .B(_0514_));
 sg13g2_xor2_1 _1635_ (.B(_0359_),
    .A(net143),
    .X(_0645_));
 sg13g2_o21ai_1 _1636_ (.B1(_0644_),
    .Y(_0078_),
    .A1(_0642_),
    .A2(_0645_));
 sg13g2_and2_1 _1637_ (.A(_0360_),
    .B(_0512_),
    .X(_0646_));
 sg13g2_o21ai_1 _1638_ (.B1(net156),
    .Y(_0647_),
    .A1(net351),
    .A2(_0646_));
 sg13g2_a21oi_1 _1639_ (.A1(net351),
    .A2(_0646_),
    .Y(_0079_),
    .B1(_0647_));
 sg13g2_a21oi_1 _1640_ (.A1(_0367_),
    .A2(_0512_),
    .Y(_0648_),
    .B1(net484));
 sg13g2_and3_2 _1641_ (.X(_0649_),
    .A(_0360_),
    .B(_0361_),
    .C(_0512_));
 sg13g2_nor3_1 _1642_ (.A(net154),
    .B(_0648_),
    .C(_0649_),
    .Y(_0080_));
 sg13g2_xnor2_1 _1643_ (.Y(_0650_),
    .A(net477),
    .B(_0649_));
 sg13g2_nor2_1 _1644_ (.A(net154),
    .B(_0650_),
    .Y(_0081_));
 sg13g2_a21oi_1 _1645_ (.A1(net477),
    .A2(_0649_),
    .Y(_0651_),
    .B1(net492));
 sg13g2_and2_1 _1646_ (.A(_0362_),
    .B(_0512_),
    .X(_0652_));
 sg13g2_nor3_1 _1647_ (.A(net154),
    .B(_0651_),
    .C(_0652_),
    .Y(_0082_));
 sg13g2_xnor2_1 _1648_ (.Y(_0653_),
    .A(net396),
    .B(_0652_));
 sg13g2_nor2_1 _1649_ (.A(net154),
    .B(_0653_),
    .Y(_0083_));
 sg13g2_nand2_1 _1650_ (.Y(_0654_),
    .A(net353),
    .B(_0514_));
 sg13g2_nand2_1 _1651_ (.Y(_0655_),
    .A(net396),
    .B(_0362_));
 sg13g2_xor2_1 _1652_ (.B(_0655_),
    .A(net353),
    .X(_0656_));
 sg13g2_o21ai_1 _1653_ (.B1(_0654_),
    .Y(_0084_),
    .A1(_0642_),
    .A2(_0656_));
 sg13g2_a21oi_1 _1654_ (.A1(_0253_),
    .A2(_0566_),
    .Y(_0085_),
    .B1(net152));
 sg13g2_nor3_1 _1655_ (.A(_0234_),
    .B(_0575_),
    .C(_0579_),
    .Y(_0657_));
 sg13g2_and2_1 _1656_ (.A(\game_inst.apple_inst.apple_x[0] ),
    .B(\game_inst.apple_inst.apple_x[1] ),
    .X(_0658_));
 sg13g2_nor3_1 _1657_ (.A(\game_inst.apple_inst.apple_x[2] ),
    .B(\game_inst.apple_inst.apple_x[3] ),
    .C(_0658_),
    .Y(_0659_));
 sg13g2_nand3_1 _1658_ (.B(\game_inst.apple_inst.apple_y[2] ),
    .C(\game_inst.apple_inst.apple_y[3] ),
    .A(net582),
    .Y(_0660_));
 sg13g2_o21ai_1 _1659_ (.B1(_0660_),
    .Y(_0661_),
    .A1(_0264_),
    .A2(_0659_));
 sg13g2_nor4_2 _1660_ (.A(net152),
    .B(_0582_),
    .C(_0657_),
    .Y(_0662_),
    .D(_0661_));
 sg13g2_nor2_1 _1661_ (.A(net406),
    .B(net110),
    .Y(_0663_));
 sg13g2_a21oi_1 _1662_ (.A1(_0259_),
    .A2(net110),
    .Y(_0086_),
    .B1(_0663_));
 sg13g2_nand2_1 _1663_ (.Y(_0664_),
    .A(net437),
    .B(net111));
 sg13g2_o21ai_1 _1664_ (.B1(_0664_),
    .Y(_0087_),
    .A1(_0246_),
    .A2(net110));
 sg13g2_nand2_1 _1665_ (.Y(_0665_),
    .A(net425),
    .B(net111));
 sg13g2_o21ai_1 _1666_ (.B1(_0665_),
    .Y(_0088_),
    .A1(_0245_),
    .A2(net110));
 sg13g2_nand2_1 _1667_ (.Y(_0666_),
    .A(net446),
    .B(net111));
 sg13g2_o21ai_1 _1668_ (.B1(_0666_),
    .Y(_0089_),
    .A1(_0244_),
    .A2(net111));
 sg13g2_nor2_1 _1669_ (.A(net426),
    .B(net110),
    .Y(_0667_));
 sg13g2_a21oi_1 _1670_ (.A1(_0264_),
    .A2(net110),
    .Y(_0090_),
    .B1(_0667_));
 sg13g2_a21oi_1 _1671_ (.A1(net381),
    .A2(_0340_),
    .Y(_0668_),
    .B1(\game_inst.apple_inst.o_ready ));
 sg13g2_nor2b_1 _1672_ (.A(net382),
    .B_N(net112),
    .Y(_0091_));
 sg13g2_o21ai_1 _1673_ (.B1(net112),
    .Y(_0669_),
    .A1(net381),
    .A2(net429));
 sg13g2_inv_1 _1674_ (.Y(_0092_),
    .A(_0669_));
 sg13g2_nor2_1 _1675_ (.A(net4),
    .B(net3),
    .Y(_0670_));
 sg13g2_nor3_1 _1676_ (.A(\game_inst.control_inst.i_head_dir[0] ),
    .B(net4),
    .C(net3),
    .Y(_0671_));
 sg13g2_o21ai_1 _1677_ (.B1(net1),
    .Y(_0672_),
    .A1(net485),
    .A2(_0671_));
 sg13g2_a21oi_1 _1678_ (.A1(net468),
    .A2(_0670_),
    .Y(_0673_),
    .B1(net485));
 sg13g2_nor2b_1 _1679_ (.A(_0673_),
    .B_N(net2),
    .Y(_0674_));
 sg13g2_nand2b_1 _1680_ (.Y(_0675_),
    .B(net2),
    .A_N(_0673_));
 sg13g2_o21ai_1 _1681_ (.B1(\game_inst.control_inst.backwards[1] ),
    .Y(_0676_),
    .A1(net2),
    .A2(net1));
 sg13g2_nand2_1 _1682_ (.Y(_0677_),
    .A(\game_inst.control_inst.backwards[1] ),
    .B(\game_inst.control_inst.i_head_dir[0] ));
 sg13g2_and3_1 _1683_ (.X(_0678_),
    .A(net3),
    .B(_0676_),
    .C(_0677_));
 sg13g2_nand2b_1 _1684_ (.Y(_0679_),
    .B(\game_inst.control_inst.backwards[1] ),
    .A_N(\game_inst.control_inst.i_head_dir[0] ));
 sg13g2_nand3_1 _1685_ (.B(_0676_),
    .C(_0679_),
    .A(net4),
    .Y(_0680_));
 sg13g2_a21oi_1 _1686_ (.A1(_0240_),
    .A2(_0680_),
    .Y(_0681_),
    .B1(_0678_));
 sg13g2_o21ai_1 _1687_ (.B1(_0672_),
    .Y(_0682_),
    .A1(_0674_),
    .A2(_0681_));
 sg13g2_and2_1 _1688_ (.A(_0672_),
    .B(_0675_),
    .X(_0683_));
 sg13g2_nand2b_1 _1689_ (.Y(_0684_),
    .B(_0680_),
    .A_N(_0678_));
 sg13g2_nor2_1 _1690_ (.A(net141),
    .B(_0684_),
    .Y(_0685_));
 sg13g2_nand2b_1 _1691_ (.Y(_0686_),
    .B(_0683_),
    .A_N(_0685_));
 sg13g2_a21o_1 _1692_ (.A2(_0683_),
    .A1(\game_inst.control_inst.dir[1] ),
    .B1(_0685_),
    .X(_0687_));
 sg13g2_xnor2_1 _1693_ (.Y(_0688_),
    .A(_0240_),
    .B(_0682_));
 sg13g2_a21o_1 _1694_ (.A2(_0688_),
    .A1(_0687_),
    .B1(net419),
    .X(_0689_));
 sg13g2_nand3_1 _1695_ (.B(_0687_),
    .C(_0688_),
    .A(net419),
    .Y(_0690_));
 sg13g2_nand3_1 _1696_ (.B(_0689_),
    .C(_0690_),
    .A(net112),
    .Y(_0691_));
 sg13g2_xor2_1 _1697_ (.B(net417),
    .A(\game_inst.apple_inst.random_inst.lfsr5[4] ),
    .X(_0692_));
 sg13g2_a21oi_1 _1698_ (.A1(net108),
    .A2(net418),
    .Y(_0693_),
    .B1(net155));
 sg13g2_o21ai_1 _1699_ (.B1(_0693_),
    .Y(_0093_),
    .A1(_0247_),
    .A2(net109));
 sg13g2_a21oi_1 _1700_ (.A1(net406),
    .A2(net109),
    .Y(_0694_),
    .B1(net155));
 sg13g2_o21ai_1 _1701_ (.B1(_0694_),
    .Y(_0094_),
    .A1(_0246_),
    .A2(net108));
 sg13g2_a21oi_1 _1702_ (.A1(net416),
    .A2(net108),
    .Y(_0695_),
    .B1(net155));
 sg13g2_o21ai_1 _1703_ (.B1(_0695_),
    .Y(_0095_),
    .A1(_0245_),
    .A2(net108));
 sg13g2_o21ai_1 _1704_ (.B1(net157),
    .Y(_0696_),
    .A1(net397),
    .A2(net108));
 sg13g2_a21oi_1 _1705_ (.A1(_0245_),
    .A2(net108),
    .Y(_0096_),
    .B1(_0696_));
 sg13g2_o21ai_1 _1706_ (.B1(net157),
    .Y(_0697_),
    .A1(\game_inst.apple_inst.random_inst.lfsr5[4] ),
    .A2(net108));
 sg13g2_a21oi_1 _1707_ (.A1(_0244_),
    .A2(net108),
    .Y(_0097_),
    .B1(_0697_));
 sg13g2_a21o_1 _1708_ (.A2(net109),
    .A1(net458),
    .B1(_0243_),
    .X(_0698_));
 sg13g2_nand3_1 _1709_ (.B(_0243_),
    .C(net109),
    .A(net458),
    .Y(_0699_));
 sg13g2_nand3_1 _1710_ (.B(_0698_),
    .C(_0699_),
    .A(net157),
    .Y(_0098_));
 sg13g2_o21ai_1 _1711_ (.B1(net157),
    .Y(_0700_),
    .A1(_0242_),
    .A2(net109));
 sg13g2_a21o_1 _1712_ (.A2(net109),
    .A1(net375),
    .B1(_0700_),
    .X(_0099_));
 sg13g2_o21ai_1 _1713_ (.B1(net157),
    .Y(_0701_),
    .A1(net415),
    .A2(_0691_));
 sg13g2_a21oi_1 _1714_ (.A1(_0242_),
    .A2(net109),
    .Y(_0100_),
    .B1(_0701_));
 sg13g2_a21oi_1 _1715_ (.A1(net415),
    .A2(_0691_),
    .Y(_0702_),
    .B1(net155));
 sg13g2_o21ai_1 _1716_ (.B1(_0702_),
    .Y(_0101_),
    .A1(_0241_),
    .A2(_0691_));
 sg13g2_a21o_1 _1717_ (.A2(net121),
    .A1(net468),
    .B1(_0494_),
    .X(_0102_));
 sg13g2_a21o_1 _1718_ (.A2(net122),
    .A1(net485),
    .B1(_0497_),
    .X(_0103_));
 sg13g2_nand2_1 _1719_ (.Y(_0703_),
    .A(net500),
    .B(net119));
 sg13g2_nor2_2 _1720_ (.A(net141),
    .B(net119),
    .Y(_0704_));
 sg13g2_nor3_1 _1721_ (.A(_0238_),
    .B(net141),
    .C(net119),
    .Y(_0705_));
 sg13g2_nor2_1 _1722_ (.A(net500),
    .B(_0496_),
    .Y(_0706_));
 sg13g2_nor2_1 _1723_ (.A(_0705_),
    .B(_0706_),
    .Y(_0707_));
 sg13g2_a21oi_1 _1724_ (.A1(_0703_),
    .A2(_0707_),
    .Y(_0104_),
    .B1(net151));
 sg13g2_nand2_2 _1725_ (.Y(_0708_),
    .A(net141),
    .B(\game_inst.control_inst.dir[0] ));
 sg13g2_and2_1 _1726_ (.A(\game_inst.head_x[1] ),
    .B(_0708_),
    .X(_0709_));
 sg13g2_xor2_1 _1727_ (.B(_0708_),
    .A(\game_inst.head_x[1] ),
    .X(_0710_));
 sg13g2_xnor2_1 _1728_ (.Y(_0711_),
    .A(_0238_),
    .B(_0710_));
 sg13g2_a22oi_1 _1729_ (.Y(_0712_),
    .B1(_0711_),
    .B2(_0495_),
    .A2(_0704_),
    .A1(net531));
 sg13g2_dfrbpq_2 _1730_ (.RESET_B(net28),
    .D(_0039_),
    .Q(\game_inst.snake_inst.pos[0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _1731_ (.RESET_B(net176),
    .D(_0040_),
    .Q(\game_inst.snake_inst.pos[3] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _1732_ (.RESET_B(net175),
    .D(_0041_),
    .Q(\game_inst.snake_inst.pos[5] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _1733_ (.RESET_B(net174),
    .D(net510),
    .Q(\game_inst.snake_inst.pos[6] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _1734_ (.RESET_B(net173),
    .D(_0043_),
    .Q(\game_inst.snake_inst.pos[7] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _1735_ (.RESET_B(net172),
    .D(_0044_),
    .Q(\game_inst.vga_inst.px[0] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1736_ (.RESET_B(net171),
    .D(_0045_),
    .Q(\game_inst.vga_inst.px[1] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1737_ (.RESET_B(net170),
    .D(net385),
    .Q(\game_inst.vga_inst.px[2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1738_ (.RESET_B(net169),
    .D(_0047_),
    .Q(\game_inst.vga_inst.px[3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1739_ (.RESET_B(net168),
    .D(_0048_),
    .Q(\game_inst.vga_inst.px[4] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _1740_ (.RESET_B(net167),
    .D(_0049_),
    .Q(\game_inst.vga_inst.px[5] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _1741_ (.RESET_B(net166),
    .D(_0050_),
    .Q(\game_inst.vga_inst.px[6] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _1742_ (.RESET_B(net165),
    .D(_0051_),
    .Q(\game_inst.vga_inst.px[7] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _1743_ (.RESET_B(net164),
    .D(_0052_),
    .Q(\game_inst.vga_inst.px[8] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _1744_ (.RESET_B(net29),
    .D(_0053_),
    .Q(\game_inst.vga_inst.px[9] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _1745_ (.RESET_B(net30),
    .D(_0000_),
    .Q(\game_inst.vga_inst.color[1] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _1746_ (.RESET_B(net47),
    .D(_0001_),
    .Q(\game_inst.vga_inst.color[2] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _1747_ (.RESET_B(net163),
    .D(net347),
    .Q(\game_inst.vga_inst.color[3] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _1748_ (.RESET_B(net162),
    .D(_0054_),
    .Q(\game_inst.sound_inst.max_counter[2] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _1749_ (.RESET_B(net160),
    .D(net577),
    .Q(\game_inst.sound_inst.max_counter[1] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _1750_ (.RESET_B(net158),
    .D(net365),
    .Q(audio),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _1751_ (.RESET_B(net106),
    .D(net434),
    .Q(\game_inst.sound_inst.mode[0] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _1752_ (.RESET_B(net104),
    .D(_0058_),
    .Q(\game_inst.sound_inst.mode[1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _1753_ (.RESET_B(net102),
    .D(net424),
    .Q(\game_inst.sound_inst.counter[0] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _1754_ (.RESET_B(net99),
    .D(_0060_),
    .Q(\game_inst.sound_inst.counter[1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _1755_ (.RESET_B(net97),
    .D(_0061_),
    .Q(\game_inst.sound_inst.counter[2] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _1756_ (.RESET_B(net95),
    .D(_0062_),
    .Q(\game_inst.sound_inst.counter[3] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _1757_ (.RESET_B(net93),
    .D(_0063_),
    .Q(\game_inst.sound_inst.max_counter[0] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _1758_ (.RESET_B(net91),
    .D(net525),
    .Q(\game_inst.sound_inst.max_counter[3] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _1759_ (.RESET_B(net88),
    .D(net472),
    .Q(\game_inst.sound_inst.phase[0] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _1760_ (.RESET_B(net86),
    .D(net392),
    .Q(\game_inst.sound_inst.phase[1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _1761_ (.RESET_B(net46),
    .D(_0067_),
    .Q(\game_inst.sound_inst.phase[2] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _1762_ (.RESET_B(net44),
    .D(_0068_),
    .Q(\game_inst.sound_inst.phase[3] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _1763_ (.RESET_B(net48),
    .D(_0069_),
    .Q(\game_inst.sound_inst.phase[4] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _1764_ (.RESET_B(net49),
    .D(net341),
    .Q(\game_inst.sound_inst.prev_pwm_base ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _1765_ (.RESET_B(net50),
    .D(\game_inst.sound_inst.vsync_pulse ),
    .Q(\game_inst.sound_inst.prev_vsync ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _1766_ (.RESET_B(net51),
    .D(net339),
    .Q(\game_inst.o_vga_hsync ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _1767_ (.RESET_B(net52),
    .D(net340),
    .Q(\game_inst.o_vga_vsync ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _1768_ (.RESET_B(net53),
    .D(_0038_),
    .Q(\game_inst.vga_inst.prev_dir[0] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _1769_ (.RESET_B(net54),
    .D(net135),
    .Q(\game_inst.vga_inst.prev_dir[1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1770_ (.RESET_B(net55),
    .D(_0032_),
    .Q(\game_inst.vga_inst.row_buffer[8][0] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _1771_ (.RESET_B(net56),
    .D(_0033_),
    .Q(\game_inst.vga_inst.row_buffer[8][1] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _1772_ (.RESET_B(net58),
    .D(_0034_),
    .Q(\game_inst.vga_inst.row_buffer[8][2] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1773_ (.RESET_B(net42),
    .D(_0035_),
    .Q(\game_inst.vga_inst.row_buffer[8][3] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _1774_ (.RESET_B(net59),
    .D(net405),
    .Q(\game_inst.o_tick ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _1775_ (.RESET_B(net60),
    .D(_0004_),
    .Q(\game_inst.vga_inst.row_buffer[1][0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1776_ (.RESET_B(net61),
    .D(net546),
    .Q(\game_inst.vga_inst.row_buffer[1][1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1777_ (.RESET_B(net62),
    .D(net563),
    .Q(\game_inst.vga_inst.row_buffer[1][2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1778_ (.RESET_B(net63),
    .D(net561),
    .Q(\game_inst.vga_inst.row_buffer[1][3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1779_ (.RESET_B(net64),
    .D(net541),
    .Q(\game_inst.vga_inst.row_buffer[2][0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1780_ (.RESET_B(net65),
    .D(_0009_),
    .Q(\game_inst.vga_inst.row_buffer[2][1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1781_ (.RESET_B(net66),
    .D(net559),
    .Q(\game_inst.vga_inst.row_buffer[2][2] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _1782_ (.RESET_B(net67),
    .D(net552),
    .Q(\game_inst.vga_inst.row_buffer[2][3] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1783_ (.RESET_B(net68),
    .D(_0012_),
    .Q(\game_inst.vga_inst.row_buffer[3][0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1784_ (.RESET_B(net69),
    .D(net537),
    .Q(\game_inst.vga_inst.row_buffer[3][1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1785_ (.RESET_B(net70),
    .D(net544),
    .Q(\game_inst.vga_inst.row_buffer[3][2] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _1786_ (.RESET_B(net71),
    .D(_0015_),
    .Q(\game_inst.vga_inst.row_buffer[3][3] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1787_ (.RESET_B(net72),
    .D(_0016_),
    .Q(\game_inst.vga_inst.row_buffer[4][0] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _1788_ (.RESET_B(net73),
    .D(_0017_),
    .Q(\game_inst.vga_inst.row_buffer[4][1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1789_ (.RESET_B(net74),
    .D(_0018_),
    .Q(\game_inst.vga_inst.row_buffer[4][2] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _1790_ (.RESET_B(net75),
    .D(_0019_),
    .Q(\game_inst.vga_inst.row_buffer[4][3] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1791_ (.RESET_B(net76),
    .D(_0020_),
    .Q(\game_inst.vga_inst.row_buffer[5][0] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1792_ (.RESET_B(net77),
    .D(_0021_),
    .Q(\game_inst.vga_inst.row_buffer[5][1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1793_ (.RESET_B(net78),
    .D(_0022_),
    .Q(\game_inst.vga_inst.row_buffer[5][2] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1794_ (.RESET_B(net79),
    .D(_0023_),
    .Q(\game_inst.vga_inst.row_buffer[5][3] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1795_ (.RESET_B(net80),
    .D(net371),
    .Q(\game_inst.vga_inst.row_buffer[6][0] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _1796_ (.RESET_B(net81),
    .D(net374),
    .Q(\game_inst.vga_inst.row_buffer[6][1] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _1797_ (.RESET_B(net82),
    .D(net362),
    .Q(\game_inst.vga_inst.row_buffer[6][2] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1798_ (.RESET_B(net83),
    .D(net368),
    .Q(\game_inst.vga_inst.row_buffer[6][3] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1799_ (.RESET_B(net84),
    .D(_0028_),
    .Q(\game_inst.vga_inst.row_buffer[7][0] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _1800_ (.RESET_B(net85),
    .D(_0029_),
    .Q(\game_inst.vga_inst.row_buffer[7][1] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _1801_ (.RESET_B(net90),
    .D(net414),
    .Q(\game_inst.vga_inst.row_buffer[7][2] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1802_ (.RESET_B(net40),
    .D(_0031_),
    .Q(\game_inst.vga_inst.row_buffer[7][3] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1803_ (.RESET_B(net39),
    .D(net456),
    .Q(\game_inst.vga_inst.row_buffer[0][0] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _1804_ (.RESET_B(net38),
    .D(net440),
    .Q(\game_inst.vga_inst.row_buffer[0][1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _1805_ (.RESET_B(net37),
    .D(net445),
    .Q(\game_inst.vga_inst.row_buffer[0][2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1806_ (.RESET_B(net101),
    .D(net448),
    .Q(\game_inst.vga_inst.row_buffer[0][3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1807_ (.RESET_B(net36),
    .D(net474),
    .Q(\game_inst.vga_inst.s_hsync ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _1808_ (.RESET_B(net35),
    .D(_0075_),
    .Q(\game_inst.vga_inst.py[0] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _1809_ (.RESET_B(net33),
    .D(net421),
    .Q(\game_inst.vga_inst.py[1] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _1810_ (.RESET_B(net31),
    .D(_0077_),
    .Q(\game_inst.vga_inst.py[2] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _1811_ (.RESET_B(net26),
    .D(_0078_),
    .Q(\game_inst.pwm_base ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _1812_ (.RESET_B(net24),
    .D(_0079_),
    .Q(\game_inst.vga_inst.py[4] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _1813_ (.RESET_B(net22),
    .D(_0080_),
    .Q(\game_inst.vga_inst.py[5] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _1814_ (.RESET_B(net20),
    .D(_0081_),
    .Q(\game_inst.vga_inst.py[6] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _1815_ (.RESET_B(net18),
    .D(_0082_),
    .Q(\game_inst.vga_inst.py[7] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _1816_ (.RESET_B(net16),
    .D(_0083_),
    .Q(\game_inst.vga_inst.py[8] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _1817_ (.RESET_B(net216),
    .D(_0084_),
    .Q(\game_inst.vga_inst.py[9] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _1818_ (.RESET_B(net14),
    .D(net354),
    .Q(\game_inst.vga_inst.s_vsync ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _1819_ (.RESET_B(net215),
    .D(_0085_),
    .Q(failure),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _1820_ (.RESET_B(net214),
    .D(net407),
    .Q(\game_inst.apple_inst.apple_x[0] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _1821_ (.RESET_B(net213),
    .D(_0087_),
    .Q(\game_inst.apple_inst.apple_x[1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _1822_ (.RESET_B(net212),
    .D(_0088_),
    .Q(\game_inst.apple_inst.apple_x[2] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _1823_ (.RESET_B(net211),
    .D(_0089_),
    .Q(\game_inst.apple_inst.apple_x[3] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _1824_ (.RESET_B(net210),
    .D(net427),
    .Q(\game_inst.apple_inst.apple_x[4] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _1825_ (.RESET_B(net209),
    .D(_0091_),
    .Q(\game_inst.apple_inst.o_ready ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _1826_ (.RESET_B(net207),
    .D(_0092_),
    .Q(\game_inst.apple_inst.test ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _1827_ (.RESET_B(net205),
    .D(_0093_),
    .Q(\game_inst.apple_inst.random_inst.lfsr5[0] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _1828_ (.RESET_B(net203),
    .D(_0094_),
    .Q(\game_inst.apple_inst.random_inst.lfsr5[1] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _1829_ (.RESET_B(net201),
    .D(_0095_),
    .Q(\game_inst.apple_inst.random_inst.lfsr5[2] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _1830_ (.RESET_B(net199),
    .D(_0096_),
    .Q(\game_inst.apple_inst.random_inst.lfsr5[3] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _1831_ (.RESET_B(net197),
    .D(net398),
    .Q(\game_inst.apple_inst.random_inst.lfsr5[4] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _1832_ (.RESET_B(net195),
    .D(_0098_),
    .Q(\game_inst.apple_inst.random_inst.lfsr4[0] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _1833_ (.RESET_B(net193),
    .D(net376),
    .Q(\game_inst.apple_inst.random_inst.lfsr4[1] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _1834_ (.RESET_B(net191),
    .D(_0100_),
    .Q(\game_inst.apple_inst.random_inst.lfsr4[2] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _1835_ (.RESET_B(net189),
    .D(_0101_),
    .Q(\game_inst.apple_inst.random_inst.lfsr4[3] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _1836_ (.RESET_B(net187),
    .D(net469),
    .Q(\game_inst.control_inst.i_head_dir[0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _1837_ (.RESET_B(net185),
    .D(net486),
    .Q(\game_inst.control_inst.backwards[1] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _1838_ (.RESET_B(net183),
    .D(net501),
    .Q(\game_inst.head_x[0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _1839_ (.RESET_B(net181),
    .D(net532),
    .Q(\game_inst.head_x[1] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _1840_ (.RESET_B(net179),
    .D(net504),
    .Q(\game_inst.head_x[2] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _1841_ (.RESET_B(net177),
    .D(net530),
    .Q(\game_inst.head_x[3] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _1842_ (.RESET_B(net159),
    .D(_0108_),
    .Q(\game_inst.head_x[4] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _1843_ (.RESET_B(net105),
    .D(net506),
    .Q(\game_inst.head_y[0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _1844_ (.RESET_B(net100),
    .D(_0110_),
    .Q(\game_inst.head_y[1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _1845_ (.RESET_B(net96),
    .D(_0111_),
    .Q(\game_inst.head_y[2] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _1846_ (.RESET_B(net92),
    .D(_0112_),
    .Q(\game_inst.head_y[3] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _1847_ (.RESET_B(net87),
    .D(_0113_),
    .Q(\game_inst.control_inst.dir[0] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _1848_ (.RESET_B(net57),
    .D(_0114_),
    .Q(\game_inst.control_inst.dir[1] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _1849_ (.RESET_B(net45),
    .D(_0115_),
    .Q(\game_inst.apple_inst.i_snake_x[0] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _1850_ (.RESET_B(net43),
    .D(_0116_),
    .Q(\game_inst.apple_inst.i_snake_x[1] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _1851_ (.RESET_B(net41),
    .D(_0117_),
    .Q(\game_inst.apple_inst.i_snake_x[2] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _1852_ (.RESET_B(net34),
    .D(_0118_),
    .Q(\game_inst.apple_inst.i_snake_x[3] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _1853_ (.RESET_B(net32),
    .D(_0119_),
    .Q(\game_inst.apple_inst.i_snake_x[4] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _1854_ (.RESET_B(net27),
    .D(_0120_),
    .Q(\game_inst.apple_inst.i_snake_valid ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _1855_ (.RESET_B(net23),
    .D(_0121_),
    .Q(\game_inst.apple_inst.i_snake_y[0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _1856_ (.RESET_B(net21),
    .D(_0122_),
    .Q(\game_inst.apple_inst.i_snake_y[1] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _1857_ (.RESET_B(net19),
    .D(net527),
    .Q(\game_inst.apple_inst.i_snake_y[2] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _1858_ (.RESET_B(net17),
    .D(net515),
    .Q(\game_inst.apple_inst.i_snake_y[3] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _1859_ (.RESET_B(net15),
    .D(_0125_),
    .Q(\game_inst.snake_inst.length[0] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _1860_ (.RESET_B(net13),
    .D(_0126_),
    .Q(\game_inst.snake_inst.length[1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _1861_ (.RESET_B(net208),
    .D(net496),
    .Q(\game_inst.snake_inst.length[2] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _1862_ (.RESET_B(net206),
    .D(net467),
    .Q(\game_inst.snake_inst.length[3] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _1863_ (.RESET_B(net204),
    .D(net452),
    .Q(\game_inst.snake_inst.length[4] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _1864_ (.RESET_B(net202),
    .D(_0130_),
    .Q(\game_inst.snake_inst.length[5] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _1865_ (.RESET_B(net200),
    .D(net412),
    .Q(\game_inst.snake_inst.length[6] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _1866_ (.RESET_B(net198),
    .D(net350),
    .Q(\game_inst.snake_inst.length[7] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _1867_ (.RESET_B(net196),
    .D(_0133_),
    .Q(\game_inst.snake_inst.pos[1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _1868_ (.RESET_B(net194),
    .D(net462),
    .Q(\game_inst.snake_inst.pos[2] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _1869_ (.RESET_B(net192),
    .D(net395),
    .Q(\game_inst.snake_inst.pos[4] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _1870_ (.RESET_B(net190),
    .D(_0136_),
    .Q(\game_inst.apple_inst.apple_y[0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _1871_ (.RESET_B(net188),
    .D(net389),
    .Q(\game_inst.apple_inst.apple_y[1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _1872_ (.RESET_B(net186),
    .D(_0138_),
    .Q(\game_inst.apple_inst.apple_y[2] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _1873_ (.RESET_B(net184),
    .D(net409),
    .Q(\game_inst.apple_inst.apple_y[3] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _1874_ (.RESET_B(net182),
    .D(_0140_),
    .Q(\game_inst.control_inst.o_start ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _1875_ (.RESET_B(net180),
    .D(net400),
    .Q(\game_inst.tickgen_inst.counter_max[1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _1876_ (.RESET_B(net161),
    .D(net489),
    .Q(\game_inst.tickgen_inst.counter_max[2] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _1877_ (.RESET_B(net103),
    .D(net513),
    .Q(\game_inst.tickgen_inst.counter_max[3] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _1878_ (.RESET_B(net94),
    .D(net403),
    .Q(\game_inst.tick ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _1879_ (.RESET_B(net25),
    .D(net358),
    .Q(\game_inst.tickgen_inst.counter[0] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _1880_ (.RESET_B(net107),
    .D(_0146_),
    .Q(\game_inst.tickgen_inst.counter[1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _1881_ (.RESET_B(net89),
    .D(_0147_),
    .Q(\game_inst.tickgen_inst.counter[2] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _1882_ (.RESET_B(net178),
    .D(net345),
    .Q(\game_inst.tickgen_inst.counter[3] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _1883_ (.RESET_B(net98),
    .D(_0003_),
    .Q(\game_inst.tickgen_inst.prev_user_input ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_tiehi _1818__14 (.L_HI(net14));
 sg13g2_tiehi _1859__15 (.L_HI(net15));
 sg13g2_tiehi _1816__16 (.L_HI(net16));
 sg13g2_tiehi _1858__17 (.L_HI(net17));
 sg13g2_tiehi _1815__18 (.L_HI(net18));
 sg13g2_tiehi _1857__19 (.L_HI(net19));
 sg13g2_tiehi _1814__20 (.L_HI(net20));
 sg13g2_tiehi _1856__21 (.L_HI(net21));
 sg13g2_tiehi _1813__22 (.L_HI(net22));
 sg13g2_tiehi _1855__23 (.L_HI(net23));
 sg13g2_tiehi _1812__24 (.L_HI(net24));
 sg13g2_tiehi _1879__25 (.L_HI(net25));
 sg13g2_tiehi _1811__26 (.L_HI(net26));
 sg13g2_tiehi _1854__27 (.L_HI(net27));
 sg13g2_tiehi _1730__28 (.L_HI(net28));
 sg13g2_tiehi _1744__29 (.L_HI(net29));
 sg13g2_tiehi _1745__30 (.L_HI(net30));
 sg13g2_tiehi _1810__31 (.L_HI(net31));
 sg13g2_tiehi _1853__32 (.L_HI(net32));
 sg13g2_tiehi _1809__33 (.L_HI(net33));
 sg13g2_tiehi _1852__34 (.L_HI(net34));
 sg13g2_tiehi _1808__35 (.L_HI(net35));
 sg13g2_tiehi _1807__36 (.L_HI(net36));
 sg13g2_tiehi _1805__37 (.L_HI(net37));
 sg13g2_tiehi _1804__38 (.L_HI(net38));
 sg13g2_tiehi _1803__39 (.L_HI(net39));
 sg13g2_tiehi _1802__40 (.L_HI(net40));
 sg13g2_tiehi _1851__41 (.L_HI(net41));
 sg13g2_tiehi _1773__42 (.L_HI(net42));
 sg13g2_tiehi _1850__43 (.L_HI(net43));
 sg13g2_tiehi _1762__44 (.L_HI(net44));
 sg13g2_tiehi _1849__45 (.L_HI(net45));
 sg13g2_tiehi _1761__46 (.L_HI(net46));
 sg13g2_tiehi _1746__47 (.L_HI(net47));
 sg13g2_tiehi _1763__48 (.L_HI(net48));
 sg13g2_tiehi _1764__49 (.L_HI(net49));
 sg13g2_tiehi _1765__50 (.L_HI(net50));
 sg13g2_tiehi _1766__51 (.L_HI(net51));
 sg13g2_tiehi _1767__52 (.L_HI(net52));
 sg13g2_tiehi _1768__53 (.L_HI(net53));
 sg13g2_tiehi _1769__54 (.L_HI(net54));
 sg13g2_tiehi _1770__55 (.L_HI(net55));
 sg13g2_tiehi _1771__56 (.L_HI(net56));
 sg13g2_tiehi _1848__57 (.L_HI(net57));
 sg13g2_tiehi _1772__58 (.L_HI(net58));
 sg13g2_tiehi _1774__59 (.L_HI(net59));
 sg13g2_tiehi _1775__60 (.L_HI(net60));
 sg13g2_tiehi _1776__61 (.L_HI(net61));
 sg13g2_tiehi _1777__62 (.L_HI(net62));
 sg13g2_tiehi _1778__63 (.L_HI(net63));
 sg13g2_tiehi _1779__64 (.L_HI(net64));
 sg13g2_tiehi _1780__65 (.L_HI(net65));
 sg13g2_tiehi _1781__66 (.L_HI(net66));
 sg13g2_tiehi _1782__67 (.L_HI(net67));
 sg13g2_tiehi _1783__68 (.L_HI(net68));
 sg13g2_tiehi _1784__69 (.L_HI(net69));
 sg13g2_tiehi _1785__70 (.L_HI(net70));
 sg13g2_tiehi _1786__71 (.L_HI(net71));
 sg13g2_tiehi _1787__72 (.L_HI(net72));
 sg13g2_tiehi _1788__73 (.L_HI(net73));
 sg13g2_tiehi _1789__74 (.L_HI(net74));
 sg13g2_tiehi _1790__75 (.L_HI(net75));
 sg13g2_tiehi _1791__76 (.L_HI(net76));
 sg13g2_tiehi _1792__77 (.L_HI(net77));
 sg13g2_tiehi _1793__78 (.L_HI(net78));
 sg13g2_tiehi _1794__79 (.L_HI(net79));
 sg13g2_tiehi _1795__80 (.L_HI(net80));
 sg13g2_tiehi _1796__81 (.L_HI(net81));
 sg13g2_tiehi _1797__82 (.L_HI(net82));
 sg13g2_tiehi _1798__83 (.L_HI(net83));
 sg13g2_tiehi _1799__84 (.L_HI(net84));
 sg13g2_tiehi _1800__85 (.L_HI(net85));
 sg13g2_tiehi _1760__86 (.L_HI(net86));
 sg13g2_tiehi _1847__87 (.L_HI(net87));
 sg13g2_tiehi _1759__88 (.L_HI(net88));
 sg13g2_tiehi _1881__89 (.L_HI(net89));
 sg13g2_tiehi _1801__90 (.L_HI(net90));
 sg13g2_tiehi _1758__91 (.L_HI(net91));
 sg13g2_tiehi _1846__92 (.L_HI(net92));
 sg13g2_tiehi _1757__93 (.L_HI(net93));
 sg13g2_tiehi _1878__94 (.L_HI(net94));
 sg13g2_tiehi _1756__95 (.L_HI(net95));
 sg13g2_tiehi _1845__96 (.L_HI(net96));
 sg13g2_tiehi _1755__97 (.L_HI(net97));
 sg13g2_tiehi _1883__98 (.L_HI(net98));
 sg13g2_tiehi _1754__99 (.L_HI(net99));
 sg13g2_tiehi _1844__100 (.L_HI(net100));
 sg13g2_tiehi _1806__101 (.L_HI(net101));
 sg13g2_tiehi _1753__102 (.L_HI(net102));
 sg13g2_tiehi _1877__103 (.L_HI(net103));
 sg13g2_tiehi _1752__104 (.L_HI(net104));
 sg13g2_tiehi _1843__105 (.L_HI(net105));
 sg13g2_tiehi _1751__106 (.L_HI(net106));
 sg13g2_tiehi _1880__107 (.L_HI(net107));
 sg13g2_tiehi _1750__108 (.L_HI(net158));
 sg13g2_tiehi _1842__109 (.L_HI(net159));
 sg13g2_tiehi _1749__110 (.L_HI(net160));
 sg13g2_tiehi _1876__111 (.L_HI(net161));
 sg13g2_tiehi _1748__112 (.L_HI(net162));
 sg13g2_tiehi _1747__113 (.L_HI(net163));
 sg13g2_tiehi _1743__114 (.L_HI(net164));
 sg13g2_tiehi _1742__115 (.L_HI(net165));
 sg13g2_tiehi _1741__116 (.L_HI(net166));
 sg13g2_tiehi _1740__117 (.L_HI(net167));
 sg13g2_tiehi _1739__118 (.L_HI(net168));
 sg13g2_tiehi _1738__119 (.L_HI(net169));
 sg13g2_tiehi _1737__120 (.L_HI(net170));
 sg13g2_tiehi _1736__121 (.L_HI(net171));
 sg13g2_tiehi _1735__122 (.L_HI(net172));
 sg13g2_tiehi _1734__123 (.L_HI(net173));
 sg13g2_tiehi _1733__124 (.L_HI(net174));
 sg13g2_tiehi _1732__125 (.L_HI(net175));
 sg13g2_tiehi _1731__126 (.L_HI(net176));
 sg13g2_tiehi _1841__127 (.L_HI(net177));
 sg13g2_tiehi _1882__128 (.L_HI(net178));
 sg13g2_tiehi _1840__129 (.L_HI(net179));
 sg13g2_tiehi _1875__130 (.L_HI(net180));
 sg13g2_tiehi _1839__131 (.L_HI(net181));
 sg13g2_tiehi _1874__132 (.L_HI(net182));
 sg13g2_tiehi _1838__133 (.L_HI(net183));
 sg13g2_tiehi _1873__134 (.L_HI(net184));
 sg13g2_tiehi _1837__135 (.L_HI(net185));
 sg13g2_tiehi _1872__136 (.L_HI(net186));
 sg13g2_tiehi _1836__137 (.L_HI(net187));
 sg13g2_tiehi _1871__138 (.L_HI(net188));
 sg13g2_tiehi _1835__139 (.L_HI(net189));
 sg13g2_tiehi _1870__140 (.L_HI(net190));
 sg13g2_tiehi _1834__141 (.L_HI(net191));
 sg13g2_tiehi _1869__142 (.L_HI(net192));
 sg13g2_tiehi _1833__143 (.L_HI(net193));
 sg13g2_tiehi _1868__144 (.L_HI(net194));
 sg13g2_tiehi _1832__145 (.L_HI(net195));
 sg13g2_tiehi _1867__146 (.L_HI(net196));
 sg13g2_tiehi _1831__147 (.L_HI(net197));
 sg13g2_tiehi _1866__148 (.L_HI(net198));
 sg13g2_tiehi _1830__149 (.L_HI(net199));
 sg13g2_tiehi _1865__150 (.L_HI(net200));
 sg13g2_tiehi _1829__151 (.L_HI(net201));
 sg13g2_tiehi _1864__152 (.L_HI(net202));
 sg13g2_tiehi _1828__153 (.L_HI(net203));
 sg13g2_tiehi _1863__154 (.L_HI(net204));
 sg13g2_tiehi _1827__155 (.L_HI(net205));
 sg13g2_tiehi _1862__156 (.L_HI(net206));
 sg13g2_tiehi _1826__157 (.L_HI(net207));
 sg13g2_tiehi _1861__158 (.L_HI(net208));
 sg13g2_tiehi _1825__159 (.L_HI(net209));
 sg13g2_tiehi _1824__160 (.L_HI(net210));
 sg13g2_tiehi _1823__161 (.L_HI(net211));
 sg13g2_tiehi _1822__162 (.L_HI(net212));
 sg13g2_tiehi _1821__163 (.L_HI(net213));
 sg13g2_tiehi _1820__164 (.L_HI(net214));
 sg13g2_tiehi _1819__165 (.L_HI(net215));
 sg13g2_tiehi _1817__166 (.L_HI(net216));
 sg13g2_tiehi tt_um_snake_game_167 (.L_HI(net217));
 sg13g2_tiehi tt_um_snake_game_168 (.L_HI(net218));
 sg13g2_tiehi tt_um_snake_game_169 (.L_HI(net219));
 sg13g2_tiehi tt_um_snake_game_170 (.L_HI(net220));
 sg13g2_tiehi tt_um_snake_game_171 (.L_HI(net221));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[0].sreg_bufhigh_172  (.L_HI(net222));
 sg13g2_tielo tt_um_snake_game_8 (.L_LO(net8));
 sg13g2_tielo tt_um_snake_game_9 (.L_LO(net9));
 sg13g2_tielo tt_um_snake_game_10 (.L_LO(net10));
 sg13g2_tielo tt_um_snake_game_11 (.L_LO(net11));
 sg13g2_tielo tt_um_snake_game_12 (.L_LO(net12));
 sg13g2_tiehi _1860__13 (.L_HI(net13));
 sg13g2_buf_1 _2049_ (.A(failure),
    .X(uio_out[0]));
 sg13g2_buf_1 _2050_ (.A(\game_inst.o_success ),
    .X(uio_out[1]));
 sg13g2_buf_1 _2051_ (.A(eat),
    .X(uio_out[2]));
 sg13g2_buf_1 _2052_ (.A(\game_inst.o_tick ),
    .X(uio_out[3]));
 sg13g2_buf_1 _2053_ (.A(audio),
    .X(uio_out[7]));
 sg13g2_buf_1 _2054_ (.A(uo_out[4]),
    .X(uo_out[0]));
 sg13g2_buf_1 _2055_ (.A(uo_out[5]),
    .X(uo_out[1]));
 sg13g2_buf_1 _2056_ (.A(uo_out[6]),
    .X(uo_out[2]));
 sg13g2_buf_1 _2057_ (.A(\game_inst.o_vga_vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _2058_ (.A(\game_inst.o_vga_hsync ),
    .X(uo_out[7]));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[0].sreg_bufhigh  (.A(net222),
    .X(\game_inst.snake_inst.shiftreg_inst.high[0] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[100].sreg_bufhigh_173  (.L_HI(net223));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[100].sreg_bufhigh  (.A(net223),
    .X(\game_inst.snake_inst.shiftreg_inst.high[100] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[101].sreg_bufhigh_174  (.L_HI(net224));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[101].sreg_bufhigh  (.A(net224),
    .X(\game_inst.snake_inst.shiftreg_inst.high[101] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[102].sreg_bufhigh_175  (.L_HI(net225));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[102].sreg_bufhigh  (.A(net225),
    .X(\game_inst.snake_inst.shiftreg_inst.high[102] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[103].sreg_bufhigh_176  (.L_HI(net226));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[103].sreg_bufhigh  (.A(net226),
    .X(\game_inst.snake_inst.shiftreg_inst.high[103] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[104].sreg_bufhigh_177  (.L_HI(net227));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[104].sreg_bufhigh  (.A(net227),
    .X(\game_inst.snake_inst.shiftreg_inst.high[104] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[105].sreg_bufhigh_178  (.L_HI(net228));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[105].sreg_bufhigh  (.A(net228),
    .X(\game_inst.snake_inst.shiftreg_inst.high[105] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[106].sreg_bufhigh_179  (.L_HI(net229));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[106].sreg_bufhigh  (.A(net229),
    .X(\game_inst.snake_inst.shiftreg_inst.high[106] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[107].sreg_bufhigh_180  (.L_HI(net230));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[107].sreg_bufhigh  (.A(net230),
    .X(\game_inst.snake_inst.shiftreg_inst.high[107] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[108].sreg_bufhigh_181  (.L_HI(net231));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[108].sreg_bufhigh  (.A(net231),
    .X(\game_inst.snake_inst.shiftreg_inst.high[108] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[109].sreg_bufhigh_182  (.L_HI(net232));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[109].sreg_bufhigh  (.A(net232),
    .X(\game_inst.snake_inst.shiftreg_inst.high[109] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[10].sreg_bufhigh_183  (.L_HI(net233));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[10].sreg_bufhigh  (.A(net233),
    .X(\game_inst.snake_inst.shiftreg_inst.high[10] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[110].sreg_bufhigh_184  (.L_HI(net234));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[110].sreg_bufhigh  (.A(net234),
    .X(\game_inst.snake_inst.shiftreg_inst.high[110] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[111].sreg_bufhigh_185  (.L_HI(net235));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[111].sreg_bufhigh  (.A(net235),
    .X(\game_inst.snake_inst.shiftreg_inst.high[111] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[112].sreg_bufhigh_186  (.L_HI(net236));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[112].sreg_bufhigh  (.A(net236),
    .X(\game_inst.snake_inst.shiftreg_inst.high[112] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[113].sreg_bufhigh_187  (.L_HI(net237));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[113].sreg_bufhigh  (.A(net237),
    .X(\game_inst.snake_inst.shiftreg_inst.high[113] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[114].sreg_bufhigh_188  (.L_HI(net238));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[114].sreg_bufhigh  (.A(net238),
    .X(\game_inst.snake_inst.shiftreg_inst.high[114] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[115].sreg_bufhigh_189  (.L_HI(net239));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[115].sreg_bufhigh  (.A(net239),
    .X(\game_inst.snake_inst.shiftreg_inst.high[115] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[116].sreg_bufhigh_190  (.L_HI(net240));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[116].sreg_bufhigh  (.A(net240),
    .X(\game_inst.snake_inst.shiftreg_inst.high[116] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[11].sreg_bufhigh_191  (.L_HI(net241));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[11].sreg_bufhigh  (.A(net241),
    .X(\game_inst.snake_inst.shiftreg_inst.high[11] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[12].sreg_bufhigh_192  (.L_HI(net242));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[12].sreg_bufhigh  (.A(net242),
    .X(\game_inst.snake_inst.shiftreg_inst.high[12] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[13].sreg_bufhigh_193  (.L_HI(net243));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[13].sreg_bufhigh  (.A(net243),
    .X(\game_inst.snake_inst.shiftreg_inst.high[13] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[14].sreg_bufhigh_194  (.L_HI(net244));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[14].sreg_bufhigh  (.A(net244),
    .X(\game_inst.snake_inst.shiftreg_inst.high[14] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[15].sreg_bufhigh_195  (.L_HI(net245));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[15].sreg_bufhigh  (.A(net245),
    .X(\game_inst.snake_inst.shiftreg_inst.high[15] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[16].sreg_bufhigh_196  (.L_HI(net246));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[16].sreg_bufhigh  (.A(net246),
    .X(\game_inst.snake_inst.shiftreg_inst.high[16] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[17].sreg_bufhigh_197  (.L_HI(net247));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[17].sreg_bufhigh  (.A(net247),
    .X(\game_inst.snake_inst.shiftreg_inst.high[17] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[18].sreg_bufhigh_198  (.L_HI(net248));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[18].sreg_bufhigh  (.A(net248),
    .X(\game_inst.snake_inst.shiftreg_inst.high[18] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[19].sreg_bufhigh_199  (.L_HI(net249));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[19].sreg_bufhigh  (.A(net249),
    .X(\game_inst.snake_inst.shiftreg_inst.high[19] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[1].sreg_bufhigh_200  (.L_HI(net250));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[1].sreg_bufhigh  (.A(net250),
    .X(\game_inst.snake_inst.shiftreg_inst.high[1] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[20].sreg_bufhigh_201  (.L_HI(net251));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[20].sreg_bufhigh  (.A(net251),
    .X(\game_inst.snake_inst.shiftreg_inst.high[20] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[21].sreg_bufhigh_202  (.L_HI(net252));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[21].sreg_bufhigh  (.A(net252),
    .X(\game_inst.snake_inst.shiftreg_inst.high[21] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[22].sreg_bufhigh_203  (.L_HI(net253));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[22].sreg_bufhigh  (.A(net253),
    .X(\game_inst.snake_inst.shiftreg_inst.high[22] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[23].sreg_bufhigh_204  (.L_HI(net254));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[23].sreg_bufhigh  (.A(net254),
    .X(\game_inst.snake_inst.shiftreg_inst.high[23] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[24].sreg_bufhigh_205  (.L_HI(net255));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[24].sreg_bufhigh  (.A(net255),
    .X(\game_inst.snake_inst.shiftreg_inst.high[24] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[25].sreg_bufhigh_206  (.L_HI(net256));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[25].sreg_bufhigh  (.A(net256),
    .X(\game_inst.snake_inst.shiftreg_inst.high[25] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[26].sreg_bufhigh_207  (.L_HI(net257));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[26].sreg_bufhigh  (.A(net257),
    .X(\game_inst.snake_inst.shiftreg_inst.high[26] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[27].sreg_bufhigh_208  (.L_HI(net258));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[27].sreg_bufhigh  (.A(net258),
    .X(\game_inst.snake_inst.shiftreg_inst.high[27] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[28].sreg_bufhigh_209  (.L_HI(net259));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[28].sreg_bufhigh  (.A(net259),
    .X(\game_inst.snake_inst.shiftreg_inst.high[28] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[29].sreg_bufhigh_210  (.L_HI(net260));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[29].sreg_bufhigh  (.A(net260),
    .X(\game_inst.snake_inst.shiftreg_inst.high[29] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[2].sreg_bufhigh_211  (.L_HI(net261));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[2].sreg_bufhigh  (.A(net261),
    .X(\game_inst.snake_inst.shiftreg_inst.high[2] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[30].sreg_bufhigh_212  (.L_HI(net262));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[30].sreg_bufhigh  (.A(net262),
    .X(\game_inst.snake_inst.shiftreg_inst.high[30] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[31].sreg_bufhigh_213  (.L_HI(net263));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[31].sreg_bufhigh  (.A(net263),
    .X(\game_inst.snake_inst.shiftreg_inst.high[31] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[32].sreg_bufhigh_214  (.L_HI(net264));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[32].sreg_bufhigh  (.A(net264),
    .X(\game_inst.snake_inst.shiftreg_inst.high[32] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[33].sreg_bufhigh_215  (.L_HI(net265));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[33].sreg_bufhigh  (.A(net265),
    .X(\game_inst.snake_inst.shiftreg_inst.high[33] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[34].sreg_bufhigh_216  (.L_HI(net266));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[34].sreg_bufhigh  (.A(net266),
    .X(\game_inst.snake_inst.shiftreg_inst.high[34] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[35].sreg_bufhigh_217  (.L_HI(net267));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[35].sreg_bufhigh  (.A(net267),
    .X(\game_inst.snake_inst.shiftreg_inst.high[35] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[36].sreg_bufhigh_218  (.L_HI(net268));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[36].sreg_bufhigh  (.A(net268),
    .X(\game_inst.snake_inst.shiftreg_inst.high[36] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[37].sreg_bufhigh_219  (.L_HI(net269));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[37].sreg_bufhigh  (.A(net269),
    .X(\game_inst.snake_inst.shiftreg_inst.high[37] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[38].sreg_bufhigh_220  (.L_HI(net270));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[38].sreg_bufhigh  (.A(net270),
    .X(\game_inst.snake_inst.shiftreg_inst.high[38] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[39].sreg_bufhigh_221  (.L_HI(net271));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[39].sreg_bufhigh  (.A(net271),
    .X(\game_inst.snake_inst.shiftreg_inst.high[39] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[3].sreg_bufhigh_222  (.L_HI(net272));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[3].sreg_bufhigh  (.A(net272),
    .X(\game_inst.snake_inst.shiftreg_inst.high[3] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[40].sreg_bufhigh_223  (.L_HI(net273));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[40].sreg_bufhigh  (.A(net273),
    .X(\game_inst.snake_inst.shiftreg_inst.high[40] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[41].sreg_bufhigh_224  (.L_HI(net274));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[41].sreg_bufhigh  (.A(net274),
    .X(\game_inst.snake_inst.shiftreg_inst.high[41] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[42].sreg_bufhigh_225  (.L_HI(net275));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[42].sreg_bufhigh  (.A(net275),
    .X(\game_inst.snake_inst.shiftreg_inst.high[42] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[43].sreg_bufhigh_226  (.L_HI(net276));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[43].sreg_bufhigh  (.A(net276),
    .X(\game_inst.snake_inst.shiftreg_inst.high[43] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[44].sreg_bufhigh_227  (.L_HI(net277));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[44].sreg_bufhigh  (.A(net277),
    .X(\game_inst.snake_inst.shiftreg_inst.high[44] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[45].sreg_bufhigh_228  (.L_HI(net278));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[45].sreg_bufhigh  (.A(net278),
    .X(\game_inst.snake_inst.shiftreg_inst.high[45] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[46].sreg_bufhigh_229  (.L_HI(net279));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[46].sreg_bufhigh  (.A(net279),
    .X(\game_inst.snake_inst.shiftreg_inst.high[46] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[47].sreg_bufhigh_230  (.L_HI(net280));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[47].sreg_bufhigh  (.A(net280),
    .X(\game_inst.snake_inst.shiftreg_inst.high[47] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[48].sreg_bufhigh_231  (.L_HI(net281));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[48].sreg_bufhigh  (.A(net281),
    .X(\game_inst.snake_inst.shiftreg_inst.high[48] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[49].sreg_bufhigh_232  (.L_HI(net282));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[49].sreg_bufhigh  (.A(net282),
    .X(\game_inst.snake_inst.shiftreg_inst.high[49] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[4].sreg_bufhigh_233  (.L_HI(net283));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[4].sreg_bufhigh  (.A(net283),
    .X(\game_inst.snake_inst.shiftreg_inst.high[4] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[50].sreg_bufhigh_234  (.L_HI(net284));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[50].sreg_bufhigh  (.A(net284),
    .X(\game_inst.snake_inst.shiftreg_inst.high[50] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[51].sreg_bufhigh_235  (.L_HI(net285));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[51].sreg_bufhigh  (.A(net285),
    .X(\game_inst.snake_inst.shiftreg_inst.high[51] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[52].sreg_bufhigh_236  (.L_HI(net286));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[52].sreg_bufhigh  (.A(net286),
    .X(\game_inst.snake_inst.shiftreg_inst.high[52] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[53].sreg_bufhigh_237  (.L_HI(net287));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[53].sreg_bufhigh  (.A(net287),
    .X(\game_inst.snake_inst.shiftreg_inst.high[53] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[54].sreg_bufhigh_238  (.L_HI(net288));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[54].sreg_bufhigh  (.A(net288),
    .X(\game_inst.snake_inst.shiftreg_inst.high[54] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[55].sreg_bufhigh_239  (.L_HI(net289));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[55].sreg_bufhigh  (.A(net289),
    .X(\game_inst.snake_inst.shiftreg_inst.high[55] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[56].sreg_bufhigh_240  (.L_HI(net290));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[56].sreg_bufhigh  (.A(net290),
    .X(\game_inst.snake_inst.shiftreg_inst.high[56] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[57].sreg_bufhigh_241  (.L_HI(net291));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[57].sreg_bufhigh  (.A(net291),
    .X(\game_inst.snake_inst.shiftreg_inst.high[57] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[58].sreg_bufhigh_242  (.L_HI(net292));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[58].sreg_bufhigh  (.A(net292),
    .X(\game_inst.snake_inst.shiftreg_inst.high[58] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[59].sreg_bufhigh_243  (.L_HI(net293));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[59].sreg_bufhigh  (.A(net293),
    .X(\game_inst.snake_inst.shiftreg_inst.high[59] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[5].sreg_bufhigh_244  (.L_HI(net294));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[5].sreg_bufhigh  (.A(net294),
    .X(\game_inst.snake_inst.shiftreg_inst.high[5] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[60].sreg_bufhigh_245  (.L_HI(net295));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[60].sreg_bufhigh  (.A(net295),
    .X(\game_inst.snake_inst.shiftreg_inst.high[60] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[61].sreg_bufhigh_246  (.L_HI(net296));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[61].sreg_bufhigh  (.A(net296),
    .X(\game_inst.snake_inst.shiftreg_inst.high[61] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[62].sreg_bufhigh_247  (.L_HI(net297));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[62].sreg_bufhigh  (.A(net297),
    .X(\game_inst.snake_inst.shiftreg_inst.high[62] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[63].sreg_bufhigh_248  (.L_HI(net298));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[63].sreg_bufhigh  (.A(net298),
    .X(\game_inst.snake_inst.shiftreg_inst.high[63] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[64].sreg_bufhigh_249  (.L_HI(net299));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[64].sreg_bufhigh  (.A(net299),
    .X(\game_inst.snake_inst.shiftreg_inst.high[64] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[65].sreg_bufhigh_250  (.L_HI(net300));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[65].sreg_bufhigh  (.A(net300),
    .X(\game_inst.snake_inst.shiftreg_inst.high[65] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[66].sreg_bufhigh_251  (.L_HI(net301));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[66].sreg_bufhigh  (.A(net301),
    .X(\game_inst.snake_inst.shiftreg_inst.high[66] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[67].sreg_bufhigh_252  (.L_HI(net302));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[67].sreg_bufhigh  (.A(net302),
    .X(\game_inst.snake_inst.shiftreg_inst.high[67] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[68].sreg_bufhigh_253  (.L_HI(net303));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[68].sreg_bufhigh  (.A(net303),
    .X(\game_inst.snake_inst.shiftreg_inst.high[68] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[69].sreg_bufhigh_254  (.L_HI(net304));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[69].sreg_bufhigh  (.A(net304),
    .X(\game_inst.snake_inst.shiftreg_inst.high[69] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[6].sreg_bufhigh_255  (.L_HI(net305));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[6].sreg_bufhigh  (.A(net305),
    .X(\game_inst.snake_inst.shiftreg_inst.high[6] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[70].sreg_bufhigh_256  (.L_HI(net306));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[70].sreg_bufhigh  (.A(net306),
    .X(\game_inst.snake_inst.shiftreg_inst.high[70] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[71].sreg_bufhigh_257  (.L_HI(net307));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[71].sreg_bufhigh  (.A(net307),
    .X(\game_inst.snake_inst.shiftreg_inst.high[71] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[72].sreg_bufhigh_258  (.L_HI(net308));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[72].sreg_bufhigh  (.A(net308),
    .X(\game_inst.snake_inst.shiftreg_inst.high[72] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[73].sreg_bufhigh_259  (.L_HI(net309));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[73].sreg_bufhigh  (.A(net309),
    .X(\game_inst.snake_inst.shiftreg_inst.high[73] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[74].sreg_bufhigh_260  (.L_HI(net310));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[74].sreg_bufhigh  (.A(net310),
    .X(\game_inst.snake_inst.shiftreg_inst.high[74] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[75].sreg_bufhigh_261  (.L_HI(net311));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[75].sreg_bufhigh  (.A(net311),
    .X(\game_inst.snake_inst.shiftreg_inst.high[75] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[76].sreg_bufhigh_262  (.L_HI(net312));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[76].sreg_bufhigh  (.A(net312),
    .X(\game_inst.snake_inst.shiftreg_inst.high[76] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[77].sreg_bufhigh_263  (.L_HI(net313));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[77].sreg_bufhigh  (.A(net313),
    .X(\game_inst.snake_inst.shiftreg_inst.high[77] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[78].sreg_bufhigh_264  (.L_HI(net314));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[78].sreg_bufhigh  (.A(net314),
    .X(\game_inst.snake_inst.shiftreg_inst.high[78] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[79].sreg_bufhigh_265  (.L_HI(net315));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[79].sreg_bufhigh  (.A(net315),
    .X(\game_inst.snake_inst.shiftreg_inst.high[79] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[7].sreg_bufhigh_266  (.L_HI(net316));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[7].sreg_bufhigh  (.A(net316),
    .X(\game_inst.snake_inst.shiftreg_inst.high[7] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[80].sreg_bufhigh_267  (.L_HI(net317));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[80].sreg_bufhigh  (.A(net317),
    .X(\game_inst.snake_inst.shiftreg_inst.high[80] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[81].sreg_bufhigh_268  (.L_HI(net318));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[81].sreg_bufhigh  (.A(net318),
    .X(\game_inst.snake_inst.shiftreg_inst.high[81] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[82].sreg_bufhigh_269  (.L_HI(net319));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[82].sreg_bufhigh  (.A(net319),
    .X(\game_inst.snake_inst.shiftreg_inst.high[82] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[83].sreg_bufhigh_270  (.L_HI(net320));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[83].sreg_bufhigh  (.A(net320),
    .X(\game_inst.snake_inst.shiftreg_inst.high[83] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[84].sreg_bufhigh_271  (.L_HI(net321));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[84].sreg_bufhigh  (.A(net321),
    .X(\game_inst.snake_inst.shiftreg_inst.high[84] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[85].sreg_bufhigh_272  (.L_HI(net322));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[85].sreg_bufhigh  (.A(net322),
    .X(\game_inst.snake_inst.shiftreg_inst.high[85] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[86].sreg_bufhigh_273  (.L_HI(net323));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[86].sreg_bufhigh  (.A(net323),
    .X(\game_inst.snake_inst.shiftreg_inst.high[86] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[87].sreg_bufhigh_274  (.L_HI(net324));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[87].sreg_bufhigh  (.A(net324),
    .X(\game_inst.snake_inst.shiftreg_inst.high[87] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[88].sreg_bufhigh_275  (.L_HI(net325));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[88].sreg_bufhigh  (.A(net325),
    .X(\game_inst.snake_inst.shiftreg_inst.high[88] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[89].sreg_bufhigh_276  (.L_HI(net326));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[89].sreg_bufhigh  (.A(net326),
    .X(\game_inst.snake_inst.shiftreg_inst.high[89] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[8].sreg_bufhigh_277  (.L_HI(net327));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[8].sreg_bufhigh  (.A(net327),
    .X(\game_inst.snake_inst.shiftreg_inst.high[8] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[90].sreg_bufhigh_278  (.L_HI(net328));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[90].sreg_bufhigh  (.A(net328),
    .X(\game_inst.snake_inst.shiftreg_inst.high[90] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[91].sreg_bufhigh_279  (.L_HI(net329));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[91].sreg_bufhigh  (.A(net329),
    .X(\game_inst.snake_inst.shiftreg_inst.high[91] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[92].sreg_bufhigh_280  (.L_HI(net330));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[92].sreg_bufhigh  (.A(net330),
    .X(\game_inst.snake_inst.shiftreg_inst.high[92] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[93].sreg_bufhigh_281  (.L_HI(net331));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[93].sreg_bufhigh  (.A(net331),
    .X(\game_inst.snake_inst.shiftreg_inst.high[93] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[94].sreg_bufhigh_282  (.L_HI(net332));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[94].sreg_bufhigh  (.A(net332),
    .X(\game_inst.snake_inst.shiftreg_inst.high[94] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[95].sreg_bufhigh_283  (.L_HI(net333));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[95].sreg_bufhigh  (.A(net333),
    .X(\game_inst.snake_inst.shiftreg_inst.high[95] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[96].sreg_bufhigh_284  (.L_HI(net334));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[96].sreg_bufhigh  (.A(net334),
    .X(\game_inst.snake_inst.shiftreg_inst.high[96] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[97].sreg_bufhigh_285  (.L_HI(net335));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[97].sreg_bufhigh  (.A(net335),
    .X(\game_inst.snake_inst.shiftreg_inst.high[97] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[98].sreg_bufhigh_286  (.L_HI(net336));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[98].sreg_bufhigh  (.A(net336),
    .X(\game_inst.snake_inst.shiftreg_inst.high[98] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[99].sreg_bufhigh_287  (.L_HI(net337));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[99].sreg_bufhigh  (.A(net337),
    .X(\game_inst.snake_inst.shiftreg_inst.high[99] [0]));
 sg13g2_tiehi \game_inst.snake_inst.shiftreg_inst.genblk1[9].sreg_bufhigh_288  (.L_HI(net338));
 sg13g2_buf_1 \game_inst.snake_inst.shiftreg_inst.genblk1[9].sreg_bufhigh  (.A(net338),
    .X(\game_inst.snake_inst.shiftreg_inst.high[9] [0]));
 sg13g2_dfrbpq_2 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[0].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[0] [0]),
    .D(net483),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[0] [0]),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[100].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[50] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[100] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[100] [0]),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[101].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[50] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[101] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[101] [0]),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[102].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[51] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[102] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[102] [0]),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[103].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[51] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[103] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[103] [0]),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[104].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[52] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[104] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[104] [0]),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[105].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[52] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[105] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[105] [0]),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[106].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[53] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[106] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[106] [0]),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[107].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[53] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[107] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[107] [0]),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[108].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[54] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[108] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[108] [0]),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[109].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[54] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[109] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[109] [0]),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[10].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[5] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[10] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[10] [0]),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[110].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[55] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[110] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[110] [0]),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[111].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[55] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[111] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[111] [0]),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[112].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[56] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[112] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[112] [0]),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[113].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[56] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[113] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[113] [0]),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[114].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[57] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[114] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[114] [0]),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[115].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[57] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[115] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[115] [0]),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[116].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[58] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[116] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[116] [0]),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[117].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[58] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[117] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[117] [0]),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[118].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[59] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[118] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[118] [0]),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[119].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[59] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[119] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[119] [0]),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[11].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[5] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[11] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[11] [0]),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[120].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[60] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[120] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[120] [0]),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[121].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[60] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[121] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[121] [0]),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[122].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[61] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[122] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[122] [0]),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[123].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[61] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[123] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[123] [0]),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[124].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[62] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[124] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[124] [0]),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[125].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[62] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[125] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[125] [0]),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[126].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[63] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[126] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[126] [0]),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[127].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[63] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[127] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[127] [0]),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[128].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[64] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[128] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[128] [0]),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[129].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[64] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[129] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[129] [0]),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[12].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[6] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[12] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[12] [0]),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[130].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[65] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[130] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[130] [0]),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[131].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[65] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[131] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[131] [0]),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[132].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[66] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[132] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[132] [0]),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[133].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[66] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[133] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[133] [0]),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[134].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[67] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[134] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[134] [0]),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[135].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[67] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[135] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[135] [0]),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[136].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[68] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[136] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[136] [0]),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[137].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[68] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[137] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[137] [0]),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[138].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[69] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[138] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[138] [0]),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[139].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[69] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[139] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[139] [0]),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[13].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[6] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[13] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[13] [0]),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[140].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[70] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[140] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[140] [0]),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[141].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[70] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[141] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[141] [0]),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[142].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[71] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[142] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[142] [0]),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[143].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[71] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[143] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[143] [0]),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[144].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[72] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[144] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[144] [0]),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[145].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[72] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[145] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[145] [0]),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[146].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[73] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[146] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[146] [0]),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[147].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[73] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[147] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[147] [0]),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[148].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[74] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[148] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[148] [0]),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[149].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[74] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[149] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[149] [0]),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[14].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[7] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[14] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[14] [0]),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[150].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[75] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[150] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[150] [0]),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[151].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[75] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[151] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[151] [0]),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[152].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[76] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[152] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[152] [0]),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[153].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[76] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[153] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[153] [0]),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[154].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[77] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[154] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[154] [0]),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[155].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[77] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[155] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[155] [0]),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[156].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[78] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[156] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[156] [0]),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[157].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[78] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[157] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[157] [0]),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[158].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[79] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[158] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[158] [0]),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[159].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[79] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[159] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[159] [0]),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[15].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[7] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[15] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[15] [0]),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[160].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[80] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[160] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[160] [0]),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[161].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[80] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[161] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[161] [0]),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[162].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[81] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[162] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[162] [0]),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[163].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[81] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[163] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[163] [0]),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[164].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[82] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[164] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[164] [0]),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[165].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[82] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[165] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[165] [0]),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[166].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[83] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[166] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[166] [0]),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[167].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[83] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[167] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[167] [0]),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[168].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[84] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[168] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[168] [0]),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[169].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[84] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[169] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[169] [0]),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[16].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[8] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[16] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[16] [0]),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[170].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[85] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[170] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[170] [0]),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[171].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[85] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[171] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[171] [0]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[172].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[86] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[172] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[172] [0]),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[173].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[86] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[173] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[173] [0]),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[174].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[87] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[174] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[174] [0]),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[175].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[87] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[175] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[175] [0]),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[176].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[88] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[176] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[176] [0]),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[177].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[88] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[177] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[177] [0]),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[178].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[89] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[178] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[178] [0]),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[179].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[89] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[179] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[179] [0]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[17].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[8] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[17] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[17] [0]),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[180].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[90] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[180] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[180] [0]),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[181].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[90] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[181] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[181] [0]),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[182].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[91] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[182] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[182] [0]),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[183].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[91] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[183] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[183] [0]),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[184].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[92] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[184] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[184] [0]),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[185].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[92] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[185] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[185] [0]),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[186].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[93] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[186] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[186] [0]),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[187].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[93] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[187] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[187] [0]),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[188].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[94] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[188] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[188] [0]),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[189].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[94] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[189] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[189] [0]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[18].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[9] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[18] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[18] [0]),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[190].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[95] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[190] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[190] [0]),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[191].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[95] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[191] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[191] [0]),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[192].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[96] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[192] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[192] [0]),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[193].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[96] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[193] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[193] [0]),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[194].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[97] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[194] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[194] [0]),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[195].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[97] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[195] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[195] [0]),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[196].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[98] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[196] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[196] [0]),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[197].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[98] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[197] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[197] [0]),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[198].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[99] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[198] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[198] [0]),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[199].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[99] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[199] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[199] [0]),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[19].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[9] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[19] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[19] [0]),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[1].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[0] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[1] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[1] [0]),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[200].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[100] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[200] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[200] [0]),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[201].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[100] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[201] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[201] [0]),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[202].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[101] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[202] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[202] [0]),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[203].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[101] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[203] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[203] [0]),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[204].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[102] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[204] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[204] [0]),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[205].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[102] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[205] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[205] [0]),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[206].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[103] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[206] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[206] [0]),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[207].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[103] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[207] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[207] [0]),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[208].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[104] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[208] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[208] [0]),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[209].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[104] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[209] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[209] [0]),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[20].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[10] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[20] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[20] [0]),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[210].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[105] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[210] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[210] [0]),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[211].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[105] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[211] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[211] [0]),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[212].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[106] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[212] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[212] [0]),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[213].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[106] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[213] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[213] [0]),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[214].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[107] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[214] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[214] [0]),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[215].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[107] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[215] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[215] [0]),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[216].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[108] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[216] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[216] [0]),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[217].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[108] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[217] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[217] [0]),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[218].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[109] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[218] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[218] [0]),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[219].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[109] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[219] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[219] [0]),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[21].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[10] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[21] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[21] [0]),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[220].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[110] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[220] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[220] [0]),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[221].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[110] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[221] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[221] [0]),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[222].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[111] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[222] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[222] [0]),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[223].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[111] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[223] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[223] [0]),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[224].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[112] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[224] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[224] [0]),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[225].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[112] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[225] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[225] [0]),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[226].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[113] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[226] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[226] [0]),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[227].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[113] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[227] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[227] [0]),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[228].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[114] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[228] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[228] [0]),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[229].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[114] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[229] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[229] [0]),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[22].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[11] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[22] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[22] [0]),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[230].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[115] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[230] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[230] [0]),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[231].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[115] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[231] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[231] [0]),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[232].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[116] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[232] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[232] [0]),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[233].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[116] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[233] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[233] [0]),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[23].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[11] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[23] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[23] [0]),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[24].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[12] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[24] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[24] [0]),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[25].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[12] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[25] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[25] [0]),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[26].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[13] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[26] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[26] [0]),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[27].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[13] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[27] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[27] [0]),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[28].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[14] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[28] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[28] [0]),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[29].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[14] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[29] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[29] [0]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[2].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[1] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[2] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[2] [0]),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[30].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[15] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[30] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[30] [0]),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[31].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[15] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[31] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[31] [0]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[32].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[16] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[32] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[32] [0]),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[33].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[16] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[33] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[33] [0]),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[34].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[17] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[34] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[34] [0]),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[35].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[17] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[35] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[35] [0]),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[36].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[18] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[36] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[36] [0]),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[37].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[18] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[37] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[37] [0]),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[38].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[19] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[38] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[38] [0]),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[39].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[19] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[39] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[39] [0]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[3].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[1] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[3] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[3] [0]),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[40].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[20] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[40] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[40] [0]),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[41].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[20] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[41] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[41] [0]),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[42].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[21] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[42] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[42] [0]),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[43].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[21] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[43] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[43] [0]),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[44].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[22] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[44] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[44] [0]),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[45].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[22] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[45] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[45] [0]),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[46].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[23] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[46] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[46] [0]),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[47].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[23] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[47] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[47] [0]),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[48].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[24] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[48] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[48] [0]),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[49].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[24] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[49] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[49] [0]),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[4].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[2] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[4] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[4] [0]),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[50].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[25] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[50] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[50] [0]),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[51].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[25] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[51] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[51] [0]),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[52].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[26] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[52] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[52] [0]),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[53].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[26] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[53] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[53] [0]),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[54].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[27] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[54] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[54] [0]),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[55].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[27] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[55] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[55] [0]),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[56].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[28] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[56] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[56] [0]),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[57].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[28] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[57] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[57] [0]),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[58].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[29] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[58] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[58] [0]),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[59].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[29] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[59] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[59] [0]),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[5].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[2] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[5] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[5] [0]),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[60].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[30] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[60] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[60] [0]),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[61].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[30] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[61] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[61] [0]),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[62].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[31] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[62] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[62] [0]),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[63].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[31] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[63] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[63] [0]),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[64].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[32] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[64] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[64] [0]),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[65].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[32] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[65] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[65] [0]),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[66].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[33] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[66] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[66] [0]),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[67].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[33] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[67] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[67] [0]),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[68].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[34] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[68] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[68] [0]),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[69].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[34] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[69] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[69] [0]),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[6].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[3] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[6] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[6] [0]),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[70].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[35] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[70] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[70] [0]),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[71].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[35] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[71] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[71] [0]),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[72].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[36] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[72] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[72] [0]),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[73].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[36] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[73] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[73] [0]),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[74].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[37] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[74] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[74] [0]),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[75].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[37] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[75] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[75] [0]),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[76].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[38] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[76] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[76] [0]),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[77].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[38] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[77] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[77] [0]),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[78].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[39] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[78] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[78] [0]),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[79].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[39] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[79] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[79] [0]),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[7].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[3] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[7] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[7] [0]),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[80].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[40] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[80] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[80] [0]),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[81].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[40] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[81] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[81] [0]),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[82].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[41] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[82] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[82] [0]),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[83].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[41] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[83] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[83] [0]),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[84].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[42] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[84] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[84] [0]),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[85].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[42] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[85] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[85] [0]),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[86].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[43] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[86] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[86] [0]),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[87].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[43] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[87] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[87] [0]),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[88].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[44] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[88] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[88] [0]),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[89].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[44] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[89] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[89] [0]),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[8].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[4] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[8] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[8] [0]),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[90].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[45] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[90] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[90] [0]),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[91].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[45] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[91] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[91] [0]),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[92].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[46] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[92] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[92] [0]),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[93].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[46] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[93] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[93] [0]),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[94].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[47] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[94] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[94] [0]),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[95].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[47] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[95] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[95] [0]),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[96].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[48] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[96] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[96] [0]),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[97].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[48] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[97] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[97] [0]),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[98].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[49] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[98] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[98] [0]),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[99].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[49] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[99] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[99] [0]),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[0].genblk1[9].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[4] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[9] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[9] [0]),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dlygate4sd3_1 dly2_0_1 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[1] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[2] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_101 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[101] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[102] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_102 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[102] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[103] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_103 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[103] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[104] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_104 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[104] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[105] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_105 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[105] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[106] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_106 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[106] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[107] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_107 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[107] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[108] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_108 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[108] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[109] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_109 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[109] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[110] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_110 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[110] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[111] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_11 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[11] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[12] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_111 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[111] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[112] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_112 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[112] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[113] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_113 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[113] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[114] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_114 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[114] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[115] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_115 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[115] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[116] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_116 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[116] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[117] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_117 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[117] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[118] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_118 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[118] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[119] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_119 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[119] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[120] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_120 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[120] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[121] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_12 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[12] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[13] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_121 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[121] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[122] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_122 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[122] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[123] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_123 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[123] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[124] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_124 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[124] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[125] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_125 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[125] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[126] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_126 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[126] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[127] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_127 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[127] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[128] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_128 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[128] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[129] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_129 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[129] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[130] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_130 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[130] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[131] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_13 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[13] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[14] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_131 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[131] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[132] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_132 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[132] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[133] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_133 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[133] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[134] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_134 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[134] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[135] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_135 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[135] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[136] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_136 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[136] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[137] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_137 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[137] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[138] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_138 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[138] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[139] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_139 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[139] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[140] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_140 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[140] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[141] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_14 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[14] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[15] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_141 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[141] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[142] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_142 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[142] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[143] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_143 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[143] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[144] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_144 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[144] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[145] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_145 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[145] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[146] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_146 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[146] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[147] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_147 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[147] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[148] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_148 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[148] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[149] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_149 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[149] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[150] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_150 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[150] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[151] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_15 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[15] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[16] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_151 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[151] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[152] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_152 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[152] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[153] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_153 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[153] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[154] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_154 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[154] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[155] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_155 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[155] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[156] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_156 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[156] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[157] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_157 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[157] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[158] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_158 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[158] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[159] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_159 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[159] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[160] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_160 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[160] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[161] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_16 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[16] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[17] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_161 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[161] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[162] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_162 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[162] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[163] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_163 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[163] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[164] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_164 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[164] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[165] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_165 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[165] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[166] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_166 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[166] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[167] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_167 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[167] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[168] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_168 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[168] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[169] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_169 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[169] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[170] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_170 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[170] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[171] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_17 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[17] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[18] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_171 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[171] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[172] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_172 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[172] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[173] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_173 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[173] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[174] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_174 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[174] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[175] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_175 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[175] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[176] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_176 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[176] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[177] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_177 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[177] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[178] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_178 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[178] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[179] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_179 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[179] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[180] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_180 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[180] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[181] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_18 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[18] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[19] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_181 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[181] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[182] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_182 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[182] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[183] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_183 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[183] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[184] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_184 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[184] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[185] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_185 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[185] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[186] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_186 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[186] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[187] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_187 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[187] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[188] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_188 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[188] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[189] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_189 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[189] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[190] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_190 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[190] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[191] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_19 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[19] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[20] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_191 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[191] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[192] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_192 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[192] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[193] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_193 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[193] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[194] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_194 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[194] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[195] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_195 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[195] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[196] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_196 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[196] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[197] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_197 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[197] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[198] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_198 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[198] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[199] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_199 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[199] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[200] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_200 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[200] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[201] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_20 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[20] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[21] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_2 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[2] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[3] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_201 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[201] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[202] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_202 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[202] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[203] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_203 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[203] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[204] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_204 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[204] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[205] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_205 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[205] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[206] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_206 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[206] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[207] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_207 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[207] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[208] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_208 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[208] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[209] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_209 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[209] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[210] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_210 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[210] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[211] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_21 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[21] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[22] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_211 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[211] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[212] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_212 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[212] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[213] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_213 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[213] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[214] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_214 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[214] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[215] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_215 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[215] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[216] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_216 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[216] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[217] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_217 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[217] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[218] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_218 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[218] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[219] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_219 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[219] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[220] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_220 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[220] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[221] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_22 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[22] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[23] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_221 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[221] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[222] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_222 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[222] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[223] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_223 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[223] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[224] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_224 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[224] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[225] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_225 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[225] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[226] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_226 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[226] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[227] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_227 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[227] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[228] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_228 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[228] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[229] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_229 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[229] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[230] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_230 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[230] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[231] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_23 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[23] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[24] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_231 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[231] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[232] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_232 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[232] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[233] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_0 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[0] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[1] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_24 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[24] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[25] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_25 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[25] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[26] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_26 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[26] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[27] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_27 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[27] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[28] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_28 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[28] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[29] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_29 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[29] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[30] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_30 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[30] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[31] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_3 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[3] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[4] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_31 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[31] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[32] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_32 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[32] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[33] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_33 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[33] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[34] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_34 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[34] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[35] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_35 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[35] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[36] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_36 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[36] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[37] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_37 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[37] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[38] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_38 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[38] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[39] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_39 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[39] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[40] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_40 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[40] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[41] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_4 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[4] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[5] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_41 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[41] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[42] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_42 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[42] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[43] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_43 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[43] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[44] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_44 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[44] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[45] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_45 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[45] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[46] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_46 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[46] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[47] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_47 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[47] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[48] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_48 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[48] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[49] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_49 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[49] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[50] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_50 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[50] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[51] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_5 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[5] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[6] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_51 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[51] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[52] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_52 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[52] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[53] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_53 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[53] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[54] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_54 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[54] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[55] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_55 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[55] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[56] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_56 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[56] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[57] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_57 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[57] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[58] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_58 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[58] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[59] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_59 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[59] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[60] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_60 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[60] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[61] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_6 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[6] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[7] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_61 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[61] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[62] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_62 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[62] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[63] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_63 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[63] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[64] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_64 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[64] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[65] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_65 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[65] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[66] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_66 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[66] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[67] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_67 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[67] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[68] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_68 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[68] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[69] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_69 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[69] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[70] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_70 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[70] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[71] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_7 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[7] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[8] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_71 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[71] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[72] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_72 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[72] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[73] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_73 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[73] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[74] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_74 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[74] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[75] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_75 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[75] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[76] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_76 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[76] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[77] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_77 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[77] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[78] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_78 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[78] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[79] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_79 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[79] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[80] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_80 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[80] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[81] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_8 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[8] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[9] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_81 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[81] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[82] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_82 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[82] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[83] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_83 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[83] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[84] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_84 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[84] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[85] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_85 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[85] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[86] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_86 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[86] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[87] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_87 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[87] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[88] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_88 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[88] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[89] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_89 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[89] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[90] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_90 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[90] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[91] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_9 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[9] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[10] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_91 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[91] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[92] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_92 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[92] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[93] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_93 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[93] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[94] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_94 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[94] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[95] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_95 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[95] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[96] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_96 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[96] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[97] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_97 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[97] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[98] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_98 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[98] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[99] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_99 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[99] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[100] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_100 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[100] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[101] [0]));
 sg13g2_dlygate4sd3_1 dly2_0_10 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[10] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[11] [0]));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[0].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[0] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[0] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[0] [0]),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[100].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[50] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[100] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[100] [0]),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[101].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[50] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[101] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[101] [0]),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[102].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[51] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[102] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[102] [0]),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[103].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[51] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[103] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[103] [0]),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[104].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[52] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[104] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[104] [0]),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[105].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[52] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[105] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[105] [0]),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[106].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[53] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[106] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[106] [0]),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[107].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[53] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[107] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[107] [0]),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[108].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[54] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[108] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[108] [0]),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[109].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[54] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[109] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[109] [0]),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[10].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[5] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[10] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[10] [0]),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[110].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[55] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[110] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[110] [0]),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[111].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[55] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[111] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[111] [0]),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[112].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[56] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[112] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[112] [0]),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[113].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[56] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[113] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[113] [0]),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[114].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[57] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[114] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[114] [0]),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[115].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[57] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[115] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[115] [0]),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[116].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[58] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[116] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[116] [0]),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[117].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[58] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[117] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[117] [0]),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[118].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[59] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[118] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[118] [0]),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[119].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[59] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[119] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[119] [0]),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[11].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[5] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[11] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[11] [0]),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[120].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[60] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[120] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[120] [0]),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[121].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[60] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[121] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[121] [0]),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[122].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[61] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[122] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[122] [0]),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[123].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[61] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[123] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[123] [0]),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[124].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[62] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[124] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[124] [0]),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[125].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[62] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[125] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[125] [0]),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[126].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[63] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[126] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[126] [0]),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[127].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[63] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[127] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[127] [0]),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[128].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[64] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[128] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[128] [0]),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[129].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[64] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[129] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[129] [0]),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[12].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[6] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[12] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[12] [0]),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[130].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[65] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[130] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[130] [0]),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[131].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[65] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[131] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[131] [0]),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[132].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[66] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[132] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[132] [0]),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[133].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[66] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[133] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[133] [0]),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[134].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[67] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[134] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[134] [0]),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[135].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[67] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[135] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[135] [0]),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[136].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[68] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[136] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[136] [0]),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[137].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[68] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[137] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[137] [0]),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[138].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[69] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[138] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[138] [0]),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[139].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[69] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[139] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[139] [0]),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[13].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[6] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[13] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[13] [0]),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[140].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[70] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[140] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[140] [0]),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[141].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[70] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[141] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[141] [0]),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[142].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[71] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[142] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[142] [0]),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[143].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[71] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[143] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[143] [0]),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[144].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[72] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[144] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[144] [0]),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[145].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[72] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[145] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[145] [0]),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[146].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[73] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[146] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[146] [0]),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[147].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[73] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[147] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[147] [0]),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[148].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[74] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[148] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[148] [0]),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[149].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[74] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[149] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[149] [0]),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[14].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[7] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[14] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[14] [0]),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[150].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[75] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[150] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[150] [0]),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[151].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[75] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[151] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[151] [0]),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[152].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[76] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[152] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[152] [0]),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[153].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[76] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[153] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[153] [0]),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[154].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[77] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[154] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[154] [0]),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[155].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[77] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[155] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[155] [0]),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[156].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[78] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[156] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[156] [0]),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[157].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[78] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[157] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[157] [0]),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[158].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[79] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[158] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[158] [0]),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[159].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[79] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[159] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[159] [0]),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[15].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[7] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[15] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[15] [0]),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[160].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[80] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[160] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[160] [0]),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[161].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[80] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[161] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[161] [0]),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[162].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[81] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[162] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[162] [0]),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[163].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[81] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[163] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[163] [0]),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[164].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[82] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[164] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[164] [0]),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[165].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[82] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[165] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[165] [0]),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[166].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[83] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[166] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[166] [0]),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[167].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[83] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[167] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[167] [0]),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[168].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[84] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[168] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[168] [0]),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[169].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[84] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[169] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[169] [0]),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[16].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[8] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[16] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[16] [0]),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[170].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[85] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[170] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[170] [0]),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[171].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[85] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[171] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[171] [0]),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[172].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[86] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[172] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[172] [0]),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[173].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[86] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[173] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[173] [0]),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[174].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[87] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[174] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[174] [0]),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[175].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[87] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[175] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[175] [0]),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[176].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[88] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[176] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[176] [0]),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[177].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[88] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[177] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[177] [0]),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[178].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[89] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[178] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[178] [0]),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[179].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[89] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[179] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[179] [0]),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[17].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[8] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[17] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[17] [0]),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[180].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[90] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[180] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[180] [0]),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[181].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[90] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[181] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[181] [0]),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[182].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[91] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[182] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[182] [0]),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[183].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[91] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[183] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[183] [0]),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[184].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[92] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[184] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[184] [0]),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[185].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[92] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[185] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[185] [0]),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[186].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[93] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[186] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[186] [0]),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[187].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[93] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[187] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[187] [0]),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[188].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[94] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[188] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[188] [0]),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[189].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[94] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[189] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[189] [0]),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[18].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[9] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[18] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[18] [0]),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[190].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[95] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[190] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[190] [0]),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[191].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[95] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[191] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[191] [0]),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[192].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[96] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[192] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[192] [0]),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[193].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[96] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[193] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[193] [0]),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[194].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[97] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[194] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[194] [0]),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[195].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[97] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[195] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[195] [0]),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[196].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[98] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[196] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[196] [0]),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[197].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[98] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[197] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[197] [0]),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[198].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[99] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[198] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[198] [0]),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[199].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[99] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[199] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[199] [0]),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[19].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[9] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[19] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[19] [0]),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[1].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[0] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[1] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[1] [0]),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[200].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[100] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[200] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[200] [0]),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[201].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[100] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[201] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[201] [0]),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[202].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[101] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[202] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[202] [0]),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[203].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[101] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[203] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[203] [0]),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[204].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[102] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[204] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[204] [0]),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[205].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[102] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[205] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[205] [0]),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[206].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[103] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[206] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[206] [0]),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[207].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[103] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[207] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[207] [0]),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[208].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[104] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[208] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[208] [0]),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[209].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[104] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[209] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[209] [0]),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[20].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[10] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[20] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[20] [0]),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[210].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[105] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[210] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[210] [0]),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[211].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[105] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[211] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[211] [0]),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[212].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[106] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[212] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[212] [0]),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[213].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[106] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[213] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[213] [0]),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[214].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[107] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[214] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[214] [0]),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[215].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[107] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[215] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[215] [0]),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[216].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[108] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[216] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[216] [0]),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[217].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[108] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[217] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[217] [0]),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[218].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[109] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[218] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[218] [0]),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[219].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[109] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[219] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[219] [0]),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[21].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[10] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[21] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[21] [0]),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[220].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[110] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[220] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[220] [0]),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[221].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[110] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[221] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[221] [0]),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[222].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[111] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[222] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[222] [0]),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[223].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[111] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[223] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[223] [0]),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[224].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[112] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[224] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[224] [0]),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[225].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[112] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[225] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[225] [0]),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[226].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[113] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[226] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[226] [0]),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[227].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[113] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[227] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[227] [0]),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[228].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[114] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[228] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[228] [0]),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[229].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[114] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[229] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[229] [0]),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[22].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[11] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[22] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[22] [0]),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[230].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[115] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[230] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[230] [0]),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[231].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[115] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[231] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[231] [0]),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[232].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[116] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[232] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[232] [0]),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[233].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[116] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[233] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[233] [0]),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[23].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[11] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[23] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[23] [0]),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[24].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[12] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[24] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[24] [0]),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[25].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[12] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[25] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[25] [0]),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[26].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[13] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[26] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[26] [0]),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[27].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[13] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[27] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[27] [0]),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[28].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[14] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[28] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[28] [0]),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[29].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[14] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[29] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[29] [0]),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[2].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[1] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[2] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[2] [0]),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[30].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[15] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[30] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[30] [0]),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[31].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[15] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[31] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[31] [0]),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[32].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[16] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[32] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[32] [0]),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[33].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[16] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[33] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[33] [0]),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[34].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[17] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[34] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[34] [0]),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[35].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[17] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[35] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[35] [0]),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[36].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[18] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[36] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[36] [0]),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[37].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[18] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[37] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[37] [0]),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[38].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[19] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[38] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[38] [0]),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[39].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[19] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[39] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[39] [0]),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[3].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[1] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[3] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[3] [0]),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[40].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[20] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[40] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[40] [0]),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[41].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[20] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[41] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[41] [0]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[42].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[21] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[42] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[42] [0]),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[43].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[21] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[43] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[43] [0]),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[44].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[22] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[44] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[44] [0]),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[45].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[22] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[45] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[45] [0]),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[46].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[23] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[46] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[46] [0]),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[47].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[23] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[47] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[47] [0]),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[48].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[24] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[48] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[48] [0]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[49].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[24] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[49] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[49] [0]),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[4].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[2] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[4] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[4] [0]),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[50].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[25] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[50] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[50] [0]),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[51].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[25] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[51] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[51] [0]),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[52].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[26] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[52] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[52] [0]),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[53].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[26] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[53] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[53] [0]),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[54].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[27] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[54] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[54] [0]),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[55].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[27] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[55] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[55] [0]),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[56].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[28] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[56] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[56] [0]),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[57].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[28] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[57] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[57] [0]),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[58].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[29] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[58] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[58] [0]),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[59].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[29] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[59] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[59] [0]),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[5].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[2] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[5] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[5] [0]),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[60].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[30] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[60] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[60] [0]),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[61].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[30] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[61] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[61] [0]),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[62].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[31] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[62] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[62] [0]),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[63].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[31] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[63] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[63] [0]),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[64].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[32] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[64] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[64] [0]),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[65].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[32] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[65] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[65] [0]),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[66].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[33] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[66] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[66] [0]),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[67].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[33] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[67] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[67] [0]),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[68].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[34] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[68] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[68] [0]),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[69].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[34] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[69] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[69] [0]),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[6].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[3] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[6] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[6] [0]),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[70].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[35] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[70] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[70] [0]),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[71].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[35] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[71] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[71] [0]),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[72].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[36] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[72] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[72] [0]),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[73].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[36] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[73] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[73] [0]),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[74].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[37] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[74] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[74] [0]),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[75].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[37] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[75] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[75] [0]),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[76].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[38] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[76] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[76] [0]),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[77].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[38] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[77] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[77] [0]),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[78].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[39] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[78] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[78] [0]),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[79].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[39] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[79] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[79] [0]),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[7].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[3] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[7] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[7] [0]),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[80].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[40] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[80] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[80] [0]),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[81].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[40] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[81] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[81] [0]),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[82].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[41] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[82] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[82] [0]),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[83].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[41] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[83] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[83] [0]),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[84].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[42] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[84] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[84] [0]),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[85].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[42] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[85] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[85] [0]),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[86].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[43] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[86] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[86] [0]),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[87].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[43] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[87] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[87] [0]),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[88].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[44] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[88] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[88] [0]),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[89].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[44] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[89] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[89] [0]),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[8].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[4] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[8] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[8] [0]),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[90].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[45] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[90] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[90] [0]),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[91].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[45] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[91] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[91] [0]),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[92].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[46] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[92] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[92] [0]),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[93].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[46] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[93] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[93] [0]),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[94].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[47] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[94] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[94] [0]),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[95].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[47] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[95] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[95] [0]),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[96].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[48] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[96] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[96] [0]),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[97].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[48] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[97] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[97] [0]),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[98].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[49] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[98] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[98] [0]),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[99].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[49] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[99] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[99] [0]),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 \game_inst.snake_inst.shiftreg_inst.genblk2[1].genblk1[9].genblk1.sreg_dff  (.RESET_B(\game_inst.snake_inst.shiftreg_inst.high[4] [0]),
    .D(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[9] [0]),
    .Q(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[9] [0]),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dlygate4sd3_1 dly2_1_1 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[1] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[2] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_101 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[101] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[102] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_102 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[102] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[103] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_103 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[103] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[104] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_104 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[104] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[105] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_105 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[105] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[106] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_106 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[106] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[107] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_107 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[107] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[108] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_108 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[108] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[109] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_109 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[109] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[110] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_110 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[110] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[111] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_11 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[11] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[12] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_111 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[111] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[112] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_112 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[112] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[113] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_113 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[113] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[114] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_114 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[114] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[115] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_115 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[115] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[116] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_116 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[116] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[117] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_117 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[117] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[118] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_118 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[118] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[119] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_119 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[119] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[120] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_120 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[120] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[121] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_12 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[12] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[13] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_121 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[121] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[122] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_122 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[122] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[123] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_123 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[123] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[124] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_124 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[124] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[125] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_125 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[125] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[126] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_126 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[126] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[127] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_127 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[127] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[128] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_128 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[128] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[129] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_129 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[129] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[130] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_130 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[130] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[131] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_13 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[13] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[14] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_131 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[131] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[132] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_132 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[132] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[133] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_133 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[133] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[134] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_134 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[134] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[135] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_135 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[135] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[136] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_136 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[136] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[137] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_137 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[137] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[138] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_138 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[138] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[139] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_139 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[139] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[140] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_140 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[140] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[141] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_14 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[14] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[15] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_141 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[141] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[142] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_142 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[142] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[143] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_143 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[143] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[144] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_144 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[144] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[145] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_145 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[145] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[146] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_146 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[146] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[147] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_147 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[147] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[148] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_148 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[148] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[149] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_149 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[149] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[150] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_150 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[150] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[151] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_15 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[15] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[16] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_151 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[151] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[152] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_152 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[152] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[153] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_153 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[153] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[154] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_154 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[154] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[155] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_155 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[155] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[156] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_156 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[156] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[157] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_157 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[157] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[158] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_158 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[158] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[159] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_159 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[159] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[160] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_160 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[160] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[161] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_16 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[16] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[17] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_161 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[161] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[162] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_162 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[162] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[163] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_163 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[163] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[164] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_164 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[164] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[165] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_165 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[165] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[166] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_166 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[166] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[167] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_167 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[167] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[168] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_168 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[168] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[169] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_169 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[169] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[170] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_170 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[170] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[171] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_17 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[17] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[18] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_171 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[171] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[172] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_172 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[172] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[173] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_173 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[173] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[174] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_174 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[174] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[175] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_175 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[175] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[176] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_176 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[176] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[177] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_177 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[177] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[178] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_178 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[178] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[179] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_179 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[179] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[180] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_180 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[180] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[181] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_18 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[18] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[19] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_181 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[181] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[182] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_182 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[182] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[183] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_183 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[183] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[184] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_184 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[184] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[185] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_185 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[185] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[186] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_186 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[186] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[187] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_187 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[187] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[188] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_188 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[188] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[189] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_189 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[189] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[190] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_190 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[190] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[191] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_19 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[19] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[20] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_191 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[191] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[192] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_192 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[192] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[193] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_193 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[193] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[194] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_194 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[194] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[195] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_195 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[195] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[196] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_196 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[196] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[197] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_197 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[197] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[198] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_198 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[198] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[199] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_199 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[199] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[200] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_200 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[200] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[201] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_20 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[20] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[21] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_2 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[2] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[3] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_201 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[201] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[202] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_202 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[202] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[203] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_203 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[203] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[204] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_204 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[204] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[205] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_205 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[205] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[206] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_206 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[206] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[207] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_207 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[207] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[208] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_208 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[208] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[209] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_209 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[209] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[210] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_210 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[210] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[211] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_21 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[21] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[22] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_211 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[211] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[212] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_212 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[212] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[213] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_213 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[213] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[214] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_214 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[214] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[215] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_215 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[215] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[216] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_216 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[216] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[217] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_217 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[217] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[218] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_218 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[218] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[219] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_219 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[219] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[220] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_220 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[220] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[221] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_22 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[22] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[23] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_221 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[221] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[222] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_222 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[222] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[223] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_223 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[223] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[224] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_224 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[224] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[225] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_225 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[225] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[226] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_226 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[226] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[227] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_227 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[227] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[228] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_228 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[228] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[229] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_229 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[229] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[230] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_230 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[230] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[231] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_23 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[23] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[24] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_231 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[231] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[232] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_232 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[232] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[233] [0]));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_dlygate4sd3_1 dly2_1_24 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[24] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[25] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_25 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[25] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[26] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_26 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[26] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[27] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_27 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[27] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[28] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_28 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[28] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[29] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_29 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[29] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[30] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_30 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[30] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[31] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_3 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[3] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[4] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_31 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[31] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[32] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_32 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[32] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[33] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_33 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[33] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[34] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_34 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[34] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[35] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_35 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[35] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[36] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_36 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[36] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[37] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_37 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[37] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[38] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_38 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[38] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[39] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_39 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[39] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[40] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_40 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[40] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[41] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_4 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[4] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[5] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_41 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[41] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[42] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_42 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[42] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[43] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_43 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[43] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[44] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_44 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[44] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[45] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_45 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[45] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[46] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_46 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[46] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[47] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_47 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[47] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[48] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_48 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[48] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[49] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_49 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[49] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[50] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_50 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[50] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[51] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_5 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[5] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[6] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_51 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[51] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[52] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_52 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[52] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[53] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_53 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[53] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[54] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_54 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[54] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[55] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_55 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[55] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[56] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_56 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[56] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[57] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_57 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[57] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[58] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_58 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[58] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[59] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_59 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[59] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[60] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_60 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[60] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[61] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_6 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[6] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[7] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_61 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[61] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[62] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_62 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[62] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[63] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_63 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[63] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[64] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_64 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[64] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[65] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_65 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[65] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[66] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_66 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[66] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[67] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_67 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[67] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[68] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_68 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[68] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[69] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_69 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[69] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[70] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_70 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[70] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[71] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_7 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[7] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[8] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_71 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[71] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[72] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_72 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[72] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[73] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_73 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[73] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[74] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_74 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[74] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[75] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_75 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[75] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[76] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_76 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[76] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[77] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_77 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[77] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[78] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_78 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[78] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[79] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_79 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[79] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[80] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_80 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[80] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[81] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_8 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[8] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[9] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_81 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[81] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[82] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_82 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[82] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[83] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_83 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[83] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[84] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_84 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[84] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[85] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_85 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[85] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[86] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_86 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[86] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[87] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_87 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[87] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[88] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_88 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[88] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[89] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_89 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[89] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[90] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_90 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[90] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[91] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_9 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[9] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[10] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_91 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[91] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[92] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_92 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[92] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[93] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_93 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[93] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[94] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_94 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[94] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[95] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_95 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[95] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[96] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_96 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[96] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[97] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_97 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[97] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[98] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_98 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[98] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[99] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_99 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[99] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[100] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_100 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[100] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[101] [0]));
 sg13g2_dlygate4sd3_1 dly2_1_10 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[10] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_w[11] [0]));
 sg13g2_fill_1 FILLER_80_312 ();
 sg13g2_fill_2 FILLER_80_310 ();
 sg13g2_fill_1 FILLER_80_282 ();
 sg13g2_fill_2 FILLER_80_280 ();
 sg13g2_fill_1 FILLER_80_274 ();
 sg13g2_fill_2 FILLER_80_220 ();
 sg13g2_fill_1 FILLER_80_215 ();
 sg13g2_fill_2 FILLER_80_213 ();
 sg13g2_fill_2 FILLER_80_180 ();
 sg13g2_fill_1 FILLER_80_166 ();
 sg13g2_fill_2 FILLER_80_164 ();
 sg13g2_fill_2 FILLER_80_116 ();
 sg13g2_fill_1 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_fill_2 FILLER_79_407 ();
 sg13g2_fill_1 FILLER_79_347 ();
 sg13g2_fill_2 FILLER_79_313 ();
 sg13g2_fill_2 FILLER_79_185 ();
 sg13g2_fill_1 FILLER_79_176 ();
 sg13g2_fill_2 FILLER_79_75 ();
 sg13g2_fill_2 FILLER_79_32 ();
 sg13g2_decap_4 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_fill_2 FILLER_78_389 ();
 sg13g2_fill_1 FILLER_78_272 ();
 sg13g2_fill_1 FILLER_78_249 ();
 sg13g2_fill_2 FILLER_78_214 ();
 sg13g2_fill_1 FILLER_78_155 ();
 sg13g2_fill_1 FILLER_78_37 ();
 sg13g2_fill_2 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_fill_1 FILLER_77_375 ();
 sg13g2_fill_2 FILLER_77_350 ();
 sg13g2_fill_2 FILLER_77_206 ();
 sg13g2_fill_1 FILLER_77_197 ();
 sg13g2_fill_1 FILLER_77_102 ();
 sg13g2_fill_1 FILLER_77_46 ();
 sg13g2_decap_4 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_76_351 ();
 sg13g2_fill_2 FILLER_76_238 ();
 sg13g2_fill_2 FILLER_76_209 ();
 sg13g2_fill_2 FILLER_76_203 ();
 sg13g2_fill_1 FILLER_76_163 ();
 sg13g2_fill_2 FILLER_76_161 ();
 sg13g2_fill_1 FILLER_76_139 ();
 sg13g2_fill_2 FILLER_76_137 ();
 sg13g2_fill_1 FILLER_76_114 ();
 sg13g2_fill_2 FILLER_76_112 ();
 sg13g2_decap_4 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_75_365 ();
 sg13g2_fill_1 FILLER_75_314 ();
 sg13g2_fill_2 FILLER_75_262 ();
 sg13g2_fill_2 FILLER_75_247 ();
 sg13g2_fill_1 FILLER_75_202 ();
 sg13g2_fill_1 FILLER_75_192 ();
 sg13g2_fill_1 FILLER_75_182 ();
 sg13g2_fill_2 FILLER_75_180 ();
 sg13g2_fill_1 FILLER_75_171 ();
 sg13g2_fill_2 FILLER_75_169 ();
 sg13g2_fill_2 FILLER_75_104 ();
 sg13g2_fill_1 FILLER_75_94 ();
 sg13g2_fill_1 FILLER_75_44 ();
 sg13g2_fill_2 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_fill_2 FILLER_74_355 ();
 sg13g2_fill_1 FILLER_74_345 ();
 sg13g2_fill_1 FILLER_74_329 ();
 sg13g2_fill_1 FILLER_74_245 ();
 sg13g2_fill_2 FILLER_74_238 ();
 sg13g2_fill_1 FILLER_74_195 ();
 sg13g2_fill_2 FILLER_74_165 ();
 sg13g2_fill_1 FILLER_74_147 ();
 sg13g2_fill_1 FILLER_74_123 ();
 sg13g2_fill_2 FILLER_74_121 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_73_407 ();
 sg13g2_fill_2 FILLER_73_327 ();
 sg13g2_fill_2 FILLER_73_281 ();
 sg13g2_fill_2 FILLER_73_271 ();
 sg13g2_fill_2 FILLER_73_244 ();
 sg13g2_fill_1 FILLER_73_210 ();
 sg13g2_fill_2 FILLER_73_208 ();
 sg13g2_fill_1 FILLER_73_122 ();
 sg13g2_fill_1 FILLER_73_111 ();
 sg13g2_decap_4 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_72_407 ();
 sg13g2_fill_1 FILLER_72_375 ();
 sg13g2_fill_1 FILLER_72_340 ();
 sg13g2_fill_1 FILLER_72_254 ();
 sg13g2_fill_1 FILLER_72_136 ();
 sg13g2_fill_2 FILLER_72_134 ();
 sg13g2_fill_1 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_fill_1 FILLER_71_377 ();
 sg13g2_fill_1 FILLER_71_320 ();
 sg13g2_fill_1 FILLER_71_222 ();
 sg13g2_fill_2 FILLER_71_174 ();
 sg13g2_fill_1 FILLER_71_131 ();
 sg13g2_fill_2 FILLER_71_129 ();
 sg13g2_fill_1 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_70_407 ();
 sg13g2_fill_1 FILLER_70_401 ();
 sg13g2_fill_2 FILLER_70_312 ();
 sg13g2_fill_1 FILLER_70_226 ();
 sg13g2_fill_2 FILLER_70_215 ();
 sg13g2_fill_2 FILLER_70_174 ();
 sg13g2_fill_1 FILLER_70_150 ();
 sg13g2_fill_2 FILLER_70_120 ();
 sg13g2_fill_1 FILLER_70_32 ();
 sg13g2_decap_4 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_fill_2 FILLER_69_378 ();
 sg13g2_fill_1 FILLER_69_360 ();
 sg13g2_fill_2 FILLER_69_349 ();
 sg13g2_fill_2 FILLER_69_326 ();
 sg13g2_fill_1 FILLER_69_180 ();
 sg13g2_fill_2 FILLER_69_173 ();
 sg13g2_fill_2 FILLER_69_164 ();
 sg13g2_fill_2 FILLER_69_151 ();
 sg13g2_fill_2 FILLER_69_144 ();
 sg13g2_fill_1 FILLER_69_139 ();
 sg13g2_fill_1 FILLER_69_69 ();
 sg13g2_fill_2 FILLER_69_67 ();
 sg13g2_fill_1 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_68_389 ();
 sg13g2_fill_2 FILLER_68_373 ();
 sg13g2_fill_2 FILLER_68_343 ();
 sg13g2_fill_2 FILLER_68_332 ();
 sg13g2_fill_1 FILLER_68_313 ();
 sg13g2_fill_2 FILLER_68_284 ();
 sg13g2_fill_2 FILLER_68_227 ();
 sg13g2_fill_1 FILLER_68_147 ();
 sg13g2_fill_2 FILLER_68_140 ();
 sg13g2_fill_2 FILLER_68_124 ();
 sg13g2_fill_1 FILLER_68_68 ();
 sg13g2_fill_2 FILLER_68_44 ();
 sg13g2_fill_2 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_67_280 ();
 sg13g2_fill_1 FILLER_67_170 ();
 sg13g2_fill_1 FILLER_67_109 ();
 sg13g2_fill_2 FILLER_67_91 ();
 sg13g2_fill_1 FILLER_67_81 ();
 sg13g2_fill_2 FILLER_67_79 ();
 sg13g2_fill_1 FILLER_67_53 ();
 sg13g2_fill_1 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_66_375 ();
 sg13g2_fill_1 FILLER_66_330 ();
 sg13g2_fill_2 FILLER_66_236 ();
 sg13g2_fill_1 FILLER_66_178 ();
 sg13g2_fill_1 FILLER_66_94 ();
 sg13g2_fill_2 FILLER_66_92 ();
 sg13g2_fill_1 FILLER_66_47 ();
 sg13g2_decap_4 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_65_388 ();
 sg13g2_fill_2 FILLER_65_329 ();
 sg13g2_fill_1 FILLER_65_323 ();
 sg13g2_fill_2 FILLER_65_288 ();
 sg13g2_fill_1 FILLER_65_275 ();
 sg13g2_fill_1 FILLER_65_220 ();
 sg13g2_fill_1 FILLER_65_210 ();
 sg13g2_fill_2 FILLER_65_195 ();
 sg13g2_fill_1 FILLER_65_189 ();
 sg13g2_fill_2 FILLER_65_177 ();
 sg13g2_fill_1 FILLER_65_171 ();
 sg13g2_fill_1 FILLER_65_151 ();
 sg13g2_fill_1 FILLER_65_127 ();
 sg13g2_fill_1 FILLER_65_98 ();
 sg13g2_fill_2 FILLER_65_25 ();
 sg13g2_decap_4 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_fill_2 FILLER_64_393 ();
 sg13g2_fill_1 FILLER_64_285 ();
 sg13g2_fill_2 FILLER_64_283 ();
 sg13g2_fill_1 FILLER_64_210 ();
 sg13g2_fill_2 FILLER_64_184 ();
 sg13g2_fill_2 FILLER_64_150 ();
 sg13g2_fill_2 FILLER_64_142 ();
 sg13g2_fill_1 FILLER_64_124 ();
 sg13g2_fill_2 FILLER_64_65 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_63_384 ();
 sg13g2_fill_1 FILLER_63_302 ();
 sg13g2_fill_2 FILLER_63_251 ();
 sg13g2_fill_1 FILLER_63_232 ();
 sg13g2_fill_1 FILLER_63_128 ();
 sg13g2_fill_1 FILLER_63_109 ();
 sg13g2_fill_1 FILLER_63_88 ();
 sg13g2_fill_1 FILLER_63_63 ();
 sg13g2_fill_1 FILLER_63_26 ();
 sg13g2_fill_1 FILLER_63_11 ();
 sg13g2_decap_4 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_fill_2 FILLER_62_394 ();
 sg13g2_fill_1 FILLER_62_384 ();
 sg13g2_fill_1 FILLER_62_324 ();
 sg13g2_fill_1 FILLER_62_286 ();
 sg13g2_fill_2 FILLER_62_240 ();
 sg13g2_fill_1 FILLER_62_235 ();
 sg13g2_fill_1 FILLER_62_170 ();
 sg13g2_fill_1 FILLER_62_161 ();
 sg13g2_fill_1 FILLER_62_133 ();
 sg13g2_fill_2 FILLER_62_110 ();
 sg13g2_fill_1 FILLER_62_96 ();
 sg13g2_fill_1 FILLER_62_36 ();
 sg13g2_fill_1 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_61_308 ();
 sg13g2_fill_2 FILLER_61_306 ();
 sg13g2_fill_1 FILLER_61_281 ();
 sg13g2_fill_2 FILLER_61_224 ();
 sg13g2_fill_1 FILLER_61_207 ();
 sg13g2_fill_1 FILLER_61_189 ();
 sg13g2_fill_1 FILLER_61_180 ();
 sg13g2_fill_2 FILLER_61_170 ();
 sg13g2_fill_1 FILLER_61_156 ();
 sg13g2_fill_1 FILLER_61_122 ();
 sg13g2_fill_1 FILLER_61_103 ();
 sg13g2_fill_1 FILLER_61_65 ();
 sg13g2_fill_2 FILLER_61_63 ();
 sg13g2_fill_2 FILLER_61_34 ();
 sg13g2_fill_1 FILLER_61_2 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_60_348 ();
 sg13g2_fill_1 FILLER_60_318 ();
 sg13g2_fill_2 FILLER_60_253 ();
 sg13g2_fill_2 FILLER_60_210 ();
 sg13g2_fill_2 FILLER_60_190 ();
 sg13g2_fill_2 FILLER_60_180 ();
 sg13g2_fill_1 FILLER_60_174 ();
 sg13g2_fill_2 FILLER_60_131 ();
 sg13g2_fill_2 FILLER_60_108 ();
 sg13g2_fill_2 FILLER_60_101 ();
 sg13g2_fill_2 FILLER_60_58 ();
 sg13g2_fill_2 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_59_381 ();
 sg13g2_fill_1 FILLER_59_375 ();
 sg13g2_fill_1 FILLER_59_357 ();
 sg13g2_fill_1 FILLER_59_316 ();
 sg13g2_fill_2 FILLER_59_314 ();
 sg13g2_fill_2 FILLER_59_255 ();
 sg13g2_fill_1 FILLER_59_168 ();
 sg13g2_fill_1 FILLER_59_105 ();
 sg13g2_fill_1 FILLER_59_34 ();
 sg13g2_fill_2 FILLER_58_357 ();
 sg13g2_fill_1 FILLER_58_320 ();
 sg13g2_fill_2 FILLER_58_296 ();
 sg13g2_fill_2 FILLER_58_289 ();
 sg13g2_fill_2 FILLER_58_265 ();
 sg13g2_fill_1 FILLER_58_244 ();
 sg13g2_fill_1 FILLER_58_231 ();
 sg13g2_fill_2 FILLER_58_184 ();
 sg13g2_fill_1 FILLER_58_138 ();
 sg13g2_fill_1 FILLER_58_107 ();
 sg13g2_fill_1 FILLER_58_60 ();
 sg13g2_fill_2 FILLER_58_58 ();
 sg13g2_fill_1 FILLER_58_25 ();
 sg13g2_fill_1 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_fill_1 FILLER_57_320 ();
 sg13g2_fill_2 FILLER_57_217 ();
 sg13g2_fill_2 FILLER_57_110 ();
 sg13g2_fill_1 FILLER_57_30 ();
 sg13g2_fill_1 FILLER_57_2 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_fill_1 FILLER_56_399 ();
 sg13g2_fill_2 FILLER_56_343 ();
 sg13g2_fill_2 FILLER_56_327 ();
 sg13g2_fill_2 FILLER_56_288 ();
 sg13g2_fill_2 FILLER_56_201 ();
 sg13g2_fill_2 FILLER_56_179 ();
 sg13g2_fill_2 FILLER_56_147 ();
 sg13g2_fill_1 FILLER_56_131 ();
 sg13g2_fill_2 FILLER_56_81 ();
 sg13g2_fill_1 FILLER_56_43 ();
 sg13g2_fill_2 FILLER_56_41 ();
 sg13g2_fill_1 FILLER_56_31 ();
 sg13g2_fill_1 FILLER_55_280 ();
 sg13g2_fill_2 FILLER_55_273 ();
 sg13g2_fill_1 FILLER_55_205 ();
 sg13g2_fill_2 FILLER_55_203 ();
 sg13g2_fill_2 FILLER_55_187 ();
 sg13g2_fill_1 FILLER_55_173 ();
 sg13g2_fill_1 FILLER_55_158 ();
 sg13g2_fill_2 FILLER_55_150 ();
 sg13g2_fill_1 FILLER_55_134 ();
 sg13g2_fill_2 FILLER_55_120 ();
 sg13g2_fill_1 FILLER_55_63 ();
 sg13g2_fill_1 FILLER_55_53 ();
 sg13g2_fill_1 FILLER_55_35 ();
 sg13g2_fill_2 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_54_407 ();
 sg13g2_fill_1 FILLER_54_337 ();
 sg13g2_fill_1 FILLER_54_318 ();
 sg13g2_fill_1 FILLER_54_257 ();
 sg13g2_fill_2 FILLER_54_239 ();
 sg13g2_fill_1 FILLER_54_174 ();
 sg13g2_fill_1 FILLER_54_152 ();
 sg13g2_fill_1 FILLER_54_140 ();
 sg13g2_fill_1 FILLER_54_121 ();
 sg13g2_fill_1 FILLER_54_104 ();
 sg13g2_fill_1 FILLER_54_89 ();
 sg13g2_fill_1 FILLER_54_65 ();
 sg13g2_fill_2 FILLER_54_63 ();
 sg13g2_fill_1 FILLER_54_2 ();
 sg13g2_fill_2 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_53_407 ();
 sg13g2_fill_1 FILLER_53_398 ();
 sg13g2_fill_2 FILLER_53_396 ();
 sg13g2_fill_2 FILLER_53_321 ();
 sg13g2_fill_1 FILLER_53_280 ();
 sg13g2_fill_2 FILLER_53_251 ();
 sg13g2_fill_2 FILLER_53_136 ();
 sg13g2_fill_1 FILLER_53_122 ();
 sg13g2_fill_1 FILLER_53_113 ();
 sg13g2_fill_2 FILLER_53_111 ();
 sg13g2_fill_1 FILLER_53_70 ();
 sg13g2_fill_2 FILLER_53_68 ();
 sg13g2_fill_1 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_fill_2 FILLER_52_406 ();
 sg13g2_fill_2 FILLER_52_348 ();
 sg13g2_fill_1 FILLER_52_307 ();
 sg13g2_fill_1 FILLER_52_292 ();
 sg13g2_fill_1 FILLER_52_251 ();
 sg13g2_fill_1 FILLER_52_244 ();
 sg13g2_fill_2 FILLER_52_215 ();
 sg13g2_fill_1 FILLER_52_205 ();
 sg13g2_fill_2 FILLER_52_168 ();
 sg13g2_fill_1 FILLER_52_135 ();
 sg13g2_fill_2 FILLER_52_32 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_decap_4 FILLER_51_403 ();
 sg13g2_fill_2 FILLER_51_397 ();
 sg13g2_fill_1 FILLER_51_277 ();
 sg13g2_fill_2 FILLER_51_266 ();
 sg13g2_fill_2 FILLER_51_216 ();
 sg13g2_fill_1 FILLER_51_113 ();
 sg13g2_fill_2 FILLER_51_81 ();
 sg13g2_fill_1 FILLER_51_2 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_50_401 ();
 sg13g2_decap_8 FILLER_50_394 ();
 sg13g2_decap_8 FILLER_50_387 ();
 sg13g2_fill_2 FILLER_50_340 ();
 sg13g2_fill_1 FILLER_50_306 ();
 sg13g2_fill_1 FILLER_50_266 ();
 sg13g2_fill_2 FILLER_50_264 ();
 sg13g2_fill_1 FILLER_50_249 ();
 sg13g2_fill_1 FILLER_50_189 ();
 sg13g2_fill_2 FILLER_50_174 ();
 sg13g2_fill_1 FILLER_50_155 ();
 sg13g2_fill_2 FILLER_50_153 ();
 sg13g2_fill_2 FILLER_50_89 ();
 sg13g2_fill_1 FILLER_50_47 ();
 sg13g2_fill_2 FILLER_50_45 ();
 sg13g2_fill_1 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_49_407 ();
 sg13g2_decap_4 FILLER_49_403 ();
 sg13g2_decap_8 FILLER_49_396 ();
 sg13g2_decap_8 FILLER_49_389 ();
 sg13g2_decap_8 FILLER_49_382 ();
 sg13g2_fill_2 FILLER_49_376 ();
 sg13g2_decap_4 FILLER_49_372 ();
 sg13g2_fill_1 FILLER_49_321 ();
 sg13g2_fill_1 FILLER_49_315 ();
 sg13g2_fill_1 FILLER_49_245 ();
 sg13g2_fill_2 FILLER_49_227 ();
 sg13g2_fill_1 FILLER_49_188 ();
 sg13g2_fill_2 FILLER_49_173 ();
 sg13g2_fill_2 FILLER_49_149 ();
 sg13g2_fill_1 FILLER_49_107 ();
 sg13g2_fill_2 FILLER_49_105 ();
 sg13g2_fill_1 FILLER_49_77 ();
 sg13g2_fill_2 FILLER_49_75 ();
 sg13g2_fill_1 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_48_407 ();
 sg13g2_decap_8 FILLER_48_400 ();
 sg13g2_decap_8 FILLER_48_393 ();
 sg13g2_decap_8 FILLER_48_386 ();
 sg13g2_decap_8 FILLER_48_379 ();
 sg13g2_decap_8 FILLER_48_372 ();
 sg13g2_decap_8 FILLER_48_365 ();
 sg13g2_fill_1 FILLER_48_317 ();
 sg13g2_fill_2 FILLER_48_224 ();
 sg13g2_fill_2 FILLER_48_124 ();
 sg13g2_fill_2 FILLER_48_18 ();
 sg13g2_decap_4 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_4 FILLER_47_405 ();
 sg13g2_decap_8 FILLER_47_398 ();
 sg13g2_decap_8 FILLER_47_391 ();
 sg13g2_decap_8 FILLER_47_384 ();
 sg13g2_decap_8 FILLER_47_377 ();
 sg13g2_decap_8 FILLER_47_370 ();
 sg13g2_decap_8 FILLER_47_363 ();
 sg13g2_decap_8 FILLER_47_356 ();
 sg13g2_fill_2 FILLER_47_300 ();
 sg13g2_fill_1 FILLER_47_286 ();
 sg13g2_fill_2 FILLER_47_284 ();
 sg13g2_fill_1 FILLER_47_248 ();
 sg13g2_fill_2 FILLER_47_233 ();
 sg13g2_fill_1 FILLER_47_223 ();
 sg13g2_fill_2 FILLER_47_208 ();
 sg13g2_fill_1 FILLER_47_192 ();
 sg13g2_decap_8 FILLER_47_185 ();
 sg13g2_fill_1 FILLER_47_157 ();
 sg13g2_decap_4 FILLER_47_149 ();
 sg13g2_fill_2 FILLER_47_119 ();
 sg13g2_decap_4 FILLER_47_115 ();
 sg13g2_decap_8 FILLER_47_108 ();
 sg13g2_fill_1 FILLER_47_23 ();
 sg13g2_decap_4 FILLER_47_19 ();
 sg13g2_decap_8 FILLER_47_12 ();
 sg13g2_decap_8 FILLER_47_5 ();
 sg13g2_fill_1 FILLER_47_0 ();
 sg13g2_decap_4 FILLER_46_405 ();
 sg13g2_decap_8 FILLER_46_398 ();
 sg13g2_decap_8 FILLER_46_391 ();
 sg13g2_decap_8 FILLER_46_371 ();
 sg13g2_decap_8 FILLER_46_364 ();
 sg13g2_decap_8 FILLER_46_344 ();
 sg13g2_fill_1 FILLER_46_309 ();
 sg13g2_fill_1 FILLER_46_282 ();
 sg13g2_decap_4 FILLER_45_333 ();
 sg13g2_fill_2 FILLER_45_18 ();
 sg13g2_decap_4 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_44_407 ();
 sg13g2_decap_4 FILLER_44_403 ();
 sg13g2_decap_8 FILLER_44_396 ();
 sg13g2_decap_8 FILLER_44_389 ();
 sg13g2_decap_8 FILLER_43_5 ();
 sg13g2_fill_1 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_42_407 ();
 sg13g2_decap_8 FILLER_42_400 ();
 sg13g2_decap_8 FILLER_42_393 ();
 sg13g2_fill_2 FILLER_42_311 ();
 sg13g2_decap_4 FILLER_42_307 ();
 sg13g2_decap_8 FILLER_42_300 ();
 sg13g2_decap_4 FILLER_42_148 ();
 sg13g2_fill_2 FILLER_41_335 ();
 sg13g2_decap_4 FILLER_41_331 ();
 sg13g2_decap_8 FILLER_41_324 ();
 sg13g2_fill_2 FILLER_41_18 ();
 sg13g2_decap_4 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_fill_1 FILLER_41_2 ();
 sg13g2_fill_2 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_fill_2 FILLER_40_406 ();
 sg13g2_decap_8 FILLER_40_399 ();
 sg13g2_fill_1 FILLER_40_72 ();
 sg13g2_decap_4 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_39_335 ();
 sg13g2_decap_4 FILLER_39_331 ();
 sg13g2_decap_8 FILLER_39_324 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_decap_8 FILLER_38_396 ();
 sg13g2_decap_8 FILLER_38_389 ();
 sg13g2_decap_8 FILLER_37_5 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_decap_8 FILLER_35_5 ();
 sg13g2_fill_1 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_4 FILLER_32_403 ();
 sg13g2_decap_8 FILLER_32_396 ();
 sg13g2_decap_8 FILLER_32_389 ();
 sg13g2_fill_2 FILLER_31_335 ();
 sg13g2_decap_4 FILLER_31_331 ();
 sg13g2_decap_8 FILLER_31_324 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_4 FILLER_30_403 ();
 sg13g2_decap_8 FILLER_30_396 ();
 sg13g2_decap_8 FILLER_30_389 ();
 sg13g2_decap_8 FILLER_29_5 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_2 FILLER_28_315 ();
 sg13g2_fill_2 FILLER_28_300 ();
 sg13g2_decap_8 FILLER_27_5 ();
 sg13g2_fill_1 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_fill_1 FILLER_23_336 ();
 sg13g2_fill_2 FILLER_23_334 ();
 sg13g2_fill_1 FILLER_23_320 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_21_5 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_20_400 ();
 sg13g2_decap_8 FILLER_20_393 ();
 sg13g2_decap_8 FILLER_19_5 ();
 sg13g2_fill_1 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_18_400 ();
 sg13g2_decap_8 FILLER_18_393 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_decap_8 FILLER_13_5 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_12_400 ();
 sg13g2_decap_8 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_11_5 ();
 sg13g2_fill_1 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_6_402 ();
 sg13g2_decap_8 FILLER_5_5 ();
 sg13g2_fill_1 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_2 FILLER_3_183 ();
 sg13g2_fill_2 FILLER_3_168 ();
 sg13g2_fill_1 FILLER_3_5 ();
 sg13g2_fill_1 FILLER_3_0 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_0_401 ();
 sg13g2_dlygate4sd3_1 hold244 (.A(\game_inst.apple_inst.apple_y[1] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold243 (.A(\game_inst.control_inst.dir[1] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold242 (.A(\game_inst.control_inst.dir[1] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold241 (.A(\game_inst.vga_inst.px[8] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold240 (.A(\game_inst.apple_inst.i_snake_y[0] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0055_),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0587_),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold237 (.A(\game_inst.sound_inst.max_counter[1] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0527_),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold235 (.A(\game_inst.vga_inst.px[9] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold234 (.A(\game_inst.apple_inst.i_snake_x[2] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0311_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0307_),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold231 (.A(\game_inst.apple_inst.apple_y[1] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold230 (.A(\game_inst.apple_inst.i_snake_x[1] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold229 (.A(\game_inst.head_y[3] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold228 (.A(\game_inst.apple_inst.i_snake_x[3] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0637_),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold226 (.A(\game_inst.snake_inst.pos[5] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0006_),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold224 (.A(\game_inst.vga_inst.row_buffer[1][2] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0007_),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold222 (.A(\game_inst.vga_inst.row_buffer[2][3] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0010_),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold220 (.A(\game_inst.vga_inst.row_buffer[3][2] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0544_),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold218 (.A(\game_inst.sound_inst.max_counter[2] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold217 (.A(\game_inst.vga_inst.row_buffer[3][1] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold216 (.A(\game_inst.vga_inst.row_buffer[4][3] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold215 (.A(\game_inst.vga_inst.row_buffer[3][0] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0011_),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold213 (.A(\game_inst.vga_inst.row_buffer[3][3] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold212 (.A(\game_inst.vga_inst.row_buffer[4][0] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold211 (.A(\game_inst.vga_inst.row_buffer[5][3] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold210 (.A(\game_inst.vga_inst.px[3] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold209 (.A(\game_inst.vga_inst.row_buffer[5][2] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0005_),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold207 (.A(\game_inst.vga_inst.row_buffer[2][1] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0014_),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold205 (.A(\game_inst.vga_inst.row_buffer[4][2] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold204 (.A(\game_inst.vga_inst.row_buffer[1][0] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0008_),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold202 (.A(\game_inst.vga_inst.row_buffer[2][0] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold201 (.A(\game_inst.vga_inst.row_buffer[5][0] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold200 (.A(\game_inst.vga_inst.row_buffer[5][1] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0013_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold198 (.A(\game_inst.vga_inst.row_buffer[4][1] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold197 (.A(\game_inst.snake_inst.pos[3] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold196 (.A(\game_inst.snake_inst.pos[1] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold195 (.A(\game_inst.head_y[1] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0105_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold193 (.A(\game_inst.head_x[1] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0107_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold191 (.A(\game_inst.head_x[3] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold190 (.A(\game_inst.head_y[2] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0123_),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold188 (.A(\game_inst.apple_inst.i_snake_y[2] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0064_),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0623_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold185 (.A(\game_inst.sound_inst.max_counter[3] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0163_),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold183 (.A(\game_inst.apple_inst.i_snake_y[1] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0617_),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold181 (.A(\game_inst.sound_inst.max_counter[0] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold180 (.A(\game_inst.snake_inst.length[0] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold179 (.A(\game_inst.vga_inst.px[3] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold178 (.A(\game_inst.apple_inst.i_snake_x[4] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0124_),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold176 (.A(\game_inst.apple_inst.i_snake_y[3] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0143_),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0208_),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold173 (.A(\game_inst.tickgen_inst.counter_max[3] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0042_),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0507_),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold170 (.A(\game_inst.snake_inst.pos[6] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold169 (.A(\game_inst.vga_inst.px[5] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0109_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold167 (.A(\game_inst.head_y[0] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0106_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold165 (.A(\game_inst.head_x[2] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold164 (.A(\game_inst.sound_inst.phase[4] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0104_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold162 (.A(\game_inst.head_x[0] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold161 (.A(\game_inst.tickgen_inst.counter[1] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold160 (.A(\game_inst.snake_inst.length[5] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold159 (.A(\game_inst.head_x[4] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0127_),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold157 (.A(\game_inst.snake_inst.length[2] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0519_),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold155 (.A(\game_inst.vga_inst.px[4] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold154 (.A(\game_inst.vga_inst.py[7] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold153 (.A(\game_inst.sound_inst.phase[3] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold152 (.A(\game_inst.sound_inst.phase[2] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0142_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0203_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold149 (.A(\game_inst.tickgen_inst.counter_max[2] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0103_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold147 (.A(\game_inst.control_inst.backwards[1] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold146 (.A(\game_inst.vga_inst.py[5] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold145 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[0] [0]),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold144 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[233] [0]),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0177_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold142 (.A(\game_inst.snake_inst.length[1] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold141 (.A(\game_inst.sound_inst.counter[3] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold140 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[233] [0]),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold139 (.A(\game_inst.vga_inst.py[6] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0281_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold137 (.A(\game_inst.vga_inst.px[6] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0036_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold135 (.A(\game_inst.vga_inst.px[7] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0065_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0626_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold132 (.A(\game_inst.sound_inst.phase[0] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0102_),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold130 (.A(\game_inst.control_inst.i_head_dir[0] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0128_),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0182_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold127 (.A(\game_inst.snake_inst.length[3] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0196_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold125 (.A(\game_inst.control_inst.o_start ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0134_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0191_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold122 (.A(\game_inst.snake_inst.pos[2] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold121 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[0] [0]),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold120 (.A(\game_inst.apple_inst.random_inst.lfsr4[3] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold119 (.A(\game_inst.apple_inst.apple_y[2] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0071_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold117 (.A(\game_inst.vga_inst.row_buffer[0][0] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold116 (.A(\game_inst.sound_inst.counter[2] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold115 (.A(\game_inst.vga_inst.py[2] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0129_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0184_),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold112 (.A(\game_inst.snake_inst.length[4] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold111 (.A(\game_inst.vga_inst.row_buffer[7][1] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0074_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold109 (.A(\game_inst.vga_inst.row_buffer[0][3] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold108 (.A(\game_inst.apple_inst.apple_x[3] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0073_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold106 (.A(\game_inst.vga_inst.row_buffer[0][2] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold105 (.A(\game_inst.vga_inst.row_buffer[7][0] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0613_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold103 (.A(\game_inst.sound_inst.counter[1] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0072_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold101 (.A(\game_inst.vga_inst.row_buffer[0][1] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold100 (.A(\game_inst.vga_inst.row_buffer[7][3] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold99 (.A(\game_inst.apple_inst.apple_x[1] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold98 (.A(\game_inst.vga_inst.px[1] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold97 (.A(\game_inst.apple_inst.i_snake_valid ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0057_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0608_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold94 (.A(\game_inst.sound_inst.mode[0] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0609_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold92 (.A(\game_inst.sound_inst.mode[1] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0340_),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold90 (.A(\game_inst.snake_inst.pos[7] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0090_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold88 (.A(\game_inst.apple_inst.random_inst.lfsr5[4] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold87 (.A(\game_inst.apple_inst.apple_x[2] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0059_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0611_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold84 (.A(\game_inst.sound_inst.counter[0] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0076_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold82 (.A(\game_inst.vga_inst.py[1] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold81 (.A(\game_inst.apple_inst.o_ready ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0692_),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold79 (.A(\game_inst.apple_inst.random_inst.lfsr5[2] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold78 (.A(\game_inst.apple_inst.random_inst.lfsr5[1] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold77 (.A(\game_inst.apple_inst.random_inst.lfsr4[2] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0030_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold75 (.A(\game_inst.vga_inst.row_buffer[7][2] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0131_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0187_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold72 (.A(\game_inst.snake_inst.length[6] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0139_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold70 (.A(\game_inst.apple_inst.apple_y[3] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0086_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold68 (.A(\game_inst.apple_inst.random_inst.lfsr5[0] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0070_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold66 (.A(\game_inst.snake_inst.pos[7] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0144_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0219_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold63 (.A(\game_inst.tick ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0141_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold61 (.A(\game_inst.tickgen_inst.counter_max[1] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0097_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold59 (.A(\game_inst.apple_inst.random_inst.lfsr5[3] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold58 (.A(\game_inst.vga_inst.py[8] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0135_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0192_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold55 (.A(\game_inst.snake_inst.pos[4] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0066_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0628_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold52 (.A(\game_inst.sound_inst.phase[1] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0137_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold50 (.A(\game_inst.apple_inst.random_inst.lfsr4[1] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0226_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold48 (.A(\game_inst.tickgen_inst.counter[2] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0046_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0517_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold45 (.A(\game_inst.vga_inst.px[2] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0668_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold43 (.A(\game_inst.apple_inst.test ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold42 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[1].sreg_q[0] [0]),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0193_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold40 (.A(\game_inst.apple_inst.apple_y[0] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold39 (.A(\game_inst.vga_inst.py[0] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0099_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold37 (.A(\game_inst.apple_inst.random_inst.lfsr4[0] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0025_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0456_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold34 (.A(\game_inst.vga_inst.row_buffer[6][1] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0024_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0454_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold31 (.A(\game_inst.vga_inst.row_buffer[6][0] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0027_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0460_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold28 (.A(\game_inst.vga_inst.row_buffer[6][3] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0056_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0597_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold25 (.A(audio),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0026_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0458_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold22 (.A(\game_inst.vga_inst.row_buffer[6][2] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold21 (.A(\game_inst.snake_inst.pos[0] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0145_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold19 (.A(\game_inst.tickgen_inst.counter[0] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold18 (.A(\game_inst.vga_inst.row_buffer[8][1] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold17 (.A(\game_inst.vga_inst.row_buffer[8][3] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0037_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold15 (.A(\game_inst.vga_inst.py[9] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold14 (.A(\game_inst.vga_inst.row_buffer[8][0] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold13 (.A(\game_inst.vga_inst.py[4] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0132_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold11 (.A(\game_inst.snake_inst.length[7] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold10 (.A(\game_inst.vga_inst.row_buffer[8][2] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0002_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold8 (.A(failure),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0148_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold6 (.A(\game_inst.tickgen_inst.counter[3] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold5 (.A(\game_inst.vga_inst.px[0] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold4 (.A(\game_inst.o_vga_vsync ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold3 (.A(\game_inst.pwm_base ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold2 (.A(\game_inst.vga_inst.s_vsync ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold1 (.A(\game_inst.vga_inst.s_hsync ),
    .X(net339));
 sg13g2_inv_2 clkload4 (.A(clknet_leaf_25_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_leaf_21_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_leaf_27_clk));
 sg13g2_inv_4 clkload1 (.A(clknet_leaf_78_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_4_15_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_dlygate4sd3_1 dly2_0_0 (.A(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_q[0] [0]),
    .X(\game_inst.snake_inst.shiftreg_inst.genblk2[0].sreg_w[1] [0]));
 sg13g2_buf_8 fanout108 (.A(net109),
    .X(net108));
 sg13g2_buf_8 fanout109 (.A(_0691_),
    .X(net109));
 sg13g2_buf_8 fanout110 (.A(net112),
    .X(net110));
 sg13g2_buf_1 fanout111 (.A(net112),
    .X(net111));
 sg13g2_buf_8 fanout112 (.A(_0662_),
    .X(net112));
 sg13g2_buf_8 fanout113 (.A(_0426_),
    .X(net113));
 sg13g2_buf_8 fanout114 (.A(_0423_),
    .X(net114));
 sg13g2_buf_8 fanout115 (.A(_0420_),
    .X(net115));
 sg13g2_buf_8 fanout116 (.A(_0344_),
    .X(net116));
 sg13g2_buf_8 fanout117 (.A(_0500_),
    .X(net117));
 sg13g2_buf_8 fanout118 (.A(_0498_),
    .X(net118));
 sg13g2_buf_8 fanout119 (.A(net120),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(net122),
    .X(net120));
 sg13g2_buf_8 fanout121 (.A(net122),
    .X(net121));
 sg13g2_buf_1 fanout122 (.A(_0492_),
    .X(net122));
 sg13g2_buf_8 fanout123 (.A(net124),
    .X(net123));
 sg13g2_buf_8 fanout124 (.A(_0324_),
    .X(net124));
 sg13g2_buf_8 fanout125 (.A(net126),
    .X(net125));
 sg13g2_buf_8 fanout126 (.A(_0324_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(net128),
    .X(net127));
 sg13g2_buf_1 fanout128 (.A(net130),
    .X(net128));
 sg13g2_buf_8 fanout129 (.A(net130),
    .X(net129));
 sg13g2_buf_8 fanout130 (.A(_0323_),
    .X(net130));
 sg13g2_buf_8 fanout131 (.A(net132),
    .X(net131));
 sg13g2_buf_8 fanout132 (.A(net133),
    .X(net132));
 sg13g2_buf_8 fanout133 (.A(_0487_),
    .X(net133));
 sg13g2_buf_8 fanout134 (.A(net135),
    .X(net134));
 sg13g2_buf_8 fanout135 (.A(net380),
    .X(net135));
 sg13g2_buf_8 fanout136 (.A(net566),
    .X(net136));
 sg13g2_buf_8 fanout137 (.A(net572),
    .X(net137));
 sg13g2_buf_8 fanout138 (.A(net568),
    .X(net138));
 sg13g2_buf_8 fanout139 (.A(\game_inst.apple_inst.i_snake_x[0] ),
    .X(net139));
 sg13g2_buf_1 fanout140 (.A(\game_inst.apple_inst.i_snake_x[0] ),
    .X(net140));
 sg13g2_buf_8 fanout141 (.A(net580),
    .X(net141));
 sg13g2_buf_8 fanout142 (.A(\game_inst.vga_inst.py[6] ),
    .X(net142));
 sg13g2_buf_8 fanout143 (.A(net341),
    .X(net143));
 sg13g2_buf_8 fanout144 (.A(net573),
    .X(net144));
 sg13g2_buf_8 fanout145 (.A(net579),
    .X(net145));
 sg13g2_buf_1 fanout146 (.A(\game_inst.vga_inst.px[8] ),
    .X(net146));
 sg13g2_buf_8 fanout147 (.A(\game_inst.vga_inst.px[7] ),
    .X(net147));
 sg13g2_buf_8 fanout148 (.A(net507),
    .X(net148));
 sg13g2_buf_8 fanout149 (.A(\game_inst.vga_inst.px[4] ),
    .X(net149));
 sg13g2_buf_8 fanout150 (.A(net151),
    .X(net150));
 sg13g2_buf_8 fanout151 (.A(net153),
    .X(net151));
 sg13g2_buf_8 fanout152 (.A(net153),
    .X(net152));
 sg13g2_buf_8 fanout153 (.A(_0488_),
    .X(net153));
 sg13g2_buf_8 fanout154 (.A(_0269_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_0269_),
    .X(net155));
 sg13g2_buf_8 fanout156 (.A(rst_n),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(rst_n),
    .X(net157));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_tielo tt_um_snake_game_7 (.L_LO(net7));
 assign uio_oe[0] = net217;
 assign uio_oe[1] = net218;
 assign uio_oe[2] = net219;
 assign uio_oe[3] = net220;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_oe[7] = net221;
 assign uio_out[4] = net10;
 assign uio_out[5] = net11;
 assign uio_out[6] = net12;
endmodule
