module tt_um_sid (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire \acc[0][0] ;
 wire \acc[0][10] ;
 wire \acc[0][11] ;
 wire \acc[0][12] ;
 wire \acc[0][13] ;
 wire \acc[0][14] ;
 wire \acc[0][15] ;
 wire \acc[0][1] ;
 wire \acc[0][2] ;
 wire \acc[0][3] ;
 wire \acc[0][4] ;
 wire \acc[0][5] ;
 wire \acc[0][6] ;
 wire \acc[0][7] ;
 wire \acc[0][8] ;
 wire \acc[0][9] ;
 wire \acc[1][0] ;
 wire \acc[1][10] ;
 wire \acc[1][11] ;
 wire \acc[1][12] ;
 wire \acc[1][13] ;
 wire \acc[1][14] ;
 wire \acc[1][15] ;
 wire \acc[1][1] ;
 wire \acc[1][2] ;
 wire \acc[1][3] ;
 wire \acc[1][4] ;
 wire \acc[1][5] ;
 wire \acc[1][6] ;
 wire \acc[1][7] ;
 wire \acc[1][8] ;
 wire \acc[1][9] ;
 wire \acc[2][0] ;
 wire \acc[2][10] ;
 wire \acc[2][11] ;
 wire \acc[2][12] ;
 wire \acc[2][13] ;
 wire \acc[2][14] ;
 wire \acc[2][15] ;
 wire \acc[2][1] ;
 wire \acc[2][2] ;
 wire \acc[2][3] ;
 wire \acc[2][4] ;
 wire \acc[2][5] ;
 wire \acc[2][6] ;
 wire \acc[2][7] ;
 wire \acc[2][8] ;
 wire \acc[2][9] ;
 wire \adsr_pre_hi[10] ;
 wire \adsr_pre_hi[11] ;
 wire \adsr_pre_hi[12] ;
 wire \adsr_pre_hi[13] ;
 wire \adsr_pre_hi[1] ;
 wire \adsr_pre_hi[2] ;
 wire \adsr_pre_hi[3] ;
 wire \adsr_pre_hi[4] ;
 wire \adsr_pre_hi[5] ;
 wire \adsr_pre_hi[6] ;
 wire \adsr_pre_hi[7] ;
 wire \adsr_pre_hi[8] ;
 wire \adsr_pre_hi[9] ;
 wire \ast[0][0] ;
 wire \ast[0][1] ;
 wire \ast[1][0] ;
 wire \ast[1][1] ;
 wire \ast[2][0] ;
 wire \ast[2][1] ;
 wire \attack_reg[0][0] ;
 wire \attack_reg[0][1] ;
 wire \attack_reg[0][2] ;
 wire \attack_reg[0][3] ;
 wire \attack_reg[0][4] ;
 wire \attack_reg[0][5] ;
 wire \attack_reg[0][6] ;
 wire \attack_reg[0][7] ;
 wire \attack_reg[1][0] ;
 wire \attack_reg[1][1] ;
 wire \attack_reg[1][2] ;
 wire \attack_reg[1][3] ;
 wire \attack_reg[1][4] ;
 wire \attack_reg[1][5] ;
 wire \attack_reg[1][6] ;
 wire \attack_reg[1][7] ;
 wire \attack_reg[2][0] ;
 wire \attack_reg[2][1] ;
 wire \attack_reg[2][2] ;
 wire \attack_reg[2][3] ;
 wire \attack_reg[2][4] ;
 wire \attack_reg[2][5] ;
 wire \attack_reg[2][6] ;
 wire \attack_reg[2][7] ;
 wire cur_gate;
 wire \env[0][0] ;
 wire \env[0][1] ;
 wire \env[0][2] ;
 wire \env[0][3] ;
 wire \env[0][4] ;
 wire \env[0][5] ;
 wire \env[0][6] ;
 wire \env[0][7] ;
 wire \env[1][0] ;
 wire \env[1][1] ;
 wire \env[1][2] ;
 wire \env[1][3] ;
 wire \env[1][4] ;
 wire \env[1][5] ;
 wire \env[1][6] ;
 wire \env[1][7] ;
 wire \env[2][0] ;
 wire \env[2][1] ;
 wire \env[2][2] ;
 wire \env[2][3] ;
 wire \env[2][4] ;
 wire \env[2][5] ;
 wire \env[2][6] ;
 wire \env[2][7] ;
 wire \freq[0][0] ;
 wire \freq[0][1] ;
 wire \freq[0][2] ;
 wire \freq[0][3] ;
 wire \freq[0][4] ;
 wire \freq[0][5] ;
 wire \freq[0][6] ;
 wire \freq[0][7] ;
 wire \freq[1][0] ;
 wire \freq[1][1] ;
 wire \freq[1][2] ;
 wire \freq[1][3] ;
 wire \freq[1][4] ;
 wire \freq[1][5] ;
 wire \freq[1][6] ;
 wire \freq[1][7] ;
 wire \freq[2][0] ;
 wire \freq[2][1] ;
 wire \freq[2][2] ;
 wire \freq[2][3] ;
 wire \freq[2][4] ;
 wire \freq[2][5] ;
 wire \freq[2][6] ;
 wire \freq[2][7] ;
 wire \gate_latch[0] ;
 wire \gate_latch[1] ;
 wire \gate_latch[2] ;
 wire \mix_acc[0] ;
 wire \mix_acc[1] ;
 wire \mix_acc[2] ;
 wire \mix_acc[3] ;
 wire \mix_acc[4] ;
 wire \mix_acc[5] ;
 wire \mix_acc[6] ;
 wire \mix_acc[7] ;
 wire \mix_acc[8] ;
 wire \mix_acc[9] ;
 wire \mix_out[0] ;
 wire \mix_out[1] ;
 wire \mix_out[2] ;
 wire \mix_out[3] ;
 wire \mix_out[4] ;
 wire \mix_out[5] ;
 wire \mix_out[6] ;
 wire \mix_out[7] ;
 wire noise_clk_d;
 wire \p_acc[0] ;
 wire \p_acc[10] ;
 wire \p_acc[11] ;
 wire \p_acc[12] ;
 wire \p_acc[13] ;
 wire \p_acc[14] ;
 wire \p_acc[15] ;
 wire \p_acc[1] ;
 wire \p_acc[2] ;
 wire \p_acc[3] ;
 wire \p_acc[4] ;
 wire \p_acc[5] ;
 wire \p_acc[6] ;
 wire \p_acc[7] ;
 wire \p_acc[8] ;
 wire \p_acc[9] ;
 wire \p_ast[0] ;
 wire \p_ast[1] ;
 wire \p_attack[0] ;
 wire \p_attack[1] ;
 wire \p_attack[2] ;
 wire \p_attack[3] ;
 wire \p_attack[4] ;
 wire \p_attack[5] ;
 wire \p_attack[6] ;
 wire \p_attack[7] ;
 wire \p_env[0] ;
 wire \p_env[1] ;
 wire \p_env[2] ;
 wire \p_env[3] ;
 wire \p_env[4] ;
 wire \p_env[5] ;
 wire \p_env[6] ;
 wire \p_env[7] ;
 wire \p_freq[0] ;
 wire \p_freq[1] ;
 wire \p_freq[2] ;
 wire \p_freq[3] ;
 wire \p_freq[4] ;
 wire \p_freq[5] ;
 wire \p_freq[6] ;
 wire \p_freq[7] ;
 wire p_gate_latch;
 wire p_prev_msb_d;
 wire \p_pw[0] ;
 wire \p_pw[1] ;
 wire \p_pw[2] ;
 wire \p_pw[3] ;
 wire \p_pw[4] ;
 wire \p_pw[5] ;
 wire \p_pw[6] ;
 wire \p_pw[7] ;
 wire p_releasing;
 wire \p_sustain[0] ;
 wire \p_sustain[1] ;
 wire \p_sustain[2] ;
 wire \p_sustain[3] ;
 wire \p_sustain[4] ;
 wire \p_sustain[5] ;
 wire \p_sustain[6] ;
 wire \p_sustain[7] ;
 wire \p_waveform[1] ;
 wire \p_waveform[2] ;
 wire \p_waveform[3] ;
 wire \p_waveform[4] ;
 wire \p_waveform[5] ;
 wire \p_waveform[6] ;
 wire \p_waveform[7] ;
 wire \prev_msb_d[0] ;
 wire \prev_msb_d[1] ;
 wire \prev_msb_d[2] ;
 wire \pw_reg[0][0] ;
 wire \pw_reg[0][1] ;
 wire \pw_reg[0][2] ;
 wire \pw_reg[0][3] ;
 wire \pw_reg[0][4] ;
 wire \pw_reg[0][5] ;
 wire \pw_reg[0][6] ;
 wire \pw_reg[0][7] ;
 wire \pw_reg[1][0] ;
 wire \pw_reg[1][1] ;
 wire \pw_reg[1][2] ;
 wire \pw_reg[1][3] ;
 wire \pw_reg[1][4] ;
 wire \pw_reg[1][5] ;
 wire \pw_reg[1][6] ;
 wire \pw_reg[1][7] ;
 wire \pw_reg[2][0] ;
 wire \pw_reg[2][1] ;
 wire \pw_reg[2][2] ;
 wire \pw_reg[2][3] ;
 wire \pw_reg[2][4] ;
 wire \pw_reg[2][5] ;
 wire \pw_reg[2][6] ;
 wire \pw_reg[2][7] ;
 wire pwm_out;
 wire \releasing[0] ;
 wire \releasing[1] ;
 wire \releasing[2] ;
 wire net1;
 wire \slot[0] ;
 wire \slot[1] ;
 wire \slot[2] ;
 wire \sustain_reg[0][0] ;
 wire \sustain_reg[0][1] ;
 wire \sustain_reg[0][2] ;
 wire \sustain_reg[0][3] ;
 wire \sustain_reg[0][4] ;
 wire \sustain_reg[0][5] ;
 wire \sustain_reg[0][6] ;
 wire \sustain_reg[0][7] ;
 wire \sustain_reg[1][0] ;
 wire \sustain_reg[1][1] ;
 wire \sustain_reg[1][2] ;
 wire \sustain_reg[1][3] ;
 wire \sustain_reg[1][4] ;
 wire \sustain_reg[1][5] ;
 wire \sustain_reg[1][6] ;
 wire \sustain_reg[1][7] ;
 wire \sustain_reg[2][0] ;
 wire \sustain_reg[2][1] ;
 wire \sustain_reg[2][2] ;
 wire \sustain_reg[2][3] ;
 wire \sustain_reg[2][4] ;
 wire \sustain_reg[2][5] ;
 wire \sustain_reg[2][6] ;
 wire \sustain_reg[2][7] ;
 wire \u_pwm.count[0] ;
 wire \u_pwm.count[1] ;
 wire \u_pwm.count[2] ;
 wire \u_pwm.count[3] ;
 wire \u_pwm.count[4] ;
 wire \u_pwm.count[5] ;
 wire \u_pwm.count[6] ;
 wire \u_pwm.count[7] ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire \waveform[0][0] ;
 wire \waveform[0][1] ;
 wire \waveform[0][2] ;
 wire \waveform[0][3] ;
 wire \waveform[0][4] ;
 wire \waveform[0][5] ;
 wire \waveform[0][6] ;
 wire \waveform[0][7] ;
 wire \waveform[1][0] ;
 wire \waveform[1][1] ;
 wire \waveform[1][2] ;
 wire \waveform[1][3] ;
 wire \waveform[1][4] ;
 wire \waveform[1][5] ;
 wire \waveform[1][6] ;
 wire \waveform[1][7] ;
 wire \waveform[2][0] ;
 wire \waveform[2][1] ;
 wire \waveform[2][2] ;
 wire \waveform[2][3] ;
 wire \waveform[2][4] ;
 wire \waveform[2][5] ;
 wire \waveform[2][6] ;
 wire \waveform[2][7] ;
 wire wr_en_d;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;

 sg13g2_inv_1 _1451_ (.Y(_1160_),
    .A(net416));
 sg13g2_inv_1 _1452_ (.Y(_1161_),
    .A(net626));
 sg13g2_inv_1 _1453_ (.Y(_1162_),
    .A(net648));
 sg13g2_inv_1 _1454_ (.Y(_1163_),
    .A(net659));
 sg13g2_inv_1 _1455_ (.Y(_1164_),
    .A(net641));
 sg13g2_inv_1 _1456_ (.Y(_1165_),
    .A(net656));
 sg13g2_inv_1 _1457_ (.Y(_1166_),
    .A(net655));
 sg13g2_inv_1 _1458_ (.Y(_1167_),
    .A(net589));
 sg13g2_inv_1 _1459_ (.Y(_1168_),
    .A(net685));
 sg13g2_inv_1 _1460_ (.Y(_1169_),
    .A(net542));
 sg13g2_inv_1 _1461_ (.Y(_1170_),
    .A(net479));
 sg13g2_inv_1 _1462_ (.Y(_1171_),
    .A(net601));
 sg13g2_inv_1 _1463_ (.Y(_1172_),
    .A(net654));
 sg13g2_inv_1 _1464_ (.Y(_1173_),
    .A(net451));
 sg13g2_inv_1 _1465_ (.Y(_1174_),
    .A(net646));
 sg13g2_inv_1 _1466_ (.Y(_1175_),
    .A(net637));
 sg13g2_inv_1 _1467_ (.Y(_1176_),
    .A(net604));
 sg13g2_inv_1 _1468_ (.Y(_1177_),
    .A(net624));
 sg13g2_inv_1 _1469_ (.Y(_1178_),
    .A(net583));
 sg13g2_inv_1 _1470_ (.Y(_1179_),
    .A(net649));
 sg13g2_inv_1 _1471_ (.Y(_1180_),
    .A(net670));
 sg13g2_inv_1 _1472_ (.Y(_1181_),
    .A(net661));
 sg13g2_inv_1 _1473_ (.Y(_1182_),
    .A(net476));
 sg13g2_inv_1 _1474_ (.Y(_1183_),
    .A(net618));
 sg13g2_inv_1 _1475_ (.Y(_1184_),
    .A(net577));
 sg13g2_inv_1 _1476_ (.Y(_1185_),
    .A(net348));
 sg13g2_inv_1 _1477_ (.Y(_1186_),
    .A(net684));
 sg13g2_inv_1 _1478_ (.Y(_1187_),
    .A(net396));
 sg13g2_inv_1 _1479_ (.Y(_1188_),
    .A(net136));
 sg13g2_inv_1 _1480_ (.Y(_1189_),
    .A(net147));
 sg13g2_inv_1 _1481_ (.Y(_1190_),
    .A(net678));
 sg13g2_inv_1 _1482_ (.Y(_1191_),
    .A(net671));
 sg13g2_inv_1 _1483_ (.Y(_1192_),
    .A(net137));
 sg13g2_inv_1 _1484_ (.Y(_1193_),
    .A(net711));
 sg13g2_inv_1 _1485_ (.Y(_1194_),
    .A(net138));
 sg13g2_inv_1 _1486_ (.Y(_1195_),
    .A(net665));
 sg13g2_inv_1 _1487_ (.Y(_1196_),
    .A(net660));
 sg13g2_inv_1 _1488_ (.Y(_1197_),
    .A(net139));
 sg13g2_inv_1 _1489_ (.Y(_1198_),
    .A(net632));
 sg13g2_inv_1 _1490_ (.Y(_1199_),
    .A(net140));
 sg13g2_inv_1 _1491_ (.Y(_1200_),
    .A(net141));
 sg13g2_inv_1 _1492_ (.Y(_1201_),
    .A(net707));
 sg13g2_inv_1 _1493_ (.Y(_1202_),
    .A(\adsr_pre_hi[5] ));
 sg13g2_inv_1 _1494_ (.Y(_0012_),
    .A(net316));
 sg13g2_inv_1 _1495_ (.Y(_1203_),
    .A(net697));
 sg13g2_inv_1 _1496_ (.Y(_1204_),
    .A(\p_attack[4] ));
 sg13g2_inv_1 _1497_ (.Y(_1205_),
    .A(net633));
 sg13g2_inv_1 _1498_ (.Y(_1206_),
    .A(net584));
 sg13g2_inv_1 _1499_ (.Y(_1207_),
    .A(net599));
 sg13g2_inv_1 _1500_ (.Y(_1208_),
    .A(net682));
 sg13g2_inv_1 _1501_ (.Y(_1209_),
    .A(net677));
 sg13g2_inv_1 _1502_ (.Y(_1210_),
    .A(\p_attack[0] ));
 sg13g2_inv_1 _1503_ (.Y(_1211_),
    .A(net691));
 sg13g2_inv_1 _1504_ (.Y(_1212_),
    .A(net726));
 sg13g2_inv_1 _1505_ (.Y(_1213_),
    .A(net640));
 sg13g2_inv_1 _1506_ (.Y(_1214_),
    .A(net609));
 sg13g2_inv_1 _1507_ (.Y(_1215_),
    .A(net135));
 sg13g2_inv_1 _1508_ (.Y(_1216_),
    .A(\p_attack[1] ));
 sg13g2_inv_1 _1509_ (.Y(_1217_),
    .A(\p_attack[2] ));
 sg13g2_inv_1 _1510_ (.Y(_1218_),
    .A(\p_attack[3] ));
 sg13g2_inv_1 _1511_ (.Y(_1219_),
    .A(net342));
 sg13g2_inv_1 _1512_ (.Y(_1220_),
    .A(net131));
 sg13g2_inv_1 _1513_ (.Y(_1221_),
    .A(net5));
 sg13g2_inv_1 _1514_ (.Y(_1222_),
    .A(net7));
 sg13g2_inv_1 _1515_ (.Y(_1223_),
    .A(net4));
 sg13g2_inv_1 _1516_ (.Y(_1224_),
    .A(net2));
 sg13g2_inv_1 _1517_ (.Y(_1225_),
    .A(net352));
 sg13g2_inv_1 _1518_ (.Y(_1226_),
    .A(net692));
 sg13g2_inv_1 _1519_ (.Y(_1227_),
    .A(\u_pwm.count[2] ));
 sg13g2_inv_1 _1520_ (.Y(_1228_),
    .A(net628));
 sg13g2_inv_1 _1521_ (.Y(_1229_),
    .A(net695));
 sg13g2_inv_1 _1522_ (.Y(_1230_),
    .A(net331));
 sg13g2_inv_1 _1523_ (.Y(_1231_),
    .A(net727));
 sg13g2_inv_1 _1524_ (.Y(_1232_),
    .A(net146));
 sg13g2_inv_1 _1525_ (.Y(_1233_),
    .A(net645));
 sg13g2_inv_1 _1526_ (.Y(_1234_),
    .A(net657));
 sg13g2_inv_1 _1527_ (.Y(_1235_),
    .A(net492));
 sg13g2_inv_1 _1528_ (.Y(_1236_),
    .A(net565));
 sg13g2_inv_1 _1529_ (.Y(_1237_),
    .A(\p_pw[3] ));
 sg13g2_inv_1 _1530_ (.Y(_1238_),
    .A(\p_pw[2] ));
 sg13g2_inv_1 _1531_ (.Y(_1239_),
    .A(net686));
 sg13g2_inv_1 _1532_ (.Y(_1240_),
    .A(net362));
 sg13g2_inv_1 _1533_ (.Y(_1241_),
    .A(net145));
 sg13g2_inv_1 _1534_ (.Y(_1242_),
    .A(net142));
 sg13g2_inv_1 _1535_ (.Y(_1243_),
    .A(net358));
 sg13g2_inv_1 _1536_ (.Y(_1244_),
    .A(net688));
 sg13g2_inv_1 _1537_ (.Y(_1245_),
    .A(net703));
 sg13g2_inv_1 _1538_ (.Y(_1246_),
    .A(net708));
 sg13g2_inv_1 _1539_ (.Y(_1247_),
    .A(net712));
 sg13g2_inv_1 _1540_ (.Y(_1248_),
    .A(net369));
 sg13g2_inv_1 _1541_ (.Y(_1249_),
    .A(net311));
 sg13g2_inv_1 _1542_ (.Y(_1250_),
    .A(net730));
 sg13g2_inv_1 _1543_ (.Y(_1251_),
    .A(net538));
 sg13g2_inv_1 _1544_ (.Y(_1252_),
    .A(net548));
 sg13g2_inv_1 _1545_ (.Y(_1253_),
    .A(net335));
 sg13g2_inv_1 _1546_ (.Y(_1254_),
    .A(net519));
 sg13g2_nand2_1 _1547_ (.Y(_1255_),
    .A(net316),
    .B(net261));
 sg13g2_xor2_1 _1548_ (.B(net261),
    .A(net733),
    .X(_0016_));
 sg13g2_nand3_1 _1549_ (.B(\adsr_pre_hi[1] ),
    .C(\adsr_pre_hi[2] ),
    .A(\adsr_pre_hi[3] ),
    .Y(_1256_));
 sg13g2_xnor2_1 _1550_ (.Y(_0017_),
    .A(net402),
    .B(_1255_));
 sg13g2_and2_1 _1551_ (.A(net257),
    .B(net402),
    .X(_1257_));
 sg13g2_nand2b_1 _1552_ (.Y(_1258_),
    .B(_1257_),
    .A_N(_1255_));
 sg13g2_xnor2_1 _1553_ (.Y(_0018_),
    .A(net257),
    .B(_1256_));
 sg13g2_nor2_1 _1554_ (.A(_1202_),
    .B(_1258_),
    .Y(_1259_));
 sg13g2_xnor2_1 _1555_ (.Y(_0019_),
    .A(net555),
    .B(_1258_));
 sg13g2_nand2_1 _1556_ (.Y(_1260_),
    .A(net314),
    .B(net555));
 sg13g2_nor2_1 _1557_ (.A(_1258_),
    .B(_1260_),
    .Y(_1261_));
 sg13g2_xor2_1 _1558_ (.B(_1259_),
    .A(net314),
    .X(_0020_));
 sg13g2_xnor2_1 _1559_ (.Y(_0021_),
    .A(_1201_),
    .B(_1261_));
 sg13g2_nand2_1 _1560_ (.Y(_1262_),
    .A(net305),
    .B(\adsr_pre_hi[7] ));
 sg13g2_nor3_1 _1561_ (.A(_1258_),
    .B(_1260_),
    .C(_1262_),
    .Y(_1263_));
 sg13g2_a21oi_1 _1562_ (.A1(\adsr_pre_hi[7] ),
    .A2(_1261_),
    .Y(_1264_),
    .B1(net305));
 sg13g2_nor2_1 _1563_ (.A(_1263_),
    .B(net306),
    .Y(_0022_));
 sg13g2_xnor2_1 _1564_ (.Y(_0023_),
    .A(_1203_),
    .B(_1263_));
 sg13g2_and3_1 _1565_ (.X(_1265_),
    .A(net278),
    .B(net697),
    .C(_1263_));
 sg13g2_a21oi_1 _1566_ (.A1(\adsr_pre_hi[9] ),
    .A2(_1263_),
    .Y(_1266_),
    .B1(net278));
 sg13g2_nor2_1 _1567_ (.A(_1265_),
    .B(net279),
    .Y(_0024_));
 sg13g2_xor2_1 _1568_ (.B(_1265_),
    .A(net360),
    .X(_0013_));
 sg13g2_nand3_1 _1569_ (.B(net360),
    .C(_1265_),
    .A(net722),
    .Y(_1267_));
 sg13g2_a21o_1 _1570_ (.A2(_1265_),
    .A1(net360),
    .B1(net722),
    .X(_1268_));
 sg13g2_and2_1 _1571_ (.A(_1267_),
    .B(net723),
    .X(_0014_));
 sg13g2_nand4_1 _1572_ (.B(\adsr_pre_hi[11] ),
    .C(\adsr_pre_hi[13] ),
    .A(\adsr_pre_hi[12] ),
    .Y(_1269_),
    .D(_1265_));
 sg13g2_xnor2_1 _1573_ (.Y(_0015_),
    .A(net259),
    .B(_1267_));
 sg13g2_nand2b_1 _1574_ (.Y(_1270_),
    .B(net729),
    .A_N(net699));
 sg13g2_o21ai_1 _1575_ (.B1(_1270_),
    .Y(_0000_),
    .A1(net699),
    .A2(net132));
 sg13g2_nand2b_1 _1576_ (.Y(_1271_),
    .B(net699),
    .A_N(net729));
 sg13g2_nand2_1 _1577_ (.Y(_0001_),
    .A(_1270_),
    .B(_1271_));
 sg13g2_and2_1 _1578_ (.A(\slot[1] ),
    .B(\slot[0] ),
    .X(_1272_));
 sg13g2_and2_1 _1579_ (.A(_1220_),
    .B(net119),
    .X(_1273_));
 sg13g2_a21o_1 _1580_ (.A2(_0001_),
    .A1(net132),
    .B1(net114),
    .X(_0002_));
 sg13g2_nand4_1 _1581_ (.B(net714),
    .C(net628),
    .A(net721),
    .Y(_1274_),
    .D(net695));
 sg13g2_nand2_1 _1582_ (.Y(_1275_),
    .A(net719),
    .B(net364));
 sg13g2_nor4_1 _1583_ (.A(net668),
    .B(_1226_),
    .C(_1274_),
    .D(_1275_),
    .Y(_1276_));
 sg13g2_nor2_1 _1584_ (.A(net668),
    .B(_1276_),
    .Y(_0004_));
 sg13g2_xnor2_1 _1585_ (.Y(_1277_),
    .A(net668),
    .B(net719));
 sg13g2_nor2_1 _1586_ (.A(_1276_),
    .B(_1277_),
    .Y(_0005_));
 sg13g2_and3_1 _1587_ (.X(_1278_),
    .A(net668),
    .B(net719),
    .C(net364));
 sg13g2_a21oi_1 _1588_ (.A1(\u_pwm.count[0] ),
    .A2(\u_pwm.count[1] ),
    .Y(_1279_),
    .B1(net364));
 sg13g2_nor3_1 _1589_ (.A(_1276_),
    .B(_1278_),
    .C(net365),
    .Y(_0006_));
 sg13g2_nor2_1 _1590_ (.A(net692),
    .B(_1278_),
    .Y(_1280_));
 sg13g2_and2_1 _1591_ (.A(net692),
    .B(_1278_),
    .X(_1281_));
 sg13g2_nor3_1 _1592_ (.A(_1276_),
    .B(net693),
    .C(_1281_),
    .Y(_0007_));
 sg13g2_nor2_1 _1593_ (.A(net714),
    .B(_1281_),
    .Y(_1282_));
 sg13g2_and2_1 _1594_ (.A(net714),
    .B(_1281_),
    .X(_1283_));
 sg13g2_nor3_1 _1595_ (.A(_1276_),
    .B(net715),
    .C(_1283_),
    .Y(_0008_));
 sg13g2_xnor2_1 _1596_ (.Y(_1284_),
    .A(net721),
    .B(_1283_));
 sg13g2_nor2_1 _1597_ (.A(_1276_),
    .B(_1284_),
    .Y(_0009_));
 sg13g2_nand3_1 _1598_ (.B(net628),
    .C(_1283_),
    .A(\u_pwm.count[5] ),
    .Y(_1285_));
 sg13g2_inv_1 _1599_ (.Y(_1286_),
    .A(_1285_));
 sg13g2_a21oi_1 _1600_ (.A1(\u_pwm.count[5] ),
    .A2(_1283_),
    .Y(_1287_),
    .B1(net628));
 sg13g2_nor3_1 _1601_ (.A(_1276_),
    .B(_1286_),
    .C(net629),
    .Y(_0010_));
 sg13g2_nand3b_1 _1602_ (.B(_1285_),
    .C(net695),
    .Y(_1288_),
    .A_N(_1276_));
 sg13g2_o21ai_1 _1603_ (.B1(_1288_),
    .Y(_0011_),
    .A1(net695),
    .A2(_1285_));
 sg13g2_nand2b_1 _1604_ (.Y(_1289_),
    .B(\mix_out[1] ),
    .A_N(\u_pwm.count[1] ));
 sg13g2_nand2b_1 _1605_ (.Y(_1290_),
    .B(\mix_out[0] ),
    .A_N(\u_pwm.count[0] ));
 sg13g2_nand2b_1 _1606_ (.Y(_1291_),
    .B(\u_pwm.count[1] ),
    .A_N(\mix_out[1] ));
 sg13g2_o21ai_1 _1607_ (.B1(_1291_),
    .Y(_1292_),
    .A1(_1227_),
    .A2(\mix_out[2] ));
 sg13g2_a21oi_1 _1608_ (.A1(_1289_),
    .A2(_1290_),
    .Y(_1293_),
    .B1(_1292_));
 sg13g2_a221oi_1 _1609_ (.B2(_1227_),
    .C1(_1293_),
    .B1(net392),
    .A1(_1226_),
    .Y(_1294_),
    .A2(net519));
 sg13g2_a221oi_1 _1610_ (.B2(net692),
    .C1(_1294_),
    .B1(_1254_),
    .A1(net714),
    .Y(_1295_),
    .A2(_1253_));
 sg13g2_nand2b_1 _1611_ (.Y(_1296_),
    .B(net548),
    .A_N(\u_pwm.count[5] ));
 sg13g2_o21ai_1 _1612_ (.B1(_1296_),
    .Y(_1297_),
    .A1(net714),
    .A2(_1253_));
 sg13g2_a22oi_1 _1613_ (.Y(_1298_),
    .B1(_1252_),
    .B2(net721),
    .A2(_1251_),
    .A1(net628));
 sg13g2_o21ai_1 _1614_ (.B1(_1298_),
    .Y(_1299_),
    .A1(_1295_),
    .A2(_1297_));
 sg13g2_a22oi_1 _1615_ (.Y(_1300_),
    .B1(net538),
    .B2(_1228_),
    .A2(net730),
    .A1(_1229_));
 sg13g2_a22oi_1 _1616_ (.Y(_0003_),
    .B1(_1299_),
    .B2(_1300_),
    .A2(_1250_),
    .A1(net695));
 sg13g2_nand2_1 _1617_ (.Y(_1301_),
    .A(net589),
    .B(\p_freq[7] ));
 sg13g2_nand2_1 _1618_ (.Y(_1302_),
    .A(\p_acc[6] ),
    .B(\p_freq[6] ));
 sg13g2_inv_1 _1619_ (.Y(_1303_),
    .A(_1302_));
 sg13g2_nand2_1 _1620_ (.Y(_1304_),
    .A(_1169_),
    .B(_1170_));
 sg13g2_nand2_1 _1621_ (.Y(_1305_),
    .A(_1302_),
    .B(_1304_));
 sg13g2_nand2_1 _1622_ (.Y(_1306_),
    .A(\p_acc[5] ),
    .B(\p_freq[5] ));
 sg13g2_xnor2_1 _1623_ (.Y(_1307_),
    .A(\p_acc[5] ),
    .B(\p_freq[5] ));
 sg13g2_nand2_1 _1624_ (.Y(_1308_),
    .A(net451),
    .B(\p_freq[4] ));
 sg13g2_inv_1 _1625_ (.Y(_1309_),
    .A(_1308_));
 sg13g2_nand2_1 _1626_ (.Y(_1310_),
    .A(_1173_),
    .B(_1174_));
 sg13g2_nand2_1 _1627_ (.Y(_1311_),
    .A(_1308_),
    .B(_1310_));
 sg13g2_nand2_1 _1628_ (.Y(_1312_),
    .A(\p_acc[3] ),
    .B(\p_freq[3] ));
 sg13g2_nand2_1 _1629_ (.Y(_1313_),
    .A(\p_acc[2] ),
    .B(\p_freq[2] ));
 sg13g2_inv_1 _1630_ (.Y(_1314_),
    .A(_1313_));
 sg13g2_nand2_1 _1631_ (.Y(_1315_),
    .A(_1177_),
    .B(_1178_));
 sg13g2_nand2_1 _1632_ (.Y(_1316_),
    .A(_1313_),
    .B(_1315_));
 sg13g2_nand2_1 _1633_ (.Y(_1317_),
    .A(\p_acc[1] ),
    .B(\p_freq[1] ));
 sg13g2_xnor2_1 _1634_ (.Y(_1318_),
    .A(\p_acc[1] ),
    .B(\p_freq[1] ));
 sg13g2_nand2_1 _1635_ (.Y(_1319_),
    .A(\p_acc[0] ),
    .B(net476));
 sg13g2_o21ai_1 _1636_ (.B1(_1317_),
    .Y(_1320_),
    .A1(_1318_),
    .A2(_1319_));
 sg13g2_a21oi_1 _1637_ (.A1(_1315_),
    .A2(_1320_),
    .Y(_1321_),
    .B1(_1314_));
 sg13g2_xnor2_1 _1638_ (.Y(_1322_),
    .A(\p_acc[3] ),
    .B(\p_freq[3] ));
 sg13g2_or2_1 _1639_ (.X(_1323_),
    .B(_1322_),
    .A(_1321_));
 sg13g2_o21ai_1 _1640_ (.B1(_1312_),
    .Y(_1324_),
    .A1(_1321_),
    .A2(_1322_));
 sg13g2_nand2b_1 _1641_ (.Y(_1325_),
    .B(_1324_),
    .A_N(_1311_));
 sg13g2_a21oi_1 _1642_ (.A1(_1310_),
    .A2(_1324_),
    .Y(_1326_),
    .B1(_1309_));
 sg13g2_or2_1 _1643_ (.X(_1327_),
    .B(_1326_),
    .A(_1307_));
 sg13g2_o21ai_1 _1644_ (.B1(_1306_),
    .Y(_1328_),
    .A1(_1307_),
    .A2(_1326_));
 sg13g2_nand2b_1 _1645_ (.Y(_1329_),
    .B(_1328_),
    .A_N(_1305_));
 sg13g2_a21oi_1 _1646_ (.A1(_1304_),
    .A2(_1328_),
    .Y(_1330_),
    .B1(_1303_));
 sg13g2_xnor2_1 _1647_ (.Y(_1331_),
    .A(\p_acc[7] ),
    .B(\p_freq[7] ));
 sg13g2_o21ai_1 _1648_ (.B1(_1301_),
    .Y(_1332_),
    .A1(_1330_),
    .A2(_1331_));
 sg13g2_nand2_1 _1649_ (.Y(_1333_),
    .A(\p_acc[8] ),
    .B(_1332_));
 sg13g2_and4_1 _1650_ (.A(net641),
    .B(\p_acc[9] ),
    .C(\p_acc[8] ),
    .D(_1332_),
    .X(_1334_));
 sg13g2_nand4_1 _1651_ (.B(\p_acc[9] ),
    .C(\p_acc[8] ),
    .A(\p_acc[10] ),
    .Y(_1335_),
    .D(_1332_));
 sg13g2_nand3_1 _1652_ (.B(\p_acc[11] ),
    .C(_1334_),
    .A(\p_acc[12] ),
    .Y(_1336_));
 sg13g2_nor4_1 _1653_ (.A(_1161_),
    .B(_1162_),
    .C(_1163_),
    .D(_1335_),
    .Y(_1337_));
 sg13g2_a21o_1 _1654_ (.A2(_1337_),
    .A1(net618),
    .B1(net577),
    .X(_1338_));
 sg13g2_nor2_1 _1655_ (.A(\slot[1] ),
    .B(net699),
    .Y(_1339_));
 sg13g2_or2_1 _1656_ (.X(_1340_),
    .B(net699),
    .A(\slot[1] ));
 sg13g2_nand2b_1 _1657_ (.Y(_1341_),
    .B(\slot[1] ),
    .A_N(\acc[1][15] ));
 sg13g2_o21ai_1 _1658_ (.B1(_1341_),
    .Y(_1342_),
    .A1(\acc[0][15] ),
    .A2(_1271_));
 sg13g2_a21oi_1 _1659_ (.A1(_1185_),
    .A2(_1339_),
    .Y(_1343_),
    .B1(_1342_));
 sg13g2_nor2_1 _1660_ (.A(p_prev_msb_d),
    .B(_1187_),
    .Y(_1344_));
 sg13g2_a21oi_1 _1661_ (.A1(_1343_),
    .A2(_1344_),
    .Y(_1345_),
    .B1(net416));
 sg13g2_nand3_1 _1662_ (.B(net577),
    .C(_1337_),
    .A(net618),
    .Y(_1346_));
 sg13g2_nand3_1 _1663_ (.B(net34),
    .C(_1346_),
    .A(_1338_),
    .Y(_1347_));
 sg13g2_nand2_1 _1664_ (.Y(_1348_),
    .A(\p_pw[7] ),
    .B(_1347_));
 sg13g2_xnor2_1 _1665_ (.Y(_1349_),
    .A(\p_acc[9] ),
    .B(_1333_));
 sg13g2_nand2_1 _1666_ (.Y(_1350_),
    .A(net35),
    .B(_1349_));
 sg13g2_nand3_1 _1667_ (.B(net35),
    .C(_1349_),
    .A(_1239_),
    .Y(_1351_));
 sg13g2_o21ai_1 _1668_ (.B1(net35),
    .Y(_1352_),
    .A1(\p_acc[8] ),
    .A2(_1332_));
 sg13g2_nand2b_1 _1669_ (.Y(_1353_),
    .B(_1333_),
    .A_N(_1352_));
 sg13g2_and2_1 _1670_ (.A(\p_pw[0] ),
    .B(_1353_),
    .X(_1354_));
 sg13g2_a21oi_1 _1671_ (.A1(net35),
    .A2(_1349_),
    .Y(_1355_),
    .B1(_1239_));
 sg13g2_o21ai_1 _1672_ (.B1(_1164_),
    .Y(_1356_),
    .A1(_1165_),
    .A2(_1333_));
 sg13g2_nand3_1 _1673_ (.B(net35),
    .C(_1356_),
    .A(_1335_),
    .Y(_1357_));
 sg13g2_a221oi_1 _1674_ (.B2(\p_pw[2] ),
    .C1(_1355_),
    .B1(_1357_),
    .A1(_1351_),
    .Y(_1358_),
    .A2(_1354_));
 sg13g2_xnor2_1 _1675_ (.Y(_1359_),
    .A(_1163_),
    .B(net642));
 sg13g2_nand2_1 _1676_ (.Y(_1360_),
    .A(net34),
    .B(net643));
 sg13g2_nand3_1 _1677_ (.B(net34),
    .C(_1359_),
    .A(_1237_),
    .Y(_1361_));
 sg13g2_o21ai_1 _1678_ (.B1(_1361_),
    .Y(_1362_),
    .A1(\p_pw[2] ),
    .A2(_1357_));
 sg13g2_o21ai_1 _1679_ (.B1(_1162_),
    .Y(_1363_),
    .A1(_1163_),
    .A2(_1335_));
 sg13g2_nand3_1 _1680_ (.B(net34),
    .C(_1363_),
    .A(_1336_),
    .Y(_1364_));
 sg13g2_a22oi_1 _1681_ (.Y(_1365_),
    .B1(_1364_),
    .B2(\p_pw[4] ),
    .A2(_1360_),
    .A1(\p_pw[3] ));
 sg13g2_o21ai_1 _1682_ (.B1(_1365_),
    .Y(_1366_),
    .A1(_1358_),
    .A2(_1362_));
 sg13g2_nor2_1 _1683_ (.A(\p_pw[4] ),
    .B(_1364_),
    .Y(_1367_));
 sg13g2_xnor2_1 _1684_ (.Y(_1368_),
    .A(\p_acc[13] ),
    .B(_1336_));
 sg13g2_and2_1 _1685_ (.A(net34),
    .B(_1368_),
    .X(_1369_));
 sg13g2_nand2_1 _1686_ (.Y(_1370_),
    .A(net34),
    .B(_1368_));
 sg13g2_a21oi_1 _1687_ (.A1(_1235_),
    .A2(_1369_),
    .Y(_1371_),
    .B1(_1367_));
 sg13g2_xnor2_1 _1688_ (.Y(_1372_),
    .A(_1183_),
    .B(_1337_));
 sg13g2_nand2_1 _1689_ (.Y(_1373_),
    .A(net34),
    .B(_1372_));
 sg13g2_a21oi_1 _1690_ (.A1(net34),
    .A2(_1372_),
    .Y(_1374_),
    .B1(_1234_));
 sg13g2_a221oi_1 _1691_ (.B2(_1366_),
    .C1(_1374_),
    .B1(_1371_),
    .A1(\p_pw[5] ),
    .Y(_1375_),
    .A2(_1370_));
 sg13g2_nand3_1 _1692_ (.B(net35),
    .C(_1372_),
    .A(_1234_),
    .Y(_1376_));
 sg13g2_o21ai_1 _1693_ (.B1(_1376_),
    .Y(_1377_),
    .A1(\p_pw[7] ),
    .A2(_1347_));
 sg13g2_o21ai_1 _1694_ (.B1(_1348_),
    .Y(_1378_),
    .A1(_1375_),
    .A2(_1377_));
 sg13g2_nand2_1 _1695_ (.Y(_1379_),
    .A(net144),
    .B(net31));
 sg13g2_nor4_1 _1696_ (.A(\p_waveform[4] ),
    .B(net146),
    .C(net145),
    .D(net142),
    .Y(_1380_));
 sg13g2_or2_1 _1697_ (.X(_1381_),
    .B(_1380_),
    .A(\p_waveform[4] ));
 sg13g2_a221oi_1 _1698_ (.B2(net146),
    .C1(_1381_),
    .B1(_1353_),
    .A1(_0032_),
    .Y(_1382_),
    .A2(net142));
 sg13g2_inv_1 _1699_ (.Y(_1383_),
    .A(_1382_));
 sg13g2_a21oi_1 _1700_ (.A1(net143),
    .A2(net30),
    .Y(_1384_),
    .B1(_1383_));
 sg13g2_nor2_1 _1701_ (.A(_1189_),
    .B(net342),
    .Y(_1385_));
 sg13g2_nor2_1 _1702_ (.A(net139),
    .B(net140),
    .Y(_1386_));
 sg13g2_nor3_1 _1703_ (.A(net139),
    .B(net140),
    .C(net141),
    .Y(_1387_));
 sg13g2_and2_1 _1704_ (.A(_1198_),
    .B(_1387_),
    .X(_1388_));
 sg13g2_nand2_1 _1705_ (.Y(_1389_),
    .A(_1196_),
    .B(_1388_));
 sg13g2_or2_1 _1706_ (.X(_1390_),
    .B(net137),
    .A(net136));
 sg13g2_nor2_1 _1707_ (.A(net136),
    .B(net138),
    .Y(_1391_));
 sg13g2_nor3_1 _1708_ (.A(net136),
    .B(net137),
    .C(net138),
    .Y(_1392_));
 sg13g2_nor2_1 _1709_ (.A(net138),
    .B(_1389_),
    .Y(_1393_));
 sg13g2_nor3_1 _1710_ (.A(net137),
    .B(net138),
    .C(_1389_),
    .Y(_1394_));
 sg13g2_nand2_1 _1711_ (.Y(_1395_),
    .A(_1188_),
    .B(_1394_));
 sg13g2_nor2b_1 _1712_ (.A(_1385_),
    .B_N(_1395_),
    .Y(_1396_));
 sg13g2_nand2_1 _1713_ (.Y(_1397_),
    .A(\p_env[4] ),
    .B(\p_env[3] ));
 sg13g2_o21ai_1 _1714_ (.B1(_1392_),
    .Y(_1398_),
    .A1(_1386_),
    .A2(_1397_));
 sg13g2_nand3_1 _1715_ (.B(\p_env[3] ),
    .C(net140),
    .A(net139),
    .Y(_1399_));
 sg13g2_nor4_1 _1716_ (.A(net136),
    .B(\p_env[6] ),
    .C(\p_env[5] ),
    .D(\p_env[4] ),
    .Y(_1400_));
 sg13g2_a21oi_1 _1717_ (.A1(_1399_),
    .A2(_1400_),
    .Y(_1401_),
    .B1(\p_sustain[4] ));
 sg13g2_nor2_1 _1718_ (.A(_1398_),
    .B(_1401_),
    .Y(_1402_));
 sg13g2_o21ai_1 _1719_ (.B1(_1212_),
    .Y(_1403_),
    .A1(_1398_),
    .A2(_1401_));
 sg13g2_o21ai_1 _1720_ (.B1(net139),
    .Y(_1404_),
    .A1(net140),
    .A2(net141));
 sg13g2_inv_1 _1721_ (.Y(_1405_),
    .A(_1404_));
 sg13g2_o21ai_1 _1722_ (.B1(_1391_),
    .Y(_1406_),
    .A1(_1397_),
    .A2(_1404_));
 sg13g2_and2_1 _1723_ (.A(_1390_),
    .B(_1406_),
    .X(_1407_));
 sg13g2_nand2_1 _1724_ (.Y(_1408_),
    .A(_1390_),
    .B(_1406_));
 sg13g2_and2_1 _1725_ (.A(\p_env[5] ),
    .B(\p_env[4] ),
    .X(_1409_));
 sg13g2_a21o_1 _1726_ (.A2(net140),
    .A1(net139),
    .B1(\p_env[3] ),
    .X(_1410_));
 sg13g2_a21oi_1 _1727_ (.A1(_1409_),
    .A2(_1410_),
    .Y(_1411_),
    .B1(_1390_));
 sg13g2_or2_1 _1728_ (.X(_1412_),
    .B(_1411_),
    .A(\p_sustain[4] ));
 sg13g2_nand2_1 _1729_ (.Y(_1413_),
    .A(_1403_),
    .B(_1412_));
 sg13g2_nand4_1 _1730_ (.B(_1403_),
    .C(_1408_),
    .A(\p_sustain[6] ),
    .Y(_1414_),
    .D(_1412_));
 sg13g2_nor2_1 _1731_ (.A(\p_sustain[7] ),
    .B(net130),
    .Y(_1415_));
 sg13g2_nor2_1 _1732_ (.A(_1208_),
    .B(\p_ast[0] ),
    .Y(_1416_));
 sg13g2_a21oi_1 _1733_ (.A1(_1399_),
    .A2(_1400_),
    .Y(_1417_),
    .B1(\p_attack[4] ));
 sg13g2_a21o_1 _1734_ (.A2(_1400_),
    .A1(_1399_),
    .B1(\p_attack[4] ),
    .X(_1418_));
 sg13g2_nor2_1 _1735_ (.A(_1398_),
    .B(_1417_),
    .Y(_1419_));
 sg13g2_nor2_1 _1736_ (.A(\p_attack[5] ),
    .B(_1419_),
    .Y(_1420_));
 sg13g2_a21o_1 _1737_ (.A2(\p_attack[5] ),
    .A1(\p_attack[4] ),
    .B1(_1411_),
    .X(_1421_));
 sg13g2_nand3_1 _1738_ (.B(_1408_),
    .C(_1421_),
    .A(\p_attack[6] ),
    .Y(_1422_));
 sg13g2_o21ai_1 _1739_ (.B1(_1206_),
    .Y(_1423_),
    .A1(_1420_),
    .A2(_1422_));
 sg13g2_nor2_1 _1740_ (.A(\p_ast[1] ),
    .B(_1209_),
    .Y(_1424_));
 sg13g2_nand2_1 _1741_ (.Y(_1425_),
    .A(_1208_),
    .B(\p_ast[0] ));
 sg13g2_a221oi_1 _1742_ (.B2(\p_attack[3] ),
    .C1(net135),
    .B1(_1424_),
    .A1(net112),
    .Y(_1426_),
    .A2(_1423_));
 sg13g2_a21oi_1 _1743_ (.A1(_1414_),
    .A2(_1415_),
    .Y(_1427_),
    .B1(_1426_));
 sg13g2_nor2b_1 _1744_ (.A(_1269_),
    .B_N(_1427_),
    .Y(_1428_));
 sg13g2_and2_1 _1745_ (.A(\p_attack[7] ),
    .B(\p_attack[6] ),
    .X(_1429_));
 sg13g2_nand2_1 _1746_ (.Y(_1430_),
    .A(\p_attack[7] ),
    .B(\p_attack[6] ));
 sg13g2_a21oi_1 _1747_ (.A1(\p_attack[5] ),
    .A2(_1429_),
    .Y(_1431_),
    .B1(\p_attack[4] ));
 sg13g2_nand2_1 _1748_ (.Y(_1432_),
    .A(_1398_),
    .B(_1431_));
 sg13g2_and3_1 _1749_ (.X(_1433_),
    .A(\p_attack[4] ),
    .B(_1399_),
    .C(_1400_));
 sg13g2_nand3_1 _1750_ (.B(_1399_),
    .C(_1400_),
    .A(\p_attack[4] ),
    .Y(_1434_));
 sg13g2_or4_1 _1751_ (.A(_1398_),
    .B(_1417_),
    .C(_1429_),
    .D(_1433_),
    .X(_1435_));
 sg13g2_a21o_1 _1752_ (.A2(_1429_),
    .A1(\p_attack[5] ),
    .B1(_1411_),
    .X(_1436_));
 sg13g2_nand3_1 _1753_ (.B(_1435_),
    .C(_1436_),
    .A(_1432_),
    .Y(_1437_));
 sg13g2_a21o_1 _1754_ (.A2(_1435_),
    .A1(_1432_),
    .B1(_1411_),
    .X(_1438_));
 sg13g2_nand3_1 _1755_ (.B(_1437_),
    .C(_1438_),
    .A(_1408_),
    .Y(_1439_));
 sg13g2_nor2_1 _1756_ (.A(\p_attack[4] ),
    .B(_1408_),
    .Y(_1440_));
 sg13g2_nor2b_1 _1757_ (.A(_1440_),
    .B_N(net112),
    .Y(_1441_));
 sg13g2_a221oi_1 _1758_ (.B2(_1441_),
    .C1(net135),
    .B1(_1439_),
    .A1(\p_attack[0] ),
    .Y(_1442_),
    .A2(_1424_));
 sg13g2_nor2_1 _1759_ (.A(_1213_),
    .B(_1214_),
    .Y(_1443_));
 sg13g2_nand3_1 _1760_ (.B(_1399_),
    .C(_1400_),
    .A(\p_sustain[4] ),
    .Y(_1444_));
 sg13g2_nor2b_1 _1761_ (.A(_1443_),
    .B_N(_1444_),
    .Y(_1445_));
 sg13g2_a21oi_1 _1762_ (.A1(\p_sustain[5] ),
    .A2(_1443_),
    .Y(_1446_),
    .B1(\p_sustain[4] ));
 sg13g2_a22oi_1 _1763_ (.Y(_1447_),
    .B1(_1446_),
    .B2(_1398_),
    .A2(_1445_),
    .A1(_1402_));
 sg13g2_nand2b_1 _1764_ (.Y(_1448_),
    .B(_1411_),
    .A_N(_1447_));
 sg13g2_a21oi_1 _1765_ (.A1(\p_sustain[5] ),
    .A2(_1443_),
    .Y(_1449_),
    .B1(_1411_));
 sg13g2_a21oi_1 _1766_ (.A1(_1447_),
    .A2(_1449_),
    .Y(_1450_),
    .B1(_1407_));
 sg13g2_a221oi_1 _1767_ (.B2(_1450_),
    .C1(net130),
    .B1(_1448_),
    .A1(\p_sustain[4] ),
    .Y(_0349_),
    .A2(_1407_));
 sg13g2_nor2_1 _1768_ (.A(_1442_),
    .B(_0349_),
    .Y(_0350_));
 sg13g2_nand4_1 _1769_ (.B(_1418_),
    .C(_1430_),
    .A(_1398_),
    .Y(_0351_),
    .D(_1434_));
 sg13g2_xnor2_1 _1770_ (.Y(_0352_),
    .A(_1205_),
    .B(_1417_));
 sg13g2_nand3b_1 _1771_ (.B(_0351_),
    .C(_1430_),
    .Y(_0353_),
    .A_N(_0352_));
 sg13g2_nand2b_1 _1772_ (.Y(_0354_),
    .B(_0352_),
    .A_N(_0351_));
 sg13g2_a21oi_1 _1773_ (.A1(_0353_),
    .A2(_0354_),
    .Y(_0355_),
    .B1(_1438_));
 sg13g2_and3_1 _1774_ (.X(_0356_),
    .A(_1438_),
    .B(_0353_),
    .C(_0354_));
 sg13g2_nor3_1 _1775_ (.A(_1407_),
    .B(_0355_),
    .C(_0356_),
    .Y(_0357_));
 sg13g2_o21ai_1 _1776_ (.B1(net112),
    .Y(_0358_),
    .A1(\p_attack[5] ),
    .A2(_1408_));
 sg13g2_nand2_1 _1777_ (.Y(_0359_),
    .A(\p_attack[1] ),
    .B(_1424_));
 sg13g2_o21ai_1 _1778_ (.B1(_0359_),
    .Y(_0360_),
    .A1(_0357_),
    .A2(_0358_));
 sg13g2_nor2_1 _1779_ (.A(\p_sustain[5] ),
    .B(_1443_),
    .Y(_0361_));
 sg13g2_nand2b_1 _1780_ (.Y(_0362_),
    .B(_1446_),
    .A_N(_1411_));
 sg13g2_xnor2_1 _1781_ (.Y(_0363_),
    .A(_0361_),
    .B(_0362_));
 sg13g2_nor2b_1 _1782_ (.A(_1402_),
    .B_N(_1445_),
    .Y(_0364_));
 sg13g2_a21oi_1 _1783_ (.A1(_0363_),
    .A2(_0364_),
    .Y(_0365_),
    .B1(_1407_));
 sg13g2_o21ai_1 _1784_ (.B1(_0365_),
    .Y(_0366_),
    .A1(_0363_),
    .A2(_0364_));
 sg13g2_a21oi_1 _1785_ (.A1(_1212_),
    .A2(_1407_),
    .Y(_0367_),
    .B1(net130));
 sg13g2_a22oi_1 _1786_ (.Y(_0368_),
    .B1(_0366_),
    .B2(_0367_),
    .A2(_0360_),
    .A1(net130));
 sg13g2_o21ai_1 _1787_ (.B1(\adsr_pre_hi[3] ),
    .Y(_0369_),
    .A1(\adsr_pre_hi[5] ),
    .A2(_0368_));
 sg13g2_a21oi_1 _1788_ (.A1(_1203_),
    .A2(_0350_),
    .Y(_0370_),
    .B1(_1262_));
 sg13g2_nand3_1 _1789_ (.B(\adsr_pre_hi[5] ),
    .C(_1257_),
    .A(\adsr_pre_hi[6] ),
    .Y(_0371_));
 sg13g2_a21oi_1 _1790_ (.A1(_1201_),
    .A2(_0350_),
    .Y(_0372_),
    .B1(_0371_));
 sg13g2_o21ai_1 _1791_ (.B1(_0372_),
    .Y(_0373_),
    .A1(_0368_),
    .A2(_0370_));
 sg13g2_o21ai_1 _1792_ (.B1(_1214_),
    .Y(_0374_),
    .A1(_1407_),
    .A2(_1413_));
 sg13g2_nand2_1 _1793_ (.Y(_0375_),
    .A(_1414_),
    .B(_0374_));
 sg13g2_nor2_1 _1794_ (.A(_1215_),
    .B(_1443_),
    .Y(_0376_));
 sg13g2_a21oi_1 _1795_ (.A1(_1411_),
    .A2(_1420_),
    .Y(_0377_),
    .B1(_1407_));
 sg13g2_xnor2_1 _1796_ (.Y(_0378_),
    .A(\p_attack[6] ),
    .B(_1421_));
 sg13g2_nand3_1 _1797_ (.B(_0377_),
    .C(_0378_),
    .A(_1430_),
    .Y(_0379_));
 sg13g2_o21ai_1 _1798_ (.B1(_1416_),
    .Y(_0380_),
    .A1(\p_attack[6] ),
    .A2(_0377_));
 sg13g2_nand2b_1 _1799_ (.Y(_0381_),
    .B(_0379_),
    .A_N(_0380_));
 sg13g2_a21oi_1 _1800_ (.A1(\p_attack[2] ),
    .A2(_1424_),
    .Y(_0382_),
    .B1(net135));
 sg13g2_a22oi_1 _1801_ (.Y(_0383_),
    .B1(_0381_),
    .B2(_0382_),
    .A2(_0376_),
    .A1(_0375_));
 sg13g2_nor2_1 _1802_ (.A(_1255_),
    .B(_1427_),
    .Y(_0384_));
 sg13g2_o21ai_1 _1803_ (.B1(_0384_),
    .Y(_0385_),
    .A1(_1257_),
    .A2(_0368_));
 sg13g2_a221oi_1 _1804_ (.B2(_0383_),
    .C1(_0385_),
    .B1(_0373_),
    .A1(_0350_),
    .Y(_0386_),
    .A2(_0369_));
 sg13g2_nor2_1 _1805_ (.A(_1428_),
    .B(_0386_),
    .Y(_0387_));
 sg13g2_nor2b_1 _1806_ (.A(net32),
    .B_N(_1396_),
    .Y(_0388_));
 sg13g2_xnor2_1 _1807_ (.Y(_0389_),
    .A(_1194_),
    .B(_1389_));
 sg13g2_a21oi_1 _1808_ (.A1(_0388_),
    .A2(_0389_),
    .Y(_0390_),
    .B1(net130));
 sg13g2_o21ai_1 _1809_ (.B1(_0390_),
    .Y(_0391_),
    .A1(net138),
    .A2(_0388_));
 sg13g2_nor2_1 _1810_ (.A(\p_ast[1] ),
    .B(\p_ast[0] ),
    .Y(_0392_));
 sg13g2_nor2_1 _1811_ (.A(net134),
    .B(_0392_),
    .Y(_0393_));
 sg13g2_or2_1 _1812_ (.X(_0394_),
    .B(_0392_),
    .A(net134));
 sg13g2_nand3_1 _1813_ (.B(net141),
    .C(_1409_),
    .A(\p_env[6] ),
    .Y(_0395_));
 sg13g2_nor3_1 _1814_ (.A(_1188_),
    .B(_1399_),
    .C(_0395_),
    .Y(_0396_));
 sg13g2_nand2b_1 _1815_ (.Y(_0397_),
    .B(net147),
    .A_N(_0396_));
 sg13g2_nor3_1 _1816_ (.A(_1197_),
    .B(_1199_),
    .C(_1200_),
    .Y(_0398_));
 sg13g2_o21ai_1 _1817_ (.B1(_0398_),
    .Y(_0399_),
    .A1(_1428_),
    .A2(_0386_));
 sg13g2_nor3_1 _1818_ (.A(_1397_),
    .B(_0397_),
    .C(_0399_),
    .Y(_0400_));
 sg13g2_xnor2_1 _1819_ (.Y(_0401_),
    .A(_1194_),
    .B(_0400_));
 sg13g2_nor2_1 _1820_ (.A(net147),
    .B(_1208_),
    .Y(_0402_));
 sg13g2_a22oi_1 _1821_ (.Y(_0403_),
    .B1(_1195_),
    .B2(\p_env[4] ),
    .A2(\p_env[5] ),
    .A1(_1193_));
 sg13g2_a221oi_1 _1822_ (.B2(_1194_),
    .C1(_0403_),
    .B1(\p_sustain[1] ),
    .A1(\p_sustain[2] ),
    .Y(_0404_),
    .A2(_1192_));
 sg13g2_a221oi_1 _1823_ (.B2(\p_env[6] ),
    .C1(_0404_),
    .B1(_1191_),
    .A1(net136),
    .Y(_0405_),
    .A2(_1190_));
 sg13g2_a21oi_1 _1824_ (.A1(_1188_),
    .A2(\p_sustain[3] ),
    .Y(_0406_),
    .B1(_0405_));
 sg13g2_nor2b_1 _1825_ (.A(net33),
    .B_N(_0406_),
    .Y(_0407_));
 sg13g2_o21ai_1 _1826_ (.B1(_0406_),
    .Y(_0408_),
    .A1(_1428_),
    .A2(_0386_));
 sg13g2_nor3_1 _1827_ (.A(_1189_),
    .B(_1208_),
    .C(_0389_),
    .Y(_0409_));
 sg13g2_nor2_1 _1828_ (.A(_1208_),
    .B(_1209_),
    .Y(_0410_));
 sg13g2_nand2_1 _1829_ (.Y(_0411_),
    .A(net147),
    .B(_0410_));
 sg13g2_inv_1 _1830_ (.Y(_0412_),
    .A(_0411_));
 sg13g2_a22oi_1 _1831_ (.Y(_0413_),
    .B1(_0412_),
    .B2(net737),
    .A2(net112),
    .A1(net138));
 sg13g2_a22oi_1 _1832_ (.Y(_0414_),
    .B1(_0407_),
    .B2(_0409_),
    .A2(_0402_),
    .A1(net138));
 sg13g2_o21ai_1 _1833_ (.B1(_0414_),
    .Y(_0415_),
    .A1(_0407_),
    .A2(_0413_));
 sg13g2_a21oi_1 _1834_ (.A1(_1424_),
    .A2(_0401_),
    .Y(_0416_),
    .B1(_0415_));
 sg13g2_o21ai_1 _1835_ (.B1(_0391_),
    .Y(_0417_),
    .A1(_0394_),
    .A2(_0416_));
 sg13g2_and2_1 _1836_ (.A(net28),
    .B(net26),
    .X(_0418_));
 sg13g2_nand2_1 _1837_ (.Y(_0419_),
    .A(net28),
    .B(net26));
 sg13g2_nor3_1 _1838_ (.A(\p_env[2] ),
    .B(_1428_),
    .C(_0386_),
    .Y(_0420_));
 sg13g2_nor2_1 _1839_ (.A(_1425_),
    .B(_0396_),
    .Y(_0421_));
 sg13g2_nor2_1 _1840_ (.A(_1425_),
    .B(_0397_),
    .Y(_0422_));
 sg13g2_nand2_1 _1841_ (.Y(_0423_),
    .A(net147),
    .B(_0421_));
 sg13g2_a21oi_1 _1842_ (.A1(\p_env[1] ),
    .A2(net141),
    .Y(_0424_),
    .B1(\p_env[2] ));
 sg13g2_nor3_1 _1843_ (.A(_0420_),
    .B(_0423_),
    .C(_0424_),
    .Y(_0425_));
 sg13g2_nor3_1 _1844_ (.A(_1387_),
    .B(_1405_),
    .C(net32),
    .Y(_0426_));
 sg13g2_nor2_1 _1845_ (.A(_0406_),
    .B(_0411_),
    .Y(_0427_));
 sg13g2_or2_1 _1846_ (.X(_0428_),
    .B(_0402_),
    .A(_1424_));
 sg13g2_nor2b_1 _1847_ (.A(_0406_),
    .B_N(net112),
    .Y(_0429_));
 sg13g2_a21o_1 _1848_ (.A2(_0428_),
    .A1(_0397_),
    .B1(_0429_),
    .X(_0430_));
 sg13g2_a21oi_1 _1849_ (.A1(net139),
    .A2(_0430_),
    .Y(_0431_),
    .B1(_0427_));
 sg13g2_o21ai_1 _1850_ (.B1(_0431_),
    .Y(_0432_),
    .A1(_0411_),
    .A2(_0426_));
 sg13g2_nand3_1 _1851_ (.B(net112),
    .C(_0406_),
    .A(net147),
    .Y(_0433_));
 sg13g2_inv_1 _1852_ (.Y(_0434_),
    .A(_0433_));
 sg13g2_nor3_1 _1853_ (.A(_0420_),
    .B(_0426_),
    .C(_0433_),
    .Y(_0435_));
 sg13g2_a21o_1 _1854_ (.A2(_0425_),
    .A1(_0399_),
    .B1(_0435_),
    .X(_0436_));
 sg13g2_o21ai_1 _1855_ (.B1(_0393_),
    .Y(_0437_),
    .A1(_0432_),
    .A2(_0436_));
 sg13g2_nand2_1 _1856_ (.Y(_0438_),
    .A(net134),
    .B(_1396_));
 sg13g2_or3_1 _1857_ (.A(_0420_),
    .B(_0426_),
    .C(_0438_),
    .X(_0439_));
 sg13g2_nand3_1 _1858_ (.B(net134),
    .C(_1385_),
    .A(net139),
    .Y(_0440_));
 sg13g2_nand3_1 _1859_ (.B(_0439_),
    .C(_0440_),
    .A(_0437_),
    .Y(_0441_));
 sg13g2_nand2_1 _1860_ (.Y(_0442_),
    .A(\p_waveform[2] ),
    .B(_1343_));
 sg13g2_xor2_1 _1861_ (.B(_0442_),
    .A(_1347_),
    .X(_0443_));
 sg13g2_xor2_1 _1862_ (.B(_0443_),
    .A(_1357_),
    .X(_0444_));
 sg13g2_a221oi_1 _1863_ (.B2(net146),
    .C1(_1380_),
    .B1(_1360_),
    .A1(_0035_),
    .Y(_0445_),
    .A2(net142));
 sg13g2_inv_1 _1864_ (.Y(_0446_),
    .A(_0445_));
 sg13g2_a221oi_1 _1865_ (.B2(\p_waveform[4] ),
    .C1(_0446_),
    .B1(_0444_),
    .A1(net144),
    .Y(_0447_),
    .A2(net31));
 sg13g2_nand2_1 _1866_ (.Y(_0448_),
    .A(net24),
    .B(net23));
 sg13g2_xnor2_1 _1867_ (.Y(_0449_),
    .A(_1350_),
    .B(_0443_));
 sg13g2_a221oi_1 _1868_ (.B2(net146),
    .C1(_1380_),
    .B1(_1357_),
    .A1(_0034_),
    .Y(_0450_),
    .A2(net142));
 sg13g2_o21ai_1 _1869_ (.B1(_0450_),
    .Y(_0451_),
    .A1(_1231_),
    .A2(_0449_));
 sg13g2_a21oi_1 _1870_ (.A1(net143),
    .A2(net30),
    .Y(_0452_),
    .B1(_0451_));
 sg13g2_and3_1 _1871_ (.X(_0453_),
    .A(\p_env[4] ),
    .B(_0397_),
    .C(_0428_));
 sg13g2_o21ai_1 _1872_ (.B1(_1196_),
    .Y(_0454_),
    .A1(_1198_),
    .A2(_0399_));
 sg13g2_o21ai_1 _1873_ (.B1(_0421_),
    .Y(_0455_),
    .A1(_1397_),
    .A2(_0399_));
 sg13g2_nand2b_1 _1874_ (.Y(_0456_),
    .B(_0454_),
    .A_N(_0455_));
 sg13g2_xnor2_1 _1875_ (.Y(_0457_),
    .A(_1196_),
    .B(_1388_));
 sg13g2_inv_1 _1876_ (.Y(_0458_),
    .A(_0457_));
 sg13g2_mux2_1 _1877_ (.A0(_0457_),
    .A1(\p_sustain[0] ),
    .S(_0408_),
    .X(_0459_));
 sg13g2_mux2_1 _1878_ (.A0(_0457_),
    .A1(\p_env[4] ),
    .S(_0408_),
    .X(_0460_));
 sg13g2_a22oi_1 _1879_ (.Y(_0461_),
    .B1(_0460_),
    .B2(net112),
    .A2(_0459_),
    .A1(_0410_));
 sg13g2_a21oi_1 _1880_ (.A1(_0456_),
    .A2(_0461_),
    .Y(_0462_),
    .B1(_1189_));
 sg13g2_o21ai_1 _1881_ (.B1(_0393_),
    .Y(_0463_),
    .A1(_0453_),
    .A2(_0462_));
 sg13g2_a21oi_1 _1882_ (.A1(_0388_),
    .A2(_0458_),
    .Y(_0464_),
    .B1(net130));
 sg13g2_o21ai_1 _1883_ (.B1(_0464_),
    .Y(_0465_),
    .A1(\p_env[4] ),
    .A2(_0388_));
 sg13g2_nand2_1 _1884_ (.Y(_0466_),
    .A(_0463_),
    .B(_0465_));
 sg13g2_xnor2_1 _1885_ (.Y(_0467_),
    .A(\p_env[3] ),
    .B(_0399_));
 sg13g2_nor2_1 _1886_ (.A(_1198_),
    .B(_1387_),
    .Y(_0468_));
 sg13g2_nor3_1 _1887_ (.A(_1388_),
    .B(net32),
    .C(_0468_),
    .Y(_0469_));
 sg13g2_a21o_1 _1888_ (.A2(net32),
    .A1(_1198_),
    .B1(_0433_),
    .X(_0470_));
 sg13g2_a21o_1 _1889_ (.A2(_0470_),
    .A1(_0411_),
    .B1(_0469_),
    .X(_0471_));
 sg13g2_a221oi_1 _1890_ (.B2(_0422_),
    .C1(_0427_),
    .B1(_0467_),
    .A1(\p_env[3] ),
    .Y(_0472_),
    .A2(_0430_));
 sg13g2_a21oi_1 _1891_ (.A1(_0471_),
    .A2(_0472_),
    .Y(_0473_),
    .B1(_0394_));
 sg13g2_a21oi_1 _1892_ (.A1(_1198_),
    .A2(net32),
    .Y(_0474_),
    .B1(_0438_));
 sg13g2_nor2b_1 _1893_ (.A(_0469_),
    .B_N(_0474_),
    .Y(_0475_));
 sg13g2_nand3_1 _1894_ (.B(net134),
    .C(_1385_),
    .A(\p_env[3] ),
    .Y(_0476_));
 sg13g2_nor2_1 _1895_ (.A(_0473_),
    .B(_0475_),
    .Y(_0477_));
 sg13g2_nand2_1 _1896_ (.Y(_0478_),
    .A(_0476_),
    .B(_0477_));
 sg13g2_xnor2_1 _1897_ (.Y(_0479_),
    .A(_1353_),
    .B(_0443_));
 sg13g2_a221oi_1 _1898_ (.B2(net146),
    .C1(_1380_),
    .B1(_1350_),
    .A1(_0033_),
    .Y(_0480_),
    .A2(net142));
 sg13g2_o21ai_1 _1899_ (.B1(_0480_),
    .Y(_0481_),
    .A1(_1231_),
    .A2(_0479_));
 sg13g2_a21oi_1 _1900_ (.A1(net143),
    .A2(net30),
    .Y(_0482_),
    .B1(_0481_));
 sg13g2_nand2_1 _1901_ (.Y(_0483_),
    .A(net19),
    .B(_0482_));
 sg13g2_a221oi_1 _1902_ (.B2(_0477_),
    .C1(_0451_),
    .B1(_0476_),
    .A1(net143),
    .Y(_0484_),
    .A2(net30));
 sg13g2_a221oi_1 _1903_ (.B2(_0465_),
    .C1(_0481_),
    .B1(_0463_),
    .A1(net143),
    .Y(_0485_),
    .A2(net30));
 sg13g2_nand2_1 _1904_ (.Y(_0486_),
    .A(_0484_),
    .B(_0485_));
 sg13g2_nor2_1 _1905_ (.A(_0484_),
    .B(_0485_),
    .Y(_0487_));
 sg13g2_xor2_1 _1906_ (.B(_0485_),
    .A(_0484_),
    .X(_0488_));
 sg13g2_xnor2_1 _1907_ (.Y(_0489_),
    .A(_0448_),
    .B(_0488_));
 sg13g2_and2_1 _1908_ (.A(_0418_),
    .B(_0489_),
    .X(_0490_));
 sg13g2_nor3_1 _1909_ (.A(_1194_),
    .B(_1397_),
    .C(_0399_),
    .Y(_0491_));
 sg13g2_xnor2_1 _1910_ (.Y(_0492_),
    .A(net137),
    .B(_0491_));
 sg13g2_xnor2_1 _1911_ (.Y(_0493_),
    .A(_1192_),
    .B(_1393_));
 sg13g2_nor2_1 _1912_ (.A(net32),
    .B(_0493_),
    .Y(_0494_));
 sg13g2_a221oi_1 _1913_ (.B2(_0406_),
    .C1(_0411_),
    .B1(_0494_),
    .A1(_1191_),
    .Y(_0495_),
    .A2(_0408_));
 sg13g2_mux2_1 _1914_ (.A0(_0493_),
    .A1(net137),
    .S(net33),
    .X(_0496_));
 sg13g2_a22oi_1 _1915_ (.Y(_0497_),
    .B1(_0434_),
    .B2(_0496_),
    .A2(_0430_),
    .A1(net137));
 sg13g2_o21ai_1 _1916_ (.B1(_0497_),
    .Y(_0498_),
    .A1(_0423_),
    .A2(_0492_));
 sg13g2_o21ai_1 _1917_ (.B1(_0393_),
    .Y(_0499_),
    .A1(_0495_),
    .A2(_0498_));
 sg13g2_mux2_1 _1918_ (.A0(net137),
    .A1(_0496_),
    .S(_1396_),
    .X(_0500_));
 sg13g2_nand2_1 _1919_ (.Y(_0501_),
    .A(net134),
    .B(_0500_));
 sg13g2_nand2_1 _1920_ (.Y(_0502_),
    .A(_0499_),
    .B(_0501_));
 sg13g2_a221oi_1 _1921_ (.B2(_0501_),
    .C1(_0481_),
    .B1(_0499_),
    .A1(net143),
    .Y(_0503_),
    .A2(net30));
 sg13g2_nand2_1 _1922_ (.Y(_0504_),
    .A(_0482_),
    .B(net18));
 sg13g2_nand2_1 _1923_ (.Y(_0505_),
    .A(_0418_),
    .B(_0503_));
 sg13g2_a22oi_1 _1924_ (.Y(_0506_),
    .B1(net18),
    .B2(net28),
    .A2(_0482_),
    .A1(net26));
 sg13g2_a21oi_1 _1925_ (.A1(_0418_),
    .A2(_0503_),
    .Y(_0507_),
    .B1(_0506_));
 sg13g2_a21oi_1 _1926_ (.A1(_1360_),
    .A2(_0443_),
    .Y(_0508_),
    .B1(_1231_));
 sg13g2_o21ai_1 _1927_ (.B1(_0508_),
    .Y(_0509_),
    .A1(_1360_),
    .A2(_0443_));
 sg13g2_a221oi_1 _1928_ (.B2(net146),
    .C1(_1380_),
    .B1(_1364_),
    .A1(_0036_),
    .Y(_0510_),
    .A2(net142));
 sg13g2_nand3_1 _1929_ (.B(_0509_),
    .C(_0510_),
    .A(_1379_),
    .Y(_0511_));
 sg13g2_nand4_1 _1930_ (.B(net24),
    .C(_0509_),
    .A(_1379_),
    .Y(_0512_),
    .D(_0510_));
 sg13g2_nand2_1 _1931_ (.Y(_0513_),
    .A(net23),
    .B(net21));
 sg13g2_and3_1 _1932_ (.X(_0514_),
    .A(net23),
    .B(net21),
    .C(_0484_));
 sg13g2_a22oi_1 _1933_ (.Y(_0515_),
    .B1(net19),
    .B2(net23),
    .A2(net21),
    .A1(_0452_));
 sg13g2_or3_1 _1934_ (.A(_0512_),
    .B(_0514_),
    .C(_0515_),
    .X(_0516_));
 sg13g2_o21ai_1 _1935_ (.B1(_0512_),
    .Y(_0517_),
    .A1(_0514_),
    .A2(_0515_));
 sg13g2_nand3_1 _1936_ (.B(_0516_),
    .C(_0517_),
    .A(_0507_),
    .Y(_0518_));
 sg13g2_a21o_1 _1937_ (.A2(_0517_),
    .A1(_0516_),
    .B1(_0507_),
    .X(_0519_));
 sg13g2_nand3_1 _1938_ (.B(_0518_),
    .C(_0519_),
    .A(_0490_),
    .Y(_0520_));
 sg13g2_a21o_1 _1939_ (.A2(_0519_),
    .A1(_0518_),
    .B1(_0490_),
    .X(_0521_));
 sg13g2_o21ai_1 _1940_ (.B1(net134),
    .Y(_0522_),
    .A1(net141),
    .A2(_0388_));
 sg13g2_a21oi_1 _1941_ (.A1(net141),
    .A2(_0388_),
    .Y(_0523_),
    .B1(_0522_));
 sg13g2_nand2_1 _1942_ (.Y(_0524_),
    .A(_1200_),
    .B(_1209_));
 sg13g2_a21oi_1 _1943_ (.A1(\p_env[0] ),
    .A2(_0407_),
    .Y(_0525_),
    .B1(_1208_));
 sg13g2_o21ai_1 _1944_ (.B1(_0525_),
    .Y(_0526_),
    .A1(_0407_),
    .A2(_0524_));
 sg13g2_xnor2_1 _1945_ (.Y(_0527_),
    .A(\p_env[0] ),
    .B(net33));
 sg13g2_o21ai_1 _1946_ (.B1(_0428_),
    .Y(_0528_),
    .A1(_0397_),
    .A2(_0527_));
 sg13g2_a221oi_1 _1947_ (.B2(_0528_),
    .C1(_0394_),
    .B1(_0526_),
    .A1(_1189_),
    .Y(_0529_),
    .A2(_1200_));
 sg13g2_or2_1 _1948_ (.X(_0530_),
    .B(_0529_),
    .A(_0523_));
 sg13g2_xnor2_1 _1949_ (.Y(_0531_),
    .A(_1370_),
    .B(_0443_));
 sg13g2_a221oi_1 _1950_ (.B2(\p_waveform[5] ),
    .C1(_1380_),
    .B1(_1373_),
    .A1(_0038_),
    .Y(_0532_),
    .A2(net142));
 sg13g2_o21ai_1 _1951_ (.B1(_0532_),
    .Y(_0533_),
    .A1(_1231_),
    .A2(_0531_));
 sg13g2_a21oi_1 _1952_ (.A1(net144),
    .A2(net31),
    .Y(_0534_),
    .B1(_0533_));
 sg13g2_nand2_1 _1953_ (.Y(_0535_),
    .A(net17),
    .B(_0534_));
 sg13g2_o21ai_1 _1954_ (.B1(_0486_),
    .Y(_0536_),
    .A1(_0448_),
    .A2(_0487_));
 sg13g2_xnor2_1 _1955_ (.Y(_0537_),
    .A(net140),
    .B(net141));
 sg13g2_mux2_1 _1956_ (.A0(net140),
    .A1(_0537_),
    .S(_0388_),
    .X(_0538_));
 sg13g2_nand2b_1 _1957_ (.Y(_0539_),
    .B(_0423_),
    .A_N(_0537_));
 sg13g2_nand3_1 _1958_ (.B(_0433_),
    .C(_0537_),
    .A(_0411_),
    .Y(_0540_));
 sg13g2_a21o_1 _1959_ (.A2(_0540_),
    .A1(_0539_),
    .B1(net32),
    .X(_0541_));
 sg13g2_a22oi_1 _1960_ (.Y(_0542_),
    .B1(_0423_),
    .B2(_0433_),
    .A2(net32),
    .A1(_1199_));
 sg13g2_o21ai_1 _1961_ (.B1(_0541_),
    .Y(_0543_),
    .A1(_0412_),
    .A2(_0542_));
 sg13g2_a21oi_1 _1962_ (.A1(\p_env[1] ),
    .A2(_0430_),
    .Y(_0544_),
    .B1(_0427_));
 sg13g2_a21oi_1 _1963_ (.A1(_0543_),
    .A2(_0544_),
    .Y(_0545_),
    .B1(_0394_));
 sg13g2_a21o_1 _1964_ (.A2(_0538_),
    .A1(net134),
    .B1(_0545_),
    .X(_0546_));
 sg13g2_xor2_1 _1965_ (.B(_0443_),
    .A(_1364_),
    .X(_0547_));
 sg13g2_a21oi_1 _1966_ (.A1(_0037_),
    .A2(\p_waveform[7] ),
    .Y(_0548_),
    .B1(_1380_));
 sg13g2_o21ai_1 _1967_ (.B1(_0548_),
    .Y(_0549_),
    .A1(_1232_),
    .A2(_1369_));
 sg13g2_a221oi_1 _1968_ (.B2(\p_waveform[4] ),
    .C1(_0549_),
    .B1(_0547_),
    .A1(net145),
    .Y(_0550_),
    .A2(_1378_));
 sg13g2_nand2_1 _1969_ (.Y(_0551_),
    .A(net29),
    .B(_0550_));
 sg13g2_nand2b_1 _1970_ (.Y(_0552_),
    .B(_0536_),
    .A_N(_0551_));
 sg13g2_xor2_1 _1971_ (.B(_0551_),
    .A(_0536_),
    .X(_0553_));
 sg13g2_xor2_1 _1972_ (.B(_0553_),
    .A(_0535_),
    .X(_0554_));
 sg13g2_nand3_1 _1973_ (.B(_0521_),
    .C(_0554_),
    .A(_0520_),
    .Y(_0555_));
 sg13g2_and2_1 _1974_ (.A(_0520_),
    .B(_0555_),
    .X(_0556_));
 sg13g2_nand2_1 _1975_ (.Y(_0557_),
    .A(net24),
    .B(_0550_));
 sg13g2_nand4_1 _1976_ (.B(net21),
    .C(_0509_),
    .A(_1379_),
    .Y(_0558_),
    .D(_0510_));
 sg13g2_nand4_1 _1977_ (.B(net19),
    .C(_0509_),
    .A(_1379_),
    .Y(_0559_),
    .D(_0510_));
 sg13g2_xor2_1 _1978_ (.B(_0559_),
    .A(_0513_),
    .X(_0560_));
 sg13g2_nand2b_1 _1979_ (.Y(_0561_),
    .B(_0560_),
    .A_N(_0557_));
 sg13g2_xnor2_1 _1980_ (.Y(_0562_),
    .A(_0557_),
    .B(_0560_));
 sg13g2_nand2_1 _1981_ (.Y(_0563_),
    .A(net26),
    .B(_0452_));
 sg13g2_xnor2_1 _1982_ (.Y(_0564_),
    .A(_1188_),
    .B(_1394_));
 sg13g2_nor2_1 _1983_ (.A(net136),
    .B(net147),
    .Y(_0565_));
 sg13g2_nor4_1 _1984_ (.A(_1190_),
    .B(_1208_),
    .C(_1209_),
    .D(_0565_),
    .Y(_0566_));
 sg13g2_a21oi_1 _1985_ (.A1(\p_env[7] ),
    .A2(net112),
    .Y(_0567_),
    .B1(_0566_));
 sg13g2_nor3_1 _1986_ (.A(_1399_),
    .B(net33),
    .C(_0395_),
    .Y(_0568_));
 sg13g2_nor2_1 _1987_ (.A(\p_env[7] ),
    .B(_0568_),
    .Y(_0569_));
 sg13g2_nor3_1 _1988_ (.A(_1425_),
    .B(_0565_),
    .C(_0569_),
    .Y(_0570_));
 sg13g2_nand2_1 _1989_ (.Y(_0571_),
    .A(\p_env[7] ),
    .B(_0402_));
 sg13g2_nand4_1 _1990_ (.B(\p_ast[1] ),
    .C(_0407_),
    .A(cur_gate),
    .Y(_0572_),
    .D(_0564_));
 sg13g2_o21ai_1 _1991_ (.B1(_0571_),
    .Y(_0573_),
    .A1(_0407_),
    .A2(_0567_));
 sg13g2_nand2b_1 _1992_ (.Y(_0574_),
    .B(_0572_),
    .A_N(_0573_));
 sg13g2_o21ai_1 _1993_ (.B1(_0393_),
    .Y(_0575_),
    .A1(_0570_),
    .A2(_0574_));
 sg13g2_a21oi_1 _1994_ (.A1(_1394_),
    .A2(_0388_),
    .Y(_0576_),
    .B1(net130));
 sg13g2_nand2_1 _1995_ (.Y(_0577_),
    .A(net136),
    .B(_0576_));
 sg13g2_nand2_1 _1996_ (.Y(_0578_),
    .A(_0575_),
    .B(_0577_));
 sg13g2_a221oi_1 _1997_ (.B2(_0577_),
    .C1(_0481_),
    .B1(_0575_),
    .A1(net143),
    .Y(_0579_),
    .A2(net30));
 sg13g2_a221oi_1 _1998_ (.B2(_0577_),
    .C1(_1383_),
    .B1(_0575_),
    .A1(net143),
    .Y(_0580_),
    .A2(net30));
 sg13g2_nand2_1 _1999_ (.Y(_0581_),
    .A(_0503_),
    .B(_0580_));
 sg13g2_nor2_1 _2000_ (.A(_0503_),
    .B(_0580_),
    .Y(_0582_));
 sg13g2_xor2_1 _2001_ (.B(_0580_),
    .A(_0503_),
    .X(_0583_));
 sg13g2_xnor2_1 _2002_ (.Y(_0584_),
    .A(_0563_),
    .B(_0583_));
 sg13g2_nor2b_1 _2003_ (.A(_0505_),
    .B_N(_0584_),
    .Y(_0585_));
 sg13g2_xnor2_1 _2004_ (.Y(_0586_),
    .A(_0505_),
    .B(_0584_));
 sg13g2_xnor2_1 _2005_ (.Y(_0587_),
    .A(_0562_),
    .B(_0586_));
 sg13g2_nor2_1 _2006_ (.A(_0518_),
    .B(_0587_),
    .Y(_0588_));
 sg13g2_xor2_1 _2007_ (.B(_0587_),
    .A(_0518_),
    .X(_0589_));
 sg13g2_xnor2_1 _2008_ (.Y(_0590_),
    .A(_1373_),
    .B(_0443_));
 sg13g2_a221oi_1 _2009_ (.B2(net146),
    .C1(_1380_),
    .B1(_1347_),
    .A1(_0039_),
    .Y(_0591_),
    .A2(\p_waveform[7] ));
 sg13g2_o21ai_1 _2010_ (.B1(_0591_),
    .Y(_0592_),
    .A1(_1231_),
    .A2(_0590_));
 sg13g2_a21oi_1 _2011_ (.A1(net144),
    .A2(net31),
    .Y(_0593_),
    .B1(_0592_));
 sg13g2_nand2_1 _2012_ (.Y(_0594_),
    .A(net17),
    .B(_0593_));
 sg13g2_nand2b_1 _2013_ (.Y(_0595_),
    .B(_0516_),
    .A_N(_0514_));
 sg13g2_nand2_1 _2014_ (.Y(_0596_),
    .A(_0534_),
    .B(net29));
 sg13g2_nand2b_1 _2015_ (.Y(_0597_),
    .B(_0595_),
    .A_N(_0596_));
 sg13g2_xor2_1 _2016_ (.B(_0596_),
    .A(_0595_),
    .X(_0598_));
 sg13g2_xor2_1 _2017_ (.B(_0598_),
    .A(_0594_),
    .X(_0599_));
 sg13g2_xnor2_1 _2018_ (.Y(_0600_),
    .A(_0589_),
    .B(_0599_));
 sg13g2_nor2_1 _2019_ (.A(_0556_),
    .B(_0600_),
    .Y(_0601_));
 sg13g2_o21ai_1 _2020_ (.B1(_0552_),
    .Y(_0602_),
    .A1(_0535_),
    .A2(_0553_));
 sg13g2_xor2_1 _2021_ (.B(_0600_),
    .A(_0556_),
    .X(_0603_));
 sg13g2_and2_1 _2022_ (.A(_0602_),
    .B(_0603_),
    .X(_0604_));
 sg13g2_a21oi_1 _2023_ (.A1(_0602_),
    .A2(_0603_),
    .Y(_0605_),
    .B1(_0601_));
 sg13g2_o21ai_1 _2024_ (.B1(_0597_),
    .Y(_0606_),
    .A1(_0594_),
    .A2(_0598_));
 sg13g2_a21oi_1 _2025_ (.A1(_0589_),
    .A2(_0599_),
    .Y(_0607_),
    .B1(_0588_));
 sg13g2_o21ai_1 _2026_ (.B1(_0561_),
    .Y(_0608_),
    .A1(_0513_),
    .A2(_0559_));
 sg13g2_nand2_1 _2027_ (.Y(_0609_),
    .A(net29),
    .B(_0593_));
 sg13g2_nor2b_1 _2028_ (.A(_0609_),
    .B_N(_0608_),
    .Y(_0610_));
 sg13g2_xor2_1 _2029_ (.B(_0609_),
    .A(_0608_),
    .X(_0611_));
 sg13g2_a21oi_1 _2030_ (.A1(_0562_),
    .A2(_0586_),
    .Y(_0612_),
    .B1(_0585_));
 sg13g2_nand2_1 _2031_ (.Y(_0613_),
    .A(net24),
    .B(_0534_));
 sg13g2_nand2_1 _2032_ (.Y(_0614_),
    .A(net21),
    .B(_0550_));
 sg13g2_nand2_1 _2033_ (.Y(_0615_),
    .A(net19),
    .B(_0550_));
 sg13g2_xor2_1 _2034_ (.B(_0615_),
    .A(_0558_),
    .X(_0616_));
 sg13g2_nand2b_1 _2035_ (.Y(_0617_),
    .B(_0616_),
    .A_N(_0613_));
 sg13g2_xnor2_1 _2036_ (.Y(_0618_),
    .A(_0613_),
    .B(_0616_));
 sg13g2_o21ai_1 _2037_ (.B1(_0581_),
    .Y(_0619_),
    .A1(_0563_),
    .A2(_0582_));
 sg13g2_and2_1 _2038_ (.A(net27),
    .B(net23),
    .X(_0620_));
 sg13g2_nand2_1 _2039_ (.Y(_0621_),
    .A(_0452_),
    .B(net16));
 sg13g2_a221oi_1 _2040_ (.B2(_0501_),
    .C1(_0451_),
    .B1(_0499_),
    .A1(net144),
    .Y(_0622_),
    .A2(net31));
 sg13g2_xor2_1 _2041_ (.B(_0622_),
    .A(_0579_),
    .X(_0623_));
 sg13g2_nand2_1 _2042_ (.Y(_0624_),
    .A(_0620_),
    .B(_0623_));
 sg13g2_xor2_1 _2043_ (.B(_0623_),
    .A(_0620_),
    .X(_0625_));
 sg13g2_and2_1 _2044_ (.A(_0619_),
    .B(_0625_),
    .X(_0626_));
 sg13g2_xor2_1 _2045_ (.B(_0625_),
    .A(_0619_),
    .X(_0627_));
 sg13g2_xnor2_1 _2046_ (.Y(_0628_),
    .A(_0618_),
    .B(_0627_));
 sg13g2_xor2_1 _2047_ (.B(_0628_),
    .A(_0612_),
    .X(_0629_));
 sg13g2_nand2b_1 _2048_ (.Y(_0630_),
    .B(_0629_),
    .A_N(_0611_));
 sg13g2_xnor2_1 _2049_ (.Y(_0631_),
    .A(_0611_),
    .B(_0629_));
 sg13g2_nor2b_1 _2050_ (.A(_0607_),
    .B_N(_0631_),
    .Y(_0632_));
 sg13g2_xnor2_1 _2051_ (.Y(_0633_),
    .A(_0607_),
    .B(_0631_));
 sg13g2_xnor2_1 _2052_ (.Y(_0634_),
    .A(_0606_),
    .B(_0633_));
 sg13g2_nor2_1 _2053_ (.A(_0605_),
    .B(_0634_),
    .Y(_0635_));
 sg13g2_or3_1 _2054_ (.A(_0601_),
    .B(_0604_),
    .C(_0634_),
    .X(_0636_));
 sg13g2_nand2b_1 _2055_ (.Y(_0637_),
    .B(_0634_),
    .A_N(_0605_));
 sg13g2_and2_1 _2056_ (.A(_0636_),
    .B(_0637_),
    .X(_0638_));
 sg13g2_xnor2_1 _2057_ (.Y(_0639_),
    .A(_0602_),
    .B(_0603_));
 sg13g2_xnor2_1 _2058_ (.Y(_0640_),
    .A(_0419_),
    .B(_0489_));
 sg13g2_nand2_1 _2059_ (.Y(_0641_),
    .A(net17),
    .B(_0550_));
 sg13g2_nand2_1 _2060_ (.Y(_0642_),
    .A(net28),
    .B(net19));
 sg13g2_nand2_1 _2061_ (.Y(_0643_),
    .A(net28),
    .B(net21));
 sg13g2_nand3_1 _2062_ (.B(net19),
    .C(_0485_),
    .A(net28),
    .Y(_0644_));
 sg13g2_nand2_1 _2063_ (.Y(_0645_),
    .A(net24),
    .B(_0452_));
 sg13g2_a22oi_1 _2064_ (.Y(_0646_),
    .B1(net20),
    .B2(_0482_),
    .A2(net22),
    .A1(net28));
 sg13g2_xor2_1 _2065_ (.B(_0643_),
    .A(_0483_),
    .X(_0647_));
 sg13g2_o21ai_1 _2066_ (.B1(_0644_),
    .Y(_0648_),
    .A1(_0645_),
    .A2(_0646_));
 sg13g2_nand2b_1 _2067_ (.Y(_0649_),
    .B(net29),
    .A_N(_0511_));
 sg13g2_nand2b_1 _2068_ (.Y(_0650_),
    .B(_0648_),
    .A_N(_0649_));
 sg13g2_xor2_1 _2069_ (.B(_0649_),
    .A(_0648_),
    .X(_0651_));
 sg13g2_xor2_1 _2070_ (.B(_0651_),
    .A(_0641_),
    .X(_0652_));
 sg13g2_and2_1 _2071_ (.A(_0640_),
    .B(_0652_),
    .X(_0653_));
 sg13g2_a21o_1 _2072_ (.A2(_0521_),
    .A1(_0520_),
    .B1(_0554_),
    .X(_0654_));
 sg13g2_and2_1 _2073_ (.A(_0555_),
    .B(_0654_),
    .X(_0655_));
 sg13g2_nand3_1 _2074_ (.B(_0653_),
    .C(_0654_),
    .A(_0555_),
    .Y(_0656_));
 sg13g2_o21ai_1 _2075_ (.B1(_0650_),
    .Y(_0657_),
    .A1(_0641_),
    .A2(_0651_));
 sg13g2_a21o_1 _2076_ (.A2(_0654_),
    .A1(_0555_),
    .B1(_0653_),
    .X(_0658_));
 sg13g2_and3_1 _2077_ (.X(_0659_),
    .A(_0656_),
    .B(_0657_),
    .C(_0658_));
 sg13g2_a21oi_1 _2078_ (.A1(_0653_),
    .A2(_0655_),
    .Y(_0660_),
    .B1(_0659_));
 sg13g2_and2_1 _2079_ (.A(_0639_),
    .B(_0660_),
    .X(_0661_));
 sg13g2_or2_1 _2080_ (.X(_0662_),
    .B(_0660_),
    .A(_0639_));
 sg13g2_a21oi_1 _2081_ (.A1(_0656_),
    .A2(_0658_),
    .Y(_0663_),
    .B1(_0657_));
 sg13g2_nand2_1 _2082_ (.Y(_0664_),
    .A(net23),
    .B(net29));
 sg13g2_nand2_1 _2083_ (.Y(_0665_),
    .A(net28),
    .B(net24));
 sg13g2_nand2_1 _2084_ (.Y(_0666_),
    .A(net24),
    .B(_0482_));
 sg13g2_or2_1 _2085_ (.X(_0667_),
    .B(_0665_),
    .A(_0483_));
 sg13g2_nor2_1 _2086_ (.A(_0664_),
    .B(_0667_),
    .Y(_0668_));
 sg13g2_nand2b_1 _2087_ (.Y(_0669_),
    .B(net17),
    .A_N(_0511_));
 sg13g2_xor2_1 _2088_ (.B(_0667_),
    .A(_0664_),
    .X(_0670_));
 sg13g2_nor2b_1 _2089_ (.A(_0669_),
    .B_N(_0670_),
    .Y(_0671_));
 sg13g2_nor2_1 _2090_ (.A(_0668_),
    .B(_0671_),
    .Y(_0672_));
 sg13g2_inv_1 _2091_ (.Y(_0673_),
    .A(_0672_));
 sg13g2_xnor2_1 _2092_ (.Y(_0674_),
    .A(_0645_),
    .B(_0647_));
 sg13g2_xnor2_1 _2093_ (.Y(_0675_),
    .A(_0669_),
    .B(_0670_));
 sg13g2_nand2_1 _2094_ (.Y(_0676_),
    .A(_0674_),
    .B(_0675_));
 sg13g2_xnor2_1 _2095_ (.Y(_0677_),
    .A(_0640_),
    .B(_0652_));
 sg13g2_nor2_1 _2096_ (.A(_0676_),
    .B(_0677_),
    .Y(_0678_));
 sg13g2_xor2_1 _2097_ (.B(_0677_),
    .A(_0676_),
    .X(_0679_));
 sg13g2_xor2_1 _2098_ (.B(_0675_),
    .A(_0674_),
    .X(_0680_));
 sg13g2_nand2_1 _2099_ (.Y(_0681_),
    .A(_0452_),
    .B(net17));
 sg13g2_nor2_1 _2100_ (.A(_0664_),
    .B(_0681_),
    .Y(_0682_));
 sg13g2_nand2_1 _2101_ (.Y(_0683_),
    .A(_0680_),
    .B(_0682_));
 sg13g2_xor2_1 _2102_ (.B(_0666_),
    .A(_0642_),
    .X(_0684_));
 sg13g2_a22oi_1 _2103_ (.Y(_0685_),
    .B1(net29),
    .B2(_0452_),
    .A2(net17),
    .A1(net23));
 sg13g2_nor2_1 _2104_ (.A(_0682_),
    .B(_0685_),
    .Y(_0686_));
 sg13g2_nand2_1 _2105_ (.Y(_0687_),
    .A(_0684_),
    .B(_0686_));
 sg13g2_inv_1 _2106_ (.Y(_0688_),
    .A(_0687_));
 sg13g2_nand2_1 _2107_ (.Y(_0689_),
    .A(_0482_),
    .B(net29));
 sg13g2_or2_1 _2108_ (.X(_0690_),
    .B(_0681_),
    .A(_0665_));
 sg13g2_nor2_1 _2109_ (.A(_0689_),
    .B(_0690_),
    .Y(_0691_));
 sg13g2_nor2_1 _2110_ (.A(_0684_),
    .B(_0686_),
    .Y(_0692_));
 sg13g2_a22oi_1 _2111_ (.Y(_0693_),
    .B1(net17),
    .B2(_1382_),
    .A2(net25),
    .A1(_1384_));
 sg13g2_a221oi_1 _2112_ (.B2(_0681_),
    .C1(_0692_),
    .B1(_0693_),
    .A1(_0689_),
    .Y(_0694_),
    .A2(_0690_));
 sg13g2_nor3_1 _2113_ (.A(_0688_),
    .B(_0691_),
    .C(_0694_),
    .Y(_0695_));
 sg13g2_nand2_1 _2114_ (.Y(_0696_),
    .A(_0688_),
    .B(_0691_));
 sg13g2_nor2_1 _2115_ (.A(_0680_),
    .B(_0682_),
    .Y(_0697_));
 sg13g2_a21oi_1 _2116_ (.A1(_0673_),
    .A2(_0679_),
    .Y(_0698_),
    .B1(_0678_));
 sg13g2_nor3_1 _2117_ (.A(_0659_),
    .B(_0663_),
    .C(_0698_),
    .Y(_0699_));
 sg13g2_xnor2_1 _2118_ (.Y(_0700_),
    .A(_0673_),
    .B(_0679_));
 sg13g2_a221oi_1 _2119_ (.B2(_0697_),
    .C1(_0700_),
    .B1(_0696_),
    .A1(_0683_),
    .Y(_0701_),
    .A2(_0695_));
 sg13g2_o21ai_1 _2120_ (.B1(_0698_),
    .Y(_0702_),
    .A1(_0659_),
    .A2(_0663_));
 sg13g2_o21ai_1 _2121_ (.B1(_0702_),
    .Y(_0703_),
    .A1(_0699_),
    .A2(_0701_));
 sg13g2_a21o_1 _2122_ (.A2(_0703_),
    .A1(_0662_),
    .B1(_0661_),
    .X(_0704_));
 sg13g2_a221oi_1 _2123_ (.B2(_0703_),
    .C1(_0661_),
    .B1(_0662_),
    .A1(_0636_),
    .Y(_0705_),
    .A2(_0637_));
 sg13g2_xnor2_1 _2124_ (.Y(_0706_),
    .A(_0638_),
    .B(_0704_));
 sg13g2_nand2_1 _2125_ (.Y(_0707_),
    .A(net358),
    .B(_1340_));
 sg13g2_xnor2_1 _2126_ (.Y(_0708_),
    .A(_0706_),
    .B(_0707_));
 sg13g2_or3_1 _2127_ (.A(net131),
    .B(net119),
    .C(_0708_),
    .X(_0709_));
 sg13g2_o21ai_1 _2128_ (.B1(_0709_),
    .Y(_0303_),
    .A1(_1220_),
    .A2(_1243_));
 sg13g2_a21oi_1 _2129_ (.A1(_0606_),
    .A2(_0633_),
    .Y(_0710_),
    .B1(_0632_));
 sg13g2_o21ai_1 _2130_ (.B1(_0630_),
    .Y(_0711_),
    .A1(_0612_),
    .A2(_0628_));
 sg13g2_o21ai_1 _2131_ (.B1(_0617_),
    .Y(_0712_),
    .A1(_0558_),
    .A2(_0615_));
 sg13g2_a21oi_1 _2132_ (.A1(_0618_),
    .A2(_0627_),
    .Y(_0713_),
    .B1(_0626_));
 sg13g2_nand2_1 _2133_ (.Y(_0714_),
    .A(net24),
    .B(_0593_));
 sg13g2_nand2_1 _2134_ (.Y(_0715_),
    .A(net19),
    .B(_0534_));
 sg13g2_xor2_1 _2135_ (.B(_0715_),
    .A(_0614_),
    .X(_0716_));
 sg13g2_nand2b_1 _2136_ (.Y(_0717_),
    .B(_0716_),
    .A_N(_0714_));
 sg13g2_xnor2_1 _2137_ (.Y(_0718_),
    .A(_0714_),
    .B(_0716_));
 sg13g2_o21ai_1 _2138_ (.B1(_0624_),
    .Y(_0719_),
    .A1(_0504_),
    .A2(_0621_));
 sg13g2_nand2b_1 _2139_ (.Y(_0720_),
    .B(net26),
    .A_N(_0511_));
 sg13g2_nand2_1 _2140_ (.Y(_0721_),
    .A(net23),
    .B(net16));
 sg13g2_nand2_1 _2141_ (.Y(_0722_),
    .A(_0447_),
    .B(net18));
 sg13g2_xor2_1 _2142_ (.B(_0722_),
    .A(_0621_),
    .X(_0723_));
 sg13g2_nand2b_1 _2143_ (.Y(_0724_),
    .B(_0723_),
    .A_N(_0720_));
 sg13g2_xnor2_1 _2144_ (.Y(_0725_),
    .A(_0720_),
    .B(_0723_));
 sg13g2_and2_1 _2145_ (.A(_0719_),
    .B(_0725_),
    .X(_0726_));
 sg13g2_xor2_1 _2146_ (.B(_0725_),
    .A(_0719_),
    .X(_0727_));
 sg13g2_xnor2_1 _2147_ (.Y(_0728_),
    .A(_0718_),
    .B(_0727_));
 sg13g2_nor2_1 _2148_ (.A(_0713_),
    .B(_0728_),
    .Y(_0729_));
 sg13g2_xor2_1 _2149_ (.B(_0728_),
    .A(_0713_),
    .X(_0730_));
 sg13g2_xnor2_1 _2150_ (.Y(_0731_),
    .A(_0712_),
    .B(_0730_));
 sg13g2_nor2b_1 _2151_ (.A(_0731_),
    .B_N(_0711_),
    .Y(_0732_));
 sg13g2_xnor2_1 _2152_ (.Y(_0733_),
    .A(_0711_),
    .B(_0731_));
 sg13g2_xnor2_1 _2153_ (.Y(_0734_),
    .A(_0610_),
    .B(_0733_));
 sg13g2_or2_1 _2154_ (.X(_0735_),
    .B(_0734_),
    .A(_0710_));
 sg13g2_xor2_1 _2155_ (.B(_0734_),
    .A(_0710_),
    .X(_0736_));
 sg13g2_or3_1 _2156_ (.A(_0635_),
    .B(_0705_),
    .C(_0736_),
    .X(_0737_));
 sg13g2_o21ai_1 _2157_ (.B1(_0736_),
    .Y(_0738_),
    .A1(_0635_),
    .A2(_0705_));
 sg13g2_and2_1 _2158_ (.A(_0737_),
    .B(_0738_),
    .X(_0739_));
 sg13g2_nand3_1 _2159_ (.B(_0737_),
    .C(_0738_),
    .A(net688),
    .Y(_0740_));
 sg13g2_a21oi_1 _2160_ (.A1(_0737_),
    .A2(_0738_),
    .Y(_0741_),
    .B1(net688));
 sg13g2_xnor2_1 _2161_ (.Y(_0742_),
    .A(_1244_),
    .B(_0739_));
 sg13g2_or2_1 _2162_ (.X(_0743_),
    .B(_0706_),
    .A(_1243_));
 sg13g2_nor2_1 _2163_ (.A(net132),
    .B(_1271_),
    .Y(_0744_));
 sg13g2_nand2b_1 _2164_ (.Y(_0745_),
    .B(_1220_),
    .A_N(_1270_));
 sg13g2_a21oi_1 _2165_ (.A1(_1270_),
    .A2(_1271_),
    .Y(_0746_),
    .B1(net132));
 sg13g2_inv_1 _2166_ (.Y(_0747_),
    .A(_0746_));
 sg13g2_xnor2_1 _2167_ (.Y(_0748_),
    .A(_0742_),
    .B(_0743_));
 sg13g2_a221oi_1 _2168_ (.B2(_0748_),
    .C1(net131),
    .B1(_0746_),
    .A1(_1339_),
    .Y(_0749_),
    .A2(_0739_));
 sg13g2_a21oi_1 _2169_ (.A1(net131),
    .A2(_1244_),
    .Y(_0304_),
    .B1(_0749_));
 sg13g2_a21oi_1 _2170_ (.A1(_0712_),
    .A2(_0730_),
    .Y(_0750_),
    .B1(_0729_));
 sg13g2_o21ai_1 _2171_ (.B1(_0717_),
    .Y(_0751_),
    .A1(_0614_),
    .A2(_0715_));
 sg13g2_a21oi_1 _2172_ (.A1(_0718_),
    .A2(_0727_),
    .Y(_0752_),
    .B1(_0726_));
 sg13g2_nand2_1 _2173_ (.Y(_0753_),
    .A(net21),
    .B(_0593_));
 sg13g2_nor2_1 _2174_ (.A(_0715_),
    .B(_0753_),
    .Y(_0754_));
 sg13g2_or2_1 _2175_ (.X(_0755_),
    .B(_0753_),
    .A(_0715_));
 sg13g2_a22oi_1 _2176_ (.Y(_0756_),
    .B1(_0593_),
    .B2(net19),
    .A2(_0534_),
    .A1(net21));
 sg13g2_or2_1 _2177_ (.X(_0757_),
    .B(_0756_),
    .A(_0754_));
 sg13g2_o21ai_1 _2178_ (.B1(_0724_),
    .Y(_0758_),
    .A1(_0621_),
    .A2(_0722_));
 sg13g2_nand2_1 _2179_ (.Y(_0759_),
    .A(net26),
    .B(_0550_));
 sg13g2_nor2b_1 _2180_ (.A(_0511_),
    .B_N(net16),
    .Y(_0760_));
 sg13g2_nand2b_1 _2181_ (.Y(_0761_),
    .B(net18),
    .A_N(_0511_));
 sg13g2_xor2_1 _2182_ (.B(_0761_),
    .A(_0721_),
    .X(_0762_));
 sg13g2_nand2b_1 _2183_ (.Y(_0763_),
    .B(_0762_),
    .A_N(_0759_));
 sg13g2_xnor2_1 _2184_ (.Y(_0764_),
    .A(_0759_),
    .B(_0762_));
 sg13g2_nand2_1 _2185_ (.Y(_0765_),
    .A(_0758_),
    .B(_0764_));
 sg13g2_xnor2_1 _2186_ (.Y(_0766_),
    .A(_0758_),
    .B(_0764_));
 sg13g2_xnor2_1 _2187_ (.Y(_0767_),
    .A(_0757_),
    .B(_0766_));
 sg13g2_nor2_1 _2188_ (.A(_0752_),
    .B(_0767_),
    .Y(_0768_));
 sg13g2_xor2_1 _2189_ (.B(_0767_),
    .A(_0752_),
    .X(_0769_));
 sg13g2_xnor2_1 _2190_ (.Y(_0770_),
    .A(_0751_),
    .B(_0769_));
 sg13g2_or2_1 _2191_ (.X(_0771_),
    .B(_0770_),
    .A(_0750_));
 sg13g2_xor2_1 _2192_ (.B(_0770_),
    .A(_0750_),
    .X(_0772_));
 sg13g2_a21oi_1 _2193_ (.A1(_0610_),
    .A2(_0733_),
    .Y(_0773_),
    .B1(_0732_));
 sg13g2_nand2b_1 _2194_ (.Y(_0774_),
    .B(_0772_),
    .A_N(_0773_));
 sg13g2_xor2_1 _2195_ (.B(_0773_),
    .A(_0772_),
    .X(_0775_));
 sg13g2_a21oi_1 _2196_ (.A1(_0735_),
    .A2(_0738_),
    .Y(_0776_),
    .B1(_0775_));
 sg13g2_a21o_1 _2197_ (.A2(_0738_),
    .A1(_0735_),
    .B1(_0775_),
    .X(_0777_));
 sg13g2_and3_1 _2198_ (.X(_0778_),
    .A(_0735_),
    .B(_0738_),
    .C(_0775_));
 sg13g2_nor3_1 _2199_ (.A(_1245_),
    .B(_0776_),
    .C(_0778_),
    .Y(_0779_));
 sg13g2_o21ai_1 _2200_ (.B1(_1245_),
    .Y(_0780_),
    .A1(_0776_),
    .A2(_0778_));
 sg13g2_nand2b_1 _2201_ (.Y(_0781_),
    .B(_0780_),
    .A_N(_0779_));
 sg13g2_o21ai_1 _2202_ (.B1(_0740_),
    .Y(_0782_),
    .A1(_0741_),
    .A2(_0743_));
 sg13g2_nand2b_1 _2203_ (.Y(_0783_),
    .B(_0781_),
    .A_N(_0782_));
 sg13g2_nand2b_1 _2204_ (.Y(_0784_),
    .B(_0782_),
    .A_N(_0781_));
 sg13g2_nand3_1 _2205_ (.B(_0783_),
    .C(_0784_),
    .A(_0746_),
    .Y(_0785_));
 sg13g2_nor3_1 _2206_ (.A(_1340_),
    .B(_0776_),
    .C(_0778_),
    .Y(_0786_));
 sg13g2_nor2_1 _2207_ (.A(net131),
    .B(_0786_),
    .Y(_0787_));
 sg13g2_a22oi_1 _2208_ (.Y(_0305_),
    .B1(_0785_),
    .B2(_0787_),
    .A2(_1245_),
    .A1(net131));
 sg13g2_a21oi_1 _2209_ (.A1(_0780_),
    .A2(_0782_),
    .Y(_0788_),
    .B1(_0779_));
 sg13g2_a21oi_1 _2210_ (.A1(_0751_),
    .A2(_0769_),
    .Y(_0789_),
    .B1(_0768_));
 sg13g2_o21ai_1 _2211_ (.B1(_0765_),
    .Y(_0790_),
    .A1(_0757_),
    .A2(_0766_));
 sg13g2_o21ai_1 _2212_ (.B1(_0763_),
    .Y(_0791_),
    .A1(_0721_),
    .A2(_0761_));
 sg13g2_nand2_1 _2213_ (.Y(_0792_),
    .A(net26),
    .B(_0534_));
 sg13g2_nand2_1 _2214_ (.Y(_0793_),
    .A(_0550_),
    .B(net16));
 sg13g2_nand2_1 _2215_ (.Y(_0794_),
    .A(net18),
    .B(_0550_));
 sg13g2_nor2_1 _2216_ (.A(_0761_),
    .B(_0793_),
    .Y(_0795_));
 sg13g2_xnor2_1 _2217_ (.Y(_0796_),
    .A(_0760_),
    .B(_0794_));
 sg13g2_nor2b_1 _2218_ (.A(_0792_),
    .B_N(_0796_),
    .Y(_0797_));
 sg13g2_xnor2_1 _2219_ (.Y(_0798_),
    .A(_0792_),
    .B(_0796_));
 sg13g2_nand2_1 _2220_ (.Y(_0799_),
    .A(_0791_),
    .B(_0798_));
 sg13g2_xnor2_1 _2221_ (.Y(_0800_),
    .A(_0791_),
    .B(_0798_));
 sg13g2_xor2_1 _2222_ (.B(_0800_),
    .A(_0753_),
    .X(_0801_));
 sg13g2_and2_1 _2223_ (.A(_0790_),
    .B(_0801_),
    .X(_0802_));
 sg13g2_xnor2_1 _2224_ (.Y(_0803_),
    .A(_0790_),
    .B(_0801_));
 sg13g2_nor2_1 _2225_ (.A(_0755_),
    .B(_0803_),
    .Y(_0804_));
 sg13g2_xor2_1 _2226_ (.B(_0803_),
    .A(_0755_),
    .X(_0805_));
 sg13g2_nor2b_1 _2227_ (.A(_0789_),
    .B_N(_0805_),
    .Y(_0806_));
 sg13g2_xor2_1 _2228_ (.B(_0805_),
    .A(_0789_),
    .X(_0807_));
 sg13g2_and2_1 _2229_ (.A(_0771_),
    .B(_0807_),
    .X(_0808_));
 sg13g2_or2_1 _2230_ (.X(_0809_),
    .B(_0807_),
    .A(_0771_));
 sg13g2_nand2b_1 _2231_ (.Y(_0810_),
    .B(_0809_),
    .A_N(_0808_));
 sg13g2_nand3_1 _2232_ (.B(_0777_),
    .C(_0810_),
    .A(_0774_),
    .Y(_0811_));
 sg13g2_a21o_1 _2233_ (.A2(_0777_),
    .A1(_0774_),
    .B1(_0810_),
    .X(_0812_));
 sg13g2_nand2_1 _2234_ (.Y(_0813_),
    .A(_0811_),
    .B(_0812_));
 sg13g2_nand3_1 _2235_ (.B(_0811_),
    .C(_0812_),
    .A(net724),
    .Y(_0814_));
 sg13g2_a21oi_1 _2236_ (.A1(_0811_),
    .A2(_0812_),
    .Y(_0815_),
    .B1(net724));
 sg13g2_xnor2_1 _2237_ (.Y(_0816_),
    .A(net724),
    .B(_0813_));
 sg13g2_nand2b_1 _2238_ (.Y(_0817_),
    .B(_0816_),
    .A_N(_0788_));
 sg13g2_nor2b_1 _2239_ (.A(_0816_),
    .B_N(_0788_),
    .Y(_0818_));
 sg13g2_nand3b_1 _2240_ (.B(_0746_),
    .C(_0817_),
    .Y(_0819_),
    .A_N(_0818_));
 sg13g2_o21ai_1 _2241_ (.B1(_0819_),
    .Y(_0820_),
    .A1(_1340_),
    .A2(_0813_));
 sg13g2_mux2_1 _2242_ (.A0(net724),
    .A1(_0820_),
    .S(_1220_),
    .X(_0306_));
 sg13g2_nand2_1 _2243_ (.Y(_0821_),
    .A(net26),
    .B(_0593_));
 sg13g2_nand2_1 _2244_ (.Y(_0822_),
    .A(_0534_),
    .B(net16));
 sg13g2_nand2_1 _2245_ (.Y(_0823_),
    .A(net18),
    .B(_0534_));
 sg13g2_nor2_1 _2246_ (.A(_0793_),
    .B(_0823_),
    .Y(_0824_));
 sg13g2_xor2_1 _2247_ (.B(_0823_),
    .A(_0793_),
    .X(_0825_));
 sg13g2_nor2b_1 _2248_ (.A(_0821_),
    .B_N(_0825_),
    .Y(_0826_));
 sg13g2_xnor2_1 _2249_ (.Y(_0827_),
    .A(_0821_),
    .B(_0825_));
 sg13g2_o21ai_1 _2250_ (.B1(_0827_),
    .Y(_0828_),
    .A1(_0795_),
    .A2(_0797_));
 sg13g2_or3_1 _2251_ (.A(_0795_),
    .B(_0797_),
    .C(_0827_),
    .X(_0829_));
 sg13g2_and2_1 _2252_ (.A(_0828_),
    .B(_0829_),
    .X(_0830_));
 sg13g2_o21ai_1 _2253_ (.B1(_0799_),
    .Y(_0831_),
    .A1(_0753_),
    .A2(_0800_));
 sg13g2_nand2_1 _2254_ (.Y(_0832_),
    .A(_0830_),
    .B(_0831_));
 sg13g2_xor2_1 _2255_ (.B(_0831_),
    .A(_0830_),
    .X(_0833_));
 sg13g2_o21ai_1 _2256_ (.B1(_0833_),
    .Y(_0834_),
    .A1(_0802_),
    .A2(_0804_));
 sg13g2_or3_1 _2257_ (.A(_0802_),
    .B(_0804_),
    .C(_0833_),
    .X(_0835_));
 sg13g2_and2_1 _2258_ (.A(_0834_),
    .B(_0835_),
    .X(_0836_));
 sg13g2_and2_1 _2259_ (.A(_0806_),
    .B(_0836_),
    .X(_0837_));
 sg13g2_xnor2_1 _2260_ (.Y(_0838_),
    .A(_0806_),
    .B(_0836_));
 sg13g2_and2_1 _2261_ (.A(_0774_),
    .B(_0809_),
    .X(_0839_));
 sg13g2_a21oi_1 _2262_ (.A1(_0777_),
    .A2(_0839_),
    .Y(_0840_),
    .B1(_0808_));
 sg13g2_a221oi_1 _2263_ (.B2(_0777_),
    .C1(_0838_),
    .B1(_0839_),
    .A1(_0771_),
    .Y(_0841_),
    .A2(_0807_));
 sg13g2_xor2_1 _2264_ (.B(_0840_),
    .A(_0838_),
    .X(_0842_));
 sg13g2_inv_1 _2265_ (.Y(_0843_),
    .A(_0842_));
 sg13g2_nor2_1 _2266_ (.A(_1246_),
    .B(_0842_),
    .Y(_0844_));
 sg13g2_nand2_1 _2267_ (.Y(_0845_),
    .A(_1246_),
    .B(_0842_));
 sg13g2_nor2b_1 _2268_ (.A(_0844_),
    .B_N(_0845_),
    .Y(_0846_));
 sg13g2_o21ai_1 _2269_ (.B1(_0814_),
    .Y(_0847_),
    .A1(_0788_),
    .A2(_0815_));
 sg13g2_a21oi_1 _2270_ (.A1(_0846_),
    .A2(_0847_),
    .Y(_0848_),
    .B1(_0747_));
 sg13g2_o21ai_1 _2271_ (.B1(_0848_),
    .Y(_0849_),
    .A1(_0846_),
    .A2(_0847_));
 sg13g2_nor2_1 _2272_ (.A(net133),
    .B(_1340_),
    .Y(_0850_));
 sg13g2_a22oi_1 _2273_ (.Y(_0851_),
    .B1(_0843_),
    .B2(net76),
    .A2(net708),
    .A1(net131));
 sg13g2_nand2_1 _2274_ (.Y(_0307_),
    .A(_0849_),
    .B(net709));
 sg13g2_nor2_1 _2275_ (.A(_0837_),
    .B(_0841_),
    .Y(_0852_));
 sg13g2_nand2_1 _2276_ (.Y(_0853_),
    .A(net18),
    .B(_0593_));
 sg13g2_xor2_1 _2277_ (.B(_0853_),
    .A(_0822_),
    .X(_0854_));
 sg13g2_o21ai_1 _2278_ (.B1(_0854_),
    .Y(_0855_),
    .A1(_0824_),
    .A2(_0826_));
 sg13g2_or3_1 _2279_ (.A(_0824_),
    .B(_0826_),
    .C(_0854_),
    .X(_0856_));
 sg13g2_nand2_1 _2280_ (.Y(_0857_),
    .A(_0855_),
    .B(_0856_));
 sg13g2_nand2_1 _2281_ (.Y(_0858_),
    .A(_0828_),
    .B(_0832_));
 sg13g2_a21oi_1 _2282_ (.A1(_0828_),
    .A2(_0832_),
    .Y(_0859_),
    .B1(_0857_));
 sg13g2_nand2b_1 _2283_ (.Y(_0860_),
    .B(_0858_),
    .A_N(_0857_));
 sg13g2_xor2_1 _2284_ (.B(_0858_),
    .A(_0857_),
    .X(_0861_));
 sg13g2_nor2_1 _2285_ (.A(_0834_),
    .B(_0861_),
    .Y(_0862_));
 sg13g2_nand2_1 _2286_ (.Y(_0863_),
    .A(_0834_),
    .B(_0861_));
 sg13g2_nor2b_1 _2287_ (.A(_0862_),
    .B_N(_0863_),
    .Y(_0864_));
 sg13g2_xnor2_1 _2288_ (.Y(_0865_),
    .A(_0852_),
    .B(_0864_));
 sg13g2_nand2_1 _2289_ (.Y(_0866_),
    .A(\mix_acc[5] ),
    .B(_0865_));
 sg13g2_xnor2_1 _2290_ (.Y(_0867_),
    .A(net728),
    .B(_0865_));
 sg13g2_a21oi_1 _2291_ (.A1(_0845_),
    .A2(_0847_),
    .Y(_0868_),
    .B1(_0844_));
 sg13g2_xnor2_1 _2292_ (.Y(_0869_),
    .A(_0867_),
    .B(_0868_));
 sg13g2_a22oi_1 _2293_ (.Y(_0870_),
    .B1(net76),
    .B2(_0865_),
    .A2(net728),
    .A1(net131));
 sg13g2_o21ai_1 _2294_ (.B1(_0870_),
    .Y(_0308_),
    .A1(_0747_),
    .A2(_0869_));
 sg13g2_or2_1 _2295_ (.X(_0871_),
    .B(_0862_),
    .A(_0837_));
 sg13g2_o21ai_1 _2296_ (.B1(_0863_),
    .Y(_0872_),
    .A1(_0841_),
    .A2(_0871_));
 sg13g2_nand2_1 _2297_ (.Y(_0873_),
    .A(net16),
    .B(_0593_));
 sg13g2_nor2b_1 _2298_ (.A(_0873_),
    .B_N(_0823_),
    .Y(_0874_));
 sg13g2_nand2_1 _2299_ (.Y(_0875_),
    .A(_0855_),
    .B(_0860_));
 sg13g2_xnor2_1 _2300_ (.Y(_0876_),
    .A(_0874_),
    .B(_0875_));
 sg13g2_xor2_1 _2301_ (.B(_0876_),
    .A(_0872_),
    .X(_0877_));
 sg13g2_xnor2_1 _2302_ (.Y(_0878_),
    .A(net712),
    .B(_0877_));
 sg13g2_inv_1 _2303_ (.Y(_0879_),
    .A(_0878_));
 sg13g2_o21ai_1 _2304_ (.B1(_0866_),
    .Y(_0880_),
    .A1(_0867_),
    .A2(_0868_));
 sg13g2_and2_1 _2305_ (.A(_0879_),
    .B(_0880_),
    .X(_0881_));
 sg13g2_nor2_1 _2306_ (.A(_0747_),
    .B(_0881_),
    .Y(_0882_));
 sg13g2_o21ai_1 _2307_ (.B1(_0882_),
    .Y(_0883_),
    .A1(_0879_),
    .A2(_0880_));
 sg13g2_a21oi_1 _2308_ (.A1(_1339_),
    .A2(_0877_),
    .Y(_0884_),
    .B1(net132));
 sg13g2_a22oi_1 _2309_ (.Y(_0309_),
    .B1(_0883_),
    .B2(_0884_),
    .A2(_1247_),
    .A1(net133));
 sg13g2_a21oi_1 _2310_ (.A1(_0823_),
    .A2(_0855_),
    .Y(_0885_),
    .B1(_0873_));
 sg13g2_a21oi_1 _2311_ (.A1(_0859_),
    .A2(_0874_),
    .Y(_0886_),
    .B1(_0885_));
 sg13g2_o21ai_1 _2312_ (.B1(_0886_),
    .Y(_0887_),
    .A1(_0872_),
    .A2(_0876_));
 sg13g2_xnor2_1 _2313_ (.Y(_0888_),
    .A(_1248_),
    .B(_0887_));
 sg13g2_a21o_1 _2314_ (.A2(_0877_),
    .A1(net712),
    .B1(_0881_),
    .X(_0889_));
 sg13g2_nand3_1 _2315_ (.B(_0880_),
    .C(_0888_),
    .A(_0879_),
    .Y(_0890_));
 sg13g2_and3_1 _2316_ (.X(_0891_),
    .A(net712),
    .B(_0877_),
    .C(_0888_));
 sg13g2_nor2_1 _2317_ (.A(_0747_),
    .B(_0891_),
    .Y(_0892_));
 sg13g2_and2_1 _2318_ (.A(_0890_),
    .B(_0892_),
    .X(_0893_));
 sg13g2_o21ai_1 _2319_ (.B1(_0893_),
    .Y(_0894_),
    .A1(_0888_),
    .A2(_0889_));
 sg13g2_a21oi_1 _2320_ (.A1(_1339_),
    .A2(_0887_),
    .Y(_0895_),
    .B1(net132));
 sg13g2_a22oi_1 _2321_ (.Y(_0310_),
    .B1(_0894_),
    .B2(_0895_),
    .A2(_1248_),
    .A1(net132));
 sg13g2_nand2_1 _2322_ (.Y(_0896_),
    .A(net132),
    .B(net311));
 sg13g2_a21oi_1 _2323_ (.A1(net369),
    .A2(_0887_),
    .Y(_0897_),
    .B1(_0891_));
 sg13g2_nand3_1 _2324_ (.B(_0890_),
    .C(_0897_),
    .A(_1249_),
    .Y(_0898_));
 sg13g2_a21oi_1 _2325_ (.A1(_0890_),
    .A2(net370),
    .Y(_0899_),
    .B1(_1249_));
 sg13g2_nand2_1 _2326_ (.Y(_0900_),
    .A(_0746_),
    .B(_0898_));
 sg13g2_o21ai_1 _2327_ (.B1(net312),
    .Y(_0311_),
    .A1(_0899_),
    .A2(_0900_));
 sg13g2_and3_1 _2328_ (.X(_0901_),
    .A(_1220_),
    .B(net318),
    .C(_0899_));
 sg13g2_a21oi_1 _2329_ (.A1(_1220_),
    .A2(net371),
    .Y(_0902_),
    .B1(net318));
 sg13g2_nand2_1 _2330_ (.Y(_0903_),
    .A(_1220_),
    .B(_1270_));
 sg13g2_nand3_1 _2331_ (.B(_1270_),
    .C(_1271_),
    .A(_1220_),
    .Y(_0904_));
 sg13g2_inv_1 _2332_ (.Y(_0905_),
    .A(net38));
 sg13g2_nor3_1 _2333_ (.A(_0901_),
    .B(_0902_),
    .C(_0905_),
    .Y(_0312_));
 sg13g2_nor2_1 _2334_ (.A(net372),
    .B(net113),
    .Y(_0906_));
 sg13g2_a21oi_1 _2335_ (.A1(_1245_),
    .A2(net113),
    .Y(_0313_),
    .B1(_0906_));
 sg13g2_mux2_1 _2336_ (.A0(net652),
    .A1(\mix_acc[3] ),
    .S(net113),
    .X(_0314_));
 sg13g2_nor2_1 _2337_ (.A(net392),
    .B(net113),
    .Y(_0907_));
 sg13g2_a21oi_1 _2338_ (.A1(_1246_),
    .A2(net113),
    .Y(_0315_),
    .B1(_0907_));
 sg13g2_nand2_1 _2339_ (.Y(_0908_),
    .A(net734),
    .B(net113));
 sg13g2_o21ai_1 _2340_ (.B1(_0908_),
    .Y(_0316_),
    .A1(_1254_),
    .A2(net113));
 sg13g2_nor2_1 _2341_ (.A(net335),
    .B(net113),
    .Y(_0909_));
 sg13g2_a21oi_1 _2342_ (.A1(_1247_),
    .A2(net114),
    .Y(_0317_),
    .B1(_0909_));
 sg13g2_nor2_1 _2343_ (.A(net548),
    .B(net114),
    .Y(_0910_));
 sg13g2_a21oi_1 _2344_ (.A1(_1248_),
    .A2(net114),
    .Y(_0318_),
    .B1(_0910_));
 sg13g2_nor2_1 _2345_ (.A(net538),
    .B(net114),
    .Y(_0911_));
 sg13g2_a21oi_1 _2346_ (.A1(_1249_),
    .A2(net114),
    .Y(_0319_),
    .B1(_0911_));
 sg13g2_nand2_1 _2347_ (.Y(_0912_),
    .A(net318),
    .B(net114));
 sg13g2_o21ai_1 _2348_ (.B1(_0912_),
    .Y(_0320_),
    .A1(_1250_),
    .A2(_1273_));
 sg13g2_nor2_1 _2349_ (.A(net621),
    .B(net89),
    .Y(_0913_));
 sg13g2_nand2_1 _2350_ (.Y(_0914_),
    .A(_1181_),
    .B(_1182_));
 sg13g2_nand3_1 _2351_ (.B(net36),
    .C(_0914_),
    .A(_1319_),
    .Y(_0915_));
 sg13g2_a21oi_1 _2352_ (.A1(net89),
    .A2(_0915_),
    .Y(_0321_),
    .B1(_0913_));
 sg13g2_nor2_1 _2353_ (.A(net403),
    .B(net87),
    .Y(_0916_));
 sg13g2_xor2_1 _2354_ (.B(_1319_),
    .A(_1318_),
    .X(_0917_));
 sg13g2_nand2_1 _2355_ (.Y(_0918_),
    .A(net36),
    .B(_0917_));
 sg13g2_a21oi_1 _2356_ (.A1(net87),
    .A2(_0918_),
    .Y(_0322_),
    .B1(_0916_));
 sg13g2_nor2_1 _2357_ (.A(net376),
    .B(net89),
    .Y(_0919_));
 sg13g2_xnor2_1 _2358_ (.Y(_0920_),
    .A(_1316_),
    .B(_1320_));
 sg13g2_nand2_1 _2359_ (.Y(_0921_),
    .A(net36),
    .B(_0920_));
 sg13g2_a21oi_1 _2360_ (.A1(net89),
    .A2(_0921_),
    .Y(_0323_),
    .B1(_0919_));
 sg13g2_nand2_1 _2361_ (.Y(_0922_),
    .A(_1321_),
    .B(_1322_));
 sg13g2_nand3_1 _2362_ (.B(net36),
    .C(_0922_),
    .A(_1323_),
    .Y(_0923_));
 sg13g2_nor2_1 _2363_ (.A(net354),
    .B(net89),
    .Y(_0924_));
 sg13g2_a21oi_1 _2364_ (.A1(net89),
    .A2(_0923_),
    .Y(_0324_),
    .B1(_0924_));
 sg13g2_nand2b_1 _2365_ (.Y(_0925_),
    .B(_1311_),
    .A_N(_1324_));
 sg13g2_nand3_1 _2366_ (.B(net36),
    .C(_0925_),
    .A(_1325_),
    .Y(_0926_));
 sg13g2_nor2_1 _2367_ (.A(net464),
    .B(net87),
    .Y(_0927_));
 sg13g2_a21oi_1 _2368_ (.A1(net87),
    .A2(_0926_),
    .Y(_0325_),
    .B1(_0927_));
 sg13g2_nand2_1 _2369_ (.Y(_0928_),
    .A(_1307_),
    .B(_1326_));
 sg13g2_nand3_1 _2370_ (.B(net36),
    .C(_0928_),
    .A(_1327_),
    .Y(_0929_));
 sg13g2_nor2_1 _2371_ (.A(net329),
    .B(net87),
    .Y(_0930_));
 sg13g2_a21oi_1 _2372_ (.A1(net87),
    .A2(_0929_),
    .Y(_0326_),
    .B1(_0930_));
 sg13g2_nor2_1 _2373_ (.A(net356),
    .B(net83),
    .Y(_0931_));
 sg13g2_nand2b_1 _2374_ (.Y(_0932_),
    .B(_1305_),
    .A_N(_1328_));
 sg13g2_nand3_1 _2375_ (.B(net36),
    .C(_0932_),
    .A(_1329_),
    .Y(_0933_));
 sg13g2_a21oi_1 _2376_ (.A1(net83),
    .A2(_0933_),
    .Y(_0327_),
    .B1(_0931_));
 sg13g2_a221oi_1 _2377_ (.B2(_1344_),
    .C1(\p_waveform[3] ),
    .B1(_1343_),
    .A1(_1330_),
    .Y(_0934_),
    .A2(_1331_));
 sg13g2_o21ai_1 _2378_ (.B1(_0934_),
    .Y(_0935_),
    .A1(_1330_),
    .A2(_1331_));
 sg13g2_nor2_1 _2379_ (.A(net327),
    .B(net83),
    .Y(_0936_));
 sg13g2_a21oi_1 _2380_ (.A1(net83),
    .A2(_0935_),
    .Y(_0328_),
    .B1(_0936_));
 sg13g2_nor2_1 _2381_ (.A(net466),
    .B(net83),
    .Y(_0937_));
 sg13g2_a21oi_1 _2382_ (.A1(_1353_),
    .A2(net82),
    .Y(_0329_),
    .B1(_0937_));
 sg13g2_nor2_1 _2383_ (.A(net346),
    .B(net82),
    .Y(_0938_));
 sg13g2_a21oi_1 _2384_ (.A1(_1350_),
    .A2(net82),
    .Y(_0330_),
    .B1(_0938_));
 sg13g2_nor2_1 _2385_ (.A(net400),
    .B(net82),
    .Y(_0939_));
 sg13g2_a21oi_1 _2386_ (.A1(_1357_),
    .A2(net82),
    .Y(_0331_),
    .B1(_0939_));
 sg13g2_nor2_1 _2387_ (.A(net247),
    .B(net78),
    .Y(_0940_));
 sg13g2_a21oi_1 _2388_ (.A1(_1360_),
    .A2(net78),
    .Y(_0332_),
    .B1(_0940_));
 sg13g2_nor2_1 _2389_ (.A(net394),
    .B(net77),
    .Y(_0941_));
 sg13g2_a21oi_1 _2390_ (.A1(_1364_),
    .A2(net77),
    .Y(_0333_),
    .B1(_0941_));
 sg13g2_nor2_1 _2391_ (.A(net337),
    .B(net77),
    .Y(_0942_));
 sg13g2_a21oi_1 _2392_ (.A1(_1370_),
    .A2(net77),
    .Y(_0334_),
    .B1(_0942_));
 sg13g2_nor2_1 _2393_ (.A(net382),
    .B(net78),
    .Y(_0943_));
 sg13g2_a21oi_1 _2394_ (.A1(_1373_),
    .A2(net78),
    .Y(_0335_),
    .B1(_0943_));
 sg13g2_nor2_1 _2395_ (.A(net705),
    .B(net78),
    .Y(_0944_));
 sg13g2_a21oi_1 _2396_ (.A1(_1347_),
    .A2(net78),
    .Y(_0336_),
    .B1(_0944_));
 sg13g2_nor2_1 _2397_ (.A(net333),
    .B(net109),
    .Y(_0945_));
 sg13g2_a21oi_1 _2398_ (.A1(net109),
    .A2(_0915_),
    .Y(_0337_),
    .B1(_0945_));
 sg13g2_nor2_1 _2399_ (.A(net386),
    .B(net108),
    .Y(_0946_));
 sg13g2_a21oi_1 _2400_ (.A1(net108),
    .A2(_0918_),
    .Y(_0338_),
    .B1(_0946_));
 sg13g2_nor2_1 _2401_ (.A(net384),
    .B(net108),
    .Y(_0947_));
 sg13g2_a21oi_1 _2402_ (.A1(net108),
    .A2(_0921_),
    .Y(_0339_),
    .B1(_0947_));
 sg13g2_nor2_1 _2403_ (.A(net414),
    .B(net109),
    .Y(_0948_));
 sg13g2_a21oi_1 _2404_ (.A1(net109),
    .A2(_0923_),
    .Y(_0340_),
    .B1(_0948_));
 sg13g2_nor2_1 _2405_ (.A(net444),
    .B(net108),
    .Y(_0949_));
 sg13g2_a21oi_1 _2406_ (.A1(net108),
    .A2(_0926_),
    .Y(_0341_),
    .B1(_0949_));
 sg13g2_nor2_1 _2407_ (.A(net388),
    .B(net108),
    .Y(_0950_));
 sg13g2_a21oi_1 _2408_ (.A1(net108),
    .A2(_0929_),
    .Y(_0342_),
    .B1(_0950_));
 sg13g2_nor2_1 _2409_ (.A(net344),
    .B(net110),
    .Y(_0951_));
 sg13g2_a21oi_1 _2410_ (.A1(net110),
    .A2(_0933_),
    .Y(_0343_),
    .B1(_0951_));
 sg13g2_nor2_1 _2411_ (.A(net374),
    .B(net110),
    .Y(_0952_));
 sg13g2_a21oi_1 _2412_ (.A1(net110),
    .A2(_0935_),
    .Y(_0344_),
    .B1(_0952_));
 sg13g2_nor2_1 _2413_ (.A(net442),
    .B(net110),
    .Y(_0953_));
 sg13g2_a21oi_1 _2414_ (.A1(_1353_),
    .A2(net110),
    .Y(_0345_),
    .B1(_0953_));
 sg13g2_nor2_1 _2415_ (.A(net367),
    .B(net103),
    .Y(_0954_));
 sg13g2_a21oi_1 _2416_ (.A1(_1350_),
    .A2(net103),
    .Y(_0346_),
    .B1(_0954_));
 sg13g2_nor2_1 _2417_ (.A(net350),
    .B(net103),
    .Y(_0955_));
 sg13g2_a21oi_1 _2418_ (.A1(_1357_),
    .A2(net103),
    .Y(_0347_),
    .B1(_0955_));
 sg13g2_nor2_1 _2419_ (.A(net522),
    .B(net103),
    .Y(_0956_));
 sg13g2_a21oi_1 _2420_ (.A1(_1360_),
    .A2(net103),
    .Y(_0348_),
    .B1(_0956_));
 sg13g2_nor2_1 _2421_ (.A(net412),
    .B(net104),
    .Y(_0957_));
 sg13g2_a21oi_1 _2422_ (.A1(_1364_),
    .A2(net104),
    .Y(_0040_),
    .B1(_0957_));
 sg13g2_nor2_1 _2423_ (.A(net410),
    .B(net103),
    .Y(_0958_));
 sg13g2_a21oi_1 _2424_ (.A1(_1370_),
    .A2(net103),
    .Y(_0041_),
    .B1(_0958_));
 sg13g2_nor2_1 _2425_ (.A(net390),
    .B(net104),
    .Y(_0959_));
 sg13g2_a21oi_1 _2426_ (.A1(_1373_),
    .A2(net104),
    .Y(_0042_),
    .B1(_0959_));
 sg13g2_nor2_1 _2427_ (.A(net675),
    .B(net104),
    .Y(_0960_));
 sg13g2_a21oi_1 _2428_ (.A1(_1347_),
    .A2(net104),
    .Y(_0043_),
    .B1(_0960_));
 sg13g2_nand2_1 _2429_ (.Y(_0961_),
    .A(net302),
    .B(net100));
 sg13g2_o21ai_1 _2430_ (.B1(net303),
    .Y(_0044_),
    .A1(net100),
    .A2(_0915_));
 sg13g2_nand2_1 _2431_ (.Y(_0962_),
    .A(net287),
    .B(net99));
 sg13g2_o21ai_1 _2432_ (.B1(net288),
    .Y(_0045_),
    .A1(net99),
    .A2(_0918_));
 sg13g2_nand2_1 _2433_ (.Y(_0963_),
    .A(net275),
    .B(net99));
 sg13g2_o21ai_1 _2434_ (.B1(net276),
    .Y(_0046_),
    .A1(net99),
    .A2(_0921_));
 sg13g2_nand2_1 _2435_ (.Y(_0964_),
    .A(net293),
    .B(net100));
 sg13g2_o21ai_1 _2436_ (.B1(net294),
    .Y(_0047_),
    .A1(net100),
    .A2(_0923_));
 sg13g2_nand2_1 _2437_ (.Y(_0965_),
    .A(net284),
    .B(net99));
 sg13g2_o21ai_1 _2438_ (.B1(net285),
    .Y(_0048_),
    .A1(net99),
    .A2(_0926_));
 sg13g2_nand2_1 _2439_ (.Y(_0966_),
    .A(net263),
    .B(net99));
 sg13g2_o21ai_1 _2440_ (.B1(net264),
    .Y(_0049_),
    .A1(net99),
    .A2(_0929_));
 sg13g2_nand2_1 _2441_ (.Y(_0967_),
    .A(net272),
    .B(net101));
 sg13g2_o21ai_1 _2442_ (.B1(net273),
    .Y(_0050_),
    .A1(net101),
    .A2(_0933_));
 sg13g2_nand2_1 _2443_ (.Y(_0968_),
    .A(net308),
    .B(net101));
 sg13g2_o21ai_1 _2444_ (.B1(net309),
    .Y(_0051_),
    .A1(net101),
    .A2(_0935_));
 sg13g2_nand2_1 _2445_ (.Y(_0969_),
    .A(net281),
    .B(net101));
 sg13g2_o21ai_1 _2446_ (.B1(net282),
    .Y(_0052_),
    .A1(_1353_),
    .A2(net101));
 sg13g2_nand2_1 _2447_ (.Y(_0970_),
    .A(net269),
    .B(net95));
 sg13g2_o21ai_1 _2448_ (.B1(net270),
    .Y(_0053_),
    .A1(_1350_),
    .A2(net95));
 sg13g2_nand2_1 _2449_ (.Y(_0971_),
    .A(net320),
    .B(net95));
 sg13g2_o21ai_1 _2450_ (.B1(_0971_),
    .Y(_0054_),
    .A1(_1357_),
    .A2(net95));
 sg13g2_nand2_1 _2451_ (.Y(_0972_),
    .A(net290),
    .B(net95));
 sg13g2_o21ai_1 _2452_ (.B1(net291),
    .Y(_0055_),
    .A1(_1360_),
    .A2(net95));
 sg13g2_nand2_1 _2453_ (.Y(_0973_),
    .A(net325),
    .B(net96));
 sg13g2_o21ai_1 _2454_ (.B1(_0973_),
    .Y(_0056_),
    .A1(_1364_),
    .A2(net96));
 sg13g2_nand2_1 _2455_ (.Y(_0974_),
    .A(net299),
    .B(net95));
 sg13g2_o21ai_1 _2456_ (.B1(net300),
    .Y(_0057_),
    .A1(_1370_),
    .A2(net95));
 sg13g2_nand2_1 _2457_ (.Y(_0975_),
    .A(net322),
    .B(net96));
 sg13g2_o21ai_1 _2458_ (.B1(_0975_),
    .Y(_0058_),
    .A1(_1373_),
    .A2(net96));
 sg13g2_nand2_1 _2459_ (.Y(_0976_),
    .A(net348),
    .B(net96));
 sg13g2_o21ai_1 _2460_ (.B1(_0976_),
    .Y(_0059_),
    .A1(_1347_),
    .A2(net96));
 sg13g2_mux2_1 _2461_ (.A0(net620),
    .A1(net17),
    .S(net75),
    .X(_0060_));
 sg13g2_mux2_1 _2462_ (.A0(net625),
    .A1(net29),
    .S(net75),
    .X(_0061_));
 sg13g2_mux2_1 _2463_ (.A0(net598),
    .A1(net25),
    .S(net80),
    .X(_0062_));
 sg13g2_mux2_1 _2464_ (.A0(net590),
    .A1(net20),
    .S(net75),
    .X(_0063_));
 sg13g2_mux2_1 _2465_ (.A0(net434),
    .A1(net22),
    .S(net75),
    .X(_0064_));
 sg13g2_mux2_1 _2466_ (.A0(net569),
    .A1(net27),
    .S(net80),
    .X(_0065_));
 sg13g2_mux2_1 _2467_ (.A0(net458),
    .A1(net18),
    .S(net79),
    .X(_0066_));
 sg13g2_mux2_1 _2468_ (.A0(net537),
    .A1(net16),
    .S(net80),
    .X(_0067_));
 sg13g2_mux2_1 _2469_ (.A0(net588),
    .A1(_0530_),
    .S(net105),
    .X(_0068_));
 sg13g2_mux2_1 _2470_ (.A0(net602),
    .A1(_0546_),
    .S(net105),
    .X(_0069_));
 sg13g2_mux2_1 _2471_ (.A0(net567),
    .A1(net25),
    .S(net105),
    .X(_0070_));
 sg13g2_mux2_1 _2472_ (.A0(net503),
    .A1(net20),
    .S(net105),
    .X(_0071_));
 sg13g2_mux2_1 _2473_ (.A0(net468),
    .A1(net22),
    .S(net105),
    .X(_0072_));
 sg13g2_mux2_1 _2474_ (.A0(net543),
    .A1(net27),
    .S(net105),
    .X(_0073_));
 sg13g2_mux2_1 _2475_ (.A0(net424),
    .A1(_0502_),
    .S(net105),
    .X(_0074_));
 sg13g2_mux2_1 _2476_ (.A0(net550),
    .A1(net16),
    .S(net105),
    .X(_0075_));
 sg13g2_mux2_1 _2477_ (.A0(_0530_),
    .A1(net447),
    .S(net97),
    .X(_0076_));
 sg13g2_mux2_1 _2478_ (.A0(_0546_),
    .A1(net574),
    .S(net97),
    .X(_0077_));
 sg13g2_mux2_1 _2479_ (.A0(net25),
    .A1(net420),
    .S(net97),
    .X(_0078_));
 sg13g2_mux2_1 _2480_ (.A0(net20),
    .A1(net427),
    .S(net97),
    .X(_0079_));
 sg13g2_mux2_1 _2481_ (.A0(net22),
    .A1(net408),
    .S(net97),
    .X(_0080_));
 sg13g2_mux2_1 _2482_ (.A0(net27),
    .A1(net409),
    .S(net97),
    .X(_0081_));
 sg13g2_mux2_1 _2483_ (.A0(_0502_),
    .A1(net647),
    .S(net97),
    .X(_0082_));
 sg13g2_mux2_1 _2484_ (.A0(_0578_),
    .A1(net525),
    .S(net97),
    .X(_0083_));
 sg13g2_a21oi_1 _2485_ (.A1(cur_gate),
    .A2(_0396_),
    .Y(_0977_),
    .B1(\p_ast[1] ));
 sg13g2_a21oi_1 _2486_ (.A1(cur_gate),
    .A2(_0429_),
    .Y(_0978_),
    .B1(_0977_));
 sg13g2_nor2_1 _2487_ (.A(_0392_),
    .B(_0978_),
    .Y(_0979_));
 sg13g2_and2_1 _2488_ (.A(_1385_),
    .B(_0392_),
    .X(_0980_));
 sg13g2_nor4_1 _2489_ (.A(net135),
    .B(_0410_),
    .C(_0979_),
    .D(_0980_),
    .Y(_0981_));
 sg13g2_a21oi_1 _2490_ (.A1(\p_ast[0] ),
    .A2(_1395_),
    .Y(_0982_),
    .B1(_1385_));
 sg13g2_a21oi_1 _2491_ (.A1(net135),
    .A2(_0982_),
    .Y(_0983_),
    .B1(_0981_));
 sg13g2_mux2_1 _2492_ (.A0(net594),
    .A1(_0983_),
    .S(net79),
    .X(_0084_));
 sg13g2_nor2_1 _2493_ (.A(net507),
    .B(net79),
    .Y(_0984_));
 sg13g2_nor2_1 _2494_ (.A(_0394_),
    .B(_0977_),
    .Y(_0985_));
 sg13g2_a21oi_1 _2495_ (.A1(\p_ast[1] ),
    .A2(_1396_),
    .Y(_0986_),
    .B1(_0985_));
 sg13g2_a21oi_1 _2496_ (.A1(net79),
    .A2(_0986_),
    .Y(_0085_),
    .B1(_0984_));
 sg13g2_mux2_1 _2497_ (.A0(net531),
    .A1(_0983_),
    .S(net106),
    .X(_0086_));
 sg13g2_nor2_1 _2498_ (.A(net540),
    .B(net106),
    .Y(_0987_));
 sg13g2_a21oi_1 _2499_ (.A1(net106),
    .A2(_0986_),
    .Y(_0087_),
    .B1(_0987_));
 sg13g2_mux2_1 _2500_ (.A0(_0983_),
    .A1(net616),
    .S(net98),
    .X(_0088_));
 sg13g2_nand2_1 _2501_ (.Y(_0988_),
    .A(net266),
    .B(net98));
 sg13g2_o21ai_1 _2502_ (.B1(net267),
    .Y(_0089_),
    .A1(net98),
    .A2(_0986_));
 sg13g2_nor2_1 _2503_ (.A(net381),
    .B(net85),
    .Y(_0989_));
 sg13g2_a21oi_1 _2504_ (.A1(_1189_),
    .A2(net85),
    .Y(_0090_),
    .B1(_0989_));
 sg13g2_nor2_1 _2505_ (.A(net475),
    .B(net111),
    .Y(_0990_));
 sg13g2_a21oi_1 _2506_ (.A1(_1189_),
    .A2(net111),
    .Y(_0091_),
    .B1(_0990_));
 sg13g2_nand2_1 _2507_ (.Y(_0991_),
    .A(net324),
    .B(net102));
 sg13g2_o21ai_1 _2508_ (.B1(_0991_),
    .Y(_0092_),
    .A1(_1189_),
    .A2(net102));
 sg13g2_o21ai_1 _2509_ (.B1(_0438_),
    .Y(_0992_),
    .A1(net147),
    .A2(_0394_));
 sg13g2_mux2_1 _2510_ (.A0(net586),
    .A1(_0992_),
    .S(net80),
    .X(_0093_));
 sg13g2_mux2_1 _2511_ (.A0(net560),
    .A1(_0992_),
    .S(net106),
    .X(_0094_));
 sg13g2_mux2_1 _2512_ (.A0(_0992_),
    .A1(net500),
    .S(net98),
    .X(_0095_));
 sg13g2_nand2_1 _2513_ (.Y(_0993_),
    .A(\acc[0][15] ),
    .B(net104));
 sg13g2_o21ai_1 _2514_ (.B1(_0993_),
    .Y(_0096_),
    .A1(_1225_),
    .A2(net104));
 sg13g2_mux2_1 _2515_ (.A0(\acc[1][15] ),
    .A1(net529),
    .S(net96),
    .X(_0097_));
 sg13g2_nor2_1 _2516_ (.A(net501),
    .B(net76),
    .Y(_0994_));
 sg13g2_a21oi_1 _2517_ (.A1(_1185_),
    .A2(net76),
    .Y(_0098_),
    .B1(_0994_));
 sg13g2_nor2b_1 _2518_ (.A(net481),
    .B_N(net247),
    .Y(_0995_));
 sg13g2_xor2_1 _2519_ (.B(_0038_),
    .A(_0039_),
    .X(_0996_));
 sg13g2_nor2_1 _2520_ (.A(net339),
    .B(net116),
    .Y(_0997_));
 sg13g2_a21oi_1 _2521_ (.A1(net116),
    .A2(_0996_),
    .Y(_0099_),
    .B1(net340));
 sg13g2_mux2_1 _2522_ (.A0(net405),
    .A1(net339),
    .S(net116),
    .X(_0100_));
 sg13g2_mux2_1 _2523_ (.A0(net398),
    .A1(net405),
    .S(net115),
    .X(_0101_));
 sg13g2_mux2_1 _2524_ (.A0(_0028_),
    .A1(net398),
    .S(net115),
    .X(_0102_));
 sg13g2_mux2_1 _2525_ (.A0(net570),
    .A1(_0028_),
    .S(net115),
    .X(_0103_));
 sg13g2_mux2_1 _2526_ (.A0(net639),
    .A1(net570),
    .S(net115),
    .X(_0104_));
 sg13g2_mux2_1 _2527_ (.A0(net418),
    .A1(_0030_),
    .S(net115),
    .X(_0105_));
 sg13g2_mux2_1 _2528_ (.A0(net430),
    .A1(net418),
    .S(net115),
    .X(_0106_));
 sg13g2_mux2_1 _2529_ (.A0(net679),
    .A1(net430),
    .S(net115),
    .X(_0107_));
 sg13g2_mux2_1 _2530_ (.A0(net680),
    .A1(net679),
    .S(net115),
    .X(_0108_));
 sg13g2_mux2_1 _2531_ (.A0(net666),
    .A1(_0034_),
    .S(net116),
    .X(_0109_));
 sg13g2_mux2_1 _2532_ (.A0(net674),
    .A1(net666),
    .S(net116),
    .X(_0110_));
 sg13g2_mux2_1 _2533_ (.A0(net662),
    .A1(_0036_),
    .S(net116),
    .X(_0111_));
 sg13g2_mux2_1 _2534_ (.A0(net664),
    .A1(net662),
    .S(net116),
    .X(_0112_));
 sg13g2_mux2_1 _2535_ (.A0(net702),
    .A1(net664),
    .S(net116),
    .X(_0113_));
 sg13g2_a21oi_1 _2536_ (.A1(net621),
    .A2(net124),
    .Y(_0998_),
    .B1(net65));
 sg13g2_a22oi_1 _2537_ (.Y(_0999_),
    .B1(net43),
    .B2(net302),
    .A2(net88),
    .A1(net333));
 sg13g2_a22oi_1 _2538_ (.Y(_0114_),
    .B1(_0998_),
    .B2(_0999_),
    .A2(net65),
    .A1(_1181_));
 sg13g2_a21oi_1 _2539_ (.A1(net403),
    .A2(net124),
    .Y(_1000_),
    .B1(net64));
 sg13g2_a22oi_1 _2540_ (.Y(_1001_),
    .B1(net43),
    .B2(net287),
    .A2(net87),
    .A1(net386));
 sg13g2_a22oi_1 _2541_ (.Y(_0115_),
    .B1(_1000_),
    .B2(_1001_),
    .A2(net64),
    .A1(_1179_));
 sg13g2_a21oi_1 _2542_ (.A1(net376),
    .A2(net124),
    .Y(_1002_),
    .B1(net63));
 sg13g2_a22oi_1 _2543_ (.Y(_1003_),
    .B1(net43),
    .B2(net275),
    .A2(net89),
    .A1(net384));
 sg13g2_a22oi_1 _2544_ (.Y(_0116_),
    .B1(_1002_),
    .B2(_1003_),
    .A2(net63),
    .A1(_1177_));
 sg13g2_a21oi_1 _2545_ (.A1(net354),
    .A2(net125),
    .Y(_1004_),
    .B1(net63));
 sg13g2_a22oi_1 _2546_ (.Y(_1005_),
    .B1(net43),
    .B2(net293),
    .A2(net89),
    .A1(net414));
 sg13g2_a22oi_1 _2547_ (.Y(_0117_),
    .B1(_1004_),
    .B2(_1005_),
    .A2(net63),
    .A1(_1175_));
 sg13g2_a21oi_1 _2548_ (.A1(\acc[0][4] ),
    .A2(net124),
    .Y(_1006_),
    .B1(net64));
 sg13g2_a22oi_1 _2549_ (.Y(_1007_),
    .B1(net43),
    .B2(net284),
    .A2(net88),
    .A1(net444));
 sg13g2_a22oi_1 _2550_ (.Y(_0118_),
    .B1(_1006_),
    .B2(_1007_),
    .A2(net64),
    .A1(_1173_));
 sg13g2_a21oi_1 _2551_ (.A1(net329),
    .A2(net124),
    .Y(_1008_),
    .B1(net64));
 sg13g2_a22oi_1 _2552_ (.Y(_1009_),
    .B1(net43),
    .B2(net263),
    .A2(net87),
    .A1(net388));
 sg13g2_a22oi_1 _2553_ (.Y(_0119_),
    .B1(_1008_),
    .B2(_1009_),
    .A2(net64),
    .A1(_1171_));
 sg13g2_a21oi_1 _2554_ (.A1(net356),
    .A2(net120),
    .Y(_1010_),
    .B1(net61));
 sg13g2_a22oi_1 _2555_ (.Y(_1011_),
    .B1(net41),
    .B2(net272),
    .A2(net83),
    .A1(net344));
 sg13g2_a22oi_1 _2556_ (.Y(_0120_),
    .B1(_1010_),
    .B2(_1011_),
    .A2(net61),
    .A1(_1169_));
 sg13g2_a21oi_1 _2557_ (.A1(net327),
    .A2(net121),
    .Y(_1012_),
    .B1(net61));
 sg13g2_a22oi_1 _2558_ (.Y(_1013_),
    .B1(net41),
    .B2(net308),
    .A2(net83),
    .A1(net374));
 sg13g2_a22oi_1 _2559_ (.Y(_0121_),
    .B1(_1012_),
    .B2(_1013_),
    .A2(net61),
    .A1(_1167_));
 sg13g2_a21oi_1 _2560_ (.A1(net466),
    .A2(net121),
    .Y(_1014_),
    .B1(net61));
 sg13g2_a22oi_1 _2561_ (.Y(_1015_),
    .B1(net41),
    .B2(net281),
    .A2(net82),
    .A1(net442));
 sg13g2_a22oi_1 _2562_ (.Y(_0122_),
    .B1(_1014_),
    .B2(_1015_),
    .A2(net61),
    .A1(_1166_));
 sg13g2_a21oi_1 _2563_ (.A1(net346),
    .A2(net120),
    .Y(_1016_),
    .B1(net50));
 sg13g2_a22oi_1 _2564_ (.Y(_1017_),
    .B1(net37),
    .B2(net269),
    .A2(net82),
    .A1(net367));
 sg13g2_a22oi_1 _2565_ (.Y(_0123_),
    .B1(_1016_),
    .B2(_1017_),
    .A2(net50),
    .A1(_1165_));
 sg13g2_a21oi_1 _2566_ (.A1(net400),
    .A2(net120),
    .Y(_1018_),
    .B1(net50));
 sg13g2_a22oi_1 _2567_ (.Y(_1019_),
    .B1(net37),
    .B2(net320),
    .A2(net82),
    .A1(net350));
 sg13g2_a22oi_1 _2568_ (.Y(_0124_),
    .B1(_1018_),
    .B2(_1019_),
    .A2(net50),
    .A1(_1164_));
 sg13g2_a21oi_1 _2569_ (.A1(net247),
    .A2(net117),
    .Y(_1020_),
    .B1(net50));
 sg13g2_a22oi_1 _2570_ (.Y(_1021_),
    .B1(net37),
    .B2(net290),
    .A2(net77),
    .A1(net522));
 sg13g2_a22oi_1 _2571_ (.Y(_0125_),
    .B1(_1020_),
    .B2(_1021_),
    .A2(net50),
    .A1(_1163_));
 sg13g2_a21oi_1 _2572_ (.A1(net394),
    .A2(net117),
    .Y(_1022_),
    .B1(net51));
 sg13g2_a22oi_1 _2573_ (.Y(_1023_),
    .B1(net37),
    .B2(net325),
    .A2(net77),
    .A1(net412));
 sg13g2_a22oi_1 _2574_ (.Y(_0126_),
    .B1(_1022_),
    .B2(_1023_),
    .A2(net51),
    .A1(_1162_));
 sg13g2_a21oi_1 _2575_ (.A1(net337),
    .A2(net117),
    .Y(_1024_),
    .B1(net50));
 sg13g2_a22oi_1 _2576_ (.Y(_1025_),
    .B1(net37),
    .B2(net299),
    .A2(net77),
    .A1(net410));
 sg13g2_a22oi_1 _2577_ (.Y(_0127_),
    .B1(_1024_),
    .B2(_1025_),
    .A2(net50),
    .A1(_1161_));
 sg13g2_a21oi_1 _2578_ (.A1(net382),
    .A2(net117),
    .Y(_1026_),
    .B1(net55));
 sg13g2_a22oi_1 _2579_ (.Y(_1027_),
    .B1(net38),
    .B2(net322),
    .A2(net78),
    .A1(net390));
 sg13g2_a22oi_1 _2580_ (.Y(_0128_),
    .B1(_1026_),
    .B2(_1027_),
    .A2(net55),
    .A1(_1183_));
 sg13g2_a21oi_1 _2581_ (.A1(\acc[0][15] ),
    .A2(net117),
    .Y(_1028_),
    .B1(net55));
 sg13g2_a22oi_1 _2582_ (.Y(_1029_),
    .B1(net38),
    .B2(net348),
    .A2(net78),
    .A1(\acc[1][15] ));
 sg13g2_a22oi_1 _2583_ (.Y(_0129_),
    .B1(_1028_),
    .B2(_1029_),
    .A2(net55),
    .A1(_1184_));
 sg13g2_a21oi_1 _2584_ (.A1(\freq[0][0] ),
    .A2(net126),
    .Y(_1030_),
    .B1(net65));
 sg13g2_a22oi_1 _2585_ (.Y(_1031_),
    .B1(net47),
    .B2(\freq[2][0] ),
    .A2(net91),
    .A1(\freq[1][0] ));
 sg13g2_a22oi_1 _2586_ (.Y(_0130_),
    .B1(_1030_),
    .B2(_1031_),
    .A2(net65),
    .A1(_1182_));
 sg13g2_a21oi_1 _2587_ (.A1(net509),
    .A2(net124),
    .Y(_1032_),
    .B1(net66));
 sg13g2_a22oi_1 _2588_ (.Y(_1033_),
    .B1(net43),
    .B2(net470),
    .A2(net90),
    .A1(net478));
 sg13g2_a22oi_1 _2589_ (.Y(_0131_),
    .B1(_1032_),
    .B2(_1033_),
    .A2(net66),
    .A1(_1180_));
 sg13g2_a21oi_1 _2590_ (.A1(net482),
    .A2(net125),
    .Y(_1034_),
    .B1(net63));
 sg13g2_a22oi_1 _2591_ (.Y(_1035_),
    .B1(net43),
    .B2(net579),
    .A2(net90),
    .A1(net545));
 sg13g2_a22oi_1 _2592_ (.Y(_0132_),
    .B1(_1034_),
    .B2(_1035_),
    .A2(net63),
    .A1(_1178_));
 sg13g2_a21oi_1 _2593_ (.A1(net561),
    .A2(net125),
    .Y(_1036_),
    .B1(net63));
 sg13g2_a22oi_1 _2594_ (.Y(_1037_),
    .B1(net44),
    .B2(net457),
    .A2(net90),
    .A1(net510));
 sg13g2_a22oi_1 _2595_ (.Y(_0133_),
    .B1(_1036_),
    .B2(_1037_),
    .A2(net63),
    .A1(_1176_));
 sg13g2_a21oi_1 _2596_ (.A1(net607),
    .A2(net125),
    .Y(_1038_),
    .B1(net65));
 sg13g2_a22oi_1 _2597_ (.Y(_1039_),
    .B1(net44),
    .B2(net619),
    .A2(net90),
    .A1(net581));
 sg13g2_a22oi_1 _2598_ (.Y(_0134_),
    .B1(_1038_),
    .B2(_1039_),
    .A2(net65),
    .A1(_1174_));
 sg13g2_a21oi_1 _2599_ (.A1(net554),
    .A2(net126),
    .Y(_1040_),
    .B1(net70));
 sg13g2_a22oi_1 _2600_ (.Y(_1041_),
    .B1(net47),
    .B2(net528),
    .A2(net92),
    .A1(net455));
 sg13g2_a22oi_1 _2601_ (.Y(_0135_),
    .B1(_1040_),
    .B2(_1041_),
    .A2(net70),
    .A1(_1172_));
 sg13g2_a21oi_1 _2602_ (.A1(\freq[0][6] ),
    .A2(net124),
    .Y(_1042_),
    .B1(net64));
 sg13g2_a22oi_1 _2603_ (.Y(_1043_),
    .B1(net44),
    .B2(\freq[2][6] ),
    .A2(net88),
    .A1(\freq[1][6] ));
 sg13g2_a22oi_1 _2604_ (.Y(_0136_),
    .B1(_1042_),
    .B2(_1043_),
    .A2(net64),
    .A1(_1170_));
 sg13g2_a21oi_1 _2605_ (.A1(net576),
    .A2(net125),
    .Y(_1044_),
    .B1(net66));
 sg13g2_a22oi_1 _2606_ (.Y(_1045_),
    .B1(net44),
    .B2(net557),
    .A2(net90),
    .A1(net580));
 sg13g2_a22oi_1 _2607_ (.Y(_0137_),
    .B1(_1044_),
    .B2(_1045_),
    .A2(net66),
    .A1(_1168_));
 sg13g2_a21oi_1 _2608_ (.A1(net552),
    .A2(net122),
    .Y(_1046_),
    .B1(net58));
 sg13g2_a22oi_1 _2609_ (.Y(_1047_),
    .B1(net39),
    .B2(net593),
    .A2(net85),
    .A1(net553));
 sg13g2_a22oi_1 _2610_ (.Y(_0138_),
    .B1(_1046_),
    .B2(_1047_),
    .A2(net58),
    .A1(_1189_));
 sg13g2_a21oi_1 _2611_ (.A1(\waveform[0][1] ),
    .A2(net121),
    .Y(_1048_),
    .B1(net62));
 sg13g2_a22oi_1 _2612_ (.Y(_1049_),
    .B1(net41),
    .B2(\waveform[2][1] ),
    .A2(net83),
    .A1(\waveform[1][1] ));
 sg13g2_a22oi_1 _2613_ (.Y(_0139_),
    .B1(_1048_),
    .B2(_1049_),
    .A2(net62),
    .A1(_1187_));
 sg13g2_a21oi_1 _2614_ (.A1(\waveform[0][2] ),
    .A2(net120),
    .Y(_1050_),
    .B1(net51));
 sg13g2_a22oi_1 _2615_ (.Y(_1051_),
    .B1(net37),
    .B2(\waveform[2][2] ),
    .A2(net84),
    .A1(\waveform[1][2] ));
 sg13g2_a22oi_1 _2616_ (.Y(_0140_),
    .B1(_1050_),
    .B2(_1051_),
    .A2(net51),
    .A1(_1230_));
 sg13g2_a21oi_1 _2617_ (.A1(\waveform[0][3] ),
    .A2(net121),
    .Y(_1052_),
    .B1(net61));
 sg13g2_a22oi_1 _2618_ (.Y(_1053_),
    .B1(net41),
    .B2(\waveform[2][3] ),
    .A2(net84),
    .A1(\waveform[1][3] ));
 sg13g2_a22oi_1 _2619_ (.Y(_0141_),
    .B1(_1052_),
    .B2(_1053_),
    .A2(net61),
    .A1(_1160_));
 sg13g2_a21oi_1 _2620_ (.A1(net627),
    .A2(net117),
    .Y(_1054_),
    .B1(net52));
 sg13g2_a22oi_1 _2621_ (.Y(_1055_),
    .B1(net37),
    .B2(net536),
    .A2(net77),
    .A1(net613));
 sg13g2_a22oi_1 _2622_ (.Y(_0142_),
    .B1(_1054_),
    .B2(_1055_),
    .A2(net52),
    .A1(_1231_));
 sg13g2_a21oi_1 _2623_ (.A1(net425),
    .A2(net117),
    .Y(_1056_),
    .B1(net52));
 sg13g2_a22oi_1 _2624_ (.Y(_1057_),
    .B1(net37),
    .B2(net556),
    .A2(net81),
    .A1(net502));
 sg13g2_a22oi_1 _2625_ (.Y(_0143_),
    .B1(_1056_),
    .B2(_1057_),
    .A2(net52),
    .A1(_1232_));
 sg13g2_a21oi_1 _2626_ (.A1(net533),
    .A2(net118),
    .Y(_1058_),
    .B1(net58));
 sg13g2_a22oi_1 _2627_ (.Y(_1059_),
    .B1(net40),
    .B2(net518),
    .A2(net79),
    .A1(net631));
 sg13g2_a22oi_1 _2628_ (.Y(_0144_),
    .B1(_1058_),
    .B2(_1059_),
    .A2(net58),
    .A1(_1241_));
 sg13g2_a21oi_1 _2629_ (.A1(net517),
    .A2(net117),
    .Y(_1060_),
    .B1(net52));
 sg13g2_a22oi_1 _2630_ (.Y(_1061_),
    .B1(net38),
    .B2(net597),
    .A2(net79),
    .A1(net453));
 sg13g2_a22oi_1 _2631_ (.Y(_0145_),
    .B1(_1060_),
    .B2(_1061_),
    .A2(net52),
    .A1(_1242_));
 sg13g2_a21oi_1 _2632_ (.A1(\pw_reg[0][0] ),
    .A2(net122),
    .Y(_1062_),
    .B1(net68));
 sg13g2_a22oi_1 _2633_ (.Y(_1063_),
    .B1(net46),
    .B2(\pw_reg[2][0] ),
    .A2(net86),
    .A1(\pw_reg[1][0] ));
 sg13g2_a22oi_1 _2634_ (.Y(_0146_),
    .B1(_1062_),
    .B2(_1063_),
    .A2(net68),
    .A1(_1240_));
 sg13g2_a21oi_1 _2635_ (.A1(net484),
    .A2(net124),
    .Y(_1064_),
    .B1(net62));
 sg13g2_a22oi_1 _2636_ (.Y(_1065_),
    .B1(net41),
    .B2(net407),
    .A2(net88),
    .A1(net596));
 sg13g2_a22oi_1 _2637_ (.Y(_0147_),
    .B1(_1064_),
    .B2(_1065_),
    .A2(net62),
    .A1(_1239_));
 sg13g2_a21oi_1 _2638_ (.A1(net738),
    .A2(net121),
    .Y(_1066_),
    .B1(net62));
 sg13g2_a22oi_1 _2639_ (.Y(_1067_),
    .B1(net41),
    .B2(net244),
    .A2(net88),
    .A1(\pw_reg[1][2] ));
 sg13g2_a22oi_1 _2640_ (.Y(_0148_),
    .B1(_1066_),
    .B2(net245),
    .A2(net62),
    .A1(_1238_));
 sg13g2_a21oi_1 _2641_ (.A1(\pw_reg[0][3] ),
    .A2(net120),
    .Y(_1068_),
    .B1(net52));
 sg13g2_a22oi_1 _2642_ (.Y(_1069_),
    .B1(net41),
    .B2(net439),
    .A2(net84),
    .A1(\pw_reg[1][3] ));
 sg13g2_a22oi_1 _2643_ (.Y(_0149_),
    .B1(_1068_),
    .B2(net440),
    .A2(net52),
    .A1(_1237_));
 sg13g2_a21oi_1 _2644_ (.A1(net516),
    .A2(net120),
    .Y(_1070_),
    .B1(net62));
 sg13g2_a22oi_1 _2645_ (.Y(_1071_),
    .B1(net42),
    .B2(net432),
    .A2(net84),
    .A1(net564));
 sg13g2_a22oi_1 _2646_ (.Y(_0150_),
    .B1(_1070_),
    .B2(_1071_),
    .A2(net67),
    .A1(_1236_));
 sg13g2_a21oi_1 _2647_ (.A1(net487),
    .A2(net120),
    .Y(_1072_),
    .B1(net53));
 sg13g2_a22oi_1 _2648_ (.Y(_1073_),
    .B1(net42),
    .B2(\pw_reg[2][5] ),
    .A2(net84),
    .A1(\pw_reg[1][5] ));
 sg13g2_a22oi_1 _2649_ (.Y(_0151_),
    .B1(_1072_),
    .B2(_1073_),
    .A2(net53),
    .A1(_1235_));
 sg13g2_a21oi_1 _2650_ (.A1(net496),
    .A2(net121),
    .Y(_1074_),
    .B1(net67));
 sg13g2_a22oi_1 _2651_ (.Y(_1075_),
    .B1(net42),
    .B2(net615),
    .A2(net84),
    .A1(net505));
 sg13g2_a22oi_1 _2652_ (.Y(_0152_),
    .B1(_1074_),
    .B2(_1075_),
    .A2(net67),
    .A1(_1234_));
 sg13g2_a21oi_1 _2653_ (.A1(net456),
    .A2(net120),
    .Y(_1076_),
    .B1(net53));
 sg13g2_a22oi_1 _2654_ (.Y(_1077_),
    .B1(net42),
    .B2(net572),
    .A2(net85),
    .A1(net612));
 sg13g2_a22oi_1 _2655_ (.Y(_0153_),
    .B1(_1076_),
    .B2(_1077_),
    .A2(net53),
    .A1(_1233_));
 sg13g2_a21oi_1 _2656_ (.A1(net620),
    .A2(net119),
    .Y(_1078_),
    .B1(net56));
 sg13g2_a22oi_1 _2657_ (.Y(_1079_),
    .B1(net39),
    .B2(net447),
    .A2(net75),
    .A1(net588));
 sg13g2_a22oi_1 _2658_ (.Y(_0154_),
    .B1(_1078_),
    .B2(_1079_),
    .A2(net56),
    .A1(_1200_));
 sg13g2_a21oi_1 _2659_ (.A1(net625),
    .A2(net119),
    .Y(_1080_),
    .B1(net56));
 sg13g2_a22oi_1 _2660_ (.Y(_1081_),
    .B1(net39),
    .B2(net574),
    .A2(net75),
    .A1(net602));
 sg13g2_a22oi_1 _2661_ (.Y(_0155_),
    .B1(_1080_),
    .B2(_1081_),
    .A2(net56),
    .A1(_1199_));
 sg13g2_a21oi_1 _2662_ (.A1(net598),
    .A2(net118),
    .Y(_1082_),
    .B1(net57));
 sg13g2_a22oi_1 _2663_ (.Y(_1083_),
    .B1(net39),
    .B2(net420),
    .A2(net75),
    .A1(net567));
 sg13g2_a22oi_1 _2664_ (.Y(_0156_),
    .B1(_1082_),
    .B2(_1083_),
    .A2(net57),
    .A1(_1197_));
 sg13g2_a21oi_1 _2665_ (.A1(net590),
    .A2(net119),
    .Y(_1084_),
    .B1(net56));
 sg13g2_a22oi_1 _2666_ (.Y(_1085_),
    .B1(net39),
    .B2(net427),
    .A2(net75),
    .A1(net503));
 sg13g2_a22oi_1 _2667_ (.Y(_0157_),
    .B1(_1084_),
    .B2(_1085_),
    .A2(net56),
    .A1(_1198_));
 sg13g2_a21oi_1 _2668_ (.A1(net434),
    .A2(net119),
    .Y(_1086_),
    .B1(net56));
 sg13g2_a22oi_1 _2669_ (.Y(_1087_),
    .B1(net39),
    .B2(net408),
    .A2(net76),
    .A1(net468));
 sg13g2_a22oi_1 _2670_ (.Y(_0158_),
    .B1(_1086_),
    .B2(_1087_),
    .A2(net56),
    .A1(_1196_));
 sg13g2_a21oi_1 _2671_ (.A1(net569),
    .A2(net118),
    .Y(_1088_),
    .B1(net57));
 sg13g2_a22oi_1 _2672_ (.Y(_1089_),
    .B1(net39),
    .B2(net409),
    .A2(net80),
    .A1(net543));
 sg13g2_a22oi_1 _2673_ (.Y(_0159_),
    .B1(_1088_),
    .B2(net736),
    .A2(net57),
    .A1(_1194_));
 sg13g2_a21oi_1 _2674_ (.A1(net458),
    .A2(net118),
    .Y(_1090_),
    .B1(net58));
 sg13g2_a22oi_1 _2675_ (.Y(_1091_),
    .B1(net40),
    .B2(net647),
    .A2(net79),
    .A1(net424));
 sg13g2_a22oi_1 _2676_ (.Y(_0160_),
    .B1(_1090_),
    .B2(_1091_),
    .A2(net58),
    .A1(_1192_));
 sg13g2_a21oi_1 _2677_ (.A1(net537),
    .A2(net118),
    .Y(_1092_),
    .B1(net57));
 sg13g2_a22oi_1 _2678_ (.Y(_1093_),
    .B1(net39),
    .B2(net525),
    .A2(net80),
    .A1(net550));
 sg13g2_a22oi_1 _2679_ (.Y(_0161_),
    .B1(_1092_),
    .B2(_1093_),
    .A2(net57),
    .A1(_1188_));
 sg13g2_a21oi_1 _2680_ (.A1(net594),
    .A2(net118),
    .Y(_1094_),
    .B1(net60));
 sg13g2_a22oi_1 _2681_ (.Y(_1095_),
    .B1(net40),
    .B2(net616),
    .A2(net85),
    .A1(net531));
 sg13g2_a22oi_1 _2682_ (.Y(_0162_),
    .B1(_1094_),
    .B2(_1095_),
    .A2(net60),
    .A1(_1209_));
 sg13g2_a21oi_1 _2683_ (.A1(net507),
    .A2(net118),
    .Y(_1096_),
    .B1(net58));
 sg13g2_a22oi_1 _2684_ (.Y(_1097_),
    .B1(net40),
    .B2(net266),
    .A2(net79),
    .A1(net540));
 sg13g2_a22oi_1 _2685_ (.Y(_0163_),
    .B1(_1096_),
    .B2(_1097_),
    .A2(net58),
    .A1(_1208_));
 sg13g2_a21oi_1 _2686_ (.A1(\gate_latch[0] ),
    .A2(net122),
    .Y(_1098_),
    .B1(net60));
 sg13g2_a22oi_1 _2687_ (.Y(_1099_),
    .B1(net46),
    .B2(net324),
    .A2(net85),
    .A1(\gate_latch[1] ));
 sg13g2_a22oi_1 _2688_ (.Y(_0164_),
    .B1(_1098_),
    .B2(_1099_),
    .A2(net60),
    .A1(_1219_));
 sg13g2_a21oi_1 _2689_ (.A1(net586),
    .A2(net118),
    .Y(_1100_),
    .B1(net60));
 sg13g2_a22oi_1 _2690_ (.Y(_1101_),
    .B1(net40),
    .B2(net500),
    .A2(net80),
    .A1(net560));
 sg13g2_a22oi_1 _2691_ (.Y(_0165_),
    .B1(_1100_),
    .B2(_1101_),
    .A2(net60),
    .A1(net130));
 sg13g2_a21oi_1 _2692_ (.A1(net539),
    .A2(net126),
    .Y(_1102_),
    .B1(net72));
 sg13g2_a22oi_1 _2693_ (.Y(_1103_),
    .B1(net47),
    .B2(net296),
    .A2(net91),
    .A1(\attack_reg[1][0] ));
 sg13g2_a22oi_1 _2694_ (.Y(_0166_),
    .B1(_1102_),
    .B2(net297),
    .A2(net71),
    .A1(_1210_));
 sg13g2_a21oi_1 _2695_ (.A1(net251),
    .A2(net126),
    .Y(_1104_),
    .B1(net70));
 sg13g2_a22oi_1 _2696_ (.Y(_1105_),
    .B1(net47),
    .B2(net587),
    .A2(net91),
    .A1(net499));
 sg13g2_a22oi_1 _2697_ (.Y(_0167_),
    .B1(net252),
    .B2(_1105_),
    .A2(net70),
    .A1(_1216_));
 sg13g2_a21oi_1 _2698_ (.A1(net248),
    .A2(net126),
    .Y(_1106_),
    .B1(net70));
 sg13g2_a22oi_1 _2699_ (.Y(_1107_),
    .B1(net47),
    .B2(net573),
    .A2(net91),
    .A1(net614));
 sg13g2_a22oi_1 _2700_ (.Y(_0168_),
    .B1(net249),
    .B2(_1107_),
    .A2(net70),
    .A1(_1217_));
 sg13g2_a21oi_1 _2701_ (.A1(net254),
    .A2(net126),
    .Y(_1108_),
    .B1(net70));
 sg13g2_a22oi_1 _2702_ (.Y(_1109_),
    .B1(net47),
    .B2(net515),
    .A2(net91),
    .A1(net494));
 sg13g2_a22oi_1 _2703_ (.Y(_0169_),
    .B1(net255),
    .B2(_1109_),
    .A2(net70),
    .A1(_1218_));
 sg13g2_a21oi_1 _2704_ (.A1(\attack_reg[0][4] ),
    .A2(net127),
    .Y(_1110_),
    .B1(net71));
 sg13g2_a22oi_1 _2705_ (.Y(_1111_),
    .B1(net47),
    .B2(net378),
    .A2(net91),
    .A1(\attack_reg[1][4] ));
 sg13g2_a22oi_1 _2706_ (.Y(_0170_),
    .B1(_1110_),
    .B2(net379),
    .A2(net71),
    .A1(_1204_));
 sg13g2_a21oi_1 _2707_ (.A1(net450),
    .A2(net127),
    .Y(_1112_),
    .B1(net71));
 sg13g2_a22oi_1 _2708_ (.Y(_1113_),
    .B1(net47),
    .B2(net460),
    .A2(net91),
    .A1(net459));
 sg13g2_a22oi_1 _2709_ (.Y(_0171_),
    .B1(_1112_),
    .B2(_1113_),
    .A2(net71),
    .A1(_1205_));
 sg13g2_a21oi_1 _2710_ (.A1(net429),
    .A2(net127),
    .Y(_1114_),
    .B1(net71));
 sg13g2_a22oi_1 _2711_ (.Y(_1115_),
    .B1(net48),
    .B2(net527),
    .A2(net91),
    .A1(net546));
 sg13g2_a22oi_1 _2712_ (.Y(_0172_),
    .B1(_1114_),
    .B2(_1115_),
    .A2(net72),
    .A1(_1207_));
 sg13g2_a21oi_1 _2713_ (.A1(net521),
    .A2(net127),
    .Y(_1116_),
    .B1(net71));
 sg13g2_a22oi_1 _2714_ (.Y(_1117_),
    .B1(net48),
    .B2(net483),
    .A2(net92),
    .A1(\attack_reg[1][7] ));
 sg13g2_a22oi_1 _2715_ (.Y(_0173_),
    .B1(_1116_),
    .B2(_1117_),
    .A2(net71),
    .A1(_1206_));
 sg13g2_a21oi_1 _2716_ (.A1(net490),
    .A2(net122),
    .Y(_1118_),
    .B1(net68));
 sg13g2_a22oi_1 _2717_ (.Y(_1119_),
    .B1(net46),
    .B2(net611),
    .A2(net86),
    .A1(net514));
 sg13g2_a22oi_1 _2718_ (.Y(_0174_),
    .B1(_1118_),
    .B2(_1119_),
    .A2(net68),
    .A1(_1195_));
 sg13g2_a21oi_1 _2719_ (.A1(net506),
    .A2(net122),
    .Y(_1120_),
    .B1(net68));
 sg13g2_a22oi_1 _2720_ (.Y(_1121_),
    .B1(net46),
    .B2(net644),
    .A2(net86),
    .A1(net600));
 sg13g2_a22oi_1 _2721_ (.Y(_0175_),
    .B1(_1120_),
    .B2(_1121_),
    .A2(net68),
    .A1(_1193_));
 sg13g2_a21oi_1 _2722_ (.A1(net606),
    .A2(net122),
    .Y(_1122_),
    .B1(net59));
 sg13g2_a22oi_1 _2723_ (.Y(_1123_),
    .B1(net46),
    .B2(net512),
    .A2(net85),
    .A1(net638));
 sg13g2_a22oi_1 _2724_ (.Y(_0176_),
    .B1(_1122_),
    .B2(_1123_),
    .A2(net59),
    .A1(_1191_));
 sg13g2_a21oi_1 _2725_ (.A1(net610),
    .A2(net122),
    .Y(_1124_),
    .B1(net59));
 sg13g2_a22oi_1 _2726_ (.Y(_1125_),
    .B1(net46),
    .B2(net549),
    .A2(net85),
    .A1(net524));
 sg13g2_a22oi_1 _2727_ (.Y(_0177_),
    .B1(_1124_),
    .B2(_1125_),
    .A2(net59),
    .A1(_1190_));
 sg13g2_a21oi_1 _2728_ (.A1(net568),
    .A2(net126),
    .Y(_1126_),
    .B1(net68));
 sg13g2_a22oi_1 _2729_ (.Y(_1127_),
    .B1(net46),
    .B2(net473),
    .A2(net86),
    .A1(net474));
 sg13g2_a22oi_1 _2730_ (.Y(_0178_),
    .B1(_1126_),
    .B2(_1127_),
    .A2(net68),
    .A1(_1211_));
 sg13g2_a21oi_1 _2731_ (.A1(net650),
    .A2(net122),
    .Y(_1128_),
    .B1(net69));
 sg13g2_a22oi_1 _2732_ (.Y(_1129_),
    .B1(net46),
    .B2(net422),
    .A2(net86),
    .A1(net635));
 sg13g2_a22oi_1 _2733_ (.Y(_0179_),
    .B1(_1128_),
    .B2(_1129_),
    .A2(net69),
    .A1(_1212_));
 sg13g2_a21oi_1 _2734_ (.A1(net435),
    .A2(net126),
    .Y(_1130_),
    .B1(net69));
 sg13g2_a22oi_1 _2735_ (.Y(_1131_),
    .B1(net48),
    .B2(net495),
    .A2(net92),
    .A1(net608));
 sg13g2_a22oi_1 _2736_ (.Y(_0180_),
    .B1(_1130_),
    .B2(_1131_),
    .A2(net69),
    .A1(_1214_));
 sg13g2_a21oi_1 _2737_ (.A1(net437),
    .A2(net123),
    .Y(_1132_),
    .B1(net69));
 sg13g2_a22oi_1 _2738_ (.Y(_1133_),
    .B1(net48),
    .B2(net582),
    .A2(net86),
    .A1(net605));
 sg13g2_a22oi_1 _2739_ (.Y(_0181_),
    .B1(_1132_),
    .B2(_1133_),
    .A2(net69),
    .A1(_1213_));
 sg13g2_a21oi_1 _2740_ (.A1(_1225_),
    .A2(net76),
    .Y(_1134_),
    .B1(_1273_));
 sg13g2_o21ai_1 _2741_ (.B1(_1134_),
    .Y(_1135_),
    .A1(net529),
    .A2(net76));
 sg13g2_a21oi_1 _2742_ (.A1(net501),
    .A2(net119),
    .Y(_1136_),
    .B1(net55));
 sg13g2_a22oi_1 _2743_ (.Y(_0182_),
    .B1(_1135_),
    .B2(_1136_),
    .A2(net55),
    .A1(_1186_));
 sg13g2_nor3_1 _2744_ (.A(net5),
    .B(net471),
    .C(_1222_),
    .Y(_1137_));
 sg13g2_nand2b_1 _2745_ (.Y(_1138_),
    .B(_1137_),
    .A_N(net6));
 sg13g2_nor4_1 _2746_ (.A(net4),
    .B(net2),
    .C(net3),
    .D(_1138_),
    .Y(_1139_));
 sg13g2_mux2_1 _2747_ (.A0(net488),
    .A1(net151),
    .S(_1139_),
    .X(_0183_));
 sg13g2_mux2_1 _2748_ (.A0(net509),
    .A1(net149),
    .S(_1139_),
    .X(_0184_));
 sg13g2_mux2_1 _2749_ (.A0(net482),
    .A1(net162),
    .S(_1139_),
    .X(_0185_));
 sg13g2_mux2_1 _2750_ (.A0(net561),
    .A1(net161),
    .S(_1139_),
    .X(_0186_));
 sg13g2_mux2_1 _2751_ (.A0(net607),
    .A1(net158),
    .S(_1139_),
    .X(_0187_));
 sg13g2_mux2_1 _2752_ (.A0(net554),
    .A1(net157),
    .S(_1139_),
    .X(_0188_));
 sg13g2_mux2_1 _2753_ (.A0(net489),
    .A1(net154),
    .S(_1139_),
    .X(_0189_));
 sg13g2_mux2_1 _2754_ (.A0(net576),
    .A1(net152),
    .S(_1139_),
    .X(_0190_));
 sg13g2_or4_1 _2755_ (.A(_1221_),
    .B(net6),
    .C(net471),
    .D(_1222_),
    .X(_1140_));
 sg13g2_nor4_1 _2756_ (.A(net4),
    .B(net2),
    .C(net3),
    .D(_1140_),
    .Y(_1141_));
 sg13g2_mux2_1 _2757_ (.A0(net534),
    .A1(net151),
    .S(_1141_),
    .X(_0191_));
 sg13g2_mux2_1 _2758_ (.A0(net478),
    .A1(net149),
    .S(_1141_),
    .X(_0192_));
 sg13g2_mux2_1 _2759_ (.A0(net545),
    .A1(net163),
    .S(_1141_),
    .X(_0193_));
 sg13g2_mux2_1 _2760_ (.A0(net510),
    .A1(net161),
    .S(_1141_),
    .X(_0194_));
 sg13g2_mux2_1 _2761_ (.A0(net581),
    .A1(net158),
    .S(_1141_),
    .X(_0195_));
 sg13g2_mux2_1 _2762_ (.A0(net455),
    .A1(net157),
    .S(_1141_),
    .X(_0196_));
 sg13g2_mux2_1 _2763_ (.A0(net491),
    .A1(net154),
    .S(_1141_),
    .X(_0197_));
 sg13g2_mux2_1 _2764_ (.A0(net580),
    .A1(net153),
    .S(_1141_),
    .X(_0198_));
 sg13g2_nand2_1 _2765_ (.Y(_1142_),
    .A(net6),
    .B(_1137_));
 sg13g2_or4_1 _2766_ (.A(net4),
    .B(net2),
    .C(net3),
    .D(_1142_),
    .X(_1143_));
 sg13g2_mux2_1 _2767_ (.A0(net151),
    .A1(net547),
    .S(_1143_),
    .X(_0199_));
 sg13g2_mux2_1 _2768_ (.A0(net149),
    .A1(net470),
    .S(_1143_),
    .X(_0200_));
 sg13g2_mux2_1 _2769_ (.A0(net163),
    .A1(net579),
    .S(_1143_),
    .X(_0201_));
 sg13g2_mux2_1 _2770_ (.A0(net161),
    .A1(net457),
    .S(_1143_),
    .X(_0202_));
 sg13g2_mux2_1 _2771_ (.A0(net158),
    .A1(net619),
    .S(_1143_),
    .X(_0203_));
 sg13g2_mux2_1 _2772_ (.A0(net157),
    .A1(net528),
    .S(_1143_),
    .X(_0204_));
 sg13g2_mux2_1 _2773_ (.A0(net154),
    .A1(net562),
    .S(_1143_),
    .X(_0205_));
 sg13g2_mux2_1 _2774_ (.A0(net153),
    .A1(net557),
    .S(_1143_),
    .X(_0206_));
 sg13g2_nand3_1 _2775_ (.B(_1224_),
    .C(net3),
    .A(net4),
    .Y(_1144_));
 sg13g2_nor2_1 _2776_ (.A(_1138_),
    .B(_1144_),
    .Y(_1145_));
 sg13g2_mux2_1 _2777_ (.A0(net552),
    .A1(net150),
    .S(_1145_),
    .X(_0207_));
 sg13g2_mux2_1 _2778_ (.A0(net513),
    .A1(net148),
    .S(_1145_),
    .X(_0208_));
 sg13g2_mux2_1 _2779_ (.A0(net462),
    .A1(net162),
    .S(_1145_),
    .X(_0209_));
 sg13g2_mux2_1 _2780_ (.A0(net592),
    .A1(net160),
    .S(_1145_),
    .X(_0210_));
 sg13g2_mux2_1 _2781_ (.A0(net627),
    .A1(net159),
    .S(_1145_),
    .X(_0211_));
 sg13g2_mux2_1 _2782_ (.A0(net425),
    .A1(net156),
    .S(_1145_),
    .X(_0212_));
 sg13g2_mux2_1 _2783_ (.A0(net533),
    .A1(net155),
    .S(_1145_),
    .X(_0213_));
 sg13g2_mux2_1 _2784_ (.A0(net517),
    .A1(net152),
    .S(_1145_),
    .X(_0214_));
 sg13g2_nor2_1 _2785_ (.A(_1140_),
    .B(_1144_),
    .Y(_1146_));
 sg13g2_mux2_1 _2786_ (.A0(net553),
    .A1(net150),
    .S(_1146_),
    .X(_0215_));
 sg13g2_mux2_1 _2787_ (.A0(net421),
    .A1(net148),
    .S(_1146_),
    .X(_0216_));
 sg13g2_mux2_1 _2788_ (.A0(net485),
    .A1(net162),
    .S(_1146_),
    .X(_0217_));
 sg13g2_mux2_1 _2789_ (.A0(net636),
    .A1(net160),
    .S(_1146_),
    .X(_0218_));
 sg13g2_mux2_1 _2790_ (.A0(net613),
    .A1(net159),
    .S(_1146_),
    .X(_0219_));
 sg13g2_mux2_1 _2791_ (.A0(net502),
    .A1(net156),
    .S(_1146_),
    .X(_0220_));
 sg13g2_mux2_1 _2792_ (.A0(net631),
    .A1(net155),
    .S(_1146_),
    .X(_0221_));
 sg13g2_mux2_1 _2793_ (.A0(net453),
    .A1(net152),
    .S(_1146_),
    .X(_0222_));
 sg13g2_nor2_1 _2794_ (.A(_1142_),
    .B(_1144_),
    .Y(_1147_));
 sg13g2_mux2_1 _2795_ (.A0(net593),
    .A1(net150),
    .S(_1147_),
    .X(_0223_));
 sg13g2_mux2_1 _2796_ (.A0(net469),
    .A1(net148),
    .S(_1147_),
    .X(_0224_));
 sg13g2_mux2_1 _2797_ (.A0(net535),
    .A1(net162),
    .S(_1147_),
    .X(_0225_));
 sg13g2_mux2_1 _2798_ (.A0(net511),
    .A1(net160),
    .S(_1147_),
    .X(_0226_));
 sg13g2_mux2_1 _2799_ (.A0(net536),
    .A1(net159),
    .S(_1147_),
    .X(_0227_));
 sg13g2_mux2_1 _2800_ (.A0(net556),
    .A1(net156),
    .S(_1147_),
    .X(_0228_));
 sg13g2_mux2_1 _2801_ (.A0(net518),
    .A1(net155),
    .S(_1147_),
    .X(_0229_));
 sg13g2_mux2_1 _2802_ (.A0(net597),
    .A1(net152),
    .S(_1147_),
    .X(_0230_));
 sg13g2_nand3_1 _2803_ (.B(_1224_),
    .C(net3),
    .A(_1223_),
    .Y(_1148_));
 sg13g2_or2_1 _2804_ (.X(_1149_),
    .B(_1148_),
    .A(_1138_));
 sg13g2_mux2_1 _2805_ (.A0(net150),
    .A1(net446),
    .S(_1149_),
    .X(_0231_));
 sg13g2_mux2_1 _2806_ (.A0(net148),
    .A1(net484),
    .S(_1149_),
    .X(_0232_));
 sg13g2_mux2_1 _2807_ (.A0(net162),
    .A1(net486),
    .S(_1149_),
    .X(_0233_));
 sg13g2_mux2_1 _2808_ (.A0(net160),
    .A1(net498),
    .S(_1149_),
    .X(_0234_));
 sg13g2_mux2_1 _2809_ (.A0(net159),
    .A1(net516),
    .S(_1149_),
    .X(_0235_));
 sg13g2_mux2_1 _2810_ (.A0(net156),
    .A1(net487),
    .S(_1149_),
    .X(_0236_));
 sg13g2_mux2_1 _2811_ (.A0(net155),
    .A1(net496),
    .S(_1149_),
    .X(_0237_));
 sg13g2_mux2_1 _2812_ (.A0(net152),
    .A1(net456),
    .S(_1149_),
    .X(_0238_));
 sg13g2_nor2_1 _2813_ (.A(_1140_),
    .B(_1148_),
    .Y(_1150_));
 sg13g2_mux2_1 _2814_ (.A0(net448),
    .A1(net150),
    .S(_1150_),
    .X(_0239_));
 sg13g2_mux2_1 _2815_ (.A0(net596),
    .A1(net148),
    .S(_1150_),
    .X(_0240_));
 sg13g2_mux2_1 _2816_ (.A0(net544),
    .A1(net163),
    .S(_1150_),
    .X(_0241_));
 sg13g2_mux2_1 _2817_ (.A0(net558),
    .A1(net160),
    .S(_1150_),
    .X(_0242_));
 sg13g2_mux2_1 _2818_ (.A0(net564),
    .A1(net159),
    .S(_1150_),
    .X(_0243_));
 sg13g2_mux2_1 _2819_ (.A0(net497),
    .A1(net156),
    .S(_1150_),
    .X(_0244_));
 sg13g2_mux2_1 _2820_ (.A0(net505),
    .A1(net155),
    .S(_1150_),
    .X(_0245_));
 sg13g2_mux2_1 _2821_ (.A0(net612),
    .A1(net152),
    .S(_1150_),
    .X(_0246_));
 sg13g2_nor2_1 _2822_ (.A(_1142_),
    .B(_1148_),
    .Y(_1151_));
 sg13g2_mux2_1 _2823_ (.A0(net566),
    .A1(net151),
    .S(_1151_),
    .X(_0247_));
 sg13g2_mux2_1 _2824_ (.A0(net407),
    .A1(net148),
    .S(_1151_),
    .X(_0248_));
 sg13g2_mux2_1 _2825_ (.A0(net244),
    .A1(net163),
    .S(_1151_),
    .X(_0249_));
 sg13g2_mux2_1 _2826_ (.A0(net439),
    .A1(net161),
    .S(_1151_),
    .X(_0250_));
 sg13g2_mux2_1 _2827_ (.A0(net432),
    .A1(net159),
    .S(_1151_),
    .X(_0251_));
 sg13g2_mux2_1 _2828_ (.A0(net559),
    .A1(net156),
    .S(_1151_),
    .X(_0252_));
 sg13g2_mux2_1 _2829_ (.A0(net615),
    .A1(net155),
    .S(_1151_),
    .X(_0253_));
 sg13g2_mux2_1 _2830_ (.A0(net572),
    .A1(net152),
    .S(_1151_),
    .X(_0254_));
 sg13g2_nor3_1 _2831_ (.A(_1223_),
    .B(net2),
    .C(net3),
    .Y(_1152_));
 sg13g2_nand2b_1 _2832_ (.Y(_1153_),
    .B(_1152_),
    .A_N(_1138_));
 sg13g2_mux2_1 _2833_ (.A0(net151),
    .A1(net539),
    .S(_1153_),
    .X(_0255_));
 sg13g2_mux2_1 _2834_ (.A0(net149),
    .A1(net251),
    .S(_1153_),
    .X(_0256_));
 sg13g2_mux2_1 _2835_ (.A0(net163),
    .A1(net248),
    .S(_1153_),
    .X(_0257_));
 sg13g2_mux2_1 _2836_ (.A0(net161),
    .A1(net254),
    .S(_1153_),
    .X(_0258_));
 sg13g2_mux2_1 _2837_ (.A0(net158),
    .A1(net563),
    .S(_1153_),
    .X(_0259_));
 sg13g2_mux2_1 _2838_ (.A0(net157),
    .A1(net450),
    .S(_1153_),
    .X(_0260_));
 sg13g2_mux2_1 _2839_ (.A0(net154),
    .A1(net429),
    .S(_1153_),
    .X(_0261_));
 sg13g2_mux2_1 _2840_ (.A0(net153),
    .A1(net521),
    .S(_1153_),
    .X(_0262_));
 sg13g2_nor2b_1 _2841_ (.A(_1140_),
    .B_N(_1152_),
    .Y(_1154_));
 sg13g2_mux2_1 _2842_ (.A0(net472),
    .A1(net151),
    .S(_1154_),
    .X(_0263_));
 sg13g2_mux2_1 _2843_ (.A0(net499),
    .A1(net149),
    .S(_1154_),
    .X(_0264_));
 sg13g2_mux2_1 _2844_ (.A0(net614),
    .A1(net163),
    .S(_1154_),
    .X(_0265_));
 sg13g2_mux2_1 _2845_ (.A0(net494),
    .A1(net161),
    .S(_1154_),
    .X(_0266_));
 sg13g2_mux2_1 _2846_ (.A0(net551),
    .A1(net158),
    .S(_1154_),
    .X(_0267_));
 sg13g2_mux2_1 _2847_ (.A0(net459),
    .A1(net157),
    .S(_1154_),
    .X(_0268_));
 sg13g2_mux2_1 _2848_ (.A0(net546),
    .A1(net154),
    .S(_1154_),
    .X(_0269_));
 sg13g2_mux2_1 _2849_ (.A0(net634),
    .A1(net153),
    .S(_1154_),
    .X(_0270_));
 sg13g2_nand3_1 _2850_ (.B(_1137_),
    .C(_1152_),
    .A(net6),
    .Y(_1155_));
 sg13g2_mux2_1 _2851_ (.A0(net151),
    .A1(net296),
    .S(_1155_),
    .X(_0271_));
 sg13g2_mux2_1 _2852_ (.A0(net149),
    .A1(net587),
    .S(_1155_),
    .X(_0272_));
 sg13g2_mux2_1 _2853_ (.A0(net163),
    .A1(net573),
    .S(_1155_),
    .X(_0273_));
 sg13g2_mux2_1 _2854_ (.A0(net161),
    .A1(net515),
    .S(_1155_),
    .X(_0274_));
 sg13g2_mux2_1 _2855_ (.A0(net158),
    .A1(net378),
    .S(_1155_),
    .X(_0275_));
 sg13g2_mux2_1 _2856_ (.A0(net157),
    .A1(net460),
    .S(_1155_),
    .X(_0276_));
 sg13g2_mux2_1 _2857_ (.A0(net155),
    .A1(net527),
    .S(_1155_),
    .X(_0277_));
 sg13g2_mux2_1 _2858_ (.A0(net153),
    .A1(net483),
    .S(_1155_),
    .X(_0278_));
 sg13g2_nand3b_1 _2859_ (.B(net2),
    .C(net4),
    .Y(_1156_),
    .A_N(net3));
 sg13g2_nor2_1 _2860_ (.A(_1138_),
    .B(_1156_),
    .Y(_1157_));
 sg13g2_mux2_1 _2861_ (.A0(net490),
    .A1(net150),
    .S(_1157_),
    .X(_0279_));
 sg13g2_mux2_1 _2862_ (.A0(net506),
    .A1(net148),
    .S(_1157_),
    .X(_0280_));
 sg13g2_mux2_1 _2863_ (.A0(net606),
    .A1(net162),
    .S(_1157_),
    .X(_0281_));
 sg13g2_mux2_1 _2864_ (.A0(net610),
    .A1(net160),
    .S(_1157_),
    .X(_0282_));
 sg13g2_mux2_1 _2865_ (.A0(net568),
    .A1(net158),
    .S(_1157_),
    .X(_0283_));
 sg13g2_mux2_1 _2866_ (.A0(net650),
    .A1(net156),
    .S(_1157_),
    .X(_0284_));
 sg13g2_mux2_1 _2867_ (.A0(net435),
    .A1(net154),
    .S(_1157_),
    .X(_0285_));
 sg13g2_mux2_1 _2868_ (.A0(net437),
    .A1(net152),
    .S(_1157_),
    .X(_0286_));
 sg13g2_nor2_1 _2869_ (.A(_1140_),
    .B(_1156_),
    .Y(_1158_));
 sg13g2_mux2_1 _2870_ (.A0(net514),
    .A1(net150),
    .S(_1158_),
    .X(_0287_));
 sg13g2_mux2_1 _2871_ (.A0(net600),
    .A1(net148),
    .S(_1158_),
    .X(_0288_));
 sg13g2_mux2_1 _2872_ (.A0(net638),
    .A1(net162),
    .S(_1158_),
    .X(_0289_));
 sg13g2_mux2_1 _2873_ (.A0(net524),
    .A1(net160),
    .S(_1158_),
    .X(_0290_));
 sg13g2_mux2_1 _2874_ (.A0(net474),
    .A1(net158),
    .S(_1158_),
    .X(_0291_));
 sg13g2_mux2_1 _2875_ (.A0(net635),
    .A1(net156),
    .S(_1158_),
    .X(_0292_));
 sg13g2_mux2_1 _2876_ (.A0(net608),
    .A1(net154),
    .S(_1158_),
    .X(_0293_));
 sg13g2_mux2_1 _2877_ (.A0(net605),
    .A1(net153),
    .S(_1158_),
    .X(_0294_));
 sg13g2_nor2_1 _2878_ (.A(_1142_),
    .B(_1156_),
    .Y(_1159_));
 sg13g2_mux2_1 _2879_ (.A0(net611),
    .A1(net150),
    .S(_1159_),
    .X(_0295_));
 sg13g2_mux2_1 _2880_ (.A0(net644),
    .A1(net149),
    .S(_1159_),
    .X(_0296_));
 sg13g2_mux2_1 _2881_ (.A0(net512),
    .A1(net162),
    .S(_1159_),
    .X(_0297_));
 sg13g2_mux2_1 _2882_ (.A0(net549),
    .A1(net160),
    .S(_1159_),
    .X(_0298_));
 sg13g2_mux2_1 _2883_ (.A0(net473),
    .A1(net159),
    .S(_1159_),
    .X(_0299_));
 sg13g2_mux2_1 _2884_ (.A0(net422),
    .A1(net157),
    .S(_1159_),
    .X(_0300_));
 sg13g2_mux2_1 _2885_ (.A0(net495),
    .A1(net154),
    .S(_1159_),
    .X(_0301_));
 sg13g2_mux2_1 _2886_ (.A0(net582),
    .A1(net153),
    .S(_1159_),
    .X(_0302_));
 sg13g2_dfrbpq_1 _2887_ (.RESET_B(net166),
    .D(net359),
    .Q(\mix_acc[0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2888_ (.RESET_B(net166),
    .D(net689),
    .Q(\mix_acc[1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2889_ (.RESET_B(net166),
    .D(net704),
    .Q(\mix_acc[2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2890_ (.RESET_B(net164),
    .D(net725),
    .Q(\mix_acc[3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2891_ (.RESET_B(net164),
    .D(net710),
    .Q(\mix_acc[4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2892_ (.RESET_B(net166),
    .D(_0308_),
    .Q(\mix_acc[5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2893_ (.RESET_B(net165),
    .D(net718),
    .Q(\mix_acc[6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2894_ (.RESET_B(net168),
    .D(net713),
    .Q(\mix_acc[7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2895_ (.RESET_B(net167),
    .D(net313),
    .Q(\mix_acc[8] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2896_ (.RESET_B(net167),
    .D(_0312_),
    .Q(\mix_acc[9] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2897_ (.RESET_B(net164),
    .D(net373),
    .Q(\mix_out[0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2898_ (.RESET_B(net164),
    .D(net653),
    .Q(\mix_out[1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2899_ (.RESET_B(net164),
    .D(net393),
    .Q(\mix_out[2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2900_ (.RESET_B(net165),
    .D(net520),
    .Q(\mix_out[3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2901_ (.RESET_B(net165),
    .D(net336),
    .Q(\mix_out[4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2902_ (.RESET_B(net167),
    .D(_0318_),
    .Q(\mix_out[5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2903_ (.RESET_B(net167),
    .D(_0319_),
    .Q(\mix_out[6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2904_ (.RESET_B(net167),
    .D(net319),
    .Q(\mix_out[7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2905_ (.RESET_B(net210),
    .D(net622),
    .Q(\acc[0][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2906_ (.RESET_B(net202),
    .D(net404),
    .Q(\acc[0][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2907_ (.RESET_B(net208),
    .D(net377),
    .Q(\acc[0][2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2908_ (.RESET_B(net207),
    .D(net355),
    .Q(\acc[0][3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2909_ (.RESET_B(net203),
    .D(net465),
    .Q(\acc[0][4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2910_ (.RESET_B(net202),
    .D(net330),
    .Q(\acc[0][5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2911_ (.RESET_B(net202),
    .D(net357),
    .Q(\acc[0][6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2912_ (.RESET_B(net189),
    .D(net328),
    .Q(\acc[0][7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2913_ (.RESET_B(net188),
    .D(net467),
    .Q(\acc[0][8] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2914_ (.RESET_B(net184),
    .D(net347),
    .Q(\acc[0][9] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2915_ (.RESET_B(net185),
    .D(net401),
    .Q(\acc[0][10] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2916_ (.RESET_B(net174),
    .D(_0332_),
    .Q(\acc[0][11] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2917_ (.RESET_B(net184),
    .D(net395),
    .Q(\acc[0][12] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2918_ (.RESET_B(net174),
    .D(net338),
    .Q(\acc[0][13] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2919_ (.RESET_B(net174),
    .D(net383),
    .Q(\acc[0][14] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2920_ (.RESET_B(net171),
    .D(net706),
    .Q(\acc[0][15] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2921_ (.RESET_B(net205),
    .D(net334),
    .Q(\acc[1][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2922_ (.RESET_B(net203),
    .D(net387),
    .Q(\acc[1][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2923_ (.RESET_B(net208),
    .D(net385),
    .Q(\acc[1][2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2924_ (.RESET_B(net207),
    .D(net415),
    .Q(\acc[1][3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2925_ (.RESET_B(net203),
    .D(net445),
    .Q(\acc[1][4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2926_ (.RESET_B(net202),
    .D(net389),
    .Q(\acc[1][5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2927_ (.RESET_B(net189),
    .D(net345),
    .Q(\acc[1][6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2928_ (.RESET_B(net189),
    .D(net375),
    .Q(\acc[1][7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2929_ (.RESET_B(net188),
    .D(net443),
    .Q(\acc[1][8] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2930_ (.RESET_B(net184),
    .D(net368),
    .Q(\acc[1][9] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2931_ (.RESET_B(net185),
    .D(net351),
    .Q(\acc[1][10] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2932_ (.RESET_B(net174),
    .D(net523),
    .Q(\acc[1][11] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2933_ (.RESET_B(net184),
    .D(net413),
    .Q(\acc[1][12] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2934_ (.RESET_B(net175),
    .D(net411),
    .Q(\acc[1][13] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2935_ (.RESET_B(net174),
    .D(net391),
    .Q(\acc[1][14] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2936_ (.RESET_B(net171),
    .D(net676),
    .Q(\acc[1][15] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2937_ (.RESET_B(net205),
    .D(net304),
    .Q(\acc[2][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2938_ (.RESET_B(net203),
    .D(net289),
    .Q(\acc[2][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2939_ (.RESET_B(net208),
    .D(net277),
    .Q(\acc[2][2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2940_ (.RESET_B(net207),
    .D(net295),
    .Q(\acc[2][3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2941_ (.RESET_B(net203),
    .D(net286),
    .Q(\acc[2][4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2942_ (.RESET_B(net202),
    .D(net265),
    .Q(\acc[2][5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2943_ (.RESET_B(net189),
    .D(net274),
    .Q(\acc[2][6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2944_ (.RESET_B(net189),
    .D(net310),
    .Q(\acc[2][7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2945_ (.RESET_B(net188),
    .D(net283),
    .Q(\acc[2][8] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2946_ (.RESET_B(net184),
    .D(net271),
    .Q(\acc[2][9] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2947_ (.RESET_B(net185),
    .D(net321),
    .Q(\acc[2][10] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2948_ (.RESET_B(net175),
    .D(net292),
    .Q(\acc[2][11] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2949_ (.RESET_B(net184),
    .D(net326),
    .Q(\acc[2][12] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2950_ (.RESET_B(net175),
    .D(net301),
    .Q(\acc[2][13] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2951_ (.RESET_B(net174),
    .D(net323),
    .Q(\acc[2][14] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2952_ (.RESET_B(net171),
    .D(net349),
    .Q(\acc[2][15] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2953_ (.RESET_B(net169),
    .D(_0060_),
    .Q(\env[0][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2954_ (.RESET_B(net169),
    .D(_0061_),
    .Q(\env[0][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2955_ (.RESET_B(net178),
    .D(_0062_),
    .Q(\env[0][2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2956_ (.RESET_B(net169),
    .D(net591),
    .Q(\env[0][3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2957_ (.RESET_B(net178),
    .D(_0064_),
    .Q(\env[0][4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2958_ (.RESET_B(net180),
    .D(_0065_),
    .Q(\env[0][5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2959_ (.RESET_B(net180),
    .D(_0066_),
    .Q(\env[0][6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2960_ (.RESET_B(net180),
    .D(_0067_),
    .Q(\env[0][7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2961_ (.RESET_B(net169),
    .D(_0068_),
    .Q(\env[1][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2962_ (.RESET_B(net169),
    .D(net603),
    .Q(\env[1][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2963_ (.RESET_B(net178),
    .D(_0070_),
    .Q(\env[1][2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2964_ (.RESET_B(net170),
    .D(net504),
    .Q(\env[1][3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2965_ (.RESET_B(net178),
    .D(_0072_),
    .Q(\env[1][4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2966_ (.RESET_B(net178),
    .D(_0073_),
    .Q(\env[1][5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2967_ (.RESET_B(net180),
    .D(_0074_),
    .Q(\env[1][6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2968_ (.RESET_B(net178),
    .D(_0075_),
    .Q(\env[1][7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2969_ (.RESET_B(net169),
    .D(_0076_),
    .Q(\env[2][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2970_ (.RESET_B(net169),
    .D(net575),
    .Q(\env[2][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2971_ (.RESET_B(net179),
    .D(_0078_),
    .Q(\env[2][2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2972_ (.RESET_B(net169),
    .D(net428),
    .Q(\env[2][3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2973_ (.RESET_B(net178),
    .D(_0080_),
    .Q(\env[2][4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2974_ (.RESET_B(net178),
    .D(_0081_),
    .Q(\env[2][5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2975_ (.RESET_B(net180),
    .D(_0082_),
    .Q(\env[2][6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2976_ (.RESET_B(net180),
    .D(net526),
    .Q(\env[2][7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2977_ (.RESET_B(net195),
    .D(net595),
    .Q(\ast[0][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2978_ (.RESET_B(net193),
    .D(net508),
    .Q(\ast[0][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2979_ (.RESET_B(net195),
    .D(net532),
    .Q(\ast[1][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2980_ (.RESET_B(net193),
    .D(net541),
    .Q(\ast[1][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2981_ (.RESET_B(net195),
    .D(net617),
    .Q(\ast[2][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2982_ (.RESET_B(net193),
    .D(net268),
    .Q(\ast[2][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2983_ (.RESET_B(net195),
    .D(_0090_),
    .Q(\gate_latch[0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2984_ (.RESET_B(net195),
    .D(_0091_),
    .Q(\gate_latch[1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2985_ (.RESET_B(net195),
    .D(_0092_),
    .Q(\gate_latch[2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2986_ (.RESET_B(net182),
    .D(_0093_),
    .Q(\releasing[0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2987_ (.RESET_B(net182),
    .D(_0094_),
    .Q(\releasing[1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2988_ (.RESET_B(net182),
    .D(_0095_),
    .Q(\releasing[2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2989_ (.RESET_B(net171),
    .D(net353),
    .Q(\prev_msb_d[0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2990_ (.RESET_B(net171),
    .D(net530),
    .Q(\prev_msb_d[1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2991_ (.RESET_B(net171),
    .D(_0098_),
    .Q(\prev_msb_d[2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2992_ (.RESET_B(net172),
    .D(net341),
    .Q(_0025_),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2993_ (.RESET_B(net172),
    .D(net406),
    .Q(_0026_),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2994_ (.RESET_B(net172),
    .D(_0101_),
    .Q(_0027_),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2995_ (.RESET_B(net172),
    .D(net399),
    .Q(_0028_),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2996_ (.RESET_B(net171),
    .D(net571),
    .Q(_0029_),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2997_ (.RESET_B(net173),
    .D(_0104_),
    .Q(_0030_),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2998_ (.RESET_B(net173),
    .D(net419),
    .Q(_0031_),
    .CLK(clk));
 sg13g2_dfrbpq_1 _2999_ (.RESET_B(net173),
    .D(net431),
    .Q(_0032_),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3000_ (.RESET_B(net173),
    .D(_0107_),
    .Q(_0033_),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3001_ (.RESET_B(net173),
    .D(_0108_),
    .Q(_0034_),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3002_ (.RESET_B(net173),
    .D(net667),
    .Q(_0035_),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3003_ (.RESET_B(net183),
    .D(_0110_),
    .Q(_0036_),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3004_ (.RESET_B(net176),
    .D(net663),
    .Q(_0037_),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3005_ (.RESET_B(net176),
    .D(_0112_),
    .Q(_0038_),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3006_ (.RESET_B(net176),
    .D(_0113_),
    .Q(_0039_),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3007_ (.RESET_B(net210),
    .D(_0114_),
    .Q(\p_acc[0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3008_ (.RESET_B(net203),
    .D(_0115_),
    .Q(\p_acc[1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3009_ (.RESET_B(net208),
    .D(_0116_),
    .Q(\p_acc[2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3010_ (.RESET_B(net207),
    .D(_0117_),
    .Q(\p_acc[3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3011_ (.RESET_B(net207),
    .D(net452),
    .Q(\p_acc[4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3012_ (.RESET_B(net202),
    .D(_0119_),
    .Q(\p_acc[5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3013_ (.RESET_B(net202),
    .D(_0120_),
    .Q(\p_acc[6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3014_ (.RESET_B(net189),
    .D(_0121_),
    .Q(\p_acc[7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3015_ (.RESET_B(net188),
    .D(_0122_),
    .Q(\p_acc[8] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3016_ (.RESET_B(net185),
    .D(_0123_),
    .Q(\p_acc[9] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3017_ (.RESET_B(net185),
    .D(_0124_),
    .Q(\p_acc[10] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3018_ (.RESET_B(net175),
    .D(_0125_),
    .Q(\p_acc[11] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3019_ (.RESET_B(net184),
    .D(_0126_),
    .Q(\p_acc[12] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3020_ (.RESET_B(net175),
    .D(_0127_),
    .Q(\p_acc[13] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3021_ (.RESET_B(net174),
    .D(_0128_),
    .Q(\p_acc[14] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3022_ (.RESET_B(net172),
    .D(net578),
    .Q(\p_acc[15] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3023_ (.RESET_B(net210),
    .D(net477),
    .Q(\p_freq[0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3024_ (.RESET_B(net205),
    .D(_0131_),
    .Q(\p_freq[1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3025_ (.RESET_B(net208),
    .D(_0132_),
    .Q(\p_freq[2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3026_ (.RESET_B(net210),
    .D(_0133_),
    .Q(\p_freq[3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3027_ (.RESET_B(net207),
    .D(_0134_),
    .Q(\p_freq[4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3028_ (.RESET_B(net212),
    .D(_0135_),
    .Q(\p_freq[5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3029_ (.RESET_B(net202),
    .D(net480),
    .Q(\p_freq[6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3030_ (.RESET_B(net209),
    .D(_0137_),
    .Q(\p_freq[7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3031_ (.RESET_B(net193),
    .D(_0138_),
    .Q(cur_gate),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3032_ (.RESET_B(net192),
    .D(net397),
    .Q(\p_waveform[1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3033_ (.RESET_B(net186),
    .D(net332),
    .Q(\p_waveform[2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3034_ (.RESET_B(net188),
    .D(net417),
    .Q(\p_waveform[3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3035_ (.RESET_B(net176),
    .D(_0142_),
    .Q(\p_waveform[4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3036_ (.RESET_B(net176),
    .D(_0143_),
    .Q(\p_waveform[5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3037_ (.RESET_B(net181),
    .D(_0144_),
    .Q(\p_waveform[6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3038_ (.RESET_B(net176),
    .D(_0145_),
    .Q(\p_waveform[7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3039_ (.RESET_B(net197),
    .D(net363),
    .Q(\p_pw[0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3040_ (.RESET_B(net204),
    .D(_0147_),
    .Q(\p_pw[1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3041_ (.RESET_B(net190),
    .D(net246),
    .Q(\p_pw[2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3042_ (.RESET_B(net186),
    .D(net441),
    .Q(\p_pw[3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3043_ (.RESET_B(net186),
    .D(_0150_),
    .Q(\p_pw[4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3044_ (.RESET_B(net186),
    .D(net493),
    .Q(\p_pw[5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3045_ (.RESET_B(net190),
    .D(_0152_),
    .Q(\p_pw[6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3046_ (.RESET_B(net186),
    .D(_0153_),
    .Q(\p_pw[7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3047_ (.RESET_B(net179),
    .D(_0154_),
    .Q(\p_env[0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3048_ (.RESET_B(net170),
    .D(_0155_),
    .Q(\p_env[1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3049_ (.RESET_B(net179),
    .D(_0156_),
    .Q(\p_env[2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3050_ (.RESET_B(net179),
    .D(_0157_),
    .Q(\p_env[3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3051_ (.RESET_B(net179),
    .D(_0158_),
    .Q(\p_env[4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3052_ (.RESET_B(net180),
    .D(_0159_),
    .Q(\p_env[5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3053_ (.RESET_B(net181),
    .D(_0160_),
    .Q(\p_env[6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3054_ (.RESET_B(net180),
    .D(_0161_),
    .Q(\p_env[7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3055_ (.RESET_B(net195),
    .D(_0162_),
    .Q(\p_ast[0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3056_ (.RESET_B(net193),
    .D(_0163_),
    .Q(\p_ast[1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3057_ (.RESET_B(net195),
    .D(net343),
    .Q(p_gate_latch),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3058_ (.RESET_B(net182),
    .D(_0165_),
    .Q(p_releasing),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3059_ (.RESET_B(net217),
    .D(net298),
    .Q(\p_attack[0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3060_ (.RESET_B(net212),
    .D(net253),
    .Q(\p_attack[1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3061_ (.RESET_B(net213),
    .D(net250),
    .Q(\p_attack[2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3062_ (.RESET_B(net212),
    .D(net256),
    .Q(\p_attack[3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3063_ (.RESET_B(net218),
    .D(net380),
    .Q(\p_attack[4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3064_ (.RESET_B(net217),
    .D(_0171_),
    .Q(\p_attack[5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3065_ (.RESET_B(net218),
    .D(_0172_),
    .Q(\p_attack[6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3066_ (.RESET_B(net214),
    .D(net585),
    .Q(\p_attack[7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3067_ (.RESET_B(net196),
    .D(_0174_),
    .Q(\p_sustain[0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3068_ (.RESET_B(net197),
    .D(_0175_),
    .Q(\p_sustain[1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3069_ (.RESET_B(net193),
    .D(_0176_),
    .Q(\p_sustain[2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3070_ (.RESET_B(net194),
    .D(_0177_),
    .Q(\p_sustain[3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3071_ (.RESET_B(net198),
    .D(_0178_),
    .Q(\p_sustain[4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3072_ (.RESET_B(net199),
    .D(_0179_),
    .Q(\p_sustain[5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3073_ (.RESET_B(net214),
    .D(_0180_),
    .Q(\p_sustain[6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3074_ (.RESET_B(net199),
    .D(_0181_),
    .Q(\p_sustain[7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3075_ (.RESET_B(net171),
    .D(_0182_),
    .Q(p_prev_msb_d),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3076_ (.RESET_B(net209),
    .D(_0183_),
    .Q(\freq[0][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3077_ (.RESET_B(net205),
    .D(_0184_),
    .Q(\freq[0][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3078_ (.RESET_B(net208),
    .D(_0185_),
    .Q(\freq[0][2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3079_ (.RESET_B(net207),
    .D(_0186_),
    .Q(\freq[0][3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3080_ (.RESET_B(net207),
    .D(_0187_),
    .Q(\freq[0][4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3081_ (.RESET_B(net212),
    .D(_0188_),
    .Q(\freq[0][5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3082_ (.RESET_B(net204),
    .D(_0189_),
    .Q(\freq[0][6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3083_ (.RESET_B(net209),
    .D(_0190_),
    .Q(\freq[0][7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3084_ (.RESET_B(net215),
    .D(_0191_),
    .Q(\freq[1][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3085_ (.RESET_B(net210),
    .D(_0192_),
    .Q(\freq[1][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3086_ (.RESET_B(net209),
    .D(_0193_),
    .Q(\freq[1][2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3087_ (.RESET_B(net210),
    .D(_0194_),
    .Q(\freq[1][3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3088_ (.RESET_B(net209),
    .D(_0195_),
    .Q(\freq[1][4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3089_ (.RESET_B(net212),
    .D(_0196_),
    .Q(\freq[1][5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3090_ (.RESET_B(net205),
    .D(_0197_),
    .Q(\freq[1][6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3091_ (.RESET_B(net211),
    .D(_0198_),
    .Q(\freq[1][7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3092_ (.RESET_B(net215),
    .D(_0199_),
    .Q(\freq[2][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3093_ (.RESET_B(net210),
    .D(_0200_),
    .Q(\freq[2][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3094_ (.RESET_B(net209),
    .D(_0201_),
    .Q(\freq[2][2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3095_ (.RESET_B(net209),
    .D(_0202_),
    .Q(\freq[2][3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3096_ (.RESET_B(net209),
    .D(_0203_),
    .Q(\freq[2][4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3097_ (.RESET_B(net212),
    .D(_0204_),
    .Q(\freq[2][5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3098_ (.RESET_B(net205),
    .D(_0205_),
    .Q(\freq[2][6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3099_ (.RESET_B(net211),
    .D(_0206_),
    .Q(\freq[2][7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3100_ (.RESET_B(net194),
    .D(_0207_),
    .Q(\waveform[0][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3101_ (.RESET_B(net190),
    .D(_0208_),
    .Q(\waveform[0][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3102_ (.RESET_B(net184),
    .D(net463),
    .Q(\waveform[0][2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3103_ (.RESET_B(net188),
    .D(_0210_),
    .Q(\waveform[0][3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3104_ (.RESET_B(net176),
    .D(_0211_),
    .Q(\waveform[0][4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3105_ (.RESET_B(net176),
    .D(net426),
    .Q(\waveform[0][5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3106_ (.RESET_B(net181),
    .D(_0213_),
    .Q(\waveform[0][6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3107_ (.RESET_B(net177),
    .D(_0214_),
    .Q(\waveform[0][7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3108_ (.RESET_B(net194),
    .D(_0215_),
    .Q(\waveform[1][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3109_ (.RESET_B(net190),
    .D(_0216_),
    .Q(\waveform[1][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3110_ (.RESET_B(net185),
    .D(_0217_),
    .Q(\waveform[1][2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3111_ (.RESET_B(net188),
    .D(_0218_),
    .Q(\waveform[1][3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3112_ (.RESET_B(net177),
    .D(_0219_),
    .Q(\waveform[1][4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3113_ (.RESET_B(net186),
    .D(_0220_),
    .Q(\waveform[1][5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3114_ (.RESET_B(net193),
    .D(_0221_),
    .Q(\waveform[1][6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3115_ (.RESET_B(net181),
    .D(net454),
    .Q(\waveform[1][7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3116_ (.RESET_B(net194),
    .D(_0223_),
    .Q(\waveform[2][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3117_ (.RESET_B(net204),
    .D(_0224_),
    .Q(\waveform[2][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3118_ (.RESET_B(net185),
    .D(_0225_),
    .Q(\waveform[2][2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3119_ (.RESET_B(net188),
    .D(_0226_),
    .Q(\waveform[2][3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3120_ (.RESET_B(net177),
    .D(_0227_),
    .Q(\waveform[2][4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3121_ (.RESET_B(net186),
    .D(_0228_),
    .Q(\waveform[2][5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3122_ (.RESET_B(net193),
    .D(_0229_),
    .Q(\waveform[2][6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3123_ (.RESET_B(net181),
    .D(_0230_),
    .Q(\waveform[2][7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3124_ (.RESET_B(net197),
    .D(_0231_),
    .Q(\pw_reg[0][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3125_ (.RESET_B(net204),
    .D(_0232_),
    .Q(\pw_reg[0][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3126_ (.RESET_B(net198),
    .D(_0233_),
    .Q(\pw_reg[0][2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3127_ (.RESET_B(net186),
    .D(_0234_),
    .Q(\pw_reg[0][3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3128_ (.RESET_B(net187),
    .D(_0235_),
    .Q(\pw_reg[0][4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3129_ (.RESET_B(net187),
    .D(_0236_),
    .Q(\pw_reg[0][5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3130_ (.RESET_B(net190),
    .D(_0237_),
    .Q(\pw_reg[0][6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3131_ (.RESET_B(net187),
    .D(_0238_),
    .Q(\pw_reg[0][7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3132_ (.RESET_B(net198),
    .D(net449),
    .Q(\pw_reg[1][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3133_ (.RESET_B(net204),
    .D(_0240_),
    .Q(\pw_reg[1][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3134_ (.RESET_B(net204),
    .D(_0241_),
    .Q(\pw_reg[1][2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3135_ (.RESET_B(net190),
    .D(_0242_),
    .Q(\pw_reg[1][3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3136_ (.RESET_B(net191),
    .D(_0243_),
    .Q(\pw_reg[1][4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3137_ (.RESET_B(net191),
    .D(_0244_),
    .Q(\pw_reg[1][5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3138_ (.RESET_B(net190),
    .D(_0245_),
    .Q(\pw_reg[1][6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3139_ (.RESET_B(net197),
    .D(_0246_),
    .Q(\pw_reg[1][7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3140_ (.RESET_B(net198),
    .D(_0247_),
    .Q(\pw_reg[2][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3141_ (.RESET_B(net204),
    .D(_0248_),
    .Q(\pw_reg[2][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3142_ (.RESET_B(net204),
    .D(_0249_),
    .Q(\pw_reg[2][2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3143_ (.RESET_B(net190),
    .D(_0250_),
    .Q(\pw_reg[2][3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3144_ (.RESET_B(net191),
    .D(net433),
    .Q(\pw_reg[2][4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3145_ (.RESET_B(net191),
    .D(_0252_),
    .Q(\pw_reg[2][5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3146_ (.RESET_B(net191),
    .D(_0253_),
    .Q(\pw_reg[2][6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3147_ (.RESET_B(net197),
    .D(_0254_),
    .Q(\pw_reg[2][7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3148_ (.RESET_B(net216),
    .D(_0255_),
    .Q(\attack_reg[0][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3149_ (.RESET_B(net213),
    .D(_0256_),
    .Q(\attack_reg[0][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3150_ (.RESET_B(net212),
    .D(_0257_),
    .Q(\attack_reg[0][2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3151_ (.RESET_B(net212),
    .D(_0258_),
    .Q(\attack_reg[0][3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3152_ (.RESET_B(net218),
    .D(_0259_),
    .Q(\attack_reg[0][4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3153_ (.RESET_B(net218),
    .D(_0260_),
    .Q(\attack_reg[0][5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3154_ (.RESET_B(net216),
    .D(_0261_),
    .Q(\attack_reg[0][6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3155_ (.RESET_B(net214),
    .D(_0262_),
    .Q(\attack_reg[0][7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3156_ (.RESET_B(net216),
    .D(_0263_),
    .Q(\attack_reg[1][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3157_ (.RESET_B(net215),
    .D(_0264_),
    .Q(\attack_reg[1][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3158_ (.RESET_B(net215),
    .D(_0265_),
    .Q(\attack_reg[1][2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3159_ (.RESET_B(net216),
    .D(_0266_),
    .Q(\attack_reg[1][3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3160_ (.RESET_B(net218),
    .D(_0267_),
    .Q(\attack_reg[1][4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3161_ (.RESET_B(net217),
    .D(_0268_),
    .Q(\attack_reg[1][5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3162_ (.RESET_B(net216),
    .D(_0269_),
    .Q(\attack_reg[1][6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3163_ (.RESET_B(net215),
    .D(_0270_),
    .Q(\attack_reg[1][7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3164_ (.RESET_B(net216),
    .D(_0271_),
    .Q(\attack_reg[2][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3165_ (.RESET_B(net215),
    .D(_0272_),
    .Q(\attack_reg[2][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3166_ (.RESET_B(net215),
    .D(_0273_),
    .Q(\attack_reg[2][2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3167_ (.RESET_B(net216),
    .D(_0274_),
    .Q(\attack_reg[2][3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3168_ (.RESET_B(net218),
    .D(_0275_),
    .Q(\attack_reg[2][4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3169_ (.RESET_B(net217),
    .D(net461),
    .Q(\attack_reg[2][5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3170_ (.RESET_B(net218),
    .D(_0277_),
    .Q(\attack_reg[2][6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3171_ (.RESET_B(net215),
    .D(_0278_),
    .Q(\attack_reg[2][7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3172_ (.RESET_B(net196),
    .D(_0279_),
    .Q(\sustain_reg[0][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3173_ (.RESET_B(net201),
    .D(_0280_),
    .Q(\sustain_reg[0][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3174_ (.RESET_B(net194),
    .D(_0281_),
    .Q(\sustain_reg[0][2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3175_ (.RESET_B(net194),
    .D(_0282_),
    .Q(\sustain_reg[0][3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3176_ (.RESET_B(net213),
    .D(_0283_),
    .Q(\sustain_reg[0][4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3177_ (.RESET_B(net199),
    .D(_0284_),
    .Q(\sustain_reg[0][5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3178_ (.RESET_B(net213),
    .D(net436),
    .Q(\sustain_reg[0][6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3179_ (.RESET_B(net200),
    .D(net438),
    .Q(\sustain_reg[0][7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3180_ (.RESET_B(net197),
    .D(_0287_),
    .Q(\sustain_reg[1][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3181_ (.RESET_B(net201),
    .D(_0288_),
    .Q(\sustain_reg[1][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3182_ (.RESET_B(net198),
    .D(_0289_),
    .Q(\sustain_reg[1][2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3183_ (.RESET_B(net197),
    .D(_0290_),
    .Q(\sustain_reg[1][3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3184_ (.RESET_B(net213),
    .D(_0291_),
    .Q(\sustain_reg[1][4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3185_ (.RESET_B(net199),
    .D(_0292_),
    .Q(\sustain_reg[1][5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3186_ (.RESET_B(net214),
    .D(_0293_),
    .Q(\sustain_reg[1][6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3187_ (.RESET_B(net200),
    .D(_0294_),
    .Q(\sustain_reg[1][7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3188_ (.RESET_B(net198),
    .D(_0295_),
    .Q(\sustain_reg[2][0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3189_ (.RESET_B(net201),
    .D(_0296_),
    .Q(\sustain_reg[2][1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3190_ (.RESET_B(net198),
    .D(_0297_),
    .Q(\sustain_reg[2][2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3191_ (.RESET_B(net197),
    .D(_0298_),
    .Q(\sustain_reg[2][3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3192_ (.RESET_B(net213),
    .D(_0299_),
    .Q(\sustain_reg[2][4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3193_ (.RESET_B(net199),
    .D(net423),
    .Q(\sustain_reg[2][5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3194_ (.RESET_B(net214),
    .D(_0301_),
    .Q(\sustain_reg[2][6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3195_ (.RESET_B(net200),
    .D(_0302_),
    .Q(\sustain_reg[2][7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3196_ (.RESET_B(net174),
    .D(net247),
    .Q(noise_clk_d),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3197_ (.RESET_B(net217),
    .D(net317),
    .Q(\adsr_pre_hi[1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3198_ (.RESET_B(net217),
    .D(net262),
    .Q(\adsr_pre_hi[2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3199_ (.RESET_B(net217),
    .D(_0017_),
    .Q(\adsr_pre_hi[3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3200_ (.RESET_B(net217),
    .D(net258),
    .Q(\adsr_pre_hi[4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3201_ (.RESET_B(net214),
    .D(_0019_),
    .Q(\adsr_pre_hi[5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3202_ (.RESET_B(net220),
    .D(net315),
    .Q(\adsr_pre_hi[6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3203_ (.RESET_B(net214),
    .D(_0021_),
    .Q(\adsr_pre_hi[7] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3204_ (.RESET_B(net214),
    .D(net307),
    .Q(\adsr_pre_hi[8] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3205_ (.RESET_B(net200),
    .D(net698),
    .Q(\adsr_pre_hi[9] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3206_ (.RESET_B(net200),
    .D(net280),
    .Q(\adsr_pre_hi[10] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3207_ (.RESET_B(net199),
    .D(net361),
    .Q(\adsr_pre_hi[11] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3208_ (.RESET_B(net199),
    .D(_0014_),
    .Q(\adsr_pre_hi[12] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3209_ (.RESET_B(net199),
    .D(net260),
    .Q(\adsr_pre_hi[13] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3210_ (.RESET_B(net167),
    .D(net700),
    .Q(\slot[0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3211_ (.RESET_B(net168),
    .D(_0001_),
    .Q(\slot[1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3212_ (.RESET_B(net168),
    .D(_0002_),
    .Q(\slot[2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3213_ (.RESET_B(net216),
    .D(net7),
    .Q(wr_en_d),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3214_ (.RESET_B(net189),
    .D(net731),
    .Q(pwm_out),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3215_ (.RESET_B(net164),
    .D(net669),
    .Q(\u_pwm.count[0] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3216_ (.RESET_B(net164),
    .D(net720),
    .Q(\u_pwm.count[1] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3217_ (.RESET_B(net164),
    .D(net366),
    .Q(\u_pwm.count[2] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3218_ (.RESET_B(net165),
    .D(net694),
    .Q(\u_pwm.count[3] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3219_ (.RESET_B(net165),
    .D(net716),
    .Q(\u_pwm.count[4] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3220_ (.RESET_B(net167),
    .D(_0009_),
    .Q(\u_pwm.count[5] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3221_ (.RESET_B(net167),
    .D(net630),
    .Q(\u_pwm.count[6] ),
    .CLK(clk));
 sg13g2_dfrbpq_1 _3222_ (.RESET_B(net168),
    .D(net696),
    .Q(\u_pwm.count[7] ),
    .CLK(clk));
 sg13g2_tielo tt_um_sid_222 (.L_LO(net222));
 sg13g2_tielo tt_um_sid_223 (.L_LO(net223));
 sg13g2_tielo tt_um_sid_224 (.L_LO(net224));
 sg13g2_tielo tt_um_sid_225 (.L_LO(net225));
 sg13g2_tielo tt_um_sid_226 (.L_LO(net226));
 sg13g2_tielo tt_um_sid_227 (.L_LO(net227));
 sg13g2_tielo tt_um_sid_228 (.L_LO(net228));
 sg13g2_tielo tt_um_sid_229 (.L_LO(net229));
 sg13g2_tielo tt_um_sid_230 (.L_LO(net230));
 sg13g2_tielo tt_um_sid_231 (.L_LO(net231));
 sg13g2_tielo tt_um_sid_232 (.L_LO(net232));
 sg13g2_tielo tt_um_sid_233 (.L_LO(net233));
 sg13g2_tielo tt_um_sid_234 (.L_LO(net234));
 sg13g2_tielo tt_um_sid_235 (.L_LO(net235));
 sg13g2_tielo tt_um_sid_236 (.L_LO(net236));
 sg13g2_tielo tt_um_sid_237 (.L_LO(net237));
 sg13g2_tielo tt_um_sid_238 (.L_LO(net238));
 sg13g2_tielo tt_um_sid_239 (.L_LO(net239));
 sg13g2_tielo tt_um_sid_240 (.L_LO(net240));
 sg13g2_tielo tt_um_sid_241 (.L_LO(net241));
 sg13g2_tielo tt_um_sid_242 (.L_LO(net242));
 sg13g2_tielo tt_um_sid_243 (.L_LO(net243));
 sg13g2_dlygate4sd3_1 hold244 (.A(\pw_reg[2][2] ),
    .X(net244));
 sg13g2_buf_1 _3246_ (.A(pwm_out),
    .X(uo_out[0]));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[7]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[0]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[1]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[2]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[3]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[4]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[5]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[6]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[7]),
    .X(net15));
 sg13g2_buf_1 fanout16 (.A(_0578_),
    .X(net16));
 sg13g2_buf_1 fanout17 (.A(_0530_),
    .X(net17));
 sg13g2_buf_1 fanout18 (.A(_0502_),
    .X(net18));
 sg13g2_buf_1 fanout19 (.A(_0478_),
    .X(net19));
 sg13g2_buf_1 fanout20 (.A(_0478_),
    .X(net20));
 sg13g2_buf_1 fanout21 (.A(_0466_),
    .X(net21));
 sg13g2_buf_1 fanout22 (.A(_0466_),
    .X(net22));
 sg13g2_buf_1 fanout23 (.A(_0447_),
    .X(net23));
 sg13g2_buf_1 fanout24 (.A(net25),
    .X(net24));
 sg13g2_buf_1 fanout25 (.A(_0441_),
    .X(net25));
 sg13g2_buf_1 fanout26 (.A(_0417_),
    .X(net26));
 sg13g2_buf_1 fanout27 (.A(_0417_),
    .X(net27));
 sg13g2_buf_1 fanout28 (.A(_1384_),
    .X(net28));
 sg13g2_buf_1 fanout29 (.A(_0546_),
    .X(net29));
 sg13g2_buf_1 fanout30 (.A(net31),
    .X(net30));
 sg13g2_buf_1 fanout31 (.A(_1378_),
    .X(net31));
 sg13g2_buf_1 fanout32 (.A(net33),
    .X(net32));
 sg13g2_buf_1 fanout33 (.A(_0387_),
    .X(net33));
 sg13g2_buf_1 fanout34 (.A(net35),
    .X(net34));
 sg13g2_buf_1 fanout35 (.A(net36),
    .X(net35));
 sg13g2_buf_1 fanout36 (.A(_1345_),
    .X(net36));
 sg13g2_buf_1 fanout37 (.A(net38),
    .X(net37));
 sg13g2_buf_1 fanout38 (.A(net49),
    .X(net38));
 sg13g2_buf_1 fanout39 (.A(net49),
    .X(net39));
 sg13g2_buf_1 fanout40 (.A(net49),
    .X(net40));
 sg13g2_buf_1 fanout41 (.A(net45),
    .X(net41));
 sg13g2_buf_1 fanout42 (.A(net45),
    .X(net42));
 sg13g2_buf_1 fanout43 (.A(net45),
    .X(net43));
 sg13g2_buf_1 fanout44 (.A(net45),
    .X(net44));
 sg13g2_buf_1 fanout45 (.A(net49),
    .X(net45));
 sg13g2_buf_1 fanout46 (.A(net48),
    .X(net46));
 sg13g2_buf_1 fanout47 (.A(net48),
    .X(net47));
 sg13g2_buf_1 fanout48 (.A(net49),
    .X(net48));
 sg13g2_buf_1 fanout49 (.A(_0904_),
    .X(net49));
 sg13g2_buf_1 fanout50 (.A(net54),
    .X(net50));
 sg13g2_buf_1 fanout51 (.A(net54),
    .X(net51));
 sg13g2_buf_1 fanout52 (.A(net54),
    .X(net52));
 sg13g2_buf_1 fanout53 (.A(net54),
    .X(net53));
 sg13g2_buf_1 fanout54 (.A(net55),
    .X(net54));
 sg13g2_buf_1 fanout55 (.A(net74),
    .X(net55));
 sg13g2_buf_1 fanout56 (.A(net57),
    .X(net56));
 sg13g2_buf_1 fanout57 (.A(net74),
    .X(net57));
 sg13g2_buf_1 fanout58 (.A(net60),
    .X(net58));
 sg13g2_buf_1 fanout59 (.A(net60),
    .X(net59));
 sg13g2_buf_1 fanout60 (.A(net74),
    .X(net60));
 sg13g2_buf_1 fanout61 (.A(net62),
    .X(net61));
 sg13g2_buf_1 fanout62 (.A(net67),
    .X(net62));
 sg13g2_buf_1 fanout63 (.A(net65),
    .X(net63));
 sg13g2_buf_1 fanout64 (.A(net65),
    .X(net64));
 sg13g2_buf_1 fanout65 (.A(net67),
    .X(net65));
 sg13g2_buf_1 fanout66 (.A(net67),
    .X(net66));
 sg13g2_buf_1 fanout67 (.A(net73),
    .X(net67));
 sg13g2_buf_1 fanout68 (.A(net73),
    .X(net68));
 sg13g2_buf_1 fanout69 (.A(net73),
    .X(net69));
 sg13g2_buf_1 fanout70 (.A(net72),
    .X(net70));
 sg13g2_buf_1 fanout71 (.A(net72),
    .X(net71));
 sg13g2_buf_1 fanout72 (.A(net73),
    .X(net72));
 sg13g2_buf_1 fanout73 (.A(net74),
    .X(net73));
 sg13g2_buf_1 fanout74 (.A(_0903_),
    .X(net74));
 sg13g2_buf_1 fanout75 (.A(net76),
    .X(net75));
 sg13g2_buf_1 fanout76 (.A(net94),
    .X(net76));
 sg13g2_buf_1 fanout77 (.A(net81),
    .X(net77));
 sg13g2_buf_1 fanout78 (.A(net81),
    .X(net78));
 sg13g2_buf_1 fanout79 (.A(net80),
    .X(net79));
 sg13g2_buf_1 fanout80 (.A(net81),
    .X(net80));
 sg13g2_buf_1 fanout81 (.A(net94),
    .X(net81));
 sg13g2_buf_1 fanout82 (.A(net84),
    .X(net82));
 sg13g2_buf_1 fanout83 (.A(net84),
    .X(net83));
 sg13g2_buf_1 fanout84 (.A(net94),
    .X(net84));
 sg13g2_buf_1 fanout85 (.A(net86),
    .X(net85));
 sg13g2_buf_1 fanout86 (.A(net94),
    .X(net86));
 sg13g2_buf_1 fanout87 (.A(net88),
    .X(net87));
 sg13g2_buf_1 fanout88 (.A(net93),
    .X(net88));
 sg13g2_buf_1 fanout89 (.A(net93),
    .X(net89));
 sg13g2_buf_1 fanout90 (.A(net93),
    .X(net90));
 sg13g2_buf_1 fanout91 (.A(net92),
    .X(net91));
 sg13g2_buf_1 fanout92 (.A(net93),
    .X(net92));
 sg13g2_buf_1 fanout93 (.A(net94),
    .X(net93));
 sg13g2_buf_1 fanout94 (.A(_0850_),
    .X(net94));
 sg13g2_buf_1 fanout95 (.A(net96),
    .X(net95));
 sg13g2_buf_1 fanout96 (.A(net102),
    .X(net96));
 sg13g2_buf_1 fanout97 (.A(net102),
    .X(net97));
 sg13g2_buf_1 fanout98 (.A(net102),
    .X(net98));
 sg13g2_buf_1 fanout99 (.A(net100),
    .X(net99));
 sg13g2_buf_1 fanout100 (.A(net101),
    .X(net100));
 sg13g2_buf_1 fanout101 (.A(net102),
    .X(net101));
 sg13g2_buf_1 fanout102 (.A(_0745_),
    .X(net102));
 sg13g2_buf_1 fanout103 (.A(net107),
    .X(net103));
 sg13g2_buf_1 fanout104 (.A(net107),
    .X(net104));
 sg13g2_buf_1 fanout105 (.A(net107),
    .X(net105));
 sg13g2_buf_1 fanout106 (.A(net107),
    .X(net106));
 sg13g2_buf_1 fanout107 (.A(net111),
    .X(net107));
 sg13g2_buf_1 fanout108 (.A(net109),
    .X(net108));
 sg13g2_buf_1 fanout109 (.A(net110),
    .X(net109));
 sg13g2_buf_1 fanout110 (.A(net111),
    .X(net110));
 sg13g2_buf_1 fanout111 (.A(_0744_),
    .X(net111));
 sg13g2_buf_1 fanout112 (.A(_1416_),
    .X(net112));
 sg13g2_buf_1 fanout113 (.A(net114),
    .X(net113));
 sg13g2_buf_1 fanout114 (.A(_1273_),
    .X(net114));
 sg13g2_buf_1 fanout115 (.A(_0995_),
    .X(net115));
 sg13g2_buf_1 fanout116 (.A(_0995_),
    .X(net116));
 sg13g2_buf_1 fanout117 (.A(net129),
    .X(net117));
 sg13g2_buf_1 fanout118 (.A(net119),
    .X(net118));
 sg13g2_buf_1 fanout119 (.A(net129),
    .X(net119));
 sg13g2_buf_1 fanout120 (.A(net123),
    .X(net120));
 sg13g2_buf_1 fanout121 (.A(net123),
    .X(net121));
 sg13g2_buf_1 fanout122 (.A(net123),
    .X(net122));
 sg13g2_buf_1 fanout123 (.A(net129),
    .X(net123));
 sg13g2_buf_1 fanout124 (.A(net128),
    .X(net124));
 sg13g2_buf_1 fanout125 (.A(net128),
    .X(net125));
 sg13g2_buf_1 fanout126 (.A(net128),
    .X(net126));
 sg13g2_buf_1 fanout127 (.A(net128),
    .X(net127));
 sg13g2_buf_1 fanout128 (.A(net129),
    .X(net128));
 sg13g2_buf_1 fanout129 (.A(_1272_),
    .X(net129));
 sg13g2_buf_1 fanout130 (.A(_1215_),
    .X(net130));
 sg13g2_buf_1 fanout131 (.A(net133),
    .X(net131));
 sg13g2_buf_1 fanout132 (.A(net133),
    .X(net132));
 sg13g2_buf_1 fanout133 (.A(net717),
    .X(net133));
 sg13g2_buf_1 fanout134 (.A(net135),
    .X(net134));
 sg13g2_buf_1 fanout135 (.A(net739),
    .X(net135));
 sg13g2_buf_1 fanout136 (.A(net687),
    .X(net136));
 sg13g2_buf_1 fanout137 (.A(net672),
    .X(net137));
 sg13g2_buf_1 fanout138 (.A(net681),
    .X(net138));
 sg13g2_buf_1 fanout139 (.A(net658),
    .X(net139));
 sg13g2_buf_1 fanout140 (.A(net673),
    .X(net140));
 sg13g2_buf_1 fanout141 (.A(net623),
    .X(net141));
 sg13g2_buf_1 fanout142 (.A(net651),
    .X(net142));
 sg13g2_buf_1 fanout143 (.A(net144),
    .X(net143));
 sg13g2_buf_1 fanout144 (.A(net145),
    .X(net144));
 sg13g2_buf_1 fanout145 (.A(net683),
    .X(net145));
 sg13g2_buf_1 fanout146 (.A(net690),
    .X(net146));
 sg13g2_buf_1 fanout147 (.A(net701),
    .X(net147));
 sg13g2_buf_1 fanout148 (.A(net149),
    .X(net148));
 sg13g2_buf_1 fanout149 (.A(net9),
    .X(net149));
 sg13g2_buf_1 fanout150 (.A(net151),
    .X(net150));
 sg13g2_buf_1 fanout151 (.A(net8),
    .X(net151));
 sg13g2_buf_1 fanout152 (.A(net15),
    .X(net152));
 sg13g2_buf_1 fanout153 (.A(net15),
    .X(net153));
 sg13g2_buf_1 fanout154 (.A(net155),
    .X(net154));
 sg13g2_buf_1 fanout155 (.A(net14),
    .X(net155));
 sg13g2_buf_1 fanout156 (.A(net157),
    .X(net156));
 sg13g2_buf_1 fanout157 (.A(net13),
    .X(net157));
 sg13g2_buf_1 fanout158 (.A(net159),
    .X(net158));
 sg13g2_buf_1 fanout159 (.A(net12),
    .X(net159));
 sg13g2_buf_1 fanout160 (.A(net161),
    .X(net160));
 sg13g2_buf_1 fanout161 (.A(net11),
    .X(net161));
 sg13g2_buf_1 fanout162 (.A(net10),
    .X(net162));
 sg13g2_buf_1 fanout163 (.A(net10),
    .X(net163));
 sg13g2_buf_1 fanout164 (.A(net166),
    .X(net164));
 sg13g2_buf_1 fanout165 (.A(net166),
    .X(net165));
 sg13g2_buf_1 fanout166 (.A(net170),
    .X(net166));
 sg13g2_buf_1 fanout167 (.A(net168),
    .X(net167));
 sg13g2_buf_1 fanout168 (.A(net170),
    .X(net168));
 sg13g2_buf_1 fanout169 (.A(net170),
    .X(net169));
 sg13g2_buf_1 fanout170 (.A(net1),
    .X(net170));
 sg13g2_buf_1 fanout171 (.A(net173),
    .X(net171));
 sg13g2_buf_1 fanout172 (.A(net173),
    .X(net172));
 sg13g2_buf_1 fanout173 (.A(net183),
    .X(net173));
 sg13g2_buf_1 fanout174 (.A(net177),
    .X(net174));
 sg13g2_buf_1 fanout175 (.A(net177),
    .X(net175));
 sg13g2_buf_1 fanout176 (.A(net177),
    .X(net176));
 sg13g2_buf_1 fanout177 (.A(net183),
    .X(net177));
 sg13g2_buf_1 fanout178 (.A(net183),
    .X(net178));
 sg13g2_buf_1 fanout179 (.A(net183),
    .X(net179));
 sg13g2_buf_1 fanout180 (.A(net182),
    .X(net180));
 sg13g2_buf_1 fanout181 (.A(net182),
    .X(net181));
 sg13g2_buf_1 fanout182 (.A(net183),
    .X(net182));
 sg13g2_buf_1 fanout183 (.A(net1),
    .X(net183));
 sg13g2_buf_1 fanout184 (.A(net187),
    .X(net184));
 sg13g2_buf_1 fanout185 (.A(net187),
    .X(net185));
 sg13g2_buf_1 fanout186 (.A(net187),
    .X(net186));
 sg13g2_buf_1 fanout187 (.A(net192),
    .X(net187));
 sg13g2_buf_1 fanout188 (.A(net189),
    .X(net188));
 sg13g2_buf_1 fanout189 (.A(net192),
    .X(net189));
 sg13g2_buf_1 fanout190 (.A(net191),
    .X(net190));
 sg13g2_buf_1 fanout191 (.A(net192),
    .X(net191));
 sg13g2_buf_1 fanout192 (.A(net221),
    .X(net192));
 sg13g2_buf_1 fanout193 (.A(net196),
    .X(net193));
 sg13g2_buf_1 fanout194 (.A(net196),
    .X(net194));
 sg13g2_buf_1 fanout195 (.A(net196),
    .X(net195));
 sg13g2_buf_1 fanout196 (.A(net221),
    .X(net196));
 sg13g2_buf_1 fanout197 (.A(net198),
    .X(net197));
 sg13g2_buf_1 fanout198 (.A(net201),
    .X(net198));
 sg13g2_buf_1 fanout199 (.A(net201),
    .X(net199));
 sg13g2_buf_1 fanout200 (.A(net201),
    .X(net200));
 sg13g2_buf_1 fanout201 (.A(net221),
    .X(net201));
 sg13g2_buf_1 fanout202 (.A(net206),
    .X(net202));
 sg13g2_buf_1 fanout203 (.A(net206),
    .X(net203));
 sg13g2_buf_1 fanout204 (.A(net206),
    .X(net204));
 sg13g2_buf_1 fanout205 (.A(net206),
    .X(net205));
 sg13g2_buf_1 fanout206 (.A(net221),
    .X(net206));
 sg13g2_buf_1 fanout207 (.A(net211),
    .X(net207));
 sg13g2_buf_1 fanout208 (.A(net211),
    .X(net208));
 sg13g2_buf_1 fanout209 (.A(net210),
    .X(net209));
 sg13g2_buf_1 fanout210 (.A(net211),
    .X(net210));
 sg13g2_buf_1 fanout211 (.A(net221),
    .X(net211));
 sg13g2_buf_1 fanout212 (.A(net213),
    .X(net212));
 sg13g2_buf_1 fanout213 (.A(net220),
    .X(net213));
 sg13g2_buf_1 fanout214 (.A(net220),
    .X(net214));
 sg13g2_buf_1 fanout215 (.A(net219),
    .X(net215));
 sg13g2_buf_1 fanout216 (.A(net219),
    .X(net216));
 sg13g2_buf_1 fanout217 (.A(net219),
    .X(net217));
 sg13g2_buf_1 fanout218 (.A(net219),
    .X(net218));
 sg13g2_buf_1 fanout219 (.A(net220),
    .X(net219));
 sg13g2_buf_1 fanout220 (.A(net221),
    .X(net220));
 sg13g2_buf_1 fanout221 (.A(net1),
    .X(net221));
 sg13g2_tielo tt_um_sid (.L_LO(net));
 sg13g2_dlygate4sd3_1 hold245 (.A(_1067_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0148_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold247 (.A(net732),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold248 (.A(\attack_reg[0][2] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold249 (.A(_1106_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0168_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold251 (.A(\attack_reg[0][1] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold252 (.A(_1104_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0167_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold254 (.A(\attack_reg[0][3] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold255 (.A(_1108_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0169_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold257 (.A(\adsr_pre_hi[4] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0018_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold259 (.A(\adsr_pre_hi[13] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0015_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold261 (.A(\adsr_pre_hi[2] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0016_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold263 (.A(\acc[2][5] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0966_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold265 (.A(_0049_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold266 (.A(\ast[2][1] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0988_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0089_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold269 (.A(\acc[2][9] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0970_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0053_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold272 (.A(\acc[2][6] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0967_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold274 (.A(_0050_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold275 (.A(\acc[2][2] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold276 (.A(_0963_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0046_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold278 (.A(\adsr_pre_hi[10] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold279 (.A(_1266_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0024_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold281 (.A(\acc[2][8] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0969_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0052_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold284 (.A(\acc[2][4] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0965_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0048_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold287 (.A(\acc[2][1] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0962_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0045_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold290 (.A(\acc[2][11] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold291 (.A(_0972_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0055_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold293 (.A(\acc[2][3] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold294 (.A(_0964_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0047_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold296 (.A(\attack_reg[2][0] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold297 (.A(_1103_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0166_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold299 (.A(\acc[2][13] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0974_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold301 (.A(_0057_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold302 (.A(\acc[2][0] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0961_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0044_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold305 (.A(\adsr_pre_hi[8] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold306 (.A(_1264_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold307 (.A(_0022_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold308 (.A(\acc[2][7] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0968_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold310 (.A(_0051_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold311 (.A(\mix_acc[8] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold312 (.A(_0896_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold313 (.A(_0311_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold314 (.A(\adsr_pre_hi[6] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold315 (.A(_0020_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold316 (.A(\adsr_pre_hi[1] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0012_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold318 (.A(\mix_acc[9] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold319 (.A(_0320_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold320 (.A(\acc[2][10] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold321 (.A(_0054_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold322 (.A(\acc[2][14] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold323 (.A(_0058_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold324 (.A(\gate_latch[2] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold325 (.A(\acc[2][12] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold326 (.A(_0056_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold327 (.A(\acc[0][7] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold328 (.A(_0328_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold329 (.A(\acc[0][5] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold330 (.A(_0326_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold331 (.A(\p_waveform[2] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold332 (.A(_0140_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold333 (.A(\acc[1][0] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold334 (.A(_0337_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold335 (.A(\mix_out[4] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold336 (.A(_0317_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold337 (.A(\acc[0][13] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold338 (.A(_0334_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold339 (.A(_0025_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0997_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold341 (.A(_0099_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold342 (.A(p_gate_latch),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold343 (.A(_0164_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold344 (.A(\acc[1][6] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold345 (.A(_0343_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold346 (.A(\acc[0][9] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold347 (.A(_0330_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold348 (.A(\acc[2][15] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold349 (.A(_0059_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold350 (.A(\acc[1][10] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold351 (.A(_0347_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold352 (.A(\prev_msb_d[0] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold353 (.A(_0096_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold354 (.A(\acc[0][3] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold355 (.A(_0324_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold356 (.A(\acc[0][6] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold357 (.A(_0327_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold358 (.A(\mix_acc[0] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold359 (.A(_0303_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold360 (.A(\adsr_pre_hi[11] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold361 (.A(_0013_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold362 (.A(\p_pw[0] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold363 (.A(_0146_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold364 (.A(\u_pwm.count[2] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold365 (.A(_1279_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold366 (.A(_0006_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold367 (.A(\acc[1][9] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold368 (.A(_0346_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold369 (.A(\mix_acc[7] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold370 (.A(_0897_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold371 (.A(_0899_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold372 (.A(\mix_out[0] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0313_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold374 (.A(\acc[1][7] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold375 (.A(_0344_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold376 (.A(\acc[0][2] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold377 (.A(_0323_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold378 (.A(\attack_reg[2][4] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold379 (.A(_1111_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold380 (.A(_0170_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold381 (.A(\gate_latch[0] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold382 (.A(\acc[0][14] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold383 (.A(_0335_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold384 (.A(\acc[1][2] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold385 (.A(_0339_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold386 (.A(\acc[1][1] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold387 (.A(_0338_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold388 (.A(\acc[1][5] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold389 (.A(_0342_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold390 (.A(\acc[1][14] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold391 (.A(_0042_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold392 (.A(\mix_out[2] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold393 (.A(_0315_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold394 (.A(\acc[0][12] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold395 (.A(_0333_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold396 (.A(\p_waveform[1] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold397 (.A(_0139_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold398 (.A(_0027_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0102_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold400 (.A(\acc[0][10] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0331_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold402 (.A(\adsr_pre_hi[3] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold403 (.A(\acc[0][1] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold404 (.A(_0322_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold405 (.A(_0026_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold406 (.A(_0100_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold407 (.A(\pw_reg[2][1] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold408 (.A(\env[2][4] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold409 (.A(net735),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold410 (.A(\acc[1][13] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold411 (.A(_0041_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold412 (.A(\acc[1][12] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold413 (.A(_0040_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold414 (.A(\acc[1][3] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold415 (.A(_0340_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold416 (.A(\p_waveform[3] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold417 (.A(_0141_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold418 (.A(_0031_),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold419 (.A(_0105_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold420 (.A(\env[2][2] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold421 (.A(\waveform[1][1] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold422 (.A(\sustain_reg[2][5] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0300_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold424 (.A(\env[1][6] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold425 (.A(\waveform[0][5] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold426 (.A(_0212_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold427 (.A(\env[2][3] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold428 (.A(_0079_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold429 (.A(\attack_reg[0][6] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold430 (.A(_0032_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold431 (.A(_0106_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold432 (.A(\pw_reg[2][4] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold433 (.A(_0251_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold434 (.A(\env[0][4] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold435 (.A(\sustain_reg[0][6] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold436 (.A(_0285_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold437 (.A(\sustain_reg[0][7] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold438 (.A(_0286_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold439 (.A(\pw_reg[2][3] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold440 (.A(_1069_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold441 (.A(_0149_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold442 (.A(\acc[1][8] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold443 (.A(_0345_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold444 (.A(\acc[1][4] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold445 (.A(_0341_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold446 (.A(\pw_reg[0][0] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold447 (.A(\env[2][0] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold448 (.A(\pw_reg[1][0] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold449 (.A(_0239_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold450 (.A(\attack_reg[0][5] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold451 (.A(\p_acc[4] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold452 (.A(_0118_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold453 (.A(\waveform[1][7] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold454 (.A(_0222_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold455 (.A(\freq[1][5] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold456 (.A(\pw_reg[0][7] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold457 (.A(\freq[2][3] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold458 (.A(\env[0][6] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold459 (.A(\attack_reg[1][5] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold460 (.A(\attack_reg[2][5] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold461 (.A(_0276_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold462 (.A(\waveform[0][2] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold463 (.A(_0209_),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold464 (.A(\acc[0][4] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold465 (.A(_0325_),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold466 (.A(\acc[0][8] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold467 (.A(_0329_),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold468 (.A(\env[1][4] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold469 (.A(\waveform[2][1] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold470 (.A(\freq[2][1] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold471 (.A(wr_en_d),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold472 (.A(\attack_reg[1][0] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold473 (.A(\sustain_reg[2][4] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold474 (.A(\sustain_reg[1][4] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold475 (.A(\gate_latch[1] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold476 (.A(\p_freq[0] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold477 (.A(_0130_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold478 (.A(\freq[1][1] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold479 (.A(\p_freq[6] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold480 (.A(_0136_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold481 (.A(noise_clk_d),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold482 (.A(\freq[0][2] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold483 (.A(\attack_reg[2][7] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold484 (.A(\pw_reg[0][1] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold485 (.A(\waveform[1][2] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold486 (.A(\pw_reg[0][2] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold487 (.A(\pw_reg[0][5] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold488 (.A(\freq[0][0] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold489 (.A(\freq[0][6] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold490 (.A(\sustain_reg[0][0] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold491 (.A(\freq[1][6] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold492 (.A(\p_pw[5] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold493 (.A(_0151_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold494 (.A(\attack_reg[1][3] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold495 (.A(\sustain_reg[2][6] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold496 (.A(\pw_reg[0][6] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold497 (.A(\pw_reg[1][5] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold498 (.A(\pw_reg[0][3] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold499 (.A(\attack_reg[1][1] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold500 (.A(\releasing[2] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold501 (.A(\prev_msb_d[2] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold502 (.A(\waveform[1][5] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold503 (.A(\env[1][3] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold504 (.A(_0071_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold505 (.A(\pw_reg[1][6] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold506 (.A(\sustain_reg[0][1] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold507 (.A(\ast[0][1] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold508 (.A(_0085_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold509 (.A(\freq[0][1] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold510 (.A(\freq[1][3] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold511 (.A(\waveform[2][3] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold512 (.A(\sustain_reg[2][2] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold513 (.A(\waveform[0][1] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold514 (.A(\sustain_reg[1][0] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold515 (.A(\attack_reg[2][3] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold516 (.A(\pw_reg[0][4] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold517 (.A(\waveform[0][7] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold518 (.A(\waveform[2][6] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold519 (.A(\mix_out[3] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold520 (.A(_0316_),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold521 (.A(\attack_reg[0][7] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold522 (.A(\acc[1][11] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold523 (.A(_0348_),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold524 (.A(\sustain_reg[1][3] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold525 (.A(\env[2][7] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold526 (.A(_0083_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold527 (.A(\attack_reg[2][6] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold528 (.A(\freq[2][5] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold529 (.A(\prev_msb_d[1] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold530 (.A(_0097_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold531 (.A(\ast[1][0] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold532 (.A(_0086_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold533 (.A(\waveform[0][6] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold534 (.A(\freq[1][0] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold535 (.A(\waveform[2][2] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold536 (.A(\waveform[2][4] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold537 (.A(\env[0][7] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold538 (.A(\mix_out[6] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold539 (.A(\attack_reg[0][0] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold540 (.A(\ast[1][1] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold541 (.A(_0087_),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold542 (.A(\p_acc[6] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold543 (.A(\env[1][5] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold544 (.A(\pw_reg[1][2] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold545 (.A(\freq[1][2] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold546 (.A(\attack_reg[1][6] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold547 (.A(\freq[2][0] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold548 (.A(\mix_out[5] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold549 (.A(\sustain_reg[2][3] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold550 (.A(\env[1][7] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold551 (.A(\attack_reg[1][4] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold552 (.A(\waveform[0][0] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold553 (.A(\waveform[1][0] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold554 (.A(\freq[0][5] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold555 (.A(\adsr_pre_hi[5] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold556 (.A(\waveform[2][5] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold557 (.A(\freq[2][7] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold558 (.A(\pw_reg[1][3] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold559 (.A(\pw_reg[2][5] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold560 (.A(\releasing[1] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold561 (.A(\freq[0][3] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold562 (.A(\freq[2][6] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold563 (.A(\attack_reg[0][4] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold564 (.A(\pw_reg[1][4] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold565 (.A(\p_pw[4] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold566 (.A(\pw_reg[2][0] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold567 (.A(\env[1][2] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold568 (.A(\sustain_reg[0][4] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold569 (.A(\env[0][5] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold570 (.A(_0029_),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold571 (.A(_0103_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold572 (.A(\pw_reg[2][7] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold573 (.A(\attack_reg[2][2] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold574 (.A(\env[2][1] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold575 (.A(_0077_),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold576 (.A(\freq[0][7] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold577 (.A(\p_acc[15] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold578 (.A(_0129_),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold579 (.A(\freq[2][2] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold580 (.A(\freq[1][7] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold581 (.A(\freq[1][4] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold582 (.A(\sustain_reg[2][7] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold583 (.A(\p_freq[2] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold584 (.A(\p_attack[7] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold585 (.A(_0173_),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold586 (.A(\releasing[0] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold587 (.A(\attack_reg[2][1] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold588 (.A(\env[1][0] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold589 (.A(\p_acc[7] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold590 (.A(\env[0][3] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold591 (.A(_0063_),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold592 (.A(\waveform[0][3] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold593 (.A(\waveform[2][0] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold594 (.A(\ast[0][0] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold595 (.A(_0084_),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold596 (.A(\pw_reg[1][1] ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold597 (.A(\waveform[2][7] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold598 (.A(\env[0][2] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold599 (.A(\p_attack[6] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold600 (.A(\sustain_reg[1][1] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold601 (.A(\p_acc[5] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold602 (.A(\env[1][1] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold603 (.A(_0069_),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold604 (.A(\p_freq[3] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold605 (.A(\sustain_reg[1][7] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold606 (.A(\sustain_reg[0][2] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold607 (.A(\freq[0][4] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold608 (.A(\sustain_reg[1][6] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold609 (.A(\p_sustain[6] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold610 (.A(\sustain_reg[0][3] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold611 (.A(\sustain_reg[2][0] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold612 (.A(\pw_reg[1][7] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold613 (.A(\waveform[1][4] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold614 (.A(\attack_reg[1][2] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold615 (.A(\pw_reg[2][6] ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold616 (.A(\ast[2][0] ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold617 (.A(_0088_),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold618 (.A(\p_acc[14] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold619 (.A(\freq[2][4] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold620 (.A(\env[0][0] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold621 (.A(\acc[0][0] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold622 (.A(_0321_),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold623 (.A(\p_env[0] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold624 (.A(\p_acc[2] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold625 (.A(\env[0][1] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold626 (.A(\p_acc[13] ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold627 (.A(\waveform[0][4] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold628 (.A(\u_pwm.count[6] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold629 (.A(_1287_),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold630 (.A(_0010_),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold631 (.A(\waveform[1][6] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold632 (.A(\p_env[3] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold633 (.A(\p_attack[5] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold634 (.A(\attack_reg[1][7] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold635 (.A(\sustain_reg[1][5] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold636 (.A(\waveform[1][3] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold637 (.A(\p_acc[3] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold638 (.A(\sustain_reg[1][2] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold639 (.A(_0030_),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold640 (.A(\p_sustain[7] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold641 (.A(\p_acc[10] ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold642 (.A(_1334_),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold643 (.A(_1359_),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold644 (.A(\sustain_reg[2][1] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold645 (.A(\p_pw[7] ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold646 (.A(\p_freq[4] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold647 (.A(\env[2][6] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold648 (.A(\p_acc[12] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold649 (.A(\p_acc[1] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold650 (.A(\sustain_reg[0][5] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold651 (.A(\p_waveform[7] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold652 (.A(\mix_out[1] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold653 (.A(_0314_),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold654 (.A(\p_freq[5] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold655 (.A(\p_acc[8] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold656 (.A(\p_acc[9] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold657 (.A(\p_pw[6] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold658 (.A(\p_env[2] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold659 (.A(\p_acc[11] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold660 (.A(\p_env[4] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold661 (.A(\p_acc[0] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold662 (.A(_0037_),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold663 (.A(_0111_),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold664 (.A(_0038_),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold665 (.A(\p_sustain[0] ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold666 (.A(_0035_),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold667 (.A(_0109_),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold668 (.A(\u_pwm.count[0] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold669 (.A(_0004_),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold670 (.A(\p_freq[1] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold671 (.A(\p_sustain[2] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold672 (.A(\p_env[6] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold673 (.A(\p_env[1] ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold674 (.A(_0036_),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold675 (.A(\acc[1][15] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold676 (.A(_0043_),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold677 (.A(\p_ast[0] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold678 (.A(\p_sustain[3] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold679 (.A(_0033_),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold680 (.A(_0034_),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold681 (.A(\p_env[5] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold682 (.A(\p_ast[1] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold683 (.A(\p_waveform[6] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold684 (.A(p_prev_msb_d),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold685 (.A(\p_freq[7] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold686 (.A(\p_pw[1] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold687 (.A(\p_env[7] ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold688 (.A(\mix_acc[1] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold689 (.A(_0304_),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold690 (.A(\p_waveform[5] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold691 (.A(\p_sustain[4] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold692 (.A(\u_pwm.count[3] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold693 (.A(_1280_),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold694 (.A(_0007_),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold695 (.A(\u_pwm.count[7] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold696 (.A(_0011_),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold697 (.A(\adsr_pre_hi[9] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold698 (.A(_0023_),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold699 (.A(\slot[0] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold700 (.A(_0000_),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold701 (.A(cur_gate),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold702 (.A(_0039_),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold703 (.A(\mix_acc[2] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold704 (.A(_0305_),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold705 (.A(\acc[0][15] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold706 (.A(_0336_),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold707 (.A(\adsr_pre_hi[7] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold708 (.A(\mix_acc[4] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold709 (.A(_0851_),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold710 (.A(_0307_),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold711 (.A(\p_sustain[1] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold712 (.A(\mix_acc[6] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold713 (.A(_0310_),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold714 (.A(\u_pwm.count[4] ),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold715 (.A(_1282_),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold716 (.A(_0008_),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold717 (.A(\slot[2] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold718 (.A(_0309_),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold719 (.A(\u_pwm.count[1] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold720 (.A(_0005_),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold721 (.A(\u_pwm.count[5] ),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold722 (.A(\adsr_pre_hi[12] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold723 (.A(_1268_),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold724 (.A(\mix_acc[3] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold725 (.A(_0306_),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold726 (.A(\p_sustain[5] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold727 (.A(\p_waveform[4] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold728 (.A(\mix_acc[5] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold729 (.A(\slot[1] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold730 (.A(\mix_out[7] ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold731 (.A(_0003_),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold732 (.A(\acc[0][11] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold733 (.A(\adsr_pre_hi[1] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold734 (.A(\mix_acc[5] ),
    .X(net734));
 sg13g2_antennanp ANTENNA_1 (.A(ui_in[1]));
 sg13g2_antennanp ANTENNA_2 (.A(ui_in[2]));
 sg13g2_dlygate4sd3_1 hold735 (.A(\env[2][5] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold736 (.A(_1089_),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold737 (.A(\p_sustain[1] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold738 (.A(\pw_reg[0][2] ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold739 (.A(p_releasing),
    .X(net739));
 sg13g2_antennanp ANTENNA_3 (.A(_1264_));
 sg13g2_antennanp ANTENNA_4 (.A(_1432_));
 sg13g2_antennanp ANTENNA_5 (.A(uio_in[1]));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_4 FILLER_0_413 ();
 sg13g2_fill_2 FILLER_0_417 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_4 FILLER_1_413 ();
 sg13g2_fill_2 FILLER_1_417 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_fill_1 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_155 ();
 sg13g2_decap_8 FILLER_2_162 ();
 sg13g2_decap_8 FILLER_2_169 ();
 sg13g2_fill_2 FILLER_2_176 ();
 sg13g2_decap_8 FILLER_2_181 ();
 sg13g2_decap_4 FILLER_2_188 ();
 sg13g2_fill_1 FILLER_2_192 ();
 sg13g2_decap_8 FILLER_2_198 ();
 sg13g2_decap_8 FILLER_2_205 ();
 sg13g2_fill_2 FILLER_2_212 ();
 sg13g2_decap_8 FILLER_2_219 ();
 sg13g2_decap_8 FILLER_2_226 ();
 sg13g2_decap_8 FILLER_2_233 ();
 sg13g2_decap_8 FILLER_2_240 ();
 sg13g2_decap_8 FILLER_2_247 ();
 sg13g2_decap_8 FILLER_2_254 ();
 sg13g2_decap_8 FILLER_2_261 ();
 sg13g2_decap_8 FILLER_2_268 ();
 sg13g2_decap_8 FILLER_2_275 ();
 sg13g2_decap_8 FILLER_2_282 ();
 sg13g2_decap_8 FILLER_2_289 ();
 sg13g2_decap_8 FILLER_2_296 ();
 sg13g2_decap_8 FILLER_2_303 ();
 sg13g2_decap_8 FILLER_2_310 ();
 sg13g2_decap_8 FILLER_2_317 ();
 sg13g2_decap_8 FILLER_2_324 ();
 sg13g2_decap_8 FILLER_2_331 ();
 sg13g2_decap_8 FILLER_2_338 ();
 sg13g2_decap_8 FILLER_2_345 ();
 sg13g2_decap_8 FILLER_2_352 ();
 sg13g2_decap_8 FILLER_2_359 ();
 sg13g2_decap_8 FILLER_2_366 ();
 sg13g2_decap_8 FILLER_2_373 ();
 sg13g2_decap_8 FILLER_2_380 ();
 sg13g2_decap_8 FILLER_2_387 ();
 sg13g2_decap_8 FILLER_2_394 ();
 sg13g2_decap_8 FILLER_2_401 ();
 sg13g2_decap_8 FILLER_2_408 ();
 sg13g2_decap_4 FILLER_2_415 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_4 FILLER_3_126 ();
 sg13g2_fill_2 FILLER_3_130 ();
 sg13g2_fill_1 FILLER_3_156 ();
 sg13g2_decap_4 FILLER_3_166 ();
 sg13g2_fill_2 FILLER_3_181 ();
 sg13g2_decap_4 FILLER_3_199 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_4 FILLER_3_413 ();
 sg13g2_fill_2 FILLER_3_417 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_fill_1 FILLER_4_112 ();
 sg13g2_fill_1 FILLER_4_122 ();
 sg13g2_fill_1 FILLER_4_135 ();
 sg13g2_fill_1 FILLER_4_191 ();
 sg13g2_decap_8 FILLER_4_247 ();
 sg13g2_decap_8 FILLER_4_254 ();
 sg13g2_decap_8 FILLER_4_261 ();
 sg13g2_decap_8 FILLER_4_268 ();
 sg13g2_decap_8 FILLER_4_275 ();
 sg13g2_decap_8 FILLER_4_282 ();
 sg13g2_decap_8 FILLER_4_289 ();
 sg13g2_decap_8 FILLER_4_296 ();
 sg13g2_decap_8 FILLER_4_303 ();
 sg13g2_decap_8 FILLER_4_310 ();
 sg13g2_decap_8 FILLER_4_317 ();
 sg13g2_decap_8 FILLER_4_324 ();
 sg13g2_decap_8 FILLER_4_331 ();
 sg13g2_decap_8 FILLER_4_338 ();
 sg13g2_decap_8 FILLER_4_345 ();
 sg13g2_decap_8 FILLER_4_352 ();
 sg13g2_decap_8 FILLER_4_359 ();
 sg13g2_decap_8 FILLER_4_366 ();
 sg13g2_decap_8 FILLER_4_373 ();
 sg13g2_decap_8 FILLER_4_380 ();
 sg13g2_decap_8 FILLER_4_387 ();
 sg13g2_decap_8 FILLER_4_394 ();
 sg13g2_decap_8 FILLER_4_401 ();
 sg13g2_decap_8 FILLER_4_408 ();
 sg13g2_decap_4 FILLER_4_415 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_4 FILLER_5_105 ();
 sg13g2_fill_1 FILLER_5_140 ();
 sg13g2_fill_2 FILLER_5_204 ();
 sg13g2_fill_2 FILLER_5_221 ();
 sg13g2_decap_8 FILLER_5_256 ();
 sg13g2_decap_8 FILLER_5_263 ();
 sg13g2_decap_8 FILLER_5_270 ();
 sg13g2_fill_2 FILLER_5_277 ();
 sg13g2_fill_1 FILLER_5_279 ();
 sg13g2_decap_8 FILLER_5_285 ();
 sg13g2_decap_8 FILLER_5_292 ();
 sg13g2_decap_8 FILLER_5_299 ();
 sg13g2_decap_8 FILLER_5_306 ();
 sg13g2_decap_8 FILLER_5_313 ();
 sg13g2_decap_8 FILLER_5_320 ();
 sg13g2_decap_8 FILLER_5_327 ();
 sg13g2_decap_8 FILLER_5_334 ();
 sg13g2_decap_8 FILLER_5_341 ();
 sg13g2_decap_8 FILLER_5_348 ();
 sg13g2_decap_8 FILLER_5_355 ();
 sg13g2_decap_8 FILLER_5_362 ();
 sg13g2_decap_8 FILLER_5_369 ();
 sg13g2_decap_8 FILLER_5_376 ();
 sg13g2_decap_8 FILLER_5_383 ();
 sg13g2_decap_8 FILLER_5_390 ();
 sg13g2_decap_8 FILLER_5_397 ();
 sg13g2_decap_8 FILLER_5_404 ();
 sg13g2_decap_8 FILLER_5_411 ();
 sg13g2_fill_1 FILLER_5_418 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_fill_2 FILLER_6_98 ();
 sg13g2_fill_1 FILLER_6_100 ();
 sg13g2_fill_1 FILLER_6_191 ();
 sg13g2_fill_2 FILLER_6_209 ();
 sg13g2_decap_8 FILLER_6_267 ();
 sg13g2_fill_1 FILLER_6_274 ();
 sg13g2_decap_8 FILLER_6_295 ();
 sg13g2_decap_8 FILLER_6_302 ();
 sg13g2_decap_8 FILLER_6_309 ();
 sg13g2_decap_8 FILLER_6_316 ();
 sg13g2_decap_8 FILLER_6_323 ();
 sg13g2_decap_8 FILLER_6_330 ();
 sg13g2_decap_8 FILLER_6_337 ();
 sg13g2_decap_8 FILLER_6_344 ();
 sg13g2_decap_8 FILLER_6_351 ();
 sg13g2_decap_8 FILLER_6_358 ();
 sg13g2_decap_8 FILLER_6_365 ();
 sg13g2_decap_8 FILLER_6_372 ();
 sg13g2_decap_8 FILLER_6_379 ();
 sg13g2_decap_8 FILLER_6_386 ();
 sg13g2_decap_8 FILLER_6_393 ();
 sg13g2_decap_8 FILLER_6_400 ();
 sg13g2_decap_8 FILLER_6_407 ();
 sg13g2_decap_4 FILLER_6_414 ();
 sg13g2_fill_1 FILLER_6_418 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_4 FILLER_7_91 ();
 sg13g2_fill_1 FILLER_7_208 ();
 sg13g2_fill_2 FILLER_7_252 ();
 sg13g2_fill_1 FILLER_7_254 ();
 sg13g2_fill_1 FILLER_7_263 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_4 FILLER_7_413 ();
 sg13g2_fill_2 FILLER_7_417 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_fill_1 FILLER_8_98 ();
 sg13g2_fill_2 FILLER_8_140 ();
 sg13g2_fill_2 FILLER_8_156 ();
 sg13g2_fill_2 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_237 ();
 sg13g2_decap_4 FILLER_8_244 ();
 sg13g2_fill_1 FILLER_8_248 ();
 sg13g2_decap_8 FILLER_8_298 ();
 sg13g2_decap_8 FILLER_8_305 ();
 sg13g2_decap_8 FILLER_8_312 ();
 sg13g2_decap_8 FILLER_8_319 ();
 sg13g2_decap_8 FILLER_8_326 ();
 sg13g2_decap_8 FILLER_8_333 ();
 sg13g2_decap_8 FILLER_8_340 ();
 sg13g2_decap_8 FILLER_8_347 ();
 sg13g2_decap_8 FILLER_8_354 ();
 sg13g2_decap_8 FILLER_8_361 ();
 sg13g2_decap_8 FILLER_8_368 ();
 sg13g2_decap_8 FILLER_8_375 ();
 sg13g2_decap_8 FILLER_8_382 ();
 sg13g2_decap_8 FILLER_8_389 ();
 sg13g2_decap_8 FILLER_8_396 ();
 sg13g2_decap_8 FILLER_8_403 ();
 sg13g2_decap_8 FILLER_8_410 ();
 sg13g2_fill_2 FILLER_8_417 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_fill_1 FILLER_9_120 ();
 sg13g2_fill_1 FILLER_9_151 ();
 sg13g2_fill_1 FILLER_9_235 ();
 sg13g2_fill_2 FILLER_9_249 ();
 sg13g2_fill_1 FILLER_9_251 ();
 sg13g2_decap_8 FILLER_9_260 ();
 sg13g2_decap_8 FILLER_9_267 ();
 sg13g2_decap_4 FILLER_9_274 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_4 FILLER_9_413 ();
 sg13g2_fill_2 FILLER_9_417 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_4 FILLER_10_98 ();
 sg13g2_fill_1 FILLER_10_102 ();
 sg13g2_fill_1 FILLER_10_217 ();
 sg13g2_fill_1 FILLER_10_241 ();
 sg13g2_fill_1 FILLER_10_260 ();
 sg13g2_decap_4 FILLER_10_269 ();
 sg13g2_fill_1 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_278 ();
 sg13g2_decap_4 FILLER_10_285 ();
 sg13g2_fill_2 FILLER_10_299 ();
 sg13g2_decap_8 FILLER_10_306 ();
 sg13g2_decap_8 FILLER_10_313 ();
 sg13g2_decap_8 FILLER_10_320 ();
 sg13g2_decap_8 FILLER_10_327 ();
 sg13g2_decap_8 FILLER_10_334 ();
 sg13g2_decap_8 FILLER_10_341 ();
 sg13g2_decap_8 FILLER_10_348 ();
 sg13g2_decap_8 FILLER_10_355 ();
 sg13g2_decap_8 FILLER_10_362 ();
 sg13g2_decap_8 FILLER_10_369 ();
 sg13g2_decap_8 FILLER_10_376 ();
 sg13g2_decap_8 FILLER_10_383 ();
 sg13g2_decap_8 FILLER_10_390 ();
 sg13g2_decap_8 FILLER_10_397 ();
 sg13g2_decap_8 FILLER_10_404 ();
 sg13g2_decap_8 FILLER_10_411 ();
 sg13g2_fill_1 FILLER_10_418 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_4 FILLER_11_91 ();
 sg13g2_fill_2 FILLER_11_95 ();
 sg13g2_fill_1 FILLER_11_124 ();
 sg13g2_fill_1 FILLER_11_178 ();
 sg13g2_fill_2 FILLER_11_196 ();
 sg13g2_decap_4 FILLER_11_207 ();
 sg13g2_fill_1 FILLER_11_211 ();
 sg13g2_decap_8 FILLER_11_215 ();
 sg13g2_fill_2 FILLER_11_248 ();
 sg13g2_fill_1 FILLER_11_250 ();
 sg13g2_fill_2 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_316 ();
 sg13g2_decap_8 FILLER_11_323 ();
 sg13g2_decap_8 FILLER_11_330 ();
 sg13g2_decap_8 FILLER_11_337 ();
 sg13g2_decap_8 FILLER_11_344 ();
 sg13g2_decap_8 FILLER_11_351 ();
 sg13g2_decap_8 FILLER_11_358 ();
 sg13g2_decap_8 FILLER_11_365 ();
 sg13g2_decap_8 FILLER_11_372 ();
 sg13g2_decap_8 FILLER_11_379 ();
 sg13g2_decap_8 FILLER_11_386 ();
 sg13g2_decap_8 FILLER_11_393 ();
 sg13g2_decap_8 FILLER_11_400 ();
 sg13g2_decap_8 FILLER_11_407 ();
 sg13g2_decap_4 FILLER_11_414 ();
 sg13g2_fill_1 FILLER_11_418 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_4 FILLER_12_98 ();
 sg13g2_fill_1 FILLER_12_102 ();
 sg13g2_fill_1 FILLER_12_187 ();
 sg13g2_decap_8 FILLER_12_199 ();
 sg13g2_fill_1 FILLER_12_215 ();
 sg13g2_decap_4 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_236 ();
 sg13g2_decap_4 FILLER_12_243 ();
 sg13g2_fill_1 FILLER_12_270 ();
 sg13g2_fill_2 FILLER_12_299 ();
 sg13g2_fill_1 FILLER_12_301 ();
 sg13g2_fill_2 FILLER_12_307 ();
 sg13g2_fill_1 FILLER_12_309 ();
 sg13g2_decap_8 FILLER_12_314 ();
 sg13g2_decap_8 FILLER_12_321 ();
 sg13g2_decap_8 FILLER_12_328 ();
 sg13g2_decap_8 FILLER_12_335 ();
 sg13g2_decap_8 FILLER_12_342 ();
 sg13g2_decap_8 FILLER_12_349 ();
 sg13g2_decap_8 FILLER_12_356 ();
 sg13g2_decap_8 FILLER_12_363 ();
 sg13g2_decap_8 FILLER_12_370 ();
 sg13g2_decap_8 FILLER_12_377 ();
 sg13g2_decap_8 FILLER_12_384 ();
 sg13g2_decap_8 FILLER_12_391 ();
 sg13g2_decap_8 FILLER_12_398 ();
 sg13g2_decap_8 FILLER_12_405 ();
 sg13g2_decap_8 FILLER_12_412 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_4 FILLER_13_98 ();
 sg13g2_fill_2 FILLER_13_102 ();
 sg13g2_fill_1 FILLER_13_146 ();
 sg13g2_fill_2 FILLER_13_152 ();
 sg13g2_fill_1 FILLER_13_225 ();
 sg13g2_decap_4 FILLER_13_231 ();
 sg13g2_fill_1 FILLER_13_235 ();
 sg13g2_fill_2 FILLER_13_249 ();
 sg13g2_fill_1 FILLER_13_251 ();
 sg13g2_decap_8 FILLER_13_256 ();
 sg13g2_decap_8 FILLER_13_263 ();
 sg13g2_fill_2 FILLER_13_275 ();
 sg13g2_fill_2 FILLER_13_289 ();
 sg13g2_fill_1 FILLER_13_291 ();
 sg13g2_fill_1 FILLER_13_305 ();
 sg13g2_decap_8 FILLER_13_319 ();
 sg13g2_decap_8 FILLER_13_326 ();
 sg13g2_decap_8 FILLER_13_333 ();
 sg13g2_decap_8 FILLER_13_340 ();
 sg13g2_decap_8 FILLER_13_347 ();
 sg13g2_decap_8 FILLER_13_354 ();
 sg13g2_decap_8 FILLER_13_361 ();
 sg13g2_decap_8 FILLER_13_368 ();
 sg13g2_decap_8 FILLER_13_375 ();
 sg13g2_decap_8 FILLER_13_382 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_decap_8 FILLER_13_403 ();
 sg13g2_decap_8 FILLER_13_410 ();
 sg13g2_fill_2 FILLER_13_417 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_4 FILLER_14_98 ();
 sg13g2_fill_1 FILLER_14_141 ();
 sg13g2_fill_1 FILLER_14_148 ();
 sg13g2_fill_2 FILLER_14_159 ();
 sg13g2_fill_2 FILLER_14_222 ();
 sg13g2_fill_1 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_229 ();
 sg13g2_fill_2 FILLER_14_236 ();
 sg13g2_fill_1 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_251 ();
 sg13g2_decap_8 FILLER_14_258 ();
 sg13g2_fill_1 FILLER_14_265 ();
 sg13g2_decap_4 FILLER_14_270 ();
 sg13g2_fill_2 FILLER_14_274 ();
 sg13g2_fill_2 FILLER_14_284 ();
 sg13g2_fill_1 FILLER_14_286 ();
 sg13g2_decap_8 FILLER_14_300 ();
 sg13g2_fill_1 FILLER_14_311 ();
 sg13g2_decap_8 FILLER_14_320 ();
 sg13g2_decap_8 FILLER_14_327 ();
 sg13g2_decap_8 FILLER_14_334 ();
 sg13g2_decap_8 FILLER_14_341 ();
 sg13g2_decap_8 FILLER_14_348 ();
 sg13g2_decap_8 FILLER_14_355 ();
 sg13g2_decap_8 FILLER_14_362 ();
 sg13g2_decap_8 FILLER_14_369 ();
 sg13g2_decap_8 FILLER_14_376 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_8 FILLER_14_404 ();
 sg13g2_decap_8 FILLER_14_411 ();
 sg13g2_fill_1 FILLER_14_418 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_fill_2 FILLER_15_91 ();
 sg13g2_fill_2 FILLER_15_196 ();
 sg13g2_fill_1 FILLER_15_213 ();
 sg13g2_decap_4 FILLER_15_234 ();
 sg13g2_fill_1 FILLER_15_238 ();
 sg13g2_fill_1 FILLER_15_243 ();
 sg13g2_fill_2 FILLER_15_265 ();
 sg13g2_fill_1 FILLER_15_267 ();
 sg13g2_fill_1 FILLER_15_276 ();
 sg13g2_fill_1 FILLER_15_290 ();
 sg13g2_decap_8 FILLER_15_327 ();
 sg13g2_decap_8 FILLER_15_334 ();
 sg13g2_decap_4 FILLER_15_341 ();
 sg13g2_fill_1 FILLER_15_345 ();
 sg13g2_decap_4 FILLER_15_356 ();
 sg13g2_fill_1 FILLER_15_360 ();
 sg13g2_decap_8 FILLER_15_370 ();
 sg13g2_decap_8 FILLER_15_377 ();
 sg13g2_decap_8 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_8 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_15_412 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_fill_2 FILLER_16_91 ();
 sg13g2_fill_2 FILLER_16_139 ();
 sg13g2_fill_2 FILLER_16_213 ();
 sg13g2_fill_1 FILLER_16_215 ();
 sg13g2_fill_1 FILLER_16_220 ();
 sg13g2_fill_2 FILLER_16_239 ();
 sg13g2_fill_1 FILLER_16_294 ();
 sg13g2_decap_4 FILLER_16_332 ();
 sg13g2_decap_8 FILLER_16_389 ();
 sg13g2_decap_8 FILLER_16_396 ();
 sg13g2_decap_8 FILLER_16_403 ();
 sg13g2_decap_8 FILLER_16_410 ();
 sg13g2_fill_2 FILLER_16_417 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_fill_2 FILLER_17_98 ();
 sg13g2_fill_2 FILLER_17_192 ();
 sg13g2_fill_1 FILLER_17_216 ();
 sg13g2_fill_2 FILLER_17_225 ();
 sg13g2_fill_1 FILLER_17_240 ();
 sg13g2_fill_2 FILLER_17_278 ();
 sg13g2_fill_1 FILLER_17_280 ();
 sg13g2_fill_2 FILLER_17_285 ();
 sg13g2_fill_1 FILLER_17_287 ();
 sg13g2_fill_2 FILLER_17_309 ();
 sg13g2_fill_1 FILLER_17_311 ();
 sg13g2_fill_2 FILLER_17_320 ();
 sg13g2_fill_1 FILLER_17_322 ();
 sg13g2_fill_1 FILLER_17_337 ();
 sg13g2_fill_2 FILLER_17_357 ();
 sg13g2_fill_1 FILLER_17_359 ();
 sg13g2_decap_8 FILLER_17_397 ();
 sg13g2_decap_8 FILLER_17_404 ();
 sg13g2_decap_8 FILLER_17_411 ();
 sg13g2_fill_1 FILLER_17_418 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_4 FILLER_18_105 ();
 sg13g2_fill_2 FILLER_18_154 ();
 sg13g2_fill_2 FILLER_18_222 ();
 sg13g2_fill_1 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_253 ();
 sg13g2_decap_8 FILLER_18_260 ();
 sg13g2_fill_2 FILLER_18_267 ();
 sg13g2_fill_2 FILLER_18_297 ();
 sg13g2_fill_2 FILLER_18_303 ();
 sg13g2_decap_8 FILLER_18_400 ();
 sg13g2_decap_8 FILLER_18_407 ();
 sg13g2_decap_4 FILLER_18_414 ();
 sg13g2_fill_1 FILLER_18_418 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_4 FILLER_19_112 ();
 sg13g2_fill_1 FILLER_19_116 ();
 sg13g2_fill_1 FILLER_19_153 ();
 sg13g2_fill_1 FILLER_19_198 ();
 sg13g2_fill_1 FILLER_19_203 ();
 sg13g2_fill_2 FILLER_19_214 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_fill_1 FILLER_19_252 ();
 sg13g2_fill_2 FILLER_19_257 ();
 sg13g2_fill_1 FILLER_19_259 ();
 sg13g2_fill_1 FILLER_19_264 ();
 sg13g2_fill_2 FILLER_19_283 ();
 sg13g2_fill_1 FILLER_19_303 ();
 sg13g2_decap_8 FILLER_19_412 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_fill_1 FILLER_20_112 ();
 sg13g2_fill_2 FILLER_20_143 ();
 sg13g2_fill_2 FILLER_20_172 ();
 sg13g2_fill_2 FILLER_20_203 ();
 sg13g2_fill_1 FILLER_20_205 ();
 sg13g2_fill_2 FILLER_20_228 ();
 sg13g2_fill_2 FILLER_20_235 ();
 sg13g2_fill_2 FILLER_20_250 ();
 sg13g2_fill_2 FILLER_20_266 ();
 sg13g2_fill_2 FILLER_20_273 ();
 sg13g2_fill_1 FILLER_20_275 ();
 sg13g2_fill_2 FILLER_20_299 ();
 sg13g2_fill_1 FILLER_20_301 ();
 sg13g2_fill_2 FILLER_20_312 ();
 sg13g2_decap_4 FILLER_20_413 ();
 sg13g2_fill_2 FILLER_20_417 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_fill_1 FILLER_21_112 ();
 sg13g2_fill_1 FILLER_21_164 ();
 sg13g2_fill_1 FILLER_21_177 ();
 sg13g2_fill_2 FILLER_21_233 ();
 sg13g2_fill_2 FILLER_21_251 ();
 sg13g2_fill_1 FILLER_21_253 ();
 sg13g2_fill_1 FILLER_21_278 ();
 sg13g2_fill_2 FILLER_21_290 ();
 sg13g2_fill_1 FILLER_21_292 ();
 sg13g2_fill_2 FILLER_21_309 ();
 sg13g2_fill_1 FILLER_21_311 ();
 sg13g2_decap_8 FILLER_21_406 ();
 sg13g2_decap_4 FILLER_21_413 ();
 sg13g2_fill_2 FILLER_21_417 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_4 FILLER_22_105 ();
 sg13g2_fill_2 FILLER_22_109 ();
 sg13g2_fill_2 FILLER_22_141 ();
 sg13g2_fill_1 FILLER_22_295 ();
 sg13g2_fill_2 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_411 ();
 sg13g2_fill_1 FILLER_22_418 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_fill_1 FILLER_23_119 ();
 sg13g2_fill_1 FILLER_23_260 ();
 sg13g2_decap_4 FILLER_23_266 ();
 sg13g2_decap_4 FILLER_23_275 ();
 sg13g2_fill_1 FILLER_23_300 ();
 sg13g2_fill_2 FILLER_23_369 ();
 sg13g2_decap_8 FILLER_23_407 ();
 sg13g2_decap_4 FILLER_23_414 ();
 sg13g2_fill_1 FILLER_23_418 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_fill_2 FILLER_24_112 ();
 sg13g2_fill_1 FILLER_24_114 ();
 sg13g2_fill_1 FILLER_24_174 ();
 sg13g2_fill_1 FILLER_24_246 ();
 sg13g2_decap_8 FILLER_24_260 ();
 sg13g2_decap_4 FILLER_24_267 ();
 sg13g2_fill_2 FILLER_24_271 ();
 sg13g2_fill_2 FILLER_24_299 ();
 sg13g2_fill_1 FILLER_24_369 ();
 sg13g2_decap_8 FILLER_24_407 ();
 sg13g2_decap_4 FILLER_24_414 ();
 sg13g2_fill_1 FILLER_24_418 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_fill_2 FILLER_25_105 ();
 sg13g2_fill_1 FILLER_25_107 ();
 sg13g2_fill_2 FILLER_25_181 ();
 sg13g2_fill_1 FILLER_25_220 ();
 sg13g2_fill_2 FILLER_25_230 ();
 sg13g2_fill_1 FILLER_25_264 ();
 sg13g2_decap_4 FILLER_25_269 ();
 sg13g2_fill_1 FILLER_25_303 ();
 sg13g2_decap_8 FILLER_25_408 ();
 sg13g2_decap_4 FILLER_25_415 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_fill_1 FILLER_26_134 ();
 sg13g2_fill_2 FILLER_26_199 ();
 sg13g2_fill_2 FILLER_26_238 ();
 sg13g2_fill_1 FILLER_26_286 ();
 sg13g2_fill_2 FILLER_26_292 ();
 sg13g2_fill_1 FILLER_26_310 ();
 sg13g2_fill_1 FILLER_26_321 ();
 sg13g2_fill_1 FILLER_26_342 ();
 sg13g2_fill_1 FILLER_26_380 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_8 FILLER_26_403 ();
 sg13g2_decap_8 FILLER_26_410 ();
 sg13g2_fill_2 FILLER_26_417 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_4 FILLER_27_105 ();
 sg13g2_fill_2 FILLER_27_109 ();
 sg13g2_fill_2 FILLER_27_192 ();
 sg13g2_fill_1 FILLER_27_236 ();
 sg13g2_fill_2 FILLER_27_247 ();
 sg13g2_fill_2 FILLER_27_310 ();
 sg13g2_fill_1 FILLER_27_312 ();
 sg13g2_fill_2 FILLER_27_334 ();
 sg13g2_fill_2 FILLER_27_351 ();
 sg13g2_fill_2 FILLER_27_360 ();
 sg13g2_fill_1 FILLER_27_385 ();
 sg13g2_decap_4 FILLER_27_413 ();
 sg13g2_fill_2 FILLER_27_417 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_fill_1 FILLER_28_187 ();
 sg13g2_fill_2 FILLER_28_297 ();
 sg13g2_decap_8 FILLER_28_406 ();
 sg13g2_decap_4 FILLER_28_413 ();
 sg13g2_fill_2 FILLER_28_417 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_fill_2 FILLER_29_161 ();
 sg13g2_fill_1 FILLER_29_190 ();
 sg13g2_fill_1 FILLER_29_274 ();
 sg13g2_fill_1 FILLER_29_330 ();
 sg13g2_fill_1 FILLER_29_379 ();
 sg13g2_fill_2 FILLER_29_390 ();
 sg13g2_decap_8 FILLER_29_410 ();
 sg13g2_fill_2 FILLER_29_417 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_4 FILLER_30_98 ();
 sg13g2_fill_2 FILLER_30_102 ();
 sg13g2_fill_2 FILLER_30_194 ();
 sg13g2_fill_2 FILLER_30_253 ();
 sg13g2_fill_2 FILLER_30_264 ();
 sg13g2_fill_2 FILLER_30_389 ();
 sg13g2_fill_1 FILLER_30_391 ();
 sg13g2_decap_8 FILLER_30_404 ();
 sg13g2_decap_8 FILLER_30_411 ();
 sg13g2_fill_1 FILLER_30_418 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_fill_1 FILLER_31_98 ();
 sg13g2_fill_1 FILLER_31_126 ();
 sg13g2_fill_1 FILLER_31_142 ();
 sg13g2_fill_2 FILLER_31_189 ();
 sg13g2_fill_1 FILLER_31_255 ();
 sg13g2_fill_2 FILLER_31_308 ();
 sg13g2_fill_2 FILLER_31_315 ();
 sg13g2_fill_2 FILLER_31_396 ();
 sg13g2_decap_8 FILLER_31_410 ();
 sg13g2_fill_2 FILLER_31_417 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_fill_2 FILLER_32_98 ();
 sg13g2_fill_1 FILLER_32_100 ();
 sg13g2_fill_2 FILLER_32_153 ();
 sg13g2_fill_2 FILLER_32_291 ();
 sg13g2_fill_1 FILLER_32_293 ();
 sg13g2_fill_2 FILLER_32_321 ();
 sg13g2_fill_1 FILLER_32_362 ();
 sg13g2_fill_2 FILLER_32_402 ();
 sg13g2_fill_1 FILLER_32_404 ();
 sg13g2_fill_2 FILLER_32_417 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_fill_2 FILLER_33_91 ();
 sg13g2_fill_1 FILLER_33_93 ();
 sg13g2_fill_1 FILLER_33_225 ();
 sg13g2_fill_1 FILLER_33_255 ();
 sg13g2_fill_2 FILLER_33_266 ();
 sg13g2_fill_1 FILLER_33_337 ();
 sg13g2_fill_2 FILLER_33_385 ();
 sg13g2_fill_1 FILLER_33_387 ();
 sg13g2_fill_2 FILLER_33_416 ();
 sg13g2_fill_1 FILLER_33_418 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_4 FILLER_34_91 ();
 sg13g2_fill_2 FILLER_34_95 ();
 sg13g2_fill_1 FILLER_34_244 ();
 sg13g2_fill_2 FILLER_34_359 ();
 sg13g2_fill_2 FILLER_34_380 ();
 sg13g2_fill_1 FILLER_34_382 ();
 sg13g2_fill_2 FILLER_34_395 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_fill_1 FILLER_35_91 ();
 sg13g2_fill_1 FILLER_35_149 ();
 sg13g2_fill_1 FILLER_35_387 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_4 FILLER_36_91 ();
 sg13g2_fill_1 FILLER_36_95 ();
 sg13g2_fill_1 FILLER_36_186 ();
 sg13g2_fill_1 FILLER_36_229 ();
 sg13g2_fill_2 FILLER_36_286 ();
 sg13g2_fill_2 FILLER_36_324 ();
 sg13g2_fill_2 FILLER_36_346 ();
 sg13g2_fill_2 FILLER_36_363 ();
 sg13g2_fill_2 FILLER_36_416 ();
 sg13g2_fill_1 FILLER_36_418 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_fill_1 FILLER_37_98 ();
 sg13g2_fill_1 FILLER_37_187 ();
 sg13g2_fill_1 FILLER_37_213 ();
 sg13g2_fill_2 FILLER_37_273 ();
 sg13g2_fill_2 FILLER_37_347 ();
 sg13g2_fill_1 FILLER_37_349 ();
 sg13g2_fill_2 FILLER_37_417 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_4 FILLER_38_98 ();
 sg13g2_fill_2 FILLER_38_102 ();
 sg13g2_fill_2 FILLER_38_145 ();
 sg13g2_fill_1 FILLER_38_255 ();
 sg13g2_fill_2 FILLER_38_337 ();
 sg13g2_fill_1 FILLER_38_339 ();
 sg13g2_fill_2 FILLER_38_369 ();
 sg13g2_fill_2 FILLER_38_417 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_fill_2 FILLER_39_91 ();
 sg13g2_fill_2 FILLER_39_133 ();
 sg13g2_fill_1 FILLER_39_144 ();
 sg13g2_fill_2 FILLER_39_190 ();
 sg13g2_fill_2 FILLER_39_264 ();
 sg13g2_fill_2 FILLER_39_304 ();
 sg13g2_fill_1 FILLER_39_306 ();
 sg13g2_fill_1 FILLER_39_393 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_fill_1 FILLER_40_178 ();
 sg13g2_fill_2 FILLER_40_297 ();
 sg13g2_fill_2 FILLER_40_352 ();
 sg13g2_fill_2 FILLER_40_359 ();
 sg13g2_fill_2 FILLER_40_371 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_fill_2 FILLER_41_105 ();
 sg13g2_fill_1 FILLER_41_107 ();
 sg13g2_fill_1 FILLER_41_350 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_fill_2 FILLER_42_105 ();
 sg13g2_fill_2 FILLER_42_148 ();
 sg13g2_fill_2 FILLER_42_357 ();
 sg13g2_fill_2 FILLER_42_364 ();
 sg13g2_fill_2 FILLER_42_417 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_fill_2 FILLER_43_105 ();
 sg13g2_fill_1 FILLER_43_116 ();
 sg13g2_fill_2 FILLER_43_253 ();
 sg13g2_fill_2 FILLER_43_356 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_fill_2 FILLER_44_98 ();
 sg13g2_fill_2 FILLER_44_125 ();
 sg13g2_fill_2 FILLER_44_243 ();
 sg13g2_fill_1 FILLER_44_263 ();
 sg13g2_fill_1 FILLER_44_274 ();
 sg13g2_fill_2 FILLER_44_293 ();
 sg13g2_fill_1 FILLER_44_367 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_4 FILLER_45_91 ();
 sg13g2_fill_2 FILLER_45_95 ();
 sg13g2_fill_1 FILLER_45_143 ();
 sg13g2_fill_2 FILLER_45_195 ();
 sg13g2_fill_1 FILLER_45_264 ();
 sg13g2_fill_2 FILLER_45_275 ();
 sg13g2_fill_1 FILLER_45_307 ();
 sg13g2_fill_1 FILLER_45_418 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_4 FILLER_46_98 ();
 sg13g2_fill_1 FILLER_46_148 ();
 sg13g2_fill_2 FILLER_46_215 ();
 sg13g2_fill_1 FILLER_46_217 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_fill_1 FILLER_47_105 ();
 sg13g2_fill_1 FILLER_47_171 ();
 sg13g2_fill_1 FILLER_47_303 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_4 FILLER_48_98 ();
 sg13g2_fill_1 FILLER_48_102 ();
 sg13g2_fill_1 FILLER_48_139 ();
 sg13g2_fill_1 FILLER_48_173 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_fill_2 FILLER_49_91 ();
 sg13g2_fill_1 FILLER_49_120 ();
 sg13g2_fill_2 FILLER_49_186 ();
 sg13g2_fill_1 FILLER_49_198 ();
 sg13g2_fill_1 FILLER_49_236 ();
 sg13g2_fill_1 FILLER_49_243 ();
 sg13g2_fill_2 FILLER_49_263 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_fill_2 FILLER_50_84 ();
 sg13g2_fill_2 FILLER_50_198 ();
 sg13g2_fill_1 FILLER_50_367 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_fill_2 FILLER_51_91 ();
 sg13g2_fill_1 FILLER_51_93 ();
 sg13g2_fill_1 FILLER_51_177 ();
 sg13g2_fill_2 FILLER_51_292 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_fill_1 FILLER_52_179 ();
 sg13g2_fill_1 FILLER_52_335 ();
 sg13g2_fill_1 FILLER_52_418 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_fill_2 FILLER_53_114 ();
 sg13g2_fill_2 FILLER_53_170 ();
 sg13g2_fill_1 FILLER_53_205 ();
 sg13g2_fill_1 FILLER_53_228 ();
 sg13g2_fill_2 FILLER_53_262 ();
 sg13g2_fill_1 FILLER_53_316 ();
 sg13g2_fill_2 FILLER_53_377 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_fill_2 FILLER_54_166 ();
 sg13g2_fill_1 FILLER_54_226 ();
 sg13g2_fill_1 FILLER_54_281 ();
 sg13g2_fill_1 FILLER_54_418 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_fill_1 FILLER_55_98 ();
 sg13g2_fill_1 FILLER_55_130 ();
 sg13g2_fill_1 FILLER_55_152 ();
 sg13g2_fill_1 FILLER_55_289 ();
 sg13g2_fill_1 FILLER_55_360 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_fill_2 FILLER_56_327 ();
 sg13g2_fill_1 FILLER_56_400 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_fill_1 FILLER_57_139 ();
 sg13g2_fill_1 FILLER_57_161 ();
 sg13g2_fill_2 FILLER_57_171 ();
 sg13g2_fill_1 FILLER_57_209 ();
 sg13g2_fill_2 FILLER_57_292 ();
 sg13g2_fill_1 FILLER_57_371 ();
 sg13g2_fill_1 FILLER_57_418 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_fill_2 FILLER_58_91 ();
 sg13g2_fill_1 FILLER_58_93 ();
 sg13g2_fill_2 FILLER_58_161 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_4 FILLER_59_84 ();
 sg13g2_fill_2 FILLER_59_88 ();
 sg13g2_fill_2 FILLER_59_171 ();
 sg13g2_fill_2 FILLER_59_223 ();
 sg13g2_fill_1 FILLER_59_241 ();
 sg13g2_fill_2 FILLER_59_307 ();
 sg13g2_fill_2 FILLER_59_318 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_4 FILLER_60_77 ();
 sg13g2_fill_1 FILLER_60_124 ();
 sg13g2_fill_1 FILLER_60_245 ();
 sg13g2_fill_1 FILLER_60_346 ();
 sg13g2_fill_1 FILLER_60_385 ();
 sg13g2_fill_2 FILLER_60_417 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_fill_2 FILLER_61_77 ();
 sg13g2_fill_1 FILLER_61_143 ();
 sg13g2_fill_2 FILLER_61_267 ();
 sg13g2_fill_1 FILLER_61_371 ();
 sg13g2_fill_2 FILLER_61_388 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_4 FILLER_62_70 ();
 sg13g2_fill_1 FILLER_62_74 ();
 sg13g2_fill_1 FILLER_62_327 ();
 sg13g2_fill_1 FILLER_62_391 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_fill_2 FILLER_63_77 ();
 sg13g2_fill_1 FILLER_63_79 ();
 sg13g2_fill_2 FILLER_63_288 ();
 sg13g2_fill_1 FILLER_63_383 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_4 FILLER_64_77 ();
 sg13g2_fill_1 FILLER_64_159 ();
 sg13g2_fill_1 FILLER_64_236 ();
 sg13g2_fill_1 FILLER_64_255 ();
 sg13g2_fill_1 FILLER_64_409 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_fill_2 FILLER_65_70 ();
 sg13g2_fill_2 FILLER_65_180 ();
 sg13g2_fill_2 FILLER_65_258 ();
 sg13g2_fill_1 FILLER_65_367 ();
 sg13g2_fill_2 FILLER_65_400 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_4 FILLER_66_70 ();
 sg13g2_fill_2 FILLER_66_74 ();
 sg13g2_fill_1 FILLER_66_229 ();
 sg13g2_fill_1 FILLER_66_257 ();
 sg13g2_fill_1 FILLER_66_274 ();
 sg13g2_fill_2 FILLER_66_389 ();
 sg13g2_fill_2 FILLER_66_408 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_fill_2 FILLER_67_70 ();
 sg13g2_fill_1 FILLER_67_175 ();
 sg13g2_fill_1 FILLER_67_222 ();
 sg13g2_fill_2 FILLER_67_383 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_fill_1 FILLER_68_70 ();
 sg13g2_fill_1 FILLER_68_239 ();
 sg13g2_fill_2 FILLER_68_390 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_4 FILLER_69_63 ();
 sg13g2_fill_2 FILLER_69_67 ();
 sg13g2_fill_1 FILLER_69_284 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_4 FILLER_70_63 ();
 sg13g2_fill_2 FILLER_70_67 ();
 sg13g2_fill_2 FILLER_70_197 ();
 sg13g2_fill_1 FILLER_70_228 ();
 sg13g2_fill_1 FILLER_70_389 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_fill_1 FILLER_71_130 ();
 sg13g2_fill_1 FILLER_71_260 ();
 sg13g2_fill_1 FILLER_71_383 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_fill_2 FILLER_72_70 ();
 sg13g2_fill_1 FILLER_72_72 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_fill_1 FILLER_73_70 ();
 sg13g2_fill_1 FILLER_73_164 ();
 sg13g2_fill_1 FILLER_73_228 ();
 sg13g2_fill_2 FILLER_73_259 ();
 sg13g2_fill_1 FILLER_73_409 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_4 FILLER_74_70 ();
 sg13g2_fill_1 FILLER_74_74 ();
 sg13g2_fill_1 FILLER_74_156 ();
 sg13g2_fill_2 FILLER_74_166 ();
 sg13g2_fill_1 FILLER_74_195 ();
 sg13g2_fill_2 FILLER_74_260 ();
 sg13g2_fill_2 FILLER_74_336 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_4 FILLER_75_70 ();
 sg13g2_fill_1 FILLER_75_74 ();
 sg13g2_fill_1 FILLER_75_232 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_fill_2 FILLER_76_63 ();
 sg13g2_fill_1 FILLER_76_65 ();
 sg13g2_fill_2 FILLER_76_210 ();
 sg13g2_fill_1 FILLER_76_418 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_fill_2 FILLER_77_63 ();
 sg13g2_fill_1 FILLER_77_65 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_4 FILLER_78_49 ();
 sg13g2_fill_2 FILLER_78_53 ();
 sg13g2_fill_1 FILLER_78_240 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_4 FILLER_79_49 ();
 sg13g2_fill_1 FILLER_79_53 ();
 sg13g2_fill_2 FILLER_79_155 ();
 sg13g2_fill_2 FILLER_79_417 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_4 FILLER_80_35 ();
 sg13g2_fill_2 FILLER_80_156 ();
 sg13g2_fill_2 FILLER_80_238 ();
 assign uio_oe[0] = net;
 assign uio_oe[1] = net222;
 assign uio_oe[2] = net223;
 assign uio_oe[3] = net224;
 assign uio_oe[4] = net225;
 assign uio_oe[5] = net226;
 assign uio_oe[6] = net227;
 assign uio_oe[7] = net228;
 assign uio_out[0] = net229;
 assign uio_out[1] = net230;
 assign uio_out[2] = net231;
 assign uio_out[3] = net232;
 assign uio_out[4] = net233;
 assign uio_out[5] = net234;
 assign uio_out[6] = net235;
 assign uio_out[7] = net236;
 assign uo_out[1] = net237;
 assign uo_out[2] = net238;
 assign uo_out[3] = net239;
 assign uo_out[4] = net240;
 assign uo_out[5] = net241;
 assign uo_out[6] = net242;
 assign uo_out[7] = net243;
endmodule
