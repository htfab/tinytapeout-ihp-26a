module tt_um_aksp_mbist_mbisr (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire clknet_0_clk;
 wire done;
 wire fail;
 wire \u_top.bist_fail_addr[0] ;
 wire \u_top.bist_fail_addr[1] ;
 wire \u_top.bist_fail_addr[2] ;
 wire \u_top.bist_fail_addr[3] ;
 wire \u_top.bist_fail_addr[4] ;
 wire \u_top.bist_fail_valid ;
 wire \u_top.bist_mem_addr[0] ;
 wire \u_top.bist_mem_addr[1] ;
 wire \u_top.bist_mem_addr[2] ;
 wire \u_top.bist_mem_addr[3] ;
 wire \u_top.bist_mem_addr[4] ;
 wire \u_top.bist_mem_en ;
 wire \u_top.bist_mem_rdata[0] ;
 wire \u_top.bist_mem_wdata[0] ;
 wire \u_top.bist_mem_we ;
 wire \u_top.u_mbisr.inserted ;
 wire \u_top.u_mbist.addr[0] ;
 wire \u_top.u_mbist.addr[1] ;
 wire \u_top.u_mbist.addr[2] ;
 wire \u_top.u_mbist.addr[3] ;
 wire \u_top.u_mbist.addr[4] ;
 wire \u_top.u_mbist.read_addr[0] ;
 wire \u_top.u_mbist.read_addr[1] ;
 wire \u_top.u_mbist.read_addr[2] ;
 wire \u_top.u_mbist.read_addr[3] ;
 wire \u_top.u_mbist.read_addr[4] ;
 wire \u_top.u_mbist.read_phase ;
 wire \u_top.u_mbist.state[1] ;
 wire \u_top.u_mbist.state[2] ;
 wire \u_top.u_mbist.state[3] ;
 wire \u_top.u_mbist.state[4] ;
 wire \u_top.u_mbist.state[5] ;
 wire \u_top.u_mbist.state[6] ;
 wire \u_top.u_mbist.state[7] ;
 wire \u_top.u_mbist.state[8] ;
 wire \u_top.u_memory.mem_array[0][0] ;
 wire \u_top.u_memory.mem_array[10][0] ;
 wire \u_top.u_memory.mem_array[11][0] ;
 wire \u_top.u_memory.mem_array[12][0] ;
 wire \u_top.u_memory.mem_array[13][0] ;
 wire \u_top.u_memory.mem_array[14][0] ;
 wire \u_top.u_memory.mem_array[15][0] ;
 wire \u_top.u_memory.mem_array[16][0] ;
 wire \u_top.u_memory.mem_array[17][0] ;
 wire \u_top.u_memory.mem_array[18][0] ;
 wire \u_top.u_memory.mem_array[19][0] ;
 wire \u_top.u_memory.mem_array[1][0] ;
 wire \u_top.u_memory.mem_array[20][0] ;
 wire \u_top.u_memory.mem_array[21][0] ;
 wire \u_top.u_memory.mem_array[22][0] ;
 wire \u_top.u_memory.mem_array[23][0] ;
 wire \u_top.u_memory.mem_array[24][0] ;
 wire \u_top.u_memory.mem_array[25][0] ;
 wire \u_top.u_memory.mem_array[26][0] ;
 wire \u_top.u_memory.mem_array[27][0] ;
 wire \u_top.u_memory.mem_array[28][0] ;
 wire \u_top.u_memory.mem_array[29][0] ;
 wire \u_top.u_memory.mem_array[2][0] ;
 wire \u_top.u_memory.mem_array[30][0] ;
 wire \u_top.u_memory.mem_array[31][0] ;
 wire \u_top.u_memory.mem_array[3][0] ;
 wire \u_top.u_memory.mem_array[4][0] ;
 wire \u_top.u_memory.mem_array[5][0] ;
 wire \u_top.u_memory.mem_array[6][0] ;
 wire \u_top.u_memory.mem_array[7][0] ;
 wire \u_top.u_memory.mem_array[8][0] ;
 wire \u_top.u_memory.mem_array[9][0] ;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net1;
 wire net2;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire [0:0] _406_;
 wire [0:0] \u_top.u_mbisr.repair_valid[0] ;
 wire [0:0] \u_top.u_mbisr.repair_valid[1] ;

 sg13g2_inv_1 _407_ (.Y(_082_),
    .A(net64));
 sg13g2_inv_1 _408_ (.Y(_083_),
    .A(_363_));
 sg13g2_inv_1 _409_ (.Y(_084_),
    .A(net192));
 sg13g2_inv_2 _410_ (.Y(_085_),
    .A(net213));
 sg13g2_inv_1 _411_ (.Y(_086_),
    .A(net79));
 sg13g2_inv_2 _412_ (.Y(_087_),
    .A(net78));
 sg13g2_inv_1 _413_ (.Y(_088_),
    .A(\u_top.bist_mem_addr[3] ));
 sg13g2_inv_1 _414_ (.Y(_089_),
    .A(net232));
 sg13g2_inv_1 _415_ (.Y(_090_),
    .A(net86));
 sg13g2_inv_2 _416_ (.Y(_091_),
    .A(net217));
 sg13g2_inv_1 _417_ (.Y(_092_),
    .A(net209));
 sg13g2_inv_1 _418_ (.Y(_093_),
    .A(\u_top.bist_fail_valid ));
 sg13g2_inv_1 _419_ (.Y(_094_),
    .A(net202));
 sg13g2_inv_1 _420_ (.Y(_095_),
    .A(net81));
 sg13g2_inv_1 _421_ (.Y(_096_),
    .A(net105));
 sg13g2_inv_1 _422_ (.Y(_097_),
    .A(net148));
 sg13g2_inv_1 _423_ (.Y(_098_),
    .A(net158));
 sg13g2_nand2b_1 _424_ (.Y(_099_),
    .B(net227),
    .A_N(net99));
 sg13g2_nand2b_1 _425_ (.Y(_010_),
    .B(_099_),
    .A_N(net1));
 sg13g2_nor2b_1 _426_ (.A(net227),
    .B_N(net1),
    .Y(_100_));
 sg13g2_and3_1 _427_ (.X(_101_),
    .A(net202),
    .B(net231),
    .C(net225));
 sg13g2_and3_1 _428_ (.X(_102_),
    .A(net81),
    .B(net238),
    .C(_101_));
 sg13g2_nand3_1 _429_ (.B(net228),
    .C(_101_),
    .A(net81),
    .Y(_103_));
 sg13g2_a21o_1 _430_ (.A2(_103_),
    .A1(net165),
    .B1(_100_),
    .X(_004_));
 sg13g2_nor4_1 _431_ (.A(net150),
    .B(net81),
    .C(net169),
    .D(\u_top.u_mbist.addr[4] ),
    .Y(_104_));
 sg13g2_nand3_1 _432_ (.B(_094_),
    .C(_104_),
    .A(net80),
    .Y(_105_));
 sg13g2_a21o_1 _433_ (.A2(_105_),
    .A1(net217),
    .B1(net84),
    .X(_005_));
 sg13g2_and2_1 _434_ (.A(net80),
    .B(_102_),
    .X(_106_));
 sg13g2_nand2_1 _435_ (.Y(_107_),
    .A(net80),
    .B(_102_));
 sg13g2_a21o_1 _436_ (.A2(_107_),
    .A1(\u_top.u_mbist.state[7] ),
    .B1(net156),
    .X(_006_));
 sg13g2_a21o_1 _437_ (.A2(_107_),
    .A1(net82),
    .B1(net188),
    .X(_007_));
 sg13g2_a22oi_1 _438_ (.Y(_108_),
    .B1(_106_),
    .B2(net82),
    .A2(net99),
    .A1(net1));
 sg13g2_inv_1 _439_ (.Y(_003_),
    .A(_108_));
 sg13g2_nor2_1 _440_ (.A(_091_),
    .B(_105_),
    .Y(_002_));
 sg13g2_a21oi_1 _441_ (.A1(net82),
    .A2(_107_),
    .Y(_109_),
    .B1(_100_));
 sg13g2_o21ai_1 _442_ (.B1(_109_),
    .Y(_406_[0]),
    .A1(net82),
    .A2(_099_));
 sg13g2_nor2_2 _443_ (.A(net204),
    .B(net82),
    .Y(_110_));
 sg13g2_nor2_1 _444_ (.A(net223),
    .B(net217),
    .Y(_111_));
 sg13g2_nand2_2 _445_ (.Y(_112_),
    .A(_091_),
    .B(_110_));
 sg13g2_nand2_1 _446_ (.Y(_113_),
    .A(net80),
    .B(_112_));
 sg13g2_xnor2_1 _447_ (.Y(_114_),
    .A(net192),
    .B(_110_));
 sg13g2_nor2_1 _448_ (.A(_113_),
    .B(_114_),
    .Y(_008_));
 sg13g2_and2_1 _449_ (.A(net165),
    .B(_102_),
    .X(_001_));
 sg13g2_and2_1 _450_ (.A(net204),
    .B(_106_),
    .X(_000_));
 sg13g2_nor2_1 _451_ (.A(_364_),
    .B(net79),
    .Y(_115_));
 sg13g2_nand2_1 _452_ (.Y(_116_),
    .A(_366_),
    .B(\u_top.bist_mem_addr[3] ));
 sg13g2_nor2_1 _453_ (.A(_366_),
    .B(\u_top.bist_mem_addr[3] ),
    .Y(_117_));
 sg13g2_o21ai_1 _454_ (.B1(\u_top.u_mbisr.repair_valid[0] [0]),
    .Y(_118_),
    .A1(_365_),
    .A2(net78));
 sg13g2_xnor2_1 _455_ (.Y(_119_),
    .A(_367_),
    .B(\u_top.bist_mem_addr[4] ));
 sg13g2_nor3_1 _456_ (.A(_115_),
    .B(_117_),
    .C(_119_),
    .Y(_120_));
 sg13g2_a22oi_1 _457_ (.Y(_121_),
    .B1(net79),
    .B2(_364_),
    .A2(\u_top.bist_mem_addr[0] ),
    .A1(_363_));
 sg13g2_a221oi_1 _458_ (.B2(_365_),
    .C1(_118_),
    .B1(net78),
    .A1(_083_),
    .Y(_122_),
    .A2(_085_));
 sg13g2_and4_1 _459_ (.A(_116_),
    .B(_120_),
    .C(_121_),
    .D(_122_),
    .X(_123_));
 sg13g2_nand4_1 _460_ (.B(_120_),
    .C(_121_),
    .A(_116_),
    .Y(_124_),
    .D(_122_));
 sg13g2_xor2_1 _461_ (.B(\u_top.bist_mem_addr[4] ),
    .A(_362_),
    .X(_125_));
 sg13g2_xor2_1 _462_ (.B(\u_top.bist_mem_addr[0] ),
    .A(_358_),
    .X(_126_));
 sg13g2_xnor2_1 _463_ (.Y(_127_),
    .A(_361_),
    .B(\u_top.bist_mem_addr[3] ));
 sg13g2_o21ai_1 _464_ (.B1(_126_),
    .Y(_128_),
    .A1(_360_),
    .A2(net78));
 sg13g2_o21ai_1 _465_ (.B1(\u_top.u_mbisr.repair_valid[1] [0]),
    .Y(_129_),
    .A1(_359_),
    .A2(net79));
 sg13g2_a22oi_1 _466_ (.Y(_130_),
    .B1(\u_top.bist_mem_addr[2] ),
    .B2(_360_),
    .A2(net79),
    .A1(_359_));
 sg13g2_nand2_1 _467_ (.Y(_131_),
    .A(_125_),
    .B(_130_));
 sg13g2_nor4_1 _468_ (.A(_127_),
    .B(_128_),
    .C(_129_),
    .D(_131_),
    .Y(_132_));
 sg13g2_nor3_2 _469_ (.A(\u_top.bist_mem_addr[4] ),
    .B(_123_),
    .C(net68),
    .Y(_133_));
 sg13g2_and3_1 _470_ (.X(_134_),
    .A(_087_),
    .B(\u_top.bist_mem_addr[3] ),
    .C(_133_));
 sg13g2_nand3_1 _471_ (.B(\u_top.bist_mem_addr[3] ),
    .C(_133_),
    .A(_087_),
    .Y(_135_));
 sg13g2_and3_2 _472_ (.X(_136_),
    .A(\u_top.bist_mem_we ),
    .B(\u_top.bist_mem_en ),
    .C(net86));
 sg13g2_or2_1 _473_ (.X(_137_),
    .B(_132_),
    .A(net79));
 sg13g2_or3_1 _474_ (.A(net79),
    .B(_123_),
    .C(net68),
    .X(_138_));
 sg13g2_nor4_2 _475_ (.A(\u_top.bist_mem_addr[0] ),
    .B(net79),
    .C(_123_),
    .Y(_139_),
    .D(net68));
 sg13g2_nand2_2 _476_ (.Y(_140_),
    .A(_136_),
    .B(net67));
 sg13g2_or2_1 _477_ (.X(_141_),
    .B(_140_),
    .A(_135_));
 sg13g2_nand3_1 _478_ (.B(net114),
    .C(_141_),
    .A(net86),
    .Y(_142_));
 sg13g2_o21ai_1 _479_ (.B1(_142_),
    .Y(_011_),
    .A1(net73),
    .A2(_141_));
 sg13g2_a21oi_1 _480_ (.A1(\u_top.bist_mem_addr[0] ),
    .A2(_124_),
    .Y(_143_),
    .B1(net68));
 sg13g2_a21o_2 _481_ (.A2(_124_),
    .A1(\u_top.bist_mem_addr[0] ),
    .B1(net68),
    .X(_144_));
 sg13g2_and2_1 _482_ (.A(_137_),
    .B(_144_),
    .X(_145_));
 sg13g2_and2_1 _483_ (.A(_136_),
    .B(_145_),
    .X(_146_));
 sg13g2_nand2_2 _484_ (.Y(_147_),
    .A(_136_),
    .B(_145_));
 sg13g2_nand2_1 _485_ (.Y(_148_),
    .A(_134_),
    .B(_146_));
 sg13g2_nand3_1 _486_ (.B(net138),
    .C(_148_),
    .A(net97),
    .Y(_149_));
 sg13g2_o21ai_1 _487_ (.B1(_149_),
    .Y(_012_),
    .A1(net73),
    .A2(_148_));
 sg13g2_nand3_1 _488_ (.B(\u_top.bist_mem_addr[3] ),
    .C(_133_),
    .A(net78),
    .Y(_150_));
 sg13g2_or2_1 _489_ (.X(_151_),
    .B(_150_),
    .A(_140_));
 sg13g2_nand3_1 _490_ (.B(net103),
    .C(_151_),
    .A(net85),
    .Y(_152_));
 sg13g2_o21ai_1 _491_ (.B1(_152_),
    .Y(_013_),
    .A1(net72),
    .A2(_151_));
 sg13g2_nor4_2 _492_ (.A(_085_),
    .B(\u_top.bist_mem_addr[1] ),
    .C(_123_),
    .Y(_153_),
    .D(net68));
 sg13g2_nand2_2 _493_ (.Y(_154_),
    .A(_136_),
    .B(net66));
 sg13g2_or2_1 _494_ (.X(_155_),
    .B(_154_),
    .A(_150_));
 sg13g2_nand3_1 _495_ (.B(net111),
    .C(_155_),
    .A(net85),
    .Y(_156_));
 sg13g2_o21ai_1 _496_ (.B1(_156_),
    .Y(_014_),
    .A1(net72),
    .A2(_155_));
 sg13g2_nor3_2 _497_ (.A(\u_top.bist_mem_addr[3] ),
    .B(_123_),
    .C(net68),
    .Y(_157_));
 sg13g2_nor2_1 _498_ (.A(_133_),
    .B(_157_),
    .Y(_158_));
 sg13g2_nor3_1 _499_ (.A(net78),
    .B(_123_),
    .C(net68),
    .Y(_159_));
 sg13g2_nand2_2 _500_ (.Y(_160_),
    .A(_158_),
    .B(_159_));
 sg13g2_or2_1 _501_ (.X(_161_),
    .B(_160_),
    .A(_147_));
 sg13g2_nand3_1 _502_ (.B(net125),
    .C(_161_),
    .A(net91),
    .Y(_162_));
 sg13g2_o21ai_1 _503_ (.B1(_162_),
    .Y(_015_),
    .A1(net74),
    .A2(_161_));
 sg13g2_and3_2 _504_ (.X(_163_),
    .A(_087_),
    .B(_089_),
    .C(_157_));
 sg13g2_nand2b_1 _505_ (.Y(_164_),
    .B(_163_),
    .A_N(_140_));
 sg13g2_nand3_1 _506_ (.B(net141),
    .C(_164_),
    .A(net92),
    .Y(_165_));
 sg13g2_o21ai_1 _507_ (.B1(_165_),
    .Y(_016_),
    .A1(net75),
    .A2(_164_));
 sg13g2_nand3_1 _508_ (.B(_137_),
    .C(_144_),
    .A(\u_top.u_memory.mem_array[3][0] ),
    .Y(_166_));
 sg13g2_and2_1 _509_ (.A(_138_),
    .B(_143_),
    .X(_167_));
 sg13g2_nand3_1 _510_ (.B(_138_),
    .C(_143_),
    .A(\u_top.u_memory.mem_array[2][0] ),
    .Y(_168_));
 sg13g2_a22oi_1 _511_ (.Y(_169_),
    .B1(net66),
    .B2(\u_top.u_memory.mem_array[1][0] ),
    .A2(net67),
    .A1(\u_top.u_memory.mem_array[0][0] ));
 sg13g2_nand3_1 _512_ (.B(_168_),
    .C(_169_),
    .A(_166_),
    .Y(_170_));
 sg13g2_nand3_1 _513_ (.B(_089_),
    .C(_157_),
    .A(net78),
    .Y(_171_));
 sg13g2_inv_1 _514_ (.Y(_172_),
    .A(_171_));
 sg13g2_nand3_1 _515_ (.B(_138_),
    .C(_143_),
    .A(\u_top.u_memory.mem_array[6][0] ),
    .Y(_173_));
 sg13g2_nand3_1 _516_ (.B(_137_),
    .C(_144_),
    .A(\u_top.u_memory.mem_array[7][0] ),
    .Y(_174_));
 sg13g2_a22oi_1 _517_ (.Y(_175_),
    .B1(net66),
    .B2(\u_top.u_memory.mem_array[5][0] ),
    .A2(net67),
    .A1(\u_top.u_memory.mem_array[4][0] ));
 sg13g2_nand3_1 _518_ (.B(_174_),
    .C(_175_),
    .A(_173_),
    .Y(_176_));
 sg13g2_nor3_2 _519_ (.A(_133_),
    .B(_157_),
    .C(_159_),
    .Y(_177_));
 sg13g2_nand3_1 _520_ (.B(_137_),
    .C(_144_),
    .A(\u_top.u_memory.mem_array[31][0] ),
    .Y(_178_));
 sg13g2_nand2_1 _521_ (.Y(_179_),
    .A(\u_top.u_memory.mem_array[29][0] ),
    .B(net66));
 sg13g2_nand2_1 _522_ (.Y(_180_),
    .A(\u_top.u_memory.mem_array[28][0] ),
    .B(net67));
 sg13g2_nand3_1 _523_ (.B(_138_),
    .C(_143_),
    .A(\u_top.u_memory.mem_array[30][0] ),
    .Y(_181_));
 sg13g2_nand4_1 _524_ (.B(_179_),
    .C(_180_),
    .A(_178_),
    .Y(_182_),
    .D(_181_));
 sg13g2_nand3_1 _525_ (.B(\u_top.bist_mem_addr[4] ),
    .C(_157_),
    .A(_087_),
    .Y(_183_));
 sg13g2_a22oi_1 _526_ (.Y(_184_),
    .B1(net66),
    .B2(net126),
    .A2(_145_),
    .A1(\u_top.u_memory.mem_array[19][0] ));
 sg13g2_a22oi_1 _527_ (.Y(_185_),
    .B1(_167_),
    .B2(net112),
    .A2(net67),
    .A1(net132));
 sg13g2_a21oi_1 _528_ (.A1(_184_),
    .A2(_185_),
    .Y(_186_),
    .B1(_183_));
 sg13g2_nand2b_1 _529_ (.Y(_187_),
    .B(net206),
    .A_N(\u_top.bist_mem_we ));
 sg13g2_a22oi_1 _530_ (.Y(_188_),
    .B1(net66),
    .B2(\u_top.u_memory.mem_array[25][0] ),
    .A2(net67),
    .A1(\u_top.u_memory.mem_array[24][0] ));
 sg13g2_a22oi_1 _531_ (.Y(_189_),
    .B1(_167_),
    .B2(\u_top.u_memory.mem_array[26][0] ),
    .A2(_145_),
    .A1(\u_top.u_memory.mem_array[27][0] ));
 sg13g2_a21o_1 _532_ (.A2(_189_),
    .A1(_188_),
    .B1(_160_),
    .X(_190_));
 sg13g2_a22oi_1 _533_ (.Y(_191_),
    .B1(net66),
    .B2(net111),
    .A2(_145_),
    .A1(net116));
 sg13g2_a22oi_1 _534_ (.Y(_192_),
    .B1(_167_),
    .B2(net101),
    .A2(net67),
    .A1(net103));
 sg13g2_a21oi_1 _535_ (.A1(_191_),
    .A2(_192_),
    .Y(_193_),
    .B1(_150_));
 sg13g2_nand3_1 _536_ (.B(\u_top.bist_mem_addr[4] ),
    .C(_157_),
    .A(net78),
    .Y(_194_));
 sg13g2_a22oi_1 _537_ (.Y(_195_),
    .B1(_145_),
    .B2(\u_top.u_memory.mem_array[23][0] ),
    .A2(_139_),
    .A1(\u_top.u_memory.mem_array[20][0] ));
 sg13g2_a22oi_1 _538_ (.Y(_196_),
    .B1(_167_),
    .B2(\u_top.u_memory.mem_array[22][0] ),
    .A2(_153_),
    .A1(\u_top.u_memory.mem_array[21][0] ));
 sg13g2_a21o_1 _539_ (.A2(_196_),
    .A1(_195_),
    .B1(_194_),
    .X(_197_));
 sg13g2_a22oi_1 _540_ (.Y(_198_),
    .B1(net66),
    .B2(net134),
    .A2(net67),
    .A1(net114));
 sg13g2_a22oi_1 _541_ (.Y(_199_),
    .B1(_167_),
    .B2(net109),
    .A2(_145_),
    .A1(net138));
 sg13g2_a21oi_1 _542_ (.A1(_198_),
    .A2(_199_),
    .Y(_200_),
    .B1(_135_));
 sg13g2_nor3_1 _543_ (.A(_186_),
    .B(_193_),
    .C(_200_),
    .Y(_201_));
 sg13g2_a21oi_1 _544_ (.A1(_172_),
    .A2(_176_),
    .Y(_202_),
    .B1(_187_));
 sg13g2_a22oi_1 _545_ (.Y(_203_),
    .B1(_177_),
    .B2(_182_),
    .A2(_170_),
    .A1(_163_));
 sg13g2_and4_1 _546_ (.A(_190_),
    .B(_197_),
    .C(_202_),
    .D(_203_),
    .X(_204_));
 sg13g2_a221oi_1 _547_ (.B2(_204_),
    .C1(_090_),
    .B1(_201_),
    .A1(_084_),
    .Y(_017_),
    .A2(net207));
 sg13g2_and2_1 _548_ (.A(_136_),
    .B(_167_),
    .X(_205_));
 sg13g2_nand2_1 _549_ (.Y(_206_),
    .A(_163_),
    .B(_205_));
 sg13g2_nand3_1 _550_ (.B(net173),
    .C(_206_),
    .A(net92),
    .Y(_207_));
 sg13g2_o21ai_1 _551_ (.B1(_207_),
    .Y(_018_),
    .A1(net74),
    .A2(_206_));
 sg13g2_nand2_1 _552_ (.Y(_208_),
    .A(_177_),
    .B(_205_));
 sg13g2_nand3_1 _553_ (.B(net131),
    .C(_208_),
    .A(net92),
    .Y(_209_));
 sg13g2_o21ai_1 _554_ (.B1(_209_),
    .Y(_019_),
    .A1(net76),
    .A2(_208_));
 sg13g2_nand2_1 _555_ (.Y(_210_),
    .A(\u_top.u_mbist.addr[0] ),
    .B(_112_));
 sg13g2_nor3_1 _556_ (.A(\u_top.u_mbist.state[4] ),
    .B(\u_top.u_mbist.state[3] ),
    .C(_112_),
    .Y(_211_));
 sg13g2_or3_1 _557_ (.A(net188),
    .B(net156),
    .C(_112_),
    .X(_212_));
 sg13g2_and2_1 _558_ (.A(_113_),
    .B(_212_),
    .X(_213_));
 sg13g2_nor2_1 _559_ (.A(net83),
    .B(_212_),
    .Y(_214_));
 sg13g2_o21ai_1 _560_ (.B1(_113_),
    .Y(_215_),
    .A1(net84),
    .A2(_212_));
 sg13g2_a22oi_1 _561_ (.Y(_020_),
    .B1(_215_),
    .B2(_096_),
    .A2(_213_),
    .A1(_210_));
 sg13g2_nand2_1 _562_ (.Y(_216_),
    .A(net150),
    .B(_112_));
 sg13g2_a22oi_1 _563_ (.Y(_021_),
    .B1(net151),
    .B2(_213_),
    .A2(_215_),
    .A1(_097_));
 sg13g2_nand2_1 _564_ (.Y(_217_),
    .A(net169),
    .B(_112_));
 sg13g2_a22oi_1 _565_ (.Y(_022_),
    .B1(net170),
    .B2(_213_),
    .A2(_215_),
    .A1(_098_));
 sg13g2_a21oi_1 _566_ (.A1(net81),
    .A2(_112_),
    .Y(_218_),
    .B1(_211_));
 sg13g2_nand2_1 _567_ (.Y(_219_),
    .A(net62),
    .B(_215_));
 sg13g2_o21ai_1 _568_ (.B1(_219_),
    .Y(_023_),
    .A1(_215_),
    .A2(_218_));
 sg13g2_a21oi_1 _569_ (.A1(\u_top.u_mbist.addr[4] ),
    .A2(_112_),
    .Y(_220_),
    .B1(_211_));
 sg13g2_nand2_1 _570_ (.Y(_221_),
    .A(net129),
    .B(_215_));
 sg13g2_o21ai_1 _571_ (.B1(_221_),
    .Y(_024_),
    .A1(_215_),
    .A2(_220_));
 sg13g2_or2_1 _572_ (.X(_222_),
    .B(_171_),
    .A(_140_));
 sg13g2_nand3_1 _573_ (.B(net107),
    .C(_222_),
    .A(net91),
    .Y(_223_));
 sg13g2_o21ai_1 _574_ (.B1(_223_),
    .Y(_025_),
    .A1(net76),
    .A2(_222_));
 sg13g2_or2_1 _575_ (.X(_224_),
    .B(_171_),
    .A(_154_));
 sg13g2_nand3_1 _576_ (.B(net123),
    .C(_224_),
    .A(net91),
    .Y(_225_));
 sg13g2_o21ai_1 _577_ (.B1(_225_),
    .Y(_026_),
    .A1(net77),
    .A2(_224_));
 sg13g2_nand2_1 _578_ (.Y(_226_),
    .A(_172_),
    .B(_205_));
 sg13g2_nand3_1 _579_ (.B(net144),
    .C(_226_),
    .A(net93),
    .Y(_227_));
 sg13g2_o21ai_1 _580_ (.B1(_227_),
    .Y(_027_),
    .A1(net76),
    .A2(_226_));
 sg13g2_nand2b_1 _581_ (.Y(_228_),
    .B(_205_),
    .A_N(_183_));
 sg13g2_nand3_1 _582_ (.B(net112),
    .C(_228_),
    .A(net85),
    .Y(_229_));
 sg13g2_o21ai_1 _583_ (.B1(_229_),
    .Y(_028_),
    .A1(net72),
    .A2(_228_));
 sg13g2_nand2_1 _584_ (.Y(_230_),
    .A(_134_),
    .B(_205_));
 sg13g2_nand3_1 _585_ (.B(net109),
    .C(_230_),
    .A(net91),
    .Y(_231_));
 sg13g2_o21ai_1 _586_ (.B1(_231_),
    .Y(_029_),
    .A1(net73),
    .A2(_230_));
 sg13g2_nand2b_1 _587_ (.Y(_232_),
    .B(_177_),
    .A_N(_140_));
 sg13g2_nand3_1 _588_ (.B(net155),
    .C(_232_),
    .A(net93),
    .Y(_233_));
 sg13g2_o21ai_1 _589_ (.B1(_233_),
    .Y(_030_),
    .A1(net74),
    .A2(_232_));
 sg13g2_or2_1 _590_ (.X(_234_),
    .B(_183_),
    .A(_140_));
 sg13g2_nand3_1 _591_ (.B(net132),
    .C(_234_),
    .A(net85),
    .Y(_235_));
 sg13g2_o21ai_1 _592_ (.B1(_235_),
    .Y(_031_),
    .A1(net72),
    .A2(_234_));
 sg13g2_or2_1 _593_ (.X(_236_),
    .B(_154_),
    .A(_135_));
 sg13g2_nand3_1 _594_ (.B(net134),
    .C(_236_),
    .A(net86),
    .Y(_237_));
 sg13g2_o21ai_1 _595_ (.B1(_237_),
    .Y(_032_),
    .A1(net73),
    .A2(_236_));
 sg13g2_nand2b_1 _596_ (.Y(_238_),
    .B(_205_),
    .A_N(_150_));
 sg13g2_nand3_1 _597_ (.B(net101),
    .C(_238_),
    .A(net85),
    .Y(_239_));
 sg13g2_o21ai_1 _598_ (.B1(_239_),
    .Y(_033_),
    .A1(net72),
    .A2(_238_));
 sg13g2_or2_1 _599_ (.X(_240_),
    .B(_194_),
    .A(_147_));
 sg13g2_nand3_1 _600_ (.B(net119),
    .C(_240_),
    .A(net92),
    .Y(_241_));
 sg13g2_o21ai_1 _601_ (.B1(_241_),
    .Y(_034_),
    .A1(net74),
    .A2(_240_));
 sg13g2_or2_1 _602_ (.X(_242_),
    .B(_160_),
    .A(_140_));
 sg13g2_nand3_1 _603_ (.B(net121),
    .C(_242_),
    .A(net91),
    .Y(_243_));
 sg13g2_o21ai_1 _604_ (.B1(_243_),
    .Y(_035_),
    .A1(net74),
    .A2(_242_));
 sg13g2_nand2b_1 _605_ (.Y(_244_),
    .B(_177_),
    .A_N(_154_));
 sg13g2_nand3_1 _606_ (.B(net179),
    .C(_244_),
    .A(net93),
    .Y(_245_));
 sg13g2_o21ai_1 _607_ (.B1(_245_),
    .Y(_036_),
    .A1(net74),
    .A2(_244_));
 sg13g2_nor2_1 _608_ (.A(_147_),
    .B(_183_),
    .Y(_246_));
 sg13g2_nand2_1 _609_ (.Y(_247_),
    .A(net64),
    .B(_246_));
 sg13g2_nand2_1 _610_ (.Y(_248_),
    .A(net85),
    .B(\u_top.u_memory.mem_array[19][0] ));
 sg13g2_o21ai_1 _611_ (.B1(net65),
    .Y(_037_),
    .A1(_246_),
    .A2(_248_));
 sg13g2_or2_1 _612_ (.X(_249_),
    .B(_160_),
    .A(_154_));
 sg13g2_nand3_1 _613_ (.B(net140),
    .C(_249_),
    .A(net91),
    .Y(_250_));
 sg13g2_o21ai_1 _614_ (.B1(_250_),
    .Y(_038_),
    .A1(net74),
    .A2(_249_));
 sg13g2_nand2b_1 _615_ (.Y(_251_),
    .B(_205_),
    .A_N(_160_));
 sg13g2_nand3_1 _616_ (.B(net128),
    .C(_251_),
    .A(net91),
    .Y(_252_));
 sg13g2_o21ai_1 _617_ (.B1(_252_),
    .Y(_039_),
    .A1(net74),
    .A2(_251_));
 sg13g2_nor3_2 _618_ (.A(net234),
    .B(net209),
    .C(_093_),
    .Y(_253_));
 sg13g2_or2_1 _619_ (.X(_040_),
    .B(_253_),
    .A(net234));
 sg13g2_nor2_1 _620_ (.A(_367_),
    .B(net190),
    .Y(_254_));
 sg13g2_a221oi_1 _621_ (.B2(net163),
    .C1(_254_),
    .B1(net181),
    .A1(net184),
    .Y(_255_),
    .A2(net171));
 sg13g2_or2_1 _622_ (.X(_256_),
    .B(net171),
    .A(net184));
 sg13g2_o21ai_1 _623_ (.B1(_256_),
    .Y(_257_),
    .A1(net199),
    .A2(net153));
 sg13g2_a221oi_1 _624_ (.B2(net153),
    .C1(_257_),
    .B1(net199),
    .A1(_367_),
    .Y(_258_),
    .A2(net190));
 sg13g2_xnor2_1 _625_ (.Y(_259_),
    .A(_366_),
    .B(net174));
 sg13g2_o21ai_1 _626_ (.B1(\u_top.u_mbisr.repair_valid[0] [0]),
    .Y(_260_),
    .A1(net181),
    .A2(net163));
 sg13g2_nor2_1 _627_ (.A(_259_),
    .B(_260_),
    .Y(_261_));
 sg13g2_nand3_1 _628_ (.B(_258_),
    .C(_261_),
    .A(_255_),
    .Y(_262_));
 sg13g2_nand2_1 _629_ (.Y(_263_),
    .A(\u_top.bist_fail_addr[4] ),
    .B(_362_));
 sg13g2_xnor2_1 _630_ (.Y(_264_),
    .A(\u_top.bist_fail_addr[1] ),
    .B(_359_));
 sg13g2_xnor2_1 _631_ (.Y(_265_),
    .A(\u_top.bist_fail_addr[3] ),
    .B(_361_));
 sg13g2_a22oi_1 _632_ (.Y(_266_),
    .B1(_358_),
    .B2(\u_top.bist_fail_addr[0] ),
    .A2(_360_),
    .A1(\u_top.bist_fail_addr[2] ));
 sg13g2_o21ai_1 _633_ (.B1(_266_),
    .Y(_267_),
    .A1(net171),
    .A2(_360_));
 sg13g2_o21ai_1 _634_ (.B1(\u_top.u_mbisr.repair_valid[1] [0]),
    .Y(_268_),
    .A1(\u_top.bist_fail_addr[4] ),
    .A2(_362_));
 sg13g2_o21ai_1 _635_ (.B1(_263_),
    .Y(_269_),
    .A1(\u_top.bist_fail_addr[0] ),
    .A2(_358_));
 sg13g2_nor4_1 _636_ (.A(_264_),
    .B(_265_),
    .C(_268_),
    .D(_269_),
    .Y(_270_));
 sg13g2_nor2b_1 _637_ (.A(_267_),
    .B_N(_270_),
    .Y(_271_));
 sg13g2_nor2_1 _638_ (.A(net221),
    .B(net209),
    .Y(_272_));
 sg13g2_o21ai_1 _639_ (.B1(\u_top.bist_fail_valid ),
    .Y(_273_),
    .A1(\u_top.u_mbisr.repair_valid[0] [0]),
    .A2(net209));
 sg13g2_nor3_1 _640_ (.A(_271_),
    .B(_272_),
    .C(_273_),
    .Y(_274_));
 sg13g2_a22oi_1 _641_ (.Y(_041_),
    .B1(_262_),
    .B2(_274_),
    .A2(_093_),
    .A1(_092_));
 sg13g2_and2_1 _642_ (.A(\u_top.bist_fail_valid ),
    .B(_272_),
    .X(_275_));
 sg13g2_nor2_1 _643_ (.A(net196),
    .B(net69),
    .Y(_276_));
 sg13g2_a21oi_1 _644_ (.A1(net153),
    .A2(net69),
    .Y(_042_),
    .B1(net197));
 sg13g2_nor2_1 _645_ (.A(_359_),
    .B(net69),
    .Y(_277_));
 sg13g2_a21oi_1 _646_ (.A1(net163),
    .A2(net69),
    .Y(_043_),
    .B1(_277_));
 sg13g2_nor2_1 _647_ (.A(_360_),
    .B(net69),
    .Y(_278_));
 sg13g2_a21oi_1 _648_ (.A1(net171),
    .A2(net69),
    .Y(_044_),
    .B1(_278_));
 sg13g2_nor2_1 _649_ (.A(net176),
    .B(net69),
    .Y(_279_));
 sg13g2_a21oi_1 _650_ (.A1(net174),
    .A2(net69),
    .Y(_045_),
    .B1(net177));
 sg13g2_nor2_1 _651_ (.A(net193),
    .B(_275_),
    .Y(_280_));
 sg13g2_a21oi_1 _652_ (.A1(net190),
    .A2(_275_),
    .Y(_046_),
    .B1(net194));
 sg13g2_nor2_1 _653_ (.A(net199),
    .B(net70),
    .Y(_281_));
 sg13g2_a21oi_1 _654_ (.A1(net153),
    .A2(net70),
    .Y(_047_),
    .B1(net200));
 sg13g2_nor2_1 _655_ (.A(net181),
    .B(net70),
    .Y(_282_));
 sg13g2_a21oi_1 _656_ (.A1(net163),
    .A2(net70),
    .Y(_048_),
    .B1(net182));
 sg13g2_nor2_1 _657_ (.A(net184),
    .B(net70),
    .Y(_283_));
 sg13g2_a21oi_1 _658_ (.A1(net171),
    .A2(net70),
    .Y(_049_),
    .B1(net185));
 sg13g2_nor2_1 _659_ (.A(_366_),
    .B(net70),
    .Y(_284_));
 sg13g2_a21oi_1 _660_ (.A1(net174),
    .A2(net70),
    .Y(_050_),
    .B1(_284_));
 sg13g2_nor2_1 _661_ (.A(_367_),
    .B(_253_),
    .Y(_285_));
 sg13g2_a21oi_1 _662_ (.A1(net190),
    .A2(_253_),
    .Y(_051_),
    .B1(_285_));
 sg13g2_nand2b_1 _663_ (.Y(_286_),
    .B(_205_),
    .A_N(_194_));
 sg13g2_nand3_1 _664_ (.B(net142),
    .C(_286_),
    .A(net92),
    .Y(_287_));
 sg13g2_o21ai_1 _665_ (.B1(_287_),
    .Y(_052_),
    .A1(net75),
    .A2(_286_));
 sg13g2_or2_1 _666_ (.X(_288_),
    .B(_194_),
    .A(_154_));
 sg13g2_nand3_1 _667_ (.B(net146),
    .C(_288_),
    .A(net92),
    .Y(_289_));
 sg13g2_o21ai_1 _668_ (.B1(_289_),
    .Y(_053_),
    .A1(net75),
    .A2(_288_));
 sg13g2_or2_1 _669_ (.X(_290_),
    .B(_194_),
    .A(_140_));
 sg13g2_nand3_1 _670_ (.B(net136),
    .C(_290_),
    .A(net92),
    .Y(_291_));
 sg13g2_o21ai_1 _671_ (.B1(_291_),
    .Y(_054_),
    .A1(net75),
    .A2(_290_));
 sg13g2_nand2b_1 _672_ (.Y(_292_),
    .B(_163_),
    .A_N(_154_));
 sg13g2_nand3_1 _673_ (.B(net122),
    .C(_292_),
    .A(net92),
    .Y(_293_));
 sg13g2_o21ai_1 _674_ (.B1(_293_),
    .Y(_055_),
    .A1(net75),
    .A2(_292_));
 sg13g2_nand2_1 _675_ (.Y(_294_),
    .A(_146_),
    .B(_163_));
 sg13g2_nand3_1 _676_ (.B(net118),
    .C(_294_),
    .A(net93),
    .Y(_295_));
 sg13g2_o21ai_1 _677_ (.B1(_295_),
    .Y(_056_),
    .A1(net76),
    .A2(_294_));
 sg13g2_nand2_1 _678_ (.Y(_296_),
    .A(_146_),
    .B(_172_));
 sg13g2_nand3_1 _679_ (.B(net180),
    .C(_296_),
    .A(net93),
    .Y(_297_));
 sg13g2_o21ai_1 _680_ (.B1(_297_),
    .Y(_057_),
    .A1(net76),
    .A2(_296_));
 sg13g2_nand2_1 _681_ (.Y(_298_),
    .A(_146_),
    .B(_177_));
 sg13g2_nand3_1 _682_ (.B(net187),
    .C(_298_),
    .A(net93),
    .Y(_299_));
 sg13g2_o21ai_1 _683_ (.B1(_299_),
    .Y(_058_),
    .A1(net76),
    .A2(_298_));
 sg13g2_or2_1 _684_ (.X(_300_),
    .B(net227),
    .A(net1));
 sg13g2_nor4_1 _685_ (.A(\u_top.u_mbist.state[5] ),
    .B(net239),
    .C(\u_top.u_mbist.state[3] ),
    .D(net84),
    .Y(_301_));
 sg13g2_nand3_1 _686_ (.B(_111_),
    .C(net240),
    .A(net227),
    .Y(_302_));
 sg13g2_o21ai_1 _687_ (.B1(_300_),
    .Y(_303_),
    .A1(net82),
    .A2(_302_));
 sg13g2_nor3_2 _688_ (.A(\u_top.u_mbist.state[7] ),
    .B(\u_top.u_mbist.state[5] ),
    .C(net82),
    .Y(_304_));
 sg13g2_nor2_1 _689_ (.A(_103_),
    .B(net71),
    .Y(_305_));
 sg13g2_a21oi_1 _690_ (.A1(_091_),
    .A2(_110_),
    .Y(_306_),
    .B1(net80));
 sg13g2_or4_1 _691_ (.A(_002_),
    .B(_303_),
    .C(_305_),
    .D(_306_),
    .X(_307_));
 sg13g2_inv_1 _692_ (.Y(_308_),
    .A(_307_));
 sg13g2_nand2_1 _693_ (.Y(_309_),
    .A(net202),
    .B(_307_));
 sg13g2_nor2_1 _694_ (.A(net83),
    .B(_094_),
    .Y(_310_));
 sg13g2_nand2_2 _695_ (.Y(_311_),
    .A(_091_),
    .B(net71));
 sg13g2_o21ai_1 _696_ (.B1(_308_),
    .Y(_312_),
    .A1(net83),
    .A2(_311_));
 sg13g2_o21ai_1 _697_ (.B1(_309_),
    .Y(_059_),
    .A1(_310_),
    .A2(_312_));
 sg13g2_nand2_1 _698_ (.Y(_313_),
    .A(net150),
    .B(_307_));
 sg13g2_and2_1 _699_ (.A(\u_top.u_mbist.addr[1] ),
    .B(net71),
    .X(_314_));
 sg13g2_xor2_1 _700_ (.B(_304_),
    .A(net150),
    .X(_315_));
 sg13g2_xnor2_1 _701_ (.Y(_316_),
    .A(_094_),
    .B(_315_));
 sg13g2_nor2_1 _702_ (.A(net83),
    .B(_316_),
    .Y(_317_));
 sg13g2_o21ai_1 _703_ (.B1(_313_),
    .Y(_060_),
    .A1(_312_),
    .A2(_317_));
 sg13g2_nand2_1 _704_ (.Y(_318_),
    .A(net169),
    .B(_307_));
 sg13g2_a21oi_1 _705_ (.A1(net202),
    .A2(_315_),
    .Y(_319_),
    .B1(_314_));
 sg13g2_nand2_1 _706_ (.Y(_320_),
    .A(\u_top.u_mbist.addr[2] ),
    .B(net71));
 sg13g2_xnor2_1 _707_ (.Y(_321_),
    .A(net225),
    .B(net71));
 sg13g2_xor2_1 _708_ (.B(_321_),
    .A(_319_),
    .X(_322_));
 sg13g2_nor2_1 _709_ (.A(net83),
    .B(net226),
    .Y(_323_));
 sg13g2_o21ai_1 _710_ (.B1(_318_),
    .Y(_061_),
    .A1(_312_),
    .A2(_323_));
 sg13g2_o21ai_1 _711_ (.B1(_320_),
    .Y(_324_),
    .A1(_319_),
    .A2(_321_));
 sg13g2_nand2_1 _712_ (.Y(_325_),
    .A(net81),
    .B(net71));
 sg13g2_xnor2_1 _713_ (.Y(_326_),
    .A(net81),
    .B(net71));
 sg13g2_xnor2_1 _714_ (.Y(_327_),
    .A(_324_),
    .B(_326_));
 sg13g2_nor2_1 _715_ (.A(net83),
    .B(_327_),
    .Y(_328_));
 sg13g2_nand2_1 _716_ (.Y(_329_),
    .A(net81),
    .B(_307_));
 sg13g2_o21ai_1 _717_ (.B1(_329_),
    .Y(_062_),
    .A1(_312_),
    .A2(_328_));
 sg13g2_o21ai_1 _718_ (.B1(_325_),
    .Y(_330_),
    .A1(_101_),
    .A2(net71));
 sg13g2_a21oi_1 _719_ (.A1(_095_),
    .A2(_324_),
    .Y(_331_),
    .B1(_330_));
 sg13g2_xor2_1 _720_ (.B(_331_),
    .A(net228),
    .X(_332_));
 sg13g2_nor2_1 _721_ (.A(net83),
    .B(_332_),
    .Y(_333_));
 sg13g2_nand2_1 _722_ (.Y(_334_),
    .A(net228),
    .B(_307_));
 sg13g2_o21ai_1 _723_ (.B1(_334_),
    .Y(_063_),
    .A1(_312_),
    .A2(_333_));
 sg13g2_or2_1 _724_ (.X(_335_),
    .B(_150_),
    .A(_147_));
 sg13g2_nand3_1 _725_ (.B(net116),
    .C(_335_),
    .A(net85),
    .Y(_336_));
 sg13g2_o21ai_1 _726_ (.B1(_336_),
    .Y(_064_),
    .A1(net72),
    .A2(_335_));
 sg13g2_or2_1 _727_ (.X(_337_),
    .B(_183_),
    .A(_154_));
 sg13g2_nand3_1 _728_ (.B(net126),
    .C(_337_),
    .A(net85),
    .Y(_338_));
 sg13g2_o21ai_1 _729_ (.B1(_338_),
    .Y(_065_),
    .A1(net72),
    .A2(_337_));
 sg13g2_a21o_1 _730_ (.A2(_214_),
    .A1(net211),
    .B1(_306_),
    .X(_066_));
 sg13g2_or2_1 _731_ (.X(_067_),
    .B(_275_),
    .A(net221));
 sg13g2_a21o_1 _732_ (.A2(done),
    .A1(_009_),
    .B1(net99),
    .X(_068_));
 sg13g2_nand2_1 _733_ (.Y(_339_),
    .A(net202),
    .B(_311_));
 sg13g2_nor3_1 _734_ (.A(\u_top.u_mbist.state[5] ),
    .B(net84),
    .C(_212_),
    .Y(_340_));
 sg13g2_a21o_2 _735_ (.A2(net80),
    .A1(net82),
    .B1(_340_),
    .X(_341_));
 sg13g2_nor2_1 _736_ (.A(net188),
    .B(_311_),
    .Y(_342_));
 sg13g2_nor2_2 _737_ (.A(_341_),
    .B(_342_),
    .Y(_343_));
 sg13g2_a22oi_1 _738_ (.Y(_069_),
    .B1(_343_),
    .B2(_339_),
    .A2(_341_),
    .A1(_085_));
 sg13g2_nand2_1 _739_ (.Y(_344_),
    .A(net150),
    .B(_311_));
 sg13g2_a22oi_1 _740_ (.Y(_070_),
    .B1(_343_),
    .B2(_344_),
    .A2(_341_),
    .A1(_086_));
 sg13g2_nand2_1 _741_ (.Y(_345_),
    .A(net169),
    .B(_311_));
 sg13g2_a22oi_1 _742_ (.Y(_071_),
    .B1(_343_),
    .B2(_345_),
    .A2(_341_),
    .A1(_087_));
 sg13g2_nand2_1 _743_ (.Y(_346_),
    .A(net160),
    .B(_311_));
 sg13g2_a22oi_1 _744_ (.Y(_072_),
    .B1(_343_),
    .B2(net161),
    .A2(_341_),
    .A1(_088_));
 sg13g2_nand2_1 _745_ (.Y(_347_),
    .A(net228),
    .B(_311_));
 sg13g2_a22oi_1 _746_ (.Y(_073_),
    .B1(_343_),
    .B2(_347_),
    .A2(_341_),
    .A1(_089_));
 sg13g2_o21ai_1 _747_ (.B1(_300_),
    .Y(_348_),
    .A1(net80),
    .A2(_111_));
 sg13g2_nor2b_1 _748_ (.A(_348_),
    .B_N(_302_),
    .Y(_349_));
 sg13g2_o21ai_1 _749_ (.B1(_349_),
    .Y(_350_),
    .A1(net204),
    .A2(net83));
 sg13g2_o21ai_1 _750_ (.B1(_350_),
    .Y(_074_),
    .A1(net72),
    .A2(_349_));
 sg13g2_nand2_1 _751_ (.Y(_351_),
    .A(\u_top.bist_mem_rdata[0] ),
    .B(\u_top.u_mbist.state[6] ));
 sg13g2_and2_1 _752_ (.A(_008_),
    .B(_351_),
    .X(_352_));
 sg13g2_or2_1 _753_ (.X(_075_),
    .B(_352_),
    .A(net167));
 sg13g2_a21oi_1 _754_ (.A1(\u_top.u_mbist.state[8] ),
    .A2(net80),
    .Y(_353_),
    .B1(_303_));
 sg13g2_mux2_1 _755_ (.A0(net215),
    .A1(_215_),
    .S(_353_),
    .X(_076_));
 sg13g2_nand2_2 _756_ (.Y(_354_),
    .A(net96),
    .B(_352_));
 sg13g2_nand2_1 _757_ (.Y(_355_),
    .A(net153),
    .B(_354_));
 sg13g2_o21ai_1 _758_ (.B1(_355_),
    .Y(_077_),
    .A1(_096_),
    .A2(_354_));
 sg13g2_nand2_1 _759_ (.Y(_356_),
    .A(\u_top.bist_fail_addr[1] ),
    .B(_354_));
 sg13g2_o21ai_1 _760_ (.B1(_356_),
    .Y(_078_),
    .A1(_097_),
    .A2(_354_));
 sg13g2_nand2_1 _761_ (.Y(_357_),
    .A(\u_top.bist_fail_addr[2] ),
    .B(_354_));
 sg13g2_o21ai_1 _762_ (.B1(_357_),
    .Y(_079_),
    .A1(_098_),
    .A2(_354_));
 sg13g2_mux2_1 _763_ (.A0(net62),
    .A1(net174),
    .S(_354_),
    .X(_080_));
 sg13g2_mux2_1 _764_ (.A0(net129),
    .A1(net190),
    .S(_354_),
    .X(_081_));
 sg13g2_dfrbpq_1 _765_ (.RESET_B(net30),
    .D(net115),
    .Q(\u_top.u_memory.mem_array[8][0] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _766_ (.RESET_B(net57),
    .D(net139),
    .Q(\u_top.u_memory.mem_array[11][0] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _767_ (.RESET_B(net56),
    .D(net104),
    .Q(\u_top.u_memory.mem_array[12][0] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _768_ (.RESET_B(net55),
    .D(_014_),
    .Q(\u_top.u_memory.mem_array[13][0] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _769_ (.RESET_B(net54),
    .D(_015_),
    .Q(\u_top.u_memory.mem_array[27][0] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _770_ (.RESET_B(net53),
    .D(_016_),
    .Q(\u_top.u_memory.mem_array[0][0] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_2 _771_ (.RESET_B(net52),
    .D(net208),
    .Q(\u_top.bist_mem_rdata[0] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_1 _772_ (.RESET_B(net51),
    .D(_018_),
    .Q(\u_top.u_memory.mem_array[2][0] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_2 _773_ (.RESET_B(net88),
    .D(_010_),
    .Q(_009_),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_1 _774_ (.RESET_B(net88),
    .D(_003_),
    .Q(\u_top.u_mbist.state[1] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_1 _775_ (.RESET_B(net90),
    .D(net205),
    .Q(\u_top.u_mbist.state[2] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_2 _776_ (.RESET_B(net88),
    .D(net166),
    .Q(\u_top.u_mbist.state[3] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_2 _777_ (.RESET_B(net89),
    .D(net218),
    .Q(\u_top.u_mbist.state[4] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _778_ (.RESET_B(net90),
    .D(_004_),
    .Q(\u_top.u_mbist.state[5] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_2 _779_ (.RESET_B(net89),
    .D(net220),
    .Q(\u_top.u_mbist.state[6] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_2 _780_ (.RESET_B(net90),
    .D(net157),
    .Q(\u_top.u_mbist.state[7] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_1 _781_ (.RESET_B(net88),
    .D(net189),
    .Q(\u_top.u_mbist.state[8] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_1 _782_ (.RESET_B(net50),
    .D(_019_),
    .Q(\u_top.u_memory.mem_array[30][0] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_1 _783_ (.RESET_B(net89),
    .D(net106),
    .Q(\u_top.u_mbist.read_addr[0] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_1 _784_ (.RESET_B(net96),
    .D(net152),
    .Q(\u_top.u_mbist.read_addr[1] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_1 _785_ (.RESET_B(net89),
    .D(_022_),
    .Q(\u_top.u_mbist.read_addr[2] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_1 _786_ (.RESET_B(net89),
    .D(net63),
    .Q(\u_top.u_mbist.read_addr[3] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_1 _787_ (.RESET_B(net90),
    .D(net130),
    .Q(\u_top.u_mbist.read_addr[4] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_1 _788_ (.RESET_B(net49),
    .D(net108),
    .Q(\u_top.u_memory.mem_array[4][0] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_1 _789_ (.RESET_B(net48),
    .D(net124),
    .Q(\u_top.u_memory.mem_array[5][0] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_1 _790_ (.RESET_B(net47),
    .D(net145),
    .Q(\u_top.u_memory.mem_array[6][0] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_1 _791_ (.RESET_B(net46),
    .D(net113),
    .Q(\u_top.u_memory.mem_array[18][0] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _792_ (.RESET_B(net45),
    .D(net110),
    .Q(\u_top.u_memory.mem_array[10][0] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _793_ (.RESET_B(net43),
    .D(_030_),
    .Q(\u_top.u_memory.mem_array[28][0] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _794_ (.RESET_B(net42),
    .D(net133),
    .Q(\u_top.u_memory.mem_array[16][0] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _795_ (.RESET_B(net40),
    .D(net135),
    .Q(\u_top.u_memory.mem_array[9][0] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_1 _796_ (.RESET_B(net39),
    .D(net102),
    .Q(\u_top.u_memory.mem_array[14][0] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _797_ (.RESET_B(net37),
    .D(net120),
    .Q(\u_top.u_memory.mem_array[23][0] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_1 _798_ (.RESET_B(net36),
    .D(_035_),
    .Q(\u_top.u_memory.mem_array[24][0] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _799_ (.RESET_B(net34),
    .D(_036_),
    .Q(\u_top.u_memory.mem_array[29][0] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _800_ (.RESET_B(net32),
    .D(net98),
    .Q(\u_top.u_memory.mem_array[19][0] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_1 _801_ (.RESET_B(net29),
    .D(_038_),
    .Q(\u_top.u_memory.mem_array[25][0] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _802_ (.RESET_B(net27),
    .D(_039_),
    .Q(\u_top.u_memory.mem_array[26][0] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _803_ (.RESET_B(net94),
    .D(net235),
    .Q(\u_top.u_mbisr.repair_valid[0] [0]),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _804_ (.RESET_B(net95),
    .D(net210),
    .Q(\u_top.u_mbisr.inserted ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _805_ (.RESET_B(net94),
    .D(net198),
    .Q(_358_),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _806_ (.RESET_B(net94),
    .D(net164),
    .Q(_359_),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _807_ (.RESET_B(net94),
    .D(net172),
    .Q(_360_),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _808_ (.RESET_B(net95),
    .D(net178),
    .Q(_361_),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_2 _809_ (.RESET_B(net95),
    .D(net195),
    .Q(_362_),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _810_ (.RESET_B(net94),
    .D(net201),
    .Q(_363_),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _811_ (.RESET_B(net94),
    .D(net183),
    .Q(_364_),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _812_ (.RESET_B(net94),
    .D(net186),
    .Q(_365_),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _813_ (.RESET_B(net96),
    .D(net175),
    .Q(_366_),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _814_ (.RESET_B(net94),
    .D(net191),
    .Q(_367_),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_1 _815_ (.RESET_B(net44),
    .D(net143),
    .Q(\u_top.u_memory.mem_array[22][0] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _816_ (.RESET_B(net41),
    .D(net147),
    .Q(\u_top.u_memory.mem_array[21][0] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _817_ (.RESET_B(net38),
    .D(net137),
    .Q(\u_top.u_memory.mem_array[20][0] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _818_ (.RESET_B(net35),
    .D(_055_),
    .Q(\u_top.u_memory.mem_array[1][0] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _819_ (.RESET_B(net31),
    .D(_056_),
    .Q(\u_top.u_memory.mem_array[3][0] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_1 _820_ (.RESET_B(net26),
    .D(_057_),
    .Q(\u_top.u_memory.mem_array[7][0] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_1 _821_ (.RESET_B(net24),
    .D(_058_),
    .Q(\u_top.u_memory.mem_array[31][0] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_2 _822_ (.RESET_B(net89),
    .D(net203),
    .Q(\u_top.u_mbist.addr[0] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _823_ (.RESET_B(net88),
    .D(_060_),
    .Q(\u_top.u_mbist.addr[1] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _824_ (.RESET_B(net87),
    .D(_061_),
    .Q(\u_top.u_mbist.addr[2] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_1 _825_ (.RESET_B(net88),
    .D(_062_),
    .Q(\u_top.u_mbist.addr[3] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _826_ (.RESET_B(net88),
    .D(_063_),
    .Q(\u_top.u_mbist.addr[4] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_1 _827_ (.RESET_B(net60),
    .D(net117),
    .Q(\u_top.u_memory.mem_array[15][0] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _828_ (.RESET_B(net58),
    .D(net127),
    .Q(\u_top.u_memory.mem_array[17][0] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _829_ (.RESET_B(net90),
    .D(net212),
    .Q(\u_top.u_mbist.read_phase ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_2 _830_ (.RESET_B(net95),
    .D(net222),
    .Q(\u_top.u_mbisr.repair_valid[1] [0]),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_1 _831_ (.RESET_B(net86),
    .D(_406_[0]),
    .Q(\u_top.bist_mem_en ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_1 _832_ (.RESET_B(net88),
    .D(net100),
    .Q(done),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_2 _833_ (.RESET_B(net96),
    .D(net214),
    .Q(\u_top.bist_mem_addr[0] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _834_ (.RESET_B(net96),
    .D(net230),
    .Q(\u_top.bist_mem_addr[1] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _835_ (.RESET_B(net91),
    .D(net237),
    .Q(\u_top.bist_mem_addr[2] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _836_ (.RESET_B(net89),
    .D(net162),
    .Q(\u_top.bist_mem_addr[3] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _837_ (.RESET_B(net96),
    .D(net233),
    .Q(\u_top.bist_mem_addr[4] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_1 _838_ (.RESET_B(net96),
    .D(_008_),
    .Q(\u_top.bist_fail_valid ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_1 _839_ (.RESET_B(net87),
    .D(_074_),
    .Q(\u_top.bist_mem_wdata[0] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_1 _840_ (.RESET_B(net90),
    .D(net168),
    .Q(fail),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_1 _841_ (.RESET_B(net89),
    .D(net216),
    .Q(\u_top.bist_mem_we ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _842_ (.RESET_B(net33),
    .D(net154),
    .Q(\u_top.bist_fail_addr[0] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_2 _843_ (.RESET_B(net28),
    .D(net149),
    .Q(\u_top.bist_fail_addr[1] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_2 _844_ (.RESET_B(net25),
    .D(net159),
    .Q(\u_top.bist_fail_addr[2] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_2 _845_ (.RESET_B(net61),
    .D(_080_),
    .Q(\u_top.bist_fail_addr[3] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _846_ (.RESET_B(net59),
    .D(_081_),
    .Q(\u_top.bist_fail_addr[4] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_tiehi _844__25 (.L_HI(net25));
 sg13g2_tiehi _820__26 (.L_HI(net26));
 sg13g2_tiehi _802__27 (.L_HI(net27));
 sg13g2_tiehi _843__28 (.L_HI(net28));
 sg13g2_tiehi _801__29 (.L_HI(net29));
 sg13g2_tiehi _765__30 (.L_HI(net30));
 sg13g2_tiehi _819__31 (.L_HI(net31));
 sg13g2_tiehi _800__32 (.L_HI(net32));
 sg13g2_tiehi _842__33 (.L_HI(net33));
 sg13g2_tiehi _799__34 (.L_HI(net34));
 sg13g2_tiehi _818__35 (.L_HI(net35));
 sg13g2_tiehi _798__36 (.L_HI(net36));
 sg13g2_tiehi _797__37 (.L_HI(net37));
 sg13g2_tiehi _817__38 (.L_HI(net38));
 sg13g2_tiehi _796__39 (.L_HI(net39));
 sg13g2_tiehi _795__40 (.L_HI(net40));
 sg13g2_tiehi _816__41 (.L_HI(net41));
 sg13g2_tiehi _794__42 (.L_HI(net42));
 sg13g2_tiehi _793__43 (.L_HI(net43));
 sg13g2_tiehi _815__44 (.L_HI(net44));
 sg13g2_tiehi _792__45 (.L_HI(net45));
 sg13g2_tiehi _791__46 (.L_HI(net46));
 sg13g2_tiehi _790__47 (.L_HI(net47));
 sg13g2_tiehi _789__48 (.L_HI(net48));
 sg13g2_tiehi _788__49 (.L_HI(net49));
 sg13g2_tiehi _782__50 (.L_HI(net50));
 sg13g2_tiehi _772__51 (.L_HI(net51));
 sg13g2_tiehi _771__52 (.L_HI(net52));
 sg13g2_tiehi _770__53 (.L_HI(net53));
 sg13g2_tiehi _769__54 (.L_HI(net54));
 sg13g2_tiehi _768__55 (.L_HI(net55));
 sg13g2_tiehi _767__56 (.L_HI(net56));
 sg13g2_tiehi _766__57 (.L_HI(net57));
 sg13g2_tiehi _828__58 (.L_HI(net58));
 sg13g2_tiehi _846__59 (.L_HI(net59));
 sg13g2_tiehi _827__60 (.L_HI(net60));
 sg13g2_tiehi _845__61 (.L_HI(net61));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_aksp_mbist_mbisr_3 (.L_LO(net3));
 sg13g2_tielo tt_um_aksp_mbist_mbisr_4 (.L_LO(net4));
 sg13g2_tielo tt_um_aksp_mbist_mbisr_5 (.L_LO(net5));
 sg13g2_tielo tt_um_aksp_mbist_mbisr_6 (.L_LO(net6));
 sg13g2_tielo tt_um_aksp_mbist_mbisr_7 (.L_LO(net7));
 sg13g2_tielo tt_um_aksp_mbist_mbisr_8 (.L_LO(net8));
 sg13g2_tielo tt_um_aksp_mbist_mbisr_9 (.L_LO(net9));
 sg13g2_tielo tt_um_aksp_mbist_mbisr_10 (.L_LO(net10));
 sg13g2_tielo tt_um_aksp_mbist_mbisr_11 (.L_LO(net11));
 sg13g2_tielo tt_um_aksp_mbist_mbisr_12 (.L_LO(net12));
 sg13g2_tielo tt_um_aksp_mbist_mbisr_13 (.L_LO(net13));
 sg13g2_tielo tt_um_aksp_mbist_mbisr_14 (.L_LO(net14));
 sg13g2_tielo tt_um_aksp_mbist_mbisr_15 (.L_LO(net15));
 sg13g2_tielo tt_um_aksp_mbist_mbisr_16 (.L_LO(net16));
 sg13g2_tielo tt_um_aksp_mbist_mbisr_17 (.L_LO(net17));
 sg13g2_tielo tt_um_aksp_mbist_mbisr_18 (.L_LO(net18));
 sg13g2_tielo tt_um_aksp_mbist_mbisr_19 (.L_LO(net19));
 sg13g2_tielo tt_um_aksp_mbist_mbisr_20 (.L_LO(net20));
 sg13g2_tielo tt_um_aksp_mbist_mbisr_21 (.L_LO(net21));
 sg13g2_tielo tt_um_aksp_mbist_mbisr_22 (.L_LO(net22));
 sg13g2_tielo tt_um_aksp_mbist_mbisr_23 (.L_LO(net23));
 sg13g2_tiehi _821__24 (.L_HI(net24));
 sg13g2_buf_1 _907_ (.A(done),
    .X(uo_out[0]));
 sg13g2_buf_1 _908_ (.A(fail),
    .X(uo_out[1]));
 sg13g2_buf_8 fanout66 (.A(_153_),
    .X(net66));
 sg13g2_buf_8 fanout67 (.A(_139_),
    .X(net67));
 sg13g2_buf_8 fanout68 (.A(_132_),
    .X(net68));
 sg13g2_buf_8 fanout69 (.A(_275_),
    .X(net69));
 sg13g2_buf_8 fanout70 (.A(_253_),
    .X(net70));
 sg13g2_buf_8 fanout71 (.A(_304_),
    .X(net71));
 sg13g2_buf_8 fanout72 (.A(net77),
    .X(net72));
 sg13g2_buf_1 fanout73 (.A(net77),
    .X(net73));
 sg13g2_buf_8 fanout74 (.A(net76),
    .X(net74));
 sg13g2_buf_1 fanout75 (.A(net76),
    .X(net75));
 sg13g2_buf_8 fanout76 (.A(net77),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_082_),
    .X(net77));
 sg13g2_buf_8 fanout78 (.A(net236),
    .X(net78));
 sg13g2_buf_8 fanout79 (.A(net229),
    .X(net79));
 sg13g2_buf_8 fanout80 (.A(net211),
    .X(net80));
 sg13g2_buf_8 fanout81 (.A(net160),
    .X(net81));
 sg13g2_buf_8 fanout82 (.A(net224),
    .X(net82));
 sg13g2_buf_8 fanout83 (.A(net219),
    .X(net83));
 sg13g2_buf_1 fanout84 (.A(net219),
    .X(net84));
 sg13g2_buf_8 fanout85 (.A(net87),
    .X(net85));
 sg13g2_buf_1 fanout86 (.A(net87),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(rst_n),
    .X(net87));
 sg13g2_buf_8 fanout88 (.A(net90),
    .X(net88));
 sg13g2_buf_8 fanout89 (.A(net90),
    .X(net89));
 sg13g2_buf_8 fanout90 (.A(rst_n),
    .X(net90));
 sg13g2_buf_8 fanout91 (.A(net97),
    .X(net91));
 sg13g2_buf_8 fanout92 (.A(net93),
    .X(net92));
 sg13g2_buf_8 fanout93 (.A(net97),
    .X(net93));
 sg13g2_buf_8 fanout94 (.A(net97),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(net96),
    .X(net95));
 sg13g2_buf_8 fanout96 (.A(net97),
    .X(net96));
 sg13g2_buf_8 fanout97 (.A(rst_n),
    .X(net97));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_tielo tt_um_aksp_mbist_mbisr_2 (.L_LO(net2));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_2_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_4_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_12_0_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\u_top.u_mbist.read_addr[3] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold2 (.A(_023_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold3 (.A(\u_top.bist_mem_wdata[0] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold4 (.A(_247_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold5 (.A(_037_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold6 (.A(\u_top.u_mbist.state[1] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold7 (.A(_068_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold8 (.A(\u_top.u_memory.mem_array[14][0] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold9 (.A(_033_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold10 (.A(\u_top.u_memory.mem_array[12][0] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold11 (.A(_013_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold12 (.A(\u_top.u_mbist.read_addr[0] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold13 (.A(_020_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold14 (.A(\u_top.u_memory.mem_array[4][0] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold15 (.A(_025_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold16 (.A(\u_top.u_memory.mem_array[10][0] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold17 (.A(_029_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold18 (.A(\u_top.u_memory.mem_array[13][0] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold19 (.A(\u_top.u_memory.mem_array[18][0] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold20 (.A(_028_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold21 (.A(\u_top.u_memory.mem_array[8][0] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold22 (.A(_011_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold23 (.A(\u_top.u_memory.mem_array[15][0] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold24 (.A(_064_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold25 (.A(\u_top.u_memory.mem_array[3][0] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold26 (.A(\u_top.u_memory.mem_array[23][0] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold27 (.A(_034_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold28 (.A(\u_top.u_memory.mem_array[24][0] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold29 (.A(\u_top.u_memory.mem_array[1][0] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold30 (.A(\u_top.u_memory.mem_array[5][0] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold31 (.A(_026_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold32 (.A(\u_top.u_memory.mem_array[27][0] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold33 (.A(\u_top.u_memory.mem_array[17][0] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold34 (.A(_065_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold35 (.A(\u_top.u_memory.mem_array[26][0] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold36 (.A(\u_top.u_mbist.read_addr[4] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold37 (.A(_024_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold38 (.A(\u_top.u_memory.mem_array[30][0] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold39 (.A(\u_top.u_memory.mem_array[16][0] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold40 (.A(_031_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold41 (.A(\u_top.u_memory.mem_array[9][0] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold42 (.A(_032_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold43 (.A(\u_top.u_memory.mem_array[20][0] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold44 (.A(_054_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold45 (.A(\u_top.u_memory.mem_array[11][0] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold46 (.A(_012_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold47 (.A(\u_top.u_memory.mem_array[25][0] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold48 (.A(\u_top.u_memory.mem_array[0][0] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold49 (.A(\u_top.u_memory.mem_array[22][0] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold50 (.A(_052_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold51 (.A(\u_top.u_memory.mem_array[6][0] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold52 (.A(_027_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold53 (.A(\u_top.u_memory.mem_array[21][0] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold54 (.A(_053_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold55 (.A(\u_top.u_mbist.read_addr[1] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold56 (.A(_078_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold57 (.A(\u_top.u_mbist.addr[1] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold58 (.A(_216_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold59 (.A(_021_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold60 (.A(\u_top.bist_fail_addr[0] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold61 (.A(_077_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold62 (.A(\u_top.u_memory.mem_array[28][0] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold63 (.A(\u_top.u_mbist.state[3] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold64 (.A(_006_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold65 (.A(\u_top.u_mbist.read_addr[2] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold66 (.A(_079_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold67 (.A(\u_top.u_mbist.addr[3] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold68 (.A(_346_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold69 (.A(_072_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold70 (.A(\u_top.bist_fail_addr[1] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold71 (.A(_043_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold72 (.A(\u_top.u_mbist.state[5] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold73 (.A(_001_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold74 (.A(fail),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold75 (.A(_075_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold76 (.A(\u_top.u_mbist.addr[2] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold77 (.A(_217_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold78 (.A(\u_top.bist_fail_addr[2] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold79 (.A(_044_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold80 (.A(\u_top.u_memory.mem_array[2][0] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold81 (.A(\u_top.bist_fail_addr[3] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold82 (.A(_050_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold83 (.A(_361_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold84 (.A(_279_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold85 (.A(_045_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold86 (.A(\u_top.u_memory.mem_array[29][0] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold87 (.A(\u_top.u_memory.mem_array[7][0] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold88 (.A(_364_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold89 (.A(_282_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold90 (.A(_048_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold91 (.A(_365_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold92 (.A(_283_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold93 (.A(_049_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold94 (.A(\u_top.u_memory.mem_array[31][0] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold95 (.A(\u_top.u_mbist.state[4] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold96 (.A(_007_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold97 (.A(\u_top.bist_fail_addr[4] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold98 (.A(_051_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold99 (.A(\u_top.bist_mem_rdata[0] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold100 (.A(_362_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold101 (.A(_280_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold102 (.A(_046_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold103 (.A(_358_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold104 (.A(_276_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold105 (.A(_042_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold106 (.A(_363_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold107 (.A(_281_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold108 (.A(_047_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold109 (.A(\u_top.u_mbist.addr[0] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold110 (.A(_059_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold111 (.A(\u_top.u_mbist.state[7] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold112 (.A(_000_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold113 (.A(\u_top.bist_mem_en ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold114 (.A(_187_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold115 (.A(_017_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold116 (.A(\u_top.u_mbisr.inserted ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold117 (.A(_041_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold118 (.A(\u_top.u_mbist.read_phase ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold119 (.A(_066_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold120 (.A(\u_top.bist_mem_addr[0] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold121 (.A(_069_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold122 (.A(\u_top.bist_mem_we ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold123 (.A(_076_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold124 (.A(\u_top.u_mbist.state[6] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold125 (.A(_002_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold126 (.A(\u_top.u_mbist.state[2] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold127 (.A(_005_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold128 (.A(\u_top.u_mbisr.repair_valid[1] [0]),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold129 (.A(_067_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold130 (.A(\u_top.u_mbist.state[7] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold131 (.A(\u_top.u_mbist.state[8] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold132 (.A(\u_top.u_mbist.addr[2] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold133 (.A(_322_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold134 (.A(_009_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold135 (.A(\u_top.u_mbist.addr[4] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold136 (.A(\u_top.bist_mem_addr[1] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold137 (.A(_070_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold138 (.A(\u_top.u_mbist.addr[1] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold139 (.A(\u_top.bist_mem_addr[4] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold140 (.A(_073_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold141 (.A(\u_top.u_mbisr.repair_valid[0] [0]),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold142 (.A(_040_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold143 (.A(\u_top.bist_mem_addr[2] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold144 (.A(_071_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold145 (.A(\u_top.u_mbist.addr[4] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold146 (.A(\u_top.u_mbist.state[4] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold147 (.A(_301_),
    .X(net240));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_4 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_253 ();
 sg13g2_decap_8 FILLER_15_260 ();
 sg13g2_decap_8 FILLER_15_267 ();
 sg13g2_decap_8 FILLER_15_274 ();
 sg13g2_fill_2 FILLER_15_281 ();
 sg13g2_fill_1 FILLER_15_283 ();
 sg13g2_fill_1 FILLER_15_288 ();
 sg13g2_fill_1 FILLER_15_294 ();
 sg13g2_decap_4 FILLER_15_300 ();
 sg13g2_fill_2 FILLER_15_304 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_334 ();
 sg13g2_decap_8 FILLER_15_341 ();
 sg13g2_decap_8 FILLER_15_348 ();
 sg13g2_decap_8 FILLER_15_355 ();
 sg13g2_decap_8 FILLER_15_362 ();
 sg13g2_decap_8 FILLER_15_369 ();
 sg13g2_decap_8 FILLER_15_376 ();
 sg13g2_decap_8 FILLER_15_383 ();
 sg13g2_decap_8 FILLER_15_390 ();
 sg13g2_decap_8 FILLER_15_397 ();
 sg13g2_decap_4 FILLER_15_404 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_4 FILLER_16_189 ();
 sg13g2_fill_1 FILLER_16_193 ();
 sg13g2_decap_8 FILLER_16_198 ();
 sg13g2_decap_8 FILLER_16_205 ();
 sg13g2_decap_8 FILLER_16_212 ();
 sg13g2_decap_4 FILLER_16_219 ();
 sg13g2_fill_1 FILLER_16_223 ();
 sg13g2_decap_8 FILLER_16_228 ();
 sg13g2_decap_8 FILLER_16_235 ();
 sg13g2_fill_2 FILLER_16_242 ();
 sg13g2_fill_1 FILLER_16_244 ();
 sg13g2_decap_8 FILLER_16_272 ();
 sg13g2_fill_2 FILLER_16_333 ();
 sg13g2_fill_1 FILLER_16_335 ();
 sg13g2_decap_8 FILLER_16_345 ();
 sg13g2_decap_8 FILLER_16_352 ();
 sg13g2_decap_8 FILLER_16_359 ();
 sg13g2_decap_8 FILLER_16_366 ();
 sg13g2_decap_8 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_fill_1 FILLER_17_126 ();
 sg13g2_fill_2 FILLER_17_131 ();
 sg13g2_fill_1 FILLER_17_133 ();
 sg13g2_decap_4 FILLER_17_139 ();
 sg13g2_fill_1 FILLER_17_148 ();
 sg13g2_fill_1 FILLER_17_154 ();
 sg13g2_fill_2 FILLER_17_186 ();
 sg13g2_fill_1 FILLER_17_188 ();
 sg13g2_decap_8 FILLER_17_207 ();
 sg13g2_decap_4 FILLER_17_214 ();
 sg13g2_fill_1 FILLER_17_218 ();
 sg13g2_fill_2 FILLER_17_261 ();
 sg13g2_fill_2 FILLER_17_276 ();
 sg13g2_fill_1 FILLER_17_287 ();
 sg13g2_fill_1 FILLER_17_307 ();
 sg13g2_fill_1 FILLER_17_322 ();
 sg13g2_fill_2 FILLER_17_332 ();
 sg13g2_decap_8 FILLER_17_361 ();
 sg13g2_decap_8 FILLER_17_368 ();
 sg13g2_decap_8 FILLER_17_375 ();
 sg13g2_decap_8 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_4 FILLER_17_403 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_fill_2 FILLER_18_119 ();
 sg13g2_fill_1 FILLER_18_121 ();
 sg13g2_fill_1 FILLER_18_149 ();
 sg13g2_fill_2 FILLER_18_159 ();
 sg13g2_decap_4 FILLER_18_170 ();
 sg13g2_fill_1 FILLER_18_188 ();
 sg13g2_decap_8 FILLER_18_216 ();
 sg13g2_decap_8 FILLER_18_223 ();
 sg13g2_fill_1 FILLER_18_230 ();
 sg13g2_fill_1 FILLER_18_246 ();
 sg13g2_fill_2 FILLER_18_261 ();
 sg13g2_fill_1 FILLER_18_263 ();
 sg13g2_fill_2 FILLER_18_291 ();
 sg13g2_fill_1 FILLER_18_293 ();
 sg13g2_fill_2 FILLER_18_303 ();
 sg13g2_fill_1 FILLER_18_305 ();
 sg13g2_fill_2 FILLER_18_340 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_fill_2 FILLER_19_105 ();
 sg13g2_fill_2 FILLER_19_144 ();
 sg13g2_fill_1 FILLER_19_152 ();
 sg13g2_fill_2 FILLER_19_157 ();
 sg13g2_decap_8 FILLER_19_195 ();
 sg13g2_decap_8 FILLER_19_202 ();
 sg13g2_fill_2 FILLER_19_209 ();
 sg13g2_fill_1 FILLER_19_211 ();
 sg13g2_decap_8 FILLER_19_255 ();
 sg13g2_decap_8 FILLER_19_262 ();
 sg13g2_decap_8 FILLER_19_269 ();
 sg13g2_fill_2 FILLER_19_286 ();
 sg13g2_fill_1 FILLER_19_288 ();
 sg13g2_decap_4 FILLER_19_330 ();
 sg13g2_fill_2 FILLER_19_352 ();
 sg13g2_fill_1 FILLER_19_354 ();
 sg13g2_decap_8 FILLER_19_372 ();
 sg13g2_decap_8 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_19_386 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_fill_2 FILLER_20_105 ();
 sg13g2_fill_1 FILLER_20_107 ();
 sg13g2_decap_4 FILLER_20_144 ();
 sg13g2_fill_2 FILLER_20_161 ();
 sg13g2_fill_1 FILLER_20_163 ();
 sg13g2_fill_2 FILLER_20_174 ();
 sg13g2_fill_1 FILLER_20_176 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_fill_1 FILLER_20_189 ();
 sg13g2_fill_2 FILLER_20_195 ();
 sg13g2_decap_4 FILLER_20_201 ();
 sg13g2_fill_2 FILLER_20_214 ();
 sg13g2_fill_1 FILLER_20_216 ();
 sg13g2_decap_8 FILLER_20_221 ();
 sg13g2_decap_4 FILLER_20_228 ();
 sg13g2_fill_2 FILLER_20_237 ();
 sg13g2_fill_1 FILLER_20_239 ();
 sg13g2_decap_8 FILLER_20_255 ();
 sg13g2_fill_1 FILLER_20_262 ();
 sg13g2_fill_2 FILLER_20_290 ();
 sg13g2_decap_4 FILLER_20_322 ();
 sg13g2_fill_2 FILLER_20_326 ();
 sg13g2_decap_8 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_fill_2 FILLER_21_105 ();
 sg13g2_fill_1 FILLER_21_190 ();
 sg13g2_fill_2 FILLER_21_245 ();
 sg13g2_fill_1 FILLER_21_247 ();
 sg13g2_fill_1 FILLER_21_273 ();
 sg13g2_fill_2 FILLER_21_288 ();
 sg13g2_fill_1 FILLER_21_290 ();
 sg13g2_decap_8 FILLER_21_306 ();
 sg13g2_fill_2 FILLER_21_322 ();
 sg13g2_fill_1 FILLER_21_324 ();
 sg13g2_decap_8 FILLER_21_330 ();
 sg13g2_decap_8 FILLER_21_347 ();
 sg13g2_decap_8 FILLER_21_354 ();
 sg13g2_fill_2 FILLER_21_370 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_fill_2 FILLER_22_109 ();
 sg13g2_fill_1 FILLER_22_111 ();
 sg13g2_fill_2 FILLER_22_125 ();
 sg13g2_fill_2 FILLER_22_177 ();
 sg13g2_fill_2 FILLER_22_184 ();
 sg13g2_fill_2 FILLER_22_195 ();
 sg13g2_fill_1 FILLER_22_197 ();
 sg13g2_decap_8 FILLER_22_206 ();
 sg13g2_decap_8 FILLER_22_213 ();
 sg13g2_fill_2 FILLER_22_220 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_fill_2 FILLER_22_243 ();
 sg13g2_fill_2 FILLER_22_254 ();
 sg13g2_fill_1 FILLER_22_326 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_fill_1 FILLER_23_98 ();
 sg13g2_fill_1 FILLER_23_148 ();
 sg13g2_fill_2 FILLER_23_176 ();
 sg13g2_fill_1 FILLER_23_178 ();
 sg13g2_fill_1 FILLER_23_188 ();
 sg13g2_fill_1 FILLER_23_222 ();
 sg13g2_fill_2 FILLER_23_241 ();
 sg13g2_decap_8 FILLER_23_248 ();
 sg13g2_fill_1 FILLER_23_255 ();
 sg13g2_fill_1 FILLER_23_261 ();
 sg13g2_decap_4 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_297 ();
 sg13g2_decap_4 FILLER_23_304 ();
 sg13g2_fill_1 FILLER_23_313 ();
 sg13g2_decap_8 FILLER_23_324 ();
 sg13g2_decap_8 FILLER_23_331 ();
 sg13g2_fill_1 FILLER_23_353 ();
 sg13g2_fill_2 FILLER_23_367 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_fill_2 FILLER_24_91 ();
 sg13g2_fill_1 FILLER_24_93 ();
 sg13g2_fill_2 FILLER_24_121 ();
 sg13g2_decap_4 FILLER_24_158 ();
 sg13g2_fill_1 FILLER_24_171 ();
 sg13g2_decap_4 FILLER_24_247 ();
 sg13g2_decap_8 FILLER_24_296 ();
 sg13g2_decap_8 FILLER_24_303 ();
 sg13g2_fill_2 FILLER_24_310 ();
 sg13g2_fill_2 FILLER_24_327 ();
 sg13g2_fill_1 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_400 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_fill_1 FILLER_25_112 ();
 sg13g2_fill_2 FILLER_25_204 ();
 sg13g2_fill_1 FILLER_25_244 ();
 sg13g2_fill_2 FILLER_25_250 ();
 sg13g2_fill_2 FILLER_25_257 ();
 sg13g2_fill_1 FILLER_25_259 ();
 sg13g2_fill_2 FILLER_25_277 ();
 sg13g2_decap_4 FILLER_25_288 ();
 sg13g2_fill_2 FILLER_25_292 ();
 sg13g2_fill_2 FILLER_25_299 ();
 sg13g2_fill_1 FILLER_25_301 ();
 sg13g2_decap_4 FILLER_25_324 ();
 sg13g2_fill_1 FILLER_25_328 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_fill_1 FILLER_26_112 ();
 sg13g2_fill_2 FILLER_26_118 ();
 sg13g2_fill_1 FILLER_26_120 ();
 sg13g2_decap_8 FILLER_26_125 ();
 sg13g2_fill_2 FILLER_26_226 ();
 sg13g2_fill_1 FILLER_26_228 ();
 sg13g2_fill_2 FILLER_26_247 ();
 sg13g2_decap_8 FILLER_26_262 ();
 sg13g2_decap_4 FILLER_26_269 ();
 sg13g2_fill_2 FILLER_26_273 ();
 sg13g2_fill_1 FILLER_26_306 ();
 sg13g2_decap_8 FILLER_26_325 ();
 sg13g2_fill_2 FILLER_26_332 ();
 sg13g2_fill_1 FILLER_26_352 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_fill_1 FILLER_27_112 ();
 sg13g2_fill_2 FILLER_27_141 ();
 sg13g2_fill_1 FILLER_27_143 ();
 sg13g2_fill_2 FILLER_27_153 ();
 sg13g2_fill_2 FILLER_27_168 ();
 sg13g2_fill_1 FILLER_27_170 ();
 sg13g2_fill_2 FILLER_27_212 ();
 sg13g2_fill_1 FILLER_27_214 ();
 sg13g2_fill_2 FILLER_27_242 ();
 sg13g2_fill_1 FILLER_27_248 ();
 sg13g2_decap_8 FILLER_27_265 ();
 sg13g2_decap_8 FILLER_27_272 ();
 sg13g2_fill_1 FILLER_27_279 ();
 sg13g2_decap_8 FILLER_27_310 ();
 sg13g2_decap_8 FILLER_27_330 ();
 sg13g2_fill_2 FILLER_27_337 ();
 sg13g2_fill_1 FILLER_27_339 ();
 sg13g2_fill_1 FILLER_27_353 ();
 sg13g2_fill_2 FILLER_27_376 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_4 FILLER_28_84 ();
 sg13g2_fill_1 FILLER_28_96 ();
 sg13g2_fill_2 FILLER_28_118 ();
 sg13g2_fill_1 FILLER_28_120 ();
 sg13g2_decap_8 FILLER_28_130 ();
 sg13g2_decap_8 FILLER_28_137 ();
 sg13g2_fill_2 FILLER_28_144 ();
 sg13g2_decap_8 FILLER_28_153 ();
 sg13g2_decap_8 FILLER_28_160 ();
 sg13g2_fill_1 FILLER_28_167 ();
 sg13g2_fill_2 FILLER_28_205 ();
 sg13g2_fill_2 FILLER_28_291 ();
 sg13g2_decap_4 FILLER_28_306 ();
 sg13g2_fill_2 FILLER_28_310 ();
 sg13g2_decap_8 FILLER_28_326 ();
 sg13g2_fill_2 FILLER_28_333 ();
 sg13g2_fill_1 FILLER_28_335 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_fill_1 FILLER_29_125 ();
 sg13g2_fill_2 FILLER_29_135 ();
 sg13g2_fill_1 FILLER_29_137 ();
 sg13g2_fill_1 FILLER_29_157 ();
 sg13g2_decap_8 FILLER_29_186 ();
 sg13g2_decap_8 FILLER_29_233 ();
 sg13g2_fill_1 FILLER_29_246 ();
 sg13g2_decap_4 FILLER_29_262 ();
 sg13g2_fill_1 FILLER_29_266 ();
 sg13g2_decap_4 FILLER_29_304 ();
 sg13g2_decap_4 FILLER_29_334 ();
 sg13g2_fill_1 FILLER_29_347 ();
 sg13g2_decap_8 FILLER_29_402 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_fill_2 FILLER_30_77 ();
 sg13g2_fill_1 FILLER_30_84 ();
 sg13g2_fill_1 FILLER_30_93 ();
 sg13g2_fill_2 FILLER_30_99 ();
 sg13g2_fill_1 FILLER_30_101 ();
 sg13g2_fill_1 FILLER_30_108 ();
 sg13g2_fill_2 FILLER_30_127 ();
 sg13g2_fill_2 FILLER_30_137 ();
 sg13g2_decap_4 FILLER_30_164 ();
 sg13g2_fill_2 FILLER_30_168 ();
 sg13g2_fill_1 FILLER_30_188 ();
 sg13g2_fill_2 FILLER_30_193 ();
 sg13g2_fill_2 FILLER_30_199 ();
 sg13g2_decap_8 FILLER_30_235 ();
 sg13g2_decap_8 FILLER_30_242 ();
 sg13g2_fill_1 FILLER_30_249 ();
 sg13g2_decap_4 FILLER_30_256 ();
 sg13g2_fill_1 FILLER_30_260 ();
 sg13g2_decap_8 FILLER_30_270 ();
 sg13g2_fill_2 FILLER_30_286 ();
 sg13g2_decap_4 FILLER_30_291 ();
 sg13g2_decap_8 FILLER_30_299 ();
 sg13g2_decap_4 FILLER_30_306 ();
 sg13g2_fill_1 FILLER_30_327 ();
 sg13g2_fill_2 FILLER_30_346 ();
 sg13g2_fill_2 FILLER_30_353 ();
 sg13g2_fill_1 FILLER_30_369 ();
 sg13g2_fill_2 FILLER_30_379 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_fill_2 FILLER_31_49 ();
 sg13g2_fill_1 FILLER_31_51 ();
 sg13g2_fill_2 FILLER_31_141 ();
 sg13g2_fill_1 FILLER_31_143 ();
 sg13g2_decap_4 FILLER_31_251 ();
 sg13g2_fill_1 FILLER_31_255 ();
 sg13g2_decap_4 FILLER_31_284 ();
 sg13g2_fill_1 FILLER_31_288 ();
 sg13g2_fill_2 FILLER_31_298 ();
 sg13g2_fill_1 FILLER_31_317 ();
 sg13g2_fill_1 FILLER_31_322 ();
 sg13g2_decap_4 FILLER_31_332 ();
 sg13g2_fill_1 FILLER_31_336 ();
 sg13g2_fill_2 FILLER_31_361 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_fill_1 FILLER_32_63 ();
 sg13g2_fill_2 FILLER_32_109 ();
 sg13g2_fill_1 FILLER_32_129 ();
 sg13g2_decap_4 FILLER_32_162 ();
 sg13g2_fill_1 FILLER_32_166 ();
 sg13g2_fill_2 FILLER_32_171 ();
 sg13g2_fill_1 FILLER_32_173 ();
 sg13g2_fill_1 FILLER_32_211 ();
 sg13g2_decap_4 FILLER_32_247 ();
 sg13g2_fill_2 FILLER_32_264 ();
 sg13g2_fill_1 FILLER_32_266 ();
 sg13g2_decap_4 FILLER_32_308 ();
 sg13g2_fill_2 FILLER_32_312 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_fill_1 FILLER_33_86 ();
 sg13g2_fill_2 FILLER_33_140 ();
 sg13g2_fill_2 FILLER_33_151 ();
 sg13g2_fill_1 FILLER_33_158 ();
 sg13g2_fill_2 FILLER_33_187 ();
 sg13g2_fill_2 FILLER_33_212 ();
 sg13g2_fill_2 FILLER_33_337 ();
 sg13g2_fill_2 FILLER_33_377 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_fill_1 FILLER_34_77 ();
 sg13g2_fill_2 FILLER_34_101 ();
 sg13g2_fill_2 FILLER_34_129 ();
 sg13g2_fill_1 FILLER_34_146 ();
 sg13g2_fill_1 FILLER_34_176 ();
 sg13g2_fill_2 FILLER_34_244 ();
 sg13g2_decap_4 FILLER_34_258 ();
 sg13g2_decap_4 FILLER_34_266 ();
 sg13g2_fill_1 FILLER_34_270 ();
 sg13g2_decap_8 FILLER_34_306 ();
 sg13g2_fill_2 FILLER_34_313 ();
 sg13g2_fill_2 FILLER_34_329 ();
 sg13g2_fill_1 FILLER_34_331 ();
 sg13g2_fill_1 FILLER_34_355 ();
 sg13g2_fill_1 FILLER_34_396 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_fill_2 FILLER_35_49 ();
 sg13g2_fill_1 FILLER_35_84 ();
 sg13g2_fill_1 FILLER_35_118 ();
 sg13g2_fill_1 FILLER_35_151 ();
 sg13g2_fill_2 FILLER_35_194 ();
 sg13g2_fill_2 FILLER_35_250 ();
 sg13g2_fill_2 FILLER_35_292 ();
 sg13g2_fill_1 FILLER_35_294 ();
 sg13g2_fill_2 FILLER_35_351 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_fill_2 FILLER_36_42 ();
 sg13g2_fill_2 FILLER_36_245 ();
 sg13g2_fill_1 FILLER_36_256 ();
 sg13g2_decap_8 FILLER_36_273 ();
 sg13g2_fill_2 FILLER_36_335 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_fill_2 FILLER_37_67 ();
 sg13g2_fill_1 FILLER_37_69 ();
 sg13g2_fill_2 FILLER_37_79 ();
 sg13g2_fill_2 FILLER_37_110 ();
 sg13g2_fill_2 FILLER_37_158 ();
 sg13g2_fill_1 FILLER_37_160 ();
 sg13g2_fill_1 FILLER_37_178 ();
 sg13g2_fill_2 FILLER_37_219 ();
 sg13g2_fill_2 FILLER_37_248 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_fill_1 FILLER_38_42 ();
 sg13g2_fill_2 FILLER_38_86 ();
 sg13g2_fill_1 FILLER_38_88 ();
 sg13g2_fill_1 FILLER_38_122 ();
 sg13g2_fill_2 FILLER_38_144 ();
 sg13g2_fill_2 FILLER_38_159 ();
 sg13g2_fill_1 FILLER_38_205 ();
 sg13g2_fill_1 FILLER_38_210 ();
 sg13g2_fill_1 FILLER_38_217 ();
 sg13g2_fill_1 FILLER_38_254 ();
 sg13g2_fill_1 FILLER_38_272 ();
 sg13g2_fill_2 FILLER_38_282 ();
 sg13g2_decap_4 FILLER_38_297 ();
 sg13g2_fill_2 FILLER_38_319 ();
 sg13g2_fill_1 FILLER_38_335 ();
 sg13g2_fill_2 FILLER_38_364 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
 assign uo_out[2] = net18;
 assign uo_out[3] = net19;
 assign uo_out[4] = net20;
 assign uo_out[5] = net21;
 assign uo_out[6] = net22;
 assign uo_out[7] = net23;
endmodule
