module tt_um_brmurrell3_m31_accel (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire busy;
 wire mac_mode;
 wire \mul_accum[0] ;
 wire \mul_accum[10] ;
 wire \mul_accum[11] ;
 wire \mul_accum[12] ;
 wire \mul_accum[13] ;
 wire \mul_accum[14] ;
 wire \mul_accum[15] ;
 wire \mul_accum[16] ;
 wire \mul_accum[17] ;
 wire \mul_accum[18] ;
 wire \mul_accum[19] ;
 wire \mul_accum[1] ;
 wire \mul_accum[20] ;
 wire \mul_accum[21] ;
 wire \mul_accum[22] ;
 wire \mul_accum[23] ;
 wire \mul_accum[24] ;
 wire \mul_accum[25] ;
 wire \mul_accum[26] ;
 wire \mul_accum[27] ;
 wire \mul_accum[28] ;
 wire \mul_accum[29] ;
 wire \mul_accum[2] ;
 wire \mul_accum[30] ;
 wire \mul_accum[31] ;
 wire \mul_accum[32] ;
 wire \mul_accum[33] ;
 wire \mul_accum[34] ;
 wire \mul_accum[35] ;
 wire \mul_accum[36] ;
 wire \mul_accum[37] ;
 wire \mul_accum[38] ;
 wire \mul_accum[39] ;
 wire \mul_accum[3] ;
 wire \mul_accum[40] ;
 wire \mul_accum[41] ;
 wire \mul_accum[42] ;
 wire \mul_accum[43] ;
 wire \mul_accum[44] ;
 wire \mul_accum[45] ;
 wire \mul_accum[46] ;
 wire \mul_accum[47] ;
 wire \mul_accum[48] ;
 wire \mul_accum[49] ;
 wire \mul_accum[4] ;
 wire \mul_accum[50] ;
 wire \mul_accum[51] ;
 wire \mul_accum[52] ;
 wire \mul_accum[53] ;
 wire \mul_accum[54] ;
 wire \mul_accum[55] ;
 wire \mul_accum[56] ;
 wire \mul_accum[57] ;
 wire \mul_accum[58] ;
 wire \mul_accum[59] ;
 wire \mul_accum[5] ;
 wire \mul_accum[60] ;
 wire \mul_accum[61] ;
 wire \mul_accum[6] ;
 wire \mul_accum[7] ;
 wire \mul_accum[8] ;
 wire \mul_accum[9] ;
 wire \mul_b_shift[0] ;
 wire \mul_b_shift[10] ;
 wire \mul_b_shift[11] ;
 wire \mul_b_shift[12] ;
 wire \mul_b_shift[13] ;
 wire \mul_b_shift[14] ;
 wire \mul_b_shift[15] ;
 wire \mul_b_shift[16] ;
 wire \mul_b_shift[17] ;
 wire \mul_b_shift[18] ;
 wire \mul_b_shift[19] ;
 wire \mul_b_shift[1] ;
 wire \mul_b_shift[20] ;
 wire \mul_b_shift[21] ;
 wire \mul_b_shift[22] ;
 wire \mul_b_shift[23] ;
 wire \mul_b_shift[24] ;
 wire \mul_b_shift[25] ;
 wire \mul_b_shift[26] ;
 wire \mul_b_shift[27] ;
 wire \mul_b_shift[28] ;
 wire \mul_b_shift[29] ;
 wire \mul_b_shift[2] ;
 wire \mul_b_shift[30] ;
 wire \mul_b_shift[3] ;
 wire \mul_b_shift[4] ;
 wire \mul_b_shift[5] ;
 wire \mul_b_shift[6] ;
 wire \mul_b_shift[7] ;
 wire \mul_b_shift[8] ;
 wire \mul_b_shift[9] ;
 wire \mul_counter[0] ;
 wire \mul_counter[1] ;
 wire \mul_counter[2] ;
 wire \mul_counter[3] ;
 wire \mul_counter[4] ;
 wire \mul_operand_r[0] ;
 wire \mul_operand_r[10] ;
 wire \mul_operand_r[11] ;
 wire \mul_operand_r[12] ;
 wire \mul_operand_r[13] ;
 wire \mul_operand_r[14] ;
 wire \mul_operand_r[15] ;
 wire \mul_operand_r[16] ;
 wire \mul_operand_r[17] ;
 wire \mul_operand_r[18] ;
 wire \mul_operand_r[19] ;
 wire \mul_operand_r[1] ;
 wire \mul_operand_r[20] ;
 wire \mul_operand_r[21] ;
 wire \mul_operand_r[22] ;
 wire \mul_operand_r[23] ;
 wire \mul_operand_r[24] ;
 wire \mul_operand_r[25] ;
 wire \mul_operand_r[26] ;
 wire \mul_operand_r[27] ;
 wire \mul_operand_r[28] ;
 wire \mul_operand_r[29] ;
 wire \mul_operand_r[2] ;
 wire \mul_operand_r[30] ;
 wire \mul_operand_r[3] ;
 wire \mul_operand_r[4] ;
 wire \mul_operand_r[5] ;
 wire \mul_operand_r[6] ;
 wire \mul_operand_r[7] ;
 wire \mul_operand_r[8] ;
 wire \mul_operand_r[9] ;
 wire \read_counter[0] ;
 wire \read_counter[1] ;
 wire reducing;
 wire \reg_a[0] ;
 wire \reg_a[10] ;
 wire \reg_a[11] ;
 wire \reg_a[12] ;
 wire \reg_a[13] ;
 wire \reg_a[14] ;
 wire \reg_a[15] ;
 wire \reg_a[16] ;
 wire \reg_a[17] ;
 wire \reg_a[18] ;
 wire \reg_a[19] ;
 wire \reg_a[1] ;
 wire \reg_a[20] ;
 wire \reg_a[21] ;
 wire \reg_a[22] ;
 wire \reg_a[23] ;
 wire \reg_a[24] ;
 wire \reg_a[25] ;
 wire \reg_a[26] ;
 wire \reg_a[27] ;
 wire \reg_a[28] ;
 wire \reg_a[29] ;
 wire \reg_a[2] ;
 wire \reg_a[30] ;
 wire \reg_a[31] ;
 wire \reg_a[3] ;
 wire \reg_a[4] ;
 wire \reg_a[5] ;
 wire \reg_a[6] ;
 wire \reg_a[7] ;
 wire \reg_a[8] ;
 wire \reg_a[9] ;
 wire \reg_b[0] ;
 wire \reg_b[10] ;
 wire \reg_b[11] ;
 wire \reg_b[12] ;
 wire \reg_b[13] ;
 wire \reg_b[14] ;
 wire \reg_b[15] ;
 wire \reg_b[16] ;
 wire \reg_b[17] ;
 wire \reg_b[18] ;
 wire \reg_b[19] ;
 wire \reg_b[1] ;
 wire \reg_b[20] ;
 wire \reg_b[21] ;
 wire \reg_b[22] ;
 wire \reg_b[23] ;
 wire \reg_b[24] ;
 wire \reg_b[25] ;
 wire \reg_b[26] ;
 wire \reg_b[27] ;
 wire \reg_b[28] ;
 wire \reg_b[29] ;
 wire \reg_b[2] ;
 wire \reg_b[30] ;
 wire \reg_b[31] ;
 wire \reg_b[3] ;
 wire \reg_b[4] ;
 wire \reg_b[5] ;
 wire \reg_b[6] ;
 wire \reg_b[7] ;
 wire \reg_b[8] ;
 wire \reg_b[9] ;
 wire \reg_c[0] ;
 wire \reg_c[10] ;
 wire \reg_c[11] ;
 wire \reg_c[12] ;
 wire \reg_c[13] ;
 wire \reg_c[14] ;
 wire \reg_c[15] ;
 wire \reg_c[16] ;
 wire \reg_c[17] ;
 wire \reg_c[18] ;
 wire \reg_c[19] ;
 wire \reg_c[1] ;
 wire \reg_c[20] ;
 wire \reg_c[21] ;
 wire \reg_c[22] ;
 wire \reg_c[23] ;
 wire \reg_c[24] ;
 wire \reg_c[25] ;
 wire \reg_c[26] ;
 wire \reg_c[27] ;
 wire \reg_c[28] ;
 wire \reg_c[29] ;
 wire \reg_c[2] ;
 wire \reg_c[30] ;
 wire \reg_c[31] ;
 wire \reg_c[3] ;
 wire \reg_c[4] ;
 wire \reg_c[5] ;
 wire \reg_c[6] ;
 wire \reg_c[7] ;
 wire \reg_c[8] ;
 wire \reg_c[9] ;
 wire clknet_leaf_0_clk;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;

 sg13g2_inv_4 _2367_ (.A(\reg_a[25] ),
    .Y(_1922_));
 sg13g2_inv_2 _2368_ (.Y(_1923_),
    .A(\reg_a[17] ));
 sg13g2_inv_1 _2369_ (.Y(_1924_),
    .A(net729));
 sg13g2_inv_2 _2370_ (.Y(_1925_),
    .A(\reg_a[9] ));
 sg13g2_inv_1 _2371_ (.Y(_1926_),
    .A(net731));
 sg13g2_inv_2 _2372_ (.Y(_1927_),
    .A(\reg_a[18] ));
 sg13g2_inv_4 _2373_ (.A(net385),
    .Y(_1928_));
 sg13g2_inv_4 _2374_ (.A(net382),
    .Y(_1929_));
 sg13g2_inv_4 _2375_ (.A(\reg_a[19] ),
    .Y(_1930_));
 sg13g2_inv_4 _2376_ (.A(\reg_a[11] ),
    .Y(_1931_));
 sg13g2_inv_2 _2377_ (.Y(_1932_),
    .A(\reg_a[4] ));
 sg13g2_inv_4 _2378_ (.A(net381),
    .Y(_1933_));
 sg13g2_inv_2 _2379_ (.Y(_1934_),
    .A(\reg_a[6] ));
 sg13g2_inv_4 _2380_ (.A(net390),
    .Y(_1935_));
 sg13g2_inv_2 _2381_ (.Y(_1936_),
    .A(\reg_a[14] ));
 sg13g2_inv_2 _2382_ (.Y(_1937_),
    .A(\reg_a[15] ));
 sg13g2_inv_4 _2383_ (.A(\reg_b[15] ),
    .Y(_1938_));
 sg13g2_inv_1 _2384_ (.Y(_1939_),
    .A(net11));
 sg13g2_inv_4 _2385_ (.A(net706),
    .Y(_1940_));
 sg13g2_inv_1 _2386_ (.Y(_1941_),
    .A(\mul_accum[7] ));
 sg13g2_inv_1 _2387_ (.Y(_1942_),
    .A(\mul_accum[9] ));
 sg13g2_inv_1 _2388_ (.Y(_1943_),
    .A(net255));
 sg13g2_inv_1 _2389_ (.Y(_1944_),
    .A(\mul_accum[24] ));
 sg13g2_inv_1 _2390_ (.Y(_1945_),
    .A(net205));
 sg13g2_inv_1 _2391_ (.Y(_1946_),
    .A(net253));
 sg13g2_inv_1 _2392_ (.Y(_1947_),
    .A(\mul_accum[36] ));
 sg13g2_inv_1 _2393_ (.Y(_1948_),
    .A(\mul_accum[37] ));
 sg13g2_inv_1 _2394_ (.Y(_1949_),
    .A(\mul_accum[38] ));
 sg13g2_inv_1 _2395_ (.Y(_1950_),
    .A(\mul_accum[40] ));
 sg13g2_inv_1 _2396_ (.Y(_1951_),
    .A(\mul_accum[41] ));
 sg13g2_inv_1 _2397_ (.Y(_1952_),
    .A(\mul_accum[42] ));
 sg13g2_inv_1 _2398_ (.Y(_1953_),
    .A(\mul_accum[43] ));
 sg13g2_inv_1 _2399_ (.Y(_1954_),
    .A(net270));
 sg13g2_inv_1 _2400_ (.Y(_1955_),
    .A(\mul_accum[48] ));
 sg13g2_inv_1 _2401_ (.Y(_1956_),
    .A(\mul_accum[49] ));
 sg13g2_inv_1 _2402_ (.Y(_1957_),
    .A(net263));
 sg13g2_inv_1 _2403_ (.Y(_1958_),
    .A(net153));
 sg13g2_inv_2 _2404_ (.Y(_1959_),
    .A(net203));
 sg13g2_inv_2 _2405_ (.Y(_1960_),
    .A(net246));
 sg13g2_inv_1 _2406_ (.Y(_1961_),
    .A(net274));
 sg13g2_inv_2 _2407_ (.Y(_1962_),
    .A(net1));
 sg13g2_inv_1 _2408_ (.Y(_1963_),
    .A(net3));
 sg13g2_inv_2 _2409_ (.Y(_1964_),
    .A(net716));
 sg13g2_nand2_1 _2410_ (.Y(_1965_),
    .A(net721),
    .B(net719));
 sg13g2_nor2_2 _2411_ (.A(net10),
    .B(net765),
    .Y(_1966_));
 sg13g2_nor2b_1 _2412_ (.A(net765),
    .B_N(net10),
    .Y(_1967_));
 sg13g2_nand2_1 _2413_ (.Y(_1968_),
    .A(\reg_b[24] ),
    .B(net755));
 sg13g2_a22oi_1 _2414_ (.Y(_1969_),
    .B1(net761),
    .B2(net735),
    .A2(\reg_c[24] ),
    .A1(net764));
 sg13g2_a21oi_1 _2415_ (.A1(_1968_),
    .A2(_1969_),
    .Y(_1970_),
    .B1(net699));
 sg13g2_a22oi_1 _2416_ (.Y(_1971_),
    .B1(net758),
    .B2(\reg_a[16] ),
    .A2(\reg_c[16] ),
    .A1(net763));
 sg13g2_nand2_1 _2417_ (.Y(_1972_),
    .A(net719),
    .B(_1971_));
 sg13g2_a21oi_1 _2418_ (.A1(\reg_b[16] ),
    .A2(net751),
    .Y(_1973_),
    .B1(_1972_));
 sg13g2_nand2_1 _2419_ (.Y(_1974_),
    .A(net744),
    .B(net759));
 sg13g2_nor2_1 _2420_ (.A(net721),
    .B(_1973_),
    .Y(_1975_));
 sg13g2_a22oi_1 _2421_ (.Y(_1976_),
    .B1(net749),
    .B2(\reg_b[8] ),
    .A2(\reg_c[8] ),
    .A1(net762));
 sg13g2_a21oi_1 _2422_ (.A1(_1974_),
    .A2(_1976_),
    .Y(_1977_),
    .B1(net719));
 sg13g2_nor3_1 _2423_ (.A(_1970_),
    .B(_1975_),
    .C(_1977_),
    .Y(_1978_));
 sg13g2_nand2_1 _2424_ (.Y(_1979_),
    .A(\reg_b[0] ),
    .B(net750));
 sg13g2_or2_1 _2425_ (.X(_1980_),
    .B(net719),
    .A(net301));
 sg13g2_a221oi_1 _2426_ (.B2(\reg_a[0] ),
    .C1(net698),
    .B1(net757),
    .A1(\reg_c[0] ),
    .Y(_1981_),
    .A2(net762));
 sg13g2_a21oi_2 _2427_ (.B1(_1978_),
    .Y(uo_out[0]),
    .A2(_1981_),
    .A1(_1979_));
 sg13g2_nand2_1 _2428_ (.Y(_1982_),
    .A(\reg_b[1] ),
    .B(net750));
 sg13g2_a221oi_1 _2429_ (.B2(net747),
    .C1(net698),
    .B1(net757),
    .A1(net762),
    .Y(_1983_),
    .A2(\reg_c[1] ));
 sg13g2_a22oi_1 _2430_ (.Y(_1984_),
    .B1(net757),
    .B2(\reg_a[9] ),
    .A2(\reg_c[9] ),
    .A1(net762));
 sg13g2_nand2_1 _2431_ (.Y(_1985_),
    .A(net721),
    .B(_1984_));
 sg13g2_a21oi_1 _2432_ (.A1(net731),
    .A2(net751),
    .Y(_1986_),
    .B1(_1985_));
 sg13g2_nor2_1 _2433_ (.A(net719),
    .B(_1986_),
    .Y(_1987_));
 sg13g2_nand2b_2 _2434_ (.Y(_1988_),
    .B(net720),
    .A_N(\read_counter[0] ));
 sg13g2_nand2_1 _2435_ (.Y(_1989_),
    .A(net729),
    .B(net751));
 sg13g2_a22oi_1 _2436_ (.Y(_1990_),
    .B1(net758),
    .B2(\reg_a[17] ),
    .A2(\reg_c[17] ),
    .A1(net763));
 sg13g2_a21oi_1 _2437_ (.A1(_1989_),
    .A2(_1990_),
    .Y(_1991_),
    .B1(_1988_));
 sg13g2_nand2_1 _2438_ (.Y(_1992_),
    .A(net724),
    .B(net755));
 sg13g2_a22oi_1 _2439_ (.Y(_1993_),
    .B1(net760),
    .B2(\reg_a[25] ),
    .A2(\reg_c[25] ),
    .A1(net764));
 sg13g2_a21oi_1 _2440_ (.A1(_1992_),
    .A2(_1993_),
    .Y(_1994_),
    .B1(net699));
 sg13g2_nor3_1 _2441_ (.A(_1987_),
    .B(_1991_),
    .C(_1994_),
    .Y(_1995_));
 sg13g2_a21oi_2 _2442_ (.B1(_1995_),
    .Y(uo_out[1]),
    .A2(_1983_),
    .A1(_1982_));
 sg13g2_a22oi_1 _2443_ (.Y(_1996_),
    .B1(net748),
    .B2(\reg_b[2] ),
    .A2(\reg_c[2] ),
    .A1(net762));
 sg13g2_a21oi_1 _2444_ (.A1(net746),
    .A2(net757),
    .Y(_1997_),
    .B1(net698));
 sg13g2_nand2_1 _2445_ (.Y(_1998_),
    .A(net333),
    .B(net754));
 sg13g2_a22oi_1 _2446_ (.Y(_1999_),
    .B1(net761),
    .B2(net734),
    .A2(\reg_c[26] ),
    .A1(net764));
 sg13g2_a21oi_1 _2447_ (.A1(_1998_),
    .A2(_1999_),
    .Y(_2000_),
    .B1(net699));
 sg13g2_a22oi_1 _2448_ (.Y(_2001_),
    .B1(net758),
    .B2(net743),
    .A2(\reg_c[10] ),
    .A1(net763));
 sg13g2_nand2_1 _2449_ (.Y(_2002_),
    .A(net721),
    .B(_2001_));
 sg13g2_a21oi_1 _2450_ (.A1(\reg_b[10] ),
    .A2(net751),
    .Y(_2003_),
    .B1(_2002_));
 sg13g2_nor2_1 _2451_ (.A(net719),
    .B(_2003_),
    .Y(_2004_));
 sg13g2_nand2_1 _2452_ (.Y(_2005_),
    .A(\reg_a[18] ),
    .B(net760));
 sg13g2_a22oi_1 _2453_ (.Y(_2006_),
    .B1(net753),
    .B2(net728),
    .A2(\reg_c[18] ),
    .A1(net766));
 sg13g2_a21oi_1 _2454_ (.A1(_2005_),
    .A2(_2006_),
    .Y(_2007_),
    .B1(_1988_));
 sg13g2_nor3_1 _2455_ (.A(_2000_),
    .B(_2004_),
    .C(_2007_),
    .Y(_2008_));
 sg13g2_a21oi_2 _2456_ (.B1(_2008_),
    .Y(uo_out[2]),
    .A2(_1997_),
    .A1(_1996_));
 sg13g2_nand2_1 _2457_ (.Y(_2009_),
    .A(\reg_a[19] ),
    .B(net758));
 sg13g2_a22oi_1 _2458_ (.Y(_2010_),
    .B1(net753),
    .B2(net727),
    .A2(\reg_c[19] ),
    .A1(net763));
 sg13g2_a21oi_1 _2459_ (.A1(_2009_),
    .A2(_2010_),
    .Y(_2011_),
    .B1(_1988_));
 sg13g2_a22oi_1 _2460_ (.Y(_2012_),
    .B1(net758),
    .B2(\reg_a[11] ),
    .A2(\reg_c[11] ),
    .A1(net763));
 sg13g2_nand2_1 _2461_ (.Y(_2013_),
    .A(net721),
    .B(_2012_));
 sg13g2_a21oi_1 _2462_ (.A1(\reg_b[11] ),
    .A2(net751),
    .Y(_2014_),
    .B1(_2013_));
 sg13g2_nor2_1 _2463_ (.A(net719),
    .B(_2014_),
    .Y(_2015_));
 sg13g2_nand2_1 _2464_ (.Y(_2016_),
    .A(\reg_a[27] ),
    .B(net760));
 sg13g2_a22oi_1 _2465_ (.Y(_2017_),
    .B1(net756),
    .B2(net723),
    .A2(\reg_c[27] ),
    .A1(net764));
 sg13g2_a21oi_1 _2466_ (.A1(_2016_),
    .A2(_2017_),
    .Y(_2018_),
    .B1(net699));
 sg13g2_nor3_1 _2467_ (.A(_2011_),
    .B(_2015_),
    .C(_2018_),
    .Y(_2019_));
 sg13g2_a22oi_1 _2468_ (.Y(_2020_),
    .B1(net748),
    .B2(\reg_b[3] ),
    .A2(\reg_c[3] ),
    .A1(net762));
 sg13g2_a21oi_1 _2469_ (.A1(\reg_a[3] ),
    .A2(net757),
    .Y(_2021_),
    .B1(net698));
 sg13g2_a21oi_2 _2470_ (.B1(_2019_),
    .Y(uo_out[3]),
    .A2(_2021_),
    .A1(_2020_));
 sg13g2_nand2_1 _2471_ (.Y(_2022_),
    .A(\reg_b[4] ),
    .B(net748));
 sg13g2_a221oi_1 _2472_ (.B2(\reg_a[4] ),
    .C1(net698),
    .B1(net757),
    .A1(net762),
    .Y(_2023_),
    .A2(\reg_c[4] ));
 sg13g2_nand2_1 _2473_ (.Y(_2024_),
    .A(net733),
    .B(net760));
 sg13g2_a22oi_1 _2474_ (.Y(_2025_),
    .B1(net754),
    .B2(\reg_b[28] ),
    .A2(\reg_c[28] ),
    .A1(net764));
 sg13g2_a21oi_1 _2475_ (.A1(_2024_),
    .A2(_2025_),
    .Y(_2026_),
    .B1(net699));
 sg13g2_nand2_1 _2476_ (.Y(_2027_),
    .A(\reg_b[20] ),
    .B(net753));
 sg13g2_a22oi_1 _2477_ (.Y(_2028_),
    .B1(net761),
    .B2(\reg_a[20] ),
    .A2(\reg_c[20] ),
    .A1(net766));
 sg13g2_a21oi_1 _2478_ (.A1(_2027_),
    .A2(_2028_),
    .Y(_2029_),
    .B1(_1988_));
 sg13g2_a22oi_1 _2479_ (.Y(_2030_),
    .B1(net758),
    .B2(net742),
    .A2(\reg_c[12] ),
    .A1(net767));
 sg13g2_nand2_1 _2480_ (.Y(_2031_),
    .A(net721),
    .B(_2030_));
 sg13g2_a21oi_1 _2481_ (.A1(\reg_b[12] ),
    .A2(net751),
    .Y(_2032_),
    .B1(_2031_));
 sg13g2_nor2_1 _2482_ (.A(net719),
    .B(_2032_),
    .Y(_2033_));
 sg13g2_nor3_1 _2483_ (.A(_2026_),
    .B(_2029_),
    .C(_2033_),
    .Y(_2034_));
 sg13g2_a21oi_2 _2484_ (.B1(_2034_),
    .Y(uo_out[4]),
    .A2(_2023_),
    .A1(_2022_));
 sg13g2_nand2_1 _2485_ (.Y(_2035_),
    .A(\reg_a[5] ),
    .B(net759));
 sg13g2_a221oi_1 _2486_ (.B2(\reg_b[5] ),
    .C1(net698),
    .B1(net749),
    .A1(net762),
    .Y(_2036_),
    .A2(\reg_c[5] ));
 sg13g2_a22oi_1 _2487_ (.Y(_2037_),
    .B1(net751),
    .B2(net730),
    .A2(\reg_c[13] ),
    .A1(net767));
 sg13g2_nand2_1 _2488_ (.Y(_2038_),
    .A(net721),
    .B(_2037_));
 sg13g2_a21oi_1 _2489_ (.A1(\reg_a[13] ),
    .A2(net758),
    .Y(_2039_),
    .B1(_2038_));
 sg13g2_nor2_1 _2490_ (.A(net720),
    .B(_2039_),
    .Y(_2040_));
 sg13g2_nand2_1 _2491_ (.Y(_2041_),
    .A(net726),
    .B(net753));
 sg13g2_a22oi_1 _2492_ (.Y(_2042_),
    .B1(net761),
    .B2(net739),
    .A2(\reg_c[21] ),
    .A1(net766));
 sg13g2_a21oi_1 _2493_ (.A1(_2041_),
    .A2(_2042_),
    .Y(_2043_),
    .B1(_1988_));
 sg13g2_nand2_1 _2494_ (.Y(_2044_),
    .A(\reg_a[29] ),
    .B(net761));
 sg13g2_a22oi_1 _2495_ (.Y(_2045_),
    .B1(net754),
    .B2(net722),
    .A2(\reg_c[29] ),
    .A1(net764));
 sg13g2_a21oi_1 _2496_ (.A1(_2044_),
    .A2(_2045_),
    .Y(_2046_),
    .B1(net699));
 sg13g2_nor3_1 _2497_ (.A(_2040_),
    .B(_2043_),
    .C(_2046_),
    .Y(_2047_));
 sg13g2_a21oi_2 _2498_ (.B1(_2047_),
    .Y(uo_out[5]),
    .A2(_2036_),
    .A1(_2035_));
 sg13g2_a22oi_1 _2499_ (.Y(_2048_),
    .B1(net757),
    .B2(\reg_a[6] ),
    .A2(\reg_c[6] ),
    .A1(net763));
 sg13g2_a21oi_1 _2500_ (.A1(\reg_b[6] ),
    .A2(net749),
    .Y(_2049_),
    .B1(net698));
 sg13g2_a22oi_1 _2501_ (.Y(_2050_),
    .B1(net759),
    .B2(\reg_a[14] ),
    .A2(\reg_c[14] ),
    .A1(net767));
 sg13g2_nand2_1 _2502_ (.Y(_2051_),
    .A(\read_counter[0] ),
    .B(_2050_));
 sg13g2_a21oi_1 _2503_ (.A1(\reg_b[14] ),
    .A2(net753),
    .Y(_2052_),
    .B1(_2051_));
 sg13g2_nor2_1 _2504_ (.A(net720),
    .B(_2052_),
    .Y(_2053_));
 sg13g2_nand2_1 _2505_ (.Y(_2054_),
    .A(\reg_b[22] ),
    .B(net753));
 sg13g2_a22oi_1 _2506_ (.Y(_2055_),
    .B1(net761),
    .B2(net738),
    .A2(\reg_c[22] ),
    .A1(net766));
 sg13g2_a21oi_1 _2507_ (.A1(_2054_),
    .A2(_2055_),
    .Y(_2056_),
    .B1(_1988_));
 sg13g2_nand2_1 _2508_ (.Y(_2057_),
    .A(\reg_a[30] ),
    .B(net760));
 sg13g2_a22oi_1 _2509_ (.Y(_2058_),
    .B1(net755),
    .B2(\reg_b[30] ),
    .A2(\reg_c[30] ),
    .A1(net764));
 sg13g2_a21oi_1 _2510_ (.A1(_2057_),
    .A2(_2058_),
    .Y(_2059_),
    .B1(net699));
 sg13g2_nor3_1 _2511_ (.A(_2053_),
    .B(_2056_),
    .C(_2059_),
    .Y(_2060_));
 sg13g2_a21oi_2 _2512_ (.B1(_2060_),
    .Y(uo_out[6]),
    .A2(_2049_),
    .A1(_2048_));
 sg13g2_a22oi_1 _2513_ (.Y(_2061_),
    .B1(net749),
    .B2(\reg_b[7] ),
    .A2(\reg_c[7] ),
    .A1(net763));
 sg13g2_a21oi_1 _2514_ (.A1(net745),
    .A2(net757),
    .Y(_2062_),
    .B1(net698));
 sg13g2_and2_1 _2515_ (.A(net37),
    .B(net754),
    .X(_2063_));
 sg13g2_a221oi_1 _2516_ (.B2(\reg_a[31] ),
    .C1(_2063_),
    .B1(net761),
    .A1(net764),
    .Y(_2064_),
    .A2(\reg_c[31] ));
 sg13g2_o21ai_1 _2517_ (.B1(_1980_),
    .Y(_2065_),
    .A1(_1965_),
    .A2(_2064_));
 sg13g2_nand2_1 _2518_ (.Y(_2066_),
    .A(net736),
    .B(net760));
 sg13g2_a22oi_1 _2519_ (.Y(_2067_),
    .B1(net753),
    .B2(net725),
    .A2(\reg_c[23] ),
    .A1(net766));
 sg13g2_a21oi_1 _2520_ (.A1(_2066_),
    .A2(_2067_),
    .Y(_2068_),
    .B1(_1988_));
 sg13g2_nand2_1 _2521_ (.Y(_2069_),
    .A(\reg_a[15] ),
    .B(net759));
 sg13g2_a22oi_1 _2522_ (.Y(_2070_),
    .B1(net753),
    .B2(\reg_b[15] ),
    .A2(\reg_c[15] ),
    .A1(net766));
 sg13g2_a21oi_1 _2523_ (.A1(_2069_),
    .A2(_2070_),
    .Y(_2071_),
    .B1(net720));
 sg13g2_nor3_1 _2524_ (.A(_2065_),
    .B(_2068_),
    .C(_2071_),
    .Y(_2072_));
 sg13g2_a21oi_2 _2525_ (.B1(_2072_),
    .Y(uo_out[7]),
    .A2(_2062_),
    .A1(_2061_));
 sg13g2_nor3_1 _2526_ (.A(net721),
    .B(_1939_),
    .C(net9),
    .Y(_0000_));
 sg13g2_nand3_1 _2527_ (.B(net699),
    .C(_1980_),
    .A(net11),
    .Y(_2073_));
 sg13g2_nor2_1 _2528_ (.A(net9),
    .B(_2073_),
    .Y(_0001_));
 sg13g2_nor4_1 _2529_ (.A(net209),
    .B(net30),
    .C(net28),
    .D(net38),
    .Y(_2074_));
 sg13g2_nor2b_1 _2530_ (.A(net27),
    .B_N(_2074_),
    .Y(_2075_));
 sg13g2_nand2b_1 _2531_ (.Y(_2076_),
    .B(_2074_),
    .A_N(\mul_counter[0] ));
 sg13g2_nor2_1 _2532_ (.A(net704),
    .B(net684),
    .Y(_2077_));
 sg13g2_inv_2 _2533_ (.Y(busy),
    .A(net653));
 sg13g2_nor3_1 _2534_ (.A(net11),
    .B(net9),
    .C(busy),
    .Y(_2078_));
 sg13g2_nand3b_1 _2535_ (.B(net765),
    .C(net591),
    .Y(_2079_),
    .A_N(net10));
 sg13g2_nor2_1 _2536_ (.A(\reg_c[8] ),
    .B(net584),
    .Y(_2080_));
 sg13g2_nand2_1 _2537_ (.Y(_2081_),
    .A(net765),
    .B(net591));
 sg13g2_nor2_2 _2538_ (.A(net10),
    .B(_2081_),
    .Y(_2082_));
 sg13g2_nor2_1 _2539_ (.A(net159),
    .B(net565),
    .Y(_2083_));
 sg13g2_nor3_1 _2540_ (.A(net2),
    .B(net4),
    .C(_1963_),
    .Y(_2084_));
 sg13g2_and2_1 _2541_ (.A(_1962_),
    .B(_2084_),
    .X(_2085_));
 sg13g2_nor2b_2 _2542_ (.A(net705),
    .B_N(net9),
    .Y(_2086_));
 sg13g2_and3_1 _2543_ (.X(_2087_),
    .A(net696),
    .B(_2085_),
    .C(_2086_));
 sg13g2_nor3_1 _2544_ (.A(_2080_),
    .B(_2083_),
    .C(net640),
    .Y(_0066_));
 sg13g2_nor2_1 _2545_ (.A(\reg_c[9] ),
    .B(net584),
    .Y(_2088_));
 sg13g2_nor2_1 _2546_ (.A(net71),
    .B(net565),
    .Y(_2089_));
 sg13g2_nor3_1 _2547_ (.A(net640),
    .B(_2088_),
    .C(_2089_),
    .Y(_0077_));
 sg13g2_nor2_1 _2548_ (.A(\reg_c[10] ),
    .B(net584),
    .Y(_2090_));
 sg13g2_nor2_1 _2549_ (.A(net172),
    .B(net565),
    .Y(_2091_));
 sg13g2_nor3_1 _2550_ (.A(net640),
    .B(_2090_),
    .C(_2091_),
    .Y(_0088_));
 sg13g2_nor2_1 _2551_ (.A(\reg_c[11] ),
    .B(net584),
    .Y(_2092_));
 sg13g2_nor2_1 _2552_ (.A(net78),
    .B(net566),
    .Y(_2093_));
 sg13g2_nor3_1 _2553_ (.A(net641),
    .B(_2092_),
    .C(_2093_),
    .Y(_0091_));
 sg13g2_nor2_1 _2554_ (.A(\reg_c[12] ),
    .B(net584),
    .Y(_2094_));
 sg13g2_nor2_1 _2555_ (.A(net126),
    .B(net565),
    .Y(_2095_));
 sg13g2_nor3_1 _2556_ (.A(net640),
    .B(_2094_),
    .C(_2095_),
    .Y(_0092_));
 sg13g2_nor2_1 _2557_ (.A(net182),
    .B(net584),
    .Y(_2096_));
 sg13g2_nor2_1 _2558_ (.A(net196),
    .B(net565),
    .Y(_2097_));
 sg13g2_nor3_1 _2559_ (.A(net641),
    .B(_2096_),
    .C(_2097_),
    .Y(_0093_));
 sg13g2_nor2_1 _2560_ (.A(\reg_c[14] ),
    .B(net585),
    .Y(_2098_));
 sg13g2_nor2_1 _2561_ (.A(net113),
    .B(net566),
    .Y(_2099_));
 sg13g2_nor3_1 _2562_ (.A(net641),
    .B(_2098_),
    .C(_2099_),
    .Y(_0094_));
 sg13g2_nor2_1 _2563_ (.A(\reg_c[15] ),
    .B(net585),
    .Y(_2100_));
 sg13g2_nor2_1 _2564_ (.A(net142),
    .B(net566),
    .Y(_2101_));
 sg13g2_nor3_1 _2565_ (.A(net642),
    .B(_2100_),
    .C(_2101_),
    .Y(_0095_));
 sg13g2_nor2_1 _2566_ (.A(net225),
    .B(net585),
    .Y(_2102_));
 sg13g2_nor2_1 _2567_ (.A(net278),
    .B(net565),
    .Y(_2103_));
 sg13g2_nor3_1 _2568_ (.A(net642),
    .B(_2102_),
    .C(_2103_),
    .Y(_0096_));
 sg13g2_nor2_1 _2569_ (.A(\reg_c[17] ),
    .B(net584),
    .Y(_2104_));
 sg13g2_nor2_1 _2570_ (.A(net115),
    .B(net565),
    .Y(_2105_));
 sg13g2_nor3_1 _2571_ (.A(net640),
    .B(_2104_),
    .C(_2105_),
    .Y(_0097_));
 sg13g2_nor2_1 _2572_ (.A(net232),
    .B(net585),
    .Y(_2106_));
 sg13g2_nor2_1 _2573_ (.A(net248),
    .B(net566),
    .Y(_2107_));
 sg13g2_nor3_1 _2574_ (.A(net642),
    .B(_2106_),
    .C(_2107_),
    .Y(_0067_));
 sg13g2_nor2_1 _2575_ (.A(net212),
    .B(net585),
    .Y(_2108_));
 sg13g2_nor2_1 _2576_ (.A(net233),
    .B(net565),
    .Y(_2109_));
 sg13g2_nor3_1 _2577_ (.A(net642),
    .B(_2108_),
    .C(_2109_),
    .Y(_0068_));
 sg13g2_nor2_1 _2578_ (.A(net201),
    .B(net584),
    .Y(_2110_));
 sg13g2_nor2_1 _2579_ (.A(net216),
    .B(net566),
    .Y(_2111_));
 sg13g2_nor3_1 _2580_ (.A(net642),
    .B(_2110_),
    .C(_2111_),
    .Y(_0069_));
 sg13g2_nor2_1 _2581_ (.A(\reg_c[21] ),
    .B(net585),
    .Y(_2112_));
 sg13g2_nor2_1 _2582_ (.A(net182),
    .B(net566),
    .Y(_2113_));
 sg13g2_nor3_1 _2583_ (.A(net650),
    .B(_2112_),
    .C(_2113_),
    .Y(_0070_));
 sg13g2_nor2_1 _2584_ (.A(net184),
    .B(net588),
    .Y(_2114_));
 sg13g2_nor2_1 _2585_ (.A(net219),
    .B(net569),
    .Y(_2115_));
 sg13g2_nor3_1 _2586_ (.A(net650),
    .B(_2114_),
    .C(_2115_),
    .Y(_0071_));
 sg13g2_nor2_1 _2587_ (.A(net146),
    .B(net588),
    .Y(_2116_));
 sg13g2_nor2_1 _2588_ (.A(net187),
    .B(net569),
    .Y(_2117_));
 sg13g2_nor3_1 _2589_ (.A(net650),
    .B(_2116_),
    .C(_2117_),
    .Y(_0072_));
 sg13g2_nor2_1 _2590_ (.A(\reg_c[24] ),
    .B(net588),
    .Y(_2118_));
 sg13g2_nor2_1 _2591_ (.A(net225),
    .B(net569),
    .Y(_2119_));
 sg13g2_nor3_1 _2592_ (.A(net650),
    .B(_2118_),
    .C(_2119_),
    .Y(_0073_));
 sg13g2_nor2_1 _2593_ (.A(net177),
    .B(net586),
    .Y(_2120_));
 sg13g2_nor2_1 _2594_ (.A(net269),
    .B(net569),
    .Y(_2121_));
 sg13g2_nor3_1 _2595_ (.A(net648),
    .B(_2120_),
    .C(_2121_),
    .Y(_0074_));
 sg13g2_nor2_1 _2596_ (.A(net220),
    .B(net587),
    .Y(_2122_));
 sg13g2_nor2_1 _2597_ (.A(net232),
    .B(net568),
    .Y(_2123_));
 sg13g2_nor3_1 _2598_ (.A(net649),
    .B(_2122_),
    .C(_2123_),
    .Y(_0075_));
 sg13g2_nor2_1 _2599_ (.A(\reg_c[27] ),
    .B(net587),
    .Y(_2124_));
 sg13g2_nor2_1 _2600_ (.A(net212),
    .B(net568),
    .Y(_2125_));
 sg13g2_nor3_1 _2601_ (.A(net649),
    .B(_2124_),
    .C(_2125_),
    .Y(_0076_));
 sg13g2_nor2_1 _2602_ (.A(net150),
    .B(net586),
    .Y(_2126_));
 sg13g2_nor2_1 _2603_ (.A(net201),
    .B(net567),
    .Y(_2127_));
 sg13g2_nor3_1 _2604_ (.A(net648),
    .B(_2126_),
    .C(_2127_),
    .Y(_0078_));
 sg13g2_nor2_1 _2605_ (.A(net156),
    .B(net586),
    .Y(_2128_));
 sg13g2_nor2_1 _2606_ (.A(net202),
    .B(net567),
    .Y(_2129_));
 sg13g2_nor3_1 _2607_ (.A(net648),
    .B(_2128_),
    .C(_2129_),
    .Y(_0079_));
 sg13g2_nor2_1 _2608_ (.A(net139),
    .B(net586),
    .Y(_2130_));
 sg13g2_nor2_1 _2609_ (.A(net184),
    .B(net567),
    .Y(_2131_));
 sg13g2_nor3_1 _2610_ (.A(net649),
    .B(_2130_),
    .C(_2131_),
    .Y(_0080_));
 sg13g2_nor2_1 _2611_ (.A(\reg_c[31] ),
    .B(net587),
    .Y(_2132_));
 sg13g2_nor2_1 _2612_ (.A(net146),
    .B(net568),
    .Y(_2133_));
 sg13g2_nor3_1 _2613_ (.A(net651),
    .B(_2132_),
    .C(_2133_),
    .Y(_0081_));
 sg13g2_nor2_1 _2614_ (.A(net1),
    .B(net587),
    .Y(_2134_));
 sg13g2_nor2_1 _2615_ (.A(net231),
    .B(net567),
    .Y(_2135_));
 sg13g2_nor3_1 _2616_ (.A(net649),
    .B(_2134_),
    .C(_2135_),
    .Y(_0082_));
 sg13g2_nor2_1 _2617_ (.A(net2),
    .B(net586),
    .Y(_2136_));
 sg13g2_nor2_1 _2618_ (.A(net177),
    .B(net567),
    .Y(_2137_));
 sg13g2_nor3_1 _2619_ (.A(net648),
    .B(_2136_),
    .C(_2137_),
    .Y(_0083_));
 sg13g2_nor2_1 _2620_ (.A(net3),
    .B(net587),
    .Y(_2138_));
 sg13g2_nor2_1 _2621_ (.A(net220),
    .B(net568),
    .Y(_2139_));
 sg13g2_nor3_1 _2622_ (.A(net649),
    .B(_2138_),
    .C(_2139_),
    .Y(_0084_));
 sg13g2_nor2_1 _2623_ (.A(net4),
    .B(net587),
    .Y(_2140_));
 sg13g2_nor2_1 _2624_ (.A(net236),
    .B(net568),
    .Y(_2141_));
 sg13g2_nor3_1 _2625_ (.A(net649),
    .B(_2140_),
    .C(_2141_),
    .Y(_0085_));
 sg13g2_nor2_1 _2626_ (.A(net5),
    .B(net586),
    .Y(_2142_));
 sg13g2_nor2_1 _2627_ (.A(net150),
    .B(net567),
    .Y(_2143_));
 sg13g2_nor3_1 _2628_ (.A(net645),
    .B(_2142_),
    .C(_2143_),
    .Y(_0086_));
 sg13g2_nor2_1 _2629_ (.A(net6),
    .B(net586),
    .Y(_2144_));
 sg13g2_nor2_1 _2630_ (.A(net156),
    .B(net567),
    .Y(_2145_));
 sg13g2_nor3_1 _2631_ (.A(net648),
    .B(_2144_),
    .C(_2145_),
    .Y(_0087_));
 sg13g2_nor2_1 _2632_ (.A(net7),
    .B(net586),
    .Y(_2146_));
 sg13g2_nor2_1 _2633_ (.A(net139),
    .B(net567),
    .Y(_2147_));
 sg13g2_nor3_1 _2634_ (.A(net648),
    .B(_2146_),
    .C(_2147_),
    .Y(_0089_));
 sg13g2_nor2_1 _2635_ (.A(net8),
    .B(net587),
    .Y(_2148_));
 sg13g2_nor2_1 _2636_ (.A(net155),
    .B(net568),
    .Y(_2149_));
 sg13g2_nor3_1 _2637_ (.A(net649),
    .B(_2148_),
    .C(_2149_),
    .Y(_0090_));
 sg13g2_and2_1 _2638_ (.A(net754),
    .B(net592),
    .X(_2150_));
 sg13g2_nand2_2 _2639_ (.Y(_2151_),
    .A(net748),
    .B(net589));
 sg13g2_nand2_1 _2640_ (.Y(_2152_),
    .A(net249),
    .B(net580));
 sg13g2_nand3_1 _2641_ (.B(net750),
    .C(net589),
    .A(\reg_b[8] ),
    .Y(_2153_));
 sg13g2_a21oi_1 _2642_ (.A1(_2152_),
    .A2(_2153_),
    .Y(_0034_),
    .B1(net644));
 sg13g2_nand2_1 _2643_ (.Y(_2154_),
    .A(net256),
    .B(net580));
 sg13g2_nand3_1 _2644_ (.B(net750),
    .C(net589),
    .A(net731),
    .Y(_2155_));
 sg13g2_a21oi_1 _2645_ (.A1(_2154_),
    .A2(_2155_),
    .Y(_0045_),
    .B1(net644));
 sg13g2_nand2_1 _2646_ (.Y(_2156_),
    .A(net260),
    .B(net580));
 sg13g2_nand3_1 _2647_ (.B(net750),
    .C(net589),
    .A(\reg_b[10] ),
    .Y(_2157_));
 sg13g2_a21oi_1 _2648_ (.A1(_2156_),
    .A2(_2157_),
    .Y(_0056_),
    .B1(net644));
 sg13g2_nand2_1 _2649_ (.Y(_2158_),
    .A(net322),
    .B(net579));
 sg13g2_nand3_1 _2650_ (.B(net748),
    .C(net590),
    .A(\reg_b[11] ),
    .Y(_2159_));
 sg13g2_a21oi_1 _2651_ (.A1(_2158_),
    .A2(_2159_),
    .Y(_0059_),
    .B1(net641));
 sg13g2_nand2_1 _2652_ (.Y(_2160_),
    .A(net318),
    .B(net579));
 sg13g2_nand3_1 _2653_ (.B(net748),
    .C(net590),
    .A(\reg_b[12] ),
    .Y(_2161_));
 sg13g2_a21oi_1 _2654_ (.A1(_2160_),
    .A2(_2161_),
    .Y(_0060_),
    .B1(net640));
 sg13g2_nand2_1 _2655_ (.Y(_2162_),
    .A(net358),
    .B(net579));
 sg13g2_nand3_1 _2656_ (.B(net748),
    .C(net590),
    .A(net730),
    .Y(_2163_));
 sg13g2_a21oi_1 _2657_ (.A1(_2162_),
    .A2(_2163_),
    .Y(_0061_),
    .B1(net641));
 sg13g2_nand2_1 _2658_ (.Y(_2164_),
    .A(net345),
    .B(net579));
 sg13g2_nand3_1 _2659_ (.B(net748),
    .C(net590),
    .A(\reg_b[14] ),
    .Y(_2165_));
 sg13g2_a21oi_1 _2660_ (.A1(_2164_),
    .A2(_2165_),
    .Y(_0062_),
    .B1(net640));
 sg13g2_nand2_1 _2661_ (.Y(_2166_),
    .A(net347),
    .B(net579));
 sg13g2_nand3_1 _2662_ (.B(net752),
    .C(net590),
    .A(net262),
    .Y(_2167_));
 sg13g2_a21oi_1 _2663_ (.A1(_2166_),
    .A2(_2167_),
    .Y(_0063_),
    .B1(net641));
 sg13g2_nand2_1 _2664_ (.Y(_2168_),
    .A(net311),
    .B(net579));
 sg13g2_nand3_1 _2665_ (.B(net750),
    .C(net589),
    .A(\reg_b[16] ),
    .Y(_2169_));
 sg13g2_a21oi_1 _2666_ (.A1(_2168_),
    .A2(_2169_),
    .Y(_0064_),
    .B1(net640));
 sg13g2_nand2_1 _2667_ (.Y(_2170_),
    .A(net731),
    .B(net580));
 sg13g2_nand2b_1 _2668_ (.Y(_2171_),
    .B(net589),
    .A_N(_1989_));
 sg13g2_a21oi_1 _2669_ (.A1(_2170_),
    .A2(_2171_),
    .Y(_0065_),
    .B1(net644));
 sg13g2_nand2_1 _2670_ (.Y(_2172_),
    .A(net327),
    .B(net579));
 sg13g2_nand3_1 _2671_ (.B(net752),
    .C(net589),
    .A(net728),
    .Y(_2173_));
 sg13g2_a21oi_1 _2672_ (.A1(_2172_),
    .A2(_2173_),
    .Y(_0035_),
    .B1(net642));
 sg13g2_nand2_1 _2673_ (.Y(_2174_),
    .A(net343),
    .B(net579));
 sg13g2_nand3_1 _2674_ (.B(net751),
    .C(net589),
    .A(net727),
    .Y(_2175_));
 sg13g2_a21oi_1 _2675_ (.A1(_2174_),
    .A2(_2175_),
    .Y(_0036_),
    .B1(net643));
 sg13g2_nand2_1 _2676_ (.Y(_2176_),
    .A(net338),
    .B(net580));
 sg13g2_nand2b_1 _2677_ (.Y(_2177_),
    .B(net591),
    .A_N(_2027_));
 sg13g2_a21oi_1 _2678_ (.A1(_2176_),
    .A2(_2177_),
    .Y(_0037_),
    .B1(net642));
 sg13g2_nand2_1 _2679_ (.Y(_2178_),
    .A(net730),
    .B(net580));
 sg13g2_nand2b_1 _2680_ (.Y(_2179_),
    .B(net591),
    .A_N(_2041_));
 sg13g2_a21oi_1 _2681_ (.A1(_2178_),
    .A2(_2179_),
    .Y(_0038_),
    .B1(net642));
 sg13g2_nand2_1 _2682_ (.Y(_2180_),
    .A(net353),
    .B(net583));
 sg13g2_nand2b_1 _2683_ (.Y(_2181_),
    .B(net592),
    .A_N(_2054_));
 sg13g2_a21oi_1 _2684_ (.A1(_2180_),
    .A2(_2181_),
    .Y(_0039_),
    .B1(net647));
 sg13g2_nand2_1 _2685_ (.Y(_2182_),
    .A(net262),
    .B(net583));
 sg13g2_nand3_1 _2686_ (.B(net756),
    .C(net591),
    .A(net725),
    .Y(_2183_));
 sg13g2_a21oi_1 _2687_ (.A1(_2182_),
    .A2(_2183_),
    .Y(_0040_),
    .B1(net650));
 sg13g2_nand2_1 _2688_ (.Y(_2184_),
    .A(net340),
    .B(net583));
 sg13g2_nand2b_1 _2689_ (.Y(_2185_),
    .B(net591),
    .A_N(_1968_));
 sg13g2_a21oi_1 _2690_ (.A1(_2184_),
    .A2(_2185_),
    .Y(_0041_),
    .B1(net650));
 sg13g2_nand2_1 _2691_ (.Y(_2186_),
    .A(net729),
    .B(net582));
 sg13g2_nand2b_1 _2692_ (.Y(_2187_),
    .B(net592),
    .A_N(_1992_));
 sg13g2_a21oi_1 _2693_ (.A1(_2186_),
    .A2(_2187_),
    .Y(_0042_),
    .B1(net647));
 sg13g2_nand2_1 _2694_ (.Y(_2188_),
    .A(net728),
    .B(net583));
 sg13g2_nand2b_1 _2695_ (.Y(_2189_),
    .B(net591),
    .A_N(_1998_));
 sg13g2_a21oi_1 _2696_ (.A1(_2188_),
    .A2(_2189_),
    .Y(_0043_),
    .B1(net650));
 sg13g2_nand2_1 _2697_ (.Y(_2190_),
    .A(net727),
    .B(net583));
 sg13g2_nand3_1 _2698_ (.B(net756),
    .C(net593),
    .A(net723),
    .Y(_2191_));
 sg13g2_a21oi_1 _2699_ (.A1(_2190_),
    .A2(_2191_),
    .Y(_0044_),
    .B1(net648));
 sg13g2_nand2_1 _2700_ (.Y(_2192_),
    .A(net351),
    .B(net581));
 sg13g2_nand3_1 _2701_ (.B(net754),
    .C(net592),
    .A(net349),
    .Y(_2193_));
 sg13g2_a21oi_1 _2702_ (.A1(_2192_),
    .A2(_2193_),
    .Y(_0046_),
    .B1(net646));
 sg13g2_nand2_1 _2703_ (.Y(_2194_),
    .A(net726),
    .B(net582));
 sg13g2_nand3_1 _2704_ (.B(net754),
    .C(net592),
    .A(net722),
    .Y(_2195_));
 sg13g2_a21oi_1 _2705_ (.A1(_2194_),
    .A2(_2195_),
    .Y(_0047_),
    .B1(net646));
 sg13g2_nand2_1 _2706_ (.Y(_2196_),
    .A(net355),
    .B(net582));
 sg13g2_nand3_1 _2707_ (.B(net754),
    .C(net592),
    .A(net283),
    .Y(_2197_));
 sg13g2_a21oi_1 _2708_ (.A1(_2196_),
    .A2(_2197_),
    .Y(_0048_),
    .B1(net646));
 sg13g2_a22oi_1 _2709_ (.Y(_2198_),
    .B1(net583),
    .B2(net123),
    .A2(net591),
    .A1(_2063_));
 sg13g2_nor2_1 _2710_ (.A(net648),
    .B(_2198_),
    .Y(_0049_));
 sg13g2_nor2_1 _2711_ (.A(net1),
    .B(net581),
    .Y(_2199_));
 sg13g2_nor2_1 _2712_ (.A(net348),
    .B(_2150_),
    .Y(_2200_));
 sg13g2_nor3_1 _2713_ (.A(net645),
    .B(_2199_),
    .C(_2200_),
    .Y(_0050_));
 sg13g2_nor2_1 _2714_ (.A(net2),
    .B(net581),
    .Y(_2201_));
 sg13g2_nor2_1 _2715_ (.A(net724),
    .B(_2150_),
    .Y(_2202_));
 sg13g2_nor3_1 _2716_ (.A(net645),
    .B(_2201_),
    .C(_2202_),
    .Y(_0051_));
 sg13g2_nor2_1 _2717_ (.A(net3),
    .B(net581),
    .Y(_2203_));
 sg13g2_nor2_1 _2718_ (.A(net333),
    .B(_2150_),
    .Y(_2204_));
 sg13g2_nor3_1 _2719_ (.A(net645),
    .B(_2203_),
    .C(_2204_),
    .Y(_0052_));
 sg13g2_nor2_1 _2720_ (.A(net4),
    .B(net581),
    .Y(_2205_));
 sg13g2_nor2_1 _2721_ (.A(net723),
    .B(_2150_),
    .Y(_2206_));
 sg13g2_nor3_1 _2722_ (.A(net645),
    .B(_2205_),
    .C(_2206_),
    .Y(_0053_));
 sg13g2_nor2_1 _2723_ (.A(net5),
    .B(net581),
    .Y(_2207_));
 sg13g2_nor2_1 _2724_ (.A(net349),
    .B(_2150_),
    .Y(_2208_));
 sg13g2_nor3_1 _2725_ (.A(net645),
    .B(_2207_),
    .C(_2208_),
    .Y(_0054_));
 sg13g2_nor2_1 _2726_ (.A(net6),
    .B(net581),
    .Y(_2209_));
 sg13g2_nor2_1 _2727_ (.A(net120),
    .B(_2150_),
    .Y(_2210_));
 sg13g2_nor3_1 _2728_ (.A(net645),
    .B(_2209_),
    .C(_2210_),
    .Y(_0055_));
 sg13g2_nor2_1 _2729_ (.A(net7),
    .B(net581),
    .Y(_2211_));
 sg13g2_nor2_1 _2730_ (.A(net283),
    .B(_2150_),
    .Y(_2212_));
 sg13g2_nor3_1 _2731_ (.A(net645),
    .B(_2211_),
    .C(_2212_),
    .Y(_0057_));
 sg13g2_nor2_1 _2732_ (.A(net8),
    .B(net582),
    .Y(_2213_));
 sg13g2_nor2_1 _2733_ (.A(net37),
    .B(_2150_),
    .Y(_2214_));
 sg13g2_nor3_1 _2734_ (.A(net646),
    .B(_2213_),
    .C(_2214_),
    .Y(_0058_));
 sg13g2_nand2_1 _2735_ (.Y(_2215_),
    .A(\mul_accum[30] ),
    .B(\mul_accum[61] ));
 sg13g2_nor2_1 _2736_ (.A(\mul_accum[30] ),
    .B(\mul_accum[61] ),
    .Y(_2216_));
 sg13g2_xor2_1 _2737_ (.B(\mul_accum[61] ),
    .A(\mul_accum[30] ),
    .X(_2217_));
 sg13g2_or2_1 _2738_ (.X(_2218_),
    .B(\mul_accum[60] ),
    .A(\mul_accum[29] ));
 sg13g2_and2_1 _2739_ (.A(\mul_accum[29] ),
    .B(\mul_accum[60] ),
    .X(_2219_));
 sg13g2_and2_1 _2740_ (.A(\mul_accum[28] ),
    .B(\mul_accum[59] ),
    .X(_2220_));
 sg13g2_xor2_1 _2741_ (.B(\mul_accum[58] ),
    .A(\mul_accum[27] ),
    .X(_2221_));
 sg13g2_and2_1 _2742_ (.A(\mul_accum[26] ),
    .B(\mul_accum[57] ),
    .X(_2222_));
 sg13g2_xnor2_1 _2743_ (.Y(_2223_),
    .A(\mul_accum[26] ),
    .B(\mul_accum[57] ));
 sg13g2_inv_1 _2744_ (.Y(_2224_),
    .A(_2223_));
 sg13g2_nand2_1 _2745_ (.Y(_2225_),
    .A(_2221_),
    .B(_2224_));
 sg13g2_nor2_1 _2746_ (.A(\mul_accum[25] ),
    .B(\mul_accum[56] ),
    .Y(_2226_));
 sg13g2_a22oi_1 _2747_ (.Y(_2227_),
    .B1(\mul_accum[56] ),
    .B2(\mul_accum[25] ),
    .A2(\mul_accum[55] ),
    .A1(\mul_accum[24] ));
 sg13g2_and2_1 _2748_ (.A(\mul_accum[22] ),
    .B(\mul_accum[53] ),
    .X(_2228_));
 sg13g2_xor2_1 _2749_ (.B(\mul_accum[53] ),
    .A(\mul_accum[22] ),
    .X(_2229_));
 sg13g2_inv_1 _2750_ (.Y(_2230_),
    .A(_2229_));
 sg13g2_xnor2_1 _2751_ (.Y(_2231_),
    .A(\mul_accum[23] ),
    .B(\mul_accum[54] ));
 sg13g2_inv_1 _2752_ (.Y(_2232_),
    .A(_2231_));
 sg13g2_nor2_1 _2753_ (.A(\mul_accum[21] ),
    .B(\mul_accum[52] ),
    .Y(_2233_));
 sg13g2_nand2_1 _2754_ (.Y(_2234_),
    .A(\mul_accum[20] ),
    .B(\mul_accum[51] ));
 sg13g2_a22oi_1 _2755_ (.Y(_2235_),
    .B1(\mul_accum[52] ),
    .B2(\mul_accum[21] ),
    .A2(\mul_accum[51] ),
    .A1(\mul_accum[20] ));
 sg13g2_nor4_1 _2756_ (.A(_2230_),
    .B(_2231_),
    .C(_2233_),
    .D(_2235_),
    .Y(_2236_));
 sg13g2_a21oi_1 _2757_ (.A1(\mul_accum[23] ),
    .A2(\mul_accum[54] ),
    .Y(_2237_),
    .B1(_2228_));
 sg13g2_a21oi_1 _2758_ (.A1(_1943_),
    .A2(_1959_),
    .Y(_2238_),
    .B1(_2237_));
 sg13g2_nor2_1 _2759_ (.A(_2236_),
    .B(_2238_),
    .Y(_2239_));
 sg13g2_xor2_1 _2760_ (.B(\mul_accum[51] ),
    .A(\mul_accum[20] ),
    .X(_2240_));
 sg13g2_xnor2_1 _2761_ (.Y(_2241_),
    .A(\mul_accum[21] ),
    .B(\mul_accum[52] ));
 sg13g2_inv_1 _2762_ (.Y(_2242_),
    .A(_2241_));
 sg13g2_nand4_1 _2763_ (.B(_2232_),
    .C(_2240_),
    .A(_2229_),
    .Y(_2243_),
    .D(_2242_));
 sg13g2_and2_1 _2764_ (.A(\mul_accum[18] ),
    .B(\mul_accum[49] ),
    .X(_2244_));
 sg13g2_or2_1 _2765_ (.X(_2245_),
    .B(\mul_accum[49] ),
    .A(\mul_accum[18] ));
 sg13g2_xnor2_1 _2766_ (.Y(_2246_),
    .A(\mul_accum[18] ),
    .B(\mul_accum[49] ));
 sg13g2_nand2_1 _2767_ (.Y(_2247_),
    .A(\mul_accum[19] ),
    .B(\mul_accum[50] ));
 sg13g2_xnor2_1 _2768_ (.Y(_2248_),
    .A(\mul_accum[19] ),
    .B(\mul_accum[50] ));
 sg13g2_nor2_1 _2769_ (.A(_2246_),
    .B(_2248_),
    .Y(_2249_));
 sg13g2_nand2_1 _2770_ (.Y(_2250_),
    .A(\mul_accum[17] ),
    .B(\mul_accum[48] ));
 sg13g2_and2_1 _2771_ (.A(\mul_accum[16] ),
    .B(\mul_accum[47] ),
    .X(_2251_));
 sg13g2_nand2_1 _2772_ (.Y(_2252_),
    .A(\mul_accum[16] ),
    .B(\mul_accum[47] ));
 sg13g2_nor2_1 _2773_ (.A(\mul_accum[17] ),
    .B(\mul_accum[48] ),
    .Y(_2253_));
 sg13g2_or2_1 _2774_ (.X(_2254_),
    .B(\mul_accum[48] ),
    .A(\mul_accum[17] ));
 sg13g2_o21ai_1 _2775_ (.B1(_2250_),
    .Y(_2255_),
    .A1(_2252_),
    .A2(_2253_));
 sg13g2_nand2_1 _2776_ (.Y(_2256_),
    .A(_2249_),
    .B(_2255_));
 sg13g2_o21ai_1 _2777_ (.B1(_2244_),
    .Y(_2257_),
    .A1(\mul_accum[19] ),
    .A2(\mul_accum[50] ));
 sg13g2_nand3_1 _2778_ (.B(_2256_),
    .C(_2257_),
    .A(_2247_),
    .Y(_2258_));
 sg13g2_inv_1 _2779_ (.Y(_2259_),
    .A(_2258_));
 sg13g2_nand2_1 _2780_ (.Y(_2260_),
    .A(\mul_accum[15] ),
    .B(\mul_accum[46] ));
 sg13g2_nor2_1 _2781_ (.A(\mul_accum[15] ),
    .B(\mul_accum[46] ),
    .Y(_2261_));
 sg13g2_xor2_1 _2782_ (.B(\mul_accum[46] ),
    .A(\mul_accum[15] ),
    .X(_2262_));
 sg13g2_nand2_1 _2783_ (.Y(_2263_),
    .A(\mul_accum[14] ),
    .B(\mul_accum[45] ));
 sg13g2_inv_1 _2784_ (.Y(_2264_),
    .A(_2263_));
 sg13g2_xor2_1 _2785_ (.B(\mul_accum[45] ),
    .A(\mul_accum[14] ),
    .X(_2265_));
 sg13g2_and2_1 _2786_ (.A(_2262_),
    .B(_2265_),
    .X(_2266_));
 sg13g2_or2_1 _2787_ (.X(_2267_),
    .B(\mul_accum[44] ),
    .A(\mul_accum[13] ));
 sg13g2_nand2_1 _2788_ (.Y(_2268_),
    .A(\mul_accum[12] ),
    .B(\mul_accum[43] ));
 sg13g2_a22oi_1 _2789_ (.Y(_2269_),
    .B1(\mul_accum[44] ),
    .B2(\mul_accum[13] ),
    .A2(\mul_accum[43] ),
    .A1(\mul_accum[12] ));
 sg13g2_xnor2_1 _2790_ (.Y(_2270_),
    .A(\mul_accum[13] ),
    .B(\mul_accum[44] ));
 sg13g2_xnor2_1 _2791_ (.Y(_2271_),
    .A(\mul_accum[12] ),
    .B(\mul_accum[43] ));
 sg13g2_nor2_1 _2792_ (.A(_2270_),
    .B(_2271_),
    .Y(_2272_));
 sg13g2_or2_1 _2793_ (.X(_2273_),
    .B(\mul_accum[42] ),
    .A(\mul_accum[11] ));
 sg13g2_a22oi_1 _2794_ (.Y(_2274_),
    .B1(\mul_accum[42] ),
    .B2(\mul_accum[11] ),
    .A2(\mul_accum[41] ),
    .A1(\mul_accum[10] ));
 sg13g2_inv_1 _2795_ (.Y(_2275_),
    .A(_2274_));
 sg13g2_nand2_1 _2796_ (.Y(_2276_),
    .A(_2273_),
    .B(_2275_));
 sg13g2_xnor2_1 _2797_ (.Y(_2277_),
    .A(\mul_accum[10] ),
    .B(\mul_accum[41] ));
 sg13g2_xor2_1 _2798_ (.B(\mul_accum[42] ),
    .A(\mul_accum[11] ),
    .X(_2278_));
 sg13g2_nand2b_1 _2799_ (.Y(_2279_),
    .B(_2278_),
    .A_N(_2277_));
 sg13g2_nand2_1 _2800_ (.Y(_2280_),
    .A(\mul_accum[8] ),
    .B(\mul_accum[39] ));
 sg13g2_a22oi_1 _2801_ (.Y(_2281_),
    .B1(\mul_accum[40] ),
    .B2(\mul_accum[9] ),
    .A2(\mul_accum[39] ),
    .A1(\mul_accum[8] ));
 sg13g2_nor2_1 _2802_ (.A(\mul_accum[9] ),
    .B(\mul_accum[40] ),
    .Y(_2282_));
 sg13g2_or3_1 _2803_ (.A(_2279_),
    .B(_2281_),
    .C(_2282_),
    .X(_2283_));
 sg13g2_nand2_1 _2804_ (.Y(_2284_),
    .A(_2266_),
    .B(_2267_));
 sg13g2_nor2_1 _2805_ (.A(_2269_),
    .B(_2284_),
    .Y(_2285_));
 sg13g2_nand2_1 _2806_ (.Y(_2286_),
    .A(_2266_),
    .B(_2272_));
 sg13g2_a21oi_1 _2807_ (.A1(_2276_),
    .A2(_2283_),
    .Y(_2287_),
    .B1(_2286_));
 sg13g2_o21ai_1 _2808_ (.B1(_2260_),
    .Y(_2288_),
    .A1(_2261_),
    .A2(_2263_));
 sg13g2_nor3_2 _2809_ (.A(_2285_),
    .B(_2287_),
    .C(_2288_),
    .Y(_2289_));
 sg13g2_xnor2_1 _2810_ (.Y(_2290_),
    .A(\mul_accum[6] ),
    .B(\mul_accum[37] ));
 sg13g2_nor2_1 _2811_ (.A(\mul_accum[5] ),
    .B(\mul_accum[36] ),
    .Y(_2291_));
 sg13g2_nand2_1 _2812_ (.Y(_2292_),
    .A(\mul_accum[5] ),
    .B(\mul_accum[36] ));
 sg13g2_or2_1 _2813_ (.X(_2293_),
    .B(\mul_accum[34] ),
    .A(\mul_accum[3] ));
 sg13g2_nand2_1 _2814_ (.Y(_2294_),
    .A(\mul_accum[1] ),
    .B(\mul_accum[32] ));
 sg13g2_nand2_1 _2815_ (.Y(_2295_),
    .A(\mul_accum[0] ),
    .B(\mul_accum[31] ));
 sg13g2_nor2_1 _2816_ (.A(\mul_accum[1] ),
    .B(\mul_accum[32] ),
    .Y(_2296_));
 sg13g2_xor2_1 _2817_ (.B(\mul_accum[32] ),
    .A(\mul_accum[1] ),
    .X(_2297_));
 sg13g2_o21ai_1 _2818_ (.B1(_2294_),
    .Y(_2298_),
    .A1(_2295_),
    .A2(_2296_));
 sg13g2_xnor2_1 _2819_ (.Y(_2299_),
    .A(\mul_accum[2] ),
    .B(\mul_accum[33] ));
 sg13g2_nor2b_1 _2820_ (.A(_2299_),
    .B_N(_2298_),
    .Y(_2300_));
 sg13g2_a21oi_1 _2821_ (.A1(\mul_accum[2] ),
    .A2(\mul_accum[33] ),
    .Y(_2301_),
    .B1(_2300_));
 sg13g2_and3_1 _2822_ (.X(_2302_),
    .A(\mul_accum[2] ),
    .B(\mul_accum[33] ),
    .C(_2293_));
 sg13g2_xnor2_1 _2823_ (.Y(_2303_),
    .A(\mul_accum[3] ),
    .B(\mul_accum[34] ));
 sg13g2_nor2_1 _2824_ (.A(_2299_),
    .B(_2303_),
    .Y(_2304_));
 sg13g2_a221oi_1 _2825_ (.B2(_2304_),
    .C1(_2302_),
    .B1(_2298_),
    .A1(\mul_accum[3] ),
    .Y(_2305_),
    .A2(\mul_accum[34] ));
 sg13g2_xnor2_1 _2826_ (.Y(_2306_),
    .A(\mul_accum[4] ),
    .B(\mul_accum[35] ));
 sg13g2_nor2_1 _2827_ (.A(_2305_),
    .B(_2306_),
    .Y(_2307_));
 sg13g2_a21oi_1 _2828_ (.A1(\mul_accum[4] ),
    .A2(\mul_accum[35] ),
    .Y(_2308_),
    .B1(_2307_));
 sg13g2_a22oi_1 _2829_ (.Y(_2309_),
    .B1(\mul_accum[36] ),
    .B2(\mul_accum[5] ),
    .A2(\mul_accum[35] ),
    .A1(\mul_accum[4] ));
 sg13g2_a21oi_1 _2830_ (.A1(_2292_),
    .A2(_2308_),
    .Y(_2310_),
    .B1(_2291_));
 sg13g2_nor2b_1 _2831_ (.A(_2290_),
    .B_N(_2310_),
    .Y(_2311_));
 sg13g2_a21o_1 _2832_ (.A2(\mul_accum[37] ),
    .A1(\mul_accum[6] ),
    .B1(_2311_),
    .X(_2312_));
 sg13g2_a22oi_1 _2833_ (.Y(_2313_),
    .B1(\mul_accum[38] ),
    .B2(\mul_accum[7] ),
    .A2(\mul_accum[37] ),
    .A1(\mul_accum[6] ));
 sg13g2_a21oi_1 _2834_ (.A1(_1941_),
    .A2(_1949_),
    .Y(_2314_),
    .B1(_2313_));
 sg13g2_xnor2_1 _2835_ (.Y(_2315_),
    .A(\mul_accum[7] ),
    .B(\mul_accum[38] ));
 sg13g2_nor2_1 _2836_ (.A(_2290_),
    .B(_2315_),
    .Y(_2316_));
 sg13g2_or4_1 _2837_ (.A(_2290_),
    .B(_2291_),
    .C(_2309_),
    .D(_2315_),
    .X(_2317_));
 sg13g2_nor2b_1 _2838_ (.A(_2291_),
    .B_N(_2292_),
    .Y(_2318_));
 sg13g2_nand3b_1 _2839_ (.B(_2316_),
    .C(_2318_),
    .Y(_2319_),
    .A_N(_2306_));
 sg13g2_o21ai_1 _2840_ (.B1(_2317_),
    .Y(_2320_),
    .A1(_2305_),
    .A2(_2319_));
 sg13g2_nor2_1 _2841_ (.A(_2314_),
    .B(_2320_),
    .Y(_2321_));
 sg13g2_xor2_1 _2842_ (.B(\mul_accum[39] ),
    .A(\mul_accum[8] ),
    .X(_2322_));
 sg13g2_xor2_1 _2843_ (.B(\mul_accum[40] ),
    .A(\mul_accum[9] ),
    .X(_2323_));
 sg13g2_nand2_1 _2844_ (.Y(_2324_),
    .A(_2322_),
    .B(_2323_));
 sg13g2_nor3_1 _2845_ (.A(_2279_),
    .B(_2286_),
    .C(_2324_),
    .Y(_2325_));
 sg13g2_o21ai_1 _2846_ (.B1(_2325_),
    .Y(_2326_),
    .A1(_2314_),
    .A2(_2320_));
 sg13g2_nand2_1 _2847_ (.Y(_2327_),
    .A(_2289_),
    .B(_2326_));
 sg13g2_xor2_1 _2848_ (.B(\mul_accum[47] ),
    .A(\mul_accum[16] ),
    .X(_2328_));
 sg13g2_nand2_1 _2849_ (.Y(_2329_),
    .A(_2250_),
    .B(_2254_));
 sg13g2_nand4_1 _2850_ (.B(_2250_),
    .C(_2254_),
    .A(_2249_),
    .Y(_2330_),
    .D(_2328_));
 sg13g2_a21oi_1 _2851_ (.A1(_2289_),
    .A2(_2326_),
    .Y(_2331_),
    .B1(_2330_));
 sg13g2_o21ai_1 _2852_ (.B1(_2239_),
    .Y(_2332_),
    .A1(_2243_),
    .A2(_2259_));
 sg13g2_or2_1 _2853_ (.X(_2333_),
    .B(_2330_),
    .A(_2243_));
 sg13g2_a21oi_1 _2854_ (.A1(_2289_),
    .A2(_2326_),
    .Y(_2334_),
    .B1(_2333_));
 sg13g2_xor2_1 _2855_ (.B(\mul_accum[55] ),
    .A(\mul_accum[24] ),
    .X(_2335_));
 sg13g2_inv_1 _2856_ (.Y(_2336_),
    .A(_2335_));
 sg13g2_o21ai_1 _2857_ (.B1(_2335_),
    .Y(_2337_),
    .A1(_2332_),
    .A2(_2334_));
 sg13g2_a21oi_1 _2858_ (.A1(_2227_),
    .A2(_2337_),
    .Y(_2338_),
    .B1(_2226_));
 sg13g2_or3_1 _2859_ (.A(_2225_),
    .B(_2226_),
    .C(_2227_),
    .X(_2339_));
 sg13g2_xnor2_1 _2860_ (.Y(_2340_),
    .A(\mul_accum[25] ),
    .B(\mul_accum[56] ));
 sg13g2_nor3_1 _2861_ (.A(_2225_),
    .B(_2336_),
    .C(_2340_),
    .Y(_2341_));
 sg13g2_o21ai_1 _2862_ (.B1(_2341_),
    .Y(_2342_),
    .A1(_2332_),
    .A2(_2334_));
 sg13g2_a21oi_1 _2863_ (.A1(\mul_accum[27] ),
    .A2(\mul_accum[58] ),
    .Y(_2343_),
    .B1(_2222_));
 sg13g2_inv_1 _2864_ (.Y(_2344_),
    .A(_2343_));
 sg13g2_o21ai_1 _2865_ (.B1(_2344_),
    .Y(_2345_),
    .A1(\mul_accum[27] ),
    .A2(\mul_accum[58] ));
 sg13g2_nand3_1 _2866_ (.B(_2342_),
    .C(_2345_),
    .A(_2339_),
    .Y(_2346_));
 sg13g2_xor2_1 _2867_ (.B(\mul_accum[59] ),
    .A(\mul_accum[28] ),
    .X(_2347_));
 sg13g2_a21oi_1 _2868_ (.A1(_2346_),
    .A2(_2347_),
    .Y(_2348_),
    .B1(_2220_));
 sg13g2_xor2_1 _2869_ (.B(\mul_accum[60] ),
    .A(\mul_accum[29] ),
    .X(_2349_));
 sg13g2_and2_1 _2870_ (.A(_2347_),
    .B(_2349_),
    .X(_2350_));
 sg13g2_a221oi_1 _2871_ (.B2(_2350_),
    .C1(_2219_),
    .B1(_2346_),
    .A1(_2218_),
    .Y(_2351_),
    .A2(_2220_));
 sg13g2_xnor2_1 _2872_ (.Y(_2352_),
    .A(_2217_),
    .B(_2351_));
 sg13g2_xor2_1 _2873_ (.B(_2349_),
    .A(_2348_),
    .X(_2353_));
 sg13g2_xnor2_1 _2874_ (.Y(_2354_),
    .A(_2346_),
    .B(_2347_));
 sg13g2_a21oi_1 _2875_ (.A1(_2224_),
    .A2(_2338_),
    .Y(_2355_),
    .B1(_2222_));
 sg13g2_xor2_1 _2876_ (.B(_2355_),
    .A(_2221_),
    .X(_2356_));
 sg13g2_xnor2_1 _2877_ (.Y(_2357_),
    .A(_2221_),
    .B(_2355_));
 sg13g2_xnor2_1 _2878_ (.Y(_2358_),
    .A(_2223_),
    .B(_2338_));
 sg13g2_or3_1 _2879_ (.A(_2332_),
    .B(_2334_),
    .C(_2335_),
    .X(_2359_));
 sg13g2_and2_1 _2880_ (.A(_2337_),
    .B(_2359_),
    .X(_2360_));
 sg13g2_o21ai_1 _2881_ (.B1(_2337_),
    .Y(_2361_),
    .A1(_1944_),
    .A2(_1960_));
 sg13g2_xnor2_1 _2882_ (.Y(_2362_),
    .A(_2340_),
    .B(_2361_));
 sg13g2_nand2_1 _2883_ (.Y(_2363_),
    .A(_2360_),
    .B(_2362_));
 sg13g2_o21ai_1 _2884_ (.B1(_2240_),
    .Y(_2364_),
    .A1(_2258_),
    .A2(_2331_));
 sg13g2_a21oi_1 _2885_ (.A1(_2235_),
    .A2(_2364_),
    .Y(_2365_),
    .B1(_2233_));
 sg13g2_xnor2_1 _2886_ (.Y(_2366_),
    .A(_2229_),
    .B(_2365_));
 sg13g2_inv_1 _2887_ (.Y(_0229_),
    .A(_2366_));
 sg13g2_a21oi_1 _2888_ (.A1(_2229_),
    .A2(_2365_),
    .Y(_0230_),
    .B1(_2228_));
 sg13g2_xnor2_1 _2889_ (.Y(_0231_),
    .A(_2231_),
    .B(_0230_));
 sg13g2_nand2b_1 _2890_ (.Y(_0232_),
    .B(_0229_),
    .A_N(_0231_));
 sg13g2_or3_1 _2891_ (.A(_2240_),
    .B(_2258_),
    .C(_2331_),
    .X(_0233_));
 sg13g2_nand2_2 _2892_ (.Y(_0234_),
    .A(_2364_),
    .B(_0233_));
 sg13g2_nand2_1 _2893_ (.Y(_0235_),
    .A(_2234_),
    .B(_2364_));
 sg13g2_xnor2_1 _2894_ (.Y(_0236_),
    .A(_2241_),
    .B(_0235_));
 sg13g2_nor2b_2 _2895_ (.A(_0234_),
    .B_N(_0236_),
    .Y(_0237_));
 sg13g2_inv_2 _2896_ (.Y(_0238_),
    .A(_0237_));
 sg13g2_xor2_1 _2897_ (.B(_2315_),
    .A(_2312_),
    .X(_0239_));
 sg13g2_xor2_1 _2898_ (.B(_2303_),
    .A(_2301_),
    .X(_0240_));
 sg13g2_o21ai_1 _2899_ (.B1(_2215_),
    .Y(_0241_),
    .A1(_2216_),
    .A2(_2351_));
 sg13g2_xor2_1 _2900_ (.B(\mul_accum[31] ),
    .A(\mul_accum[0] ),
    .X(_0242_));
 sg13g2_xnor2_1 _2901_ (.Y(_0243_),
    .A(_2295_),
    .B(_2297_));
 sg13g2_nand3_1 _2902_ (.B(_0242_),
    .C(_0243_),
    .A(_0241_),
    .Y(_0244_));
 sg13g2_xor2_1 _2903_ (.B(_2299_),
    .A(_2298_),
    .X(_0245_));
 sg13g2_inv_1 _2904_ (.Y(_0246_),
    .A(_0245_));
 sg13g2_nand4_1 _2905_ (.B(_0242_),
    .C(_0243_),
    .A(_0241_),
    .Y(_0247_),
    .D(_0246_));
 sg13g2_and2_1 _2906_ (.A(_0240_),
    .B(_0246_),
    .X(_0248_));
 sg13g2_nand4_1 _2907_ (.B(_0242_),
    .C(_0243_),
    .A(_0241_),
    .Y(_0249_),
    .D(_0248_));
 sg13g2_xnor2_1 _2908_ (.Y(_0250_),
    .A(_2308_),
    .B(_2318_));
 sg13g2_xor2_1 _2909_ (.B(_2310_),
    .A(_2290_),
    .X(_0251_));
 sg13g2_xnor2_1 _2910_ (.Y(_0252_),
    .A(_2305_),
    .B(_2306_));
 sg13g2_nor2_1 _2911_ (.A(_0251_),
    .B(_0252_),
    .Y(_0253_));
 sg13g2_nand2_1 _2912_ (.Y(_0254_),
    .A(_0250_),
    .B(_0253_));
 sg13g2_nor2_1 _2913_ (.A(net562),
    .B(_0254_),
    .Y(_0255_));
 sg13g2_or2_1 _2914_ (.X(_0256_),
    .B(_0254_),
    .A(_0239_));
 sg13g2_inv_1 _2915_ (.Y(_0257_),
    .A(net564));
 sg13g2_nor2_1 _2916_ (.A(net562),
    .B(net564),
    .Y(_0258_));
 sg13g2_o21ai_1 _2917_ (.B1(_2322_),
    .Y(_0259_),
    .A1(_2314_),
    .A2(_2320_));
 sg13g2_a21oi_1 _2918_ (.A1(_2281_),
    .A2(_0259_),
    .Y(_0260_),
    .B1(_2282_));
 sg13g2_a221oi_1 _2919_ (.B2(_0259_),
    .C1(_2277_),
    .B1(_2281_),
    .A1(_1942_),
    .Y(_0261_),
    .A2(_1950_));
 sg13g2_o21ai_1 _2920_ (.B1(_2273_),
    .Y(_0262_),
    .A1(_2275_),
    .A2(_0261_));
 sg13g2_o21ai_1 _2921_ (.B1(_2269_),
    .Y(_0263_),
    .A1(_2271_),
    .A2(_0262_));
 sg13g2_and3_2 _2922_ (.X(_0264_),
    .A(_2265_),
    .B(_2267_),
    .C(_0263_));
 sg13g2_a21oi_1 _2923_ (.A1(_2267_),
    .A2(_0263_),
    .Y(_0265_),
    .B1(_2265_));
 sg13g2_nor2_1 _2924_ (.A(_0264_),
    .B(_0265_),
    .Y(_0266_));
 sg13g2_xor2_1 _2925_ (.B(_0262_),
    .A(_2271_),
    .X(_0267_));
 sg13g2_xor2_1 _2926_ (.B(_2322_),
    .A(_2321_),
    .X(_0268_));
 sg13g2_nand2_1 _2927_ (.Y(_0269_),
    .A(_2280_),
    .B(_0259_));
 sg13g2_xnor2_1 _2928_ (.Y(_0270_),
    .A(_2323_),
    .B(_0269_));
 sg13g2_nor2_1 _2929_ (.A(_0268_),
    .B(_0270_),
    .Y(_0271_));
 sg13g2_xnor2_1 _2930_ (.Y(_0272_),
    .A(_2277_),
    .B(_0260_));
 sg13g2_nand2_2 _2931_ (.Y(_0273_),
    .A(_0271_),
    .B(_0272_));
 sg13g2_a21oi_1 _2932_ (.A1(\mul_accum[10] ),
    .A2(\mul_accum[41] ),
    .Y(_0274_),
    .B1(_0261_));
 sg13g2_xnor2_1 _2933_ (.Y(_0275_),
    .A(_2278_),
    .B(_0274_));
 sg13g2_nor2b_1 _2934_ (.A(_0273_),
    .B_N(_0275_),
    .Y(_0276_));
 sg13g2_nand2_1 _2935_ (.Y(_0277_),
    .A(_0267_),
    .B(_0275_));
 sg13g2_nor4_1 _2936_ (.A(_0264_),
    .B(_0265_),
    .C(_0273_),
    .D(_0277_),
    .Y(_0278_));
 sg13g2_or3_1 _2937_ (.A(_2262_),
    .B(_2264_),
    .C(_0264_),
    .X(_0279_));
 sg13g2_o21ai_1 _2938_ (.B1(_2262_),
    .Y(_0280_),
    .A1(_2264_),
    .A2(_0264_));
 sg13g2_nand2_1 _2939_ (.Y(_0281_),
    .A(_0279_),
    .B(_0280_));
 sg13g2_o21ai_1 _2940_ (.B1(_2268_),
    .Y(_0282_),
    .A1(_2271_),
    .A2(_0262_));
 sg13g2_xnor2_1 _2941_ (.Y(_0283_),
    .A(_2270_),
    .B(_0282_));
 sg13g2_nand3_1 _2942_ (.B(_0280_),
    .C(_0283_),
    .A(_0279_),
    .Y(_0284_));
 sg13g2_nand4_1 _2943_ (.B(_0279_),
    .C(_0280_),
    .A(_0278_),
    .Y(_0285_),
    .D(_0283_));
 sg13g2_nor3_1 _2944_ (.A(net563),
    .B(net564),
    .C(_0285_),
    .Y(_0286_));
 sg13g2_xnor2_1 _2945_ (.Y(_0287_),
    .A(_2327_),
    .B(_2328_));
 sg13g2_nor4_2 _2946_ (.A(net563),
    .B(net564),
    .C(_0285_),
    .Y(_0288_),
    .D(_0287_));
 sg13g2_a21oi_1 _2947_ (.A1(_2327_),
    .A2(_2328_),
    .Y(_0289_),
    .B1(_2251_));
 sg13g2_o21ai_1 _2948_ (.B1(_2250_),
    .Y(_0290_),
    .A1(_2253_),
    .A2(_0289_));
 sg13g2_a21oi_1 _2949_ (.A1(_2245_),
    .A2(_0290_),
    .Y(_0291_),
    .B1(_2244_));
 sg13g2_xor2_1 _2950_ (.B(_0291_),
    .A(_2248_),
    .X(_0292_));
 sg13g2_xor2_1 _2951_ (.B(_0290_),
    .A(_2246_),
    .X(_0293_));
 sg13g2_xnor2_1 _2952_ (.Y(_0294_),
    .A(_2329_),
    .B(_0289_));
 sg13g2_inv_1 _2953_ (.Y(_0295_),
    .A(_0294_));
 sg13g2_nor2_1 _2954_ (.A(_0293_),
    .B(_0294_),
    .Y(_0296_));
 sg13g2_nand3_1 _2955_ (.B(_0292_),
    .C(_0296_),
    .A(_0288_),
    .Y(_0297_));
 sg13g2_nor3_1 _2956_ (.A(_0232_),
    .B(_0238_),
    .C(_0297_),
    .Y(_0298_));
 sg13g2_nor2b_1 _2957_ (.A(_2363_),
    .B_N(_0298_),
    .Y(_0299_));
 sg13g2_nand3_1 _2958_ (.B(_2358_),
    .C(_0299_),
    .A(_2357_),
    .Y(_0300_));
 sg13g2_nor2_1 _2959_ (.A(_2354_),
    .B(_0300_),
    .Y(_0301_));
 sg13g2_nand3b_1 _2960_ (.B(_0292_),
    .C(_0296_),
    .Y(_0302_),
    .A_N(_0287_));
 sg13g2_nor4_2 _2961_ (.A(net563),
    .B(net564),
    .C(_0285_),
    .Y(_0303_),
    .D(_0302_));
 sg13g2_or4_1 _2962_ (.A(net563),
    .B(_0256_),
    .C(_0285_),
    .D(_0302_),
    .X(_0304_));
 sg13g2_nor3_1 _2963_ (.A(_0232_),
    .B(_0238_),
    .C(_0304_),
    .Y(_0305_));
 sg13g2_nor4_2 _2964_ (.A(_2363_),
    .B(_0232_),
    .C(_0238_),
    .Y(_0306_),
    .D(_0304_));
 sg13g2_nand3_1 _2965_ (.B(_2358_),
    .C(_0306_),
    .A(_2357_),
    .Y(_0307_));
 sg13g2_nor3_1 _2966_ (.A(_2353_),
    .B(_2354_),
    .C(_0307_),
    .Y(_0308_));
 sg13g2_or2_1 _2967_ (.X(_0309_),
    .B(_0308_),
    .A(_2352_));
 sg13g2_xnor2_1 _2968_ (.Y(_0310_),
    .A(_2354_),
    .B(_0307_));
 sg13g2_xor2_1 _2969_ (.B(_0306_),
    .A(_2358_),
    .X(_0311_));
 sg13g2_inv_1 _2970_ (.Y(_0312_),
    .A(_0311_));
 sg13g2_nor3_1 _2971_ (.A(_2366_),
    .B(_0238_),
    .C(_0297_),
    .Y(_0313_));
 sg13g2_nand3_1 _2972_ (.B(_0237_),
    .C(_0303_),
    .A(_0229_),
    .Y(_0314_));
 sg13g2_a21oi_2 _2973_ (.B1(_0305_),
    .Y(_0315_),
    .A2(_0314_),
    .A1(_0231_));
 sg13g2_inv_1 _2974_ (.Y(_0316_),
    .A(_0315_));
 sg13g2_nor3_1 _2975_ (.A(net562),
    .B(net564),
    .C(_0273_),
    .Y(_0317_));
 sg13g2_nor3_1 _2976_ (.A(net562),
    .B(net564),
    .C(_0268_),
    .Y(_0318_));
 sg13g2_a21oi_1 _2977_ (.A1(_0258_),
    .A2(_0271_),
    .Y(_0319_),
    .B1(_0272_));
 sg13g2_nor2_2 _2978_ (.A(_0317_),
    .B(_0319_),
    .Y(_0320_));
 sg13g2_xnor2_1 _2979_ (.Y(_0321_),
    .A(_0286_),
    .B(_0287_));
 sg13g2_nand3b_1 _2980_ (.B(_0257_),
    .C(_0276_),
    .Y(_0322_),
    .A_N(net562));
 sg13g2_nor4_2 _2981_ (.A(net562),
    .B(net564),
    .C(_0273_),
    .Y(_0323_),
    .D(_0277_));
 sg13g2_xnor2_1 _2982_ (.Y(_0324_),
    .A(_0267_),
    .B(_0322_));
 sg13g2_nor2_1 _2983_ (.A(net562),
    .B(_0252_),
    .Y(_0325_));
 sg13g2_nand2_1 _2984_ (.Y(_0326_),
    .A(_0250_),
    .B(_0325_));
 sg13g2_xor2_1 _2985_ (.B(_0325_),
    .A(_0250_),
    .X(_0327_));
 sg13g2_xnor2_1 _2986_ (.Y(_0328_),
    .A(_0239_),
    .B(_0255_));
 sg13g2_xnor2_1 _2987_ (.Y(_0329_),
    .A(_0240_),
    .B(_0247_));
 sg13g2_xnor2_1 _2988_ (.Y(_0330_),
    .A(_0244_),
    .B(_0246_));
 sg13g2_xor2_1 _2989_ (.B(_0242_),
    .A(_0241_),
    .X(_0331_));
 sg13g2_and4_1 _2990_ (.A(_0243_),
    .B(_0253_),
    .C(_0271_),
    .D(_0275_),
    .X(_0332_));
 sg13g2_and2_1 _2991_ (.A(_2360_),
    .B(_0332_),
    .X(_0333_));
 sg13g2_nor3_1 _2992_ (.A(_2366_),
    .B(_0293_),
    .C(_0294_),
    .Y(_0334_));
 sg13g2_nand4_1 _2993_ (.B(_0237_),
    .C(_0333_),
    .A(_2362_),
    .Y(_0335_),
    .D(_0334_));
 sg13g2_nor4_2 _2994_ (.A(_2353_),
    .B(_2356_),
    .C(_0284_),
    .Y(_0336_),
    .D(_0335_));
 sg13g2_and4_1 _2995_ (.A(_0329_),
    .B(_0330_),
    .C(_0331_),
    .D(_0336_),
    .X(_0337_));
 sg13g2_and4_1 _2996_ (.A(_0324_),
    .B(_0327_),
    .C(_0328_),
    .D(_0337_),
    .X(_0338_));
 sg13g2_a21oi_1 _2997_ (.A1(_0288_),
    .A2(_0296_),
    .Y(_0339_),
    .B1(_0292_));
 sg13g2_a21oi_1 _2998_ (.A1(_0283_),
    .A2(_0323_),
    .Y(_0340_),
    .B1(_0266_));
 sg13g2_and3_1 _2999_ (.X(_0341_),
    .A(_0266_),
    .B(_0283_),
    .C(_0323_));
 sg13g2_nand3_1 _3000_ (.B(_0283_),
    .C(_0323_),
    .A(_0266_),
    .Y(_0342_));
 sg13g2_nor2_1 _3001_ (.A(_0340_),
    .B(_0341_),
    .Y(_0343_));
 sg13g2_inv_1 _3002_ (.Y(_0344_),
    .A(_0343_));
 sg13g2_nor4_1 _3003_ (.A(_0303_),
    .B(_0339_),
    .C(_0340_),
    .D(_0341_),
    .Y(_0345_));
 sg13g2_nand4_1 _3004_ (.B(_0321_),
    .C(_0338_),
    .A(_0320_),
    .Y(_0346_),
    .D(_0345_));
 sg13g2_nor4_2 _3005_ (.A(_0310_),
    .B(_0312_),
    .C(_0316_),
    .Y(_0347_),
    .D(_0346_));
 sg13g2_inv_1 _3006_ (.Y(_0348_),
    .A(net560));
 sg13g2_nand2_1 _3007_ (.Y(_0349_),
    .A(_0234_),
    .B(_0304_));
 sg13g2_nor2_1 _3008_ (.A(_0234_),
    .B(_0297_),
    .Y(_0350_));
 sg13g2_a21o_1 _3009_ (.A2(_0306_),
    .A1(_2358_),
    .B1(_2357_),
    .X(_0351_));
 sg13g2_or2_1 _3010_ (.X(_0352_),
    .B(_0305_),
    .A(_2360_));
 sg13g2_nand2_1 _3011_ (.Y(_0353_),
    .A(_2360_),
    .B(_0298_));
 sg13g2_and2_1 _3012_ (.A(net561),
    .B(_0348_),
    .X(_0354_));
 sg13g2_nand2_1 _3013_ (.Y(_0355_),
    .A(\reg_a[30] ),
    .B(_0354_));
 sg13g2_and2_1 _3014_ (.A(net561),
    .B(net560),
    .X(_0356_));
 sg13g2_nand2_1 _3015_ (.Y(_0357_),
    .A(net561),
    .B(net560));
 sg13g2_a21o_1 _3016_ (.A2(_0242_),
    .A1(_0241_),
    .B1(_0243_),
    .X(_0358_));
 sg13g2_and2_1 _3017_ (.A(_0244_),
    .B(_0358_),
    .X(_0359_));
 sg13g2_nand2_1 _3018_ (.Y(_0360_),
    .A(net553),
    .B(_0359_));
 sg13g2_nand3_1 _3019_ (.B(net553),
    .C(_0359_),
    .A(net747),
    .Y(_0361_));
 sg13g2_nand2_1 _3020_ (.Y(_0362_),
    .A(_0331_),
    .B(net555));
 sg13g2_nand3_1 _3021_ (.B(_0331_),
    .C(net554),
    .A(\reg_a[0] ),
    .Y(_0363_));
 sg13g2_a21oi_1 _3022_ (.A1(net553),
    .A2(_0359_),
    .Y(_0364_),
    .B1(net747));
 sg13g2_xor2_1 _3023_ (.B(_0360_),
    .A(net747),
    .X(_0365_));
 sg13g2_o21ai_1 _3024_ (.B1(_0361_),
    .Y(_0366_),
    .A1(_0363_),
    .A2(_0364_));
 sg13g2_and2_1 _3025_ (.A(_0330_),
    .B(net553),
    .X(_0367_));
 sg13g2_nand2_1 _3026_ (.Y(_0368_),
    .A(net746),
    .B(_0367_));
 sg13g2_xnor2_1 _3027_ (.Y(_0369_),
    .A(net746),
    .B(_0367_));
 sg13g2_nand2b_1 _3028_ (.Y(_0370_),
    .B(_0366_),
    .A_N(_0369_));
 sg13g2_nand2_2 _3029_ (.Y(_0371_),
    .A(_0329_),
    .B(net553));
 sg13g2_nor2_1 _3030_ (.A(_1928_),
    .B(_0371_),
    .Y(_0372_));
 sg13g2_a21oi_1 _3031_ (.A1(net746),
    .A2(_0367_),
    .Y(_0373_),
    .B1(_0372_));
 sg13g2_a22oi_1 _3032_ (.Y(_0374_),
    .B1(_0373_),
    .B2(_0370_),
    .A2(_0371_),
    .A1(_1928_));
 sg13g2_nand2_1 _3033_ (.Y(_0375_),
    .A(_0328_),
    .B(net555));
 sg13g2_nand3_1 _3034_ (.B(_0328_),
    .C(net554),
    .A(net745),
    .Y(_0376_));
 sg13g2_a21o_1 _3035_ (.A2(net554),
    .A1(_0328_),
    .B1(net745),
    .X(_0377_));
 sg13g2_and2_1 _3036_ (.A(_0376_),
    .B(_0377_),
    .X(_0378_));
 sg13g2_a21oi_1 _3037_ (.A1(_0251_),
    .A2(_0326_),
    .Y(_0379_),
    .B1(_0255_));
 sg13g2_and2_1 _3038_ (.A(net553),
    .B(_0379_),
    .X(_0380_));
 sg13g2_nand2_1 _3039_ (.Y(_0381_),
    .A(net554),
    .B(_0379_));
 sg13g2_nand2_1 _3040_ (.Y(_0382_),
    .A(\reg_a[6] ),
    .B(_0380_));
 sg13g2_xnor2_1 _3041_ (.Y(_0383_),
    .A(_1934_),
    .B(_0380_));
 sg13g2_xnor2_1 _3042_ (.Y(_0384_),
    .A(\reg_a[6] ),
    .B(_0380_));
 sg13g2_nand2_1 _3043_ (.Y(_0385_),
    .A(net562),
    .B(_0252_));
 sg13g2_nand3b_1 _3044_ (.B(net553),
    .C(_0385_),
    .Y(_0386_),
    .A_N(_0325_));
 sg13g2_inv_1 _3045_ (.Y(_0387_),
    .A(_0386_));
 sg13g2_xnor2_1 _3046_ (.Y(_0388_),
    .A(\reg_a[4] ),
    .B(_0386_));
 sg13g2_nand3_1 _3047_ (.B(_0327_),
    .C(net553),
    .A(\reg_a[5] ),
    .Y(_0389_));
 sg13g2_a21o_1 _3048_ (.A2(net554),
    .A1(_0327_),
    .B1(\reg_a[5] ),
    .X(_0390_));
 sg13g2_and2_1 _3049_ (.A(_0389_),
    .B(_0390_),
    .X(_0391_));
 sg13g2_nand4_1 _3050_ (.B(_0383_),
    .C(_0388_),
    .A(_0378_),
    .Y(_0392_),
    .D(_0391_));
 sg13g2_a221oi_1 _3051_ (.B2(_0370_),
    .C1(_0392_),
    .B1(_0373_),
    .A1(_1928_),
    .Y(_0393_),
    .A2(_0371_));
 sg13g2_o21ai_1 _3052_ (.B1(_0389_),
    .Y(_0394_),
    .A1(_1932_),
    .A2(_0386_));
 sg13g2_and4_1 _3053_ (.A(_0378_),
    .B(_0383_),
    .C(_0390_),
    .D(_0394_),
    .X(_0395_));
 sg13g2_nand2_1 _3054_ (.Y(_0396_),
    .A(_0376_),
    .B(_0382_));
 sg13g2_a21o_1 _3055_ (.A2(_0396_),
    .A1(_0377_),
    .B1(_0395_),
    .X(_0397_));
 sg13g2_o21ai_1 _3056_ (.B1(_0322_),
    .Y(_0398_),
    .A1(_0275_),
    .A2(_0317_));
 sg13g2_a21o_2 _3057_ (.A2(net560),
    .A1(net561),
    .B1(_0398_),
    .X(_0399_));
 sg13g2_nor2_1 _3058_ (.A(_1931_),
    .B(_0399_),
    .Y(_0400_));
 sg13g2_nand2_1 _3059_ (.Y(_0401_),
    .A(_1931_),
    .B(_0399_));
 sg13g2_xnor2_1 _3060_ (.Y(_0402_),
    .A(_1931_),
    .B(_0399_));
 sg13g2_xnor2_1 _3061_ (.Y(_0403_),
    .A(_0270_),
    .B(_0318_));
 sg13g2_and2_1 _3062_ (.A(net556),
    .B(_0403_),
    .X(_0404_));
 sg13g2_a21oi_1 _3063_ (.A1(net556),
    .A2(_0403_),
    .Y(_0405_),
    .B1(\reg_a[9] ));
 sg13g2_and3_2 _3064_ (.X(_0406_),
    .A(net743),
    .B(_0320_),
    .C(net557));
 sg13g2_a21oi_1 _3065_ (.A1(_0320_),
    .A2(net557),
    .Y(_0407_),
    .B1(net743));
 sg13g2_nor2_1 _3066_ (.A(_0406_),
    .B(_0407_),
    .Y(_0408_));
 sg13g2_nor4_1 _3067_ (.A(_0402_),
    .B(_0405_),
    .C(_0406_),
    .D(_0407_),
    .Y(_0409_));
 sg13g2_nand3_1 _3068_ (.B(net556),
    .C(_0403_),
    .A(\reg_a[9] ),
    .Y(_0410_));
 sg13g2_nand2_1 _3069_ (.Y(_0411_),
    .A(_0409_),
    .B(_0410_));
 sg13g2_xnor2_1 _3070_ (.Y(_0412_),
    .A(_0258_),
    .B(_0268_));
 sg13g2_and2_1 _3071_ (.A(net556),
    .B(_0412_),
    .X(_0413_));
 sg13g2_nand3_1 _3072_ (.B(net556),
    .C(_0412_),
    .A(net744),
    .Y(_0414_));
 sg13g2_xnor2_1 _3073_ (.Y(_0415_),
    .A(net744),
    .B(_0413_));
 sg13g2_inv_1 _3074_ (.Y(_0416_),
    .A(_0415_));
 sg13g2_a21oi_1 _3075_ (.A1(_0281_),
    .A2(_0342_),
    .Y(_0417_),
    .B1(_0286_));
 sg13g2_a221oi_1 _3076_ (.B2(net561),
    .C1(_0286_),
    .B1(net560),
    .A1(_0281_),
    .Y(_0418_),
    .A2(_0342_));
 sg13g2_nand2_1 _3077_ (.Y(_0419_),
    .A(net557),
    .B(_0417_));
 sg13g2_nor2_1 _3078_ (.A(_1937_),
    .B(_0419_),
    .Y(_0420_));
 sg13g2_nand2_1 _3079_ (.Y(_0421_),
    .A(_1937_),
    .B(_0419_));
 sg13g2_xnor2_1 _3080_ (.Y(_0422_),
    .A(\reg_a[15] ),
    .B(_0418_));
 sg13g2_a21oi_2 _3081_ (.B1(_0344_),
    .Y(_0423_),
    .A2(net560),
    .A1(net561));
 sg13g2_and2_1 _3082_ (.A(\reg_a[14] ),
    .B(_0423_),
    .X(_0424_));
 sg13g2_xnor2_1 _3083_ (.Y(_0425_),
    .A(_1936_),
    .B(_0423_));
 sg13g2_nor2b_1 _3084_ (.A(_0422_),
    .B_N(_0425_),
    .Y(_0426_));
 sg13g2_and2_1 _3085_ (.A(_0324_),
    .B(net555),
    .X(_0427_));
 sg13g2_nand2_1 _3086_ (.Y(_0428_),
    .A(net742),
    .B(_0427_));
 sg13g2_xor2_1 _3087_ (.B(_0427_),
    .A(net742),
    .X(_0429_));
 sg13g2_xor2_1 _3088_ (.B(_0323_),
    .A(_0283_),
    .X(_0430_));
 sg13g2_a21oi_1 _3089_ (.A1(net557),
    .A2(_0430_),
    .Y(_0431_),
    .B1(net741));
 sg13g2_nand3_1 _3090_ (.B(net557),
    .C(_0430_),
    .A(net741),
    .Y(_0432_));
 sg13g2_nor2b_1 _3091_ (.A(_0431_),
    .B_N(_0432_),
    .Y(_0433_));
 sg13g2_nand3_1 _3092_ (.B(_0429_),
    .C(_0433_),
    .A(_0426_),
    .Y(_0434_));
 sg13g2_nor3_1 _3093_ (.A(_0411_),
    .B(_0415_),
    .C(_0434_),
    .Y(_0435_));
 sg13g2_o21ai_1 _3094_ (.B1(_0435_),
    .Y(_0436_),
    .A1(_0393_),
    .A2(_0397_));
 sg13g2_nand2_1 _3095_ (.Y(_0437_),
    .A(_0410_),
    .B(_0414_));
 sg13g2_inv_1 _3096_ (.Y(_0438_),
    .A(_0437_));
 sg13g2_or2_1 _3097_ (.X(_0439_),
    .B(_0406_),
    .A(_0400_));
 sg13g2_a22oi_1 _3098_ (.Y(_0440_),
    .B1(_0439_),
    .B2(_0401_),
    .A2(_0437_),
    .A1(_0409_));
 sg13g2_o21ai_1 _3099_ (.B1(_0432_),
    .Y(_0441_),
    .A1(_0428_),
    .A2(_0431_));
 sg13g2_a21oi_1 _3100_ (.A1(_0421_),
    .A2(_0424_),
    .Y(_0442_),
    .B1(_0420_));
 sg13g2_o21ai_1 _3101_ (.B1(_0442_),
    .Y(_0443_),
    .A1(_0434_),
    .A2(_0440_));
 sg13g2_a21oi_2 _3102_ (.B1(_0443_),
    .Y(_0444_),
    .A2(_0441_),
    .A1(_0426_));
 sg13g2_nand2_2 _3103_ (.Y(_0445_),
    .A(_0436_),
    .B(_0444_));
 sg13g2_nand3_1 _3104_ (.B(_0315_),
    .C(net559),
    .A(net736),
    .Y(_0446_));
 sg13g2_a21oi_1 _3105_ (.A1(_0315_),
    .A2(net558),
    .Y(_0447_),
    .B1(net736));
 sg13g2_a21o_1 _3106_ (.A2(net558),
    .A1(_0315_),
    .B1(net736),
    .X(_0448_));
 sg13g2_nand2_1 _3107_ (.Y(_0449_),
    .A(_0446_),
    .B(_0448_));
 sg13g2_a21oi_1 _3108_ (.A1(_0237_),
    .A2(_0303_),
    .Y(_0450_),
    .B1(_0229_));
 sg13g2_nor3_2 _3109_ (.A(_0313_),
    .B(_0356_),
    .C(_0450_),
    .Y(_0451_));
 sg13g2_nand2_1 _3110_ (.Y(_0452_),
    .A(net738),
    .B(_0451_));
 sg13g2_xnor2_1 _3111_ (.Y(_0453_),
    .A(net738),
    .B(_0451_));
 sg13g2_a21oi_1 _3112_ (.A1(_0309_),
    .A2(net560),
    .Y(_0454_),
    .B1(_0350_));
 sg13g2_xnor2_1 _3113_ (.Y(_0455_),
    .A(_0236_),
    .B(_0454_));
 sg13g2_nor2_1 _3114_ (.A(net739),
    .B(_0455_),
    .Y(_0456_));
 sg13g2_nand2_2 _3115_ (.Y(_0457_),
    .A(_0349_),
    .B(_0454_));
 sg13g2_nor2_1 _3116_ (.A(_1933_),
    .B(_0457_),
    .Y(_0458_));
 sg13g2_xnor2_1 _3117_ (.Y(_0459_),
    .A(_1933_),
    .B(_0457_));
 sg13g2_nand2_1 _3118_ (.Y(_0460_),
    .A(net739),
    .B(_0455_));
 sg13g2_or2_1 _3119_ (.X(_0461_),
    .B(_0453_),
    .A(_0449_));
 sg13g2_nand2b_1 _3120_ (.Y(_0462_),
    .B(_0460_),
    .A_N(_0456_));
 sg13g2_or3_1 _3121_ (.A(_0459_),
    .B(_0461_),
    .C(_0462_),
    .X(_0463_));
 sg13g2_or3_1 _3122_ (.A(_0303_),
    .B(_0339_),
    .C(_0356_),
    .X(_0464_));
 sg13g2_xnor2_1 _3123_ (.Y(_0465_),
    .A(\reg_a[19] ),
    .B(_0464_));
 sg13g2_nand2_1 _3124_ (.Y(_0466_),
    .A(_0288_),
    .B(_0295_));
 sg13g2_a22oi_1 _3125_ (.Y(_0467_),
    .B1(_0466_),
    .B2(_0293_),
    .A2(_0296_),
    .A1(_0288_));
 sg13g2_nand2_1 _3126_ (.Y(_0468_),
    .A(net558),
    .B(_0467_));
 sg13g2_nand3_1 _3127_ (.B(net558),
    .C(_0467_),
    .A(\reg_a[18] ),
    .Y(_0469_));
 sg13g2_a21oi_1 _3128_ (.A1(net558),
    .A2(_0467_),
    .Y(_0470_),
    .B1(\reg_a[18] ));
 sg13g2_xnor2_1 _3129_ (.Y(_0471_),
    .A(\reg_a[18] ),
    .B(_0468_));
 sg13g2_a21oi_1 _3130_ (.A1(net561),
    .A2(net560),
    .Y(_0472_),
    .B1(_0294_));
 sg13g2_mux2_1 _3131_ (.A0(_0472_),
    .A1(_0294_),
    .S(_0288_),
    .X(_0473_));
 sg13g2_or2_1 _3132_ (.X(_0474_),
    .B(_0473_),
    .A(\reg_a[17] ));
 sg13g2_and3_1 _3133_ (.X(_0475_),
    .A(_0465_),
    .B(_0471_),
    .C(_0474_));
 sg13g2_and2_1 _3134_ (.A(_0321_),
    .B(net558),
    .X(_0476_));
 sg13g2_nand2_1 _3135_ (.Y(_0477_),
    .A(net740),
    .B(_0476_));
 sg13g2_xnor2_1 _3136_ (.Y(_0478_),
    .A(net740),
    .B(_0476_));
 sg13g2_nand2_1 _3137_ (.Y(_0479_),
    .A(\reg_a[17] ),
    .B(_0473_));
 sg13g2_nand2_1 _3138_ (.Y(_0480_),
    .A(_0465_),
    .B(_0471_));
 sg13g2_nand2_1 _3139_ (.Y(_0481_),
    .A(_0474_),
    .B(_0479_));
 sg13g2_nor3_1 _3140_ (.A(_0478_),
    .B(_0480_),
    .C(_0481_),
    .Y(_0482_));
 sg13g2_nand2b_1 _3141_ (.Y(_0483_),
    .B(_0482_),
    .A_N(_0463_));
 sg13g2_a21oi_1 _3142_ (.A1(_0436_),
    .A2(_0444_),
    .Y(_0484_),
    .B1(_0483_));
 sg13g2_nand2_1 _3143_ (.Y(_0485_),
    .A(_0477_),
    .B(_0479_));
 sg13g2_a21o_1 _3144_ (.A2(_0464_),
    .A1(_1930_),
    .B1(_0469_),
    .X(_0486_));
 sg13g2_o21ai_1 _3145_ (.B1(_0486_),
    .Y(_0487_),
    .A1(_1930_),
    .A2(_0464_));
 sg13g2_a21o_1 _3146_ (.A2(_0485_),
    .A1(_0475_),
    .B1(_0487_),
    .X(_0488_));
 sg13g2_nor2b_1 _3147_ (.A(_0463_),
    .B_N(_0488_),
    .Y(_0489_));
 sg13g2_nor2b_1 _3148_ (.A(_0458_),
    .B_N(_0460_),
    .Y(_0490_));
 sg13g2_nor3_1 _3149_ (.A(_0456_),
    .B(_0461_),
    .C(_0490_),
    .Y(_0491_));
 sg13g2_o21ai_1 _3150_ (.B1(_0446_),
    .Y(_0492_),
    .A1(_0447_),
    .A2(_0452_));
 sg13g2_or3_1 _3151_ (.A(_0489_),
    .B(_0491_),
    .C(_0492_),
    .X(_0493_));
 sg13g2_nor2_1 _3152_ (.A(_0484_),
    .B(_0493_),
    .Y(_0494_));
 sg13g2_nand3_1 _3153_ (.B(_0351_),
    .C(net559),
    .A(_0307_),
    .Y(_0495_));
 sg13g2_nand2_1 _3154_ (.Y(_0496_),
    .A(_1929_),
    .B(_0495_));
 sg13g2_xnor2_1 _3155_ (.Y(_0497_),
    .A(_1929_),
    .B(_0495_));
 sg13g2_nor2_2 _3156_ (.A(_0312_),
    .B(_0356_),
    .Y(_0498_));
 sg13g2_nand2_1 _3157_ (.Y(_0499_),
    .A(net734),
    .B(_0498_));
 sg13g2_xnor2_1 _3158_ (.Y(_0500_),
    .A(net734),
    .B(_0498_));
 sg13g2_or2_1 _3159_ (.X(_0501_),
    .B(_0500_),
    .A(_0497_));
 sg13g2_a21oi_1 _3160_ (.A1(_2360_),
    .A2(_0305_),
    .Y(_0502_),
    .B1(_2362_));
 sg13g2_or3_1 _3161_ (.A(_0306_),
    .B(_0356_),
    .C(_0502_),
    .X(_0503_));
 sg13g2_nand2_1 _3162_ (.Y(_0504_),
    .A(_1922_),
    .B(_0503_));
 sg13g2_nor2_1 _3163_ (.A(_1922_),
    .B(_0503_),
    .Y(_0505_));
 sg13g2_xnor2_1 _3164_ (.Y(_0506_),
    .A(_1922_),
    .B(_0503_));
 sg13g2_and3_2 _3165_ (.X(_0507_),
    .A(_0352_),
    .B(_0353_),
    .C(net558));
 sg13g2_nand2_1 _3166_ (.Y(_0508_),
    .A(net735),
    .B(_0507_));
 sg13g2_xnor2_1 _3167_ (.Y(_0509_),
    .A(net735),
    .B(_0507_));
 sg13g2_nor3_1 _3168_ (.A(_0501_),
    .B(_0506_),
    .C(_0509_),
    .Y(_0510_));
 sg13g2_o21ai_1 _3169_ (.B1(_0510_),
    .Y(_0511_),
    .A1(_0484_),
    .A2(_0493_));
 sg13g2_o21ai_1 _3170_ (.B1(_0508_),
    .Y(_0512_),
    .A1(_1922_),
    .A2(_0503_));
 sg13g2_nand2_1 _3171_ (.Y(_0513_),
    .A(_0504_),
    .B(_0512_));
 sg13g2_nor2_1 _3172_ (.A(_0501_),
    .B(_0513_),
    .Y(_0514_));
 sg13g2_o21ai_1 _3173_ (.B1(_0499_),
    .Y(_0515_),
    .A1(_1929_),
    .A2(_0495_));
 sg13g2_a21oi_1 _3174_ (.A1(_0496_),
    .A2(_0515_),
    .Y(_0516_),
    .B1(_0514_));
 sg13g2_nand2_1 _3175_ (.Y(_0517_),
    .A(_0511_),
    .B(_0516_));
 sg13g2_a21oi_2 _3176_ (.B1(_0310_),
    .Y(_0518_),
    .A2(_0347_),
    .A1(net561));
 sg13g2_nand2_1 _3177_ (.Y(_0519_),
    .A(net733),
    .B(_0518_));
 sg13g2_xnor2_1 _3178_ (.Y(_0520_),
    .A(net733),
    .B(_0518_));
 sg13g2_xnor2_1 _3179_ (.Y(_0521_),
    .A(_2353_),
    .B(_0301_));
 sg13g2_and2_1 _3180_ (.A(net558),
    .B(_0521_),
    .X(_0522_));
 sg13g2_nor2_1 _3181_ (.A(net732),
    .B(_0522_),
    .Y(_0523_));
 sg13g2_nand2_1 _3182_ (.Y(_0524_),
    .A(net732),
    .B(_0522_));
 sg13g2_nand2b_1 _3183_ (.Y(_0525_),
    .B(_0524_),
    .A_N(_0523_));
 sg13g2_or2_1 _3184_ (.X(_0526_),
    .B(_0525_),
    .A(_0520_));
 sg13g2_a21oi_1 _3185_ (.A1(_0511_),
    .A2(_0516_),
    .Y(_0527_),
    .B1(_0526_));
 sg13g2_o21ai_1 _3186_ (.B1(_0524_),
    .Y(_0528_),
    .A1(_0519_),
    .A2(_0523_));
 sg13g2_xnor2_1 _3187_ (.Y(_0529_),
    .A(_1935_),
    .B(_0354_));
 sg13g2_o21ai_1 _3188_ (.B1(_0529_),
    .Y(_0530_),
    .A1(_0527_),
    .A2(_0528_));
 sg13g2_xor2_1 _3189_ (.B(_0362_),
    .A(\reg_a[0] ),
    .X(_0531_));
 sg13g2_a21o_2 _3190_ (.A2(_0530_),
    .A1(_0355_),
    .B1(_0531_),
    .X(_0532_));
 sg13g2_nand3_1 _3191_ (.B(_0530_),
    .C(_0531_),
    .A(_0355_),
    .Y(_0533_));
 sg13g2_nand2_1 _3192_ (.Y(_0534_),
    .A(_0532_),
    .B(_0533_));
 sg13g2_or3_1 _3193_ (.A(_0527_),
    .B(_0528_),
    .C(_0529_),
    .X(_0535_));
 sg13g2_nand2b_1 _3194_ (.Y(_0536_),
    .B(_0517_),
    .A_N(_0520_));
 sg13g2_nand2_1 _3195_ (.Y(_0537_),
    .A(_0519_),
    .B(_0536_));
 sg13g2_xnor2_1 _3196_ (.Y(_0538_),
    .A(_0525_),
    .B(_0537_));
 sg13g2_xor2_1 _3197_ (.B(_0520_),
    .A(_0517_),
    .X(_0539_));
 sg13g2_o21ai_1 _3198_ (.B1(_0508_),
    .Y(_0540_),
    .A1(_0494_),
    .A2(_0509_));
 sg13g2_o21ai_1 _3199_ (.B1(_0504_),
    .Y(_0541_),
    .A1(_0505_),
    .A2(_0540_));
 sg13g2_o21ai_1 _3200_ (.B1(_0499_),
    .Y(_0542_),
    .A1(_0500_),
    .A2(_0541_));
 sg13g2_xnor2_1 _3201_ (.Y(_0543_),
    .A(_0497_),
    .B(_0542_));
 sg13g2_xor2_1 _3202_ (.B(_0541_),
    .A(_0500_),
    .X(_0544_));
 sg13g2_xor2_1 _3203_ (.B(_0509_),
    .A(_0494_),
    .X(_0545_));
 sg13g2_xnor2_1 _3204_ (.Y(_0546_),
    .A(_0506_),
    .B(_0540_));
 sg13g2_a21oi_1 _3205_ (.A1(_0445_),
    .A2(_0482_),
    .Y(_0547_),
    .B1(_0488_));
 sg13g2_or2_1 _3206_ (.X(_0548_),
    .B(_0547_),
    .A(_0459_));
 sg13g2_a21oi_1 _3207_ (.A1(_0490_),
    .A2(_0548_),
    .Y(_0549_),
    .B1(_0456_));
 sg13g2_nand2b_1 _3208_ (.Y(_0550_),
    .B(_0549_),
    .A_N(_0453_));
 sg13g2_nand2_1 _3209_ (.Y(_0551_),
    .A(_0452_),
    .B(_0550_));
 sg13g2_xor2_1 _3210_ (.B(_0551_),
    .A(_0449_),
    .X(_0552_));
 sg13g2_xnor2_1 _3211_ (.Y(_0553_),
    .A(_0453_),
    .B(_0549_));
 sg13g2_inv_1 _3212_ (.Y(_0554_),
    .A(_0553_));
 sg13g2_xnor2_1 _3213_ (.Y(_0555_),
    .A(_0459_),
    .B(_0547_));
 sg13g2_nand2b_1 _3214_ (.Y(_0556_),
    .B(_0548_),
    .A_N(_0458_));
 sg13g2_xor2_1 _3215_ (.B(_0556_),
    .A(_0462_),
    .X(_0557_));
 sg13g2_or2_1 _3216_ (.X(_0558_),
    .B(_0557_),
    .A(_0555_));
 sg13g2_a21oi_1 _3217_ (.A1(_0436_),
    .A2(_0444_),
    .Y(_0559_),
    .B1(_0478_));
 sg13g2_a21oi_1 _3218_ (.A1(net740),
    .A2(_0476_),
    .Y(_0560_),
    .B1(_0559_));
 sg13g2_o21ai_1 _3219_ (.B1(_0474_),
    .Y(_0561_),
    .A1(_0485_),
    .A2(_0559_));
 sg13g2_o21ai_1 _3220_ (.B1(_0469_),
    .Y(_0562_),
    .A1(_0470_),
    .A2(_0561_));
 sg13g2_xor2_1 _3221_ (.B(_0562_),
    .A(_0465_),
    .X(_0563_));
 sg13g2_xor2_1 _3222_ (.B(_0561_),
    .A(_0471_),
    .X(_0564_));
 sg13g2_xnor2_1 _3223_ (.Y(_0565_),
    .A(_0481_),
    .B(_0560_));
 sg13g2_nor2_1 _3224_ (.A(_0564_),
    .B(_0565_),
    .Y(_0566_));
 sg13g2_xnor2_1 _3225_ (.Y(_0567_),
    .A(\reg_a[3] ),
    .B(_0371_));
 sg13g2_nand2_1 _3226_ (.Y(_0568_),
    .A(_0368_),
    .B(_0370_));
 sg13g2_xnor2_1 _3227_ (.Y(_0569_),
    .A(_0567_),
    .B(_0568_));
 sg13g2_xnor2_1 _3228_ (.Y(_0570_),
    .A(_0363_),
    .B(_0365_));
 sg13g2_xor2_1 _3229_ (.B(_0369_),
    .A(_0366_),
    .X(_0571_));
 sg13g2_or2_1 _3230_ (.X(_0572_),
    .B(_0570_),
    .A(_0532_));
 sg13g2_nor4_2 _3231_ (.A(_0532_),
    .B(_0569_),
    .C(_0570_),
    .Y(_0573_),
    .D(_0571_));
 sg13g2_or3_1 _3232_ (.A(_0569_),
    .B(_0571_),
    .C(_0572_),
    .X(_0574_));
 sg13g2_and2_1 _3233_ (.A(_0374_),
    .B(_0388_),
    .X(_0575_));
 sg13g2_o21ai_1 _3234_ (.B1(_0390_),
    .Y(_0576_),
    .A1(_0394_),
    .A2(_0575_));
 sg13g2_o21ai_1 _3235_ (.B1(_0382_),
    .Y(_0577_),
    .A1(_0384_),
    .A2(_0576_));
 sg13g2_xor2_1 _3236_ (.B(_0577_),
    .A(_0378_),
    .X(_0578_));
 sg13g2_xnor2_1 _3237_ (.Y(_0579_),
    .A(_0384_),
    .B(_0576_));
 sg13g2_xnor2_1 _3238_ (.Y(_0580_),
    .A(_0374_),
    .B(_0388_));
 sg13g2_a21oi_1 _3239_ (.A1(\reg_a[4] ),
    .A2(_0387_),
    .Y(_0581_),
    .B1(_0575_));
 sg13g2_xor2_1 _3240_ (.B(_0581_),
    .A(_0391_),
    .X(_0582_));
 sg13g2_nor3_1 _3241_ (.A(_0579_),
    .B(_0580_),
    .C(_0582_),
    .Y(_0583_));
 sg13g2_and2_1 _3242_ (.A(_0578_),
    .B(_0583_),
    .X(_0584_));
 sg13g2_nand2_1 _3243_ (.Y(_0585_),
    .A(_0573_),
    .B(_0584_));
 sg13g2_o21ai_1 _3244_ (.B1(_0416_),
    .Y(_0586_),
    .A1(_0393_),
    .A2(_0397_));
 sg13g2_o21ai_1 _3245_ (.B1(_0440_),
    .Y(_0587_),
    .A1(_0411_),
    .A2(_0586_));
 sg13g2_nand2_1 _3246_ (.Y(_0588_),
    .A(_0429_),
    .B(_0587_));
 sg13g2_and2_1 _3247_ (.A(_0428_),
    .B(_0588_),
    .X(_0589_));
 sg13g2_a21oi_1 _3248_ (.A1(_0432_),
    .A2(_0589_),
    .Y(_0590_),
    .B1(_0431_));
 sg13g2_a21oi_1 _3249_ (.A1(_0425_),
    .A2(_0590_),
    .Y(_0591_),
    .B1(_0424_));
 sg13g2_xor2_1 _3250_ (.B(_0591_),
    .A(_0422_),
    .X(_0592_));
 sg13g2_xnor2_1 _3251_ (.Y(_0593_),
    .A(_0425_),
    .B(_0590_));
 sg13g2_a21oi_1 _3252_ (.A1(_0438_),
    .A2(_0586_),
    .Y(_0594_),
    .B1(_0405_));
 sg13g2_xor2_1 _3253_ (.B(_0594_),
    .A(_0408_),
    .X(_0595_));
 sg13g2_or3_1 _3254_ (.A(_0393_),
    .B(_0397_),
    .C(_0416_),
    .X(_0596_));
 sg13g2_and2_1 _3255_ (.A(_0586_),
    .B(_0596_),
    .X(_0597_));
 sg13g2_nor2b_1 _3256_ (.A(_0405_),
    .B_N(_0410_),
    .Y(_0598_));
 sg13g2_nand2_1 _3257_ (.Y(_0599_),
    .A(_0414_),
    .B(_0586_));
 sg13g2_xnor2_1 _3258_ (.Y(_0600_),
    .A(_0598_),
    .B(_0599_));
 sg13g2_nand3b_1 _3259_ (.B(_0597_),
    .C(_0595_),
    .Y(_0601_),
    .A_N(_0600_));
 sg13g2_a21oi_1 _3260_ (.A1(_0408_),
    .A2(_0594_),
    .Y(_0602_),
    .B1(_0406_));
 sg13g2_xnor2_1 _3261_ (.Y(_0603_),
    .A(_0402_),
    .B(_0602_));
 sg13g2_nor2_1 _3262_ (.A(_0601_),
    .B(_0603_),
    .Y(_0604_));
 sg13g2_inv_1 _3263_ (.Y(_0605_),
    .A(_0604_));
 sg13g2_xnor2_1 _3264_ (.Y(_0606_),
    .A(_0429_),
    .B(_0587_));
 sg13g2_xor2_1 _3265_ (.B(_0589_),
    .A(_0433_),
    .X(_0607_));
 sg13g2_nor4_1 _3266_ (.A(_0593_),
    .B(_0605_),
    .C(_0606_),
    .D(_0607_),
    .Y(_0608_));
 sg13g2_nand4_1 _3267_ (.B(_0584_),
    .C(_0592_),
    .A(_0573_),
    .Y(_0609_),
    .D(_0608_));
 sg13g2_xnor2_1 _3268_ (.Y(_0610_),
    .A(_0445_),
    .B(_0478_));
 sg13g2_xor2_1 _3269_ (.B(_0478_),
    .A(_0445_),
    .X(_0611_));
 sg13g2_nor2_1 _3270_ (.A(_0609_),
    .B(_0611_),
    .Y(_0612_));
 sg13g2_nand3_1 _3271_ (.B(_0566_),
    .C(_0610_),
    .A(_0563_),
    .Y(_0613_));
 sg13g2_or2_1 _3272_ (.X(_0614_),
    .B(_0613_),
    .A(_0609_));
 sg13g2_nor2_1 _3273_ (.A(_0558_),
    .B(_0614_),
    .Y(_0615_));
 sg13g2_nand2_1 _3274_ (.Y(_0616_),
    .A(_0553_),
    .B(_0615_));
 sg13g2_nor4_1 _3275_ (.A(_0552_),
    .B(_0554_),
    .C(_0558_),
    .D(_0614_),
    .Y(_0617_));
 sg13g2_and3_2 _3276_ (.X(_0618_),
    .A(_0545_),
    .B(_0546_),
    .C(_0617_));
 sg13g2_and2_1 _3277_ (.A(_0544_),
    .B(_0618_),
    .X(_0619_));
 sg13g2_nand2_1 _3278_ (.Y(_0620_),
    .A(_0543_),
    .B(_0619_));
 sg13g2_nor2_1 _3279_ (.A(_0539_),
    .B(_0620_),
    .Y(_0621_));
 sg13g2_a22oi_1 _3280_ (.Y(_0622_),
    .B1(_0538_),
    .B2(_0621_),
    .A2(_0535_),
    .A1(_0530_));
 sg13g2_xor2_1 _3281_ (.B(_0620_),
    .A(_0539_),
    .X(_0623_));
 sg13g2_xor2_1 _3282_ (.B(_0619_),
    .A(_0543_),
    .X(_0624_));
 sg13g2_xor2_1 _3283_ (.B(_0616_),
    .A(_0552_),
    .X(_0625_));
 sg13g2_xor2_1 _3284_ (.B(_0614_),
    .A(_0555_),
    .X(_0626_));
 sg13g2_nand3_1 _3285_ (.B(_0584_),
    .C(_0604_),
    .A(_0573_),
    .Y(_0627_));
 sg13g2_nor2_1 _3286_ (.A(_0606_),
    .B(_0627_),
    .Y(_0628_));
 sg13g2_nor3_1 _3287_ (.A(_0606_),
    .B(_0607_),
    .C(_0627_),
    .Y(_0629_));
 sg13g2_nor2b_1 _3288_ (.A(_0593_),
    .B_N(_0629_),
    .Y(_0630_));
 sg13g2_xnor2_1 _3289_ (.Y(_0631_),
    .A(_0593_),
    .B(_0629_));
 sg13g2_nor3_1 _3290_ (.A(_0574_),
    .B(_0580_),
    .C(_0582_),
    .Y(_0632_));
 sg13g2_o21ai_1 _3291_ (.B1(_0582_),
    .Y(_0633_),
    .A1(_0574_),
    .A2(_0580_));
 sg13g2_nand2b_1 _3292_ (.Y(_0634_),
    .B(_0633_),
    .A_N(_0632_));
 sg13g2_nand3_1 _3293_ (.B(_0584_),
    .C(_0597_),
    .A(_0573_),
    .Y(_0635_));
 sg13g2_xnor2_1 _3294_ (.Y(_0636_),
    .A(_0585_),
    .B(_0597_));
 sg13g2_xnor2_1 _3295_ (.Y(_0637_),
    .A(_0609_),
    .B(_0610_));
 sg13g2_xnor2_1 _3296_ (.Y(_0638_),
    .A(_0606_),
    .B(_0627_));
 sg13g2_nor2_1 _3297_ (.A(_0600_),
    .B(_0635_),
    .Y(_0639_));
 sg13g2_nand2_1 _3298_ (.Y(_0640_),
    .A(_0595_),
    .B(_0639_));
 sg13g2_xnor2_1 _3299_ (.Y(_0641_),
    .A(_0595_),
    .B(_0639_));
 sg13g2_xnor2_1 _3300_ (.Y(_0642_),
    .A(_0545_),
    .B(_0617_));
 sg13g2_nand2b_1 _3301_ (.Y(_0643_),
    .B(_0632_),
    .A_N(_0579_));
 sg13g2_xnor2_1 _3302_ (.Y(_0644_),
    .A(_0579_),
    .B(_0632_));
 sg13g2_xor2_1 _3303_ (.B(_0572_),
    .A(_0571_),
    .X(_0645_));
 sg13g2_nor2_1 _3304_ (.A(_0554_),
    .B(_0557_),
    .Y(_0646_));
 sg13g2_and3_1 _3305_ (.X(_0647_),
    .A(_0563_),
    .B(_0566_),
    .C(_0637_));
 sg13g2_and4_1 _3306_ (.A(_0625_),
    .B(_0626_),
    .C(_0646_),
    .D(_0647_),
    .X(_0648_));
 sg13g2_or2_1 _3307_ (.X(_0649_),
    .B(_0641_),
    .A(_0603_));
 sg13g2_o21ai_1 _3308_ (.B1(_0569_),
    .Y(_0650_),
    .A1(_0571_),
    .A2(_0572_));
 sg13g2_nand2_1 _3309_ (.Y(_0651_),
    .A(_0574_),
    .B(_0650_));
 sg13g2_nor2_1 _3310_ (.A(_0534_),
    .B(_0570_),
    .Y(_0652_));
 sg13g2_nand4_1 _3311_ (.B(_0645_),
    .C(_0650_),
    .A(_0574_),
    .Y(_0653_),
    .D(_0652_));
 sg13g2_nor3_1 _3312_ (.A(_0580_),
    .B(_0634_),
    .C(_0653_),
    .Y(_0654_));
 sg13g2_nor2b_1 _3313_ (.A(_0600_),
    .B_N(_0636_),
    .Y(_0655_));
 sg13g2_nand4_1 _3314_ (.B(_0644_),
    .C(_0654_),
    .A(_0578_),
    .Y(_0656_),
    .D(_0655_));
 sg13g2_nor4_1 _3315_ (.A(_0607_),
    .B(_0638_),
    .C(_0649_),
    .D(_0656_),
    .Y(_0657_));
 sg13g2_and4_1 _3316_ (.A(_0592_),
    .B(_0631_),
    .C(_0648_),
    .D(_0657_),
    .X(_0658_));
 sg13g2_nand2_1 _3317_ (.Y(_0659_),
    .A(_0544_),
    .B(_0546_));
 sg13g2_nor2_1 _3318_ (.A(_0642_),
    .B(_0659_),
    .Y(_0660_));
 sg13g2_and2_1 _3319_ (.A(_0624_),
    .B(_0660_),
    .X(_0661_));
 sg13g2_nand4_1 _3320_ (.B(_0623_),
    .C(_0658_),
    .A(_0538_),
    .Y(_0662_),
    .D(_0661_));
 sg13g2_or2_1 _3321_ (.X(_0663_),
    .B(_0662_),
    .A(_0622_));
 sg13g2_inv_2 _3322_ (.Y(_0664_),
    .A(net551));
 sg13g2_o21ai_1 _3323_ (.B1(net715),
    .Y(_0665_),
    .A1(_0534_),
    .A2(_0664_));
 sg13g2_and2_1 _3324_ (.A(net704),
    .B(net696),
    .X(_0666_));
 sg13g2_nand2_1 _3325_ (.Y(_0667_),
    .A(net704),
    .B(net695));
 sg13g2_a21oi_1 _3326_ (.A1(net700),
    .A2(_0362_),
    .Y(_0668_),
    .B1(net635));
 sg13g2_nand2_1 _3327_ (.Y(_0669_),
    .A(_0665_),
    .B(_0668_));
 sg13g2_and2_1 _3328_ (.A(net760),
    .B(net592),
    .X(_0670_));
 sg13g2_nand2_1 _3329_ (.Y(_0671_),
    .A(net760),
    .B(net592));
 sg13g2_nor2_1 _3330_ (.A(net4),
    .B(net3),
    .Y(_0672_));
 sg13g2_nand2_1 _3331_ (.Y(_0673_),
    .A(net2),
    .B(_0672_));
 sg13g2_nor2_1 _3332_ (.A(net1),
    .B(_0673_),
    .Y(_0674_));
 sg13g2_nand3_1 _3333_ (.B(net2),
    .C(_0672_),
    .A(_1962_),
    .Y(_0675_));
 sg13g2_nor4_2 _3334_ (.A(_1962_),
    .B(net2),
    .C(net4),
    .Y(_0676_),
    .D(net3));
 sg13g2_nor3_2 _3335_ (.A(_2085_),
    .B(_0674_),
    .C(_0676_),
    .Y(_0677_));
 sg13g2_nor2b_2 _3336_ (.A(_0677_),
    .B_N(net9),
    .Y(_0678_));
 sg13g2_nand2b_1 _3337_ (.Y(_0679_),
    .B(net9),
    .A_N(_0677_));
 sg13g2_nor2_2 _3338_ (.A(net685),
    .B(net627),
    .Y(_0680_));
 sg13g2_nand2_2 _3339_ (.Y(_0681_),
    .A(net696),
    .B(net631));
 sg13g2_mux2_1 _3340_ (.A0(\reg_a[0] ),
    .A1(net744),
    .S(net574),
    .X(_0682_));
 sg13g2_o21ai_1 _3341_ (.B1(net636),
    .Y(_0683_),
    .A1(_0680_),
    .A2(_0682_));
 sg13g2_nand2_1 _3342_ (.Y(_0684_),
    .A(\reg_a[0] ),
    .B(\reg_b[0] ));
 sg13g2_xor2_1 _3343_ (.B(\reg_b[0] ),
    .A(\reg_a[0] ),
    .X(_0685_));
 sg13g2_inv_2 _3344_ (.Y(_0686_),
    .A(_0685_));
 sg13g2_xnor2_1 _3345_ (.Y(_0687_),
    .A(\reg_a[30] ),
    .B(\reg_b[30] ));
 sg13g2_nor2_1 _3346_ (.A(\reg_a[29] ),
    .B(net722),
    .Y(_0688_));
 sg13g2_and2_1 _3347_ (.A(net733),
    .B(\reg_b[28] ),
    .X(_0689_));
 sg13g2_xnor2_1 _3348_ (.Y(_0690_),
    .A(net733),
    .B(\reg_b[28] ));
 sg13g2_inv_1 _3349_ (.Y(_0691_),
    .A(_0690_));
 sg13g2_nor2_1 _3350_ (.A(\reg_a[27] ),
    .B(net723),
    .Y(_0692_));
 sg13g2_or2_1 _3351_ (.X(_0693_),
    .B(net724),
    .A(\reg_a[25] ));
 sg13g2_nor2_1 _3352_ (.A(\reg_a[19] ),
    .B(net727),
    .Y(_0694_));
 sg13g2_nand2_1 _3353_ (.Y(_0695_),
    .A(\reg_a[19] ),
    .B(net727));
 sg13g2_and2_1 _3354_ (.A(\reg_a[18] ),
    .B(net728),
    .X(_0696_));
 sg13g2_nand2_1 _3355_ (.Y(_0697_),
    .A(\reg_a[18] ),
    .B(net728));
 sg13g2_nand2_1 _3356_ (.Y(_0698_),
    .A(net740),
    .B(\reg_b[16] ));
 sg13g2_nor2_1 _3357_ (.A(\reg_a[15] ),
    .B(\reg_b[15] ),
    .Y(_0699_));
 sg13g2_nand2_1 _3358_ (.Y(_0700_),
    .A(\reg_a[15] ),
    .B(\reg_b[15] ));
 sg13g2_nand2_1 _3359_ (.Y(_0701_),
    .A(\reg_a[14] ),
    .B(\reg_b[14] ));
 sg13g2_xor2_1 _3360_ (.B(\reg_b[14] ),
    .A(\reg_a[14] ),
    .X(_0702_));
 sg13g2_nand2_1 _3361_ (.Y(_0703_),
    .A(net741),
    .B(net730));
 sg13g2_nor2_1 _3362_ (.A(net741),
    .B(net730),
    .Y(_0704_));
 sg13g2_nand2_1 _3363_ (.Y(_0705_),
    .A(net742),
    .B(\reg_b[12] ));
 sg13g2_o21ai_1 _3364_ (.B1(_0703_),
    .Y(_0706_),
    .A1(_0704_),
    .A2(_0705_));
 sg13g2_or2_1 _3365_ (.X(_0707_),
    .B(\reg_b[11] ),
    .A(\reg_a[11] ));
 sg13g2_nand2_1 _3366_ (.Y(_0708_),
    .A(\reg_a[11] ),
    .B(\reg_b[11] ));
 sg13g2_and2_1 _3367_ (.A(net743),
    .B(\reg_b[10] ),
    .X(_0709_));
 sg13g2_nor2_1 _3368_ (.A(\reg_a[9] ),
    .B(net731),
    .Y(_0710_));
 sg13g2_and2_1 _3369_ (.A(net744),
    .B(\reg_b[8] ),
    .X(_0711_));
 sg13g2_xor2_1 _3370_ (.B(\reg_b[8] ),
    .A(net744),
    .X(_0712_));
 sg13g2_nand2_1 _3371_ (.Y(_0713_),
    .A(net745),
    .B(\reg_b[7] ));
 sg13g2_nor2_1 _3372_ (.A(net745),
    .B(\reg_b[7] ),
    .Y(_0714_));
 sg13g2_xor2_1 _3373_ (.B(\reg_b[7] ),
    .A(net745),
    .X(_0715_));
 sg13g2_and2_1 _3374_ (.A(\reg_a[6] ),
    .B(\reg_b[6] ),
    .X(_0716_));
 sg13g2_xor2_1 _3375_ (.B(\reg_b[6] ),
    .A(\reg_a[6] ),
    .X(_0717_));
 sg13g2_xnor2_1 _3376_ (.Y(_0718_),
    .A(\reg_a[6] ),
    .B(\reg_b[6] ));
 sg13g2_nand2_1 _3377_ (.Y(_0719_),
    .A(\reg_a[5] ),
    .B(\reg_b[5] ));
 sg13g2_nor2b_1 _3378_ (.A(\reg_b[5] ),
    .B_N(\reg_a[5] ),
    .Y(_0720_));
 sg13g2_xnor2_1 _3379_ (.Y(_0721_),
    .A(\reg_a[5] ),
    .B(\reg_b[5] ));
 sg13g2_inv_1 _3380_ (.Y(_0722_),
    .A(_0721_));
 sg13g2_and2_1 _3381_ (.A(\reg_a[4] ),
    .B(\reg_b[4] ),
    .X(_0723_));
 sg13g2_nor2b_1 _3382_ (.A(\reg_b[4] ),
    .B_N(\reg_a[4] ),
    .Y(_0724_));
 sg13g2_nand2b_1 _3383_ (.Y(_0725_),
    .B(\reg_b[4] ),
    .A_N(\reg_a[4] ));
 sg13g2_nand2b_2 _3384_ (.Y(_0726_),
    .B(_0725_),
    .A_N(_0724_));
 sg13g2_nand2_1 _3385_ (.Y(_0727_),
    .A(\reg_a[3] ),
    .B(\reg_b[3] ));
 sg13g2_nor2_1 _3386_ (.A(_1928_),
    .B(\reg_b[3] ),
    .Y(_0728_));
 sg13g2_xnor2_1 _3387_ (.Y(_0729_),
    .A(\reg_a[3] ),
    .B(\reg_b[3] ));
 sg13g2_and2_1 _3388_ (.A(net746),
    .B(\reg_b[2] ),
    .X(_0730_));
 sg13g2_nand2b_1 _3389_ (.Y(_0731_),
    .B(net746),
    .A_N(\reg_b[2] ));
 sg13g2_xor2_1 _3390_ (.B(\reg_b[2] ),
    .A(net746),
    .X(_0732_));
 sg13g2_nand2_1 _3391_ (.Y(_0733_),
    .A(net747),
    .B(\reg_b[1] ));
 sg13g2_xnor2_1 _3392_ (.Y(_0734_),
    .A(net747),
    .B(\reg_b[1] ));
 sg13g2_o21ai_1 _3393_ (.B1(_0733_),
    .Y(_0735_),
    .A1(_0684_),
    .A2(_0734_));
 sg13g2_a21oi_1 _3394_ (.A1(_0732_),
    .A2(_0735_),
    .Y(_0736_),
    .B1(_0730_));
 sg13g2_o21ai_1 _3395_ (.B1(_0727_),
    .Y(_0737_),
    .A1(_0729_),
    .A2(_0736_));
 sg13g2_a21oi_1 _3396_ (.A1(_0726_),
    .A2(_0737_),
    .Y(_0738_),
    .B1(_0723_));
 sg13g2_o21ai_1 _3397_ (.B1(_0719_),
    .Y(_0739_),
    .A1(_0721_),
    .A2(_0738_));
 sg13g2_a21oi_2 _3398_ (.B1(_0716_),
    .Y(_0740_),
    .A2(_0739_),
    .A1(_0717_));
 sg13g2_o21ai_1 _3399_ (.B1(_0713_),
    .Y(_0741_),
    .A1(_0714_),
    .A2(_0740_));
 sg13g2_a21oi_1 _3400_ (.A1(_0712_),
    .A2(_0741_),
    .Y(_0742_),
    .B1(_0711_));
 sg13g2_a221oi_1 _3401_ (.B2(_0741_),
    .C1(_0711_),
    .B1(_0712_),
    .A1(\reg_a[9] ),
    .Y(_0743_),
    .A2(net731));
 sg13g2_nor2_1 _3402_ (.A(_0710_),
    .B(_0743_),
    .Y(_0744_));
 sg13g2_xor2_1 _3403_ (.B(\reg_b[10] ),
    .A(net743),
    .X(_0745_));
 sg13g2_a21oi_1 _3404_ (.A1(_0744_),
    .A2(_0745_),
    .Y(_0746_),
    .B1(_0709_));
 sg13g2_nand2_1 _3405_ (.Y(_0747_),
    .A(_0707_),
    .B(_0709_));
 sg13g2_nand2_1 _3406_ (.Y(_0748_),
    .A(_0707_),
    .B(_0708_));
 sg13g2_inv_2 _3407_ (.Y(_0749_),
    .A(_0748_));
 sg13g2_nand2_1 _3408_ (.Y(_0750_),
    .A(_0745_),
    .B(_0749_));
 sg13g2_or3_1 _3409_ (.A(_0710_),
    .B(_0743_),
    .C(_0750_),
    .X(_0751_));
 sg13g2_nand3_1 _3410_ (.B(_0747_),
    .C(_0751_),
    .A(_0708_),
    .Y(_0752_));
 sg13g2_xor2_1 _3411_ (.B(net730),
    .A(net741),
    .X(_0753_));
 sg13g2_inv_1 _3412_ (.Y(_0754_),
    .A(_0753_));
 sg13g2_xor2_1 _3413_ (.B(\reg_b[12] ),
    .A(net742),
    .X(_0755_));
 sg13g2_and2_1 _3414_ (.A(_0753_),
    .B(_0755_),
    .X(_0756_));
 sg13g2_a21o_1 _3415_ (.A2(_0756_),
    .A1(_0752_),
    .B1(_0706_),
    .X(_0757_));
 sg13g2_nand2_1 _3416_ (.Y(_0758_),
    .A(_0702_),
    .B(_0757_));
 sg13g2_nand2_1 _3417_ (.Y(_0759_),
    .A(_0701_),
    .B(_0758_));
 sg13g2_o21ai_1 _3418_ (.B1(_0700_),
    .Y(_0760_),
    .A1(_0699_),
    .A2(_0701_));
 sg13g2_nor2b_2 _3419_ (.A(_0699_),
    .B_N(_0700_),
    .Y(_0761_));
 sg13g2_and2_1 _3420_ (.A(_0702_),
    .B(_0761_),
    .X(_0762_));
 sg13g2_and2_1 _3421_ (.A(_0756_),
    .B(_0762_),
    .X(_0763_));
 sg13g2_a221oi_1 _3422_ (.B2(_0752_),
    .C1(_0760_),
    .B1(_0763_),
    .A1(_0706_),
    .Y(_0764_),
    .A2(_0762_));
 sg13g2_xnor2_1 _3423_ (.Y(_0765_),
    .A(net740),
    .B(\reg_b[16] ));
 sg13g2_o21ai_1 _3424_ (.B1(_0698_),
    .Y(_0766_),
    .A1(_0764_),
    .A2(_0765_));
 sg13g2_a21oi_1 _3425_ (.A1(_1923_),
    .A2(_1924_),
    .Y(_0767_),
    .B1(_0698_));
 sg13g2_a21oi_1 _3426_ (.A1(\reg_a[17] ),
    .A2(net729),
    .Y(_0768_),
    .B1(_0767_));
 sg13g2_xnor2_1 _3427_ (.Y(_0769_),
    .A(\reg_a[17] ),
    .B(net729));
 sg13g2_or2_1 _3428_ (.X(_0770_),
    .B(_0769_),
    .A(_0765_));
 sg13g2_o21ai_1 _3429_ (.B1(_0768_),
    .Y(_0771_),
    .A1(_0764_),
    .A2(_0770_));
 sg13g2_or2_1 _3430_ (.X(_0772_),
    .B(net728),
    .A(\reg_a[18] ));
 sg13g2_nand2_2 _3431_ (.Y(_0773_),
    .A(_0697_),
    .B(_0772_));
 sg13g2_a21oi_1 _3432_ (.A1(_0771_),
    .A2(_0772_),
    .Y(_0774_),
    .B1(_0696_));
 sg13g2_o21ai_1 _3433_ (.B1(_0695_),
    .Y(_0775_),
    .A1(_0694_),
    .A2(_0697_));
 sg13g2_nand2b_2 _3434_ (.Y(_0776_),
    .B(_0695_),
    .A_N(_0694_));
 sg13g2_nor2_1 _3435_ (.A(_0773_),
    .B(_0776_),
    .Y(_0777_));
 sg13g2_a21o_2 _3436_ (.A2(_0777_),
    .A1(_0771_),
    .B1(_0775_),
    .X(_0778_));
 sg13g2_nand2_2 _3437_ (.Y(_0779_),
    .A(\reg_a[20] ),
    .B(\reg_b[20] ));
 sg13g2_or2_1 _3438_ (.X(_0780_),
    .B(\reg_b[20] ),
    .A(\reg_a[20] ));
 sg13g2_nand2_2 _3439_ (.Y(_0781_),
    .A(_0779_),
    .B(_0780_));
 sg13g2_nand3_1 _3440_ (.B(_0779_),
    .C(_0780_),
    .A(_0778_),
    .Y(_0782_));
 sg13g2_nand2_1 _3441_ (.Y(_0783_),
    .A(net739),
    .B(net726));
 sg13g2_nand3_1 _3442_ (.B(_0782_),
    .C(_0783_),
    .A(_0779_),
    .Y(_0784_));
 sg13g2_nand2_1 _3443_ (.Y(_0785_),
    .A(net738),
    .B(\reg_b[22] ));
 sg13g2_xor2_1 _3444_ (.B(\reg_b[22] ),
    .A(net738),
    .X(_0786_));
 sg13g2_xnor2_1 _3445_ (.Y(_0787_),
    .A(\reg_a[22] ),
    .B(\reg_b[22] ));
 sg13g2_nand2_1 _3446_ (.Y(_0788_),
    .A(net736),
    .B(net725));
 sg13g2_nor2_1 _3447_ (.A(net736),
    .B(net725),
    .Y(_0789_));
 sg13g2_xor2_1 _3448_ (.B(net725),
    .A(net737),
    .X(_0790_));
 sg13g2_nor2_1 _3449_ (.A(net739),
    .B(net726),
    .Y(_0791_));
 sg13g2_or2_1 _3450_ (.X(_0792_),
    .B(net726),
    .A(\reg_a[21] ));
 sg13g2_and2_1 _3451_ (.A(_0786_),
    .B(_0790_),
    .X(_0793_));
 sg13g2_inv_1 _3452_ (.Y(_0794_),
    .A(_0793_));
 sg13g2_o21ai_1 _3453_ (.B1(_0783_),
    .Y(_0795_),
    .A1(_0779_),
    .A2(_0791_));
 sg13g2_nand2_2 _3454_ (.Y(_0796_),
    .A(_0783_),
    .B(_0792_));
 sg13g2_nor3_1 _3455_ (.A(_0781_),
    .B(_0794_),
    .C(_0796_),
    .Y(_0797_));
 sg13g2_o21ai_1 _3456_ (.B1(_0788_),
    .Y(_0798_),
    .A1(_0785_),
    .A2(_0789_));
 sg13g2_a221oi_1 _3457_ (.B2(_0778_),
    .C1(_0798_),
    .B1(_0797_),
    .A1(_0793_),
    .Y(_0799_),
    .A2(_0795_));
 sg13g2_xor2_1 _3458_ (.B(\reg_b[24] ),
    .A(net735),
    .X(_0800_));
 sg13g2_nor2b_1 _3459_ (.A(_0799_),
    .B_N(_0800_),
    .Y(_0801_));
 sg13g2_a21oi_1 _3460_ (.A1(net735),
    .A2(\reg_b[24] ),
    .Y(_0802_),
    .B1(_0801_));
 sg13g2_and3_1 _3461_ (.X(_0803_),
    .A(net735),
    .B(\reg_b[24] ),
    .C(_0693_));
 sg13g2_a21oi_1 _3462_ (.A1(\reg_a[25] ),
    .A2(net724),
    .Y(_0804_),
    .B1(_0803_));
 sg13g2_xor2_1 _3463_ (.B(net724),
    .A(\reg_a[25] ),
    .X(_0805_));
 sg13g2_nand2_1 _3464_ (.Y(_0806_),
    .A(_0800_),
    .B(_0805_));
 sg13g2_o21ai_1 _3465_ (.B1(_0804_),
    .Y(_0807_),
    .A1(_0799_),
    .A2(_0806_));
 sg13g2_and2_1 _3466_ (.A(net734),
    .B(\reg_b[26] ),
    .X(_0808_));
 sg13g2_nand2_1 _3467_ (.Y(_0809_),
    .A(\reg_a[26] ),
    .B(\reg_b[26] ));
 sg13g2_xnor2_1 _3468_ (.Y(_0810_),
    .A(\reg_a[26] ),
    .B(\reg_b[26] ));
 sg13g2_inv_1 _3469_ (.Y(_0811_),
    .A(_0810_));
 sg13g2_nand2_1 _3470_ (.Y(_0812_),
    .A(\reg_a[27] ),
    .B(net723));
 sg13g2_o21ai_1 _3471_ (.B1(_0812_),
    .Y(_0813_),
    .A1(_0692_),
    .A2(_0809_));
 sg13g2_nand2b_2 _3472_ (.Y(_0814_),
    .B(_0812_),
    .A_N(_0692_));
 sg13g2_nor2_1 _3473_ (.A(_0810_),
    .B(_0814_),
    .Y(_0815_));
 sg13g2_a21o_2 _3474_ (.A2(_0815_),
    .A1(_0807_),
    .B1(_0813_),
    .X(_0816_));
 sg13g2_a21o_1 _3475_ (.A2(_0816_),
    .A1(_0691_),
    .B1(_0689_),
    .X(_0817_));
 sg13g2_a221oi_1 _3476_ (.B2(_0816_),
    .C1(_0689_),
    .B1(_0691_),
    .A1(net732),
    .Y(_0818_),
    .A2(net722));
 sg13g2_nor3_1 _3477_ (.A(_0687_),
    .B(_0688_),
    .C(_0818_),
    .Y(_0819_));
 sg13g2_a21oi_2 _3478_ (.B1(_0819_),
    .Y(_0820_),
    .A2(\reg_b[30] ),
    .A1(\reg_a[30] ));
 sg13g2_nor2_1 _3479_ (.A(_0686_),
    .B(_0820_),
    .Y(_0821_));
 sg13g2_xnor2_1 _3480_ (.Y(_0822_),
    .A(_0685_),
    .B(_0820_));
 sg13g2_o21ai_1 _3481_ (.B1(_0687_),
    .Y(_0823_),
    .A1(_0688_),
    .A2(_0818_));
 sg13g2_nor2b_1 _3482_ (.A(_0819_),
    .B_N(_0823_),
    .Y(_0824_));
 sg13g2_xor2_1 _3483_ (.B(net722),
    .A(net732),
    .X(_0825_));
 sg13g2_xnor2_1 _3484_ (.Y(_0826_),
    .A(_0817_),
    .B(_0825_));
 sg13g2_xnor2_1 _3485_ (.Y(_0827_),
    .A(_0690_),
    .B(_0816_));
 sg13g2_a21oi_1 _3486_ (.A1(_0807_),
    .A2(_0811_),
    .Y(_0828_),
    .B1(_0808_));
 sg13g2_xnor2_1 _3487_ (.Y(_0829_),
    .A(_0814_),
    .B(_0828_));
 sg13g2_xnor2_1 _3488_ (.Y(_0830_),
    .A(_0807_),
    .B(_0810_));
 sg13g2_xor2_1 _3489_ (.B(_0805_),
    .A(_0802_),
    .X(_0831_));
 sg13g2_xor2_1 _3490_ (.B(_0800_),
    .A(_0799_),
    .X(_0832_));
 sg13g2_nand2_1 _3491_ (.Y(_0833_),
    .A(_0779_),
    .B(_0782_));
 sg13g2_nand2_1 _3492_ (.Y(_0834_),
    .A(_0784_),
    .B(_0792_));
 sg13g2_o21ai_1 _3493_ (.B1(_0785_),
    .Y(_0835_),
    .A1(_0787_),
    .A2(_0834_));
 sg13g2_xnor2_1 _3494_ (.Y(_0836_),
    .A(_0790_),
    .B(_0835_));
 sg13g2_xnor2_1 _3495_ (.Y(_0837_),
    .A(_0786_),
    .B(_0834_));
 sg13g2_xor2_1 _3496_ (.B(_0833_),
    .A(_0796_),
    .X(_0838_));
 sg13g2_inv_1 _3497_ (.Y(_0839_),
    .A(_0838_));
 sg13g2_xnor2_1 _3498_ (.Y(_0840_),
    .A(_0774_),
    .B(_0776_));
 sg13g2_xnor2_1 _3499_ (.Y(_0841_),
    .A(_0771_),
    .B(_0773_));
 sg13g2_xor2_1 _3500_ (.B(_0769_),
    .A(_0766_),
    .X(_0842_));
 sg13g2_xnor2_1 _3501_ (.Y(_0843_),
    .A(_0764_),
    .B(_0765_));
 sg13g2_xnor2_1 _3502_ (.Y(_0844_),
    .A(_0759_),
    .B(_0761_));
 sg13g2_xnor2_1 _3503_ (.Y(_0845_),
    .A(_0702_),
    .B(_0757_));
 sg13g2_nand2_1 _3504_ (.Y(_0846_),
    .A(_0752_),
    .B(_0755_));
 sg13g2_nand2_1 _3505_ (.Y(_0847_),
    .A(_0705_),
    .B(_0846_));
 sg13g2_xnor2_1 _3506_ (.Y(_0848_),
    .A(_0754_),
    .B(_0847_));
 sg13g2_inv_1 _3507_ (.Y(_0849_),
    .A(_0848_));
 sg13g2_xnor2_1 _3508_ (.Y(_0850_),
    .A(_0746_),
    .B(_0749_));
 sg13g2_inv_1 _3509_ (.Y(_0851_),
    .A(_0850_));
 sg13g2_xor2_1 _3510_ (.B(net731),
    .A(\reg_a[9] ),
    .X(_0852_));
 sg13g2_xnor2_1 _3511_ (.Y(_0853_),
    .A(_0742_),
    .B(_0852_));
 sg13g2_inv_1 _3512_ (.Y(_0854_),
    .A(_0853_));
 sg13g2_xnor2_1 _3513_ (.Y(_0855_),
    .A(_0712_),
    .B(_0741_));
 sg13g2_xnor2_1 _3514_ (.Y(_0856_),
    .A(_0715_),
    .B(_0740_));
 sg13g2_inv_1 _3515_ (.Y(_0857_),
    .A(_0856_));
 sg13g2_xnor2_1 _3516_ (.Y(_0858_),
    .A(_0718_),
    .B(_0739_));
 sg13g2_inv_1 _3517_ (.Y(_0859_),
    .A(_0858_));
 sg13g2_xor2_1 _3518_ (.B(_0734_),
    .A(_0684_),
    .X(_0860_));
 sg13g2_inv_2 _3519_ (.Y(_0861_),
    .A(_0860_));
 sg13g2_nor3_1 _3520_ (.A(_0686_),
    .B(_0820_),
    .C(_0861_),
    .Y(_0862_));
 sg13g2_inv_1 _3521_ (.Y(_0863_),
    .A(_0862_));
 sg13g2_xnor2_1 _3522_ (.Y(_0864_),
    .A(_0732_),
    .B(_0735_));
 sg13g2_nor4_1 _3523_ (.A(_0686_),
    .B(_0820_),
    .C(_0861_),
    .D(_0864_),
    .Y(_0865_));
 sg13g2_xor2_1 _3524_ (.B(_0737_),
    .A(_0726_),
    .X(_0866_));
 sg13g2_xnor2_1 _3525_ (.Y(_0867_),
    .A(_0729_),
    .B(_0736_));
 sg13g2_xnor2_1 _3526_ (.Y(_0868_),
    .A(_0721_),
    .B(_0738_));
 sg13g2_nor2_1 _3527_ (.A(_0867_),
    .B(_0868_),
    .Y(_0869_));
 sg13g2_nor3_1 _3528_ (.A(_0863_),
    .B(_0864_),
    .C(_0867_),
    .Y(_0870_));
 sg13g2_nand3_1 _3529_ (.B(_0866_),
    .C(_0869_),
    .A(_0865_),
    .Y(_0871_));
 sg13g2_nor2_1 _3530_ (.A(_0859_),
    .B(_0871_),
    .Y(_0872_));
 sg13g2_nand2_1 _3531_ (.Y(_0873_),
    .A(_0856_),
    .B(_0872_));
 sg13g2_or4_1 _3532_ (.A(_0855_),
    .B(_0857_),
    .C(_0859_),
    .D(_0871_),
    .X(_0874_));
 sg13g2_nand2b_1 _3533_ (.Y(_0875_),
    .B(_0853_),
    .A_N(_0874_));
 sg13g2_xnor2_1 _3534_ (.Y(_0876_),
    .A(_0744_),
    .B(_0745_));
 sg13g2_nor2_1 _3535_ (.A(_0875_),
    .B(_0876_),
    .Y(_0877_));
 sg13g2_or4_1 _3536_ (.A(_0851_),
    .B(_0854_),
    .C(_0874_),
    .D(_0876_),
    .X(_0878_));
 sg13g2_xor2_1 _3537_ (.B(_0755_),
    .A(_0752_),
    .X(_0879_));
 sg13g2_inv_1 _3538_ (.Y(_0880_),
    .A(_0879_));
 sg13g2_nor2_1 _3539_ (.A(_0878_),
    .B(_0880_),
    .Y(_0881_));
 sg13g2_nand2_1 _3540_ (.Y(_0882_),
    .A(_0848_),
    .B(_0881_));
 sg13g2_or4_1 _3541_ (.A(_0845_),
    .B(_0849_),
    .C(_0878_),
    .D(_0880_),
    .X(_0883_));
 sg13g2_nor2_1 _3542_ (.A(_0844_),
    .B(_0883_),
    .Y(_0884_));
 sg13g2_nor3_1 _3543_ (.A(_0843_),
    .B(_0844_),
    .C(_0883_),
    .Y(_0885_));
 sg13g2_nor4_1 _3544_ (.A(_0842_),
    .B(_0843_),
    .C(_0844_),
    .D(_0883_),
    .Y(_0886_));
 sg13g2_nand2_1 _3545_ (.Y(_0887_),
    .A(_0841_),
    .B(_0886_));
 sg13g2_nor2_1 _3546_ (.A(_0840_),
    .B(_0887_),
    .Y(_0888_));
 sg13g2_xnor2_1 _3547_ (.Y(_0889_),
    .A(_0778_),
    .B(_0781_));
 sg13g2_nand2_1 _3548_ (.Y(_0890_),
    .A(_0888_),
    .B(_0889_));
 sg13g2_nor2_1 _3549_ (.A(_0838_),
    .B(_0890_),
    .Y(_0891_));
 sg13g2_nand4_1 _3550_ (.B(_0839_),
    .C(_0888_),
    .A(_0837_),
    .Y(_0892_),
    .D(_0889_));
 sg13g2_or2_1 _3551_ (.X(_0893_),
    .B(_0892_),
    .A(_0836_));
 sg13g2_nor2_1 _3552_ (.A(_0832_),
    .B(_0893_),
    .Y(_0894_));
 sg13g2_nor3_1 _3553_ (.A(_0831_),
    .B(_0832_),
    .C(_0893_),
    .Y(_0895_));
 sg13g2_and2_1 _3554_ (.A(_0830_),
    .B(_0895_),
    .X(_0896_));
 sg13g2_nor2b_2 _3555_ (.A(_0829_),
    .B_N(_0896_),
    .Y(_0897_));
 sg13g2_nand2_1 _3556_ (.Y(_0898_),
    .A(_0827_),
    .B(_0897_));
 sg13g2_nand3b_1 _3557_ (.B(_0827_),
    .C(_0897_),
    .Y(_0899_),
    .A_N(_0826_));
 sg13g2_nor2b_1 _3558_ (.A(_0824_),
    .B_N(_0899_),
    .Y(_0900_));
 sg13g2_xnor2_1 _3559_ (.Y(_0901_),
    .A(_0827_),
    .B(_0897_));
 sg13g2_xnor2_1 _3560_ (.Y(_0902_),
    .A(_0830_),
    .B(_0895_));
 sg13g2_xor2_1 _3561_ (.B(_0893_),
    .A(_0832_),
    .X(_0903_));
 sg13g2_xnor2_1 _3562_ (.Y(_0904_),
    .A(_0837_),
    .B(_0891_));
 sg13g2_xnor2_1 _3563_ (.Y(_0905_),
    .A(_0888_),
    .B(_0889_));
 sg13g2_xnor2_1 _3564_ (.Y(_0906_),
    .A(_0841_),
    .B(_0886_));
 sg13g2_xnor2_1 _3565_ (.Y(_0907_),
    .A(_0843_),
    .B(_0884_));
 sg13g2_xnor2_1 _3566_ (.Y(_0908_),
    .A(_0845_),
    .B(_0882_));
 sg13g2_xnor2_1 _3567_ (.Y(_0909_),
    .A(_0878_),
    .B(_0880_));
 sg13g2_xor2_1 _3568_ (.B(_0876_),
    .A(_0875_),
    .X(_0910_));
 sg13g2_xnor2_1 _3569_ (.Y(_0911_),
    .A(_0855_),
    .B(_0873_));
 sg13g2_xnor2_1 _3570_ (.Y(_0912_),
    .A(_0858_),
    .B(_0871_));
 sg13g2_nand2_1 _3571_ (.Y(_0913_),
    .A(_0866_),
    .B(_0870_));
 sg13g2_xor2_1 _3572_ (.B(_0870_),
    .A(_0866_),
    .X(_0914_));
 sg13g2_xnor2_1 _3573_ (.Y(_0915_),
    .A(_0862_),
    .B(_0864_));
 sg13g2_xnor2_1 _3574_ (.Y(_0916_),
    .A(_0851_),
    .B(_0877_));
 sg13g2_xnor2_1 _3575_ (.Y(_0917_),
    .A(_0854_),
    .B(_0874_));
 sg13g2_nand3b_1 _3576_ (.B(_0848_),
    .C(_0856_),
    .Y(_0918_),
    .A_N(_0868_));
 sg13g2_or4_1 _3577_ (.A(_0842_),
    .B(_0844_),
    .C(_0861_),
    .D(_0918_),
    .X(_0919_));
 sg13g2_nor4_1 _3578_ (.A(_0829_),
    .B(_0836_),
    .C(_0838_),
    .D(_0919_),
    .Y(_0920_));
 sg13g2_nor2_1 _3579_ (.A(_0826_),
    .B(_0831_),
    .Y(_0921_));
 sg13g2_nand4_1 _3580_ (.B(_0915_),
    .C(_0920_),
    .A(_0914_),
    .Y(_0922_),
    .D(_0921_));
 sg13g2_xnor2_1 _3581_ (.Y(_0923_),
    .A(_0865_),
    .B(_0867_));
 sg13g2_nand3_1 _3582_ (.B(_0912_),
    .C(_0923_),
    .A(_0822_),
    .Y(_0924_));
 sg13g2_nor4_1 _3583_ (.A(_0911_),
    .B(_0917_),
    .C(_0922_),
    .D(_0924_),
    .Y(_0925_));
 sg13g2_nand3_1 _3584_ (.B(_0916_),
    .C(_0925_),
    .A(_0910_),
    .Y(_0926_));
 sg13g2_nor3_1 _3585_ (.A(_0908_),
    .B(_0909_),
    .C(_0926_),
    .Y(_0927_));
 sg13g2_nor3_1 _3586_ (.A(_0840_),
    .B(_0905_),
    .C(_0906_),
    .Y(_0928_));
 sg13g2_nand4_1 _3587_ (.B(_0907_),
    .C(_0927_),
    .A(_0903_),
    .Y(_0929_),
    .D(_0928_));
 sg13g2_nor4_1 _3588_ (.A(_0901_),
    .B(_0902_),
    .C(_0904_),
    .D(_0929_),
    .Y(_0930_));
 sg13g2_nand2b_2 _3589_ (.Y(_0931_),
    .B(_0930_),
    .A_N(_0900_));
 sg13g2_xor2_1 _3590_ (.B(_0887_),
    .A(_0840_),
    .X(_0932_));
 sg13g2_and2_1 _3591_ (.A(_0676_),
    .B(_0931_),
    .X(_0933_));
 sg13g2_nand2_2 _3592_ (.Y(_0934_),
    .A(_0676_),
    .B(_0931_));
 sg13g2_nand2b_1 _3593_ (.Y(_0935_),
    .B(net722),
    .A_N(net732));
 sg13g2_nor2b_1 _3594_ (.A(net722),
    .B_N(net732),
    .Y(_0936_));
 sg13g2_nand2_1 _3595_ (.Y(_0937_),
    .A(_1929_),
    .B(net723));
 sg13g2_nor2_1 _3596_ (.A(_1929_),
    .B(net723),
    .Y(_0938_));
 sg13g2_nand2_1 _3597_ (.Y(_0939_),
    .A(_1922_),
    .B(net724));
 sg13g2_nor2_1 _3598_ (.A(_1922_),
    .B(net724),
    .Y(_0940_));
 sg13g2_nand2b_1 _3599_ (.Y(_0941_),
    .B(net725),
    .A_N(net737));
 sg13g2_nor2b_1 _3600_ (.A(net725),
    .B_N(net737),
    .Y(_0942_));
 sg13g2_nand2b_1 _3601_ (.Y(_0943_),
    .B(net726),
    .A_N(\reg_a[21] ));
 sg13g2_nor2b_1 _3602_ (.A(net726),
    .B_N(net739),
    .Y(_0944_));
 sg13g2_nand2_1 _3603_ (.Y(_0945_),
    .A(_1930_),
    .B(net727));
 sg13g2_nor2_1 _3604_ (.A(_1930_),
    .B(net727),
    .Y(_0946_));
 sg13g2_nor2_1 _3605_ (.A(_1923_),
    .B(net729),
    .Y(_0947_));
 sg13g2_nand2b_1 _3606_ (.Y(_0948_),
    .B(\reg_a[14] ),
    .A_N(\reg_b[14] ));
 sg13g2_nor2_1 _3607_ (.A(_0702_),
    .B(_0761_),
    .Y(_0949_));
 sg13g2_nor2b_1 _3608_ (.A(net730),
    .B_N(net741),
    .Y(_0950_));
 sg13g2_nand2b_1 _3609_ (.Y(_0951_),
    .B(net742),
    .A_N(\reg_b[12] ));
 sg13g2_nor2_1 _3610_ (.A(_0753_),
    .B(_0951_),
    .Y(_0952_));
 sg13g2_o21ai_1 _3611_ (.B1(_0949_),
    .Y(_0953_),
    .A1(_0950_),
    .A2(_0952_));
 sg13g2_o21ai_1 _3612_ (.B1(_0953_),
    .Y(_0954_),
    .A1(_0761_),
    .A2(_0948_));
 sg13g2_nor4_1 _3613_ (.A(_0702_),
    .B(_0753_),
    .C(_0755_),
    .D(_0761_),
    .Y(_0955_));
 sg13g2_nor2b_1 _3614_ (.A(\reg_b[10] ),
    .B_N(net743),
    .Y(_0956_));
 sg13g2_nand2b_1 _3615_ (.Y(_0957_),
    .B(net744),
    .A_N(\reg_b[8] ));
 sg13g2_nor2b_1 _3616_ (.A(\reg_b[1] ),
    .B_N(net747),
    .Y(_0958_));
 sg13g2_nand2b_1 _3617_ (.Y(_0959_),
    .B(\reg_b[0] ),
    .A_N(\reg_a[0] ));
 sg13g2_a21oi_1 _3618_ (.A1(_0734_),
    .A2(_0959_),
    .Y(_0960_),
    .B1(_0958_));
 sg13g2_o21ai_1 _3619_ (.B1(_0731_),
    .Y(_0961_),
    .A1(_0732_),
    .A2(_0960_));
 sg13g2_a21o_2 _3620_ (.A2(_0961_),
    .A1(_0729_),
    .B1(_0728_),
    .X(_0962_));
 sg13g2_nor2_1 _3621_ (.A(_0715_),
    .B(_0717_),
    .Y(_0963_));
 sg13g2_nor2_1 _3622_ (.A(_0722_),
    .B(_0726_),
    .Y(_0964_));
 sg13g2_and2_1 _3623_ (.A(_0963_),
    .B(_0964_),
    .X(_0965_));
 sg13g2_nand2_1 _3624_ (.Y(_0966_),
    .A(_0963_),
    .B(_0964_));
 sg13g2_a21o_1 _3625_ (.A2(_0724_),
    .A1(_0721_),
    .B1(_0720_),
    .X(_0967_));
 sg13g2_nand2b_1 _3626_ (.Y(_0968_),
    .B(net745),
    .A_N(\reg_b[7] ));
 sg13g2_nand2b_1 _3627_ (.Y(_0969_),
    .B(\reg_a[6] ),
    .A_N(\reg_b[6] ));
 sg13g2_o21ai_1 _3628_ (.B1(_0968_),
    .Y(_0970_),
    .A1(_0715_),
    .A2(_0969_));
 sg13g2_a21oi_1 _3629_ (.A1(_0725_),
    .A2(_0962_),
    .Y(_0971_),
    .B1(_0724_));
 sg13g2_nor2_1 _3630_ (.A(_0722_),
    .B(_0971_),
    .Y(_0972_));
 sg13g2_nor2_1 _3631_ (.A(_0720_),
    .B(_0972_),
    .Y(_0973_));
 sg13g2_o21ai_1 _3632_ (.B1(_0969_),
    .Y(_0974_),
    .A1(_0717_),
    .A2(_0973_));
 sg13g2_a221oi_1 _3633_ (.B2(_0963_),
    .C1(_0970_),
    .B1(_0967_),
    .A1(_0962_),
    .Y(_0975_),
    .A2(_0965_));
 sg13g2_o21ai_1 _3634_ (.B1(_0957_),
    .Y(_0976_),
    .A1(_0712_),
    .A2(_0975_));
 sg13g2_o21ai_1 _3635_ (.B1(_0976_),
    .Y(_0977_),
    .A1(\reg_a[9] ),
    .A2(_1926_));
 sg13g2_o21ai_1 _3636_ (.B1(_0977_),
    .Y(_0978_),
    .A1(_1925_),
    .A2(net731));
 sg13g2_nor2b_1 _3637_ (.A(_0745_),
    .B_N(_0978_),
    .Y(_0979_));
 sg13g2_nor2_1 _3638_ (.A(_0956_),
    .B(_0979_),
    .Y(_0980_));
 sg13g2_nand2_1 _3639_ (.Y(_0981_),
    .A(_0748_),
    .B(_0956_));
 sg13g2_o21ai_1 _3640_ (.B1(_0981_),
    .Y(_0982_),
    .A1(_1931_),
    .A2(\reg_b[11] ));
 sg13g2_nor2_1 _3641_ (.A(_0745_),
    .B(_0749_),
    .Y(_0983_));
 sg13g2_a21oi_1 _3642_ (.A1(_0978_),
    .A2(_0983_),
    .Y(_0984_),
    .B1(_0982_));
 sg13g2_nand2_1 _3643_ (.Y(_0985_),
    .A(_0955_),
    .B(_0983_));
 sg13g2_nor2b_1 _3644_ (.A(_0985_),
    .B_N(_0978_),
    .Y(_0986_));
 sg13g2_a221oi_1 _3645_ (.B2(_0982_),
    .C1(_0954_),
    .B1(_0955_),
    .A1(\reg_a[15] ),
    .Y(_0987_),
    .A2(_1938_));
 sg13g2_inv_1 _3646_ (.Y(_0988_),
    .A(_0987_));
 sg13g2_nor2_1 _3647_ (.A(_0986_),
    .B(_0988_),
    .Y(_0989_));
 sg13g2_o21ai_1 _3648_ (.B1(_0765_),
    .Y(_0990_),
    .A1(_0986_),
    .A2(_0988_));
 sg13g2_nand2b_1 _3649_ (.Y(_0991_),
    .B(\reg_a[16] ),
    .A_N(\reg_b[16] ));
 sg13g2_nand2_1 _3650_ (.Y(_0992_),
    .A(_0990_),
    .B(_0991_));
 sg13g2_a22oi_1 _3651_ (.Y(_0993_),
    .B1(_0990_),
    .B2(_0991_),
    .A2(net729),
    .A1(_1923_));
 sg13g2_nor2_1 _3652_ (.A(_0947_),
    .B(_0993_),
    .Y(_0994_));
 sg13g2_o21ai_1 _3653_ (.B1(_0773_),
    .Y(_0995_),
    .A1(_0947_),
    .A2(_0993_));
 sg13g2_o21ai_1 _3654_ (.B1(_0995_),
    .Y(_0996_),
    .A1(_1927_),
    .A2(net728));
 sg13g2_a21o_1 _3655_ (.A2(_0996_),
    .A1(_0945_),
    .B1(_0946_),
    .X(_0997_));
 sg13g2_nor2_1 _3656_ (.A(_1933_),
    .B(\reg_b[20] ),
    .Y(_0998_));
 sg13g2_a21o_1 _3657_ (.A2(_0997_),
    .A1(_0781_),
    .B1(_0998_),
    .X(_0999_));
 sg13g2_a21o_1 _3658_ (.A2(_0999_),
    .A1(_0943_),
    .B1(_0944_),
    .X(_1000_));
 sg13g2_nor2b_1 _3659_ (.A(\reg_b[22] ),
    .B_N(net738),
    .Y(_1001_));
 sg13g2_a21o_1 _3660_ (.A2(_1000_),
    .A1(_0787_),
    .B1(_1001_),
    .X(_1002_));
 sg13g2_a21oi_1 _3661_ (.A1(_0941_),
    .A2(_1002_),
    .Y(_1003_),
    .B1(_0942_));
 sg13g2_nand2b_1 _3662_ (.Y(_1004_),
    .B(\reg_a[24] ),
    .A_N(\reg_b[24] ));
 sg13g2_o21ai_1 _3663_ (.B1(_1004_),
    .Y(_1005_),
    .A1(_0800_),
    .A2(_1003_));
 sg13g2_a21oi_1 _3664_ (.A1(_0939_),
    .A2(_1005_),
    .Y(_1006_),
    .B1(_0940_));
 sg13g2_nand2b_1 _3665_ (.Y(_1007_),
    .B(net734),
    .A_N(\reg_b[26] ));
 sg13g2_o21ai_1 _3666_ (.B1(_1007_),
    .Y(_1008_),
    .A1(_0811_),
    .A2(_1006_));
 sg13g2_a21oi_1 _3667_ (.A1(_0937_),
    .A2(_1008_),
    .Y(_1009_),
    .B1(_0938_));
 sg13g2_nand2b_1 _3668_ (.Y(_1010_),
    .B(net733),
    .A_N(\reg_b[28] ));
 sg13g2_o21ai_1 _3669_ (.B1(_1010_),
    .Y(_1011_),
    .A1(_0691_),
    .A2(_1009_));
 sg13g2_and2_1 _3670_ (.A(_0935_),
    .B(_1011_),
    .X(_1012_));
 sg13g2_o21ai_1 _3671_ (.B1(_0687_),
    .Y(_1013_),
    .A1(_0936_),
    .A2(_1012_));
 sg13g2_o21ai_1 _3672_ (.B1(_1013_),
    .Y(_1014_),
    .A1(_1935_),
    .A2(\reg_b[30] ));
 sg13g2_xnor2_1 _3673_ (.Y(_1015_),
    .A(_0685_),
    .B(_1014_));
 sg13g2_xnor2_1 _3674_ (.Y(_1016_),
    .A(_0825_),
    .B(_1011_));
 sg13g2_xnor2_1 _3675_ (.Y(_1017_),
    .A(_0690_),
    .B(_1009_));
 sg13g2_xor2_1 _3676_ (.B(_1008_),
    .A(_0814_),
    .X(_1018_));
 sg13g2_xnor2_1 _3677_ (.Y(_1019_),
    .A(_0810_),
    .B(_1006_));
 sg13g2_xor2_1 _3678_ (.B(_1005_),
    .A(_0805_),
    .X(_1020_));
 sg13g2_xnor2_1 _3679_ (.Y(_1021_),
    .A(_0800_),
    .B(_1003_));
 sg13g2_xnor2_1 _3680_ (.Y(_1022_),
    .A(_0790_),
    .B(_1002_));
 sg13g2_xnor2_1 _3681_ (.Y(_1023_),
    .A(_0796_),
    .B(_0999_));
 sg13g2_xnor2_1 _3682_ (.Y(_1024_),
    .A(_0781_),
    .B(_0997_));
 sg13g2_xor2_1 _3683_ (.B(_0996_),
    .A(_0776_),
    .X(_1025_));
 sg13g2_xor2_1 _3684_ (.B(_0994_),
    .A(_0773_),
    .X(_1026_));
 sg13g2_xnor2_1 _3685_ (.Y(_1027_),
    .A(_0769_),
    .B(_0992_));
 sg13g2_xor2_1 _3686_ (.B(_0989_),
    .A(_0765_),
    .X(_1028_));
 sg13g2_or2_1 _3687_ (.X(_1029_),
    .B(_0852_),
    .A(_0712_));
 sg13g2_nor2b_1 _3688_ (.A(_0685_),
    .B_N(_0729_),
    .Y(_1030_));
 sg13g2_nand3b_1 _3689_ (.B(_0734_),
    .C(_1030_),
    .Y(_1031_),
    .A_N(_0732_));
 sg13g2_nor4_1 _3690_ (.A(_0966_),
    .B(_0985_),
    .C(_1029_),
    .D(_1031_),
    .Y(_1032_));
 sg13g2_nand3_1 _3691_ (.B(_1028_),
    .C(_1032_),
    .A(_1027_),
    .Y(_1033_));
 sg13g2_nor2_1 _3692_ (.A(_1025_),
    .B(_1033_),
    .Y(_1034_));
 sg13g2_nand4_1 _3693_ (.B(_1024_),
    .C(_1026_),
    .A(_1023_),
    .Y(_1035_),
    .D(_1034_));
 sg13g2_xnor2_1 _3694_ (.Y(_1036_),
    .A(_0786_),
    .B(_1000_));
 sg13g2_nor3_1 _3695_ (.A(_0687_),
    .B(_0936_),
    .C(_1012_),
    .Y(_1037_));
 sg13g2_or3_1 _3696_ (.A(_1014_),
    .B(_1035_),
    .C(_1036_),
    .X(_1038_));
 sg13g2_nor2_1 _3697_ (.A(_1022_),
    .B(_1038_),
    .Y(_1039_));
 sg13g2_and2_1 _3698_ (.A(_1021_),
    .B(_1039_),
    .X(_1040_));
 sg13g2_nand2_1 _3699_ (.Y(_1041_),
    .A(_1020_),
    .B(_1040_));
 sg13g2_or2_1 _3700_ (.X(_1042_),
    .B(_1041_),
    .A(_1019_));
 sg13g2_nor2_1 _3701_ (.A(_1018_),
    .B(_1042_),
    .Y(_1043_));
 sg13g2_nand2b_1 _3702_ (.Y(_1044_),
    .B(_1043_),
    .A_N(_1017_));
 sg13g2_o21ai_1 _3703_ (.B1(_1013_),
    .Y(_1045_),
    .A1(_1016_),
    .A2(_1044_));
 sg13g2_nor2_1 _3704_ (.A(_1037_),
    .B(_1045_),
    .Y(_1046_));
 sg13g2_nand3b_1 _3705_ (.B(_0734_),
    .C(_0686_),
    .Y(_1047_),
    .A_N(_1014_));
 sg13g2_or2_1 _3706_ (.X(_1048_),
    .B(_1031_),
    .A(_1014_));
 sg13g2_or3_1 _3707_ (.A(_0722_),
    .B(_0726_),
    .C(_1048_),
    .X(_1049_));
 sg13g2_or2_1 _3708_ (.X(_1050_),
    .B(_1048_),
    .A(_0966_));
 sg13g2_nor2_2 _3709_ (.A(_1029_),
    .B(_1050_),
    .Y(_1051_));
 sg13g2_nand2_2 _3710_ (.Y(_1052_),
    .A(_0983_),
    .B(_1051_));
 sg13g2_nor3_1 _3711_ (.A(_0753_),
    .B(_0755_),
    .C(_1052_),
    .Y(_1053_));
 sg13g2_o21ai_1 _3712_ (.B1(_0951_),
    .Y(_1054_),
    .A1(_0755_),
    .A2(_0984_));
 sg13g2_a21oi_1 _3713_ (.A1(_0754_),
    .A2(_1054_),
    .Y(_1055_),
    .B1(_0950_));
 sg13g2_xnor2_1 _3714_ (.Y(_1056_),
    .A(_0702_),
    .B(_1055_));
 sg13g2_nand2_1 _3715_ (.Y(_1057_),
    .A(_1053_),
    .B(_1056_));
 sg13g2_xnor2_1 _3716_ (.Y(_1058_),
    .A(_1053_),
    .B(_1056_));
 sg13g2_nor3_1 _3717_ (.A(_0985_),
    .B(_1029_),
    .C(_1050_),
    .Y(_1059_));
 sg13g2_xnor2_1 _3718_ (.Y(_1060_),
    .A(_1028_),
    .B(_1059_));
 sg13g2_xnor2_1 _3719_ (.Y(_1061_),
    .A(_1016_),
    .B(_1044_));
 sg13g2_xor2_1 _3720_ (.B(_0984_),
    .A(_0755_),
    .X(_1062_));
 sg13g2_xnor2_1 _3721_ (.Y(_1063_),
    .A(_0753_),
    .B(_1054_));
 sg13g2_o21ai_1 _3722_ (.B1(_1063_),
    .Y(_1064_),
    .A1(_1052_),
    .A2(_1062_));
 sg13g2_nand2b_1 _3723_ (.Y(_1065_),
    .B(_1064_),
    .A_N(_1053_));
 sg13g2_xnor2_1 _3724_ (.Y(_1066_),
    .A(_1052_),
    .B(_1062_));
 sg13g2_xor2_1 _3725_ (.B(_1043_),
    .A(_1017_),
    .X(_1067_));
 sg13g2_xor2_1 _3726_ (.B(_0978_),
    .A(_0745_),
    .X(_1068_));
 sg13g2_and2_1 _3727_ (.A(_1051_),
    .B(_1068_),
    .X(_1069_));
 sg13g2_xnor2_1 _3728_ (.Y(_1070_),
    .A(_0749_),
    .B(_0980_));
 sg13g2_o21ai_1 _3729_ (.B1(_1052_),
    .Y(_1071_),
    .A1(_1069_),
    .A2(_1070_));
 sg13g2_xor2_1 _3730_ (.B(_0975_),
    .A(_0712_),
    .X(_1072_));
 sg13g2_xnor2_1 _3731_ (.Y(_1073_),
    .A(_0852_),
    .B(_0976_));
 sg13g2_o21ai_1 _3732_ (.B1(_1073_),
    .Y(_1074_),
    .A1(_1050_),
    .A2(_1072_));
 sg13g2_nor2b_1 _3733_ (.A(_1051_),
    .B_N(_1074_),
    .Y(_1075_));
 sg13g2_inv_1 _3734_ (.Y(_1076_),
    .A(_1075_));
 sg13g2_xnor2_1 _3735_ (.Y(_1077_),
    .A(_1018_),
    .B(_1042_));
 sg13g2_xnor2_1 _3736_ (.Y(_1078_),
    .A(_1051_),
    .B(_1068_));
 sg13g2_xnor2_1 _3737_ (.Y(_1079_),
    .A(_1050_),
    .B(_1072_));
 sg13g2_xnor2_1 _3738_ (.Y(_1080_),
    .A(_1019_),
    .B(_1041_));
 sg13g2_xnor2_1 _3739_ (.Y(_1081_),
    .A(_0718_),
    .B(_0973_));
 sg13g2_xnor2_1 _3740_ (.Y(_1082_),
    .A(_0715_),
    .B(_0974_));
 sg13g2_o21ai_1 _3741_ (.B1(_1082_),
    .Y(_1083_),
    .A1(_1049_),
    .A2(_1081_));
 sg13g2_nand2_1 _3742_ (.Y(_1084_),
    .A(_1050_),
    .B(_1083_));
 sg13g2_or2_1 _3743_ (.X(_1085_),
    .B(_1033_),
    .A(_1014_));
 sg13g2_nand2b_1 _3744_ (.Y(_1086_),
    .B(_1026_),
    .A_N(_1085_));
 sg13g2_nor2_1 _3745_ (.A(_1025_),
    .B(_1086_),
    .Y(_1087_));
 sg13g2_nand3_1 _3746_ (.B(_1024_),
    .C(_1087_),
    .A(_1023_),
    .Y(_1088_));
 sg13g2_nand2_1 _3747_ (.Y(_1089_),
    .A(_1036_),
    .B(_1088_));
 sg13g2_nand2_1 _3748_ (.Y(_1090_),
    .A(_1038_),
    .B(_1089_));
 sg13g2_xnor2_1 _3749_ (.Y(_1091_),
    .A(_1049_),
    .B(_1081_));
 sg13g2_xnor2_1 _3750_ (.Y(_1092_),
    .A(_0726_),
    .B(_0962_));
 sg13g2_xnor2_1 _3751_ (.Y(_1093_),
    .A(_0721_),
    .B(_0971_));
 sg13g2_o21ai_1 _3752_ (.B1(_1093_),
    .Y(_1094_),
    .A1(_1048_),
    .A2(_1092_));
 sg13g2_nand2_1 _3753_ (.Y(_1095_),
    .A(_1049_),
    .B(_1094_));
 sg13g2_xnor2_1 _3754_ (.Y(_1096_),
    .A(_1020_),
    .B(_1040_));
 sg13g2_xor2_1 _3755_ (.B(_0960_),
    .A(_0732_),
    .X(_1097_));
 sg13g2_xor2_1 _3756_ (.B(_0961_),
    .A(_0729_),
    .X(_1098_));
 sg13g2_o21ai_1 _3757_ (.B1(_1098_),
    .Y(_1099_),
    .A1(_1047_),
    .A2(_1097_));
 sg13g2_nand2_1 _3758_ (.Y(_1100_),
    .A(_1048_),
    .B(_1099_));
 sg13g2_xnor2_1 _3759_ (.Y(_1101_),
    .A(_1021_),
    .B(_1039_));
 sg13g2_o21ai_1 _3760_ (.B1(_0959_),
    .Y(_1102_),
    .A1(_0685_),
    .A2(_1014_));
 sg13g2_xnor2_1 _3761_ (.Y(_1103_),
    .A(_0734_),
    .B(_1102_));
 sg13g2_xnor2_1 _3762_ (.Y(_1104_),
    .A(_1048_),
    .B(_1092_));
 sg13g2_xnor2_1 _3763_ (.Y(_1105_),
    .A(_1025_),
    .B(_1086_));
 sg13g2_xnor2_1 _3764_ (.Y(_1106_),
    .A(_1022_),
    .B(_1038_));
 sg13g2_xnor2_1 _3765_ (.Y(_1107_),
    .A(_1047_),
    .B(_1097_));
 sg13g2_xor2_1 _3766_ (.B(_1085_),
    .A(_1026_),
    .X(_1108_));
 sg13g2_a21o_1 _3767_ (.A2(_1087_),
    .A1(_1024_),
    .B1(_1023_),
    .X(_1109_));
 sg13g2_nand2_1 _3768_ (.Y(_1110_),
    .A(_1088_),
    .B(_1109_));
 sg13g2_xnor2_1 _3769_ (.Y(_1111_),
    .A(_1024_),
    .B(_1087_));
 sg13g2_o21ai_1 _3770_ (.B1(_0948_),
    .Y(_1112_),
    .A1(_0702_),
    .A2(_1055_));
 sg13g2_xnor2_1 _3771_ (.Y(_1113_),
    .A(_0761_),
    .B(_1112_));
 sg13g2_a21o_1 _3772_ (.A2(_1113_),
    .A1(_1057_),
    .B1(_1059_),
    .X(_1114_));
 sg13g2_and2_1 _3773_ (.A(_1028_),
    .B(_1059_),
    .X(_1115_));
 sg13g2_o21ai_1 _3774_ (.B1(_1085_),
    .Y(_1116_),
    .A1(_1027_),
    .A2(_1115_));
 sg13g2_and4_1 _3775_ (.A(_1078_),
    .B(_1084_),
    .C(_1096_),
    .D(_1111_),
    .X(_1117_));
 sg13g2_nand3_1 _3776_ (.B(_1090_),
    .C(_1117_),
    .A(_1077_),
    .Y(_1118_));
 sg13g2_nand2_1 _3777_ (.Y(_1119_),
    .A(_1079_),
    .B(_1091_));
 sg13g2_nand2_1 _3778_ (.Y(_1120_),
    .A(_1101_),
    .B(_1105_));
 sg13g2_nand3_1 _3779_ (.B(_1103_),
    .C(_1107_),
    .A(_1095_),
    .Y(_1121_));
 sg13g2_nor3_1 _3780_ (.A(_1119_),
    .B(_1120_),
    .C(_1121_),
    .Y(_1122_));
 sg13g2_and2_1 _3781_ (.A(_1080_),
    .B(_1110_),
    .X(_1123_));
 sg13g2_nand4_1 _3782_ (.B(_1067_),
    .C(_1122_),
    .A(_1066_),
    .Y(_1124_),
    .D(_1123_));
 sg13g2_nand3_1 _3783_ (.B(_1071_),
    .C(_1114_),
    .A(_1060_),
    .Y(_1125_));
 sg13g2_nand2_1 _3784_ (.Y(_1126_),
    .A(_1104_),
    .B(_1108_));
 sg13g2_nand3_1 _3785_ (.B(_1100_),
    .C(_1106_),
    .A(_1015_),
    .Y(_1127_));
 sg13g2_nand2_1 _3786_ (.Y(_1128_),
    .A(_1058_),
    .B(_1065_));
 sg13g2_or4_1 _3787_ (.A(_1075_),
    .B(_1126_),
    .C(_1127_),
    .D(_1128_),
    .X(_1129_));
 sg13g2_nand3b_1 _3788_ (.B(_1116_),
    .C(_1061_),
    .Y(_1130_),
    .A_N(_1129_));
 sg13g2_nor4_1 _3789_ (.A(_1118_),
    .B(_1124_),
    .C(_1125_),
    .D(_1130_),
    .Y(_1131_));
 sg13g2_a21oi_2 _3790_ (.B1(_0675_),
    .Y(_1132_),
    .A2(_1131_),
    .A1(_1046_));
 sg13g2_a221oi_1 _3791_ (.B2(net543),
    .C1(_0681_),
    .B1(_1015_),
    .A1(_0822_),
    .Y(_1133_),
    .A2(net547));
 sg13g2_o21ai_1 _3792_ (.B1(_0669_),
    .Y(_0002_),
    .A1(_0683_),
    .A2(_1133_));
 sg13g2_nor2_1 _3793_ (.A(net715),
    .B(_0360_),
    .Y(_1134_));
 sg13g2_and2_1 _3794_ (.A(net715),
    .B(net551),
    .X(_1135_));
 sg13g2_xor2_1 _3795_ (.B(_0570_),
    .A(_0532_),
    .X(_1136_));
 sg13g2_a21oi_1 _3796_ (.A1(net541),
    .A2(_1136_),
    .Y(_1137_),
    .B1(_1134_));
 sg13g2_xnor2_1 _3797_ (.Y(_1138_),
    .A(_0821_),
    .B(_0861_));
 sg13g2_a22oi_1 _3798_ (.Y(_1139_),
    .B1(_1138_),
    .B2(net547),
    .A2(net543),
    .A1(_1103_));
 sg13g2_nand2_1 _3799_ (.Y(_1140_),
    .A(net747),
    .B(net570));
 sg13g2_o21ai_1 _3800_ (.B1(_1140_),
    .Y(_1141_),
    .A1(_1925_),
    .A2(net570));
 sg13g2_o21ai_1 _3801_ (.B1(net654),
    .Y(_1142_),
    .A1(net630),
    .A2(_1141_));
 sg13g2_a21oi_1 _3802_ (.A1(net630),
    .A2(_1139_),
    .Y(_1143_),
    .B1(_1142_));
 sg13g2_nand2_1 _3803_ (.Y(_1144_),
    .A(net688),
    .B(_1141_));
 sg13g2_o21ai_1 _3804_ (.B1(_1144_),
    .Y(_1145_),
    .A1(net636),
    .A2(_1137_));
 sg13g2_or2_1 _3805_ (.X(_0013_),
    .B(_1145_),
    .A(_1143_));
 sg13g2_a21oi_1 _3806_ (.A1(_0645_),
    .A2(net551),
    .Y(_1146_),
    .B1(net700));
 sg13g2_o21ai_1 _3807_ (.B1(net639),
    .Y(_1147_),
    .A1(net716),
    .A2(_0367_));
 sg13g2_mux2_1 _3808_ (.A0(net746),
    .A1(net743),
    .S(net574),
    .X(_1148_));
 sg13g2_a22oi_1 _3809_ (.Y(_1149_),
    .B1(_1107_),
    .B2(net543),
    .A2(net547),
    .A1(_0915_));
 sg13g2_nand2_1 _3810_ (.Y(_1150_),
    .A(net630),
    .B(_1149_));
 sg13g2_nor2_1 _3811_ (.A(net630),
    .B(_1148_),
    .Y(_1151_));
 sg13g2_nor2_1 _3812_ (.A(net634),
    .B(_1151_),
    .Y(_1152_));
 sg13g2_a22oi_1 _3813_ (.Y(_1153_),
    .B1(_1150_),
    .B2(_1152_),
    .A2(_1148_),
    .A1(net678));
 sg13g2_o21ai_1 _3814_ (.B1(_1153_),
    .Y(_0024_),
    .A1(_1146_),
    .A2(_1147_));
 sg13g2_mux2_1 _3815_ (.A0(_1928_),
    .A1(_1931_),
    .S(net574),
    .X(_1154_));
 sg13g2_o21ai_1 _3816_ (.B1(net715),
    .Y(_1155_),
    .A1(_0651_),
    .A2(_0664_));
 sg13g2_nand2_1 _3817_ (.Y(_1156_),
    .A(net700),
    .B(_0371_));
 sg13g2_nand3_1 _3818_ (.B(_1155_),
    .C(_1156_),
    .A(net704),
    .Y(_1157_));
 sg13g2_nand2_1 _3819_ (.Y(_1158_),
    .A(_0923_),
    .B(net547));
 sg13g2_a21oi_1 _3820_ (.A1(_1100_),
    .A2(net543),
    .Y(_1159_),
    .B1(net626));
 sg13g2_a221oi_1 _3821_ (.B2(_1159_),
    .C1(net704),
    .B1(_1158_),
    .A1(net626),
    .Y(_1160_),
    .A2(_1154_));
 sg13g2_nor2_1 _3822_ (.A(net685),
    .B(_1160_),
    .Y(_1161_));
 sg13g2_a22oi_1 _3823_ (.Y(_0027_),
    .B1(_1157_),
    .B2(_1161_),
    .A2(net386),
    .A1(net685));
 sg13g2_xnor2_1 _3824_ (.Y(_1162_),
    .A(_0573_),
    .B(_0580_));
 sg13g2_a221oi_1 _3825_ (.B2(_1162_),
    .C1(net635),
    .B1(net541),
    .A1(net700),
    .Y(_1163_),
    .A2(_0387_));
 sg13g2_nand2_1 _3826_ (.Y(_1164_),
    .A(net742),
    .B(net574));
 sg13g2_o21ai_1 _3827_ (.B1(_1164_),
    .Y(_1165_),
    .A1(_1932_),
    .A2(net574));
 sg13g2_nor2_1 _3828_ (.A(net630),
    .B(_1165_),
    .Y(_1166_));
 sg13g2_a221oi_1 _3829_ (.B2(net543),
    .C1(net626),
    .B1(_1104_),
    .A1(_0914_),
    .Y(_1167_),
    .A2(net547));
 sg13g2_o21ai_1 _3830_ (.B1(net654),
    .Y(_1168_),
    .A1(_1166_),
    .A2(_1167_));
 sg13g2_o21ai_1 _3831_ (.B1(_1168_),
    .Y(_1169_),
    .A1(net695),
    .A2(_1165_));
 sg13g2_nor2_1 _3832_ (.A(_1163_),
    .B(_1169_),
    .Y(_0028_));
 sg13g2_o21ai_1 _3833_ (.B1(net715),
    .Y(_1170_),
    .A1(_0634_),
    .A2(_0664_));
 sg13g2_a21oi_1 _3834_ (.A1(_0327_),
    .A2(net555),
    .Y(_1171_),
    .B1(net715));
 sg13g2_nand2_1 _3835_ (.Y(_1172_),
    .A(net639),
    .B(_1170_));
 sg13g2_nand2_1 _3836_ (.Y(_1173_),
    .A(_0868_),
    .B(_0913_));
 sg13g2_nand3_1 _3837_ (.B(net547),
    .C(_1173_),
    .A(_0871_),
    .Y(_1174_));
 sg13g2_a21oi_1 _3838_ (.A1(_1095_),
    .A2(net543),
    .Y(_1175_),
    .B1(net626));
 sg13g2_and2_1 _3839_ (.A(net741),
    .B(net574),
    .X(_1176_));
 sg13g2_a21oi_1 _3840_ (.A1(\reg_a[5] ),
    .A2(net570),
    .Y(_1177_),
    .B1(_1176_));
 sg13g2_a221oi_1 _3841_ (.B2(net626),
    .C1(net634),
    .B1(_1177_),
    .A1(_1174_),
    .Y(_1178_),
    .A2(_1175_));
 sg13g2_nor2_1 _3842_ (.A(net695),
    .B(_1177_),
    .Y(_1179_));
 sg13g2_nor2_1 _3843_ (.A(_1178_),
    .B(_1179_),
    .Y(_1180_));
 sg13g2_o21ai_1 _3844_ (.B1(_1180_),
    .Y(_0029_),
    .A1(_1171_),
    .A2(_1172_));
 sg13g2_a21o_1 _3845_ (.A2(net551),
    .A1(_0644_),
    .B1(net700),
    .X(_1181_));
 sg13g2_a21oi_1 _3846_ (.A1(net701),
    .A2(_0381_),
    .Y(_1182_),
    .B1(net635));
 sg13g2_a221oi_1 _3847_ (.B2(net543),
    .C1(net626),
    .B1(_1091_),
    .A1(_0912_),
    .Y(_1183_),
    .A2(net547));
 sg13g2_nand2_1 _3848_ (.Y(_1184_),
    .A(net388),
    .B(net574));
 sg13g2_o21ai_1 _3849_ (.B1(_1184_),
    .Y(_1185_),
    .A1(_1934_),
    .A2(net574));
 sg13g2_o21ai_1 _3850_ (.B1(net654),
    .Y(_1186_),
    .A1(net630),
    .A2(_1185_));
 sg13g2_a22oi_1 _3851_ (.Y(_1187_),
    .B1(_1185_),
    .B2(net678),
    .A2(_1182_),
    .A1(_1181_));
 sg13g2_o21ai_1 _3852_ (.B1(_1187_),
    .Y(_0030_),
    .A1(_1183_),
    .A2(_1186_));
 sg13g2_nand2b_1 _3853_ (.Y(_1188_),
    .B(_0643_),
    .A_N(_0578_));
 sg13g2_nand3_1 _3854_ (.B(net551),
    .C(_1188_),
    .A(_0585_),
    .Y(_1189_));
 sg13g2_nand2_1 _3855_ (.Y(_1190_),
    .A(net716),
    .B(_1189_));
 sg13g2_a21oi_1 _3856_ (.A1(net701),
    .A2(_0375_),
    .Y(_1191_),
    .B1(net635));
 sg13g2_xnor2_1 _3857_ (.Y(_1192_),
    .A(_0857_),
    .B(_0872_));
 sg13g2_a221oi_1 _3858_ (.B2(net547),
    .C1(net626),
    .B1(_1192_),
    .A1(_1084_),
    .Y(_1193_),
    .A2(net543));
 sg13g2_nand2_1 _3859_ (.Y(_1194_),
    .A(net745),
    .B(net570));
 sg13g2_o21ai_1 _3860_ (.B1(_1194_),
    .Y(_1195_),
    .A1(_1937_),
    .A2(net570));
 sg13g2_o21ai_1 _3861_ (.B1(net654),
    .Y(_1196_),
    .A1(net630),
    .A2(_1195_));
 sg13g2_a22oi_1 _3862_ (.Y(_1197_),
    .B1(_1195_),
    .B2(net678),
    .A2(_1191_),
    .A1(_1190_));
 sg13g2_o21ai_1 _3863_ (.B1(_1197_),
    .Y(_0031_),
    .A1(_1193_),
    .A2(_1196_));
 sg13g2_a221oi_1 _3864_ (.B2(net541),
    .C1(net635),
    .B1(_0636_),
    .A1(net700),
    .Y(_1198_),
    .A2(_0413_));
 sg13g2_mux2_1 _3865_ (.A0(net740),
    .A1(net744),
    .S(net570),
    .X(_1199_));
 sg13g2_inv_1 _3866_ (.Y(_1200_),
    .A(_1199_));
 sg13g2_nor2_1 _3867_ (.A(net695),
    .B(_1199_),
    .Y(_1201_));
 sg13g2_nand2b_1 _3868_ (.Y(_1202_),
    .B(net548),
    .A_N(_0911_));
 sg13g2_a21oi_1 _3869_ (.A1(_1079_),
    .A2(net544),
    .Y(_1203_),
    .B1(net627));
 sg13g2_a22oi_1 _3870_ (.Y(_1204_),
    .B1(_1202_),
    .B2(_1203_),
    .A2(_1200_),
    .A1(net626));
 sg13g2_nor2_1 _3871_ (.A(net634),
    .B(_1204_),
    .Y(_1205_));
 sg13g2_nor3_1 _3872_ (.A(_1198_),
    .B(_1201_),
    .C(_1205_),
    .Y(_0032_));
 sg13g2_xor2_1 _3873_ (.B(_0635_),
    .A(_0600_),
    .X(_1206_));
 sg13g2_a22oi_1 _3874_ (.Y(_1207_),
    .B1(net541),
    .B2(_1206_),
    .A2(_0404_),
    .A1(net700));
 sg13g2_nand2_1 _3875_ (.Y(_1208_),
    .A(\reg_a[17] ),
    .B(net575));
 sg13g2_o21ai_1 _3876_ (.B1(_1208_),
    .Y(_1209_),
    .A1(_1925_),
    .A2(net575));
 sg13g2_a21oi_1 _3877_ (.A1(_1076_),
    .A2(net544),
    .Y(_1210_),
    .B1(net627));
 sg13g2_o21ai_1 _3878_ (.B1(_1210_),
    .Y(_1211_),
    .A1(_0917_),
    .A2(_0934_));
 sg13g2_nor2_1 _3879_ (.A(net630),
    .B(_1209_),
    .Y(_1212_));
 sg13g2_nor2_1 _3880_ (.A(net634),
    .B(_1212_),
    .Y(_1213_));
 sg13g2_a22oi_1 _3881_ (.Y(_1214_),
    .B1(_1211_),
    .B2(_1213_),
    .A2(_1209_),
    .A1(net688));
 sg13g2_o21ai_1 _3882_ (.B1(_1214_),
    .Y(_0033_),
    .A1(net635),
    .A2(_1207_));
 sg13g2_o21ai_1 _3883_ (.B1(net715),
    .Y(_1215_),
    .A1(_0641_),
    .A2(_0664_));
 sg13g2_a21oi_1 _3884_ (.A1(_0320_),
    .A2(net557),
    .Y(_1216_),
    .B1(net716));
 sg13g2_nand2_1 _3885_ (.Y(_1217_),
    .A(net639),
    .B(_1215_));
 sg13g2_nand2_1 _3886_ (.Y(_1218_),
    .A(net743),
    .B(net570));
 sg13g2_o21ai_1 _3887_ (.B1(_1218_),
    .Y(_1219_),
    .A1(_1927_),
    .A2(net573));
 sg13g2_a22oi_1 _3888_ (.Y(_1220_),
    .B1(_1078_),
    .B2(net544),
    .A2(net548),
    .A1(_0910_));
 sg13g2_nand2_1 _3889_ (.Y(_1221_),
    .A(net631),
    .B(_1220_));
 sg13g2_nor2_1 _3890_ (.A(net631),
    .B(_1219_),
    .Y(_1222_));
 sg13g2_nor2_1 _3891_ (.A(net634),
    .B(_1222_),
    .Y(_1223_));
 sg13g2_a22oi_1 _3892_ (.Y(_1224_),
    .B1(_1221_),
    .B2(_1223_),
    .A2(_1219_),
    .A1(net678));
 sg13g2_o21ai_1 _3893_ (.B1(_1224_),
    .Y(_0003_),
    .A1(_1216_),
    .A2(_1217_));
 sg13g2_xnor2_1 _3894_ (.Y(_1225_),
    .A(_0603_),
    .B(_0640_));
 sg13g2_o21ai_1 _3895_ (.B1(net715),
    .Y(_1226_),
    .A1(_0664_),
    .A2(_1225_));
 sg13g2_a21oi_1 _3896_ (.A1(net700),
    .A2(_0399_),
    .Y(_1227_),
    .B1(net635));
 sg13g2_nand2_1 _3897_ (.Y(_1228_),
    .A(\reg_a[19] ),
    .B(net575));
 sg13g2_o21ai_1 _3898_ (.B1(_1228_),
    .Y(_1229_),
    .A1(_1931_),
    .A2(net575));
 sg13g2_nand2_1 _3899_ (.Y(_1230_),
    .A(net678),
    .B(_1229_));
 sg13g2_a221oi_1 _3900_ (.B2(net544),
    .C1(net629),
    .B1(_1071_),
    .A1(_0916_),
    .Y(_1231_),
    .A2(net548));
 sg13g2_o21ai_1 _3901_ (.B1(net654),
    .Y(_1232_),
    .A1(net631),
    .A2(_1229_));
 sg13g2_o21ai_1 _3902_ (.B1(_1230_),
    .Y(_1233_),
    .A1(_1231_),
    .A2(_1232_));
 sg13g2_a21oi_1 _3903_ (.A1(_1226_),
    .A2(_1227_),
    .Y(_1234_),
    .B1(_1233_));
 sg13g2_inv_1 _3904_ (.Y(_0004_),
    .A(_1234_));
 sg13g2_nor2_1 _3905_ (.A(_1933_),
    .B(net571),
    .Y(_1235_));
 sg13g2_a21oi_1 _3906_ (.A1(net742),
    .A2(net570),
    .Y(_1236_),
    .B1(_1235_));
 sg13g2_nand2b_1 _3907_ (.Y(_1237_),
    .B(net551),
    .A_N(_0638_));
 sg13g2_o21ai_1 _3908_ (.B1(net704),
    .Y(_1238_),
    .A1(net716),
    .A2(_0427_));
 sg13g2_a21oi_1 _3909_ (.A1(net716),
    .A2(_1237_),
    .Y(_1239_),
    .B1(_1238_));
 sg13g2_nand2b_1 _3910_ (.Y(_1240_),
    .B(net548),
    .A_N(_0909_));
 sg13g2_a21oi_1 _3911_ (.A1(_1066_),
    .A2(net544),
    .Y(_1241_),
    .B1(net627));
 sg13g2_a221oi_1 _3912_ (.B2(_1241_),
    .C1(net704),
    .B1(_1240_),
    .A1(net627),
    .Y(_1242_),
    .A2(_1236_));
 sg13g2_nor3_1 _3913_ (.A(net678),
    .B(_1239_),
    .C(_1242_),
    .Y(_1243_));
 sg13g2_a21oi_1 _3914_ (.A1(net679),
    .A2(_1236_),
    .Y(_0005_),
    .B1(_1243_));
 sg13g2_nand3_1 _3915_ (.B(net557),
    .C(_0430_),
    .A(net701),
    .Y(_1244_));
 sg13g2_xnor2_1 _3916_ (.Y(_1245_),
    .A(_0607_),
    .B(_0628_));
 sg13g2_nand2_1 _3917_ (.Y(_1246_),
    .A(net541),
    .B(_1245_));
 sg13g2_a21oi_1 _3918_ (.A1(_1244_),
    .A2(_1246_),
    .Y(_1247_),
    .B1(net636));
 sg13g2_nor2b_1 _3919_ (.A(_0881_),
    .B_N(_0931_),
    .Y(_1248_));
 sg13g2_xnor2_1 _3920_ (.Y(_1249_),
    .A(_0848_),
    .B(_1248_));
 sg13g2_a221oi_1 _3921_ (.B2(_0676_),
    .C1(net627),
    .B1(_1249_),
    .A1(_1065_),
    .Y(_1250_),
    .A2(net544));
 sg13g2_mux2_1 _3922_ (.A0(net739),
    .A1(net741),
    .S(net573),
    .X(_1251_));
 sg13g2_o21ai_1 _3923_ (.B1(net654),
    .Y(_1252_),
    .A1(net631),
    .A2(_1251_));
 sg13g2_nand2_1 _3924_ (.Y(_1253_),
    .A(net683),
    .B(_1251_));
 sg13g2_o21ai_1 _3925_ (.B1(_1253_),
    .Y(_1254_),
    .A1(_1250_),
    .A2(_1252_));
 sg13g2_or2_1 _3926_ (.X(_0006_),
    .B(_1254_),
    .A(_1247_));
 sg13g2_a22oi_1 _3927_ (.Y(_1255_),
    .B1(_0631_),
    .B2(net541),
    .A2(_0423_),
    .A1(net701));
 sg13g2_a21oi_1 _3928_ (.A1(_1058_),
    .A2(net544),
    .Y(_1256_),
    .B1(net627));
 sg13g2_o21ai_1 _3929_ (.B1(_1256_),
    .Y(_1257_),
    .A1(_0908_),
    .A2(_0934_));
 sg13g2_nand2_1 _3930_ (.Y(_1258_),
    .A(net738),
    .B(net576));
 sg13g2_o21ai_1 _3931_ (.B1(_1258_),
    .Y(_1259_),
    .A1(_1936_),
    .A2(net575));
 sg13g2_nor2_1 _3932_ (.A(net631),
    .B(_1259_),
    .Y(_1260_));
 sg13g2_nor2_1 _3933_ (.A(net634),
    .B(_1260_),
    .Y(_1261_));
 sg13g2_nand2_1 _3934_ (.Y(_1262_),
    .A(net678),
    .B(_1259_));
 sg13g2_o21ai_1 _3935_ (.B1(_1262_),
    .Y(_1263_),
    .A1(net636),
    .A2(_1255_));
 sg13g2_a21o_1 _3936_ (.A2(_1261_),
    .A1(_1257_),
    .B1(_1263_),
    .X(_0007_));
 sg13g2_o21ai_1 _3937_ (.B1(_0609_),
    .Y(_1264_),
    .A1(_0592_),
    .A2(_0630_));
 sg13g2_inv_1 _3938_ (.Y(_1265_),
    .A(_1264_));
 sg13g2_a22oi_1 _3939_ (.Y(_1266_),
    .B1(net541),
    .B2(_1265_),
    .A2(_0418_),
    .A1(net701));
 sg13g2_nand2_1 _3940_ (.Y(_1267_),
    .A(net736),
    .B(net576));
 sg13g2_o21ai_1 _3941_ (.B1(_1267_),
    .Y(_1268_),
    .A1(_1937_),
    .A2(net575));
 sg13g2_xor2_1 _3942_ (.B(_0883_),
    .A(_0844_),
    .X(_1269_));
 sg13g2_a22oi_1 _3943_ (.Y(_1270_),
    .B1(_1269_),
    .B2(net548),
    .A2(_1132_),
    .A1(_1114_));
 sg13g2_o21ai_1 _3944_ (.B1(net654),
    .Y(_1271_),
    .A1(net631),
    .A2(_1268_));
 sg13g2_a21oi_1 _3945_ (.A1(net631),
    .A2(_1270_),
    .Y(_1272_),
    .B1(_1271_));
 sg13g2_a21oi_1 _3946_ (.A1(net678),
    .A2(_1268_),
    .Y(_1273_),
    .B1(_1272_));
 sg13g2_o21ai_1 _3947_ (.B1(_1273_),
    .Y(_0008_),
    .A1(net635),
    .A2(_1266_));
 sg13g2_a21oi_1 _3948_ (.A1(_0637_),
    .A2(net552),
    .Y(_1274_),
    .B1(net703));
 sg13g2_o21ai_1 _3949_ (.B1(net639),
    .Y(_1275_),
    .A1(net717),
    .A2(_0476_));
 sg13g2_nor2_1 _3950_ (.A(_1274_),
    .B(_1275_),
    .Y(_1276_));
 sg13g2_mux2_1 _3951_ (.A0(net735),
    .A1(net740),
    .S(net571),
    .X(_1277_));
 sg13g2_nand2_1 _3952_ (.Y(_1278_),
    .A(net683),
    .B(_1277_));
 sg13g2_a221oi_1 _3953_ (.B2(net546),
    .C1(net628),
    .B1(_1060_),
    .A1(_0907_),
    .Y(_1279_),
    .A2(net549));
 sg13g2_o21ai_1 _3954_ (.B1(net653),
    .Y(_1280_),
    .A1(net633),
    .A2(_1277_));
 sg13g2_o21ai_1 _3955_ (.B1(_1278_),
    .Y(_1281_),
    .A1(_1279_),
    .A2(_1280_));
 sg13g2_or2_1 _3956_ (.X(_0009_),
    .B(_1281_),
    .A(_1276_));
 sg13g2_nor3_1 _3957_ (.A(_0565_),
    .B(_0609_),
    .C(_0611_),
    .Y(_1282_));
 sg13g2_xnor2_1 _3958_ (.Y(_1283_),
    .A(_0565_),
    .B(_0612_));
 sg13g2_a21oi_1 _3959_ (.A1(net552),
    .A2(_1283_),
    .Y(_1284_),
    .B1(net703));
 sg13g2_o21ai_1 _3960_ (.B1(net639),
    .Y(_1285_),
    .A1(net717),
    .A2(_0473_));
 sg13g2_xor2_1 _3961_ (.B(_0885_),
    .A(_0842_),
    .X(_1286_));
 sg13g2_a21oi_1 _3962_ (.A1(_1116_),
    .A2(net546),
    .Y(_1287_),
    .B1(_0681_));
 sg13g2_o21ai_1 _3963_ (.B1(_1287_),
    .Y(_1288_),
    .A1(_0934_),
    .A2(_1286_));
 sg13g2_a21oi_1 _3964_ (.A1(net379),
    .A2(net577),
    .Y(_1289_),
    .B1(_0680_));
 sg13g2_o21ai_1 _3965_ (.B1(_1289_),
    .Y(_1290_),
    .A1(_1923_),
    .A2(net576));
 sg13g2_nand3_1 _3966_ (.B(_1288_),
    .C(net380),
    .A(net637),
    .Y(_1291_));
 sg13g2_o21ai_1 _3967_ (.B1(_1291_),
    .Y(_0010_),
    .A1(_1284_),
    .A2(_1285_));
 sg13g2_nor2_1 _3968_ (.A(_1927_),
    .B(net576),
    .Y(_1292_));
 sg13g2_a21oi_1 _3969_ (.A1(net734),
    .A2(net576),
    .Y(_1293_),
    .B1(_1292_));
 sg13g2_nor2_1 _3970_ (.A(net717),
    .B(_0468_),
    .Y(_1294_));
 sg13g2_xnor2_1 _3971_ (.Y(_1295_),
    .A(_0564_),
    .B(_1282_));
 sg13g2_a21oi_1 _3972_ (.A1(net541),
    .A2(_1295_),
    .Y(_1296_),
    .B1(_1294_));
 sg13g2_nand2b_1 _3973_ (.Y(_1297_),
    .B(net705),
    .A_N(_1296_));
 sg13g2_nand2_1 _3974_ (.Y(_1298_),
    .A(_1108_),
    .B(net546));
 sg13g2_o21ai_1 _3975_ (.B1(_1298_),
    .Y(_1299_),
    .A1(_0906_),
    .A2(_0934_));
 sg13g2_nor3_1 _3976_ (.A(_0666_),
    .B(_0680_),
    .C(_1293_),
    .Y(_1300_));
 sg13g2_a21oi_1 _3977_ (.A1(_2086_),
    .A2(_1299_),
    .Y(_1301_),
    .B1(_1300_));
 sg13g2_a22oi_1 _3978_ (.Y(_0011_),
    .B1(_1297_),
    .B2(_1301_),
    .A2(net372),
    .A1(net683));
 sg13g2_nand2_1 _3979_ (.Y(_1302_),
    .A(net382),
    .B(net577));
 sg13g2_o21ai_1 _3980_ (.B1(_1302_),
    .Y(_1303_),
    .A1(_1930_),
    .A2(net576));
 sg13g2_nor2_1 _3981_ (.A(net696),
    .B(net383),
    .Y(_1304_));
 sg13g2_a21o_1 _3982_ (.A2(_0612_),
    .A1(_0566_),
    .B1(_0563_),
    .X(_1305_));
 sg13g2_nand3_1 _3983_ (.B(net552),
    .C(_1305_),
    .A(_0614_),
    .Y(_1306_));
 sg13g2_nand2_1 _3984_ (.Y(_1307_),
    .A(net703),
    .B(_0464_));
 sg13g2_nand2_1 _3985_ (.Y(_1308_),
    .A(net705),
    .B(_1307_));
 sg13g2_a21oi_1 _3986_ (.A1(net717),
    .A2(_1306_),
    .Y(_1309_),
    .B1(_1308_));
 sg13g2_a221oi_1 _3987_ (.B2(net546),
    .C1(net628),
    .B1(_1105_),
    .A1(_0932_),
    .Y(_1310_),
    .A2(net549));
 sg13g2_nor2_1 _3988_ (.A(net633),
    .B(_1303_),
    .Y(_1311_));
 sg13g2_nor3_1 _3989_ (.A(net704),
    .B(_1310_),
    .C(_1311_),
    .Y(_1312_));
 sg13g2_nor3_1 _3990_ (.A(net683),
    .B(_1309_),
    .C(_1312_),
    .Y(_1313_));
 sg13g2_nor2_1 _3991_ (.A(_1304_),
    .B(_1313_),
    .Y(_0012_));
 sg13g2_nor2_1 _3992_ (.A(net717),
    .B(_0457_),
    .Y(_1314_));
 sg13g2_a21oi_1 _3993_ (.A1(_0626_),
    .A2(net542),
    .Y(_1315_),
    .B1(_1314_));
 sg13g2_nand2_1 _3994_ (.Y(_1316_),
    .A(net733),
    .B(net577));
 sg13g2_o21ai_1 _3995_ (.B1(_1316_),
    .Y(_1317_),
    .A1(_1933_),
    .A2(net577));
 sg13g2_a21oi_1 _3996_ (.A1(_1111_),
    .A2(net546),
    .Y(_1318_),
    .B1(net628));
 sg13g2_o21ai_1 _3997_ (.B1(_1318_),
    .Y(_1319_),
    .A1(_0905_),
    .A2(_0934_));
 sg13g2_nor2_1 _3998_ (.A(net633),
    .B(_1317_),
    .Y(_1320_));
 sg13g2_nor2_1 _3999_ (.A(net634),
    .B(_1320_),
    .Y(_1321_));
 sg13g2_a22oi_1 _4000_ (.Y(_1322_),
    .B1(_1319_),
    .B2(_1321_),
    .A2(_1317_),
    .A1(net683));
 sg13g2_o21ai_1 _4001_ (.B1(_1322_),
    .Y(_0014_),
    .A1(net638),
    .A2(_1315_));
 sg13g2_o21ai_1 _4002_ (.B1(_0557_),
    .Y(_1323_),
    .A1(_0555_),
    .A2(_0614_));
 sg13g2_nand2_1 _4003_ (.Y(_1324_),
    .A(net552),
    .B(_1323_));
 sg13g2_o21ai_1 _4004_ (.B1(net718),
    .Y(_1325_),
    .A1(_0615_),
    .A2(_1324_));
 sg13g2_o21ai_1 _4005_ (.B1(_1325_),
    .Y(_1326_),
    .A1(net718),
    .A2(_0455_));
 sg13g2_mux2_1 _4006_ (.A0(net732),
    .A1(net739),
    .S(net571),
    .X(_1327_));
 sg13g2_xnor2_1 _4007_ (.Y(_1328_),
    .A(_0839_),
    .B(_0890_));
 sg13g2_a221oi_1 _4008_ (.B2(net549),
    .C1(net629),
    .B1(_1328_),
    .A1(_1110_),
    .Y(_1329_),
    .A2(net545));
 sg13g2_nor2_1 _4009_ (.A(net632),
    .B(_1327_),
    .Y(_1330_));
 sg13g2_nor2_1 _4010_ (.A(_1329_),
    .B(_1330_),
    .Y(_1331_));
 sg13g2_a22oi_1 _4011_ (.Y(_1332_),
    .B1(_1331_),
    .B2(net652),
    .A2(_1327_),
    .A1(net683));
 sg13g2_o21ai_1 _4012_ (.B1(_1332_),
    .Y(_0015_),
    .A1(net637),
    .A2(_1326_));
 sg13g2_xnor2_1 _4013_ (.Y(_1333_),
    .A(_0554_),
    .B(_0615_));
 sg13g2_a22oi_1 _4014_ (.Y(_1334_),
    .B1(net542),
    .B2(_1333_),
    .A2(_0451_),
    .A1(net702));
 sg13g2_nand2_1 _4015_ (.Y(_1335_),
    .A(net738),
    .B(net571));
 sg13g2_o21ai_1 _4016_ (.B1(_1335_),
    .Y(_1336_),
    .A1(_1935_),
    .A2(net571));
 sg13g2_nand2b_1 _4017_ (.Y(_1337_),
    .B(net549),
    .A_N(_0904_));
 sg13g2_a21oi_1 _4018_ (.A1(_1090_),
    .A2(net545),
    .Y(_1338_),
    .B1(net629));
 sg13g2_o21ai_1 _4019_ (.B1(net653),
    .Y(_1339_),
    .A1(net632),
    .A2(_1336_));
 sg13g2_a21oi_1 _4020_ (.A1(_1337_),
    .A2(_1338_),
    .Y(_1340_),
    .B1(_1339_));
 sg13g2_a21oi_1 _4021_ (.A1(net683),
    .A2(_1336_),
    .Y(_1341_),
    .B1(_1340_));
 sg13g2_o21ai_1 _4022_ (.B1(_1341_),
    .Y(_0016_),
    .A1(net637),
    .A2(_1334_));
 sg13g2_a21oi_1 _4023_ (.A1(_0625_),
    .A2(net552),
    .Y(_1342_),
    .B1(net702));
 sg13g2_a21oi_1 _4024_ (.A1(_0315_),
    .A2(net559),
    .Y(_1343_),
    .B1(net718));
 sg13g2_or3_1 _4025_ (.A(net637),
    .B(_1342_),
    .C(_1343_),
    .X(_1344_));
 sg13g2_xor2_1 _4026_ (.B(_0892_),
    .A(_0836_),
    .X(_1345_));
 sg13g2_a221oi_1 _4027_ (.B2(net550),
    .C1(_0681_),
    .B1(_1345_),
    .A1(_1106_),
    .Y(_1346_),
    .A2(net545));
 sg13g2_mux2_1 _4028_ (.A0(net237),
    .A1(net737),
    .S(net572),
    .X(_1347_));
 sg13g2_o21ai_1 _4029_ (.B1(net638),
    .Y(_1348_),
    .A1(_0680_),
    .A2(_1347_));
 sg13g2_o21ai_1 _4030_ (.B1(_1344_),
    .Y(_0017_),
    .A1(_1346_),
    .A2(_1348_));
 sg13g2_nor2b_1 _4031_ (.A(_0642_),
    .B_N(net542),
    .Y(_1349_));
 sg13g2_a21oi_1 _4032_ (.A1(net702),
    .A2(_0507_),
    .Y(_1350_),
    .B1(_1349_));
 sg13g2_a22oi_1 _4033_ (.Y(_1351_),
    .B1(_1101_),
    .B2(net545),
    .A2(net549),
    .A1(_0903_));
 sg13g2_nor2_1 _4034_ (.A(net735),
    .B(net578),
    .Y(_1352_));
 sg13g2_a21oi_1 _4035_ (.A1(_1962_),
    .A2(net578),
    .Y(_1353_),
    .B1(_1352_));
 sg13g2_o21ai_1 _4036_ (.B1(net652),
    .Y(_1354_),
    .A1(net632),
    .A2(_1353_));
 sg13g2_a21oi_1 _4037_ (.A1(net632),
    .A2(_1351_),
    .Y(_1355_),
    .B1(_1354_));
 sg13g2_a21oi_1 _4038_ (.A1(net692),
    .A2(_1353_),
    .Y(_1356_),
    .B1(_1355_));
 sg13g2_o21ai_1 _4039_ (.B1(_1356_),
    .Y(_0018_),
    .A1(net637),
    .A2(_1350_));
 sg13g2_a21o_1 _4040_ (.A2(_0617_),
    .A1(_0545_),
    .B1(_0546_),
    .X(_1357_));
 sg13g2_nand2_1 _4041_ (.Y(_1358_),
    .A(net551),
    .B(_1357_));
 sg13g2_o21ai_1 _4042_ (.B1(net717),
    .Y(_1359_),
    .A1(_0618_),
    .A2(_1358_));
 sg13g2_a21oi_1 _4043_ (.A1(net702),
    .A2(_0503_),
    .Y(_1360_),
    .B1(net637));
 sg13g2_xnor2_1 _4044_ (.Y(_1361_),
    .A(_0831_),
    .B(_0894_));
 sg13g2_a221oi_1 _4045_ (.B2(net549),
    .C1(net628),
    .B1(_1361_),
    .A1(_1096_),
    .Y(_1362_),
    .A2(net545));
 sg13g2_nor2_1 _4046_ (.A(net2),
    .B(net571),
    .Y(_1363_));
 sg13g2_a21oi_1 _4047_ (.A1(_1922_),
    .A2(net572),
    .Y(_1364_),
    .B1(_1363_));
 sg13g2_o21ai_1 _4048_ (.B1(net652),
    .Y(_1365_),
    .A1(net632),
    .A2(_1364_));
 sg13g2_a22oi_1 _4049_ (.Y(_1366_),
    .B1(_1364_),
    .B2(net683),
    .A2(_1360_),
    .A1(_1359_));
 sg13g2_o21ai_1 _4050_ (.B1(_1366_),
    .Y(_0019_),
    .A1(_1362_),
    .A2(_1365_));
 sg13g2_xor2_1 _4051_ (.B(_0618_),
    .A(_0544_),
    .X(_1367_));
 sg13g2_a21oi_1 _4052_ (.A1(net551),
    .A2(_1367_),
    .Y(_1368_),
    .B1(net702));
 sg13g2_o21ai_1 _4053_ (.B1(net639),
    .Y(_1369_),
    .A1(net717),
    .A2(_0498_));
 sg13g2_nor2_1 _4054_ (.A(_1368_),
    .B(_1369_),
    .Y(_1370_));
 sg13g2_nand2_1 _4055_ (.Y(_1371_),
    .A(net734),
    .B(net572));
 sg13g2_a21oi_1 _4056_ (.A1(net3),
    .A2(net578),
    .Y(_1372_),
    .B1(_0680_));
 sg13g2_nand2b_1 _4057_ (.Y(_1373_),
    .B(net549),
    .A_N(_0902_));
 sg13g2_a21oi_1 _4058_ (.A1(_1080_),
    .A2(net545),
    .Y(_1374_),
    .B1(_0681_));
 sg13g2_a221oi_1 _4059_ (.B2(_1374_),
    .C1(_0666_),
    .B1(_1373_),
    .A1(_1371_),
    .Y(_1375_),
    .A2(_1372_));
 sg13g2_or2_1 _4060_ (.X(_0020_),
    .B(_1375_),
    .A(_1370_));
 sg13g2_nor2_1 _4061_ (.A(net717),
    .B(_0495_),
    .Y(_1376_));
 sg13g2_a21oi_1 _4062_ (.A1(_0624_),
    .A2(net542),
    .Y(_1377_),
    .B1(_1376_));
 sg13g2_nor2_1 _4063_ (.A(net4),
    .B(net571),
    .Y(_1378_));
 sg13g2_a21oi_1 _4064_ (.A1(_1929_),
    .A2(net571),
    .Y(_1379_),
    .B1(_1378_));
 sg13g2_xnor2_1 _4065_ (.Y(_1380_),
    .A(_0829_),
    .B(_0896_));
 sg13g2_a221oi_1 _4066_ (.B2(net550),
    .C1(net628),
    .B1(_1380_),
    .A1(_1077_),
    .Y(_1381_),
    .A2(net545));
 sg13g2_o21ai_1 _4067_ (.B1(net652),
    .Y(_1382_),
    .A1(net632),
    .A2(_1379_));
 sg13g2_nor2_1 _4068_ (.A(_1381_),
    .B(_1382_),
    .Y(_1383_));
 sg13g2_a21oi_1 _4069_ (.A1(net684),
    .A2(_1379_),
    .Y(_1384_),
    .B1(_1383_));
 sg13g2_o21ai_1 _4070_ (.B1(_1384_),
    .Y(_0021_),
    .A1(net637),
    .A2(_1377_));
 sg13g2_a22oi_1 _4071_ (.Y(_1385_),
    .B1(_0623_),
    .B2(net542),
    .A2(_0518_),
    .A1(net702));
 sg13g2_mux2_1 _4072_ (.A0(net387),
    .A1(net5),
    .S(net578),
    .X(_1386_));
 sg13g2_a21oi_1 _4073_ (.A1(_1067_),
    .A2(net545),
    .Y(_1387_),
    .B1(net628));
 sg13g2_o21ai_1 _4074_ (.B1(_1387_),
    .Y(_1388_),
    .A1(_0901_),
    .A2(_0934_));
 sg13g2_nor2_1 _4075_ (.A(net632),
    .B(_1386_),
    .Y(_1389_));
 sg13g2_nor2_1 _4076_ (.A(net634),
    .B(_1389_),
    .Y(_1390_));
 sg13g2_a22oi_1 _4077_ (.Y(_1391_),
    .B1(_1388_),
    .B2(_1390_),
    .A2(_1386_),
    .A1(net692));
 sg13g2_o21ai_1 _4078_ (.B1(_1391_),
    .Y(_0022_),
    .A1(net637),
    .A2(_1385_));
 sg13g2_xor2_1 _4079_ (.B(_0621_),
    .A(_0538_),
    .X(_1392_));
 sg13g2_a21oi_1 _4080_ (.A1(net552),
    .A2(_1392_),
    .Y(_1393_),
    .B1(net702));
 sg13g2_o21ai_1 _4081_ (.B1(net639),
    .Y(_1394_),
    .A1(net718),
    .A2(_0522_));
 sg13g2_mux2_1 _4082_ (.A0(net389),
    .A1(net6),
    .S(net578),
    .X(_1395_));
 sg13g2_xor2_1 _4083_ (.B(_0898_),
    .A(_0826_),
    .X(_1396_));
 sg13g2_a221oi_1 _4084_ (.B2(net549),
    .C1(net628),
    .B1(_1396_),
    .A1(_1061_),
    .Y(_1397_),
    .A2(net546));
 sg13g2_o21ai_1 _4085_ (.B1(net652),
    .Y(_1398_),
    .A1(net633),
    .A2(_1395_));
 sg13g2_nor2_1 _4086_ (.A(_1397_),
    .B(_1398_),
    .Y(_1399_));
 sg13g2_a21oi_1 _4087_ (.A1(net684),
    .A2(_1395_),
    .Y(_1400_),
    .B1(_1399_));
 sg13g2_o21ai_1 _4088_ (.B1(_1400_),
    .Y(_0023_),
    .A1(_1393_),
    .A2(_1394_));
 sg13g2_nor2_1 _4089_ (.A(net703),
    .B(_0622_),
    .Y(_1401_));
 sg13g2_a22oi_1 _4090_ (.Y(_1402_),
    .B1(_0662_),
    .B2(_1401_),
    .A2(_0354_),
    .A1(net702));
 sg13g2_nand2b_1 _4091_ (.Y(_1403_),
    .B(net639),
    .A_N(_1402_));
 sg13g2_nand2_1 _4092_ (.Y(_1404_),
    .A(net7),
    .B(net576));
 sg13g2_o21ai_1 _4093_ (.B1(_1404_),
    .Y(_1405_),
    .A1(_1935_),
    .A2(net576));
 sg13g2_nand2_1 _4094_ (.Y(_1406_),
    .A(net684),
    .B(_1405_));
 sg13g2_nand2b_1 _4095_ (.Y(_1407_),
    .B(_0676_),
    .A_N(_0930_));
 sg13g2_nor2_1 _4096_ (.A(_0675_),
    .B(_1131_),
    .Y(_1408_));
 sg13g2_a21oi_1 _4097_ (.A1(_1046_),
    .A2(_1408_),
    .Y(_1409_),
    .B1(net628));
 sg13g2_o21ai_1 _4098_ (.B1(_1409_),
    .Y(_1410_),
    .A1(_0900_),
    .A2(_1407_));
 sg13g2_o21ai_1 _4099_ (.B1(net652),
    .Y(_1411_),
    .A1(net632),
    .A2(_1405_));
 sg13g2_nand2b_1 _4100_ (.Y(_1412_),
    .B(_1410_),
    .A_N(_1411_));
 sg13g2_nand3_1 _4101_ (.B(_1406_),
    .C(_1412_),
    .A(_1403_),
    .Y(_0025_));
 sg13g2_nor2_1 _4102_ (.A(net8),
    .B(net572),
    .Y(_1413_));
 sg13g2_nor2_1 _4103_ (.A(net237),
    .B(net578),
    .Y(_1414_));
 sg13g2_nor4_1 _4104_ (.A(_0666_),
    .B(_0680_),
    .C(_1413_),
    .D(_1414_),
    .Y(_0026_));
 sg13g2_and2_1 _4105_ (.A(net1),
    .B(_2084_),
    .X(_1415_));
 sg13g2_nand3_1 _4106_ (.B(net652),
    .C(net661),
    .A(net9),
    .Y(_1416_));
 sg13g2_o21ai_1 _4107_ (.B1(_1416_),
    .Y(_0098_),
    .A1(net703),
    .A2(net652));
 sg13g2_nand2b_1 _4108_ (.Y(_1417_),
    .B(_0673_),
    .A_N(_2084_));
 sg13g2_nand3_1 _4109_ (.B(_2086_),
    .C(_1417_),
    .A(net1),
    .Y(_1418_));
 sg13g2_and2_1 _4110_ (.A(net696),
    .B(_1418_),
    .X(_1419_));
 sg13g2_nor2_1 _4111_ (.A(net27),
    .B(net619),
    .Y(_0099_));
 sg13g2_nor3_1 _4112_ (.A(net27),
    .B(net209),
    .C(net619),
    .Y(_1420_));
 sg13g2_a21o_1 _4113_ (.A2(net209),
    .A1(net27),
    .B1(_1420_),
    .X(_0100_));
 sg13g2_nor2b_1 _4114_ (.A(net30),
    .B_N(_1420_),
    .Y(_1421_));
 sg13g2_xor2_1 _4115_ (.B(_1420_),
    .A(net30),
    .X(_0101_));
 sg13g2_nand2b_1 _4116_ (.Y(_1422_),
    .B(_1421_),
    .A_N(net28));
 sg13g2_xor2_1 _4117_ (.B(_1421_),
    .A(net28),
    .X(_0102_));
 sg13g2_nor2_1 _4118_ (.A(net692),
    .B(_1418_),
    .Y(_1423_));
 sg13g2_or2_1 _4119_ (.X(_1424_),
    .B(_1418_),
    .A(net692));
 sg13g2_a21o_1 _4120_ (.A2(_1422_),
    .A1(net38),
    .B1(net605),
    .X(_0103_));
 sg13g2_nand2_1 _4121_ (.Y(_1425_),
    .A(net34),
    .B(net621));
 sg13g2_nand3_1 _4122_ (.B(net32),
    .C(net686),
    .A(net712),
    .Y(_1426_));
 sg13g2_nand2_1 _4123_ (.Y(_0104_),
    .A(_1425_),
    .B(_1426_));
 sg13g2_nand2_1 _4124_ (.Y(_1427_),
    .A(net712),
    .B(net55));
 sg13g2_xnor2_1 _4125_ (.Y(_1428_),
    .A(net34),
    .B(_1427_));
 sg13g2_a22oi_1 _4126_ (.Y(_1429_),
    .B1(_1428_),
    .B2(net685),
    .A2(net621),
    .A1(net357));
 sg13g2_inv_1 _4127_ (.Y(_0105_),
    .A(_1429_));
 sg13g2_nand2_1 _4128_ (.Y(_1430_),
    .A(\mul_operand_r[2] ),
    .B(\mul_accum[1] ));
 sg13g2_xnor2_1 _4129_ (.Y(_1431_),
    .A(\mul_operand_r[2] ),
    .B(\mul_accum[1] ));
 sg13g2_nand2_1 _4130_ (.Y(_1432_),
    .A(net55),
    .B(net34));
 sg13g2_xnor2_1 _4131_ (.Y(_1433_),
    .A(_1431_),
    .B(_1432_));
 sg13g2_o21ai_1 _4132_ (.B1(net685),
    .Y(_1434_),
    .A1(net712),
    .A2(\mul_accum[1] ));
 sg13g2_a21oi_1 _4133_ (.A1(net712),
    .A2(_1433_),
    .Y(_1435_),
    .B1(_1434_));
 sg13g2_a21o_1 _4134_ (.A2(net621),
    .A1(net334),
    .B1(_1435_),
    .X(_0106_));
 sg13g2_and2_1 _4135_ (.A(\mul_operand_r[3] ),
    .B(\mul_accum[2] ),
    .X(_1436_));
 sg13g2_xor2_1 _4136_ (.B(\mul_accum[2] ),
    .A(\mul_operand_r[3] ),
    .X(_1437_));
 sg13g2_o21ai_1 _4137_ (.B1(_1430_),
    .Y(_1438_),
    .A1(_1431_),
    .A2(_1432_));
 sg13g2_xnor2_1 _4138_ (.Y(_1439_),
    .A(_1437_),
    .B(_1438_));
 sg13g2_o21ai_1 _4139_ (.B1(net685),
    .Y(_1440_),
    .A1(net713),
    .A2(\mul_accum[2] ));
 sg13g2_a21oi_1 _4140_ (.A1(net713),
    .A2(_1439_),
    .Y(_1441_),
    .B1(_1440_));
 sg13g2_a21o_1 _4141_ (.A2(net621),
    .A1(net331),
    .B1(_1441_),
    .X(_0107_));
 sg13g2_nand2_1 _4142_ (.Y(_1442_),
    .A(\mul_operand_r[4] ),
    .B(\mul_accum[3] ));
 sg13g2_xnor2_1 _4143_ (.Y(_1443_),
    .A(\mul_operand_r[4] ),
    .B(\mul_accum[3] ));
 sg13g2_a21oi_1 _4144_ (.A1(_1437_),
    .A2(_1438_),
    .Y(_1444_),
    .B1(_1436_));
 sg13g2_xnor2_1 _4145_ (.Y(_1445_),
    .A(_1443_),
    .B(_1444_));
 sg13g2_o21ai_1 _4146_ (.B1(net685),
    .Y(_1446_),
    .A1(net713),
    .A2(\mul_accum[3] ));
 sg13g2_a21oi_1 _4147_ (.A1(net713),
    .A2(_1445_),
    .Y(_1447_),
    .B1(_1446_));
 sg13g2_a21o_1 _4148_ (.A2(net621),
    .A1(net329),
    .B1(_1447_),
    .X(_0108_));
 sg13g2_and2_1 _4149_ (.A(\mul_operand_r[5] ),
    .B(\mul_accum[4] ),
    .X(_1448_));
 sg13g2_xor2_1 _4150_ (.B(\mul_accum[4] ),
    .A(\mul_operand_r[5] ),
    .X(_1449_));
 sg13g2_o21ai_1 _4151_ (.B1(_1442_),
    .Y(_1450_),
    .A1(_1443_),
    .A2(_1444_));
 sg13g2_xnor2_1 _4152_ (.Y(_1451_),
    .A(_1449_),
    .B(_1450_));
 sg13g2_o21ai_1 _4153_ (.B1(net685),
    .Y(_1452_),
    .A1(net712),
    .A2(net329));
 sg13g2_a21oi_1 _4154_ (.A1(net712),
    .A2(_1451_),
    .Y(_1453_),
    .B1(_1452_));
 sg13g2_a21o_1 _4155_ (.A2(net621),
    .A1(net342),
    .B1(_1453_),
    .X(_0109_));
 sg13g2_a21oi_1 _4156_ (.A1(_1449_),
    .A2(_1450_),
    .Y(_1454_),
    .B1(_1448_));
 sg13g2_nor2_1 _4157_ (.A(\mul_operand_r[6] ),
    .B(\mul_accum[5] ),
    .Y(_1455_));
 sg13g2_xnor2_1 _4158_ (.Y(_1456_),
    .A(net103),
    .B(\mul_accum[5] ));
 sg13g2_xnor2_1 _4159_ (.Y(_1457_),
    .A(_1454_),
    .B(_1456_));
 sg13g2_o21ai_1 _4160_ (.B1(net679),
    .Y(_1458_),
    .A1(net712),
    .A2(\mul_accum[5] ));
 sg13g2_a21oi_1 _4161_ (.A1(net712),
    .A2(_1457_),
    .Y(_1459_),
    .B1(_1458_));
 sg13g2_a21o_1 _4162_ (.A2(net613),
    .A1(net336),
    .B1(_1459_),
    .X(_0110_));
 sg13g2_nand2_1 _4163_ (.Y(_1460_),
    .A(net207),
    .B(net613));
 sg13g2_nand2_1 _4164_ (.Y(_1461_),
    .A(\mul_operand_r[7] ),
    .B(\mul_accum[6] ));
 sg13g2_xnor2_1 _4165_ (.Y(_1462_),
    .A(\mul_operand_r[7] ),
    .B(\mul_accum[6] ));
 sg13g2_a221oi_1 _4166_ (.B2(_1450_),
    .C1(_1448_),
    .B1(_1449_),
    .A1(\mul_operand_r[6] ),
    .Y(_1463_),
    .A2(\mul_accum[5] ));
 sg13g2_o21ai_1 _4167_ (.B1(_1462_),
    .Y(_1464_),
    .A1(_1455_),
    .A2(_1463_));
 sg13g2_or3_1 _4168_ (.A(_1455_),
    .B(_1462_),
    .C(_1463_),
    .X(_1465_));
 sg13g2_a21oi_1 _4169_ (.A1(_1464_),
    .A2(_1465_),
    .Y(_1466_),
    .B1(_1940_));
 sg13g2_o21ai_1 _4170_ (.B1(net679),
    .Y(_1467_),
    .A1(net708),
    .A2(\mul_accum[6] ));
 sg13g2_o21ai_1 _4171_ (.B1(_1460_),
    .Y(_0111_),
    .A1(_1466_),
    .A2(_1467_));
 sg13g2_and2_1 _4172_ (.A(\mul_operand_r[8] ),
    .B(\mul_accum[7] ),
    .X(_1468_));
 sg13g2_xnor2_1 _4173_ (.Y(_1469_),
    .A(\mul_operand_r[8] ),
    .B(\mul_accum[7] ));
 sg13g2_nand2_1 _4174_ (.Y(_1470_),
    .A(_1461_),
    .B(_1465_));
 sg13g2_a21oi_1 _4175_ (.A1(_1461_),
    .A2(_1465_),
    .Y(_1471_),
    .B1(_1469_));
 sg13g2_xor2_1 _4176_ (.B(_1470_),
    .A(_1469_),
    .X(_1472_));
 sg13g2_o21ai_1 _4177_ (.B1(net679),
    .Y(_1473_),
    .A1(net708),
    .A2(net207));
 sg13g2_a21oi_1 _4178_ (.A1(net708),
    .A2(_1472_),
    .Y(_1474_),
    .B1(_1473_));
 sg13g2_a21o_1 _4179_ (.A2(net611),
    .A1(net315),
    .B1(_1474_),
    .X(_0112_));
 sg13g2_and2_1 _4180_ (.A(net364),
    .B(net610),
    .X(_1475_));
 sg13g2_nand2_1 _4181_ (.Y(_1476_),
    .A(\mul_operand_r[9] ),
    .B(\mul_accum[8] ));
 sg13g2_xor2_1 _4182_ (.B(\mul_accum[8] ),
    .A(\mul_operand_r[9] ),
    .X(_1477_));
 sg13g2_nor3_1 _4183_ (.A(_1468_),
    .B(_1471_),
    .C(_1477_),
    .Y(_1478_));
 sg13g2_o21ai_1 _4184_ (.B1(_1477_),
    .Y(_1479_),
    .A1(_1468_),
    .A2(_1471_));
 sg13g2_nor2b_1 _4185_ (.A(_1478_),
    .B_N(_1479_),
    .Y(_1480_));
 sg13g2_mux2_1 _4186_ (.A0(net315),
    .A1(_1480_),
    .S(net708),
    .X(_1481_));
 sg13g2_a21o_1 _4187_ (.A2(_1481_),
    .A1(net676),
    .B1(_1475_),
    .X(_0113_));
 sg13g2_nand2_1 _4188_ (.Y(_1482_),
    .A(_1476_),
    .B(_1479_));
 sg13g2_or2_1 _4189_ (.X(_1483_),
    .B(\mul_accum[9] ),
    .A(\mul_operand_r[10] ));
 sg13g2_nand2_1 _4190_ (.Y(_1484_),
    .A(\mul_operand_r[10] ),
    .B(\mul_accum[9] ));
 sg13g2_and2_1 _4191_ (.A(_1483_),
    .B(_1484_),
    .X(_1485_));
 sg13g2_xnor2_1 _4192_ (.Y(_1486_),
    .A(_1482_),
    .B(_1485_));
 sg13g2_o21ai_1 _4193_ (.B1(net677),
    .Y(_1487_),
    .A1(net706),
    .A2(\mul_accum[9] ));
 sg13g2_a21oi_1 _4194_ (.A1(net706),
    .A2(_1486_),
    .Y(_1488_),
    .B1(_1487_));
 sg13g2_a21o_1 _4195_ (.A2(net611),
    .A1(net324),
    .B1(_1488_),
    .X(_0114_));
 sg13g2_nand2_1 _4196_ (.Y(_1489_),
    .A(net190),
    .B(net610));
 sg13g2_nand2_1 _4197_ (.Y(_1490_),
    .A(\mul_operand_r[11] ),
    .B(\mul_accum[10] ));
 sg13g2_xor2_1 _4198_ (.B(\mul_accum[10] ),
    .A(\mul_operand_r[11] ),
    .X(_1491_));
 sg13g2_nand3_1 _4199_ (.B(_1479_),
    .C(_1484_),
    .A(_1476_),
    .Y(_1492_));
 sg13g2_a21o_1 _4200_ (.A2(_1492_),
    .A1(_1483_),
    .B1(_1491_),
    .X(_1493_));
 sg13g2_nand3_1 _4201_ (.B(_1491_),
    .C(_1492_),
    .A(_1483_),
    .Y(_1494_));
 sg13g2_a21oi_1 _4202_ (.A1(_1493_),
    .A2(_1494_),
    .Y(_1495_),
    .B1(_1940_));
 sg13g2_o21ai_1 _4203_ (.B1(net676),
    .Y(_1496_),
    .A1(net707),
    .A2(\mul_accum[10] ));
 sg13g2_o21ai_1 _4204_ (.B1(_1489_),
    .Y(_0115_),
    .A1(_1495_),
    .A2(_1496_));
 sg13g2_nand2_1 _4205_ (.Y(_1497_),
    .A(_1490_),
    .B(_1494_));
 sg13g2_or2_1 _4206_ (.X(_1498_),
    .B(\mul_accum[11] ),
    .A(\mul_operand_r[12] ));
 sg13g2_nand2_1 _4207_ (.Y(_1499_),
    .A(\mul_operand_r[12] ),
    .B(\mul_accum[11] ));
 sg13g2_and2_1 _4208_ (.A(_1498_),
    .B(_1499_),
    .X(_1500_));
 sg13g2_xnor2_1 _4209_ (.Y(_1501_),
    .A(_1497_),
    .B(_1500_));
 sg13g2_o21ai_1 _4210_ (.B1(net676),
    .Y(_1502_),
    .A1(net706),
    .A2(net190));
 sg13g2_a21oi_1 _4211_ (.A1(net706),
    .A2(_1501_),
    .Y(_1503_),
    .B1(_1502_));
 sg13g2_a21o_1 _4212_ (.A2(net610),
    .A1(net302),
    .B1(_1503_),
    .X(_0116_));
 sg13g2_and2_1 _4213_ (.A(net363),
    .B(net610),
    .X(_1504_));
 sg13g2_nand2_1 _4214_ (.Y(_1505_),
    .A(\mul_operand_r[13] ),
    .B(\mul_accum[12] ));
 sg13g2_xor2_1 _4215_ (.B(\mul_accum[12] ),
    .A(\mul_operand_r[13] ),
    .X(_1506_));
 sg13g2_nand3_1 _4216_ (.B(_1494_),
    .C(_1499_),
    .A(_1490_),
    .Y(_1507_));
 sg13g2_a21oi_1 _4217_ (.A1(_1498_),
    .A2(_1507_),
    .Y(_1508_),
    .B1(_1506_));
 sg13g2_nand3_1 _4218_ (.B(_1506_),
    .C(_1507_),
    .A(_1498_),
    .Y(_1509_));
 sg13g2_nor2b_1 _4219_ (.A(_1508_),
    .B_N(_1509_),
    .Y(_1510_));
 sg13g2_mux2_1 _4220_ (.A0(net302),
    .A1(_1510_),
    .S(net706),
    .X(_1511_));
 sg13g2_a21o_1 _4221_ (.A2(_1511_),
    .A1(net676),
    .B1(_1504_),
    .X(_0117_));
 sg13g2_nand2_1 _4222_ (.Y(_1512_),
    .A(_1505_),
    .B(_1509_));
 sg13g2_or2_1 _4223_ (.X(_1513_),
    .B(\mul_accum[13] ),
    .A(\mul_operand_r[14] ));
 sg13g2_nand2_1 _4224_ (.Y(_1514_),
    .A(\mul_operand_r[14] ),
    .B(\mul_accum[13] ));
 sg13g2_and2_1 _4225_ (.A(_1513_),
    .B(_1514_),
    .X(_1515_));
 sg13g2_xnor2_1 _4226_ (.Y(_1516_),
    .A(_1512_),
    .B(_1515_));
 sg13g2_o21ai_1 _4227_ (.B1(net676),
    .Y(_1517_),
    .A1(net706),
    .A2(\mul_accum[13] ));
 sg13g2_a21oi_1 _4228_ (.A1(net706),
    .A2(_1516_),
    .Y(_1518_),
    .B1(_1517_));
 sg13g2_a21o_1 _4229_ (.A2(net612),
    .A1(net279),
    .B1(_1518_),
    .X(_0118_));
 sg13g2_nand2_1 _4230_ (.Y(_1519_),
    .A(net133),
    .B(net614));
 sg13g2_nand2_1 _4231_ (.Y(_1520_),
    .A(\mul_operand_r[15] ),
    .B(\mul_accum[14] ));
 sg13g2_xor2_1 _4232_ (.B(\mul_accum[14] ),
    .A(\mul_operand_r[15] ),
    .X(_1521_));
 sg13g2_nand3_1 _4233_ (.B(_1509_),
    .C(_1514_),
    .A(_1505_),
    .Y(_1522_));
 sg13g2_a21o_1 _4234_ (.A2(_1522_),
    .A1(_1513_),
    .B1(_1521_),
    .X(_1523_));
 sg13g2_nand3_1 _4235_ (.B(_1521_),
    .C(_1522_),
    .A(_1513_),
    .Y(_1524_));
 sg13g2_a21oi_1 _4236_ (.A1(_1523_),
    .A2(_1524_),
    .Y(_1525_),
    .B1(_1940_));
 sg13g2_o21ai_1 _4237_ (.B1(net677),
    .Y(_1526_),
    .A1(net707),
    .A2(\mul_accum[14] ));
 sg13g2_o21ai_1 _4238_ (.B1(_1519_),
    .Y(_0119_),
    .A1(_1525_),
    .A2(_1526_));
 sg13g2_nand2_1 _4239_ (.Y(_1527_),
    .A(_1520_),
    .B(_1524_));
 sg13g2_or2_1 _4240_ (.X(_1528_),
    .B(\mul_accum[15] ),
    .A(\mul_operand_r[16] ));
 sg13g2_nand2_1 _4241_ (.Y(_1529_),
    .A(\mul_operand_r[16] ),
    .B(\mul_accum[15] ));
 sg13g2_and2_1 _4242_ (.A(_1528_),
    .B(_1529_),
    .X(_1530_));
 sg13g2_xnor2_1 _4243_ (.Y(_1531_),
    .A(_1527_),
    .B(_1530_));
 sg13g2_o21ai_1 _4244_ (.B1(net680),
    .Y(_1532_),
    .A1(net707),
    .A2(net133));
 sg13g2_a21oi_1 _4245_ (.A1(net707),
    .A2(_1531_),
    .Y(_1533_),
    .B1(_1532_));
 sg13g2_a21o_1 _4246_ (.A2(net612),
    .A1(net286),
    .B1(_1533_),
    .X(_0120_));
 sg13g2_and2_1 _4247_ (.A(net360),
    .B(net612),
    .X(_1534_));
 sg13g2_nand2_1 _4248_ (.Y(_1535_),
    .A(\mul_operand_r[17] ),
    .B(\mul_accum[16] ));
 sg13g2_xor2_1 _4249_ (.B(\mul_accum[16] ),
    .A(\mul_operand_r[17] ),
    .X(_1536_));
 sg13g2_nand3_1 _4250_ (.B(_1524_),
    .C(_1529_),
    .A(_1520_),
    .Y(_1537_));
 sg13g2_a21oi_1 _4251_ (.A1(_1528_),
    .A2(_1537_),
    .Y(_1538_),
    .B1(_1536_));
 sg13g2_nand3_1 _4252_ (.B(_1536_),
    .C(_1537_),
    .A(_1528_),
    .Y(_1539_));
 sg13g2_nor2b_1 _4253_ (.A(_1538_),
    .B_N(_1539_),
    .Y(_1540_));
 sg13g2_mux2_1 _4254_ (.A0(net286),
    .A1(_1540_),
    .S(net707),
    .X(_1541_));
 sg13g2_a21o_1 _4255_ (.A2(_1541_),
    .A1(net677),
    .B1(_1534_),
    .X(_0121_));
 sg13g2_nand2_1 _4256_ (.Y(_1542_),
    .A(_1535_),
    .B(_1539_));
 sg13g2_nor2_1 _4257_ (.A(\mul_operand_r[18] ),
    .B(\mul_accum[17] ),
    .Y(_1543_));
 sg13g2_and2_1 _4258_ (.A(\mul_operand_r[18] ),
    .B(\mul_accum[17] ),
    .X(_1544_));
 sg13g2_nor2_1 _4259_ (.A(_1543_),
    .B(_1544_),
    .Y(_1545_));
 sg13g2_xnor2_1 _4260_ (.Y(_1546_),
    .A(_1542_),
    .B(_1545_));
 sg13g2_o21ai_1 _4261_ (.B1(net682),
    .Y(_1547_),
    .A1(net710),
    .A2(\mul_accum[17] ));
 sg13g2_a21oi_1 _4262_ (.A1(net710),
    .A2(_1546_),
    .Y(_1548_),
    .B1(_1547_));
 sg13g2_a21o_1 _4263_ (.A2(net617),
    .A1(net287),
    .B1(_1548_),
    .X(_0122_));
 sg13g2_nand2_1 _4264_ (.Y(_1549_),
    .A(\mul_operand_r[19] ),
    .B(\mul_accum[18] ));
 sg13g2_xnor2_1 _4265_ (.Y(_1550_),
    .A(\mul_operand_r[19] ),
    .B(\mul_accum[18] ));
 sg13g2_inv_1 _4266_ (.Y(_1551_),
    .A(_1550_));
 sg13g2_a21oi_1 _4267_ (.A1(_1535_),
    .A2(_1539_),
    .Y(_1552_),
    .B1(_1543_));
 sg13g2_nor3_1 _4268_ (.A(_1544_),
    .B(_1551_),
    .C(_1552_),
    .Y(_1553_));
 sg13g2_o21ai_1 _4269_ (.B1(_1551_),
    .Y(_1554_),
    .A1(_1544_),
    .A2(_1552_));
 sg13g2_nand2b_1 _4270_ (.Y(_1555_),
    .B(_1554_),
    .A_N(_1553_));
 sg13g2_o21ai_1 _4271_ (.B1(net682),
    .Y(_1556_),
    .A1(net710),
    .A2(\mul_accum[18] ));
 sg13g2_a21oi_1 _4272_ (.A1(net710),
    .A2(_1555_),
    .Y(_1557_),
    .B1(_1556_));
 sg13g2_a21o_1 _4273_ (.A2(net617),
    .A1(net272),
    .B1(_1557_),
    .X(_0123_));
 sg13g2_nand2_1 _4274_ (.Y(_1558_),
    .A(_1549_),
    .B(_1554_));
 sg13g2_nor2_1 _4275_ (.A(\mul_operand_r[20] ),
    .B(\mul_accum[19] ),
    .Y(_1559_));
 sg13g2_and2_1 _4276_ (.A(\mul_operand_r[20] ),
    .B(\mul_accum[19] ),
    .X(_1560_));
 sg13g2_nor2_1 _4277_ (.A(_1559_),
    .B(_1560_),
    .Y(_1561_));
 sg13g2_xnor2_1 _4278_ (.Y(_1562_),
    .A(_1558_),
    .B(_1561_));
 sg13g2_o21ai_1 _4279_ (.B1(net682),
    .Y(_1563_),
    .A1(net710),
    .A2(net272));
 sg13g2_a21oi_1 _4280_ (.A1(net710),
    .A2(_1562_),
    .Y(_1564_),
    .B1(_1563_));
 sg13g2_a21o_1 _4281_ (.A2(net617),
    .A1(net303),
    .B1(_1564_),
    .X(_0124_));
 sg13g2_nand2_1 _4282_ (.Y(_1565_),
    .A(\mul_operand_r[21] ),
    .B(\mul_accum[20] ));
 sg13g2_xor2_1 _4283_ (.B(\mul_accum[20] ),
    .A(\mul_operand_r[21] ),
    .X(_1566_));
 sg13g2_a21oi_1 _4284_ (.A1(_1549_),
    .A2(_1554_),
    .Y(_1567_),
    .B1(_1559_));
 sg13g2_nor3_1 _4285_ (.A(_1560_),
    .B(_1566_),
    .C(_1567_),
    .Y(_1568_));
 sg13g2_o21ai_1 _4286_ (.B1(_1566_),
    .Y(_1569_),
    .A1(_1560_),
    .A2(_1567_));
 sg13g2_nand2b_1 _4287_ (.Y(_1570_),
    .B(_1569_),
    .A_N(_1568_));
 sg13g2_o21ai_1 _4288_ (.B1(net682),
    .Y(_1571_),
    .A1(net710),
    .A2(\mul_accum[20] ));
 sg13g2_a21oi_1 _4289_ (.A1(net709),
    .A2(_1570_),
    .Y(_1572_),
    .B1(_1571_));
 sg13g2_a21o_1 _4290_ (.A2(net615),
    .A1(net299),
    .B1(_1572_),
    .X(_0125_));
 sg13g2_nand2_1 _4291_ (.Y(_1573_),
    .A(net157),
    .B(net615));
 sg13g2_nand2_1 _4292_ (.Y(_1574_),
    .A(_1565_),
    .B(_1569_));
 sg13g2_nor2_1 _4293_ (.A(\mul_operand_r[22] ),
    .B(\mul_accum[21] ),
    .Y(_1575_));
 sg13g2_and2_1 _4294_ (.A(\mul_operand_r[22] ),
    .B(\mul_accum[21] ),
    .X(_1576_));
 sg13g2_nor2_1 _4295_ (.A(_1575_),
    .B(_1576_),
    .Y(_1577_));
 sg13g2_xor2_1 _4296_ (.B(_1577_),
    .A(_1574_),
    .X(_1578_));
 sg13g2_nor2_1 _4297_ (.A(_1940_),
    .B(_1578_),
    .Y(_1579_));
 sg13g2_o21ai_1 _4298_ (.B1(net681),
    .Y(_1580_),
    .A1(net709),
    .A2(\mul_accum[21] ));
 sg13g2_o21ai_1 _4299_ (.B1(_1573_),
    .Y(_0126_),
    .A1(_1579_),
    .A2(_1580_));
 sg13g2_nand2_1 _4300_ (.Y(_1581_),
    .A(\mul_operand_r[23] ),
    .B(\mul_accum[22] ));
 sg13g2_xnor2_1 _4301_ (.Y(_1582_),
    .A(\mul_operand_r[23] ),
    .B(\mul_accum[22] ));
 sg13g2_inv_1 _4302_ (.Y(_1583_),
    .A(_1582_));
 sg13g2_a21oi_1 _4303_ (.A1(_1565_),
    .A2(_1569_),
    .Y(_1584_),
    .B1(_1575_));
 sg13g2_nor3_1 _4304_ (.A(_1576_),
    .B(_1583_),
    .C(_1584_),
    .Y(_1585_));
 sg13g2_o21ai_1 _4305_ (.B1(_1583_),
    .Y(_1586_),
    .A1(_1576_),
    .A2(_1584_));
 sg13g2_nand2b_1 _4306_ (.Y(_1587_),
    .B(_1586_),
    .A_N(_1585_));
 sg13g2_o21ai_1 _4307_ (.B1(net681),
    .Y(_1588_),
    .A1(net709),
    .A2(net157));
 sg13g2_a21oi_1 _4308_ (.A1(net709),
    .A2(_1587_),
    .Y(_1589_),
    .B1(_1588_));
 sg13g2_a21o_1 _4309_ (.A2(net616),
    .A1(net255),
    .B1(_1589_),
    .X(_0127_));
 sg13g2_nand2_1 _4310_ (.Y(_1590_),
    .A(_1581_),
    .B(_1586_));
 sg13g2_nor2_1 _4311_ (.A(\mul_operand_r[24] ),
    .B(\mul_accum[23] ),
    .Y(_1591_));
 sg13g2_and2_1 _4312_ (.A(\mul_operand_r[24] ),
    .B(\mul_accum[23] ),
    .X(_1592_));
 sg13g2_o21ai_1 _4313_ (.B1(_1590_),
    .Y(_1593_),
    .A1(_1591_),
    .A2(_1592_));
 sg13g2_nor3_1 _4314_ (.A(_1590_),
    .B(_1591_),
    .C(_1592_),
    .Y(_1594_));
 sg13g2_nor2_1 _4315_ (.A(_1940_),
    .B(_1594_),
    .Y(_1595_));
 sg13g2_a221oi_1 _4316_ (.B2(_1595_),
    .C1(net694),
    .B1(_1593_),
    .A1(_1940_),
    .Y(_1596_),
    .A2(_1943_));
 sg13g2_a21o_1 _4317_ (.A2(net615),
    .A1(net305),
    .B1(_1596_),
    .X(_0128_));
 sg13g2_nand2_1 _4318_ (.Y(_1597_),
    .A(\mul_operand_r[25] ),
    .B(\mul_accum[24] ));
 sg13g2_xnor2_1 _4319_ (.Y(_1598_),
    .A(\mul_operand_r[25] ),
    .B(\mul_accum[24] ));
 sg13g2_inv_1 _4320_ (.Y(_1599_),
    .A(_1598_));
 sg13g2_a21oi_1 _4321_ (.A1(_1581_),
    .A2(_1586_),
    .Y(_1600_),
    .B1(_1591_));
 sg13g2_nor3_1 _4322_ (.A(_1592_),
    .B(_1599_),
    .C(_1600_),
    .Y(_1601_));
 sg13g2_o21ai_1 _4323_ (.B1(_1599_),
    .Y(_1602_),
    .A1(_1592_),
    .A2(_1600_));
 sg13g2_nand2b_1 _4324_ (.Y(_1603_),
    .B(_1602_),
    .A_N(_1601_));
 sg13g2_o21ai_1 _4325_ (.B1(net681),
    .Y(_1604_),
    .A1(net709),
    .A2(\mul_accum[24] ));
 sg13g2_a21oi_1 _4326_ (.A1(net709),
    .A2(_1603_),
    .Y(_1605_),
    .B1(_1604_));
 sg13g2_a21o_1 _4327_ (.A2(net615),
    .A1(net281),
    .B1(_1605_),
    .X(_0129_));
 sg13g2_nand2_1 _4328_ (.Y(_1606_),
    .A(_1597_),
    .B(_1602_));
 sg13g2_nor2_1 _4329_ (.A(\mul_operand_r[26] ),
    .B(\mul_accum[25] ),
    .Y(_1607_));
 sg13g2_and2_1 _4330_ (.A(\mul_operand_r[26] ),
    .B(\mul_accum[25] ),
    .X(_1608_));
 sg13g2_nor2_1 _4331_ (.A(_1607_),
    .B(_1608_),
    .Y(_1609_));
 sg13g2_xnor2_1 _4332_ (.Y(_1610_),
    .A(_1606_),
    .B(_1609_));
 sg13g2_o21ai_1 _4333_ (.B1(net681),
    .Y(_1611_),
    .A1(net709),
    .A2(net281));
 sg13g2_a21oi_1 _4334_ (.A1(net709),
    .A2(_1610_),
    .Y(_1612_),
    .B1(_1611_));
 sg13g2_a21o_1 _4335_ (.A2(net616),
    .A1(net285),
    .B1(_1612_),
    .X(_0130_));
 sg13g2_nand2_1 _4336_ (.Y(_1613_),
    .A(\mul_operand_r[27] ),
    .B(\mul_accum[26] ));
 sg13g2_xnor2_1 _4337_ (.Y(_1614_),
    .A(\mul_operand_r[27] ),
    .B(\mul_accum[26] ));
 sg13g2_inv_1 _4338_ (.Y(_1615_),
    .A(_1614_));
 sg13g2_a21oi_1 _4339_ (.A1(_1597_),
    .A2(_1602_),
    .Y(_1616_),
    .B1(_1607_));
 sg13g2_nor3_1 _4340_ (.A(_1608_),
    .B(_1615_),
    .C(_1616_),
    .Y(_1617_));
 sg13g2_o21ai_1 _4341_ (.B1(_1615_),
    .Y(_1618_),
    .A1(_1608_),
    .A2(_1616_));
 sg13g2_nand2b_1 _4342_ (.Y(_1619_),
    .B(_1618_),
    .A_N(_1617_));
 sg13g2_o21ai_1 _4343_ (.B1(net682),
    .Y(_1620_),
    .A1(net711),
    .A2(net285));
 sg13g2_a21oi_1 _4344_ (.A1(net711),
    .A2(_1619_),
    .Y(_1621_),
    .B1(_1620_));
 sg13g2_a21o_1 _4345_ (.A2(net616),
    .A1(net313),
    .B1(_1621_),
    .X(_0131_));
 sg13g2_nand2_1 _4346_ (.Y(_1622_),
    .A(_1613_),
    .B(_1618_));
 sg13g2_nor2_1 _4347_ (.A(\mul_operand_r[28] ),
    .B(\mul_accum[27] ),
    .Y(_1623_));
 sg13g2_and2_1 _4348_ (.A(\mul_operand_r[28] ),
    .B(\mul_accum[27] ),
    .X(_1624_));
 sg13g2_nor2_1 _4349_ (.A(_1623_),
    .B(_1624_),
    .Y(_1625_));
 sg13g2_xnor2_1 _4350_ (.Y(_1626_),
    .A(_1622_),
    .B(_1625_));
 sg13g2_o21ai_1 _4351_ (.B1(net684),
    .Y(_1627_),
    .A1(net711),
    .A2(\mul_accum[27] ));
 sg13g2_a21oi_1 _4352_ (.A1(net711),
    .A2(_1626_),
    .Y(_1628_),
    .B1(_1627_));
 sg13g2_a21o_1 _4353_ (.A2(net618),
    .A1(net265),
    .B1(_1628_),
    .X(_0132_));
 sg13g2_nand2_1 _4354_ (.Y(_1629_),
    .A(net258),
    .B(net618));
 sg13g2_nand2_1 _4355_ (.Y(_1630_),
    .A(\mul_operand_r[29] ),
    .B(\mul_accum[28] ));
 sg13g2_xor2_1 _4356_ (.B(\mul_accum[28] ),
    .A(\mul_operand_r[29] ),
    .X(_1631_));
 sg13g2_a21oi_1 _4357_ (.A1(_1613_),
    .A2(_1618_),
    .Y(_1632_),
    .B1(_1623_));
 sg13g2_nor3_1 _4358_ (.A(_1624_),
    .B(_1631_),
    .C(_1632_),
    .Y(_1633_));
 sg13g2_o21ai_1 _4359_ (.B1(_1631_),
    .Y(_1634_),
    .A1(_1624_),
    .A2(_1632_));
 sg13g2_nor2b_1 _4360_ (.A(_1633_),
    .B_N(_1634_),
    .Y(_1635_));
 sg13g2_nor2_1 _4361_ (.A(_1940_),
    .B(_1635_),
    .Y(_1636_));
 sg13g2_o21ai_1 _4362_ (.B1(net684),
    .Y(_1637_),
    .A1(net711),
    .A2(\mul_accum[28] ));
 sg13g2_o21ai_1 _4363_ (.B1(_1629_),
    .Y(_0133_),
    .A1(_1636_),
    .A2(_1637_));
 sg13g2_nand2_1 _4364_ (.Y(_1638_),
    .A(_1630_),
    .B(_1634_));
 sg13g2_nand2_1 _4365_ (.Y(_1639_),
    .A(\mul_operand_r[30] ),
    .B(\mul_accum[29] ));
 sg13g2_xor2_1 _4366_ (.B(\mul_accum[29] ),
    .A(net180),
    .X(_1640_));
 sg13g2_xnor2_1 _4367_ (.Y(_1641_),
    .A(_1638_),
    .B(_1640_));
 sg13g2_o21ai_1 _4368_ (.B1(net684),
    .Y(_1642_),
    .A1(net714),
    .A2(net258));
 sg13g2_a21oi_1 _4369_ (.A1(net714),
    .A2(_1641_),
    .Y(_1643_),
    .B1(_1642_));
 sg13g2_a21o_1 _4370_ (.A2(net618),
    .A1(net361),
    .B1(_1643_),
    .X(_0134_));
 sg13g2_and3_2 _4371_ (.X(_1644_),
    .A(_1630_),
    .B(_1634_),
    .C(_1639_));
 sg13g2_o21ai_1 _4372_ (.B1(net714),
    .Y(_1645_),
    .A1(\mul_operand_r[30] ),
    .A2(\mul_accum[29] ));
 sg13g2_nor2_1 _4373_ (.A(_1644_),
    .B(_1645_),
    .Y(_1646_));
 sg13g2_xor2_1 _4374_ (.B(_1646_),
    .A(\mul_accum[30] ),
    .X(_1647_));
 sg13g2_a22oi_1 _4375_ (.Y(_1648_),
    .B1(_1647_),
    .B2(net679),
    .A2(net613),
    .A1(net267));
 sg13g2_inv_1 _4376_ (.Y(_0135_),
    .A(net268));
 sg13g2_a21oi_1 _4377_ (.A1(\mul_accum[30] ),
    .A2(_1646_),
    .Y(_1649_),
    .B1(\mul_accum[31] ));
 sg13g2_nand2_1 _4378_ (.Y(_1650_),
    .A(\mul_accum[30] ),
    .B(net267));
 sg13g2_nor3_1 _4379_ (.A(_1644_),
    .B(_1645_),
    .C(_1650_),
    .Y(_1651_));
 sg13g2_nor3_1 _4380_ (.A(net695),
    .B(_1649_),
    .C(_1651_),
    .Y(_1652_));
 sg13g2_a21o_1 _4381_ (.A2(net613),
    .A1(net205),
    .B1(_1652_),
    .X(_0136_));
 sg13g2_nor4_2 _4382_ (.A(_1945_),
    .B(_1644_),
    .C(_1645_),
    .Y(_1653_),
    .D(_1650_));
 sg13g2_xnor2_1 _4383_ (.Y(_1654_),
    .A(_1945_),
    .B(_1651_));
 sg13g2_a22oi_1 _4384_ (.Y(_1655_),
    .B1(_1654_),
    .B2(net679),
    .A2(net613),
    .A1(net352));
 sg13g2_inv_1 _4385_ (.Y(_0137_),
    .A(_1655_));
 sg13g2_nand2_1 _4386_ (.Y(_1656_),
    .A(net151),
    .B(net614));
 sg13g2_xnor2_1 _4387_ (.Y(_1657_),
    .A(\mul_accum[33] ),
    .B(_1653_));
 sg13g2_o21ai_1 _4388_ (.B1(_1656_),
    .Y(_0138_),
    .A1(net695),
    .A2(_1657_));
 sg13g2_a21oi_1 _4389_ (.A1(\mul_accum[33] ),
    .A2(_1653_),
    .Y(_1658_),
    .B1(net151));
 sg13g2_nand3_1 _4390_ (.B(net151),
    .C(_1653_),
    .A(\mul_accum[33] ),
    .Y(_1659_));
 sg13g2_nor2_1 _4391_ (.A(net695),
    .B(_1658_),
    .Y(_1660_));
 sg13g2_a22oi_1 _4392_ (.Y(_1661_),
    .B1(_1659_),
    .B2(_1660_),
    .A2(net614),
    .A1(net253));
 sg13g2_inv_1 _4393_ (.Y(_0139_),
    .A(net254));
 sg13g2_nand4_1 _4394_ (.B(net151),
    .C(net253),
    .A(\mul_accum[33] ),
    .Y(_1662_),
    .D(_1653_));
 sg13g2_a21oi_1 _4395_ (.A1(_1946_),
    .A2(_1659_),
    .Y(_1663_),
    .B1(net695));
 sg13g2_a22oi_1 _4396_ (.Y(_1664_),
    .B1(_1662_),
    .B2(_1663_),
    .A2(net613),
    .A1(net293));
 sg13g2_inv_1 _4397_ (.Y(_0140_),
    .A(net294));
 sg13g2_nor2_1 _4398_ (.A(_1947_),
    .B(_1662_),
    .Y(_1665_));
 sg13g2_xnor2_1 _4399_ (.Y(_1666_),
    .A(\mul_accum[36] ),
    .B(_1662_));
 sg13g2_a22oi_1 _4400_ (.Y(_1667_),
    .B1(_1666_),
    .B2(net679),
    .A2(net613),
    .A1(net289));
 sg13g2_inv_1 _4401_ (.Y(_0141_),
    .A(net290));
 sg13g2_nand2_1 _4402_ (.Y(_1668_),
    .A(net289),
    .B(_1665_));
 sg13g2_xnor2_1 _4403_ (.Y(_1669_),
    .A(_1948_),
    .B(_1665_));
 sg13g2_a22oi_1 _4404_ (.Y(_1670_),
    .B1(_1669_),
    .B2(net679),
    .A2(net613),
    .A1(net251));
 sg13g2_inv_1 _4405_ (.Y(_0142_),
    .A(net252));
 sg13g2_nor4_2 _4406_ (.A(_1947_),
    .B(_1948_),
    .C(_1949_),
    .Y(_1671_),
    .D(_1662_));
 sg13g2_xnor2_1 _4407_ (.Y(_1672_),
    .A(net251),
    .B(_1668_));
 sg13g2_a22oi_1 _4408_ (.Y(_1673_),
    .B1(_1672_),
    .B2(net677),
    .A2(net611),
    .A1(net350));
 sg13g2_inv_1 _4409_ (.Y(_0143_),
    .A(_1673_));
 sg13g2_nand2_1 _4410_ (.Y(_1674_),
    .A(net223),
    .B(net611));
 sg13g2_xnor2_1 _4411_ (.Y(_1675_),
    .A(\mul_accum[39] ),
    .B(_1671_));
 sg13g2_o21ai_1 _4412_ (.B1(_1674_),
    .Y(_0144_),
    .A1(net694),
    .A2(_1675_));
 sg13g2_a21oi_1 _4413_ (.A1(\mul_accum[39] ),
    .A2(_1671_),
    .Y(_1676_),
    .B1(net223));
 sg13g2_nand3_1 _4414_ (.B(net223),
    .C(_1671_),
    .A(\mul_accum[39] ),
    .Y(_1677_));
 sg13g2_nor2_1 _4415_ (.A(net694),
    .B(_1676_),
    .Y(_1678_));
 sg13g2_a22oi_1 _4416_ (.Y(_1679_),
    .B1(_1677_),
    .B2(_1678_),
    .A2(net610),
    .A1(net309));
 sg13g2_inv_1 _4417_ (.Y(_0145_),
    .A(net310));
 sg13g2_nand4_1 _4418_ (.B(net223),
    .C(net391),
    .A(\mul_accum[39] ),
    .Y(_1680_),
    .D(_1671_));
 sg13g2_a21oi_1 _4419_ (.A1(_1951_),
    .A2(_1677_),
    .Y(_1681_),
    .B1(net694));
 sg13g2_a22oi_1 _4420_ (.Y(_1682_),
    .B1(_1680_),
    .B2(_1681_),
    .A2(net610),
    .A1(net295));
 sg13g2_inv_1 _4421_ (.Y(_0146_),
    .A(net296));
 sg13g2_nor2_1 _4422_ (.A(_1952_),
    .B(_1680_),
    .Y(_1683_));
 sg13g2_xnor2_1 _4423_ (.Y(_1684_),
    .A(net295),
    .B(_1680_));
 sg13g2_a22oi_1 _4424_ (.Y(_1685_),
    .B1(_1684_),
    .B2(net676),
    .A2(net610),
    .A1(net304));
 sg13g2_inv_1 _4425_ (.Y(_0147_),
    .A(_1685_));
 sg13g2_xnor2_1 _4426_ (.Y(_1686_),
    .A(_1953_),
    .B(_1683_));
 sg13g2_a22oi_1 _4427_ (.Y(_1687_),
    .B1(_1686_),
    .B2(net676),
    .A2(net610),
    .A1(net270));
 sg13g2_inv_1 _4428_ (.Y(_0148_),
    .A(net271));
 sg13g2_a21oi_1 _4429_ (.A1(net304),
    .A2(_1683_),
    .Y(_1688_),
    .B1(net270));
 sg13g2_nor4_2 _4430_ (.A(_1952_),
    .B(_1953_),
    .C(_1954_),
    .Y(_1689_),
    .D(_1680_));
 sg13g2_nor2_1 _4431_ (.A(_1688_),
    .B(_1689_),
    .Y(_1690_));
 sg13g2_a22oi_1 _4432_ (.Y(_1691_),
    .B1(_1690_),
    .B2(net676),
    .A2(net614),
    .A1(net307));
 sg13g2_inv_1 _4433_ (.Y(_0149_),
    .A(net308));
 sg13g2_nand2_1 _4434_ (.Y(_1692_),
    .A(net188),
    .B(net612));
 sg13g2_and2_1 _4435_ (.A(net307),
    .B(_1689_),
    .X(_1693_));
 sg13g2_o21ai_1 _4436_ (.B1(net680),
    .Y(_1694_),
    .A1(\mul_accum[45] ),
    .A2(_1689_));
 sg13g2_o21ai_1 _4437_ (.B1(_1692_),
    .Y(_0150_),
    .A1(_1693_),
    .A2(_1694_));
 sg13g2_and2_1 _4438_ (.A(net188),
    .B(_1693_),
    .X(_1695_));
 sg13g2_xor2_1 _4439_ (.B(_1693_),
    .A(net188),
    .X(_1696_));
 sg13g2_a22oi_1 _4440_ (.Y(_1697_),
    .B1(_1696_),
    .B2(net677),
    .A2(net612),
    .A1(net326));
 sg13g2_inv_1 _4441_ (.Y(_0151_),
    .A(_1697_));
 sg13g2_nand4_1 _4442_ (.B(net188),
    .C(\mul_accum[47] ),
    .A(\mul_accum[45] ),
    .Y(_1698_),
    .D(_1689_));
 sg13g2_xor2_1 _4443_ (.B(_1695_),
    .A(\mul_accum[47] ),
    .X(_1699_));
 sg13g2_a22oi_1 _4444_ (.Y(_1700_),
    .B1(_1699_),
    .B2(net677),
    .A2(net612),
    .A1(net297));
 sg13g2_inv_1 _4445_ (.Y(_0152_),
    .A(net298));
 sg13g2_xnor2_1 _4446_ (.Y(_1701_),
    .A(\mul_accum[48] ),
    .B(_1698_));
 sg13g2_a22oi_1 _4447_ (.Y(_1702_),
    .B1(_1701_),
    .B2(net677),
    .A2(net617),
    .A1(net276));
 sg13g2_inv_1 _4448_ (.Y(_0153_),
    .A(net277));
 sg13g2_o21ai_1 _4449_ (.B1(_1956_),
    .Y(_1703_),
    .A1(_1955_),
    .A2(_1698_));
 sg13g2_nand4_1 _4450_ (.B(net297),
    .C(net276),
    .A(\mul_accum[47] ),
    .Y(_1704_),
    .D(_1695_));
 sg13g2_and2_1 _4451_ (.A(net682),
    .B(_1703_),
    .X(_1705_));
 sg13g2_a22oi_1 _4452_ (.Y(_1706_),
    .B1(_1704_),
    .B2(_1705_),
    .A2(net617),
    .A1(net263));
 sg13g2_inv_1 _4453_ (.Y(_0154_),
    .A(net264));
 sg13g2_nor4_2 _4454_ (.A(_1955_),
    .B(_1956_),
    .C(_1957_),
    .Y(_1707_),
    .D(_1698_));
 sg13g2_or2_1 _4455_ (.X(_1708_),
    .B(_1707_),
    .A(net694));
 sg13g2_a21oi_1 _4456_ (.A1(_1957_),
    .A2(_1704_),
    .Y(_1709_),
    .B1(_1708_));
 sg13g2_a21oi_1 _4457_ (.A1(net320),
    .A2(net617),
    .Y(_1710_),
    .B1(_1709_));
 sg13g2_inv_1 _4458_ (.Y(_0155_),
    .A(net321));
 sg13g2_nand2_1 _4459_ (.Y(_1711_),
    .A(net153),
    .B(net617));
 sg13g2_nand2_1 _4460_ (.Y(_1712_),
    .A(\mul_accum[51] ),
    .B(_1707_));
 sg13g2_xnor2_1 _4461_ (.Y(_1713_),
    .A(\mul_accum[51] ),
    .B(_1707_));
 sg13g2_o21ai_1 _4462_ (.B1(_1711_),
    .Y(_0156_),
    .A1(net694),
    .A2(_1713_));
 sg13g2_nand3_1 _4463_ (.B(net153),
    .C(_1707_),
    .A(\mul_accum[51] ),
    .Y(_1714_));
 sg13g2_a21oi_1 _4464_ (.A1(_1958_),
    .A2(_1712_),
    .Y(_1715_),
    .B1(net694));
 sg13g2_a22oi_1 _4465_ (.Y(_1716_),
    .B1(_1714_),
    .B2(_1715_),
    .A2(net615),
    .A1(net291));
 sg13g2_inv_1 _4466_ (.Y(_0157_),
    .A(net292));
 sg13g2_nand2_1 _4467_ (.Y(_1717_),
    .A(net203),
    .B(net615));
 sg13g2_nand4_1 _4468_ (.B(net153),
    .C(\mul_accum[53] ),
    .A(\mul_accum[51] ),
    .Y(_1718_),
    .D(_1707_));
 sg13g2_xor2_1 _4469_ (.B(_1714_),
    .A(\mul_accum[53] ),
    .X(_1719_));
 sg13g2_o21ai_1 _4470_ (.B1(_1717_),
    .Y(_0158_),
    .A1(net694),
    .A2(_1719_));
 sg13g2_xnor2_1 _4471_ (.Y(_1720_),
    .A(net203),
    .B(_1718_));
 sg13g2_a22oi_1 _4472_ (.Y(_1721_),
    .B1(_1720_),
    .B2(net681),
    .A2(net615),
    .A1(net246));
 sg13g2_inv_1 _4473_ (.Y(_0159_),
    .A(net247));
 sg13g2_o21ai_1 _4474_ (.B1(_1960_),
    .Y(_1722_),
    .A1(_1959_),
    .A2(_1718_));
 sg13g2_nor3_1 _4475_ (.A(_1959_),
    .B(_1960_),
    .C(_1718_),
    .Y(_1723_));
 sg13g2_nor2_1 _4476_ (.A(net697),
    .B(_1723_),
    .Y(_1724_));
 sg13g2_a22oi_1 _4477_ (.Y(_1725_),
    .B1(_1722_),
    .B2(_1724_),
    .A2(net615),
    .A1(net274));
 sg13g2_inv_1 _4478_ (.Y(_0160_),
    .A(net275));
 sg13g2_nand2_1 _4479_ (.Y(_1726_),
    .A(net197),
    .B(net616));
 sg13g2_nor4_2 _4480_ (.A(_1959_),
    .B(_1960_),
    .C(_1961_),
    .Y(_1727_),
    .D(_1718_));
 sg13g2_o21ai_1 _4481_ (.B1(net681),
    .Y(_1728_),
    .A1(\mul_accum[56] ),
    .A2(_1723_));
 sg13g2_o21ai_1 _4482_ (.B1(_1726_),
    .Y(_0161_),
    .A1(_1727_),
    .A2(_1728_));
 sg13g2_xor2_1 _4483_ (.B(_1727_),
    .A(net197),
    .X(_1729_));
 sg13g2_a22oi_1 _4484_ (.Y(_1730_),
    .B1(_1729_),
    .B2(net681),
    .A2(net616),
    .A1(net317));
 sg13g2_inv_1 _4485_ (.Y(_0162_),
    .A(_1730_));
 sg13g2_nand2_1 _4486_ (.Y(_1731_),
    .A(net46),
    .B(net616));
 sg13g2_a21oi_1 _4487_ (.A1(\mul_accum[57] ),
    .A2(_1727_),
    .Y(_1732_),
    .B1(\mul_accum[58] ));
 sg13g2_nand3_1 _4488_ (.B(\mul_accum[58] ),
    .C(_1727_),
    .A(\mul_accum[57] ),
    .Y(_1733_));
 sg13g2_nand2_1 _4489_ (.Y(_1734_),
    .A(net681),
    .B(_1733_));
 sg13g2_o21ai_1 _4490_ (.B1(_1731_),
    .Y(_0163_),
    .A1(_1732_),
    .A2(_1734_));
 sg13g2_nand2_1 _4491_ (.Y(_1735_),
    .A(net48),
    .B(net618));
 sg13g2_nand4_1 _4492_ (.B(\mul_accum[58] ),
    .C(\mul_accum[59] ),
    .A(\mul_accum[57] ),
    .Y(_1736_),
    .D(_1727_));
 sg13g2_xor2_1 _4493_ (.B(_1733_),
    .A(net46),
    .X(_1737_));
 sg13g2_o21ai_1 _4494_ (.B1(_1735_),
    .Y(_0164_),
    .A1(net697),
    .A2(_1737_));
 sg13g2_nand2_1 _4495_ (.Y(_1738_),
    .A(net35),
    .B(net618));
 sg13g2_xor2_1 _4496_ (.B(_1736_),
    .A(\mul_accum[60] ),
    .X(_1739_));
 sg13g2_o21ai_1 _4497_ (.B1(_1738_),
    .Y(_0165_),
    .A1(net697),
    .A2(_1739_));
 sg13g2_mux2_1 _4498_ (.A0(\reg_b[0] ),
    .A1(\reg_c[0] ),
    .S(net664),
    .X(_1740_));
 sg13g2_a22oi_1 _4499_ (.Y(_1741_),
    .B1(net605),
    .B2(_1740_),
    .A2(net619),
    .A1(net140));
 sg13g2_inv_1 _4500_ (.Y(_0166_),
    .A(net141));
 sg13g2_nor2b_1 _4501_ (.A(net663),
    .B_N(\reg_b[1] ),
    .Y(_1742_));
 sg13g2_a21oi_1 _4502_ (.A1(\reg_c[1] ),
    .A2(net667),
    .Y(_1743_),
    .B1(_1742_));
 sg13g2_a22oi_1 _4503_ (.Y(_1744_),
    .B1(net619),
    .B2(net52),
    .A2(net686),
    .A1(\mul_b_shift[0] ));
 sg13g2_o21ai_1 _4504_ (.B1(net53),
    .Y(_0167_),
    .A1(net595),
    .A2(_1743_));
 sg13g2_nor2b_1 _4505_ (.A(net667),
    .B_N(\reg_b[2] ),
    .Y(_1745_));
 sg13g2_a21oi_1 _4506_ (.A1(\reg_c[2] ),
    .A2(net667),
    .Y(_1746_),
    .B1(_1745_));
 sg13g2_a22oi_1 _4507_ (.Y(_1747_),
    .B1(net620),
    .B2(net57),
    .A2(net686),
    .A1(net52));
 sg13g2_o21ai_1 _4508_ (.B1(_1747_),
    .Y(_0168_),
    .A1(net594),
    .A2(_1746_));
 sg13g2_nand2b_1 _4509_ (.Y(_1748_),
    .B(net665),
    .A_N(net78));
 sg13g2_o21ai_1 _4510_ (.B1(_1748_),
    .Y(_1749_),
    .A1(\reg_b[3] ),
    .A2(net665));
 sg13g2_a22oi_1 _4511_ (.Y(_1750_),
    .B1(net619),
    .B2(net88),
    .A2(net686),
    .A1(net57));
 sg13g2_o21ai_1 _4512_ (.B1(_1750_),
    .Y(_0169_),
    .A1(net594),
    .A2(_1749_));
 sg13g2_a22oi_1 _4513_ (.Y(_1751_),
    .B1(net619),
    .B2(net82),
    .A2(net687),
    .A1(\mul_b_shift[3] ));
 sg13g2_nand2b_1 _4514_ (.Y(_1752_),
    .B(net667),
    .A_N(\reg_c[4] ));
 sg13g2_o21ai_1 _4515_ (.B1(_1752_),
    .Y(_1753_),
    .A1(\reg_b[4] ),
    .A2(net667));
 sg13g2_o21ai_1 _4516_ (.B1(net83),
    .Y(_0170_),
    .A1(net594),
    .A2(_1753_));
 sg13g2_nand2b_1 _4517_ (.Y(_1754_),
    .B(net666),
    .A_N(\reg_c[5] ));
 sg13g2_o21ai_1 _4518_ (.B1(_1754_),
    .Y(_1755_),
    .A1(\reg_b[5] ),
    .A2(net665));
 sg13g2_a22oi_1 _4519_ (.Y(_1756_),
    .B1(net619),
    .B2(net170),
    .A2(net687),
    .A1(net82));
 sg13g2_o21ai_1 _4520_ (.B1(_1756_),
    .Y(_0171_),
    .A1(net594),
    .A2(_1755_));
 sg13g2_nand2b_1 _4521_ (.Y(_1757_),
    .B(net665),
    .A_N(net113));
 sg13g2_o21ai_1 _4522_ (.B1(_1757_),
    .Y(_1758_),
    .A1(\reg_b[6] ),
    .A2(net665));
 sg13g2_a22oi_1 _4523_ (.Y(_1759_),
    .B1(net619),
    .B2(net163),
    .A2(net687),
    .A1(\mul_b_shift[5] ));
 sg13g2_o21ai_1 _4524_ (.B1(net164),
    .Y(_0172_),
    .A1(net594),
    .A2(_1758_));
 sg13g2_a22oi_1 _4525_ (.Y(_1760_),
    .B1(net620),
    .B2(net85),
    .A2(net686),
    .A1(\mul_b_shift[6] ));
 sg13g2_nand2b_1 _4526_ (.Y(_1761_),
    .B(net665),
    .A_N(\reg_c[7] ));
 sg13g2_o21ai_1 _4527_ (.B1(_1761_),
    .Y(_1762_),
    .A1(\reg_b[7] ),
    .A2(net665));
 sg13g2_o21ai_1 _4528_ (.B1(net86),
    .Y(_0173_),
    .A1(net594),
    .A2(_1762_));
 sg13g2_a22oi_1 _4529_ (.Y(_1763_),
    .B1(net620),
    .B2(net41),
    .A2(net686),
    .A1(\mul_b_shift[7] ));
 sg13g2_nand2b_1 _4530_ (.Y(_1764_),
    .B(net666),
    .A_N(\reg_c[8] ));
 sg13g2_o21ai_1 _4531_ (.B1(_1764_),
    .Y(_1765_),
    .A1(\reg_b[8] ),
    .A2(net665));
 sg13g2_o21ai_1 _4532_ (.B1(net42),
    .Y(_0174_),
    .A1(net594),
    .A2(_1765_));
 sg13g2_nand2b_1 _4533_ (.Y(_1766_),
    .B(net667),
    .A_N(net115));
 sg13g2_o21ai_1 _4534_ (.B1(_1766_),
    .Y(_1767_),
    .A1(\reg_b[9] ),
    .A2(net667));
 sg13g2_a22oi_1 _4535_ (.Y(_1768_),
    .B1(net620),
    .B2(net131),
    .A2(net686),
    .A1(net41));
 sg13g2_o21ai_1 _4536_ (.B1(_1768_),
    .Y(_0175_),
    .A1(net594),
    .A2(_1767_));
 sg13g2_a22oi_1 _4537_ (.Y(_1769_),
    .B1(net620),
    .B2(net128),
    .A2(net687),
    .A1(\mul_b_shift[9] ));
 sg13g2_nand2b_1 _4538_ (.Y(_1770_),
    .B(net666),
    .A_N(\reg_c[10] ));
 sg13g2_o21ai_1 _4539_ (.B1(_1770_),
    .Y(_1771_),
    .A1(\reg_b[10] ),
    .A2(net666));
 sg13g2_o21ai_1 _4540_ (.B1(net129),
    .Y(_0176_),
    .A1(net595),
    .A2(_1771_));
 sg13g2_a22oi_1 _4541_ (.Y(_1772_),
    .B1(net620),
    .B2(net65),
    .A2(net687),
    .A1(\mul_b_shift[10] ));
 sg13g2_nand2b_1 _4542_ (.Y(_1773_),
    .B(net668),
    .A_N(\reg_c[11] ));
 sg13g2_o21ai_1 _4543_ (.B1(_1773_),
    .Y(_1774_),
    .A1(\reg_b[11] ),
    .A2(net674));
 sg13g2_o21ai_1 _4544_ (.B1(net66),
    .Y(_0177_),
    .A1(net595),
    .A2(_1774_));
 sg13g2_a22oi_1 _4545_ (.Y(_1775_),
    .B1(net620),
    .B2(net194),
    .A2(net687),
    .A1(net65));
 sg13g2_nand2b_1 _4546_ (.Y(_1776_),
    .B(net668),
    .A_N(\reg_c[12] ));
 sg13g2_o21ai_1 _4547_ (.B1(_1776_),
    .Y(_1777_),
    .A1(\reg_b[12] ),
    .A2(net668));
 sg13g2_o21ai_1 _4548_ (.B1(_1775_),
    .Y(_0178_),
    .A1(net595),
    .A2(_1777_));
 sg13g2_a22oi_1 _4549_ (.Y(_1778_),
    .B1(net624),
    .B2(net100),
    .A2(net691),
    .A1(\mul_b_shift[12] ));
 sg13g2_nand2b_1 _4550_ (.Y(_1779_),
    .B(net668),
    .A_N(\reg_c[13] ));
 sg13g2_o21ai_1 _4551_ (.B1(_1779_),
    .Y(_1780_),
    .A1(\reg_b[13] ),
    .A2(net668));
 sg13g2_o21ai_1 _4552_ (.B1(net101),
    .Y(_0179_),
    .A1(net595),
    .A2(_1780_));
 sg13g2_nor2b_1 _4553_ (.A(net672),
    .B_N(\reg_b[14] ),
    .Y(_1781_));
 sg13g2_a21oi_1 _4554_ (.A1(\reg_c[14] ),
    .A2(net672),
    .Y(_1782_),
    .B1(_1781_));
 sg13g2_a22oi_1 _4555_ (.Y(_1783_),
    .B1(net624),
    .B2(net111),
    .A2(net691),
    .A1(net100));
 sg13g2_o21ai_1 _4556_ (.B1(_1783_),
    .Y(_0180_),
    .A1(net598),
    .A2(_1782_));
 sg13g2_nor2_1 _4557_ (.A(_1938_),
    .B(net668),
    .Y(_1784_));
 sg13g2_a21oi_1 _4558_ (.A1(\reg_c[15] ),
    .A2(net672),
    .Y(_1785_),
    .B1(_1784_));
 sg13g2_a22oi_1 _4559_ (.Y(_1786_),
    .B1(net624),
    .B2(net73),
    .A2(net691),
    .A1(\mul_b_shift[14] ));
 sg13g2_o21ai_1 _4560_ (.B1(net74),
    .Y(_0181_),
    .A1(net598),
    .A2(_1785_));
 sg13g2_nor2b_1 _4561_ (.A(net672),
    .B_N(\reg_b[16] ),
    .Y(_1787_));
 sg13g2_a21oi_1 _4562_ (.A1(net225),
    .A2(net672),
    .Y(_1788_),
    .B1(_1787_));
 sg13g2_a22oi_1 _4563_ (.Y(_1789_),
    .B1(net624),
    .B2(net238),
    .A2(net691),
    .A1(net73));
 sg13g2_o21ai_1 _4564_ (.B1(_1789_),
    .Y(_0182_),
    .A1(net598),
    .A2(_1788_));
 sg13g2_nor2b_1 _4565_ (.A(net672),
    .B_N(\reg_b[17] ),
    .Y(_1790_));
 sg13g2_a21oi_1 _4566_ (.A1(\reg_c[17] ),
    .A2(net672),
    .Y(_1791_),
    .B1(_1790_));
 sg13g2_a22oi_1 _4567_ (.Y(_1792_),
    .B1(net623),
    .B2(net108),
    .A2(net690),
    .A1(\mul_b_shift[16] ));
 sg13g2_o21ai_1 _4568_ (.B1(net109),
    .Y(_0183_),
    .A1(net598),
    .A2(_1791_));
 sg13g2_nor2b_1 _4569_ (.A(net670),
    .B_N(\reg_b[18] ),
    .Y(_1793_));
 sg13g2_a21oi_1 _4570_ (.A1(\reg_c[18] ),
    .A2(net670),
    .Y(_1794_),
    .B1(_1793_));
 sg13g2_a22oi_1 _4571_ (.Y(_1795_),
    .B1(net623),
    .B2(net121),
    .A2(net690),
    .A1(net108));
 sg13g2_o21ai_1 _4572_ (.B1(_1795_),
    .Y(_0184_),
    .A1(net597),
    .A2(_1794_));
 sg13g2_nor2b_1 _4573_ (.A(net670),
    .B_N(\reg_b[19] ),
    .Y(_1796_));
 sg13g2_a21oi_1 _4574_ (.A1(\reg_c[19] ),
    .A2(net673),
    .Y(_1797_),
    .B1(_1796_));
 sg13g2_a22oi_1 _4575_ (.Y(_1798_),
    .B1(net623),
    .B2(net178),
    .A2(net690),
    .A1(net121));
 sg13g2_o21ai_1 _4576_ (.B1(_1798_),
    .Y(_0185_),
    .A1(net597),
    .A2(_1797_));
 sg13g2_nor2b_1 _4577_ (.A(net671),
    .B_N(\reg_b[20] ),
    .Y(_1799_));
 sg13g2_a21oi_1 _4578_ (.A1(\reg_c[20] ),
    .A2(net670),
    .Y(_1800_),
    .B1(_1799_));
 sg13g2_a22oi_1 _4579_ (.Y(_1801_),
    .B1(net623),
    .B2(net105),
    .A2(net690),
    .A1(\mul_b_shift[19] ));
 sg13g2_o21ai_1 _4580_ (.B1(net106),
    .Y(_0186_),
    .A1(net597),
    .A2(_1800_));
 sg13g2_a22oi_1 _4581_ (.Y(_1802_),
    .B1(net623),
    .B2(net124),
    .A2(net690),
    .A1(net105));
 sg13g2_nand2b_1 _4582_ (.Y(_1803_),
    .B(net670),
    .A_N(\reg_c[21] ));
 sg13g2_o21ai_1 _4583_ (.B1(_1803_),
    .Y(_1804_),
    .A1(\reg_b[21] ),
    .A2(net670));
 sg13g2_o21ai_1 _4584_ (.B1(_1802_),
    .Y(_0187_),
    .A1(net596),
    .A2(_1804_));
 sg13g2_a22oi_1 _4585_ (.Y(_1805_),
    .B1(net622),
    .B2(net90),
    .A2(net690),
    .A1(\mul_b_shift[21] ));
 sg13g2_nand2b_1 _4586_ (.Y(_1806_),
    .B(net671),
    .A_N(\reg_c[22] ));
 sg13g2_o21ai_1 _4587_ (.B1(_1806_),
    .Y(_1807_),
    .A1(\reg_b[22] ),
    .A2(net671));
 sg13g2_o21ai_1 _4588_ (.B1(net91),
    .Y(_0188_),
    .A1(net597),
    .A2(_1807_));
 sg13g2_a22oi_1 _4589_ (.Y(_1808_),
    .B1(net622),
    .B2(net68),
    .A2(net689),
    .A1(\mul_b_shift[22] ));
 sg13g2_nand2b_1 _4590_ (.Y(_1809_),
    .B(net670),
    .A_N(\reg_c[23] ));
 sg13g2_o21ai_1 _4591_ (.B1(_1809_),
    .Y(_1810_),
    .A1(\reg_b[23] ),
    .A2(net670));
 sg13g2_o21ai_1 _4592_ (.B1(net69),
    .Y(_0189_),
    .A1(net597),
    .A2(_1810_));
 sg13g2_nand2b_1 _4593_ (.Y(_1811_),
    .B(net671),
    .A_N(\reg_c[24] ));
 sg13g2_o21ai_1 _4594_ (.B1(_1811_),
    .Y(_1812_),
    .A1(\reg_b[24] ),
    .A2(net671));
 sg13g2_a22oi_1 _4595_ (.Y(_1813_),
    .B1(net623),
    .B2(net144),
    .A2(net689),
    .A1(net68));
 sg13g2_o21ai_1 _4596_ (.B1(_1813_),
    .Y(_0190_),
    .A1(net596),
    .A2(_1812_));
 sg13g2_nor2b_1 _4597_ (.A(net669),
    .B_N(\reg_b[25] ),
    .Y(_1814_));
 sg13g2_a21oi_1 _4598_ (.A1(net177),
    .A2(net669),
    .Y(_1815_),
    .B1(_1814_));
 sg13g2_a22oi_1 _4599_ (.Y(_1816_),
    .B1(net622),
    .B2(net199),
    .A2(net689),
    .A1(net144));
 sg13g2_o21ai_1 _4600_ (.B1(_1816_),
    .Y(_0191_),
    .A1(net596),
    .A2(_1815_));
 sg13g2_nor2b_1 _4601_ (.A(net669),
    .B_N(\reg_b[26] ),
    .Y(_1817_));
 sg13g2_a21oi_1 _4602_ (.A1(\reg_c[26] ),
    .A2(net671),
    .Y(_1818_),
    .B1(_1817_));
 sg13g2_a22oi_1 _4603_ (.Y(_1819_),
    .B1(net622),
    .B2(net174),
    .A2(net689),
    .A1(\mul_b_shift[25] ));
 sg13g2_o21ai_1 _4604_ (.B1(net175),
    .Y(_0192_),
    .A1(net596),
    .A2(_1818_));
 sg13g2_a22oi_1 _4605_ (.Y(_1820_),
    .B1(net622),
    .B2(net117),
    .A2(net689),
    .A1(\mul_b_shift[26] ));
 sg13g2_nand2b_1 _4606_ (.Y(_1821_),
    .B(net671),
    .A_N(\reg_c[27] ));
 sg13g2_o21ai_1 _4607_ (.B1(_1821_),
    .Y(_1822_),
    .A1(\reg_b[27] ),
    .A2(net671));
 sg13g2_o21ai_1 _4608_ (.B1(net118),
    .Y(_0193_),
    .A1(net596),
    .A2(_1822_));
 sg13g2_nand2b_1 _4609_ (.Y(_1823_),
    .B(net669),
    .A_N(\reg_c[28] ));
 sg13g2_o21ai_1 _4610_ (.B1(_1823_),
    .Y(_1824_),
    .A1(\reg_b[28] ),
    .A2(net669));
 sg13g2_a22oi_1 _4611_ (.Y(_1825_),
    .B1(net622),
    .B2(net93),
    .A2(net689),
    .A1(\mul_b_shift[27] ));
 sg13g2_o21ai_1 _4612_ (.B1(net94),
    .Y(_0194_),
    .A1(net596),
    .A2(_1824_));
 sg13g2_a22oi_1 _4613_ (.Y(_1826_),
    .B1(net622),
    .B2(net98),
    .A2(net689),
    .A1(net93));
 sg13g2_nand2b_1 _4614_ (.Y(_1827_),
    .B(net669),
    .A_N(\reg_c[29] ));
 sg13g2_o21ai_1 _4615_ (.B1(_1827_),
    .Y(_1828_),
    .A1(\reg_b[29] ),
    .A2(net669));
 sg13g2_o21ai_1 _4616_ (.B1(_1826_),
    .Y(_0195_),
    .A1(net596),
    .A2(_1828_));
 sg13g2_a22oi_1 _4617_ (.Y(_1829_),
    .B1(net622),
    .B2(net714),
    .A2(net689),
    .A1(net98));
 sg13g2_nand2b_1 _4618_ (.Y(_1830_),
    .B(net673),
    .A_N(net139));
 sg13g2_o21ai_1 _4619_ (.B1(_1830_),
    .Y(_1831_),
    .A1(net283),
    .A2(net669));
 sg13g2_o21ai_1 _4620_ (.B1(_1829_),
    .Y(_0196_),
    .A1(net596),
    .A2(_1831_));
 sg13g2_nor2_1 _4621_ (.A(net32),
    .B(net605),
    .Y(_1832_));
 sg13g2_nor2b_1 _4622_ (.A(net663),
    .B_N(\reg_a[0] ),
    .Y(_1833_));
 sg13g2_a21oi_1 _4623_ (.A1(\reg_b[0] ),
    .A2(net663),
    .Y(_1834_),
    .B1(_1833_));
 sg13g2_a21oi_1 _4624_ (.A1(net605),
    .A2(_1834_),
    .Y(_0197_),
    .B1(_1832_));
 sg13g2_nor2_1 _4625_ (.A(net55),
    .B(net605),
    .Y(_1835_));
 sg13g2_nor2b_1 _4626_ (.A(net663),
    .B_N(\reg_a[1] ),
    .Y(_1836_));
 sg13g2_a21oi_1 _4627_ (.A1(\reg_b[1] ),
    .A2(net663),
    .Y(_1837_),
    .B1(_1836_));
 sg13g2_a21oi_1 _4628_ (.A1(net605),
    .A2(_1837_),
    .Y(_0198_),
    .B1(_1835_));
 sg13g2_nor2_1 _4629_ (.A(net137),
    .B(net605),
    .Y(_1838_));
 sg13g2_nor2b_1 _4630_ (.A(net663),
    .B_N(\reg_a[2] ),
    .Y(_1839_));
 sg13g2_a21oi_1 _4631_ (.A1(\reg_b[2] ),
    .A2(net663),
    .Y(_1840_),
    .B1(_1839_));
 sg13g2_a21oi_1 _4632_ (.A1(net605),
    .A2(_1840_),
    .Y(_0199_),
    .B1(_1838_));
 sg13g2_nor2_1 _4633_ (.A(net185),
    .B(net606),
    .Y(_1841_));
 sg13g2_nor2_1 _4634_ (.A(_1928_),
    .B(net655),
    .Y(_1842_));
 sg13g2_a21oi_1 _4635_ (.A1(\reg_b[3] ),
    .A2(net655),
    .Y(_1843_),
    .B1(_1842_));
 sg13g2_a21oi_1 _4636_ (.A1(net606),
    .A2(_1843_),
    .Y(_0200_),
    .B1(_1841_));
 sg13g2_nor2_1 _4637_ (.A(net161),
    .B(net603),
    .Y(_1844_));
 sg13g2_nor2_1 _4638_ (.A(_1932_),
    .B(net658),
    .Y(_1845_));
 sg13g2_a21oi_1 _4639_ (.A1(\reg_b[4] ),
    .A2(net656),
    .Y(_1846_),
    .B1(_1845_));
 sg13g2_a21oi_1 _4640_ (.A1(net604),
    .A2(_1846_),
    .Y(_0201_),
    .B1(_1844_));
 sg13g2_nor2_1 _4641_ (.A(net168),
    .B(net604),
    .Y(_1847_));
 sg13g2_nor2b_1 _4642_ (.A(net656),
    .B_N(\reg_a[5] ),
    .Y(_1848_));
 sg13g2_a21oi_1 _4643_ (.A1(\reg_b[5] ),
    .A2(net656),
    .Y(_1849_),
    .B1(_1848_));
 sg13g2_a21oi_1 _4644_ (.A1(net604),
    .A2(_1849_),
    .Y(_0202_),
    .B1(_1847_));
 sg13g2_nor2_1 _4645_ (.A(net103),
    .B(net603),
    .Y(_1850_));
 sg13g2_nor2_1 _4646_ (.A(_1934_),
    .B(net658),
    .Y(_1851_));
 sg13g2_a21oi_1 _4647_ (.A1(\reg_b[6] ),
    .A2(net658),
    .Y(_1852_),
    .B1(_1851_));
 sg13g2_a21oi_1 _4648_ (.A1(net603),
    .A2(_1852_),
    .Y(_0203_),
    .B1(_1850_));
 sg13g2_nor2_1 _4649_ (.A(net240),
    .B(net603),
    .Y(_1853_));
 sg13g2_nor2b_1 _4650_ (.A(net655),
    .B_N(\reg_a[7] ),
    .Y(_1854_));
 sg13g2_a21oi_1 _4651_ (.A1(\reg_b[7] ),
    .A2(net655),
    .Y(_1855_),
    .B1(_1854_));
 sg13g2_a21oi_1 _4652_ (.A1(net606),
    .A2(_1855_),
    .Y(_0204_),
    .B1(_1853_));
 sg13g2_nor2_1 _4653_ (.A(net227),
    .B(net606),
    .Y(_1856_));
 sg13g2_nor2b_1 _4654_ (.A(net664),
    .B_N(\reg_a[8] ),
    .Y(_1857_));
 sg13g2_a21oi_1 _4655_ (.A1(\reg_b[8] ),
    .A2(net664),
    .Y(_1858_),
    .B1(_1857_));
 sg13g2_a21oi_1 _4656_ (.A1(net606),
    .A2(_1858_),
    .Y(_0205_),
    .B1(_1856_));
 sg13g2_nor2_1 _4657_ (.A(net192),
    .B(net603),
    .Y(_1859_));
 sg13g2_mux2_1 _4658_ (.A0(_1925_),
    .A1(_1926_),
    .S(net656),
    .X(_1860_));
 sg13g2_a21oi_1 _4659_ (.A1(net603),
    .A2(_1860_),
    .Y(_0206_),
    .B1(_1859_));
 sg13g2_nor2_1 _4660_ (.A(net244),
    .B(net606),
    .Y(_1861_));
 sg13g2_nor2b_1 _4661_ (.A(net664),
    .B_N(\reg_a[10] ),
    .Y(_1862_));
 sg13g2_a21oi_1 _4662_ (.A1(\reg_b[10] ),
    .A2(net663),
    .Y(_1863_),
    .B1(_1862_));
 sg13g2_a21oi_1 _4663_ (.A1(net606),
    .A2(_1863_),
    .Y(_0207_),
    .B1(_1861_));
 sg13g2_nor2_1 _4664_ (.A(net242),
    .B(net603),
    .Y(_1864_));
 sg13g2_nor2_1 _4665_ (.A(_1931_),
    .B(net656),
    .Y(_1865_));
 sg13g2_a21oi_1 _4666_ (.A1(\reg_b[11] ),
    .A2(net655),
    .Y(_1866_),
    .B1(_1865_));
 sg13g2_a21oi_1 _4667_ (.A1(net603),
    .A2(_1866_),
    .Y(_0208_),
    .B1(_1864_));
 sg13g2_nor2_1 _4668_ (.A(net96),
    .B(net600),
    .Y(_1867_));
 sg13g2_nor2b_1 _4669_ (.A(net655),
    .B_N(\reg_a[12] ),
    .Y(_1868_));
 sg13g2_a21oi_1 _4670_ (.A1(\reg_b[12] ),
    .A2(net655),
    .Y(_1869_),
    .B1(_1868_));
 sg13g2_a21oi_1 _4671_ (.A1(net600),
    .A2(_1869_),
    .Y(_0209_),
    .B1(_1867_));
 sg13g2_nor2_1 _4672_ (.A(net50),
    .B(net600),
    .Y(_1870_));
 sg13g2_nor2b_1 _4673_ (.A(net655),
    .B_N(\reg_a[13] ),
    .Y(_1871_));
 sg13g2_a21oi_1 _4674_ (.A1(net730),
    .A2(net656),
    .Y(_1872_),
    .B1(_1871_));
 sg13g2_a21oi_1 _4675_ (.A1(net599),
    .A2(_1872_),
    .Y(_0210_),
    .B1(_1870_));
 sg13g2_nor2_1 _4676_ (.A(net39),
    .B(net599),
    .Y(_1873_));
 sg13g2_nor2_1 _4677_ (.A(_1936_),
    .B(net658),
    .Y(_1874_));
 sg13g2_a21oi_1 _4678_ (.A1(\reg_b[14] ),
    .A2(net658),
    .Y(_1875_),
    .B1(_1874_));
 sg13g2_a21oi_1 _4679_ (.A1(net599),
    .A2(_1875_),
    .Y(_0211_),
    .B1(_1873_));
 sg13g2_nor2_1 _4680_ (.A(net148),
    .B(net599),
    .Y(_1876_));
 sg13g2_mux2_1 _4681_ (.A0(_1937_),
    .A1(_1938_),
    .S(net658),
    .X(_1877_));
 sg13g2_a21oi_1 _4682_ (.A1(net600),
    .A2(_1877_),
    .Y(_0212_),
    .B1(_1876_));
 sg13g2_nor2_1 _4683_ (.A(net59),
    .B(net599),
    .Y(_1878_));
 sg13g2_nor2b_1 _4684_ (.A(net657),
    .B_N(net740),
    .Y(_1879_));
 sg13g2_a21oi_2 _4685_ (.B1(_1879_),
    .Y(_1880_),
    .A2(net657),
    .A1(\reg_b[16] ));
 sg13g2_a21oi_1 _4686_ (.A1(net599),
    .A2(_1880_),
    .Y(_0213_),
    .B1(_1878_));
 sg13g2_nor2_1 _4687_ (.A(net63),
    .B(net599),
    .Y(_1881_));
 sg13g2_nor2_1 _4688_ (.A(_1923_),
    .B(net657),
    .Y(_1882_));
 sg13g2_a21oi_2 _4689_ (.B1(_1882_),
    .Y(_1883_),
    .A2(net657),
    .A1(net729));
 sg13g2_a21oi_1 _4690_ (.A1(net599),
    .A2(_1883_),
    .Y(_0214_),
    .B1(_1881_));
 sg13g2_nor2_1 _4691_ (.A(net44),
    .B(net601),
    .Y(_1884_));
 sg13g2_nor2_1 _4692_ (.A(_1927_),
    .B(net658),
    .Y(_1885_));
 sg13g2_a21oi_2 _4693_ (.B1(_1885_),
    .Y(_1886_),
    .A2(net658),
    .A1(net728));
 sg13g2_a21oi_1 _4694_ (.A1(net601),
    .A2(_1886_),
    .Y(_0215_),
    .B1(_1884_));
 sg13g2_nor2_1 _4695_ (.A(net135),
    .B(net601),
    .Y(_1887_));
 sg13g2_nor2_1 _4696_ (.A(_1930_),
    .B(net661),
    .Y(_1888_));
 sg13g2_a21oi_2 _4697_ (.B1(_1888_),
    .Y(_1889_),
    .A2(net661),
    .A1(net727));
 sg13g2_a21oi_1 _4698_ (.A1(net601),
    .A2(_1889_),
    .Y(_0216_),
    .B1(_1887_));
 sg13g2_nor2_1 _4699_ (.A(net61),
    .B(net601),
    .Y(_1890_));
 sg13g2_nor2_1 _4700_ (.A(_1933_),
    .B(net661),
    .Y(_1891_));
 sg13g2_a21oi_2 _4701_ (.B1(_1891_),
    .Y(_1892_),
    .A2(net661),
    .A1(\reg_b[20] ));
 sg13g2_a21oi_1 _4702_ (.A1(net601),
    .A2(_1892_),
    .Y(_0217_),
    .B1(_1890_));
 sg13g2_nor2_1 _4703_ (.A(net80),
    .B(net601),
    .Y(_1893_));
 sg13g2_nor2b_1 _4704_ (.A(net662),
    .B_N(\reg_a[21] ),
    .Y(_1894_));
 sg13g2_a21oi_2 _4705_ (.B1(_1894_),
    .Y(_1895_),
    .A2(net662),
    .A1(net726));
 sg13g2_a21oi_1 _4706_ (.A1(net601),
    .A2(_1895_),
    .Y(_0218_),
    .B1(_1893_));
 sg13g2_nor2_1 _4707_ (.A(net234),
    .B(net608),
    .Y(_1896_));
 sg13g2_nor2b_1 _4708_ (.A(net662),
    .B_N(\reg_a[22] ),
    .Y(_1897_));
 sg13g2_a21oi_1 _4709_ (.A1(\reg_b[22] ),
    .A2(net662),
    .Y(_1898_),
    .B1(_1897_));
 sg13g2_a21oi_1 _4710_ (.A1(net608),
    .A2(_1898_),
    .Y(_0219_),
    .B1(_1896_));
 sg13g2_nor2_1 _4711_ (.A(net229),
    .B(net602),
    .Y(_1899_));
 sg13g2_nor2b_1 _4712_ (.A(net660),
    .B_N(net736),
    .Y(_1900_));
 sg13g2_a21oi_1 _4713_ (.A1(net725),
    .A2(net660),
    .Y(_1901_),
    .B1(_1900_));
 sg13g2_a21oi_1 _4714_ (.A1(net607),
    .A2(_1901_),
    .Y(_0220_),
    .B1(_1899_));
 sg13g2_nor2_1 _4715_ (.A(net221),
    .B(net608),
    .Y(_1902_));
 sg13g2_nor2b_1 _4716_ (.A(net662),
    .B_N(\reg_a[24] ),
    .Y(_1903_));
 sg13g2_a21oi_1 _4717_ (.A1(\reg_b[24] ),
    .A2(net662),
    .Y(_1904_),
    .B1(_1903_));
 sg13g2_a21oi_1 _4718_ (.A1(net608),
    .A2(_1904_),
    .Y(_0221_),
    .B1(_1902_));
 sg13g2_nor2_1 _4719_ (.A(net214),
    .B(net607),
    .Y(_1905_));
 sg13g2_nor2_1 _4720_ (.A(_1922_),
    .B(net659),
    .Y(_1906_));
 sg13g2_a21oi_1 _4721_ (.A1(net724),
    .A2(net659),
    .Y(_1907_),
    .B1(_1906_));
 sg13g2_a21oi_1 _4722_ (.A1(net607),
    .A2(_1907_),
    .Y(_0222_),
    .B1(_1905_));
 sg13g2_nor2_1 _4723_ (.A(net166),
    .B(net607),
    .Y(_1908_));
 sg13g2_nor2b_1 _4724_ (.A(net659),
    .B_N(net734),
    .Y(_1909_));
 sg13g2_a21oi_1 _4725_ (.A1(\reg_b[26] ),
    .A2(net659),
    .Y(_1910_),
    .B1(_1909_));
 sg13g2_a21oi_1 _4726_ (.A1(net608),
    .A2(_1910_),
    .Y(_0223_),
    .B1(_1908_));
 sg13g2_nor2_1 _4727_ (.A(net210),
    .B(net602),
    .Y(_1911_));
 sg13g2_nor2_1 _4728_ (.A(_1929_),
    .B(net661),
    .Y(_1912_));
 sg13g2_a21oi_1 _4729_ (.A1(net723),
    .A2(net661),
    .Y(_1913_),
    .B1(_1912_));
 sg13g2_a21oi_1 _4730_ (.A1(net602),
    .A2(_1913_),
    .Y(_0224_),
    .B1(_1911_));
 sg13g2_mux2_1 _4731_ (.A0(net733),
    .A1(\reg_b[28] ),
    .S(net659),
    .X(_1914_));
 sg13g2_mux2_1 _4732_ (.A0(net217),
    .A1(_1914_),
    .S(net607),
    .X(_0225_));
 sg13g2_nor2_1 _4733_ (.A(net76),
    .B(net602),
    .Y(_1915_));
 sg13g2_nor2b_1 _4734_ (.A(net659),
    .B_N(net732),
    .Y(_1916_));
 sg13g2_a21oi_1 _4735_ (.A1(net722),
    .A2(net659),
    .Y(_1917_),
    .B1(_1916_));
 sg13g2_a21oi_1 _4736_ (.A1(net607),
    .A2(_1917_),
    .Y(_0226_),
    .B1(_1915_));
 sg13g2_nor2_1 _4737_ (.A(net180),
    .B(net607),
    .Y(_1918_));
 sg13g2_nor2_1 _4738_ (.A(_1935_),
    .B(net659),
    .Y(_1919_));
 sg13g2_a21oi_1 _4739_ (.A1(\reg_b[30] ),
    .A2(net660),
    .Y(_1920_),
    .B1(_1919_));
 sg13g2_a21oi_1 _4740_ (.A1(net607),
    .A2(_1920_),
    .Y(_0227_),
    .B1(_1918_));
 sg13g2_o21ai_1 _4741_ (.B1(net686),
    .Y(_1921_),
    .A1(net705),
    .A2(_2074_));
 sg13g2_inv_1 _4742_ (.Y(_0228_),
    .A(_1921_));
 sg13g2_dfrbpq_2 _4743_ (.RESET_B(net775),
    .D(_0002_),
    .Q(\reg_a[0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _4744_ (.RESET_B(net786),
    .D(_0013_),
    .Q(\reg_a[1] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _4745_ (.RESET_B(net776),
    .D(_0024_),
    .Q(\reg_a[2] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _4746_ (.RESET_B(net786),
    .D(_0027_),
    .Q(\reg_a[3] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _4747_ (.RESET_B(net773),
    .D(_0028_),
    .Q(\reg_a[4] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _4748_ (.RESET_B(net773),
    .D(_0029_),
    .Q(\reg_a[5] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _4749_ (.RESET_B(net775),
    .D(_0030_),
    .Q(\reg_a[6] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _4750_ (.RESET_B(net775),
    .D(_0031_),
    .Q(\reg_a[7] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _4751_ (.RESET_B(net776),
    .D(_0032_),
    .Q(\reg_a[8] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _4752_ (.RESET_B(net772),
    .D(_0033_),
    .Q(\reg_a[9] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _4753_ (.RESET_B(net772),
    .D(_0003_),
    .Q(\reg_a[10] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _4754_ (.RESET_B(net775),
    .D(_0004_),
    .Q(\reg_a[11] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _4755_ (.RESET_B(net775),
    .D(_0005_),
    .Q(\reg_a[12] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _4756_ (.RESET_B(net781),
    .D(_0006_),
    .Q(\reg_a[13] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _4757_ (.RESET_B(net775),
    .D(_0007_),
    .Q(\reg_a[14] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _4758_ (.RESET_B(net781),
    .D(_0008_),
    .Q(\reg_a[15] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _4759_ (.RESET_B(net781),
    .D(_0009_),
    .Q(\reg_a[16] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _4760_ (.RESET_B(net781),
    .D(_0010_),
    .Q(\reg_a[17] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _4761_ (.RESET_B(net785),
    .D(_0011_),
    .Q(\reg_a[18] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _4762_ (.RESET_B(net785),
    .D(_0012_),
    .Q(\reg_a[19] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _4763_ (.RESET_B(net781),
    .D(_0014_),
    .Q(\reg_a[20] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _4764_ (.RESET_B(net781),
    .D(_0015_),
    .Q(\reg_a[21] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _4765_ (.RESET_B(net782),
    .D(_0016_),
    .Q(\reg_a[22] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _4766_ (.RESET_B(net781),
    .D(_0017_),
    .Q(\reg_a[23] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _4767_ (.RESET_B(net782),
    .D(_0018_),
    .Q(\reg_a[24] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _4768_ (.RESET_B(net783),
    .D(_0019_),
    .Q(\reg_a[25] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _4769_ (.RESET_B(net782),
    .D(_0020_),
    .Q(\reg_a[26] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _4770_ (.RESET_B(net783),
    .D(_0021_),
    .Q(\reg_a[27] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _4771_ (.RESET_B(net782),
    .D(_0022_),
    .Q(\reg_a[28] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _4772_ (.RESET_B(net782),
    .D(_0023_),
    .Q(\reg_a[29] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _4773_ (.RESET_B(net783),
    .D(_0025_),
    .Q(\reg_a[30] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _4774_ (.RESET_B(net796),
    .D(_0026_),
    .Q(\reg_a[31] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _4775_ (.RESET_B(net790),
    .D(net250),
    .Q(\reg_b[0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _4776_ (.RESET_B(net790),
    .D(net257),
    .Q(\reg_b[1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _4777_ (.RESET_B(net790),
    .D(net261),
    .Q(\reg_b[2] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _4778_ (.RESET_B(net791),
    .D(net323),
    .Q(\reg_b[3] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _4779_ (.RESET_B(net790),
    .D(net319),
    .Q(\reg_b[4] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _4780_ (.RESET_B(net791),
    .D(net359),
    .Q(\reg_b[5] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _4781_ (.RESET_B(net793),
    .D(net346),
    .Q(\reg_b[6] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _4782_ (.RESET_B(net793),
    .D(_0063_),
    .Q(\reg_b[7] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _4783_ (.RESET_B(net795),
    .D(net312),
    .Q(\reg_b[8] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _4784_ (.RESET_B(net795),
    .D(net374),
    .Q(\reg_b[9] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _4785_ (.RESET_B(net794),
    .D(net328),
    .Q(\reg_b[10] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _4786_ (.RESET_B(net794),
    .D(net344),
    .Q(\reg_b[11] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _4787_ (.RESET_B(net798),
    .D(net339),
    .Q(\reg_b[12] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _4788_ (.RESET_B(net798),
    .D(net366),
    .Q(\reg_b[13] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _4789_ (.RESET_B(net800),
    .D(net354),
    .Q(\reg_b[14] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _4790_ (.RESET_B(net798),
    .D(_0040_),
    .Q(\reg_b[15] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _4791_ (.RESET_B(net800),
    .D(net341),
    .Q(\reg_b[16] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _4792_ (.RESET_B(net800),
    .D(_0042_),
    .Q(\reg_b[17] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _4793_ (.RESET_B(net799),
    .D(_0043_),
    .Q(\reg_b[18] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _4794_ (.RESET_B(net803),
    .D(_0044_),
    .Q(\reg_b[19] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _4795_ (.RESET_B(net801),
    .D(_0046_),
    .Q(\reg_b[20] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _4796_ (.RESET_B(net801),
    .D(_0047_),
    .Q(\reg_b[21] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _4797_ (.RESET_B(net801),
    .D(_0048_),
    .Q(\reg_b[22] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _4798_ (.RESET_B(net803),
    .D(_0049_),
    .Q(\reg_b[23] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _4799_ (.RESET_B(net796),
    .D(_0050_),
    .Q(\reg_b[24] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _4800_ (.RESET_B(net796),
    .D(_0051_),
    .Q(\reg_b[25] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _4801_ (.RESET_B(net796),
    .D(_0052_),
    .Q(\reg_b[26] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _4802_ (.RESET_B(net796),
    .D(_0053_),
    .Q(\reg_b[27] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _4803_ (.RESET_B(net796),
    .D(_0054_),
    .Q(\reg_b[28] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _4804_ (.RESET_B(net796),
    .D(_0055_),
    .Q(\reg_b[29] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _4805_ (.RESET_B(net796),
    .D(_0057_),
    .Q(\reg_b[30] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _4806_ (.RESET_B(net801),
    .D(_0058_),
    .Q(\reg_b[31] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _4807_ (.RESET_B(net795),
    .D(net160),
    .Q(\reg_c[0] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _4808_ (.RESET_B(net795),
    .D(net72),
    .Q(\reg_c[1] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _4809_ (.RESET_B(net793),
    .D(net173),
    .Q(\reg_c[2] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _4810_ (.RESET_B(net793),
    .D(net79),
    .Q(\reg_c[3] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _4811_ (.RESET_B(net793),
    .D(net127),
    .Q(\reg_c[4] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _4812_ (.RESET_B(net793),
    .D(_0093_),
    .Q(\reg_c[5] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _4813_ (.RESET_B(net793),
    .D(net114),
    .Q(\reg_c[6] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _4814_ (.RESET_B(net794),
    .D(net143),
    .Q(\reg_c[7] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _4815_ (.RESET_B(net794),
    .D(_0096_),
    .Q(\reg_c[8] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _4816_ (.RESET_B(net795),
    .D(net116),
    .Q(\reg_c[9] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _4817_ (.RESET_B(net794),
    .D(_0067_),
    .Q(\reg_c[10] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _4818_ (.RESET_B(net794),
    .D(_0068_),
    .Q(\reg_c[11] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _4819_ (.RESET_B(net798),
    .D(_0069_),
    .Q(\reg_c[12] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _4820_ (.RESET_B(net798),
    .D(net183),
    .Q(\reg_c[13] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _4821_ (.RESET_B(net798),
    .D(_0071_),
    .Q(\reg_c[14] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _4822_ (.RESET_B(net799),
    .D(_0072_),
    .Q(\reg_c[15] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _4823_ (.RESET_B(net799),
    .D(net226),
    .Q(\reg_c[16] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _4824_ (.RESET_B(net800),
    .D(_0074_),
    .Q(\reg_c[17] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _4825_ (.RESET_B(net803),
    .D(_0075_),
    .Q(\reg_c[18] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _4826_ (.RESET_B(net803),
    .D(net213),
    .Q(\reg_c[19] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _4827_ (.RESET_B(net804),
    .D(_0078_),
    .Q(\reg_c[20] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _4828_ (.RESET_B(net804),
    .D(_0079_),
    .Q(\reg_c[21] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _4829_ (.RESET_B(net803),
    .D(_0080_),
    .Q(\reg_c[22] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _4830_ (.RESET_B(net803),
    .D(net147),
    .Q(\reg_c[23] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _4831_ (.RESET_B(net804),
    .D(_0082_),
    .Q(\reg_c[24] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _4832_ (.RESET_B(net802),
    .D(_0083_),
    .Q(\reg_c[25] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _4833_ (.RESET_B(net804),
    .D(_0084_),
    .Q(\reg_c[26] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _4834_ (.RESET_B(net804),
    .D(_0085_),
    .Q(\reg_c[27] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _4835_ (.RESET_B(net802),
    .D(_0086_),
    .Q(\reg_c[28] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _4836_ (.RESET_B(net802),
    .D(_0087_),
    .Q(\reg_c[29] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _4837_ (.RESET_B(net801),
    .D(_0089_),
    .Q(\reg_c[30] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _4838_ (.RESET_B(net803),
    .D(_0090_),
    .Q(\reg_c[31] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _4839_ (.RESET_B(net799),
    .D(_0000_),
    .Q(\read_counter[0] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _4840_ (.RESET_B(net799),
    .D(_0001_),
    .Q(\read_counter[1] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _4841_ (.RESET_B(net781),
    .D(_0098_),
    .Q(mac_mode),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _4842_ (.RESET_B(net789),
    .D(_0099_),
    .Q(\mul_counter[0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _4843_ (.RESET_B(net789),
    .D(_0100_),
    .Q(\mul_counter[1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _4844_ (.RESET_B(net789),
    .D(net31),
    .Q(\mul_counter[2] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _4845_ (.RESET_B(net789),
    .D(net29),
    .Q(\mul_counter[3] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _4846_ (.RESET_B(net789),
    .D(_0103_),
    .Q(\mul_counter[4] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _4847_ (.RESET_B(net787),
    .D(_0104_),
    .Q(\mul_accum[0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _4848_ (.RESET_B(net787),
    .D(_0105_),
    .Q(\mul_accum[1] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _4849_ (.RESET_B(net787),
    .D(net335),
    .Q(\mul_accum[2] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _4850_ (.RESET_B(net786),
    .D(net332),
    .Q(\mul_accum[3] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _4851_ (.RESET_B(net786),
    .D(net330),
    .Q(\mul_accum[4] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _4852_ (.RESET_B(net786),
    .D(_0109_),
    .Q(\mul_accum[5] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _4853_ (.RESET_B(net774),
    .D(net337),
    .Q(\mul_accum[6] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _4854_ (.RESET_B(net773),
    .D(net208),
    .Q(\mul_accum[7] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _4855_ (.RESET_B(net769),
    .D(net316),
    .Q(\mul_accum[8] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _4856_ (.RESET_B(net769),
    .D(_0113_),
    .Q(\mul_accum[9] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _4857_ (.RESET_B(net769),
    .D(net325),
    .Q(\mul_accum[10] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _4858_ (.RESET_B(net768),
    .D(net191),
    .Q(\mul_accum[11] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _4859_ (.RESET_B(net768),
    .D(_0116_),
    .Q(\mul_accum[12] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _4860_ (.RESET_B(net768),
    .D(_0117_),
    .Q(\mul_accum[13] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _4861_ (.RESET_B(net770),
    .D(net280),
    .Q(\mul_accum[14] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _4862_ (.RESET_B(net770),
    .D(net134),
    .Q(\mul_accum[15] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _4863_ (.RESET_B(net771),
    .D(_0120_),
    .Q(\mul_accum[16] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _4864_ (.RESET_B(net771),
    .D(_0121_),
    .Q(\mul_accum[17] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _4865_ (.RESET_B(net777),
    .D(net288),
    .Q(\mul_accum[18] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _4866_ (.RESET_B(net777),
    .D(net273),
    .Q(\mul_accum[19] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _4867_ (.RESET_B(net780),
    .D(_0124_),
    .Q(\mul_accum[20] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _4868_ (.RESET_B(net778),
    .D(net300),
    .Q(\mul_accum[21] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _4869_ (.RESET_B(net778),
    .D(net158),
    .Q(\mul_accum[22] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _4870_ (.RESET_B(net779),
    .D(_0127_),
    .Q(\mul_accum[23] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _4871_ (.RESET_B(net778),
    .D(net306),
    .Q(\mul_accum[24] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _4872_ (.RESET_B(net778),
    .D(net282),
    .Q(\mul_accum[25] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _4873_ (.RESET_B(net779),
    .D(_0130_),
    .Q(\mul_accum[26] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _4874_ (.RESET_B(net779),
    .D(net314),
    .Q(\mul_accum[27] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _4875_ (.RESET_B(net782),
    .D(net266),
    .Q(\mul_accum[28] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _4876_ (.RESET_B(net782),
    .D(net259),
    .Q(\mul_accum[29] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _4877_ (.RESET_B(net784),
    .D(net362),
    .Q(\mul_accum[30] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _4878_ (.RESET_B(net773),
    .D(_0135_),
    .Q(\mul_accum[31] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _4879_ (.RESET_B(net773),
    .D(net206),
    .Q(\mul_accum[32] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _4880_ (.RESET_B(net774),
    .D(_0137_),
    .Q(\mul_accum[33] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _4881_ (.RESET_B(net774),
    .D(net152),
    .Q(\mul_accum[34] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _4882_ (.RESET_B(net774),
    .D(_0139_),
    .Q(\mul_accum[35] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _4883_ (.RESET_B(net773),
    .D(_0140_),
    .Q(\mul_accum[36] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _4884_ (.RESET_B(net773),
    .D(_0141_),
    .Q(\mul_accum[37] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _4885_ (.RESET_B(net773),
    .D(_0142_),
    .Q(\mul_accum[38] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _4886_ (.RESET_B(net769),
    .D(_0143_),
    .Q(\mul_accum[39] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _4887_ (.RESET_B(net769),
    .D(net224),
    .Q(\mul_accum[40] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _4888_ (.RESET_B(net768),
    .D(_0145_),
    .Q(\mul_accum[41] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _4889_ (.RESET_B(net768),
    .D(_0146_),
    .Q(\mul_accum[42] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _4890_ (.RESET_B(net768),
    .D(_0147_),
    .Q(\mul_accum[43] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _4891_ (.RESET_B(net768),
    .D(_0148_),
    .Q(\mul_accum[44] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _4892_ (.RESET_B(net770),
    .D(_0149_),
    .Q(\mul_accum[45] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _4893_ (.RESET_B(net770),
    .D(net189),
    .Q(\mul_accum[46] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _4894_ (.RESET_B(net771),
    .D(_0151_),
    .Q(\mul_accum[47] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _4895_ (.RESET_B(net771),
    .D(_0152_),
    .Q(\mul_accum[48] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _4896_ (.RESET_B(net777),
    .D(_0153_),
    .Q(\mul_accum[49] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _4897_ (.RESET_B(net777),
    .D(_0154_),
    .Q(\mul_accum[50] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _4898_ (.RESET_B(net777),
    .D(_0155_),
    .Q(\mul_accum[51] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _4899_ (.RESET_B(net780),
    .D(net154),
    .Q(\mul_accum[52] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _4900_ (.RESET_B(net778),
    .D(_0157_),
    .Q(\mul_accum[53] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _4901_ (.RESET_B(net778),
    .D(net204),
    .Q(\mul_accum[54] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _4902_ (.RESET_B(net778),
    .D(_0159_),
    .Q(\mul_accum[55] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _4903_ (.RESET_B(net778),
    .D(_0160_),
    .Q(\mul_accum[56] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _4904_ (.RESET_B(net779),
    .D(net198),
    .Q(\mul_accum[57] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _4905_ (.RESET_B(net779),
    .D(_0162_),
    .Q(\mul_accum[58] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _4906_ (.RESET_B(net779),
    .D(net47),
    .Q(\mul_accum[59] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _4907_ (.RESET_B(net784),
    .D(net49),
    .Q(\mul_accum[60] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _4908_ (.RESET_B(net782),
    .D(net36),
    .Q(\mul_accum[61] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _4909_ (.RESET_B(net790),
    .D(_0166_),
    .Q(\mul_b_shift[0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _4910_ (.RESET_B(net790),
    .D(net54),
    .Q(\mul_b_shift[1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _4911_ (.RESET_B(net791),
    .D(net58),
    .Q(\mul_b_shift[2] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _4912_ (.RESET_B(net791),
    .D(net89),
    .Q(\mul_b_shift[3] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _4913_ (.RESET_B(net791),
    .D(net84),
    .Q(\mul_b_shift[4] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _4914_ (.RESET_B(net791),
    .D(net171),
    .Q(\mul_b_shift[5] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _4915_ (.RESET_B(net791),
    .D(net165),
    .Q(\mul_b_shift[6] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _4916_ (.RESET_B(net791),
    .D(net87),
    .Q(\mul_b_shift[7] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _4917_ (.RESET_B(net792),
    .D(net43),
    .Q(\mul_b_shift[8] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _4918_ (.RESET_B(net792),
    .D(net132),
    .Q(\mul_b_shift[9] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _4919_ (.RESET_B(net793),
    .D(net130),
    .Q(\mul_b_shift[10] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _4920_ (.RESET_B(net794),
    .D(net67),
    .Q(\mul_b_shift[11] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _4921_ (.RESET_B(net798),
    .D(net195),
    .Q(\mul_b_shift[12] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _4922_ (.RESET_B(net798),
    .D(net102),
    .Q(\mul_b_shift[13] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _4923_ (.RESET_B(net799),
    .D(net112),
    .Q(\mul_b_shift[14] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _4924_ (.RESET_B(net799),
    .D(net75),
    .Q(\mul_b_shift[15] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _4925_ (.RESET_B(net799),
    .D(net239),
    .Q(\mul_b_shift[16] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _4926_ (.RESET_B(net805),
    .D(net110),
    .Q(\mul_b_shift[17] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _4927_ (.RESET_B(net803),
    .D(net122),
    .Q(\mul_b_shift[18] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _4928_ (.RESET_B(net805),
    .D(net179),
    .Q(\mul_b_shift[19] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _4929_ (.RESET_B(net805),
    .D(net107),
    .Q(\mul_b_shift[20] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _4930_ (.RESET_B(net805),
    .D(net125),
    .Q(\mul_b_shift[21] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _4931_ (.RESET_B(net804),
    .D(net92),
    .Q(\mul_b_shift[22] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _4932_ (.RESET_B(net804),
    .D(net70),
    .Q(\mul_b_shift[23] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _4933_ (.RESET_B(net804),
    .D(net145),
    .Q(\mul_b_shift[24] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _4934_ (.RESET_B(net802),
    .D(net200),
    .Q(\mul_b_shift[25] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _4935_ (.RESET_B(net802),
    .D(net176),
    .Q(\mul_b_shift[26] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _4936_ (.RESET_B(net801),
    .D(net119),
    .Q(\mul_b_shift[27] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _4937_ (.RESET_B(net801),
    .D(net95),
    .Q(\mul_b_shift[28] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _4938_ (.RESET_B(net801),
    .D(net99),
    .Q(\mul_b_shift[29] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _4939_ (.RESET_B(net797),
    .D(net284),
    .Q(\mul_b_shift[30] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _4940_ (.RESET_B(net789),
    .D(net33),
    .Q(\mul_operand_r[0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _4941_ (.RESET_B(net789),
    .D(net56),
    .Q(\mul_operand_r[1] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _4942_ (.RESET_B(net787),
    .D(net138),
    .Q(\mul_operand_r[2] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _4943_ (.RESET_B(net787),
    .D(net186),
    .Q(\mul_operand_r[3] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _4944_ (.RESET_B(net786),
    .D(net162),
    .Q(\mul_operand_r[4] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _4945_ (.RESET_B(net786),
    .D(net169),
    .Q(\mul_operand_r[5] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _4946_ (.RESET_B(net786),
    .D(net104),
    .Q(\mul_operand_r[6] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _4947_ (.RESET_B(net787),
    .D(net241),
    .Q(\mul_operand_r[7] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _4948_ (.RESET_B(net787),
    .D(net228),
    .Q(\mul_operand_r[8] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _4949_ (.RESET_B(net788),
    .D(net193),
    .Q(\mul_operand_r[9] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _4950_ (.RESET_B(net787),
    .D(net245),
    .Q(\mul_operand_r[10] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _4951_ (.RESET_B(net788),
    .D(net243),
    .Q(\mul_operand_r[11] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _4952_ (.RESET_B(net769),
    .D(net97),
    .Q(\mul_operand_r[12] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _4953_ (.RESET_B(net768),
    .D(net51),
    .Q(\mul_operand_r[13] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _4954_ (.RESET_B(net770),
    .D(net40),
    .Q(\mul_operand_r[14] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _4955_ (.RESET_B(net770),
    .D(net149),
    .Q(\mul_operand_r[15] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _4956_ (.RESET_B(net770),
    .D(net60),
    .Q(\mul_operand_r[16] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _4957_ (.RESET_B(net770),
    .D(net64),
    .Q(\mul_operand_r[17] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _4958_ (.RESET_B(net777),
    .D(net45),
    .Q(\mul_operand_r[18] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _4959_ (.RESET_B(net777),
    .D(net136),
    .Q(\mul_operand_r[19] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _4960_ (.RESET_B(net777),
    .D(net62),
    .Q(\mul_operand_r[20] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _4961_ (.RESET_B(net779),
    .D(net81),
    .Q(\mul_operand_r[21] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _4962_ (.RESET_B(net797),
    .D(net235),
    .Q(\mul_operand_r[22] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _4963_ (.RESET_B(net784),
    .D(net230),
    .Q(\mul_operand_r[23] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _4964_ (.RESET_B(net797),
    .D(net222),
    .Q(\mul_operand_r[24] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _4965_ (.RESET_B(net783),
    .D(net215),
    .Q(\mul_operand_r[25] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _4966_ (.RESET_B(net797),
    .D(net167),
    .Q(\mul_operand_r[26] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _4967_ (.RESET_B(net783),
    .D(net211),
    .Q(\mul_operand_r[27] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _4968_ (.RESET_B(net783),
    .D(net218),
    .Q(\mul_operand_r[28] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _4969_ (.RESET_B(net783),
    .D(net77),
    .Q(\mul_operand_r[29] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _4970_ (.RESET_B(net783),
    .D(net181),
    .Q(\mul_operand_r[30] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _4971_ (.RESET_B(net789),
    .D(_0228_),
    .Q(reducing),
    .CLK(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_brmurrell3_m31_accel_13 (.L_LO(net13));
 sg13g2_tielo tt_um_brmurrell3_m31_accel_14 (.L_LO(net14));
 sg13g2_tielo tt_um_brmurrell3_m31_accel_15 (.L_LO(net15));
 sg13g2_tielo tt_um_brmurrell3_m31_accel_16 (.L_LO(net16));
 sg13g2_tielo tt_um_brmurrell3_m31_accel_17 (.L_LO(net17));
 sg13g2_tielo tt_um_brmurrell3_m31_accel_18 (.L_LO(net18));
 sg13g2_tielo tt_um_brmurrell3_m31_accel_19 (.L_LO(net19));
 sg13g2_tielo tt_um_brmurrell3_m31_accel_20 (.L_LO(net20));
 sg13g2_tielo tt_um_brmurrell3_m31_accel_21 (.L_LO(net21));
 sg13g2_tielo tt_um_brmurrell3_m31_accel_22 (.L_LO(net22));
 sg13g2_tielo tt_um_brmurrell3_m31_accel_23 (.L_LO(net23));
 sg13g2_tielo tt_um_brmurrell3_m31_accel_24 (.L_LO(net24));
 sg13g2_tielo tt_um_brmurrell3_m31_accel_25 (.L_LO(net25));
 sg13g2_tiehi tt_um_brmurrell3_m31_accel_26 (.L_HI(net26));
 sg13g2_buf_1 _4987_ (.A(busy),
    .X(uio_out[0]));
 sg13g2_buf_8 fanout541 (.A(_1135_),
    .X(net541));
 sg13g2_buf_1 fanout542 (.A(_1135_),
    .X(net542));
 sg13g2_buf_8 fanout543 (.A(net544),
    .X(net543));
 sg13g2_buf_8 fanout544 (.A(_1132_),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(net546),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(_1132_),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(net548),
    .X(net547));
 sg13g2_buf_1 fanout548 (.A(net550),
    .X(net548));
 sg13g2_buf_8 fanout549 (.A(net550),
    .X(net549));
 sg13g2_buf_1 fanout550 (.A(_0933_),
    .X(net550));
 sg13g2_buf_8 fanout551 (.A(_0663_),
    .X(net551));
 sg13g2_buf_1 fanout552 (.A(_0663_),
    .X(net552));
 sg13g2_buf_8 fanout553 (.A(net554),
    .X(net553));
 sg13g2_buf_8 fanout554 (.A(net555),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(net556),
    .X(net555));
 sg13g2_buf_1 fanout556 (.A(net557),
    .X(net556));
 sg13g2_buf_8 fanout557 (.A(net559),
    .X(net557));
 sg13g2_buf_8 fanout558 (.A(net559),
    .X(net558));
 sg13g2_buf_8 fanout559 (.A(_0357_),
    .X(net559));
 sg13g2_buf_8 fanout560 (.A(_0347_),
    .X(net560));
 sg13g2_buf_8 fanout561 (.A(_0309_),
    .X(net561));
 sg13g2_buf_8 fanout562 (.A(_0249_),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(_0249_),
    .X(net563));
 sg13g2_buf_8 fanout564 (.A(_0256_),
    .X(net564));
 sg13g2_buf_8 fanout565 (.A(net566),
    .X(net565));
 sg13g2_buf_8 fanout566 (.A(_2082_),
    .X(net566));
 sg13g2_buf_8 fanout567 (.A(net569),
    .X(net567));
 sg13g2_buf_1 fanout568 (.A(net569),
    .X(net568));
 sg13g2_buf_8 fanout569 (.A(_2082_),
    .X(net569));
 sg13g2_buf_8 fanout570 (.A(net573),
    .X(net570));
 sg13g2_buf_8 fanout571 (.A(net572),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(net573),
    .X(net572));
 sg13g2_buf_8 fanout573 (.A(_0671_),
    .X(net573));
 sg13g2_buf_8 fanout574 (.A(_0670_),
    .X(net574));
 sg13g2_buf_1 fanout575 (.A(_0670_),
    .X(net575));
 sg13g2_buf_8 fanout576 (.A(net578),
    .X(net576));
 sg13g2_buf_1 fanout577 (.A(net578),
    .X(net577));
 sg13g2_buf_8 fanout578 (.A(_0670_),
    .X(net578));
 sg13g2_buf_8 fanout579 (.A(net580),
    .X(net579));
 sg13g2_buf_8 fanout580 (.A(_2151_),
    .X(net580));
 sg13g2_buf_8 fanout581 (.A(net582),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(net583),
    .X(net582));
 sg13g2_buf_8 fanout583 (.A(_2151_),
    .X(net583));
 sg13g2_buf_8 fanout584 (.A(_2079_),
    .X(net584));
 sg13g2_buf_1 fanout585 (.A(_2079_),
    .X(net585));
 sg13g2_buf_8 fanout586 (.A(net588),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(net588),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(_2079_),
    .X(net588));
 sg13g2_buf_8 fanout589 (.A(net593),
    .X(net589));
 sg13g2_buf_1 fanout590 (.A(net593),
    .X(net590));
 sg13g2_buf_8 fanout591 (.A(net593),
    .X(net591));
 sg13g2_buf_8 fanout592 (.A(net593),
    .X(net592));
 sg13g2_buf_8 fanout593 (.A(_2078_),
    .X(net593));
 sg13g2_buf_8 fanout594 (.A(net595),
    .X(net594));
 sg13g2_buf_8 fanout595 (.A(_1424_),
    .X(net595));
 sg13g2_buf_8 fanout596 (.A(net598),
    .X(net596));
 sg13g2_buf_1 fanout597 (.A(net598),
    .X(net597));
 sg13g2_buf_8 fanout598 (.A(_1424_),
    .X(net598));
 sg13g2_buf_8 fanout599 (.A(net600),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(net609),
    .X(net600));
 sg13g2_buf_8 fanout601 (.A(net609),
    .X(net601));
 sg13g2_buf_1 fanout602 (.A(net609),
    .X(net602));
 sg13g2_buf_8 fanout603 (.A(net604),
    .X(net603));
 sg13g2_buf_1 fanout604 (.A(net609),
    .X(net604));
 sg13g2_buf_8 fanout605 (.A(net606),
    .X(net605));
 sg13g2_buf_8 fanout606 (.A(net609),
    .X(net606));
 sg13g2_buf_8 fanout607 (.A(net608),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(net609),
    .X(net608));
 sg13g2_buf_8 fanout609 (.A(_1423_),
    .X(net609));
 sg13g2_buf_8 fanout610 (.A(net612),
    .X(net610));
 sg13g2_buf_1 fanout611 (.A(net612),
    .X(net611));
 sg13g2_buf_8 fanout612 (.A(net614),
    .X(net612));
 sg13g2_buf_8 fanout613 (.A(net614),
    .X(net613));
 sg13g2_buf_8 fanout614 (.A(net625),
    .X(net614));
 sg13g2_buf_8 fanout615 (.A(net616),
    .X(net615));
 sg13g2_buf_8 fanout616 (.A(net617),
    .X(net616));
 sg13g2_buf_8 fanout617 (.A(net618),
    .X(net617));
 sg13g2_buf_8 fanout618 (.A(net625),
    .X(net618));
 sg13g2_buf_8 fanout619 (.A(net620),
    .X(net619));
 sg13g2_buf_8 fanout620 (.A(net621),
    .X(net620));
 sg13g2_buf_8 fanout621 (.A(net625),
    .X(net621));
 sg13g2_buf_8 fanout622 (.A(net624),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(net624),
    .X(net623));
 sg13g2_buf_8 fanout624 (.A(net625),
    .X(net624));
 sg13g2_buf_8 fanout625 (.A(_1419_),
    .X(net625));
 sg13g2_buf_8 fanout626 (.A(net627),
    .X(net626));
 sg13g2_buf_8 fanout627 (.A(net629),
    .X(net627));
 sg13g2_buf_8 fanout628 (.A(net629),
    .X(net628));
 sg13g2_buf_8 fanout629 (.A(_0679_),
    .X(net629));
 sg13g2_buf_8 fanout630 (.A(_0678_),
    .X(net630));
 sg13g2_buf_8 fanout631 (.A(_0678_),
    .X(net631));
 sg13g2_buf_8 fanout632 (.A(net633),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(_0678_),
    .X(net633));
 sg13g2_buf_8 fanout634 (.A(busy),
    .X(net634));
 sg13g2_buf_8 fanout635 (.A(net636),
    .X(net635));
 sg13g2_buf_8 fanout636 (.A(net638),
    .X(net636));
 sg13g2_buf_8 fanout637 (.A(net638),
    .X(net637));
 sg13g2_buf_8 fanout638 (.A(_0667_),
    .X(net638));
 sg13g2_buf_8 fanout639 (.A(_0666_),
    .X(net639));
 sg13g2_buf_8 fanout640 (.A(net643),
    .X(net640));
 sg13g2_buf_1 fanout641 (.A(net643),
    .X(net641));
 sg13g2_buf_8 fanout642 (.A(net643),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(net644),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(net651),
    .X(net644));
 sg13g2_buf_8 fanout645 (.A(net647),
    .X(net645));
 sg13g2_buf_1 fanout646 (.A(net647),
    .X(net646));
 sg13g2_buf_1 fanout647 (.A(net651),
    .X(net647));
 sg13g2_buf_8 fanout648 (.A(net649),
    .X(net648));
 sg13g2_buf_8 fanout649 (.A(net650),
    .X(net649));
 sg13g2_buf_8 fanout650 (.A(net651),
    .X(net650));
 sg13g2_buf_1 fanout651 (.A(_2087_),
    .X(net651));
 sg13g2_buf_8 fanout652 (.A(net653),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(net654),
    .X(net653));
 sg13g2_buf_8 fanout654 (.A(_2077_),
    .X(net654));
 sg13g2_buf_8 fanout655 (.A(net656),
    .X(net655));
 sg13g2_buf_8 fanout656 (.A(net657),
    .X(net656));
 sg13g2_buf_8 fanout657 (.A(net675),
    .X(net657));
 sg13g2_buf_8 fanout658 (.A(net675),
    .X(net658));
 sg13g2_buf_8 fanout659 (.A(net660),
    .X(net659));
 sg13g2_buf_1 fanout660 (.A(net661),
    .X(net660));
 sg13g2_buf_8 fanout661 (.A(net662),
    .X(net661));
 sg13g2_buf_8 fanout662 (.A(net675),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(net664),
    .X(net663));
 sg13g2_buf_1 fanout664 (.A(net674),
    .X(net664));
 sg13g2_buf_8 fanout665 (.A(net668),
    .X(net665));
 sg13g2_buf_1 fanout666 (.A(net667),
    .X(net666));
 sg13g2_buf_8 fanout667 (.A(net668),
    .X(net667));
 sg13g2_buf_8 fanout668 (.A(net674),
    .X(net668));
 sg13g2_buf_8 fanout669 (.A(net673),
    .X(net669));
 sg13g2_buf_8 fanout670 (.A(net673),
    .X(net670));
 sg13g2_buf_8 fanout671 (.A(net672),
    .X(net671));
 sg13g2_buf_8 fanout672 (.A(net673),
    .X(net672));
 sg13g2_buf_8 fanout673 (.A(net674),
    .X(net673));
 sg13g2_buf_8 fanout674 (.A(net675),
    .X(net674));
 sg13g2_buf_8 fanout675 (.A(_1415_),
    .X(net675));
 sg13g2_buf_8 fanout676 (.A(net677),
    .X(net676));
 sg13g2_buf_8 fanout677 (.A(net680),
    .X(net677));
 sg13g2_buf_8 fanout678 (.A(net680),
    .X(net678));
 sg13g2_buf_8 fanout679 (.A(net680),
    .X(net679));
 sg13g2_buf_8 fanout680 (.A(net693),
    .X(net680));
 sg13g2_buf_8 fanout681 (.A(net682),
    .X(net681));
 sg13g2_buf_8 fanout682 (.A(net693),
    .X(net682));
 sg13g2_buf_8 fanout683 (.A(net684),
    .X(net683));
 sg13g2_buf_8 fanout684 (.A(net693),
    .X(net684));
 sg13g2_buf_8 fanout685 (.A(net688),
    .X(net685));
 sg13g2_buf_8 fanout686 (.A(net687),
    .X(net686));
 sg13g2_buf_8 fanout687 (.A(net688),
    .X(net687));
 sg13g2_buf_8 fanout688 (.A(net693),
    .X(net688));
 sg13g2_buf_8 fanout689 (.A(net691),
    .X(net689));
 sg13g2_buf_1 fanout690 (.A(net691),
    .X(net690));
 sg13g2_buf_8 fanout691 (.A(net692),
    .X(net691));
 sg13g2_buf_8 fanout692 (.A(net693),
    .X(net692));
 sg13g2_buf_8 fanout693 (.A(_2076_),
    .X(net693));
 sg13g2_buf_8 fanout694 (.A(net697),
    .X(net694));
 sg13g2_buf_8 fanout695 (.A(net697),
    .X(net695));
 sg13g2_buf_8 fanout696 (.A(net697),
    .X(net696));
 sg13g2_buf_8 fanout697 (.A(_2075_),
    .X(net697));
 sg13g2_buf_2 fanout698 (.A(_1980_),
    .X(net698));
 sg13g2_buf_8 fanout699 (.A(_1965_),
    .X(net699));
 sg13g2_buf_8 fanout700 (.A(net701),
    .X(net700));
 sg13g2_buf_8 fanout701 (.A(_1964_),
    .X(net701));
 sg13g2_buf_8 fanout702 (.A(net703),
    .X(net702));
 sg13g2_buf_8 fanout703 (.A(_1964_),
    .X(net703));
 sg13g2_buf_8 fanout704 (.A(net705),
    .X(net704));
 sg13g2_buf_8 fanout705 (.A(net356),
    .X(net705));
 sg13g2_buf_8 fanout706 (.A(net707),
    .X(net706));
 sg13g2_buf_8 fanout707 (.A(net708),
    .X(net707));
 sg13g2_buf_8 fanout708 (.A(\mul_b_shift[30] ),
    .X(net708));
 sg13g2_buf_8 fanout709 (.A(net710),
    .X(net709));
 sg13g2_buf_8 fanout710 (.A(net711),
    .X(net710));
 sg13g2_buf_8 fanout711 (.A(\mul_b_shift[30] ),
    .X(net711));
 sg13g2_buf_8 fanout712 (.A(net714),
    .X(net712));
 sg13g2_buf_1 fanout713 (.A(net714),
    .X(net713));
 sg13g2_buf_8 fanout714 (.A(\mul_b_shift[30] ),
    .X(net714));
 sg13g2_buf_8 fanout715 (.A(net716),
    .X(net715));
 sg13g2_buf_8 fanout716 (.A(net377),
    .X(net716));
 sg13g2_buf_8 fanout717 (.A(net377),
    .X(net717));
 sg13g2_buf_1 fanout718 (.A(net377),
    .X(net718));
 sg13g2_buf_8 fanout719 (.A(net378),
    .X(net719));
 sg13g2_buf_1 fanout720 (.A(\read_counter[1] ),
    .X(net720));
 sg13g2_buf_8 fanout721 (.A(net301),
    .X(net721));
 sg13g2_buf_8 fanout722 (.A(net120),
    .X(net722));
 sg13g2_buf_8 fanout723 (.A(net369),
    .X(net723));
 sg13g2_buf_8 fanout724 (.A(net370),
    .X(net724));
 sg13g2_buf_8 fanout725 (.A(net123),
    .X(net725));
 sg13g2_buf_8 fanout726 (.A(net367),
    .X(net726));
 sg13g2_buf_8 fanout727 (.A(net376),
    .X(net727));
 sg13g2_buf_8 fanout728 (.A(net368),
    .X(net728));
 sg13g2_buf_8 fanout729 (.A(net375),
    .X(net729));
 sg13g2_buf_8 fanout730 (.A(net365),
    .X(net730));
 sg13g2_buf_8 fanout731 (.A(net373),
    .X(net731));
 sg13g2_buf_8 fanout732 (.A(\reg_a[29] ),
    .X(net732));
 sg13g2_buf_8 fanout733 (.A(\reg_a[28] ),
    .X(net733));
 sg13g2_buf_8 fanout734 (.A(net371),
    .X(net734));
 sg13g2_buf_8 fanout735 (.A(\reg_a[24] ),
    .X(net735));
 sg13g2_buf_8 fanout736 (.A(\reg_a[23] ),
    .X(net736));
 sg13g2_buf_1 fanout737 (.A(\reg_a[23] ),
    .X(net737));
 sg13g2_buf_8 fanout738 (.A(\reg_a[22] ),
    .X(net738));
 sg13g2_buf_8 fanout739 (.A(\reg_a[21] ),
    .X(net739));
 sg13g2_buf_8 fanout740 (.A(\reg_a[16] ),
    .X(net740));
 sg13g2_buf_8 fanout741 (.A(\reg_a[13] ),
    .X(net741));
 sg13g2_buf_8 fanout742 (.A(net384),
    .X(net742));
 sg13g2_buf_8 fanout743 (.A(\reg_a[10] ),
    .X(net743));
 sg13g2_buf_8 fanout744 (.A(\reg_a[8] ),
    .X(net744));
 sg13g2_buf_8 fanout745 (.A(\reg_a[7] ),
    .X(net745));
 sg13g2_buf_8 fanout746 (.A(\reg_a[2] ),
    .X(net746));
 sg13g2_buf_8 fanout747 (.A(\reg_a[1] ),
    .X(net747));
 sg13g2_buf_8 fanout748 (.A(net750),
    .X(net748));
 sg13g2_buf_1 fanout749 (.A(net750),
    .X(net749));
 sg13g2_buf_8 fanout750 (.A(net752),
    .X(net750));
 sg13g2_buf_8 fanout751 (.A(net752),
    .X(net751));
 sg13g2_buf_2 fanout752 (.A(_1967_),
    .X(net752));
 sg13g2_buf_8 fanout753 (.A(net756),
    .X(net753));
 sg13g2_buf_2 fanout754 (.A(net755),
    .X(net754));
 sg13g2_buf_1 fanout755 (.A(net756),
    .X(net755));
 sg13g2_buf_2 fanout756 (.A(_1967_),
    .X(net756));
 sg13g2_buf_8 fanout757 (.A(net758),
    .X(net757));
 sg13g2_buf_8 fanout758 (.A(net759),
    .X(net758));
 sg13g2_buf_8 fanout759 (.A(_1966_),
    .X(net759));
 sg13g2_buf_8 fanout760 (.A(net761),
    .X(net760));
 sg13g2_buf_8 fanout761 (.A(_1966_),
    .X(net761));
 sg13g2_buf_8 fanout762 (.A(net763),
    .X(net762));
 sg13g2_buf_8 fanout763 (.A(net767),
    .X(net763));
 sg13g2_buf_8 fanout764 (.A(net766),
    .X(net764));
 sg13g2_buf_1 fanout765 (.A(net766),
    .X(net765));
 sg13g2_buf_8 fanout766 (.A(net767),
    .X(net766));
 sg13g2_buf_8 fanout767 (.A(uio_in[3]),
    .X(net767));
 sg13g2_buf_8 fanout768 (.A(net776),
    .X(net768));
 sg13g2_buf_8 fanout769 (.A(net776),
    .X(net769));
 sg13g2_buf_8 fanout770 (.A(net772),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(net772),
    .X(net771));
 sg13g2_buf_8 fanout772 (.A(net776),
    .X(net772));
 sg13g2_buf_8 fanout773 (.A(net775),
    .X(net773));
 sg13g2_buf_2 fanout774 (.A(net775),
    .X(net774));
 sg13g2_buf_8 fanout775 (.A(net776),
    .X(net775));
 sg13g2_buf_8 fanout776 (.A(net808),
    .X(net776));
 sg13g2_buf_8 fanout777 (.A(net780),
    .X(net777));
 sg13g2_buf_8 fanout778 (.A(net779),
    .X(net778));
 sg13g2_buf_8 fanout779 (.A(net780),
    .X(net779));
 sg13g2_buf_8 fanout780 (.A(net808),
    .X(net780));
 sg13g2_buf_8 fanout781 (.A(net785),
    .X(net781));
 sg13g2_buf_8 fanout782 (.A(net784),
    .X(net782));
 sg13g2_buf_8 fanout783 (.A(net784),
    .X(net783));
 sg13g2_buf_8 fanout784 (.A(net785),
    .X(net784));
 sg13g2_buf_8 fanout785 (.A(net808),
    .X(net785));
 sg13g2_buf_8 fanout786 (.A(net788),
    .X(net786));
 sg13g2_buf_8 fanout787 (.A(net788),
    .X(net787));
 sg13g2_buf_8 fanout788 (.A(net807),
    .X(net788));
 sg13g2_buf_8 fanout789 (.A(net792),
    .X(net789));
 sg13g2_buf_8 fanout790 (.A(net792),
    .X(net790));
 sg13g2_buf_8 fanout791 (.A(net792),
    .X(net791));
 sg13g2_buf_8 fanout792 (.A(net807),
    .X(net792));
 sg13g2_buf_8 fanout793 (.A(net795),
    .X(net793));
 sg13g2_buf_8 fanout794 (.A(net795),
    .X(net794));
 sg13g2_buf_8 fanout795 (.A(net807),
    .X(net795));
 sg13g2_buf_8 fanout796 (.A(net797),
    .X(net796));
 sg13g2_buf_8 fanout797 (.A(net807),
    .X(net797));
 sg13g2_buf_8 fanout798 (.A(net800),
    .X(net798));
 sg13g2_buf_8 fanout799 (.A(net800),
    .X(net799));
 sg13g2_buf_8 fanout800 (.A(net806),
    .X(net800));
 sg13g2_buf_8 fanout801 (.A(net806),
    .X(net801));
 sg13g2_buf_8 fanout802 (.A(net806),
    .X(net802));
 sg13g2_buf_8 fanout803 (.A(net805),
    .X(net803));
 sg13g2_buf_8 fanout804 (.A(net805),
    .X(net804));
 sg13g2_buf_8 fanout805 (.A(net806),
    .X(net805));
 sg13g2_buf_8 fanout806 (.A(net807),
    .X(net806));
 sg13g2_buf_8 fanout807 (.A(net808),
    .X(net807));
 sg13g2_buf_8 fanout808 (.A(rst_n),
    .X(net808));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_tielo tt_um_brmurrell3_m31_accel_12 (.L_LO(net12));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_3_7__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_leaf_28_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\mul_counter[0] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold2 (.A(\mul_counter[3] ),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0102_),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold4 (.A(\mul_counter[2] ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0101_),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold6 (.A(\mul_operand_r[0] ),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0197_),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold8 (.A(\mul_accum[0] ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold9 (.A(\mul_accum[61] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0165_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold11 (.A(\reg_b[31] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold12 (.A(\mul_counter[4] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold13 (.A(\mul_operand_r[14] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0211_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold15 (.A(\mul_b_shift[8] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold16 (.A(_1763_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0174_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold18 (.A(\mul_operand_r[18] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0215_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold20 (.A(\mul_accum[59] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0163_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold22 (.A(\mul_accum[60] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0164_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold24 (.A(\mul_operand_r[13] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0210_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold26 (.A(\mul_b_shift[1] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold27 (.A(_1744_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0167_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold29 (.A(\mul_operand_r[1] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0198_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold31 (.A(\mul_b_shift[2] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0168_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold33 (.A(\mul_operand_r[16] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0213_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold35 (.A(\mul_operand_r[20] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0217_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold37 (.A(\mul_operand_r[17] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0214_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold39 (.A(\mul_b_shift[11] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold40 (.A(_1772_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0177_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold42 (.A(\mul_b_shift[23] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold43 (.A(_1808_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0189_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold45 (.A(\reg_c[1] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0077_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold47 (.A(\mul_b_shift[15] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold48 (.A(_1786_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0181_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold50 (.A(\mul_operand_r[29] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0226_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold52 (.A(\reg_c[3] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0091_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold54 (.A(\mul_operand_r[21] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0218_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold56 (.A(\mul_b_shift[4] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold57 (.A(_1751_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0170_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold59 (.A(\mul_b_shift[7] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold60 (.A(_1760_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0173_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold62 (.A(\mul_b_shift[3] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0169_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold64 (.A(\mul_b_shift[22] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold65 (.A(_1805_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0188_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold67 (.A(\mul_b_shift[28] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold68 (.A(_1825_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0194_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold70 (.A(\mul_operand_r[12] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0209_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold72 (.A(\mul_b_shift[29] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0195_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold74 (.A(\mul_b_shift[13] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold75 (.A(_1778_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0179_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold77 (.A(\mul_operand_r[6] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0203_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold79 (.A(\mul_b_shift[20] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold80 (.A(_1801_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0186_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold82 (.A(\mul_b_shift[17] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold83 (.A(_1792_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0183_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold85 (.A(\mul_b_shift[14] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0180_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold87 (.A(\reg_c[6] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0094_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold89 (.A(\reg_c[9] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0097_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold91 (.A(\mul_b_shift[27] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold92 (.A(_1820_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0193_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold94 (.A(\reg_b[29] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold95 (.A(\mul_b_shift[18] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0184_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold97 (.A(\reg_b[23] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold98 (.A(\mul_b_shift[21] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0187_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold100 (.A(\reg_c[4] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0092_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold102 (.A(\mul_b_shift[10] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold103 (.A(_1769_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0176_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold105 (.A(\mul_b_shift[9] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0175_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold107 (.A(\mul_accum[15] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0119_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold109 (.A(\mul_operand_r[19] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0216_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold111 (.A(\mul_operand_r[2] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0199_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold113 (.A(\reg_c[30] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold114 (.A(\mul_b_shift[0] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold115 (.A(_1741_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold116 (.A(\reg_c[7] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0095_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold118 (.A(\mul_b_shift[24] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0190_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold120 (.A(\reg_c[23] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0081_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold122 (.A(\mul_operand_r[15] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0212_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold124 (.A(\reg_c[28] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold125 (.A(\mul_accum[34] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0138_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold127 (.A(\mul_accum[52] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0156_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold129 (.A(\reg_c[31] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold130 (.A(\reg_c[29] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold131 (.A(\mul_accum[22] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0126_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold133 (.A(\reg_c[0] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0066_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold135 (.A(\mul_operand_r[4] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0201_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold137 (.A(\mul_b_shift[6] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold138 (.A(_1759_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0172_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold140 (.A(\mul_operand_r[26] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0223_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold142 (.A(\mul_operand_r[5] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0202_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold144 (.A(\mul_b_shift[5] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0171_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold146 (.A(\reg_c[2] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0088_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold148 (.A(\mul_b_shift[26] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold149 (.A(_1819_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0192_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold151 (.A(\reg_c[25] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold152 (.A(\mul_b_shift[19] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0185_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold154 (.A(\mul_operand_r[30] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0227_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold156 (.A(\reg_c[13] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0070_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold158 (.A(\reg_c[22] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold159 (.A(\mul_operand_r[3] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0200_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold161 (.A(\reg_c[15] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold162 (.A(\mul_accum[46] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0150_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold164 (.A(\mul_accum[11] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0115_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold166 (.A(\mul_operand_r[9] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0206_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold168 (.A(\mul_b_shift[12] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0178_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold170 (.A(\reg_c[5] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold171 (.A(\mul_accum[57] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0161_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold173 (.A(\mul_b_shift[25] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0191_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold175 (.A(\reg_c[20] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold176 (.A(\reg_c[21] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold177 (.A(\mul_accum[54] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0158_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold179 (.A(\mul_accum[32] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0136_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold181 (.A(\mul_accum[7] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0111_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold183 (.A(\mul_counter[1] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold184 (.A(\mul_operand_r[27] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0224_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold186 (.A(\reg_c[19] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0076_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold188 (.A(\mul_operand_r[25] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0222_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold190 (.A(\reg_c[12] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold191 (.A(\mul_operand_r[28] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0225_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold193 (.A(\reg_c[14] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold194 (.A(\reg_c[26] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold195 (.A(\mul_operand_r[24] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0221_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold197 (.A(\mul_accum[40] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0144_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold199 (.A(\reg_c[16] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0073_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold201 (.A(\mul_operand_r[8] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0205_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold203 (.A(\mul_operand_r[23] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0220_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold205 (.A(\reg_c[24] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold206 (.A(\reg_c[18] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold207 (.A(\reg_c[11] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold208 (.A(\mul_operand_r[22] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0219_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold210 (.A(\reg_c[27] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold211 (.A(\reg_a[31] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold212 (.A(\mul_b_shift[16] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0182_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold214 (.A(\mul_operand_r[7] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0204_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold216 (.A(\mul_operand_r[11] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0208_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold218 (.A(\mul_operand_r[10] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0207_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold220 (.A(\mul_accum[55] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold221 (.A(_1721_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold222 (.A(\reg_c[10] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold223 (.A(\reg_b[0] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0034_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold225 (.A(\mul_accum[38] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold226 (.A(_1670_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold227 (.A(\mul_accum[35] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold228 (.A(_1661_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold229 (.A(\mul_accum[23] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold230 (.A(\reg_b[1] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0045_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold232 (.A(\mul_accum[29] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0133_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold234 (.A(\reg_b[2] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0056_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold236 (.A(\reg_b[15] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold237 (.A(\mul_accum[50] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold238 (.A(_1706_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold239 (.A(\mul_accum[28] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0132_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold241 (.A(\mul_accum[31] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold242 (.A(_1648_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold243 (.A(\reg_c[17] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold244 (.A(\mul_accum[44] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold245 (.A(_1687_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold246 (.A(\mul_accum[19] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0123_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold248 (.A(\mul_accum[56] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold249 (.A(_1725_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold250 (.A(\mul_accum[49] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold251 (.A(_1702_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold252 (.A(\reg_c[8] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold253 (.A(\mul_accum[14] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0118_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold255 (.A(\mul_accum[25] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0129_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold257 (.A(\reg_b[30] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0196_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold259 (.A(\mul_accum[26] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold260 (.A(\mul_accum[16] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold261 (.A(\mul_accum[18] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0122_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold263 (.A(\mul_accum[37] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold264 (.A(_1667_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold265 (.A(\mul_accum[53] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold266 (.A(_1716_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold267 (.A(\mul_accum[36] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold268 (.A(_1664_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold269 (.A(\mul_accum[42] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold270 (.A(_1682_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold271 (.A(\mul_accum[48] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold272 (.A(_1700_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold273 (.A(\mul_accum[21] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold274 (.A(_0125_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold275 (.A(\read_counter[0] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold276 (.A(\mul_accum[12] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold277 (.A(\mul_accum[20] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold278 (.A(\mul_accum[43] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold279 (.A(\mul_accum[24] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0128_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold281 (.A(\mul_accum[45] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold282 (.A(_1691_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold283 (.A(\mul_accum[41] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold284 (.A(_1679_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold285 (.A(\reg_b[8] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0064_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold287 (.A(\mul_accum[27] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0131_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold289 (.A(\mul_accum[8] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0112_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold291 (.A(\mul_accum[58] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold292 (.A(\reg_b[4] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0060_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold294 (.A(\mul_accum[51] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold295 (.A(_1710_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold296 (.A(\reg_b[3] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold297 (.A(_0059_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold298 (.A(\mul_accum[10] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold299 (.A(_0114_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold300 (.A(\mul_accum[47] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold301 (.A(\reg_b[10] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0035_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold303 (.A(\mul_accum[4] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0108_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold305 (.A(\mul_accum[3] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold306 (.A(_0107_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold307 (.A(\reg_b[26] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold308 (.A(\mul_accum[2] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0106_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold310 (.A(\mul_accum[6] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0110_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold312 (.A(\reg_b[12] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold313 (.A(_0037_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold314 (.A(\reg_b[16] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold315 (.A(_0041_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold316 (.A(\mul_accum[5] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold317 (.A(\reg_b[11] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold318 (.A(_0036_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold319 (.A(\reg_b[6] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0062_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold321 (.A(\reg_b[7] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold322 (.A(\reg_b[24] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold323 (.A(\reg_b[28] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold324 (.A(\mul_accum[39] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold325 (.A(\reg_b[20] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold326 (.A(\mul_accum[33] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold327 (.A(\reg_b[14] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold328 (.A(_0039_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold329 (.A(\reg_b[22] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold330 (.A(reducing),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold331 (.A(\mul_accum[1] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold332 (.A(\reg_b[5] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold333 (.A(_0061_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold334 (.A(\mul_accum[17] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold335 (.A(\mul_accum[30] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold336 (.A(_0134_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold337 (.A(\mul_accum[13] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold338 (.A(\mul_accum[9] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold339 (.A(\reg_b[13] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0038_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold341 (.A(\reg_b[21] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold342 (.A(\reg_b[18] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold343 (.A(\reg_b[27] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold344 (.A(\reg_b[25] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold345 (.A(\reg_a[26] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold346 (.A(_1293_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold347 (.A(\reg_b[9] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0065_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold349 (.A(\reg_b[17] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold350 (.A(\reg_b[19] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold351 (.A(mac_mode),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold352 (.A(\read_counter[1] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold353 (.A(\reg_a[25] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold354 (.A(_1290_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold355 (.A(\reg_a[20] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold356 (.A(\reg_a[27] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold357 (.A(_1303_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold358 (.A(\reg_a[12] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold359 (.A(\reg_a[3] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold360 (.A(_1154_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold361 (.A(\reg_a[28] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold362 (.A(\reg_a[14] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold363 (.A(\reg_a[29] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold364 (.A(\reg_a[30] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold365 (.A(\mul_accum[41] ),
    .X(net391));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_79 ();
 sg13g2_fill_1 FILLER_0_86 ();
 sg13g2_decap_8 FILLER_0_113 ();
 sg13g2_decap_4 FILLER_0_120 ();
 sg13g2_decap_8 FILLER_0_127 ();
 sg13g2_decap_8 FILLER_0_134 ();
 sg13g2_fill_1 FILLER_0_141 ();
 sg13g2_decap_8 FILLER_0_145 ();
 sg13g2_decap_8 FILLER_0_152 ();
 sg13g2_decap_8 FILLER_0_159 ();
 sg13g2_decap_8 FILLER_0_166 ();
 sg13g2_decap_8 FILLER_0_173 ();
 sg13g2_decap_4 FILLER_0_180 ();
 sg13g2_decap_8 FILLER_0_194 ();
 sg13g2_decap_8 FILLER_0_201 ();
 sg13g2_decap_8 FILLER_0_208 ();
 sg13g2_decap_8 FILLER_0_215 ();
 sg13g2_decap_8 FILLER_0_222 ();
 sg13g2_decap_8 FILLER_0_229 ();
 sg13g2_decap_4 FILLER_0_236 ();
 sg13g2_fill_1 FILLER_0_246 ();
 sg13g2_fill_1 FILLER_0_258 ();
 sg13g2_decap_8 FILLER_0_264 ();
 sg13g2_decap_4 FILLER_0_271 ();
 sg13g2_fill_1 FILLER_0_275 ();
 sg13g2_fill_2 FILLER_0_300 ();
 sg13g2_fill_1 FILLER_0_302 ();
 sg13g2_fill_2 FILLER_0_307 ();
 sg13g2_fill_1 FILLER_0_309 ();
 sg13g2_decap_4 FILLER_0_314 ();
 sg13g2_fill_1 FILLER_0_318 ();
 sg13g2_fill_1 FILLER_0_325 ();
 sg13g2_decap_8 FILLER_0_354 ();
 sg13g2_decap_8 FILLER_0_361 ();
 sg13g2_decap_8 FILLER_0_368 ();
 sg13g2_decap_8 FILLER_0_375 ();
 sg13g2_decap_8 FILLER_0_382 ();
 sg13g2_decap_8 FILLER_0_389 ();
 sg13g2_decap_8 FILLER_0_396 ();
 sg13g2_decap_4 FILLER_0_403 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_fill_1 FILLER_1_95 ();
 sg13g2_fill_2 FILLER_1_111 ();
 sg13g2_fill_1 FILLER_1_149 ();
 sg13g2_decap_4 FILLER_1_184 ();
 sg13g2_fill_2 FILLER_1_193 ();
 sg13g2_fill_2 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_362 ();
 sg13g2_decap_8 FILLER_1_369 ();
 sg13g2_decap_8 FILLER_1_376 ();
 sg13g2_decap_8 FILLER_1_383 ();
 sg13g2_decap_8 FILLER_1_390 ();
 sg13g2_decap_8 FILLER_1_397 ();
 sg13g2_decap_4 FILLER_1_404 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_4 FILLER_2_49 ();
 sg13g2_fill_1 FILLER_2_89 ();
 sg13g2_fill_1 FILLER_2_211 ();
 sg13g2_fill_2 FILLER_2_292 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_4 FILLER_3_49 ();
 sg13g2_fill_1 FILLER_3_53 ();
 sg13g2_fill_2 FILLER_3_57 ();
 sg13g2_fill_2 FILLER_3_128 ();
 sg13g2_fill_2 FILLER_3_155 ();
 sg13g2_fill_2 FILLER_3_197 ();
 sg13g2_fill_1 FILLER_3_199 ();
 sg13g2_fill_2 FILLER_3_214 ();
 sg13g2_fill_1 FILLER_3_231 ();
 sg13g2_fill_2 FILLER_3_250 ();
 sg13g2_fill_2 FILLER_3_264 ();
 sg13g2_fill_1 FILLER_3_300 ();
 sg13g2_fill_2 FILLER_3_314 ();
 sg13g2_decap_8 FILLER_3_387 ();
 sg13g2_decap_8 FILLER_3_394 ();
 sg13g2_decap_8 FILLER_3_401 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_4 FILLER_4_56 ();
 sg13g2_fill_2 FILLER_4_77 ();
 sg13g2_fill_1 FILLER_4_79 ();
 sg13g2_fill_2 FILLER_4_104 ();
 sg13g2_fill_1 FILLER_4_106 ();
 sg13g2_fill_2 FILLER_4_127 ();
 sg13g2_fill_1 FILLER_4_144 ();
 sg13g2_fill_2 FILLER_4_154 ();
 sg13g2_fill_1 FILLER_4_181 ();
 sg13g2_fill_2 FILLER_4_255 ();
 sg13g2_fill_2 FILLER_4_270 ();
 sg13g2_fill_1 FILLER_4_272 ();
 sg13g2_fill_2 FILLER_4_363 ();
 sg13g2_decap_8 FILLER_4_398 ();
 sg13g2_decap_4 FILLER_4_405 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_4 FILLER_5_63 ();
 sg13g2_fill_1 FILLER_5_81 ();
 sg13g2_fill_2 FILLER_5_98 ();
 sg13g2_fill_1 FILLER_5_100 ();
 sg13g2_fill_2 FILLER_5_115 ();
 sg13g2_fill_1 FILLER_5_117 ();
 sg13g2_fill_2 FILLER_5_133 ();
 sg13g2_fill_2 FILLER_5_153 ();
 sg13g2_decap_8 FILLER_5_195 ();
 sg13g2_fill_1 FILLER_5_202 ();
 sg13g2_decap_4 FILLER_5_208 ();
 sg13g2_fill_2 FILLER_5_212 ();
 sg13g2_decap_4 FILLER_5_226 ();
 sg13g2_fill_2 FILLER_5_230 ();
 sg13g2_decap_4 FILLER_5_285 ();
 sg13g2_fill_1 FILLER_5_289 ();
 sg13g2_decap_4 FILLER_5_318 ();
 sg13g2_fill_1 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_395 ();
 sg13g2_decap_8 FILLER_5_402 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_4 FILLER_6_42 ();
 sg13g2_fill_2 FILLER_6_107 ();
 sg13g2_fill_1 FILLER_6_109 ();
 sg13g2_fill_2 FILLER_6_138 ();
 sg13g2_fill_1 FILLER_6_158 ();
 sg13g2_fill_2 FILLER_6_240 ();
 sg13g2_fill_1 FILLER_6_279 ();
 sg13g2_fill_2 FILLER_6_302 ();
 sg13g2_decap_4 FILLER_6_339 ();
 sg13g2_decap_4 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_391 ();
 sg13g2_decap_8 FILLER_6_398 ();
 sg13g2_decap_4 FILLER_6_405 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_fill_1 FILLER_7_42 ();
 sg13g2_fill_1 FILLER_7_89 ();
 sg13g2_fill_1 FILLER_7_156 ();
 sg13g2_fill_2 FILLER_7_199 ();
 sg13g2_fill_1 FILLER_7_201 ();
 sg13g2_fill_2 FILLER_7_230 ();
 sg13g2_fill_1 FILLER_7_232 ();
 sg13g2_fill_2 FILLER_7_320 ();
 sg13g2_fill_1 FILLER_7_322 ();
 sg13g2_fill_2 FILLER_7_337 ();
 sg13g2_decap_4 FILLER_7_344 ();
 sg13g2_fill_2 FILLER_7_348 ();
 sg13g2_decap_4 FILLER_7_355 ();
 sg13g2_fill_1 FILLER_7_359 ();
 sg13g2_fill_2 FILLER_7_373 ();
 sg13g2_fill_1 FILLER_7_375 ();
 sg13g2_decap_8 FILLER_7_395 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_fill_2 FILLER_8_42 ();
 sg13g2_fill_1 FILLER_8_44 ();
 sg13g2_decap_4 FILLER_8_52 ();
 sg13g2_decap_4 FILLER_8_123 ();
 sg13g2_fill_1 FILLER_8_151 ();
 sg13g2_fill_1 FILLER_8_162 ();
 sg13g2_fill_2 FILLER_8_168 ();
 sg13g2_fill_1 FILLER_8_170 ();
 sg13g2_fill_1 FILLER_8_184 ();
 sg13g2_decap_4 FILLER_8_229 ();
 sg13g2_fill_2 FILLER_8_233 ();
 sg13g2_fill_1 FILLER_8_239 ();
 sg13g2_fill_2 FILLER_8_244 ();
 sg13g2_fill_1 FILLER_8_270 ();
 sg13g2_fill_1 FILLER_8_280 ();
 sg13g2_fill_1 FILLER_8_290 ();
 sg13g2_decap_8 FILLER_8_303 ();
 sg13g2_decap_8 FILLER_8_316 ();
 sg13g2_decap_8 FILLER_8_323 ();
 sg13g2_decap_8 FILLER_8_349 ();
 sg13g2_decap_8 FILLER_8_356 ();
 sg13g2_fill_2 FILLER_8_381 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_fill_1 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_51 ();
 sg13g2_decap_8 FILLER_9_65 ();
 sg13g2_fill_1 FILLER_9_72 ();
 sg13g2_fill_1 FILLER_9_109 ();
 sg13g2_fill_2 FILLER_9_119 ();
 sg13g2_fill_1 FILLER_9_121 ();
 sg13g2_fill_2 FILLER_9_132 ();
 sg13g2_fill_1 FILLER_9_134 ();
 sg13g2_fill_1 FILLER_9_154 ();
 sg13g2_fill_2 FILLER_9_167 ();
 sg13g2_fill_1 FILLER_9_169 ();
 sg13g2_decap_8 FILLER_9_181 ();
 sg13g2_fill_2 FILLER_9_188 ();
 sg13g2_decap_8 FILLER_9_213 ();
 sg13g2_decap_4 FILLER_9_220 ();
 sg13g2_fill_2 FILLER_9_224 ();
 sg13g2_fill_1 FILLER_9_230 ();
 sg13g2_fill_2 FILLER_9_248 ();
 sg13g2_fill_1 FILLER_9_260 ();
 sg13g2_fill_2 FILLER_9_266 ();
 sg13g2_decap_4 FILLER_9_272 ();
 sg13g2_fill_1 FILLER_9_276 ();
 sg13g2_decap_8 FILLER_9_281 ();
 sg13g2_fill_2 FILLER_9_288 ();
 sg13g2_fill_2 FILLER_9_361 ();
 sg13g2_fill_2 FILLER_9_371 ();
 sg13g2_fill_1 FILLER_9_373 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_7 ();
 sg13g2_fill_2 FILLER_10_11 ();
 sg13g2_decap_8 FILLER_10_72 ();
 sg13g2_decap_4 FILLER_10_79 ();
 sg13g2_fill_2 FILLER_10_83 ();
 sg13g2_decap_4 FILLER_10_89 ();
 sg13g2_fill_1 FILLER_10_102 ();
 sg13g2_fill_1 FILLER_10_108 ();
 sg13g2_fill_2 FILLER_10_114 ();
 sg13g2_decap_8 FILLER_10_121 ();
 sg13g2_decap_8 FILLER_10_128 ();
 sg13g2_fill_2 FILLER_10_135 ();
 sg13g2_fill_1 FILLER_10_137 ();
 sg13g2_fill_1 FILLER_10_148 ();
 sg13g2_decap_4 FILLER_10_163 ();
 sg13g2_decap_4 FILLER_10_180 ();
 sg13g2_fill_1 FILLER_10_184 ();
 sg13g2_decap_8 FILLER_10_198 ();
 sg13g2_decap_8 FILLER_10_205 ();
 sg13g2_decap_8 FILLER_10_212 ();
 sg13g2_fill_1 FILLER_10_219 ();
 sg13g2_fill_2 FILLER_10_253 ();
 sg13g2_fill_1 FILLER_10_255 ();
 sg13g2_fill_1 FILLER_10_264 ();
 sg13g2_fill_2 FILLER_10_270 ();
 sg13g2_fill_2 FILLER_10_276 ();
 sg13g2_fill_1 FILLER_10_278 ();
 sg13g2_fill_2 FILLER_10_309 ();
 sg13g2_fill_1 FILLER_10_352 ();
 sg13g2_fill_1 FILLER_10_379 ();
 sg13g2_fill_2 FILLER_10_390 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_4 FILLER_11_14 ();
 sg13g2_fill_1 FILLER_11_18 ();
 sg13g2_decap_4 FILLER_11_68 ();
 sg13g2_fill_1 FILLER_11_72 ();
 sg13g2_fill_2 FILLER_11_90 ();
 sg13g2_fill_1 FILLER_11_99 ();
 sg13g2_fill_2 FILLER_11_117 ();
 sg13g2_fill_2 FILLER_11_139 ();
 sg13g2_decap_4 FILLER_11_217 ();
 sg13g2_fill_1 FILLER_11_231 ();
 sg13g2_fill_2 FILLER_11_243 ();
 sg13g2_decap_4 FILLER_11_258 ();
 sg13g2_decap_4 FILLER_11_298 ();
 sg13g2_fill_1 FILLER_11_302 ();
 sg13g2_fill_1 FILLER_11_323 ();
 sg13g2_fill_2 FILLER_11_334 ();
 sg13g2_fill_2 FILLER_11_346 ();
 sg13g2_fill_1 FILLER_11_348 ();
 sg13g2_fill_2 FILLER_11_375 ();
 sg13g2_fill_2 FILLER_11_390 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_55 ();
 sg13g2_fill_1 FILLER_12_62 ();
 sg13g2_fill_1 FILLER_12_89 ();
 sg13g2_fill_2 FILLER_12_104 ();
 sg13g2_fill_1 FILLER_12_144 ();
 sg13g2_fill_2 FILLER_12_165 ();
 sg13g2_fill_1 FILLER_12_167 ();
 sg13g2_decap_8 FILLER_12_239 ();
 sg13g2_decap_8 FILLER_12_250 ();
 sg13g2_decap_4 FILLER_12_257 ();
 sg13g2_decap_8 FILLER_12_275 ();
 sg13g2_fill_2 FILLER_12_287 ();
 sg13g2_decap_4 FILLER_12_302 ();
 sg13g2_fill_1 FILLER_12_306 ();
 sg13g2_decap_8 FILLER_12_318 ();
 sg13g2_decap_8 FILLER_12_325 ();
 sg13g2_fill_2 FILLER_12_332 ();
 sg13g2_decap_4 FILLER_12_337 ();
 sg13g2_fill_1 FILLER_12_394 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_fill_2 FILLER_13_21 ();
 sg13g2_fill_1 FILLER_13_23 ();
 sg13g2_fill_1 FILLER_13_32 ();
 sg13g2_fill_1 FILLER_13_56 ();
 sg13g2_fill_1 FILLER_13_62 ();
 sg13g2_fill_2 FILLER_13_78 ();
 sg13g2_fill_1 FILLER_13_89 ();
 sg13g2_fill_1 FILLER_13_123 ();
 sg13g2_decap_4 FILLER_13_156 ();
 sg13g2_decap_4 FILLER_13_227 ();
 sg13g2_fill_1 FILLER_13_231 ();
 sg13g2_fill_1 FILLER_13_263 ();
 sg13g2_fill_1 FILLER_13_268 ();
 sg13g2_decap_8 FILLER_13_278 ();
 sg13g2_decap_8 FILLER_13_285 ();
 sg13g2_decap_8 FILLER_13_292 ();
 sg13g2_decap_8 FILLER_13_299 ();
 sg13g2_decap_8 FILLER_13_306 ();
 sg13g2_decap_8 FILLER_13_313 ();
 sg13g2_fill_2 FILLER_13_320 ();
 sg13g2_fill_1 FILLER_13_322 ();
 sg13g2_fill_1 FILLER_13_333 ();
 sg13g2_decap_4 FILLER_13_342 ();
 sg13g2_fill_1 FILLER_13_346 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_fill_2 FILLER_14_14 ();
 sg13g2_fill_1 FILLER_14_16 ();
 sg13g2_decap_4 FILLER_14_20 ();
 sg13g2_fill_1 FILLER_14_63 ();
 sg13g2_decap_4 FILLER_14_80 ();
 sg13g2_fill_2 FILLER_14_84 ();
 sg13g2_decap_4 FILLER_14_98 ();
 sg13g2_fill_2 FILLER_14_147 ();
 sg13g2_fill_1 FILLER_14_171 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_fill_1 FILLER_14_249 ();
 sg13g2_decap_4 FILLER_14_278 ();
 sg13g2_fill_2 FILLER_14_282 ();
 sg13g2_fill_2 FILLER_14_301 ();
 sg13g2_decap_4 FILLER_14_311 ();
 sg13g2_decap_4 FILLER_14_357 ();
 sg13g2_fill_2 FILLER_14_361 ();
 sg13g2_fill_1 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_7 ();
 sg13g2_fill_1 FILLER_15_9 ();
 sg13g2_decap_4 FILLER_15_38 ();
 sg13g2_decap_4 FILLER_15_49 ();
 sg13g2_fill_2 FILLER_15_66 ();
 sg13g2_decap_8 FILLER_15_81 ();
 sg13g2_fill_1 FILLER_15_88 ();
 sg13g2_fill_1 FILLER_15_110 ();
 sg13g2_decap_8 FILLER_15_120 ();
 sg13g2_decap_8 FILLER_15_127 ();
 sg13g2_decap_8 FILLER_15_134 ();
 sg13g2_decap_4 FILLER_15_141 ();
 sg13g2_fill_2 FILLER_15_154 ();
 sg13g2_fill_2 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_201 ();
 sg13g2_decap_4 FILLER_15_208 ();
 sg13g2_fill_1 FILLER_15_212 ();
 sg13g2_fill_2 FILLER_15_225 ();
 sg13g2_decap_4 FILLER_15_239 ();
 sg13g2_fill_1 FILLER_15_243 ();
 sg13g2_fill_1 FILLER_15_267 ();
 sg13g2_fill_1 FILLER_15_309 ();
 sg13g2_fill_2 FILLER_15_323 ();
 sg13g2_fill_1 FILLER_15_325 ();
 sg13g2_decap_4 FILLER_15_343 ();
 sg13g2_decap_4 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_fill_2 FILLER_15_373 ();
 sg13g2_fill_1 FILLER_15_375 ();
 sg13g2_fill_2 FILLER_15_395 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_7 ();
 sg13g2_fill_2 FILLER_16_47 ();
 sg13g2_decap_8 FILLER_16_57 ();
 sg13g2_decap_8 FILLER_16_64 ();
 sg13g2_fill_2 FILLER_16_71 ();
 sg13g2_fill_1 FILLER_16_100 ();
 sg13g2_fill_2 FILLER_16_132 ();
 sg13g2_fill_2 FILLER_16_139 ();
 sg13g2_fill_1 FILLER_16_150 ();
 sg13g2_fill_2 FILLER_16_163 ();
 sg13g2_fill_1 FILLER_16_165 ();
 sg13g2_fill_1 FILLER_16_188 ();
 sg13g2_fill_1 FILLER_16_201 ();
 sg13g2_fill_2 FILLER_16_222 ();
 sg13g2_fill_1 FILLER_16_231 ();
 sg13g2_fill_2 FILLER_16_247 ();
 sg13g2_fill_1 FILLER_16_249 ();
 sg13g2_fill_1 FILLER_16_268 ();
 sg13g2_fill_2 FILLER_16_277 ();
 sg13g2_fill_1 FILLER_16_279 ();
 sg13g2_fill_2 FILLER_16_289 ();
 sg13g2_decap_8 FILLER_16_321 ();
 sg13g2_fill_2 FILLER_16_328 ();
 sg13g2_fill_1 FILLER_16_330 ();
 sg13g2_fill_2 FILLER_16_339 ();
 sg13g2_fill_1 FILLER_16_341 ();
 sg13g2_decap_4 FILLER_16_369 ();
 sg13g2_fill_1 FILLER_16_382 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_4 ();
 sg13g2_fill_2 FILLER_17_33 ();
 sg13g2_fill_1 FILLER_17_35 ();
 sg13g2_decap_4 FILLER_17_74 ();
 sg13g2_fill_2 FILLER_17_87 ();
 sg13g2_decap_4 FILLER_17_107 ();
 sg13g2_fill_1 FILLER_17_123 ();
 sg13g2_fill_2 FILLER_17_132 ();
 sg13g2_decap_8 FILLER_17_155 ();
 sg13g2_decap_4 FILLER_17_162 ();
 sg13g2_fill_1 FILLER_17_166 ();
 sg13g2_decap_4 FILLER_17_219 ();
 sg13g2_fill_1 FILLER_17_233 ();
 sg13g2_decap_8 FILLER_17_241 ();
 sg13g2_decap_8 FILLER_17_248 ();
 sg13g2_fill_1 FILLER_17_268 ();
 sg13g2_fill_2 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_fill_1 FILLER_17_379 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_fill_2 FILLER_18_14 ();
 sg13g2_fill_1 FILLER_18_16 ();
 sg13g2_fill_2 FILLER_18_38 ();
 sg13g2_fill_1 FILLER_18_40 ();
 sg13g2_decap_8 FILLER_18_96 ();
 sg13g2_decap_8 FILLER_18_103 ();
 sg13g2_decap_8 FILLER_18_110 ();
 sg13g2_fill_2 FILLER_18_117 ();
 sg13g2_fill_1 FILLER_18_119 ();
 sg13g2_fill_2 FILLER_18_134 ();
 sg13g2_fill_2 FILLER_18_144 ();
 sg13g2_fill_1 FILLER_18_146 ();
 sg13g2_fill_2 FILLER_18_175 ();
 sg13g2_fill_1 FILLER_18_177 ();
 sg13g2_fill_2 FILLER_18_191 ();
 sg13g2_decap_8 FILLER_18_216 ();
 sg13g2_decap_4 FILLER_18_223 ();
 sg13g2_fill_2 FILLER_18_227 ();
 sg13g2_decap_8 FILLER_18_234 ();
 sg13g2_decap_8 FILLER_18_241 ();
 sg13g2_fill_2 FILLER_18_248 ();
 sg13g2_decap_8 FILLER_18_255 ();
 sg13g2_decap_4 FILLER_18_262 ();
 sg13g2_fill_1 FILLER_18_266 ();
 sg13g2_decap_4 FILLER_18_273 ();
 sg13g2_fill_1 FILLER_18_277 ();
 sg13g2_fill_2 FILLER_18_282 ();
 sg13g2_decap_4 FILLER_18_297 ();
 sg13g2_fill_1 FILLER_18_301 ();
 sg13g2_fill_2 FILLER_18_322 ();
 sg13g2_fill_2 FILLER_18_353 ();
 sg13g2_fill_1 FILLER_18_355 ();
 sg13g2_fill_1 FILLER_18_371 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_4 ();
 sg13g2_fill_2 FILLER_19_27 ();
 sg13g2_fill_1 FILLER_19_35 ();
 sg13g2_fill_2 FILLER_19_70 ();
 sg13g2_fill_1 FILLER_19_72 ();
 sg13g2_decap_8 FILLER_19_90 ();
 sg13g2_decap_8 FILLER_19_97 ();
 sg13g2_decap_8 FILLER_19_104 ();
 sg13g2_decap_8 FILLER_19_111 ();
 sg13g2_decap_8 FILLER_19_118 ();
 sg13g2_decap_8 FILLER_19_125 ();
 sg13g2_decap_8 FILLER_19_132 ();
 sg13g2_decap_8 FILLER_19_139 ();
 sg13g2_decap_8 FILLER_19_146 ();
 sg13g2_fill_2 FILLER_19_153 ();
 sg13g2_fill_1 FILLER_19_196 ();
 sg13g2_fill_2 FILLER_19_205 ();
 sg13g2_fill_2 FILLER_19_217 ();
 sg13g2_fill_1 FILLER_19_224 ();
 sg13g2_fill_1 FILLER_19_230 ();
 sg13g2_decap_8 FILLER_19_240 ();
 sg13g2_decap_4 FILLER_19_247 ();
 sg13g2_fill_1 FILLER_19_251 ();
 sg13g2_decap_8 FILLER_19_265 ();
 sg13g2_decap_8 FILLER_19_272 ();
 sg13g2_decap_4 FILLER_19_279 ();
 sg13g2_fill_2 FILLER_19_283 ();
 sg13g2_fill_1 FILLER_19_301 ();
 sg13g2_fill_1 FILLER_19_333 ();
 sg13g2_fill_1 FILLER_19_383 ();
 sg13g2_fill_2 FILLER_19_393 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_57 ();
 sg13g2_decap_8 FILLER_20_64 ();
 sg13g2_decap_8 FILLER_20_94 ();
 sg13g2_decap_8 FILLER_20_101 ();
 sg13g2_fill_1 FILLER_20_108 ();
 sg13g2_fill_2 FILLER_20_118 ();
 sg13g2_decap_4 FILLER_20_128 ();
 sg13g2_fill_1 FILLER_20_137 ();
 sg13g2_decap_8 FILLER_20_155 ();
 sg13g2_decap_8 FILLER_20_162 ();
 sg13g2_decap_8 FILLER_20_169 ();
 sg13g2_decap_8 FILLER_20_176 ();
 sg13g2_decap_8 FILLER_20_183 ();
 sg13g2_decap_8 FILLER_20_190 ();
 sg13g2_fill_2 FILLER_20_197 ();
 sg13g2_fill_1 FILLER_20_199 ();
 sg13g2_decap_4 FILLER_20_203 ();
 sg13g2_fill_2 FILLER_20_207 ();
 sg13g2_fill_2 FILLER_20_222 ();
 sg13g2_decap_4 FILLER_20_252 ();
 sg13g2_fill_2 FILLER_20_256 ();
 sg13g2_decap_8 FILLER_20_268 ();
 sg13g2_decap_4 FILLER_20_279 ();
 sg13g2_fill_1 FILLER_20_291 ();
 sg13g2_fill_1 FILLER_20_312 ();
 sg13g2_decap_8 FILLER_20_318 ();
 sg13g2_decap_8 FILLER_20_325 ();
 sg13g2_fill_2 FILLER_20_332 ();
 sg13g2_decap_4 FILLER_20_338 ();
 sg13g2_decap_4 FILLER_20_347 ();
 sg13g2_fill_2 FILLER_20_370 ();
 sg13g2_fill_1 FILLER_20_372 ();
 sg13g2_fill_1 FILLER_20_382 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_39 ();
 sg13g2_decap_8 FILLER_21_47 ();
 sg13g2_decap_4 FILLER_21_54 ();
 sg13g2_fill_1 FILLER_21_58 ();
 sg13g2_decap_4 FILLER_21_72 ();
 sg13g2_fill_2 FILLER_21_76 ();
 sg13g2_fill_1 FILLER_21_138 ();
 sg13g2_fill_2 FILLER_21_158 ();
 sg13g2_fill_1 FILLER_21_160 ();
 sg13g2_decap_8 FILLER_21_165 ();
 sg13g2_decap_8 FILLER_21_172 ();
 sg13g2_decap_8 FILLER_21_179 ();
 sg13g2_decap_8 FILLER_21_186 ();
 sg13g2_fill_2 FILLER_21_193 ();
 sg13g2_decap_8 FILLER_21_199 ();
 sg13g2_fill_2 FILLER_21_206 ();
 sg13g2_fill_1 FILLER_21_232 ();
 sg13g2_fill_2 FILLER_21_253 ();
 sg13g2_fill_2 FILLER_21_290 ();
 sg13g2_decap_8 FILLER_21_305 ();
 sg13g2_decap_8 FILLER_21_312 ();
 sg13g2_decap_8 FILLER_21_319 ();
 sg13g2_decap_8 FILLER_21_326 ();
 sg13g2_decap_8 FILLER_21_333 ();
 sg13g2_decap_8 FILLER_21_340 ();
 sg13g2_fill_2 FILLER_21_347 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_4 FILLER_21_368 ();
 sg13g2_fill_2 FILLER_21_372 ();
 sg13g2_fill_1 FILLER_21_379 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_14 ();
 sg13g2_fill_1 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_50 ();
 sg13g2_decap_4 FILLER_22_57 ();
 sg13g2_fill_1 FILLER_22_61 ();
 sg13g2_decap_8 FILLER_22_75 ();
 sg13g2_fill_1 FILLER_22_82 ();
 sg13g2_fill_2 FILLER_22_125 ();
 sg13g2_fill_1 FILLER_22_127 ();
 sg13g2_fill_2 FILLER_22_151 ();
 sg13g2_fill_1 FILLER_22_153 ();
 sg13g2_fill_2 FILLER_22_170 ();
 sg13g2_fill_2 FILLER_22_191 ();
 sg13g2_fill_1 FILLER_22_193 ();
 sg13g2_fill_1 FILLER_22_202 ();
 sg13g2_fill_2 FILLER_22_216 ();
 sg13g2_fill_1 FILLER_22_218 ();
 sg13g2_fill_2 FILLER_22_224 ();
 sg13g2_fill_1 FILLER_22_226 ();
 sg13g2_fill_2 FILLER_22_246 ();
 sg13g2_fill_2 FILLER_22_269 ();
 sg13g2_decap_8 FILLER_22_296 ();
 sg13g2_decap_8 FILLER_22_303 ();
 sg13g2_decap_4 FILLER_22_310 ();
 sg13g2_decap_8 FILLER_22_335 ();
 sg13g2_fill_2 FILLER_22_342 ();
 sg13g2_fill_1 FILLER_22_344 ();
 sg13g2_fill_1 FILLER_22_376 ();
 sg13g2_fill_2 FILLER_22_402 ();
 sg13g2_fill_1 FILLER_22_404 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_7 ();
 sg13g2_decap_4 FILLER_23_11 ();
 sg13g2_fill_1 FILLER_23_28 ();
 sg13g2_fill_1 FILLER_23_53 ();
 sg13g2_decap_4 FILLER_23_59 ();
 sg13g2_fill_1 FILLER_23_63 ();
 sg13g2_fill_2 FILLER_23_69 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_fill_2 FILLER_23_84 ();
 sg13g2_fill_1 FILLER_23_108 ();
 sg13g2_fill_2 FILLER_23_121 ();
 sg13g2_fill_1 FILLER_23_181 ();
 sg13g2_fill_1 FILLER_23_205 ();
 sg13g2_decap_4 FILLER_23_285 ();
 sg13g2_fill_1 FILLER_23_308 ();
 sg13g2_decap_4 FILLER_23_339 ();
 sg13g2_decap_4 FILLER_23_356 ();
 sg13g2_fill_1 FILLER_23_385 ();
 sg13g2_fill_1 FILLER_23_390 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_44 ();
 sg13g2_fill_2 FILLER_24_80 ();
 sg13g2_decap_4 FILLER_24_90 ();
 sg13g2_fill_1 FILLER_24_94 ();
 sg13g2_decap_4 FILLER_24_101 ();
 sg13g2_decap_8 FILLER_24_109 ();
 sg13g2_decap_8 FILLER_24_116 ();
 sg13g2_decap_8 FILLER_24_123 ();
 sg13g2_decap_4 FILLER_24_130 ();
 sg13g2_fill_1 FILLER_24_134 ();
 sg13g2_fill_2 FILLER_24_143 ();
 sg13g2_fill_1 FILLER_24_145 ();
 sg13g2_fill_1 FILLER_24_170 ();
 sg13g2_fill_2 FILLER_24_184 ();
 sg13g2_fill_1 FILLER_24_186 ();
 sg13g2_decap_8 FILLER_24_205 ();
 sg13g2_decap_4 FILLER_24_212 ();
 sg13g2_decap_8 FILLER_24_233 ();
 sg13g2_decap_8 FILLER_24_240 ();
 sg13g2_decap_8 FILLER_24_247 ();
 sg13g2_fill_2 FILLER_24_254 ();
 sg13g2_fill_2 FILLER_24_269 ();
 sg13g2_fill_1 FILLER_24_271 ();
 sg13g2_fill_1 FILLER_24_276 ();
 sg13g2_fill_2 FILLER_24_281 ();
 sg13g2_fill_2 FILLER_24_317 ();
 sg13g2_fill_2 FILLER_24_327 ();
 sg13g2_fill_1 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_fill_2 FILLER_24_350 ();
 sg13g2_fill_2 FILLER_24_377 ();
 sg13g2_fill_1 FILLER_24_379 ();
 sg13g2_fill_2 FILLER_24_390 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_27 ();
 sg13g2_fill_1 FILLER_25_59 ();
 sg13g2_decap_4 FILLER_25_110 ();
 sg13g2_decap_8 FILLER_25_124 ();
 sg13g2_decap_8 FILLER_25_131 ();
 sg13g2_decap_8 FILLER_25_138 ();
 sg13g2_fill_2 FILLER_25_145 ();
 sg13g2_fill_1 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_169 ();
 sg13g2_fill_1 FILLER_25_176 ();
 sg13g2_fill_2 FILLER_25_181 ();
 sg13g2_fill_1 FILLER_25_183 ();
 sg13g2_fill_2 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_206 ();
 sg13g2_decap_8 FILLER_25_213 ();
 sg13g2_decap_4 FILLER_25_220 ();
 sg13g2_fill_1 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_241 ();
 sg13g2_decap_8 FILLER_25_248 ();
 sg13g2_decap_8 FILLER_25_255 ();
 sg13g2_fill_1 FILLER_25_262 ();
 sg13g2_decap_8 FILLER_25_270 ();
 sg13g2_decap_8 FILLER_25_277 ();
 sg13g2_decap_4 FILLER_25_292 ();
 sg13g2_fill_2 FILLER_25_296 ();
 sg13g2_fill_2 FILLER_25_315 ();
 sg13g2_fill_1 FILLER_25_317 ();
 sg13g2_decap_8 FILLER_25_340 ();
 sg13g2_fill_1 FILLER_25_347 ();
 sg13g2_fill_2 FILLER_25_361 ();
 sg13g2_fill_1 FILLER_25_363 ();
 sg13g2_fill_2 FILLER_25_373 ();
 sg13g2_fill_1 FILLER_25_375 ();
 sg13g2_fill_1 FILLER_25_394 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_38 ();
 sg13g2_decap_8 FILLER_26_51 ();
 sg13g2_decap_8 FILLER_26_58 ();
 sg13g2_decap_4 FILLER_26_65 ();
 sg13g2_fill_1 FILLER_26_69 ();
 sg13g2_fill_2 FILLER_26_75 ();
 sg13g2_fill_1 FILLER_26_101 ();
 sg13g2_decap_4 FILLER_26_130 ();
 sg13g2_fill_1 FILLER_26_134 ();
 sg13g2_fill_1 FILLER_26_144 ();
 sg13g2_decap_8 FILLER_26_150 ();
 sg13g2_decap_4 FILLER_26_157 ();
 sg13g2_decap_8 FILLER_26_165 ();
 sg13g2_fill_2 FILLER_26_175 ();
 sg13g2_fill_1 FILLER_26_177 ();
 sg13g2_decap_8 FILLER_26_204 ();
 sg13g2_decap_4 FILLER_26_211 ();
 sg13g2_fill_2 FILLER_26_215 ();
 sg13g2_fill_1 FILLER_26_230 ();
 sg13g2_decap_4 FILLER_26_247 ();
 sg13g2_fill_1 FILLER_26_264 ();
 sg13g2_decap_8 FILLER_26_275 ();
 sg13g2_decap_8 FILLER_26_282 ();
 sg13g2_fill_2 FILLER_26_323 ();
 sg13g2_fill_1 FILLER_26_325 ();
 sg13g2_fill_1 FILLER_26_347 ();
 sg13g2_fill_2 FILLER_26_364 ();
 sg13g2_fill_1 FILLER_26_366 ();
 sg13g2_fill_1 FILLER_26_388 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_28 ();
 sg13g2_fill_1 FILLER_27_30 ();
 sg13g2_fill_1 FILLER_27_43 ();
 sg13g2_decap_8 FILLER_27_60 ();
 sg13g2_decap_8 FILLER_27_67 ();
 sg13g2_decap_8 FILLER_27_74 ();
 sg13g2_fill_2 FILLER_27_81 ();
 sg13g2_fill_1 FILLER_27_83 ();
 sg13g2_fill_1 FILLER_27_101 ();
 sg13g2_fill_2 FILLER_27_133 ();
 sg13g2_fill_1 FILLER_27_143 ();
 sg13g2_fill_2 FILLER_27_160 ();
 sg13g2_fill_1 FILLER_27_162 ();
 sg13g2_fill_1 FILLER_27_168 ();
 sg13g2_fill_1 FILLER_27_185 ();
 sg13g2_decap_4 FILLER_27_202 ();
 sg13g2_decap_4 FILLER_27_211 ();
 sg13g2_fill_1 FILLER_27_215 ();
 sg13g2_fill_1 FILLER_27_220 ();
 sg13g2_fill_1 FILLER_27_250 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_fill_2 FILLER_27_287 ();
 sg13g2_fill_1 FILLER_27_289 ();
 sg13g2_decap_4 FILLER_27_305 ();
 sg13g2_fill_1 FILLER_27_309 ();
 sg13g2_fill_2 FILLER_27_328 ();
 sg13g2_fill_1 FILLER_27_330 ();
 sg13g2_fill_2 FILLER_27_375 ();
 sg13g2_fill_1 FILLER_27_377 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_29 ();
 sg13g2_decap_8 FILLER_28_85 ();
 sg13g2_decap_8 FILLER_28_92 ();
 sg13g2_decap_8 FILLER_28_99 ();
 sg13g2_fill_1 FILLER_28_106 ();
 sg13g2_fill_2 FILLER_28_126 ();
 sg13g2_fill_2 FILLER_28_141 ();
 sg13g2_fill_1 FILLER_28_151 ();
 sg13g2_fill_1 FILLER_28_160 ();
 sg13g2_fill_1 FILLER_28_198 ();
 sg13g2_fill_2 FILLER_28_207 ();
 sg13g2_fill_1 FILLER_28_209 ();
 sg13g2_fill_2 FILLER_28_228 ();
 sg13g2_fill_1 FILLER_28_234 ();
 sg13g2_fill_1 FILLER_28_247 ();
 sg13g2_fill_1 FILLER_28_257 ();
 sg13g2_fill_2 FILLER_28_267 ();
 sg13g2_fill_1 FILLER_28_269 ();
 sg13g2_fill_1 FILLER_28_281 ();
 sg13g2_fill_1 FILLER_28_298 ();
 sg13g2_fill_1 FILLER_28_307 ();
 sg13g2_fill_2 FILLER_28_322 ();
 sg13g2_fill_1 FILLER_28_324 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_50 ();
 sg13g2_fill_1 FILLER_29_80 ();
 sg13g2_fill_2 FILLER_29_91 ();
 sg13g2_fill_1 FILLER_29_106 ();
 sg13g2_fill_2 FILLER_29_120 ();
 sg13g2_fill_1 FILLER_29_122 ();
 sg13g2_decap_8 FILLER_29_131 ();
 sg13g2_decap_4 FILLER_29_138 ();
 sg13g2_fill_2 FILLER_29_142 ();
 sg13g2_fill_2 FILLER_29_172 ();
 sg13g2_fill_1 FILLER_29_174 ();
 sg13g2_decap_4 FILLER_29_197 ();
 sg13g2_decap_8 FILLER_29_242 ();
 sg13g2_decap_4 FILLER_29_249 ();
 sg13g2_fill_2 FILLER_29_266 ();
 sg13g2_fill_1 FILLER_29_268 ();
 sg13g2_fill_1 FILLER_29_273 ();
 sg13g2_fill_2 FILLER_29_279 ();
 sg13g2_fill_1 FILLER_29_281 ();
 sg13g2_fill_2 FILLER_29_318 ();
 sg13g2_fill_1 FILLER_29_320 ();
 sg13g2_decap_4 FILLER_29_338 ();
 sg13g2_fill_1 FILLER_29_342 ();
 sg13g2_decap_8 FILLER_29_347 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_29 ();
 sg13g2_fill_1 FILLER_30_44 ();
 sg13g2_fill_2 FILLER_30_65 ();
 sg13g2_fill_2 FILLER_30_119 ();
 sg13g2_fill_1 FILLER_30_121 ();
 sg13g2_fill_2 FILLER_30_127 ();
 sg13g2_fill_1 FILLER_30_134 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_fill_1 FILLER_30_147 ();
 sg13g2_fill_2 FILLER_30_152 ();
 sg13g2_fill_1 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_165 ();
 sg13g2_decap_4 FILLER_30_172 ();
 sg13g2_fill_2 FILLER_30_176 ();
 sg13g2_fill_1 FILLER_30_183 ();
 sg13g2_decap_8 FILLER_30_188 ();
 sg13g2_fill_1 FILLER_30_195 ();
 sg13g2_fill_1 FILLER_30_213 ();
 sg13g2_fill_2 FILLER_30_227 ();
 sg13g2_decap_4 FILLER_30_246 ();
 sg13g2_fill_2 FILLER_30_250 ();
 sg13g2_fill_2 FILLER_30_269 ();
 sg13g2_fill_2 FILLER_30_291 ();
 sg13g2_fill_2 FILLER_30_306 ();
 sg13g2_fill_1 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_328 ();
 sg13g2_decap_8 FILLER_30_335 ();
 sg13g2_decap_8 FILLER_30_342 ();
 sg13g2_decap_8 FILLER_30_349 ();
 sg13g2_decap_4 FILLER_30_356 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_4 FILLER_31_12 ();
 sg13g2_decap_4 FILLER_31_25 ();
 sg13g2_decap_8 FILLER_31_41 ();
 sg13g2_decap_8 FILLER_31_48 ();
 sg13g2_decap_8 FILLER_31_55 ();
 sg13g2_fill_2 FILLER_31_62 ();
 sg13g2_fill_2 FILLER_31_93 ();
 sg13g2_fill_2 FILLER_31_120 ();
 sg13g2_fill_2 FILLER_31_130 ();
 sg13g2_fill_1 FILLER_31_132 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_fill_2 FILLER_31_180 ();
 sg13g2_decap_8 FILLER_31_215 ();
 sg13g2_decap_4 FILLER_31_222 ();
 sg13g2_fill_1 FILLER_31_240 ();
 sg13g2_decap_8 FILLER_31_275 ();
 sg13g2_fill_1 FILLER_31_282 ();
 sg13g2_decap_8 FILLER_31_300 ();
 sg13g2_fill_2 FILLER_31_307 ();
 sg13g2_fill_1 FILLER_31_309 ();
 sg13g2_decap_8 FILLER_31_320 ();
 sg13g2_decap_8 FILLER_31_327 ();
 sg13g2_fill_1 FILLER_31_334 ();
 sg13g2_fill_1 FILLER_31_363 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_4 FILLER_32_14 ();
 sg13g2_fill_2 FILLER_32_18 ();
 sg13g2_fill_2 FILLER_32_35 ();
 sg13g2_fill_1 FILLER_32_37 ();
 sg13g2_decap_8 FILLER_32_59 ();
 sg13g2_decap_8 FILLER_32_66 ();
 sg13g2_decap_8 FILLER_32_73 ();
 sg13g2_fill_1 FILLER_32_110 ();
 sg13g2_fill_2 FILLER_32_133 ();
 sg13g2_fill_1 FILLER_32_135 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_fill_2 FILLER_32_147 ();
 sg13g2_fill_1 FILLER_32_149 ();
 sg13g2_fill_2 FILLER_32_153 ();
 sg13g2_fill_1 FILLER_32_155 ();
 sg13g2_decap_4 FILLER_32_161 ();
 sg13g2_fill_1 FILLER_32_193 ();
 sg13g2_decap_8 FILLER_32_231 ();
 sg13g2_decap_4 FILLER_32_238 ();
 sg13g2_fill_2 FILLER_32_242 ();
 sg13g2_fill_2 FILLER_32_258 ();
 sg13g2_decap_8 FILLER_32_273 ();
 sg13g2_fill_2 FILLER_32_285 ();
 sg13g2_fill_1 FILLER_32_287 ();
 sg13g2_decap_8 FILLER_32_292 ();
 sg13g2_fill_1 FILLER_32_299 ();
 sg13g2_decap_8 FILLER_32_310 ();
 sg13g2_decap_8 FILLER_32_317 ();
 sg13g2_decap_4 FILLER_32_324 ();
 sg13g2_decap_8 FILLER_32_341 ();
 sg13g2_fill_1 FILLER_32_348 ();
 sg13g2_decap_4 FILLER_32_364 ();
 sg13g2_fill_2 FILLER_32_368 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_29 ();
 sg13g2_fill_1 FILLER_33_31 ();
 sg13g2_fill_2 FILLER_33_56 ();
 sg13g2_fill_1 FILLER_33_58 ();
 sg13g2_decap_8 FILLER_33_95 ();
 sg13g2_decap_4 FILLER_33_102 ();
 sg13g2_fill_1 FILLER_33_106 ();
 sg13g2_fill_1 FILLER_33_116 ();
 sg13g2_decap_8 FILLER_33_131 ();
 sg13g2_decap_8 FILLER_33_138 ();
 sg13g2_decap_8 FILLER_33_173 ();
 sg13g2_decap_8 FILLER_33_180 ();
 sg13g2_decap_8 FILLER_33_187 ();
 sg13g2_decap_8 FILLER_33_194 ();
 sg13g2_fill_2 FILLER_33_201 ();
 sg13g2_fill_1 FILLER_33_203 ();
 sg13g2_decap_4 FILLER_33_217 ();
 sg13g2_fill_2 FILLER_33_221 ();
 sg13g2_decap_8 FILLER_33_251 ();
 sg13g2_decap_8 FILLER_33_289 ();
 sg13g2_decap_8 FILLER_33_296 ();
 sg13g2_decap_4 FILLER_33_303 ();
 sg13g2_fill_2 FILLER_33_340 ();
 sg13g2_fill_2 FILLER_33_370 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_fill_1 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_29 ();
 sg13g2_fill_2 FILLER_34_43 ();
 sg13g2_decap_8 FILLER_34_73 ();
 sg13g2_decap_8 FILLER_34_80 ();
 sg13g2_decap_8 FILLER_34_87 ();
 sg13g2_decap_8 FILLER_34_94 ();
 sg13g2_decap_8 FILLER_34_101 ();
 sg13g2_decap_8 FILLER_34_108 ();
 sg13g2_decap_4 FILLER_34_115 ();
 sg13g2_decap_8 FILLER_34_124 ();
 sg13g2_decap_8 FILLER_34_131 ();
 sg13g2_decap_8 FILLER_34_138 ();
 sg13g2_decap_8 FILLER_34_145 ();
 sg13g2_decap_8 FILLER_34_152 ();
 sg13g2_decap_4 FILLER_34_159 ();
 sg13g2_fill_1 FILLER_34_163 ();
 sg13g2_decap_8 FILLER_34_170 ();
 sg13g2_decap_8 FILLER_34_177 ();
 sg13g2_decap_8 FILLER_34_184 ();
 sg13g2_decap_8 FILLER_34_191 ();
 sg13g2_decap_8 FILLER_34_198 ();
 sg13g2_decap_8 FILLER_34_205 ();
 sg13g2_decap_4 FILLER_34_212 ();
 sg13g2_fill_2 FILLER_34_216 ();
 sg13g2_fill_2 FILLER_34_246 ();
 sg13g2_decap_8 FILLER_34_253 ();
 sg13g2_fill_1 FILLER_34_260 ();
 sg13g2_fill_2 FILLER_34_307 ();
 sg13g2_decap_8 FILLER_34_336 ();
 sg13g2_fill_1 FILLER_34_380 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_7 ();
 sg13g2_fill_1 FILLER_35_43 ();
 sg13g2_fill_1 FILLER_35_58 ();
 sg13g2_fill_2 FILLER_35_95 ();
 sg13g2_decap_8 FILLER_35_101 ();
 sg13g2_decap_8 FILLER_35_108 ();
 sg13g2_decap_4 FILLER_35_131 ();
 sg13g2_fill_2 FILLER_35_141 ();
 sg13g2_fill_1 FILLER_35_143 ();
 sg13g2_fill_2 FILLER_35_152 ();
 sg13g2_fill_2 FILLER_35_167 ();
 sg13g2_fill_1 FILLER_35_188 ();
 sg13g2_decap_8 FILLER_35_194 ();
 sg13g2_decap_8 FILLER_35_201 ();
 sg13g2_decap_8 FILLER_35_208 ();
 sg13g2_decap_4 FILLER_35_215 ();
 sg13g2_fill_2 FILLER_35_219 ();
 sg13g2_fill_2 FILLER_35_234 ();
 sg13g2_fill_1 FILLER_35_236 ();
 sg13g2_fill_2 FILLER_35_282 ();
 sg13g2_decap_8 FILLER_35_297 ();
 sg13g2_fill_2 FILLER_35_304 ();
 sg13g2_fill_1 FILLER_35_306 ();
 sg13g2_fill_2 FILLER_35_326 ();
 sg13g2_fill_1 FILLER_35_328 ();
 sg13g2_decap_4 FILLER_35_357 ();
 sg13g2_fill_1 FILLER_35_374 ();
 sg13g2_decap_4 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_4 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_11 ();
 sg13g2_fill_1 FILLER_36_36 ();
 sg13g2_fill_2 FILLER_36_51 ();
 sg13g2_fill_1 FILLER_36_53 ();
 sg13g2_decap_8 FILLER_36_76 ();
 sg13g2_fill_1 FILLER_36_83 ();
 sg13g2_fill_2 FILLER_36_117 ();
 sg13g2_decap_4 FILLER_36_176 ();
 sg13g2_decap_8 FILLER_36_218 ();
 sg13g2_decap_8 FILLER_36_225 ();
 sg13g2_fill_1 FILLER_36_232 ();
 sg13g2_fill_2 FILLER_36_272 ();
 sg13g2_fill_2 FILLER_36_314 ();
 sg13g2_fill_1 FILLER_36_347 ();
 sg13g2_fill_2 FILLER_36_374 ();
 sg13g2_fill_2 FILLER_37_27 ();
 sg13g2_fill_1 FILLER_37_50 ();
 sg13g2_fill_2 FILLER_37_105 ();
 sg13g2_fill_1 FILLER_37_151 ();
 sg13g2_fill_2 FILLER_37_165 ();
 sg13g2_fill_1 FILLER_37_177 ();
 sg13g2_fill_2 FILLER_37_185 ();
 sg13g2_fill_1 FILLER_37_187 ();
 sg13g2_fill_2 FILLER_37_226 ();
 sg13g2_fill_1 FILLER_37_228 ();
 sg13g2_fill_2 FILLER_37_234 ();
 sg13g2_fill_1 FILLER_37_236 ();
 sg13g2_fill_2 FILLER_37_246 ();
 sg13g2_fill_1 FILLER_37_248 ();
 sg13g2_fill_2 FILLER_37_272 ();
 sg13g2_decap_4 FILLER_37_288 ();
 sg13g2_fill_1 FILLER_37_292 ();
 sg13g2_fill_2 FILLER_37_297 ();
 sg13g2_fill_1 FILLER_37_299 ();
 sg13g2_fill_2 FILLER_37_321 ();
 sg13g2_decap_4 FILLER_37_360 ();
 sg13g2_fill_1 FILLER_37_364 ();
 sg13g2_fill_1 FILLER_37_383 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_fill_1 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_73 ();
 sg13g2_decap_8 FILLER_38_80 ();
 sg13g2_fill_1 FILLER_38_91 ();
 sg13g2_fill_2 FILLER_38_115 ();
 sg13g2_fill_2 FILLER_38_126 ();
 sg13g2_fill_1 FILLER_38_128 ();
 sg13g2_fill_1 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_142 ();
 sg13g2_decap_8 FILLER_38_149 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_fill_1 FILLER_38_160 ();
 sg13g2_fill_1 FILLER_38_176 ();
 sg13g2_fill_2 FILLER_38_208 ();
 sg13g2_fill_2 FILLER_38_269 ();
 sg13g2_fill_1 FILLER_38_271 ();
 sg13g2_fill_1 FILLER_38_366 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_7 ();
 sg13g2_fill_2 FILLER_39_35 ();
 sg13g2_fill_1 FILLER_39_37 ();
 sg13g2_fill_1 FILLER_39_85 ();
 sg13g2_fill_2 FILLER_39_101 ();
 sg13g2_fill_2 FILLER_39_116 ();
 sg13g2_fill_1 FILLER_39_123 ();
 sg13g2_decap_8 FILLER_39_132 ();
 sg13g2_decap_4 FILLER_39_139 ();
 sg13g2_fill_2 FILLER_39_147 ();
 sg13g2_fill_2 FILLER_39_159 ();
 sg13g2_fill_2 FILLER_39_181 ();
 sg13g2_decap_8 FILLER_39_191 ();
 sg13g2_decap_4 FILLER_39_198 ();
 sg13g2_fill_2 FILLER_39_211 ();
 sg13g2_fill_1 FILLER_39_213 ();
 sg13g2_fill_2 FILLER_39_228 ();
 sg13g2_fill_1 FILLER_39_230 ();
 sg13g2_fill_2 FILLER_39_240 ();
 sg13g2_fill_2 FILLER_39_257 ();
 sg13g2_fill_1 FILLER_39_259 ();
 sg13g2_fill_1 FILLER_39_280 ();
 sg13g2_decap_8 FILLER_39_348 ();
 sg13g2_fill_2 FILLER_39_355 ();
 sg13g2_fill_1 FILLER_39_363 ();
 sg13g2_decap_4 FILLER_39_369 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_fill_1 FILLER_40_14 ();
 sg13g2_decap_4 FILLER_40_27 ();
 sg13g2_fill_1 FILLER_40_46 ();
 sg13g2_fill_1 FILLER_40_65 ();
 sg13g2_fill_2 FILLER_40_103 ();
 sg13g2_fill_1 FILLER_40_105 ();
 sg13g2_fill_2 FILLER_40_111 ();
 sg13g2_fill_1 FILLER_40_113 ();
 sg13g2_fill_1 FILLER_40_119 ();
 sg13g2_fill_2 FILLER_40_134 ();
 sg13g2_fill_1 FILLER_40_136 ();
 sg13g2_fill_2 FILLER_40_156 ();
 sg13g2_fill_2 FILLER_40_168 ();
 sg13g2_fill_1 FILLER_40_170 ();
 sg13g2_fill_2 FILLER_40_177 ();
 sg13g2_fill_1 FILLER_40_179 ();
 sg13g2_fill_2 FILLER_40_225 ();
 sg13g2_fill_1 FILLER_40_227 ();
 sg13g2_fill_2 FILLER_40_237 ();
 sg13g2_fill_1 FILLER_40_239 ();
 sg13g2_fill_2 FILLER_40_250 ();
 sg13g2_fill_1 FILLER_40_252 ();
 sg13g2_fill_2 FILLER_40_258 ();
 sg13g2_fill_1 FILLER_40_273 ();
 sg13g2_fill_2 FILLER_40_284 ();
 sg13g2_fill_2 FILLER_40_310 ();
 sg13g2_fill_1 FILLER_40_312 ();
 sg13g2_fill_1 FILLER_40_318 ();
 sg13g2_decap_8 FILLER_40_338 ();
 sg13g2_decap_8 FILLER_40_345 ();
 sg13g2_fill_2 FILLER_40_352 ();
 sg13g2_fill_1 FILLER_40_362 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_fill_2 FILLER_41_21 ();
 sg13g2_fill_1 FILLER_41_23 ();
 sg13g2_fill_2 FILLER_41_45 ();
 sg13g2_fill_1 FILLER_41_47 ();
 sg13g2_fill_1 FILLER_41_80 ();
 sg13g2_fill_2 FILLER_41_94 ();
 sg13g2_fill_1 FILLER_41_113 ();
 sg13g2_fill_1 FILLER_41_147 ();
 sg13g2_fill_2 FILLER_41_158 ();
 sg13g2_fill_1 FILLER_41_160 ();
 sg13g2_fill_2 FILLER_41_204 ();
 sg13g2_fill_1 FILLER_41_206 ();
 sg13g2_fill_2 FILLER_41_211 ();
 sg13g2_fill_2 FILLER_41_226 ();
 sg13g2_fill_2 FILLER_41_256 ();
 sg13g2_fill_1 FILLER_41_258 ();
 sg13g2_fill_2 FILLER_41_271 ();
 sg13g2_fill_1 FILLER_41_273 ();
 sg13g2_fill_2 FILLER_41_279 ();
 sg13g2_fill_2 FILLER_41_291 ();
 sg13g2_fill_1 FILLER_41_293 ();
 sg13g2_fill_2 FILLER_41_299 ();
 sg13g2_fill_2 FILLER_41_307 ();
 sg13g2_fill_1 FILLER_41_309 ();
 sg13g2_fill_2 FILLER_41_323 ();
 sg13g2_decap_4 FILLER_41_334 ();
 sg13g2_fill_2 FILLER_41_338 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_2 ();
 sg13g2_decap_8 FILLER_42_80 ();
 sg13g2_decap_8 FILLER_42_115 ();
 sg13g2_fill_2 FILLER_42_134 ();
 sg13g2_fill_1 FILLER_42_142 ();
 sg13g2_fill_2 FILLER_42_152 ();
 sg13g2_fill_1 FILLER_42_154 ();
 sg13g2_decap_4 FILLER_42_163 ();
 sg13g2_fill_1 FILLER_42_167 ();
 sg13g2_decap_4 FILLER_42_186 ();
 sg13g2_decap_4 FILLER_42_246 ();
 sg13g2_fill_1 FILLER_42_250 ();
 sg13g2_fill_2 FILLER_42_281 ();
 sg13g2_fill_1 FILLER_42_283 ();
 sg13g2_fill_2 FILLER_42_288 ();
 sg13g2_fill_1 FILLER_42_290 ();
 sg13g2_fill_2 FILLER_42_308 ();
 sg13g2_fill_1 FILLER_42_310 ();
 sg13g2_decap_4 FILLER_42_319 ();
 sg13g2_decap_8 FILLER_42_327 ();
 sg13g2_decap_4 FILLER_42_334 ();
 sg13g2_fill_1 FILLER_42_338 ();
 sg13g2_fill_2 FILLER_42_344 ();
 sg13g2_decap_8 FILLER_42_354 ();
 sg13g2_fill_1 FILLER_42_361 ();
 sg13g2_fill_1 FILLER_42_380 ();
 sg13g2_fill_2 FILLER_42_395 ();
 sg13g2_fill_2 FILLER_42_406 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_fill_2 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_2 ();
 sg13g2_fill_1 FILLER_43_27 ();
 sg13g2_fill_1 FILLER_43_37 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_128 ();
 sg13g2_decap_8 FILLER_43_135 ();
 sg13g2_decap_8 FILLER_43_155 ();
 sg13g2_decap_8 FILLER_43_162 ();
 sg13g2_fill_2 FILLER_43_169 ();
 sg13g2_fill_1 FILLER_43_171 ();
 sg13g2_decap_8 FILLER_43_184 ();
 sg13g2_decap_8 FILLER_43_191 ();
 sg13g2_fill_2 FILLER_43_198 ();
 sg13g2_decap_4 FILLER_43_208 ();
 sg13g2_fill_2 FILLER_43_212 ();
 sg13g2_decap_4 FILLER_43_218 ();
 sg13g2_fill_2 FILLER_43_222 ();
 sg13g2_fill_2 FILLER_43_234 ();
 sg13g2_decap_4 FILLER_43_240 ();
 sg13g2_fill_2 FILLER_43_244 ();
 sg13g2_decap_8 FILLER_43_257 ();
 sg13g2_decap_8 FILLER_43_264 ();
 sg13g2_decap_8 FILLER_43_271 ();
 sg13g2_decap_8 FILLER_43_278 ();
 sg13g2_decap_8 FILLER_43_285 ();
 sg13g2_decap_8 FILLER_43_292 ();
 sg13g2_fill_1 FILLER_43_303 ();
 sg13g2_fill_2 FILLER_43_322 ();
 sg13g2_fill_1 FILLER_43_324 ();
 sg13g2_decap_4 FILLER_43_343 ();
 sg13g2_decap_8 FILLER_43_357 ();
 sg13g2_fill_2 FILLER_43_364 ();
 sg13g2_fill_2 FILLER_43_398 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_2 ();
 sg13g2_decap_4 FILLER_44_31 ();
 sg13g2_decap_8 FILLER_44_88 ();
 sg13g2_decap_8 FILLER_44_95 ();
 sg13g2_decap_8 FILLER_44_102 ();
 sg13g2_decap_8 FILLER_44_109 ();
 sg13g2_decap_4 FILLER_44_116 ();
 sg13g2_decap_8 FILLER_44_124 ();
 sg13g2_decap_8 FILLER_44_131 ();
 sg13g2_decap_8 FILLER_44_138 ();
 sg13g2_fill_2 FILLER_44_145 ();
 sg13g2_fill_1 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_153 ();
 sg13g2_decap_8 FILLER_44_160 ();
 sg13g2_decap_8 FILLER_44_167 ();
 sg13g2_decap_8 FILLER_44_174 ();
 sg13g2_fill_1 FILLER_44_181 ();
 sg13g2_decap_8 FILLER_44_187 ();
 sg13g2_decap_8 FILLER_44_194 ();
 sg13g2_decap_8 FILLER_44_201 ();
 sg13g2_decap_8 FILLER_44_214 ();
 sg13g2_decap_8 FILLER_44_221 ();
 sg13g2_fill_2 FILLER_44_228 ();
 sg13g2_fill_1 FILLER_44_230 ();
 sg13g2_decap_8 FILLER_44_238 ();
 sg13g2_decap_8 FILLER_44_245 ();
 sg13g2_fill_2 FILLER_44_252 ();
 sg13g2_decap_8 FILLER_44_267 ();
 sg13g2_decap_4 FILLER_44_274 ();
 sg13g2_fill_1 FILLER_44_278 ();
 sg13g2_decap_8 FILLER_44_284 ();
 sg13g2_fill_2 FILLER_44_291 ();
 sg13g2_fill_1 FILLER_44_293 ();
 sg13g2_decap_4 FILLER_44_299 ();
 sg13g2_decap_4 FILLER_44_307 ();
 sg13g2_fill_2 FILLER_44_311 ();
 sg13g2_fill_1 FILLER_44_327 ();
 sg13g2_fill_1 FILLER_44_333 ();
 sg13g2_fill_2 FILLER_44_372 ();
 sg13g2_fill_1 FILLER_44_374 ();
 sg13g2_decap_8 FILLER_44_402 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_4 FILLER_45_14 ();
 sg13g2_fill_1 FILLER_45_18 ();
 sg13g2_fill_2 FILLER_45_72 ();
 sg13g2_fill_2 FILLER_45_113 ();
 sg13g2_fill_1 FILLER_45_115 ();
 sg13g2_decap_8 FILLER_45_134 ();
 sg13g2_fill_1 FILLER_45_141 ();
 sg13g2_fill_1 FILLER_45_160 ();
 sg13g2_decap_4 FILLER_45_166 ();
 sg13g2_fill_2 FILLER_45_197 ();
 sg13g2_fill_1 FILLER_45_199 ();
 sg13g2_fill_2 FILLER_45_213 ();
 sg13g2_decap_8 FILLER_45_219 ();
 sg13g2_fill_2 FILLER_45_226 ();
 sg13g2_decap_4 FILLER_45_242 ();
 sg13g2_fill_2 FILLER_45_246 ();
 sg13g2_fill_1 FILLER_45_271 ();
 sg13g2_fill_2 FILLER_45_308 ();
 sg13g2_fill_1 FILLER_45_310 ();
 sg13g2_fill_2 FILLER_45_318 ();
 sg13g2_fill_1 FILLER_45_320 ();
 sg13g2_fill_2 FILLER_45_339 ();
 sg13g2_fill_1 FILLER_45_341 ();
 sg13g2_decap_8 FILLER_45_366 ();
 sg13g2_fill_2 FILLER_45_378 ();
 sg13g2_fill_1 FILLER_45_380 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_4 FILLER_46_14 ();
 sg13g2_fill_1 FILLER_46_18 ();
 sg13g2_fill_1 FILLER_46_40 ();
 sg13g2_decap_4 FILLER_46_45 ();
 sg13g2_fill_1 FILLER_46_127 ();
 sg13g2_fill_1 FILLER_46_144 ();
 sg13g2_fill_2 FILLER_46_219 ();
 sg13g2_fill_1 FILLER_46_221 ();
 sg13g2_fill_2 FILLER_46_248 ();
 sg13g2_fill_1 FILLER_46_261 ();
 sg13g2_decap_4 FILLER_46_270 ();
 sg13g2_fill_2 FILLER_46_303 ();
 sg13g2_fill_2 FILLER_46_326 ();
 sg13g2_decap_4 FILLER_46_341 ();
 sg13g2_decap_8 FILLER_46_361 ();
 sg13g2_fill_2 FILLER_46_368 ();
 sg13g2_fill_1 FILLER_46_370 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_4 FILLER_47_7 ();
 sg13g2_fill_1 FILLER_47_38 ();
 sg13g2_fill_2 FILLER_47_61 ();
 sg13g2_fill_2 FILLER_47_72 ();
 sg13g2_fill_2 FILLER_47_87 ();
 sg13g2_fill_1 FILLER_47_89 ();
 sg13g2_fill_1 FILLER_47_136 ();
 sg13g2_fill_2 FILLER_47_145 ();
 sg13g2_fill_1 FILLER_47_147 ();
 sg13g2_decap_4 FILLER_47_171 ();
 sg13g2_fill_2 FILLER_47_200 ();
 sg13g2_fill_1 FILLER_47_235 ();
 sg13g2_fill_2 FILLER_47_244 ();
 sg13g2_fill_1 FILLER_47_285 ();
 sg13g2_fill_1 FILLER_47_310 ();
 sg13g2_decap_8 FILLER_47_315 ();
 sg13g2_decap_8 FILLER_47_336 ();
 sg13g2_decap_8 FILLER_47_343 ();
 sg13g2_fill_2 FILLER_47_350 ();
 sg13g2_fill_1 FILLER_47_352 ();
 sg13g2_decap_4 FILLER_47_361 ();
 sg13g2_fill_2 FILLER_47_370 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_4 FILLER_48_28 ();
 sg13g2_fill_1 FILLER_48_36 ();
 sg13g2_fill_2 FILLER_48_51 ();
 sg13g2_fill_1 FILLER_48_53 ();
 sg13g2_decap_8 FILLER_48_67 ();
 sg13g2_decap_4 FILLER_48_74 ();
 sg13g2_fill_1 FILLER_48_78 ();
 sg13g2_fill_2 FILLER_48_83 ();
 sg13g2_fill_2 FILLER_48_90 ();
 sg13g2_decap_8 FILLER_48_100 ();
 sg13g2_decap_4 FILLER_48_107 ();
 sg13g2_fill_1 FILLER_48_111 ();
 sg13g2_fill_2 FILLER_48_116 ();
 sg13g2_fill_2 FILLER_48_122 ();
 sg13g2_decap_4 FILLER_48_173 ();
 sg13g2_decap_8 FILLER_48_197 ();
 sg13g2_decap_4 FILLER_48_204 ();
 sg13g2_fill_1 FILLER_48_208 ();
 sg13g2_fill_2 FILLER_48_224 ();
 sg13g2_fill_2 FILLER_48_247 ();
 sg13g2_fill_1 FILLER_48_249 ();
 sg13g2_decap_4 FILLER_48_255 ();
 sg13g2_fill_2 FILLER_48_259 ();
 sg13g2_decap_8 FILLER_48_271 ();
 sg13g2_fill_1 FILLER_48_278 ();
 sg13g2_decap_8 FILLER_48_284 ();
 sg13g2_decap_4 FILLER_48_291 ();
 sg13g2_fill_2 FILLER_48_295 ();
 sg13g2_decap_8 FILLER_48_309 ();
 sg13g2_decap_4 FILLER_48_316 ();
 sg13g2_decap_8 FILLER_48_337 ();
 sg13g2_decap_4 FILLER_48_344 ();
 sg13g2_fill_2 FILLER_48_348 ();
 sg13g2_fill_2 FILLER_48_397 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_fill_2 FILLER_49_14 ();
 sg13g2_fill_1 FILLER_49_16 ();
 sg13g2_decap_8 FILLER_49_72 ();
 sg13g2_fill_1 FILLER_49_79 ();
 sg13g2_decap_8 FILLER_49_93 ();
 sg13g2_decap_4 FILLER_49_100 ();
 sg13g2_decap_4 FILLER_49_131 ();
 sg13g2_fill_2 FILLER_49_135 ();
 sg13g2_fill_2 FILLER_49_170 ();
 sg13g2_fill_1 FILLER_49_172 ();
 sg13g2_fill_2 FILLER_49_180 ();
 sg13g2_decap_8 FILLER_49_185 ();
 sg13g2_decap_8 FILLER_49_192 ();
 sg13g2_fill_2 FILLER_49_199 ();
 sg13g2_decap_8 FILLER_49_218 ();
 sg13g2_decap_4 FILLER_49_225 ();
 sg13g2_fill_2 FILLER_49_233 ();
 sg13g2_decap_4 FILLER_49_243 ();
 sg13g2_fill_1 FILLER_49_255 ();
 sg13g2_decap_8 FILLER_49_284 ();
 sg13g2_decap_4 FILLER_49_314 ();
 sg13g2_fill_2 FILLER_49_350 ();
 sg13g2_fill_1 FILLER_49_352 ();
 sg13g2_fill_1 FILLER_49_369 ();
 sg13g2_fill_2 FILLER_49_406 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_4 FILLER_50_21 ();
 sg13g2_fill_1 FILLER_50_25 ();
 sg13g2_fill_1 FILLER_50_88 ();
 sg13g2_fill_2 FILLER_50_104 ();
 sg13g2_fill_1 FILLER_50_106 ();
 sg13g2_decap_8 FILLER_50_139 ();
 sg13g2_decap_8 FILLER_50_146 ();
 sg13g2_fill_1 FILLER_50_153 ();
 sg13g2_fill_2 FILLER_50_159 ();
 sg13g2_decap_8 FILLER_50_168 ();
 sg13g2_decap_8 FILLER_50_175 ();
 sg13g2_decap_8 FILLER_50_182 ();
 sg13g2_decap_8 FILLER_50_189 ();
 sg13g2_fill_2 FILLER_50_196 ();
 sg13g2_fill_1 FILLER_50_198 ();
 sg13g2_decap_8 FILLER_50_226 ();
 sg13g2_decap_4 FILLER_50_233 ();
 sg13g2_decap_8 FILLER_50_241 ();
 sg13g2_decap_8 FILLER_50_248 ();
 sg13g2_decap_4 FILLER_50_255 ();
 sg13g2_decap_8 FILLER_50_268 ();
 sg13g2_fill_1 FILLER_50_275 ();
 sg13g2_fill_1 FILLER_50_281 ();
 sg13g2_fill_1 FILLER_50_294 ();
 sg13g2_decap_8 FILLER_50_308 ();
 sg13g2_decap_8 FILLER_50_315 ();
 sg13g2_fill_2 FILLER_50_322 ();
 sg13g2_fill_1 FILLER_50_324 ();
 sg13g2_fill_1 FILLER_50_341 ();
 sg13g2_fill_2 FILLER_50_357 ();
 sg13g2_decap_4 FILLER_50_364 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_7 ();
 sg13g2_fill_2 FILLER_51_36 ();
 sg13g2_fill_1 FILLER_51_79 ();
 sg13g2_decap_8 FILLER_51_129 ();
 sg13g2_decap_8 FILLER_51_136 ();
 sg13g2_decap_8 FILLER_51_143 ();
 sg13g2_decap_8 FILLER_51_150 ();
 sg13g2_decap_8 FILLER_51_157 ();
 sg13g2_decap_8 FILLER_51_164 ();
 sg13g2_decap_4 FILLER_51_171 ();
 sg13g2_fill_2 FILLER_51_175 ();
 sg13g2_decap_8 FILLER_51_198 ();
 sg13g2_fill_2 FILLER_51_205 ();
 sg13g2_fill_1 FILLER_51_207 ();
 sg13g2_fill_2 FILLER_51_213 ();
 sg13g2_decap_8 FILLER_51_220 ();
 sg13g2_decap_8 FILLER_51_227 ();
 sg13g2_fill_1 FILLER_51_239 ();
 sg13g2_fill_1 FILLER_51_244 ();
 sg13g2_decap_8 FILLER_51_253 ();
 sg13g2_fill_2 FILLER_51_260 ();
 sg13g2_fill_1 FILLER_51_262 ();
 sg13g2_decap_8 FILLER_51_267 ();
 sg13g2_decap_4 FILLER_51_282 ();
 sg13g2_fill_1 FILLER_51_286 ();
 sg13g2_decap_4 FILLER_51_300 ();
 sg13g2_fill_2 FILLER_51_304 ();
 sg13g2_decap_4 FILLER_51_318 ();
 sg13g2_fill_1 FILLER_51_322 ();
 sg13g2_decap_8 FILLER_51_336 ();
 sg13g2_decap_8 FILLER_51_351 ();
 sg13g2_decap_8 FILLER_51_358 ();
 sg13g2_decap_4 FILLER_51_365 ();
 sg13g2_decap_8 FILLER_51_378 ();
 sg13g2_fill_2 FILLER_51_385 ();
 sg13g2_fill_1 FILLER_51_387 ();
 sg13g2_decap_8 FILLER_51_401 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_4 FILLER_52_14 ();
 sg13g2_fill_2 FILLER_52_18 ();
 sg13g2_fill_1 FILLER_52_29 ();
 sg13g2_decap_4 FILLER_52_39 ();
 sg13g2_fill_2 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_108 ();
 sg13g2_fill_1 FILLER_52_119 ();
 sg13g2_decap_8 FILLER_52_124 ();
 sg13g2_decap_8 FILLER_52_131 ();
 sg13g2_fill_2 FILLER_52_138 ();
 sg13g2_fill_1 FILLER_52_140 ();
 sg13g2_decap_4 FILLER_52_149 ();
 sg13g2_fill_2 FILLER_52_153 ();
 sg13g2_fill_2 FILLER_52_160 ();
 sg13g2_fill_2 FILLER_52_175 ();
 sg13g2_fill_1 FILLER_52_177 ();
 sg13g2_fill_2 FILLER_52_188 ();
 sg13g2_fill_1 FILLER_52_190 ();
 sg13g2_fill_1 FILLER_52_195 ();
 sg13g2_decap_8 FILLER_52_203 ();
 sg13g2_decap_4 FILLER_52_223 ();
 sg13g2_fill_2 FILLER_52_227 ();
 sg13g2_fill_2 FILLER_52_245 ();
 sg13g2_fill_1 FILLER_52_247 ();
 sg13g2_decap_8 FILLER_52_270 ();
 sg13g2_decap_4 FILLER_52_277 ();
 sg13g2_decap_4 FILLER_52_285 ();
 sg13g2_fill_2 FILLER_52_289 ();
 sg13g2_decap_4 FILLER_52_304 ();
 sg13g2_fill_1 FILLER_52_308 ();
 sg13g2_fill_1 FILLER_52_314 ();
 sg13g2_decap_8 FILLER_52_333 ();
 sg13g2_decap_4 FILLER_52_340 ();
 sg13g2_fill_2 FILLER_52_344 ();
 sg13g2_decap_8 FILLER_52_354 ();
 sg13g2_fill_2 FILLER_52_389 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_fill_2 FILLER_53_14 ();
 sg13g2_fill_1 FILLER_53_16 ();
 sg13g2_fill_1 FILLER_53_26 ();
 sg13g2_fill_2 FILLER_53_50 ();
 sg13g2_fill_1 FILLER_53_52 ();
 sg13g2_decap_4 FILLER_53_76 ();
 sg13g2_fill_2 FILLER_53_85 ();
 sg13g2_fill_1 FILLER_53_87 ();
 sg13g2_decap_8 FILLER_53_105 ();
 sg13g2_decap_8 FILLER_53_112 ();
 sg13g2_fill_1 FILLER_53_119 ();
 sg13g2_fill_1 FILLER_53_124 ();
 sg13g2_fill_1 FILLER_53_130 ();
 sg13g2_decap_4 FILLER_53_144 ();
 sg13g2_fill_2 FILLER_53_159 ();
 sg13g2_fill_1 FILLER_53_161 ();
 sg13g2_decap_8 FILLER_53_189 ();
 sg13g2_decap_8 FILLER_53_196 ();
 sg13g2_fill_1 FILLER_53_244 ();
 sg13g2_decap_4 FILLER_53_256 ();
 sg13g2_fill_1 FILLER_53_260 ();
 sg13g2_decap_4 FILLER_53_269 ();
 sg13g2_fill_1 FILLER_53_273 ();
 sg13g2_fill_1 FILLER_53_290 ();
 sg13g2_fill_2 FILLER_53_304 ();
 sg13g2_fill_1 FILLER_53_306 ();
 sg13g2_decap_8 FILLER_53_327 ();
 sg13g2_fill_2 FILLER_53_334 ();
 sg13g2_fill_2 FILLER_53_355 ();
 sg13g2_fill_1 FILLER_53_402 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_decap_4 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_63 ();
 sg13g2_fill_1 FILLER_54_65 ();
 sg13g2_fill_2 FILLER_54_76 ();
 sg13g2_decap_8 FILLER_54_92 ();
 sg13g2_fill_2 FILLER_54_99 ();
 sg13g2_fill_1 FILLER_54_101 ();
 sg13g2_decap_4 FILLER_54_107 ();
 sg13g2_fill_1 FILLER_54_111 ();
 sg13g2_fill_2 FILLER_54_157 ();
 sg13g2_fill_2 FILLER_54_167 ();
 sg13g2_fill_2 FILLER_54_179 ();
 sg13g2_fill_2 FILLER_54_197 ();
 sg13g2_fill_1 FILLER_54_220 ();
 sg13g2_fill_1 FILLER_54_238 ();
 sg13g2_fill_2 FILLER_54_258 ();
 sg13g2_fill_1 FILLER_54_260 ();
 sg13g2_fill_1 FILLER_54_277 ();
 sg13g2_fill_1 FILLER_54_304 ();
 sg13g2_fill_1 FILLER_54_318 ();
 sg13g2_fill_2 FILLER_54_333 ();
 sg13g2_fill_1 FILLER_54_335 ();
 sg13g2_fill_2 FILLER_54_345 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_fill_2 FILLER_55_57 ();
 sg13g2_fill_1 FILLER_55_59 ();
 sg13g2_fill_1 FILLER_55_69 ();
 sg13g2_fill_2 FILLER_55_88 ();
 sg13g2_fill_2 FILLER_55_106 ();
 sg13g2_fill_1 FILLER_55_108 ();
 sg13g2_fill_2 FILLER_55_130 ();
 sg13g2_fill_2 FILLER_55_172 ();
 sg13g2_fill_2 FILLER_55_208 ();
 sg13g2_fill_2 FILLER_55_242 ();
 sg13g2_fill_1 FILLER_55_259 ();
 sg13g2_fill_1 FILLER_55_277 ();
 sg13g2_decap_8 FILLER_55_290 ();
 sg13g2_decap_8 FILLER_55_297 ();
 sg13g2_decap_8 FILLER_55_304 ();
 sg13g2_decap_4 FILLER_55_311 ();
 sg13g2_fill_1 FILLER_55_331 ();
 sg13g2_fill_2 FILLER_55_344 ();
 sg13g2_fill_1 FILLER_55_346 ();
 sg13g2_fill_2 FILLER_56_77 ();
 sg13g2_fill_2 FILLER_56_92 ();
 sg13g2_fill_1 FILLER_56_94 ();
 sg13g2_decap_8 FILLER_56_131 ();
 sg13g2_decap_8 FILLER_56_138 ();
 sg13g2_decap_8 FILLER_56_145 ();
 sg13g2_decap_4 FILLER_56_152 ();
 sg13g2_decap_8 FILLER_56_204 ();
 sg13g2_fill_2 FILLER_56_211 ();
 sg13g2_decap_8 FILLER_56_217 ();
 sg13g2_decap_8 FILLER_56_228 ();
 sg13g2_decap_8 FILLER_56_235 ();
 sg13g2_decap_8 FILLER_56_246 ();
 sg13g2_decap_8 FILLER_56_253 ();
 sg13g2_decap_8 FILLER_56_260 ();
 sg13g2_fill_2 FILLER_56_267 ();
 sg13g2_fill_1 FILLER_56_269 ();
 sg13g2_decap_8 FILLER_56_280 ();
 sg13g2_decap_8 FILLER_56_287 ();
 sg13g2_decap_4 FILLER_56_294 ();
 sg13g2_fill_1 FILLER_56_298 ();
 sg13g2_fill_2 FILLER_56_308 ();
 sg13g2_fill_1 FILLER_56_314 ();
 sg13g2_fill_1 FILLER_56_343 ();
 sg13g2_fill_1 FILLER_56_399 ();
 sg13g2_fill_2 FILLER_57_48 ();
 sg13g2_fill_1 FILLER_57_50 ();
 sg13g2_fill_1 FILLER_57_64 ();
 sg13g2_fill_2 FILLER_57_70 ();
 sg13g2_fill_1 FILLER_57_82 ();
 sg13g2_decap_8 FILLER_57_121 ();
 sg13g2_decap_4 FILLER_57_128 ();
 sg13g2_decap_8 FILLER_57_148 ();
 sg13g2_decap_4 FILLER_57_155 ();
 sg13g2_fill_2 FILLER_57_159 ();
 sg13g2_decap_8 FILLER_57_165 ();
 sg13g2_decap_8 FILLER_57_172 ();
 sg13g2_fill_2 FILLER_57_179 ();
 sg13g2_decap_8 FILLER_57_192 ();
 sg13g2_decap_8 FILLER_57_199 ();
 sg13g2_decap_8 FILLER_57_206 ();
 sg13g2_decap_8 FILLER_57_213 ();
 sg13g2_decap_4 FILLER_57_220 ();
 sg13g2_decap_8 FILLER_57_239 ();
 sg13g2_decap_8 FILLER_57_246 ();
 sg13g2_decap_4 FILLER_57_253 ();
 sg13g2_fill_2 FILLER_57_257 ();
 sg13g2_fill_2 FILLER_57_273 ();
 sg13g2_fill_1 FILLER_57_275 ();
 sg13g2_decap_4 FILLER_57_284 ();
 sg13g2_fill_1 FILLER_57_288 ();
 sg13g2_fill_2 FILLER_57_330 ();
 sg13g2_fill_1 FILLER_57_332 ();
 sg13g2_fill_2 FILLER_57_380 ();
 sg13g2_decap_4 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_4 ();
 sg13g2_fill_1 FILLER_58_14 ();
 sg13g2_fill_2 FILLER_58_49 ();
 sg13g2_fill_2 FILLER_58_64 ();
 sg13g2_decap_8 FILLER_58_81 ();
 sg13g2_fill_2 FILLER_58_88 ();
 sg13g2_fill_1 FILLER_58_105 ();
 sg13g2_decap_8 FILLER_58_111 ();
 sg13g2_decap_8 FILLER_58_118 ();
 sg13g2_fill_2 FILLER_58_125 ();
 sg13g2_fill_2 FILLER_58_132 ();
 sg13g2_fill_1 FILLER_58_134 ();
 sg13g2_decap_4 FILLER_58_172 ();
 sg13g2_fill_1 FILLER_58_176 ();
 sg13g2_fill_2 FILLER_58_185 ();
 sg13g2_decap_8 FILLER_58_192 ();
 sg13g2_decap_8 FILLER_58_203 ();
 sg13g2_decap_4 FILLER_58_210 ();
 sg13g2_fill_2 FILLER_58_214 ();
 sg13g2_fill_2 FILLER_58_245 ();
 sg13g2_fill_1 FILLER_58_247 ();
 sg13g2_fill_2 FILLER_58_300 ();
 sg13g2_fill_2 FILLER_58_319 ();
 sg13g2_fill_1 FILLER_58_321 ();
 sg13g2_fill_2 FILLER_58_377 ();
 sg13g2_fill_2 FILLER_58_397 ();
 sg13g2_fill_1 FILLER_58_399 ();
 sg13g2_fill_2 FILLER_59_30 ();
 sg13g2_fill_2 FILLER_59_46 ();
 sg13g2_fill_1 FILLER_59_48 ();
 sg13g2_decap_8 FILLER_59_58 ();
 sg13g2_fill_2 FILLER_59_65 ();
 sg13g2_fill_1 FILLER_59_67 ();
 sg13g2_fill_2 FILLER_59_73 ();
 sg13g2_decap_8 FILLER_59_93 ();
 sg13g2_decap_4 FILLER_59_105 ();
 sg13g2_decap_4 FILLER_59_114 ();
 sg13g2_fill_1 FILLER_59_118 ();
 sg13g2_fill_1 FILLER_59_131 ();
 sg13g2_fill_1 FILLER_59_148 ();
 sg13g2_fill_2 FILLER_59_164 ();
 sg13g2_fill_1 FILLER_59_166 ();
 sg13g2_fill_2 FILLER_59_183 ();
 sg13g2_fill_1 FILLER_59_185 ();
 sg13g2_fill_2 FILLER_59_194 ();
 sg13g2_decap_8 FILLER_59_209 ();
 sg13g2_fill_2 FILLER_59_216 ();
 sg13g2_fill_1 FILLER_59_218 ();
 sg13g2_fill_2 FILLER_59_229 ();
 sg13g2_fill_1 FILLER_59_231 ();
 sg13g2_fill_1 FILLER_59_259 ();
 sg13g2_fill_2 FILLER_59_316 ();
 sg13g2_fill_2 FILLER_59_355 ();
 sg13g2_fill_1 FILLER_59_357 ();
 sg13g2_fill_1 FILLER_59_399 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_7 ();
 sg13g2_decap_4 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_120 ();
 sg13g2_decap_8 FILLER_60_127 ();
 sg13g2_fill_1 FILLER_60_134 ();
 sg13g2_decap_8 FILLER_60_140 ();
 sg13g2_fill_2 FILLER_60_147 ();
 sg13g2_fill_2 FILLER_60_168 ();
 sg13g2_decap_8 FILLER_60_217 ();
 sg13g2_decap_4 FILLER_60_224 ();
 sg13g2_decap_8 FILLER_60_237 ();
 sg13g2_decap_4 FILLER_60_244 ();
 sg13g2_fill_2 FILLER_60_248 ();
 sg13g2_decap_8 FILLER_60_269 ();
 sg13g2_fill_2 FILLER_60_276 ();
 sg13g2_fill_2 FILLER_60_295 ();
 sg13g2_fill_1 FILLER_60_297 ();
 sg13g2_fill_2 FILLER_60_351 ();
 sg13g2_decap_4 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_4 ();
 sg13g2_fill_2 FILLER_61_23 ();
 sg13g2_fill_1 FILLER_61_25 ();
 sg13g2_fill_1 FILLER_61_112 ();
 sg13g2_decap_8 FILLER_61_117 ();
 sg13g2_decap_8 FILLER_61_124 ();
 sg13g2_decap_4 FILLER_61_131 ();
 sg13g2_decap_4 FILLER_61_148 ();
 sg13g2_fill_1 FILLER_61_152 ();
 sg13g2_fill_1 FILLER_61_161 ();
 sg13g2_decap_8 FILLER_61_171 ();
 sg13g2_fill_1 FILLER_61_178 ();
 sg13g2_fill_2 FILLER_61_191 ();
 sg13g2_fill_1 FILLER_61_193 ();
 sg13g2_decap_8 FILLER_61_212 ();
 sg13g2_decap_8 FILLER_61_219 ();
 sg13g2_fill_2 FILLER_61_226 ();
 sg13g2_fill_1 FILLER_61_228 ();
 sg13g2_decap_8 FILLER_61_237 ();
 sg13g2_decap_8 FILLER_61_244 ();
 sg13g2_decap_8 FILLER_61_251 ();
 sg13g2_fill_2 FILLER_61_258 ();
 sg13g2_decap_4 FILLER_61_264 ();
 sg13g2_fill_2 FILLER_61_329 ();
 sg13g2_fill_1 FILLER_61_331 ();
 sg13g2_fill_1 FILLER_61_369 ();
 sg13g2_fill_1 FILLER_61_394 ();
 sg13g2_fill_1 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_40 ();
 sg13g2_fill_2 FILLER_62_78 ();
 sg13g2_fill_1 FILLER_62_80 ();
 sg13g2_fill_2 FILLER_62_104 ();
 sg13g2_fill_1 FILLER_62_106 ();
 sg13g2_fill_1 FILLER_62_127 ();
 sg13g2_decap_8 FILLER_62_143 ();
 sg13g2_decap_8 FILLER_62_150 ();
 sg13g2_fill_2 FILLER_62_157 ();
 sg13g2_fill_2 FILLER_62_163 ();
 sg13g2_fill_1 FILLER_62_165 ();
 sg13g2_decap_8 FILLER_62_170 ();
 sg13g2_decap_8 FILLER_62_177 ();
 sg13g2_decap_8 FILLER_62_184 ();
 sg13g2_decap_8 FILLER_62_191 ();
 sg13g2_decap_4 FILLER_62_198 ();
 sg13g2_decap_8 FILLER_62_206 ();
 sg13g2_decap_4 FILLER_62_213 ();
 sg13g2_fill_1 FILLER_62_225 ();
 sg13g2_decap_8 FILLER_62_244 ();
 sg13g2_decap_8 FILLER_62_251 ();
 sg13g2_fill_2 FILLER_62_258 ();
 sg13g2_fill_1 FILLER_62_260 ();
 sg13g2_fill_1 FILLER_62_279 ();
 sg13g2_fill_2 FILLER_62_285 ();
 sg13g2_fill_1 FILLER_62_287 ();
 sg13g2_fill_2 FILLER_62_301 ();
 sg13g2_fill_1 FILLER_62_311 ();
 sg13g2_fill_2 FILLER_62_370 ();
 sg13g2_fill_1 FILLER_62_372 ();
 sg13g2_fill_2 FILLER_62_386 ();
 sg13g2_decap_4 FILLER_63_27 ();
 sg13g2_fill_1 FILLER_63_66 ();
 sg13g2_fill_2 FILLER_63_95 ();
 sg13g2_fill_1 FILLER_63_97 ();
 sg13g2_fill_2 FILLER_63_125 ();
 sg13g2_fill_1 FILLER_63_127 ();
 sg13g2_fill_1 FILLER_63_151 ();
 sg13g2_fill_1 FILLER_63_156 ();
 sg13g2_fill_1 FILLER_63_162 ();
 sg13g2_fill_2 FILLER_63_168 ();
 sg13g2_decap_8 FILLER_63_178 ();
 sg13g2_fill_2 FILLER_63_185 ();
 sg13g2_decap_8 FILLER_63_191 ();
 sg13g2_decap_8 FILLER_63_198 ();
 sg13g2_fill_1 FILLER_63_205 ();
 sg13g2_fill_2 FILLER_63_228 ();
 sg13g2_fill_2 FILLER_63_262 ();
 sg13g2_fill_1 FILLER_63_264 ();
 sg13g2_fill_2 FILLER_63_273 ();
 sg13g2_fill_1 FILLER_63_275 ();
 sg13g2_fill_2 FILLER_63_301 ();
 sg13g2_fill_1 FILLER_63_303 ();
 sg13g2_fill_1 FILLER_63_342 ();
 sg13g2_fill_2 FILLER_63_348 ();
 sg13g2_fill_1 FILLER_63_350 ();
 sg13g2_fill_2 FILLER_63_379 ();
 sg13g2_fill_1 FILLER_63_381 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_4 FILLER_64_7 ();
 sg13g2_fill_1 FILLER_64_11 ();
 sg13g2_fill_2 FILLER_64_102 ();
 sg13g2_fill_2 FILLER_64_170 ();
 sg13g2_fill_2 FILLER_64_177 ();
 sg13g2_fill_1 FILLER_64_179 ();
 sg13g2_fill_2 FILLER_64_185 ();
 sg13g2_fill_1 FILLER_64_192 ();
 sg13g2_fill_1 FILLER_64_353 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_fill_2 FILLER_65_21 ();
 sg13g2_fill_1 FILLER_65_23 ();
 sg13g2_fill_2 FILLER_65_55 ();
 sg13g2_decap_8 FILLER_65_143 ();
 sg13g2_fill_2 FILLER_65_150 ();
 sg13g2_fill_2 FILLER_65_167 ();
 sg13g2_fill_1 FILLER_65_205 ();
 sg13g2_fill_1 FILLER_65_228 ();
 sg13g2_fill_2 FILLER_65_264 ();
 sg13g2_fill_2 FILLER_65_301 ();
 sg13g2_fill_1 FILLER_65_307 ();
 sg13g2_fill_2 FILLER_65_313 ();
 sg13g2_fill_1 FILLER_65_315 ();
 sg13g2_fill_2 FILLER_65_321 ();
 sg13g2_fill_2 FILLER_65_407 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_4 FILLER_66_21 ();
 sg13g2_fill_1 FILLER_66_25 ();
 sg13g2_fill_2 FILLER_66_77 ();
 sg13g2_fill_1 FILLER_66_120 ();
 sg13g2_fill_1 FILLER_66_127 ();
 sg13g2_fill_1 FILLER_66_160 ();
 sg13g2_fill_2 FILLER_66_174 ();
 sg13g2_fill_1 FILLER_66_176 ();
 sg13g2_fill_2 FILLER_66_193 ();
 sg13g2_fill_1 FILLER_66_195 ();
 sg13g2_fill_2 FILLER_66_206 ();
 sg13g2_fill_1 FILLER_66_208 ();
 sg13g2_fill_1 FILLER_66_223 ();
 sg13g2_fill_2 FILLER_66_239 ();
 sg13g2_fill_2 FILLER_66_268 ();
 sg13g2_fill_1 FILLER_66_270 ();
 sg13g2_fill_2 FILLER_66_292 ();
 sg13g2_fill_2 FILLER_66_304 ();
 sg13g2_fill_1 FILLER_66_306 ();
 sg13g2_fill_2 FILLER_66_312 ();
 sg13g2_fill_1 FILLER_66_314 ();
 sg13g2_fill_2 FILLER_66_379 ();
 sg13g2_fill_1 FILLER_66_381 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_fill_1 FILLER_67_21 ();
 sg13g2_fill_2 FILLER_67_58 ();
 sg13g2_fill_1 FILLER_67_60 ();
 sg13g2_fill_2 FILLER_67_76 ();
 sg13g2_fill_2 FILLER_67_87 ();
 sg13g2_fill_2 FILLER_67_102 ();
 sg13g2_fill_2 FILLER_67_140 ();
 sg13g2_decap_4 FILLER_67_169 ();
 sg13g2_decap_4 FILLER_67_177 ();
 sg13g2_fill_2 FILLER_67_181 ();
 sg13g2_fill_2 FILLER_67_210 ();
 sg13g2_fill_1 FILLER_67_223 ();
 sg13g2_fill_2 FILLER_67_235 ();
 sg13g2_fill_2 FILLER_67_249 ();
 sg13g2_fill_1 FILLER_67_251 ();
 sg13g2_fill_2 FILLER_67_274 ();
 sg13g2_fill_2 FILLER_67_294 ();
 sg13g2_fill_2 FILLER_67_309 ();
 sg13g2_fill_1 FILLER_67_344 ();
 sg13g2_fill_2 FILLER_67_350 ();
 sg13g2_fill_1 FILLER_67_395 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_fill_1 FILLER_68_21 ();
 sg13g2_fill_1 FILLER_68_49 ();
 sg13g2_fill_2 FILLER_68_59 ();
 sg13g2_fill_1 FILLER_68_61 ();
 sg13g2_fill_2 FILLER_68_113 ();
 sg13g2_fill_1 FILLER_68_115 ();
 sg13g2_fill_1 FILLER_68_121 ();
 sg13g2_fill_2 FILLER_68_140 ();
 sg13g2_fill_1 FILLER_68_155 ();
 sg13g2_decap_8 FILLER_68_177 ();
 sg13g2_fill_2 FILLER_68_184 ();
 sg13g2_fill_1 FILLER_68_186 ();
 sg13g2_decap_4 FILLER_68_197 ();
 sg13g2_fill_1 FILLER_68_250 ();
 sg13g2_fill_2 FILLER_68_265 ();
 sg13g2_fill_1 FILLER_68_267 ();
 sg13g2_fill_2 FILLER_68_281 ();
 sg13g2_fill_2 FILLER_68_309 ();
 sg13g2_fill_1 FILLER_68_311 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_fill_2 FILLER_69_14 ();
 sg13g2_fill_1 FILLER_69_49 ();
 sg13g2_fill_1 FILLER_69_74 ();
 sg13g2_fill_1 FILLER_69_135 ();
 sg13g2_fill_1 FILLER_69_149 ();
 sg13g2_fill_2 FILLER_69_169 ();
 sg13g2_fill_2 FILLER_69_216 ();
 sg13g2_fill_1 FILLER_69_218 ();
 sg13g2_fill_2 FILLER_69_227 ();
 sg13g2_fill_1 FILLER_69_239 ();
 sg13g2_fill_2 FILLER_69_378 ();
 sg13g2_fill_1 FILLER_69_380 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_4 FILLER_70_14 ();
 sg13g2_fill_1 FILLER_70_97 ();
 sg13g2_fill_2 FILLER_70_116 ();
 sg13g2_fill_1 FILLER_70_196 ();
 sg13g2_fill_2 FILLER_70_214 ();
 sg13g2_fill_2 FILLER_70_242 ();
 sg13g2_fill_2 FILLER_70_258 ();
 sg13g2_fill_1 FILLER_70_260 ();
 sg13g2_fill_2 FILLER_70_284 ();
 sg13g2_fill_1 FILLER_70_297 ();
 sg13g2_fill_2 FILLER_70_333 ();
 sg13g2_fill_1 FILLER_70_335 ();
 sg13g2_fill_2 FILLER_70_369 ();
 sg13g2_fill_1 FILLER_70_371 ();
 sg13g2_fill_2 FILLER_70_398 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_fill_2 FILLER_71_82 ();
 sg13g2_fill_1 FILLER_71_84 ();
 sg13g2_fill_2 FILLER_71_127 ();
 sg13g2_fill_1 FILLER_71_220 ();
 sg13g2_fill_1 FILLER_71_239 ();
 sg13g2_fill_2 FILLER_71_273 ();
 sg13g2_fill_1 FILLER_71_288 ();
 sg13g2_fill_1 FILLER_71_322 ();
 sg13g2_fill_1 FILLER_71_338 ();
 sg13g2_fill_2 FILLER_71_367 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_fill_2 FILLER_72_14 ();
 sg13g2_fill_1 FILLER_72_70 ();
 sg13g2_fill_1 FILLER_72_76 ();
 sg13g2_fill_1 FILLER_72_90 ();
 sg13g2_fill_1 FILLER_72_104 ();
 sg13g2_fill_2 FILLER_72_139 ();
 sg13g2_fill_1 FILLER_72_141 ();
 sg13g2_fill_1 FILLER_72_160 ();
 sg13g2_fill_2 FILLER_72_243 ();
 sg13g2_fill_1 FILLER_72_245 ();
 sg13g2_fill_2 FILLER_72_255 ();
 sg13g2_fill_1 FILLER_72_257 ();
 sg13g2_fill_2 FILLER_72_304 ();
 sg13g2_fill_1 FILLER_72_306 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_decap_4 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_4 ();
 sg13g2_fill_2 FILLER_73_76 ();
 sg13g2_fill_1 FILLER_73_132 ();
 sg13g2_fill_2 FILLER_73_146 ();
 sg13g2_fill_2 FILLER_73_194 ();
 sg13g2_fill_1 FILLER_73_196 ();
 sg13g2_fill_1 FILLER_73_219 ();
 sg13g2_fill_1 FILLER_73_327 ();
 sg13g2_fill_1 FILLER_73_341 ();
 sg13g2_fill_2 FILLER_73_360 ();
 sg13g2_fill_1 FILLER_73_362 ();
 sg13g2_fill_1 FILLER_73_408 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_7 ();
 sg13g2_fill_2 FILLER_74_82 ();
 sg13g2_fill_2 FILLER_74_107 ();
 sg13g2_fill_1 FILLER_74_109 ();
 sg13g2_fill_2 FILLER_74_194 ();
 sg13g2_fill_1 FILLER_74_196 ();
 sg13g2_fill_2 FILLER_74_215 ();
 sg13g2_fill_2 FILLER_74_221 ();
 sg13g2_fill_1 FILLER_74_261 ();
 sg13g2_fill_1 FILLER_74_329 ();
 sg13g2_fill_1 FILLER_74_335 ();
 sg13g2_fill_2 FILLER_74_364 ();
 sg13g2_fill_1 FILLER_74_366 ();
 sg13g2_fill_1 FILLER_74_389 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_4 FILLER_75_7 ();
 sg13g2_fill_2 FILLER_75_11 ();
 sg13g2_fill_1 FILLER_75_177 ();
 sg13g2_fill_2 FILLER_75_196 ();
 sg13g2_fill_1 FILLER_75_198 ();
 sg13g2_fill_2 FILLER_75_203 ();
 sg13g2_fill_1 FILLER_75_205 ();
 sg13g2_fill_2 FILLER_75_211 ();
 sg13g2_fill_2 FILLER_75_217 ();
 sg13g2_fill_1 FILLER_75_232 ();
 sg13g2_fill_1 FILLER_75_256 ();
 sg13g2_fill_1 FILLER_75_285 ();
 sg13g2_fill_2 FILLER_75_331 ();
 sg13g2_fill_1 FILLER_75_361 ();
 sg13g2_fill_1 FILLER_75_390 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_4 FILLER_76_14 ();
 sg13g2_fill_2 FILLER_76_18 ();
 sg13g2_fill_1 FILLER_76_96 ();
 sg13g2_fill_1 FILLER_76_156 ();
 sg13g2_fill_1 FILLER_76_202 ();
 sg13g2_fill_2 FILLER_76_248 ();
 sg13g2_fill_1 FILLER_76_250 ();
 sg13g2_fill_2 FILLER_76_314 ();
 sg13g2_fill_1 FILLER_76_316 ();
 sg13g2_fill_1 FILLER_76_330 ();
 sg13g2_fill_2 FILLER_76_355 ();
 sg13g2_fill_2 FILLER_76_379 ();
 sg13g2_fill_1 FILLER_76_381 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_fill_2 FILLER_77_21 ();
 sg13g2_fill_1 FILLER_77_23 ();
 sg13g2_fill_2 FILLER_77_130 ();
 sg13g2_fill_1 FILLER_77_132 ();
 sg13g2_fill_1 FILLER_77_146 ();
 sg13g2_fill_1 FILLER_77_208 ();
 sg13g2_fill_2 FILLER_77_214 ();
 sg13g2_fill_1 FILLER_77_216 ();
 sg13g2_fill_2 FILLER_77_255 ();
 sg13g2_fill_1 FILLER_77_293 ();
 sg13g2_fill_1 FILLER_77_332 ();
 sg13g2_fill_2 FILLER_77_397 ();
 sg13g2_fill_1 FILLER_77_399 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_fill_2 FILLER_78_28 ();
 sg13g2_fill_2 FILLER_78_191 ();
 sg13g2_fill_1 FILLER_78_193 ();
 sg13g2_fill_1 FILLER_78_277 ();
 sg13g2_fill_1 FILLER_78_287 ();
 sg13g2_fill_2 FILLER_78_398 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_4 FILLER_79_21 ();
 sg13g2_fill_2 FILLER_79_25 ();
 sg13g2_fill_2 FILLER_79_102 ();
 sg13g2_fill_1 FILLER_79_104 ();
 sg13g2_fill_2 FILLER_79_110 ();
 sg13g2_fill_1 FILLER_79_215 ();
 sg13g2_fill_1 FILLER_79_225 ();
 sg13g2_fill_2 FILLER_79_266 ();
 sg13g2_fill_1 FILLER_79_349 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_fill_2 FILLER_80_14 ();
 sg13g2_fill_1 FILLER_80_76 ();
 sg13g2_fill_2 FILLER_80_100 ();
 sg13g2_fill_1 FILLER_80_102 ();
 sg13g2_fill_2 FILLER_80_131 ();
 sg13g2_fill_1 FILLER_80_133 ();
 sg13g2_fill_2 FILLER_80_180 ();
 sg13g2_fill_1 FILLER_80_202 ();
 sg13g2_fill_1 FILLER_80_211 ();
 sg13g2_fill_1 FILLER_80_245 ();
 sg13g2_fill_1 FILLER_80_256 ();
 sg13g2_fill_1 FILLER_80_263 ();
 sg13g2_fill_2 FILLER_80_297 ();
 sg13g2_fill_2 FILLER_80_312 ();
 sg13g2_fill_1 FILLER_80_314 ();
 sg13g2_fill_1 FILLER_80_324 ();
 sg13g2_fill_1 FILLER_80_386 ();
 assign uio_oe[0] = net26;
 assign uio_oe[1] = net12;
 assign uio_oe[2] = net13;
 assign uio_oe[3] = net14;
 assign uio_oe[4] = net15;
 assign uio_oe[5] = net16;
 assign uio_oe[6] = net17;
 assign uio_oe[7] = net18;
 assign uio_out[1] = net19;
 assign uio_out[2] = net20;
 assign uio_out[3] = net21;
 assign uio_out[4] = net22;
 assign uio_out[5] = net23;
 assign uio_out[6] = net24;
 assign uio_out[7] = net25;
endmodule
