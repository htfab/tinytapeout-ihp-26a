module tt_um_rejunity_vga_logo (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire clknet_0_clk;
 wire \bayer_j[0] ;
 wire \bayer_j[1] ;
 wire \cos_addr[0] ;
 wire \cos_addr[1] ;
 wire \cos_addr[2] ;
 wire \cos_addr[3] ;
 wire \cos_addr[4] ;
 wire \cos_addr[5] ;
 wire \cos_addr[6] ;
 wire \cos_x_acc[0] ;
 wire \cos_x_acc[10] ;
 wire \cos_x_acc[11] ;
 wire \cos_x_acc[12] ;
 wire \cos_x_acc[13] ;
 wire \cos_x_acc[14] ;
 wire \cos_x_acc[15] ;
 wire \cos_x_acc[16] ;
 wire \cos_x_acc[17] ;
 wire \cos_x_acc[18] ;
 wire \cos_x_acc[19] ;
 wire \cos_x_acc[1] ;
 wire \cos_x_acc[20] ;
 wire \cos_x_acc[21] ;
 wire \cos_x_acc[22] ;
 wire \cos_x_acc[23] ;
 wire \cos_x_acc[24] ;
 wire \cos_x_acc[25] ;
 wire \cos_x_acc[26] ;
 wire \cos_x_acc[2] ;
 wire \cos_x_acc[3] ;
 wire \cos_x_acc[4] ;
 wire \cos_x_acc[5] ;
 wire \cos_x_acc[6] ;
 wire \cos_x_acc[7] ;
 wire \cos_x_acc[8] ;
 wire \cos_x_acc[9] ;
 wire \cos_y_acc[0] ;
 wire \cos_y_acc[10] ;
 wire \cos_y_acc[11] ;
 wire \cos_y_acc[12] ;
 wire \cos_y_acc[13] ;
 wire \cos_y_acc[14] ;
 wire \cos_y_acc[15] ;
 wire \cos_y_acc[16] ;
 wire \cos_y_acc[17] ;
 wire \cos_y_acc[18] ;
 wire \cos_y_acc[19] ;
 wire \cos_y_acc[1] ;
 wire \cos_y_acc[20] ;
 wire \cos_y_acc[21] ;
 wire \cos_y_acc[22] ;
 wire \cos_y_acc[23] ;
 wire \cos_y_acc[24] ;
 wire \cos_y_acc[25] ;
 wire \cos_y_acc[26] ;
 wire \cos_y_acc[2] ;
 wire \cos_y_acc[3] ;
 wire \cos_y_acc[4] ;
 wire \cos_y_acc[5] ;
 wire \cos_y_acc[6] ;
 wire \cos_y_acc[7] ;
 wire \cos_y_acc[8] ;
 wire \cos_y_acc[9] ;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire \sin_x_acc[0] ;
 wire \sin_x_acc[10] ;
 wire \sin_x_acc[11] ;
 wire \sin_x_acc[12] ;
 wire \sin_x_acc[13] ;
 wire \sin_x_acc[14] ;
 wire \sin_x_acc[15] ;
 wire \sin_x_acc[16] ;
 wire \sin_x_acc[17] ;
 wire \sin_x_acc[18] ;
 wire \sin_x_acc[19] ;
 wire \sin_x_acc[1] ;
 wire \sin_x_acc[20] ;
 wire \sin_x_acc[21] ;
 wire \sin_x_acc[22] ;
 wire \sin_x_acc[23] ;
 wire \sin_x_acc[24] ;
 wire \sin_x_acc[25] ;
 wire \sin_x_acc[26] ;
 wire \sin_x_acc[2] ;
 wire \sin_x_acc[3] ;
 wire \sin_x_acc[4] ;
 wire \sin_x_acc[5] ;
 wire \sin_x_acc[6] ;
 wire \sin_x_acc[7] ;
 wire \sin_x_acc[8] ;
 wire \sin_x_acc[9] ;
 wire \sin_y_acc[0] ;
 wire \sin_y_acc[10] ;
 wire \sin_y_acc[11] ;
 wire \sin_y_acc[12] ;
 wire \sin_y_acc[13] ;
 wire \sin_y_acc[14] ;
 wire \sin_y_acc[15] ;
 wire \sin_y_acc[16] ;
 wire \sin_y_acc[17] ;
 wire \sin_y_acc[18] ;
 wire \sin_y_acc[19] ;
 wire \sin_y_acc[1] ;
 wire \sin_y_acc[20] ;
 wire \sin_y_acc[21] ;
 wire \sin_y_acc[22] ;
 wire \sin_y_acc[23] ;
 wire \sin_y_acc[24] ;
 wire \sin_y_acc[25] ;
 wire \sin_y_acc[26] ;
 wire \sin_y_acc[2] ;
 wire \sin_y_acc[3] ;
 wire \sin_y_acc[4] ;
 wire \sin_y_acc[5] ;
 wire \sin_y_acc[6] ;
 wire \sin_y_acc[7] ;
 wire \sin_y_acc[8] ;
 wire \sin_y_acc[9] ;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire \y_prv[0] ;
 wire \y_prv[1] ;
 wire \y_prv[2] ;
 wire \y_prv[3] ;
 wire \y_prv[4] ;
 wire \y_prv[5] ;
 wire \y_prv[6] ;
 wire \y_prv[7] ;
 wire \y_prv[8] ;
 wire \y_prv[9] ;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net1;
 wire net2;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;

 sg13g2_inv_1 _2040_ (.Y(_1193_),
    .A(\cos_y_acc[21] ));
 sg13g2_inv_1 _2041_ (.Y(_1194_),
    .A(\cos_y_acc[19] ));
 sg13g2_inv_1 _2042_ (.Y(_1195_),
    .A(\cos_y_acc[17] ));
 sg13g2_inv_1 _2043_ (.Y(_1196_),
    .A(\cos_y_acc[16] ));
 sg13g2_inv_2 _2044_ (.Y(_1197_),
    .A(net422));
 sg13g2_inv_1 _2045_ (.Y(_1198_),
    .A(net426));
 sg13g2_inv_1 _2046_ (.Y(_1199_),
    .A(net425));
 sg13g2_inv_1 _2047_ (.Y(_1200_),
    .A(net432));
 sg13g2_inv_1 _2048_ (.Y(_1201_),
    .A(net443));
 sg13g2_inv_1 _2049_ (.Y(_1202_),
    .A(net447));
 sg13g2_inv_1 _2050_ (.Y(_1203_),
    .A(net434));
 sg13g2_inv_2 _2051_ (.Y(_1204_),
    .A(net410));
 sg13g2_inv_2 _2052_ (.Y(_1205_),
    .A(net386));
 sg13g2_inv_2 _2053_ (.Y(_1206_),
    .A(net399));
 sg13g2_inv_1 _2054_ (.Y(_1207_),
    .A(\sin_y_acc[17] ));
 sg13g2_inv_2 _2055_ (.Y(_1208_),
    .A(net339));
 sg13g2_inv_1 _2056_ (.Y(_1209_),
    .A(net446));
 sg13g2_inv_1 _2057_ (.Y(_1210_),
    .A(net373));
 sg13g2_inv_2 _2058_ (.Y(_1211_),
    .A(net381));
 sg13g2_inv_1 _2059_ (.Y(_1212_),
    .A(net423));
 sg13g2_inv_1 _2060_ (.Y(_1213_),
    .A(\sin_x_acc[3] ));
 sg13g2_inv_2 _2061_ (.Y(_1214_),
    .A(net481));
 sg13g2_inv_2 _2062_ (.Y(_1215_),
    .A(net343));
 sg13g2_inv_1 _2063_ (.Y(_1216_),
    .A(\bayer_j[1] ));
 sg13g2_inv_1 _2064_ (.Y(_1217_),
    .A(net273));
 sg13g2_inv_2 _2065_ (.Y(_1218_),
    .A(net436));
 sg13g2_inv_2 _2066_ (.Y(_1219_),
    .A(net464));
 sg13g2_inv_2 _2067_ (.Y(_1220_),
    .A(net334));
 sg13g2_inv_1 _2068_ (.Y(_1221_),
    .A(\cos_x_acc[24] ));
 sg13g2_inv_1 _2069_ (.Y(_1222_),
    .A(\sin_x_acc[25] ));
 sg13g2_inv_1 _2070_ (.Y(_1223_),
    .A(\sin_x_acc[24] ));
 sg13g2_inv_1 _2071_ (.Y(_1224_),
    .A(\sin_x_acc[4] ));
 sg13g2_inv_1 _2072_ (.Y(_1225_),
    .A(\sin_x_acc[7] ));
 sg13g2_inv_1 _2073_ (.Y(_1226_),
    .A(\sin_x_acc[10] ));
 sg13g2_inv_2 _2074_ (.Y(_1227_),
    .A(net474));
 sg13g2_inv_2 _2075_ (.Y(_1228_),
    .A(\cos_x_acc[4] ));
 sg13g2_inv_1 _2076_ (.Y(_1229_),
    .A(\cos_x_acc[9] ));
 sg13g2_inv_1 _2077_ (.Y(_1230_),
    .A(net448));
 sg13g2_inv_2 _2078_ (.Y(_1231_),
    .A(net492));
 sg13g2_inv_1 _2079_ (.Y(_1232_),
    .A(net462));
 sg13g2_inv_1 _2080_ (.Y(_1233_),
    .A(net375));
 sg13g2_inv_1 _2081_ (.Y(_1234_),
    .A(net469));
 sg13g2_inv_2 _2082_ (.Y(_1235_),
    .A(net411));
 sg13g2_inv_1 _2083_ (.Y(_1236_),
    .A(\cos_x_acc[22] ));
 sg13g2_inv_1 _2084_ (.Y(_1237_),
    .A(\hvsync_gen.vpos[2] ));
 sg13g2_inv_2 _2085_ (.Y(_1238_),
    .A(net297));
 sg13g2_inv_1 _2086_ (.Y(_1239_),
    .A(net322));
 sg13g2_inv_2 _2087_ (.Y(_1240_),
    .A(net285));
 sg13g2_inv_1 _2088_ (.Y(_1241_),
    .A(\hvsync_gen.vpos[8] ));
 sg13g2_inv_1 _2089_ (.Y(_1242_),
    .A(\hvsync_gen.hpos[5] ));
 sg13g2_inv_1 _2090_ (.Y(_1243_),
    .A(\y_prv[0] ));
 sg13g2_inv_1 _2091_ (.Y(_1244_),
    .A(\y_prv[1] ));
 sg13g2_inv_1 _2092_ (.Y(_1245_),
    .A(\y_prv[3] ));
 sg13g2_inv_1 _2093_ (.Y(_1246_),
    .A(net276));
 sg13g2_inv_1 _2094_ (.Y(_1247_),
    .A(\y_prv[8] ));
 sg13g2_inv_1 _2095_ (.Y(_1248_),
    .A(net254));
 sg13g2_nand2b_1 _2096_ (.Y(_1249_),
    .B(\cos_x_acc[18] ),
    .A_N(\sin_y_acc[18] ));
 sg13g2_xnor2_1 _2097_ (.Y(_1250_),
    .A(\sin_y_acc[18] ),
    .B(\cos_x_acc[18] ));
 sg13g2_nor2b_1 _2098_ (.A(\sin_y_acc[15] ),
    .B_N(\cos_x_acc[15] ),
    .Y(_1251_));
 sg13g2_nand2b_1 _2099_ (.Y(_1252_),
    .B(\sin_y_acc[15] ),
    .A_N(\cos_x_acc[15] ));
 sg13g2_nor2b_1 _2100_ (.A(_1251_),
    .B_N(_1252_),
    .Y(_1253_));
 sg13g2_nor2b_1 _2101_ (.A(\sin_y_acc[14] ),
    .B_N(\cos_x_acc[14] ),
    .Y(_1254_));
 sg13g2_xnor2_1 _2102_ (.Y(_1255_),
    .A(\sin_y_acc[14] ),
    .B(\cos_x_acc[14] ));
 sg13g2_and2_1 _2103_ (.A(_1253_),
    .B(_1255_),
    .X(_1256_));
 sg13g2_nor2b_1 _2104_ (.A(\sin_y_acc[12] ),
    .B_N(\cos_x_acc[12] ),
    .Y(_1257_));
 sg13g2_a21oi_1 _2105_ (.A1(_1209_),
    .A2(\cos_x_acc[13] ),
    .Y(_1258_),
    .B1(_1257_));
 sg13g2_a21oi_1 _2106_ (.A1(\sin_y_acc[13] ),
    .A2(_1232_),
    .Y(_1259_),
    .B1(_1258_));
 sg13g2_inv_1 _2107_ (.Y(_1260_),
    .A(_1259_));
 sg13g2_a221oi_1 _2108_ (.B2(_1259_),
    .C1(_1251_),
    .B1(_1256_),
    .A1(_1252_),
    .Y(_1261_),
    .A2(_1254_));
 sg13g2_xor2_1 _2109_ (.B(\cos_x_acc[12] ),
    .A(\sin_y_acc[12] ),
    .X(_1262_));
 sg13g2_xnor2_1 _2110_ (.Y(_1263_),
    .A(\sin_y_acc[13] ),
    .B(\cos_x_acc[13] ));
 sg13g2_nor2b_1 _2111_ (.A(_1262_),
    .B_N(_1263_),
    .Y(_1264_));
 sg13g2_nand2b_1 _2112_ (.Y(_1265_),
    .B(_1263_),
    .A_N(_1262_));
 sg13g2_nand2_1 _2113_ (.Y(_1266_),
    .A(_1256_),
    .B(_1264_));
 sg13g2_nor2b_1 _2114_ (.A(\sin_y_acc[7] ),
    .B_N(\cos_x_acc[7] ),
    .Y(_1267_));
 sg13g2_nand2b_1 _2115_ (.Y(_1268_),
    .B(\cos_x_acc[6] ),
    .A_N(\sin_y_acc[6] ));
 sg13g2_nor2b_1 _2116_ (.A(\cos_x_acc[6] ),
    .B_N(\sin_y_acc[6] ),
    .Y(_1269_));
 sg13g2_xnor2_1 _2117_ (.Y(_1270_),
    .A(\sin_y_acc[6] ),
    .B(\cos_x_acc[6] ));
 sg13g2_nor2b_1 _2118_ (.A(\sin_y_acc[3] ),
    .B_N(\cos_x_acc[3] ),
    .Y(_1271_));
 sg13g2_nand2_1 _2119_ (.Y(_1272_),
    .A(_1212_),
    .B(\cos_x_acc[2] ));
 sg13g2_nor2b_1 _2120_ (.A(\sin_y_acc[1] ),
    .B_N(\cos_x_acc[1] ),
    .Y(_1273_));
 sg13g2_nand2b_2 _2121_ (.Y(_1274_),
    .B(\sin_y_acc[0] ),
    .A_N(\cos_x_acc[0] ));
 sg13g2_xnor2_1 _2122_ (.Y(_1275_),
    .A(\sin_y_acc[1] ),
    .B(\cos_x_acc[1] ));
 sg13g2_a21oi_1 _2123_ (.A1(_1274_),
    .A2(_1275_),
    .Y(_1276_),
    .B1(_1273_));
 sg13g2_nor2_1 _2124_ (.A(_1212_),
    .B(\cos_x_acc[2] ),
    .Y(_1277_));
 sg13g2_xnor2_1 _2125_ (.Y(_1278_),
    .A(\sin_y_acc[2] ),
    .B(\cos_x_acc[2] ));
 sg13g2_o21ai_1 _2126_ (.B1(_1272_),
    .Y(_1279_),
    .A1(_1276_),
    .A2(_1277_));
 sg13g2_xnor2_1 _2127_ (.Y(_1280_),
    .A(\sin_y_acc[3] ),
    .B(\cos_x_acc[3] ));
 sg13g2_a21o_2 _2128_ (.A2(_1280_),
    .A1(_1279_),
    .B1(_1271_),
    .X(_1281_));
 sg13g2_nor2_1 _2129_ (.A(\sin_y_acc[4] ),
    .B(_1228_),
    .Y(_1282_));
 sg13g2_xnor2_1 _2130_ (.Y(_1283_),
    .A(\sin_y_acc[4] ),
    .B(\cos_x_acc[4] ));
 sg13g2_nor2b_1 _2131_ (.A(\sin_y_acc[5] ),
    .B_N(\cos_x_acc[5] ),
    .Y(_1284_));
 sg13g2_nand2b_1 _2132_ (.Y(_1285_),
    .B(\sin_y_acc[5] ),
    .A_N(\cos_x_acc[5] ));
 sg13g2_nor2b_1 _2133_ (.A(_1284_),
    .B_N(_1285_),
    .Y(_1286_));
 sg13g2_and2_1 _2134_ (.A(_1283_),
    .B(_1286_),
    .X(_1287_));
 sg13g2_a221oi_1 _2135_ (.B2(_1281_),
    .C1(_1284_),
    .B1(_1287_),
    .A1(_1282_),
    .Y(_1288_),
    .A2(_1285_));
 sg13g2_o21ai_1 _2136_ (.B1(_1268_),
    .Y(_1289_),
    .A1(_1269_),
    .A2(_1288_));
 sg13g2_xnor2_1 _2137_ (.Y(_1290_),
    .A(\sin_y_acc[7] ),
    .B(\cos_x_acc[7] ));
 sg13g2_a21o_2 _2138_ (.A2(_1290_),
    .A1(_1289_),
    .B1(_1267_),
    .X(_1291_));
 sg13g2_nor2_1 _2139_ (.A(\sin_y_acc[11] ),
    .B(_1231_),
    .Y(_1292_));
 sg13g2_nand2_1 _2140_ (.Y(_1293_),
    .A(\sin_y_acc[11] ),
    .B(_1231_));
 sg13g2_nor2b_1 _2141_ (.A(_1292_),
    .B_N(_1293_),
    .Y(_1294_));
 sg13g2_nor2_1 _2142_ (.A(\sin_y_acc[10] ),
    .B(_1230_),
    .Y(_1295_));
 sg13g2_xnor2_1 _2143_ (.Y(_1296_),
    .A(\sin_y_acc[10] ),
    .B(\cos_x_acc[10] ));
 sg13g2_and2_1 _2144_ (.A(_1294_),
    .B(_1296_),
    .X(_1297_));
 sg13g2_nor2b_1 _2145_ (.A(\sin_y_acc[8] ),
    .B_N(\cos_x_acc[8] ),
    .Y(_1298_));
 sg13g2_xnor2_1 _2146_ (.Y(_1299_),
    .A(\sin_y_acc[8] ),
    .B(\cos_x_acc[8] ));
 sg13g2_xnor2_1 _2147_ (.Y(_1300_),
    .A(\sin_y_acc[9] ),
    .B(\cos_x_acc[9] ));
 sg13g2_and2_1 _2148_ (.A(_1299_),
    .B(_1300_),
    .X(_1301_));
 sg13g2_and2_1 _2149_ (.A(_1297_),
    .B(_1301_),
    .X(_1302_));
 sg13g2_nand2_1 _2150_ (.Y(_1303_),
    .A(_1291_),
    .B(_1302_));
 sg13g2_a21oi_1 _2151_ (.A1(_1211_),
    .A2(\cos_x_acc[9] ),
    .Y(_1304_),
    .B1(_1298_));
 sg13g2_a21oi_1 _2152_ (.A1(\sin_y_acc[9] ),
    .A2(_1229_),
    .Y(_1305_),
    .B1(_1304_));
 sg13g2_a221oi_1 _2153_ (.B2(_1305_),
    .C1(_1292_),
    .B1(_1297_),
    .A1(_1293_),
    .Y(_1306_),
    .A2(_1295_));
 sg13g2_inv_1 _2154_ (.Y(_1307_),
    .A(_1306_));
 sg13g2_a21oi_2 _2155_ (.B1(_1307_),
    .Y(_1308_),
    .A2(_1302_),
    .A1(_1291_));
 sg13g2_and2_1 _2156_ (.A(_1261_),
    .B(_1306_),
    .X(_1309_));
 sg13g2_o21ai_1 _2157_ (.B1(_1261_),
    .Y(_1310_),
    .A1(_1266_),
    .A2(_1308_));
 sg13g2_nor2b_1 _2158_ (.A(\sin_y_acc[16] ),
    .B_N(\cos_x_acc[16] ),
    .Y(_1311_));
 sg13g2_xnor2_1 _2159_ (.Y(_1312_),
    .A(\sin_y_acc[16] ),
    .B(\cos_x_acc[16] ));
 sg13g2_xnor2_1 _2160_ (.Y(_1313_),
    .A(\sin_y_acc[17] ),
    .B(\cos_x_acc[17] ));
 sg13g2_nand2_1 _2161_ (.Y(_1314_),
    .A(_1312_),
    .B(_1313_));
 sg13g2_a221oi_1 _2162_ (.B2(_1309_),
    .C1(_1314_),
    .B1(_1303_),
    .A1(_1261_),
    .Y(_1315_),
    .A2(_1266_));
 sg13g2_o21ai_1 _2163_ (.B1(_1311_),
    .Y(_1316_),
    .A1(_1207_),
    .A2(\cos_x_acc[17] ));
 sg13g2_o21ai_1 _2164_ (.B1(_1316_),
    .Y(_1317_),
    .A1(\sin_y_acc[17] ),
    .A2(_1233_));
 sg13g2_nor2_1 _2165_ (.A(_1315_),
    .B(_1317_),
    .Y(_1318_));
 sg13g2_o21ai_1 _2166_ (.B1(_1250_),
    .Y(_1319_),
    .A1(_1315_),
    .A2(_1317_));
 sg13g2_nand2b_1 _2167_ (.Y(_1320_),
    .B(\cos_x_acc[19] ),
    .A_N(\sin_y_acc[19] ));
 sg13g2_and2_1 _2168_ (.A(_1249_),
    .B(_1320_),
    .X(_1321_));
 sg13g2_a22oi_1 _2169_ (.Y(_1322_),
    .B1(_1319_),
    .B2(_1321_),
    .A2(_1235_),
    .A1(\sin_y_acc[19] ));
 sg13g2_nor2b_1 _2170_ (.A(\sin_y_acc[21] ),
    .B_N(\cos_x_acc[21] ),
    .Y(_1323_));
 sg13g2_nand2b_1 _2171_ (.Y(_1324_),
    .B(\sin_y_acc[21] ),
    .A_N(\cos_x_acc[21] ));
 sg13g2_nor2b_2 _2172_ (.A(_1323_),
    .B_N(_1324_),
    .Y(_1325_));
 sg13g2_nor2b_1 _2173_ (.A(\sin_y_acc[20] ),
    .B_N(\cos_x_acc[20] ),
    .Y(_1326_));
 sg13g2_xnor2_1 _2174_ (.Y(_1327_),
    .A(\sin_y_acc[20] ),
    .B(\cos_x_acc[20] ));
 sg13g2_nand2_1 _2175_ (.Y(_1328_),
    .A(_1325_),
    .B(_1327_));
 sg13g2_a221oi_1 _2176_ (.B2(_1321_),
    .C1(_1328_),
    .B1(_1319_),
    .A1(\sin_y_acc[19] ),
    .Y(_1329_),
    .A2(_1235_));
 sg13g2_a21o_1 _2177_ (.A2(_1326_),
    .A1(_1324_),
    .B1(_1323_),
    .X(_1330_));
 sg13g2_xnor2_1 _2178_ (.Y(_1331_),
    .A(\sin_y_acc[22] ),
    .B(\cos_x_acc[22] ));
 sg13g2_o21ai_1 _2179_ (.B1(_1331_),
    .Y(_1332_),
    .A1(_1329_),
    .A2(_1330_));
 sg13g2_or3_1 _2180_ (.A(_1329_),
    .B(_1330_),
    .C(_1331_),
    .X(_1333_));
 sg13g2_and2_1 _2181_ (.A(_1332_),
    .B(_1333_),
    .X(_1334_));
 sg13g2_nand2_2 _2182_ (.Y(_1335_),
    .A(_1332_),
    .B(_1333_));
 sg13g2_a21oi_1 _2183_ (.A1(_1322_),
    .A2(_1327_),
    .Y(_1336_),
    .B1(_1326_));
 sg13g2_xnor2_1 _2184_ (.Y(_1337_),
    .A(_1325_),
    .B(_1336_));
 sg13g2_xor2_1 _2185_ (.B(_1336_),
    .A(_1325_),
    .X(_1338_));
 sg13g2_xor2_1 _2186_ (.B(_1327_),
    .A(_1322_),
    .X(_1339_));
 sg13g2_xnor2_1 _2187_ (.Y(_1340_),
    .A(_1322_),
    .B(_1327_));
 sg13g2_a21oi_1 _2188_ (.A1(_1337_),
    .A2(_1339_),
    .Y(_1341_),
    .B1(_1334_));
 sg13g2_nor2_1 _2189_ (.A(\cos_y_acc[15] ),
    .B(\sin_x_acc[15] ),
    .Y(_1342_));
 sg13g2_xnor2_1 _2190_ (.Y(_1343_),
    .A(\cos_y_acc[15] ),
    .B(\sin_x_acc[15] ));
 sg13g2_nand2_1 _2191_ (.Y(_1344_),
    .A(\cos_y_acc[14] ),
    .B(\sin_x_acc[14] ));
 sg13g2_xnor2_1 _2192_ (.Y(_1345_),
    .A(\cos_y_acc[14] ),
    .B(\sin_x_acc[14] ));
 sg13g2_nor2_1 _2193_ (.A(_1343_),
    .B(_1345_),
    .Y(_1346_));
 sg13g2_nand2_1 _2194_ (.Y(_1347_),
    .A(\cos_y_acc[13] ),
    .B(\sin_x_acc[13] ));
 sg13g2_a22oi_1 _2195_ (.Y(_1348_),
    .B1(\sin_x_acc[12] ),
    .B2(\cos_y_acc[12] ),
    .A2(\sin_x_acc[13] ),
    .A1(\cos_y_acc[13] ));
 sg13g2_inv_1 _2196_ (.Y(_1349_),
    .A(_1348_));
 sg13g2_nor2_1 _2197_ (.A(\cos_y_acc[13] ),
    .B(\sin_x_acc[13] ),
    .Y(_1350_));
 sg13g2_nor2_1 _2198_ (.A(_1348_),
    .B(_1350_),
    .Y(_1351_));
 sg13g2_nor2_1 _2199_ (.A(_1342_),
    .B(_1344_),
    .Y(_1352_));
 sg13g2_a221oi_1 _2200_ (.B2(_1351_),
    .C1(_1352_),
    .B1(_1346_),
    .A1(\cos_y_acc[15] ),
    .Y(_1353_),
    .A2(\sin_x_acc[15] ));
 sg13g2_nor2_1 _2201_ (.A(\cos_y_acc[12] ),
    .B(\sin_x_acc[12] ),
    .Y(_1354_));
 sg13g2_xnor2_1 _2202_ (.Y(_1355_),
    .A(\cos_y_acc[13] ),
    .B(\sin_x_acc[13] ));
 sg13g2_nor3_1 _2203_ (.A(_1349_),
    .B(_1350_),
    .C(_1354_),
    .Y(_1356_));
 sg13g2_nand2_1 _2204_ (.Y(_1357_),
    .A(_1346_),
    .B(_1356_));
 sg13g2_and2_1 _2205_ (.A(\cos_y_acc[1] ),
    .B(\sin_x_acc[1] ),
    .X(_1358_));
 sg13g2_nand2_1 _2206_ (.Y(_1359_),
    .A(\cos_y_acc[0] ),
    .B(\sin_x_acc[0] ));
 sg13g2_a22oi_1 _2207_ (.Y(_1360_),
    .B1(\sin_x_acc[0] ),
    .B2(\cos_y_acc[0] ),
    .A2(\sin_x_acc[1] ),
    .A1(\cos_y_acc[1] ));
 sg13g2_nor2_1 _2208_ (.A(\cos_y_acc[1] ),
    .B(\sin_x_acc[1] ),
    .Y(_1361_));
 sg13g2_nor2_1 _2209_ (.A(\cos_y_acc[2] ),
    .B(\sin_x_acc[2] ),
    .Y(_1362_));
 sg13g2_nor3_1 _2210_ (.A(_1360_),
    .B(_1361_),
    .C(_1362_),
    .Y(_1363_));
 sg13g2_a22oi_1 _2211_ (.Y(_1364_),
    .B1(\sin_x_acc[2] ),
    .B2(\cos_y_acc[2] ),
    .A2(\sin_x_acc[3] ),
    .A1(\cos_y_acc[3] ));
 sg13g2_nand2b_1 _2212_ (.Y(_1365_),
    .B(_1364_),
    .A_N(_1363_));
 sg13g2_a22oi_1 _2213_ (.Y(_1366_),
    .B1(\sin_x_acc[7] ),
    .B2(\cos_y_acc[7] ),
    .A2(\sin_x_acc[6] ),
    .A1(\cos_y_acc[6] ));
 sg13g2_or2_1 _2214_ (.X(_1367_),
    .B(\sin_x_acc[7] ),
    .A(\cos_y_acc[7] ));
 sg13g2_or2_1 _2215_ (.X(_1368_),
    .B(\sin_x_acc[6] ),
    .A(\cos_y_acc[6] ));
 sg13g2_and3_1 _2216_ (.X(_1369_),
    .A(_1366_),
    .B(_1367_),
    .C(_1368_));
 sg13g2_a22oi_1 _2217_ (.Y(_1370_),
    .B1(\sin_x_acc[5] ),
    .B2(\cos_y_acc[5] ),
    .A2(\sin_x_acc[4] ),
    .A1(\cos_y_acc[4] ));
 sg13g2_nor2_1 _2218_ (.A(\cos_y_acc[5] ),
    .B(\sin_x_acc[5] ),
    .Y(_1371_));
 sg13g2_a221oi_1 _2219_ (.B2(_1205_),
    .C1(_1371_),
    .B1(_1224_),
    .A1(_1206_),
    .Y(_1372_),
    .A2(_1213_));
 sg13g2_and3_1 _2220_ (.X(_1373_),
    .A(_1369_),
    .B(_1370_),
    .C(_1372_));
 sg13g2_nor2b_1 _2221_ (.A(_1366_),
    .B_N(_1367_),
    .Y(_1374_));
 sg13g2_nor2_1 _2222_ (.A(_1370_),
    .B(_1371_),
    .Y(_1375_));
 sg13g2_a221oi_1 _2223_ (.B2(_1369_),
    .C1(_1374_),
    .B1(_1375_),
    .A1(_1365_),
    .Y(_1376_),
    .A2(_1373_));
 sg13g2_and2_1 _2224_ (.A(\cos_y_acc[11] ),
    .B(\sin_x_acc[11] ),
    .X(_1377_));
 sg13g2_a22oi_1 _2225_ (.Y(_1378_),
    .B1(\sin_x_acc[11] ),
    .B2(\cos_y_acc[11] ),
    .A2(\sin_x_acc[10] ),
    .A1(\cos_y_acc[10] ));
 sg13g2_nand2_1 _2226_ (.Y(_1379_),
    .A(\cos_y_acc[9] ),
    .B(\sin_x_acc[9] ));
 sg13g2_nand2_1 _2227_ (.Y(_1380_),
    .A(\cos_y_acc[8] ),
    .B(\sin_x_acc[8] ));
 sg13g2_nand3_1 _2228_ (.B(_1379_),
    .C(_1380_),
    .A(_1378_),
    .Y(_1381_));
 sg13g2_or2_1 _2229_ (.X(_1382_),
    .B(\sin_x_acc[11] ),
    .A(\cos_y_acc[11] ));
 sg13g2_o21ai_1 _2230_ (.B1(_1382_),
    .Y(_1383_),
    .A1(\cos_y_acc[8] ),
    .A2(\sin_x_acc[8] ));
 sg13g2_nor2_1 _2231_ (.A(\cos_y_acc[10] ),
    .B(\sin_x_acc[10] ),
    .Y(_1384_));
 sg13g2_nor2_1 _2232_ (.A(\cos_y_acc[9] ),
    .B(\sin_x_acc[9] ),
    .Y(_1385_));
 sg13g2_or4_1 _2233_ (.A(_1381_),
    .B(_1383_),
    .C(_1384_),
    .D(_1385_),
    .X(_1386_));
 sg13g2_o21ai_1 _2234_ (.B1(_1378_),
    .Y(_1387_),
    .A1(_1384_),
    .A2(_1385_));
 sg13g2_nand3_1 _2235_ (.B(_1382_),
    .C(_1387_),
    .A(_1381_),
    .Y(_1388_));
 sg13g2_o21ai_1 _2236_ (.B1(_1388_),
    .Y(_1389_),
    .A1(_1376_),
    .A2(_1386_));
 sg13g2_and2_1 _2237_ (.A(_1353_),
    .B(_1388_),
    .X(_1390_));
 sg13g2_o21ai_1 _2238_ (.B1(_1390_),
    .Y(_1391_),
    .A1(_1376_),
    .A2(_1386_));
 sg13g2_nand2_1 _2239_ (.Y(_1392_),
    .A(_1353_),
    .B(_1357_));
 sg13g2_nand2_1 _2240_ (.Y(_1393_),
    .A(\cos_y_acc[16] ),
    .B(\sin_x_acc[16] ));
 sg13g2_xor2_1 _2241_ (.B(\sin_x_acc[16] ),
    .A(\cos_y_acc[16] ),
    .X(_1394_));
 sg13g2_xor2_1 _2242_ (.B(\sin_x_acc[17] ),
    .A(\cos_y_acc[17] ),
    .X(_1395_));
 sg13g2_nand4_1 _2243_ (.B(_1392_),
    .C(_1394_),
    .A(_1391_),
    .Y(_1396_),
    .D(_1395_));
 sg13g2_a21oi_1 _2244_ (.A1(_1195_),
    .A2(_1220_),
    .Y(_1397_),
    .B1(_1393_));
 sg13g2_a21oi_1 _2245_ (.A1(\cos_y_acc[17] ),
    .A2(\sin_x_acc[17] ),
    .Y(_1398_),
    .B1(_1397_));
 sg13g2_nand2_1 _2246_ (.Y(_1399_),
    .A(_1396_),
    .B(_1398_));
 sg13g2_nand2_1 _2247_ (.Y(_1400_),
    .A(\cos_y_acc[18] ),
    .B(\sin_x_acc[18] ));
 sg13g2_xnor2_1 _2248_ (.Y(_1401_),
    .A(\cos_y_acc[18] ),
    .B(\sin_x_acc[18] ));
 sg13g2_a21o_1 _2249_ (.A2(_1398_),
    .A1(_1396_),
    .B1(_1401_),
    .X(_1402_));
 sg13g2_xnor2_1 _2250_ (.Y(_1403_),
    .A(_1399_),
    .B(_1401_));
 sg13g2_nand3_1 _2251_ (.B(_1392_),
    .C(_1394_),
    .A(_1391_),
    .Y(_1404_));
 sg13g2_nand2_1 _2252_ (.Y(_1405_),
    .A(_1393_),
    .B(_1404_));
 sg13g2_xor2_1 _2253_ (.B(_1405_),
    .A(_1395_),
    .X(_1406_));
 sg13g2_or2_1 _2254_ (.X(_1407_),
    .B(_1406_),
    .A(_1403_));
 sg13g2_xor2_1 _2255_ (.B(\sin_x_acc[19] ),
    .A(\cos_y_acc[19] ),
    .X(_1408_));
 sg13g2_and3_1 _2256_ (.X(_1409_),
    .A(_1400_),
    .B(_1402_),
    .C(_1408_));
 sg13g2_a21oi_1 _2257_ (.A1(_1400_),
    .A2(_1402_),
    .Y(_1410_),
    .B1(_1408_));
 sg13g2_or2_1 _2258_ (.X(_1411_),
    .B(_1410_),
    .A(_1409_));
 sg13g2_or4_1 _2259_ (.A(_1403_),
    .B(_1406_),
    .C(_1409_),
    .D(_1410_),
    .X(_1412_));
 sg13g2_xnor2_1 _2260_ (.Y(_1413_),
    .A(_1407_),
    .B(_1411_));
 sg13g2_nand2b_1 _2261_ (.Y(_1414_),
    .B(_1408_),
    .A_N(_1401_));
 sg13g2_a21o_1 _2262_ (.A2(_1398_),
    .A1(_1396_),
    .B1(_1414_),
    .X(_1415_));
 sg13g2_a21oi_1 _2263_ (.A1(_1194_),
    .A2(_1218_),
    .Y(_1416_),
    .B1(_1400_));
 sg13g2_a21oi_1 _2264_ (.A1(\cos_y_acc[19] ),
    .A2(\sin_x_acc[19] ),
    .Y(_1417_),
    .B1(_1416_));
 sg13g2_nand2_1 _2265_ (.Y(_1418_),
    .A(_1415_),
    .B(_1417_));
 sg13g2_and2_1 _2266_ (.A(net248),
    .B(\sin_x_acc[20] ),
    .X(_1419_));
 sg13g2_nand2_1 _2267_ (.Y(_1420_),
    .A(net248),
    .B(\sin_x_acc[20] ));
 sg13g2_xnor2_1 _2268_ (.Y(_1421_),
    .A(net248),
    .B(\sin_x_acc[20] ));
 sg13g2_a21oi_1 _2269_ (.A1(_1415_),
    .A2(_1417_),
    .Y(_1422_),
    .B1(_1421_));
 sg13g2_a21o_1 _2270_ (.A2(_1417_),
    .A1(_1415_),
    .B1(_1421_),
    .X(_1423_));
 sg13g2_xnor2_1 _2271_ (.Y(_1424_),
    .A(_1418_),
    .B(_1421_));
 sg13g2_xor2_1 _2272_ (.B(_1421_),
    .A(_1418_),
    .X(_1425_));
 sg13g2_nand2_1 _2273_ (.Y(_1426_),
    .A(_1412_),
    .B(_1425_));
 sg13g2_nand2b_1 _2274_ (.Y(_1427_),
    .B(_1425_),
    .A_N(_1412_));
 sg13g2_xnor2_1 _2275_ (.Y(_1428_),
    .A(_1412_),
    .B(_1424_));
 sg13g2_and2_1 _2276_ (.A(_1413_),
    .B(_1428_),
    .X(_1429_));
 sg13g2_and2_1 _2277_ (.A(\cos_y_acc[21] ),
    .B(\sin_x_acc[21] ),
    .X(_1430_));
 sg13g2_nor2_2 _2278_ (.A(\cos_y_acc[21] ),
    .B(\sin_x_acc[21] ),
    .Y(_1431_));
 sg13g2_nor2_1 _2279_ (.A(_1430_),
    .B(_1431_),
    .Y(_1432_));
 sg13g2_nor4_1 _2280_ (.A(_1419_),
    .B(_1422_),
    .C(_1430_),
    .D(_1431_),
    .Y(_1433_));
 sg13g2_a21oi_1 _2281_ (.A1(_1420_),
    .A2(_1423_),
    .Y(_1434_),
    .B1(_1432_));
 sg13g2_nor2_2 _2282_ (.A(_1433_),
    .B(_1434_),
    .Y(_1435_));
 sg13g2_nor4_1 _2283_ (.A(_1412_),
    .B(_1424_),
    .C(_1433_),
    .D(_1434_),
    .Y(_1436_));
 sg13g2_xnor2_1 _2284_ (.Y(_1437_),
    .A(_1427_),
    .B(_1435_));
 sg13g2_xor2_1 _2285_ (.B(_1435_),
    .A(_1427_),
    .X(_1438_));
 sg13g2_xnor2_1 _2286_ (.Y(_1439_),
    .A(net247),
    .B(\sin_x_acc[22] ));
 sg13g2_inv_1 _2287_ (.Y(_1440_),
    .A(_1439_));
 sg13g2_nor3_1 _2288_ (.A(_1419_),
    .B(_1422_),
    .C(_1430_),
    .Y(_1441_));
 sg13g2_a21oi_1 _2289_ (.A1(_1420_),
    .A2(_1423_),
    .Y(_1442_),
    .B1(_1431_));
 sg13g2_nor3_1 _2290_ (.A(_1431_),
    .B(_1439_),
    .C(_1441_),
    .Y(_1443_));
 sg13g2_o21ai_1 _2291_ (.B1(_1440_),
    .Y(_1444_),
    .A1(_1430_),
    .A2(_1442_));
 sg13g2_nor3_1 _2292_ (.A(_1430_),
    .B(_1440_),
    .C(_1442_),
    .Y(_1445_));
 sg13g2_o21ai_1 _2293_ (.B1(_1439_),
    .Y(_1446_),
    .A1(_1431_),
    .A2(_1441_));
 sg13g2_nand2_1 _2294_ (.Y(_1447_),
    .A(_1444_),
    .B(_1446_));
 sg13g2_nand3b_1 _2295_ (.B(_1444_),
    .C(_1446_),
    .Y(_1448_),
    .A_N(_1436_));
 sg13g2_o21ai_1 _2296_ (.B1(_1436_),
    .Y(_1449_),
    .A1(_1443_),
    .A2(_1445_));
 sg13g2_and2_1 _2297_ (.A(_1448_),
    .B(_1449_),
    .X(_1450_));
 sg13g2_nor2_1 _2298_ (.A(_1437_),
    .B(_1450_),
    .Y(_1451_));
 sg13g2_or2_1 _2299_ (.X(_1452_),
    .B(_1450_),
    .A(_1437_));
 sg13g2_a21oi_1 _2300_ (.A1(_1429_),
    .A2(_1451_),
    .Y(_1453_),
    .B1(_1341_));
 sg13g2_xnor2_1 _2301_ (.Y(_1454_),
    .A(\sin_y_acc[19] ),
    .B(\cos_x_acc[19] ));
 sg13g2_a21oi_1 _2302_ (.A1(_1249_),
    .A2(_1319_),
    .Y(_1455_),
    .B1(_1454_));
 sg13g2_and3_2 _2303_ (.X(_1456_),
    .A(_1249_),
    .B(_1319_),
    .C(_1454_));
 sg13g2_nor2_2 _2304_ (.A(_1455_),
    .B(_1456_),
    .Y(_1457_));
 sg13g2_or2_1 _2305_ (.X(_1458_),
    .B(_1456_),
    .A(_1455_));
 sg13g2_xnor2_1 _2306_ (.Y(_1459_),
    .A(_1250_),
    .B(_1318_));
 sg13g2_xor2_1 _2307_ (.B(_1318_),
    .A(_1250_),
    .X(_1460_));
 sg13g2_a21oi_1 _2308_ (.A1(_1310_),
    .A2(_1312_),
    .Y(_1461_),
    .B1(_1311_));
 sg13g2_xor2_1 _2309_ (.B(_1461_),
    .A(_1313_),
    .X(_1462_));
 sg13g2_xor2_1 _2310_ (.B(_1312_),
    .A(_1310_),
    .X(_1463_));
 sg13g2_xnor2_1 _2311_ (.Y(_1464_),
    .A(_1310_),
    .B(_1312_));
 sg13g2_o21ai_1 _2312_ (.B1(_1260_),
    .Y(_1465_),
    .A1(_1265_),
    .A2(_1308_));
 sg13g2_a21oi_1 _2313_ (.A1(_1255_),
    .A2(_1465_),
    .Y(_1466_),
    .B1(_1254_));
 sg13g2_xor2_1 _2314_ (.B(_1466_),
    .A(_1253_),
    .X(_1467_));
 sg13g2_nand2b_1 _2315_ (.Y(_1468_),
    .B(_1463_),
    .A_N(_1467_));
 sg13g2_a21oi_1 _2316_ (.A1(_1462_),
    .A2(_1468_),
    .Y(_1469_),
    .B1(_1460_));
 sg13g2_o21ai_1 _2317_ (.B1(_1339_),
    .Y(_1470_),
    .A1(_1458_),
    .A2(_1469_));
 sg13g2_o21ai_1 _2318_ (.B1(_1460_),
    .Y(_1471_),
    .A1(_1462_),
    .A2(_1464_));
 sg13g2_nor2_1 _2319_ (.A(_1438_),
    .B(_1447_),
    .Y(_1472_));
 sg13g2_a21o_1 _2320_ (.A2(_1392_),
    .A1(_1391_),
    .B1(_1394_),
    .X(_1473_));
 sg13g2_and2_1 _2321_ (.A(_1404_),
    .B(_1473_),
    .X(_1474_));
 sg13g2_inv_2 _2322_ (.Y(_1475_),
    .A(_1474_));
 sg13g2_a21oi_1 _2323_ (.A1(_1356_),
    .A2(_1389_),
    .Y(_1476_),
    .B1(_1351_));
 sg13g2_o21ai_1 _2324_ (.B1(_1344_),
    .Y(_1477_),
    .A1(_1345_),
    .A2(_1476_));
 sg13g2_xnor2_1 _2325_ (.Y(_1478_),
    .A(_1343_),
    .B(_1477_));
 sg13g2_nand2_1 _2326_ (.Y(_1479_),
    .A(_1474_),
    .B(_1478_));
 sg13g2_nor2_1 _2327_ (.A(_1407_),
    .B(_1479_),
    .Y(_1480_));
 sg13g2_or2_1 _2328_ (.X(_1481_),
    .B(_1480_),
    .A(_1413_));
 sg13g2_o21ai_1 _2329_ (.B1(_1472_),
    .Y(_1482_),
    .A1(_1428_),
    .A2(_1481_));
 sg13g2_and2_1 _2330_ (.A(_1452_),
    .B(_1482_),
    .X(_1483_));
 sg13g2_a21oi_1 _2331_ (.A1(_1458_),
    .A2(_1471_),
    .Y(_1484_),
    .B1(_1483_));
 sg13g2_nor2_1 _2332_ (.A(_1337_),
    .B(_1470_),
    .Y(_1485_));
 sg13g2_and2_1 _2333_ (.A(_1484_),
    .B(_1485_),
    .X(_1486_));
 sg13g2_o21ai_1 _2334_ (.B1(_1341_),
    .Y(_1487_),
    .A1(_1338_),
    .A2(_1457_));
 sg13g2_nor3_1 _2335_ (.A(_1455_),
    .B(_1456_),
    .C(_1459_),
    .Y(_1488_));
 sg13g2_nor2_1 _2336_ (.A(_1337_),
    .B(_1339_),
    .Y(_1489_));
 sg13g2_and2_1 _2337_ (.A(_1488_),
    .B(_1489_),
    .X(_1490_));
 sg13g2_nand2b_1 _2338_ (.Y(_1491_),
    .B(_1406_),
    .A_N(_1403_));
 sg13g2_nand2b_1 _2339_ (.Y(_1492_),
    .B(_1475_),
    .A_N(_1491_));
 sg13g2_a21oi_1 _2340_ (.A1(_1413_),
    .A2(_1492_),
    .Y(_1493_),
    .B1(_1428_));
 sg13g2_a22oi_1 _2341_ (.Y(_1494_),
    .B1(_1450_),
    .B2(_1493_),
    .A2(_1447_),
    .A1(_1437_));
 sg13g2_and2_1 _2342_ (.A(_1403_),
    .B(_1406_),
    .X(_1495_));
 sg13g2_nand2_1 _2343_ (.Y(_1496_),
    .A(_1411_),
    .B(_1495_));
 sg13g2_nor2b_1 _2344_ (.A(_1426_),
    .B_N(_1496_),
    .Y(_1497_));
 sg13g2_nor2_1 _2345_ (.A(_1479_),
    .B(_1496_),
    .Y(_1498_));
 sg13g2_o21ai_1 _2346_ (.B1(_1438_),
    .Y(_1499_),
    .A1(_1426_),
    .A2(_1498_));
 sg13g2_nand3_1 _2347_ (.B(_1494_),
    .C(_1499_),
    .A(_1450_),
    .Y(_1500_));
 sg13g2_nor3_1 _2348_ (.A(_1487_),
    .B(_1490_),
    .C(_1500_),
    .Y(_1501_));
 sg13g2_xor2_1 _2349_ (.B(_1476_),
    .A(_1345_),
    .X(_1502_));
 sg13g2_nor2_2 _2350_ (.A(_1478_),
    .B(_1502_),
    .Y(_1503_));
 sg13g2_xnor2_1 _2351_ (.Y(_1504_),
    .A(_1403_),
    .B(_1406_));
 sg13g2_and3_2 _2352_ (.X(_1505_),
    .A(_1413_),
    .B(_1428_),
    .C(_1504_));
 sg13g2_a22oi_1 _2353_ (.Y(_1506_),
    .B1(_1505_),
    .B2(_1438_),
    .A2(_1449_),
    .A1(_1448_));
 sg13g2_and4_1 _2354_ (.A(_1438_),
    .B(_1448_),
    .C(_1449_),
    .D(_1505_),
    .X(_1507_));
 sg13g2_nand4_1 _2355_ (.B(_1448_),
    .C(_1449_),
    .A(_1438_),
    .Y(_1508_),
    .D(_1505_));
 sg13g2_nor2_2 _2356_ (.A(_1506_),
    .B(_1507_),
    .Y(_1509_));
 sg13g2_nor3_1 _2357_ (.A(_1503_),
    .B(_1506_),
    .C(_1507_),
    .Y(_1510_));
 sg13g2_xnor2_1 _2358_ (.Y(_1511_),
    .A(_1474_),
    .B(_1510_));
 sg13g2_xnor2_1 _2359_ (.Y(_1512_),
    .A(_1475_),
    .B(_1510_));
 sg13g2_nand2b_1 _2360_ (.Y(_1513_),
    .B(_1437_),
    .A_N(_1505_));
 sg13g2_nand2_1 _2361_ (.Y(_1514_),
    .A(_1475_),
    .B(_1503_));
 sg13g2_nand4_1 _2362_ (.B(_1475_),
    .C(_1495_),
    .A(_1411_),
    .Y(_1515_),
    .D(_1503_));
 sg13g2_nor2_1 _2363_ (.A(_1425_),
    .B(_1515_),
    .Y(_1516_));
 sg13g2_a21oi_1 _2364_ (.A1(_1438_),
    .A2(_1505_),
    .Y(_1517_),
    .B1(_1516_));
 sg13g2_nand2_1 _2365_ (.Y(_1518_),
    .A(_1513_),
    .B(_1517_));
 sg13g2_nor3_1 _2366_ (.A(_1425_),
    .B(_1435_),
    .C(_1515_),
    .Y(_1519_));
 sg13g2_nor3_1 _2367_ (.A(_1506_),
    .B(_1507_),
    .C(_1519_),
    .Y(_1520_));
 sg13g2_and2_1 _2368_ (.A(_1506_),
    .B(_1513_),
    .X(_1521_));
 sg13g2_a21oi_2 _2369_ (.B1(_1521_),
    .Y(_1522_),
    .A2(_1520_),
    .A1(_1518_));
 sg13g2_a21o_2 _2370_ (.A2(_1520_),
    .A1(_1518_),
    .B1(_1521_),
    .X(_1523_));
 sg13g2_nor2_1 _2371_ (.A(_1497_),
    .B(_1505_),
    .Y(_1524_));
 sg13g2_inv_1 _2372_ (.Y(_1525_),
    .A(_1524_));
 sg13g2_a21oi_1 _2373_ (.A1(_1515_),
    .A2(_1524_),
    .Y(_1526_),
    .B1(_1516_));
 sg13g2_a21o_1 _2374_ (.A2(_1524_),
    .A1(_1515_),
    .B1(_1516_),
    .X(_1527_));
 sg13g2_mux2_1 _2375_ (.A0(_1525_),
    .A1(_1527_),
    .S(_1509_),
    .X(_1528_));
 sg13g2_mux2_1 _2376_ (.A0(_1524_),
    .A1(_1526_),
    .S(_1509_),
    .X(_1529_));
 sg13g2_nand3b_1 _2377_ (.B(_1508_),
    .C(_1514_),
    .Y(_1530_),
    .A_N(_1506_));
 sg13g2_xor2_1 _2378_ (.B(_1530_),
    .A(_1406_),
    .X(_1531_));
 sg13g2_nand2_1 _2379_ (.Y(_1532_),
    .A(_1512_),
    .B(net181));
 sg13g2_nand2_1 _2380_ (.Y(_1533_),
    .A(_1523_),
    .B(_1531_));
 sg13g2_nor2_1 _2381_ (.A(_1532_),
    .B(_1533_),
    .Y(_1534_));
 sg13g2_a22oi_1 _2382_ (.Y(_1535_),
    .B1(net181),
    .B2(_1531_),
    .A2(_1523_),
    .A1(_1512_));
 sg13g2_nor2_1 _2383_ (.A(_1534_),
    .B(_1535_),
    .Y(_1536_));
 sg13g2_nand3b_1 _2384_ (.B(_1508_),
    .C(_1502_),
    .Y(_1537_),
    .A_N(_1506_));
 sg13g2_xor2_1 _2385_ (.B(_1537_),
    .A(_1478_),
    .X(_1538_));
 sg13g2_xnor2_1 _2386_ (.Y(_1539_),
    .A(_1478_),
    .B(_1537_));
 sg13g2_nor4_1 _2387_ (.A(_1511_),
    .B(_1522_),
    .C(_1528_),
    .D(_1538_),
    .Y(_1540_));
 sg13g2_xor2_1 _2388_ (.B(_1495_),
    .A(_1411_),
    .X(_1541_));
 sg13g2_inv_1 _2389_ (.Y(_1542_),
    .A(_1541_));
 sg13g2_nand3_1 _2390_ (.B(_1475_),
    .C(_1503_),
    .A(_1406_),
    .Y(_1543_));
 sg13g2_o21ai_1 _2391_ (.B1(_1541_),
    .Y(_1544_),
    .A1(_1411_),
    .A2(_1514_));
 sg13g2_and2_1 _2392_ (.A(_1515_),
    .B(_1544_),
    .X(_1545_));
 sg13g2_inv_1 _2393_ (.Y(_1546_),
    .A(_1545_));
 sg13g2_mux2_1 _2394_ (.A0(_1541_),
    .A1(_1545_),
    .S(_1509_),
    .X(_1547_));
 sg13g2_mux2_1 _2395_ (.A0(_1542_),
    .A1(_1546_),
    .S(_1509_),
    .X(_1548_));
 sg13g2_nand2_1 _2396_ (.Y(_1549_),
    .A(_1531_),
    .B(_1547_));
 sg13g2_a22oi_1 _2397_ (.Y(_1550_),
    .B1(_1539_),
    .B2(_1523_),
    .A2(net181),
    .A1(_1512_));
 sg13g2_or3_1 _2398_ (.A(_1540_),
    .B(_1549_),
    .C(_1550_),
    .X(_1551_));
 sg13g2_nor2b_1 _2399_ (.A(_1540_),
    .B_N(_1551_),
    .Y(_1552_));
 sg13g2_nor2b_1 _2400_ (.A(_1552_),
    .B_N(_1536_),
    .Y(_1553_));
 sg13g2_nor2_1 _2401_ (.A(_1538_),
    .B(_1548_),
    .Y(_1554_));
 sg13g2_nor4_1 _2402_ (.A(_1511_),
    .B(_1528_),
    .C(_1538_),
    .D(_1548_),
    .Y(_1555_));
 sg13g2_nand4_1 _2403_ (.B(net181),
    .C(_1539_),
    .A(_1512_),
    .Y(_1556_),
    .D(_1547_));
 sg13g2_nand3b_1 _2404_ (.B(_1508_),
    .C(_1543_),
    .Y(_1557_),
    .A_N(_1506_));
 sg13g2_xnor2_1 _2405_ (.Y(_1558_),
    .A(_1504_),
    .B(_1557_));
 sg13g2_nand2b_1 _2406_ (.Y(_1559_),
    .B(_1531_),
    .A_N(_1558_));
 sg13g2_a22oi_1 _2407_ (.Y(_1560_),
    .B1(_1547_),
    .B2(_1512_),
    .A2(_1539_),
    .A1(_1529_));
 sg13g2_or3_1 _2408_ (.A(_1555_),
    .B(_1559_),
    .C(_1560_),
    .X(_1561_));
 sg13g2_o21ai_1 _2409_ (.B1(_1556_),
    .Y(_1562_),
    .A1(_1559_),
    .A2(_1560_));
 sg13g2_o21ai_1 _2410_ (.B1(_1549_),
    .Y(_1563_),
    .A1(_1540_),
    .A2(_1550_));
 sg13g2_and3_1 _2411_ (.X(_1564_),
    .A(_1551_),
    .B(_1562_),
    .C(_1563_));
 sg13g2_nand3_1 _2412_ (.B(_1562_),
    .C(_1563_),
    .A(_1551_),
    .Y(_1565_));
 sg13g2_nor2_1 _2413_ (.A(_1538_),
    .B(_1558_),
    .Y(_1566_));
 sg13g2_nor2_1 _2414_ (.A(_1511_),
    .B(_1558_),
    .Y(_1567_));
 sg13g2_and2_1 _2415_ (.A(_1554_),
    .B(_1567_),
    .X(_1568_));
 sg13g2_o21ai_1 _2416_ (.B1(_1559_),
    .Y(_1569_),
    .A1(_1555_),
    .A2(_1560_));
 sg13g2_and2_1 _2417_ (.A(_1561_),
    .B(_1569_),
    .X(_1570_));
 sg13g2_nand3_1 _2418_ (.B(_1568_),
    .C(_1569_),
    .A(_1561_),
    .Y(_1571_));
 sg13g2_a21oi_1 _2419_ (.A1(_1551_),
    .A2(_1563_),
    .Y(_1572_),
    .B1(_1562_));
 sg13g2_nor3_1 _2420_ (.A(_1564_),
    .B(_1571_),
    .C(_1572_),
    .Y(_1573_));
 sg13g2_o21ai_1 _2421_ (.B1(_1565_),
    .Y(_1574_),
    .A1(_1571_),
    .A2(_1572_));
 sg13g2_xnor2_1 _2422_ (.Y(_1575_),
    .A(_1536_),
    .B(_1552_));
 sg13g2_a21oi_1 _2423_ (.A1(_1574_),
    .A2(_1575_),
    .Y(_1576_),
    .B1(_1553_));
 sg13g2_nand2b_1 _2424_ (.Y(_1577_),
    .B(_1532_),
    .A_N(_1533_));
 sg13g2_a21oi_1 _2425_ (.A1(_1532_),
    .A2(_1576_),
    .Y(_1578_),
    .B1(_1533_));
 sg13g2_nor2_1 _2426_ (.A(_1522_),
    .B(_1528_),
    .Y(_1579_));
 sg13g2_nor2_1 _2427_ (.A(_1522_),
    .B(_1558_),
    .Y(_1580_));
 sg13g2_nand2_2 _2428_ (.Y(_1581_),
    .A(_1547_),
    .B(_1558_));
 sg13g2_a21oi_1 _2429_ (.A1(net181),
    .A2(_1581_),
    .Y(_1582_),
    .B1(_1580_));
 sg13g2_a21o_1 _2430_ (.A2(_1580_),
    .A1(net181),
    .B1(_1582_),
    .X(_1583_));
 sg13g2_nand2b_1 _2431_ (.Y(_1584_),
    .B(_1578_),
    .A_N(_1583_));
 sg13g2_xnor2_1 _2432_ (.Y(_1585_),
    .A(_1255_),
    .B(_1465_));
 sg13g2_and2_1 _2433_ (.A(_1467_),
    .B(net182),
    .X(_1586_));
 sg13g2_and4_1 _2434_ (.A(_1462_),
    .B(_1464_),
    .C(_1467_),
    .D(net182),
    .X(_1587_));
 sg13g2_nor2_1 _2435_ (.A(_1334_),
    .B(_1587_),
    .Y(_1588_));
 sg13g2_xnor2_1 _2436_ (.Y(_1589_),
    .A(_1459_),
    .B(_1588_));
 sg13g2_inv_1 _2437_ (.Y(_1590_),
    .A(net179));
 sg13g2_a22oi_1 _2438_ (.Y(_1591_),
    .B1(_1488_),
    .B2(_1587_),
    .A2(_1333_),
    .A1(_1332_));
 sg13g2_xnor2_1 _2439_ (.Y(_1592_),
    .A(_1339_),
    .B(_1591_));
 sg13g2_nor2_1 _2440_ (.A(_1339_),
    .B(_1458_),
    .Y(_1593_));
 sg13g2_nand3_1 _2441_ (.B(_1488_),
    .C(_1587_),
    .A(_1340_),
    .Y(_1594_));
 sg13g2_nand3_1 _2442_ (.B(_1338_),
    .C(_1594_),
    .A(_1335_),
    .Y(_1595_));
 sg13g2_a21o_1 _2443_ (.A2(_1594_),
    .A1(_1335_),
    .B1(_1338_),
    .X(_1596_));
 sg13g2_and2_1 _2444_ (.A(_1595_),
    .B(_1596_),
    .X(_1597_));
 sg13g2_inv_1 _2445_ (.Y(_1598_),
    .A(_1597_));
 sg13g2_nor2_1 _2446_ (.A(net180),
    .B(_1597_),
    .Y(_1599_));
 sg13g2_nand2_1 _2447_ (.Y(_1600_),
    .A(_1590_),
    .B(_1599_));
 sg13g2_a22oi_1 _2448_ (.Y(_1601_),
    .B1(_1460_),
    .B2(_1587_),
    .A2(_1333_),
    .A1(_1332_));
 sg13g2_xnor2_1 _2449_ (.Y(_1602_),
    .A(_1458_),
    .B(_1601_));
 sg13g2_xnor2_1 _2450_ (.Y(_1603_),
    .A(_1457_),
    .B(_1601_));
 sg13g2_nand2_1 _2451_ (.Y(_1604_),
    .A(net180),
    .B(_1597_));
 sg13g2_o21ai_1 _2452_ (.B1(_1589_),
    .Y(_1605_),
    .A1(net180),
    .A2(_1603_));
 sg13g2_nand2_1 _2453_ (.Y(_1606_),
    .A(net179),
    .B(_1603_));
 sg13g2_inv_1 _2454_ (.Y(_1607_),
    .A(_1606_));
 sg13g2_nand3_1 _2455_ (.B(_1604_),
    .C(_1605_),
    .A(_1600_),
    .Y(_1608_));
 sg13g2_xor2_1 _2456_ (.B(_1583_),
    .A(_1578_),
    .X(_1609_));
 sg13g2_o21ai_1 _2457_ (.B1(_1584_),
    .Y(_1610_),
    .A1(_1608_),
    .A2(_1609_));
 sg13g2_nand3b_1 _2458_ (.B(_1603_),
    .C(_1604_),
    .Y(_1611_),
    .A_N(_1599_));
 sg13g2_xnor2_1 _2459_ (.Y(_1612_),
    .A(_1523_),
    .B(_1528_));
 sg13g2_a22oi_1 _2460_ (.Y(_1613_),
    .B1(_1612_),
    .B2(_1547_),
    .A2(_1580_),
    .A1(net181));
 sg13g2_a21oi_1 _2461_ (.A1(_1600_),
    .A2(_1611_),
    .Y(_1614_),
    .B1(_1613_));
 sg13g2_nand3_1 _2462_ (.B(_1611_),
    .C(_1613_),
    .A(_1600_),
    .Y(_1615_));
 sg13g2_nand2b_1 _2463_ (.Y(_1616_),
    .B(_1615_),
    .A_N(_1614_));
 sg13g2_nor2b_1 _2464_ (.A(_1616_),
    .B_N(_1610_),
    .Y(_1617_));
 sg13g2_xor2_1 _2465_ (.B(_1616_),
    .A(_1610_),
    .X(_1618_));
 sg13g2_a21o_1 _2466_ (.A2(_1547_),
    .A1(net181),
    .B1(_1558_),
    .X(_1619_));
 sg13g2_a21oi_1 _2467_ (.A1(_1528_),
    .A2(_1548_),
    .Y(_1620_),
    .B1(_1619_));
 sg13g2_xor2_1 _2468_ (.B(_1577_),
    .A(_1576_),
    .X(_1621_));
 sg13g2_and2_1 _2469_ (.A(_1620_),
    .B(_1621_),
    .X(_1622_));
 sg13g2_xnor2_1 _2470_ (.Y(_1623_),
    .A(_1592_),
    .B(_1602_));
 sg13g2_nor2_1 _2471_ (.A(net179),
    .B(_1623_),
    .Y(_1624_));
 sg13g2_xor2_1 _2472_ (.B(_1621_),
    .A(_1620_),
    .X(_1625_));
 sg13g2_a21oi_1 _2473_ (.A1(_1624_),
    .A2(_1625_),
    .Y(_1626_),
    .B1(_1622_));
 sg13g2_xnor2_1 _2474_ (.Y(_1627_),
    .A(_1608_),
    .B(_1609_));
 sg13g2_nor2_1 _2475_ (.A(_1626_),
    .B(_1627_),
    .Y(_1628_));
 sg13g2_a21oi_1 _2476_ (.A1(_1464_),
    .A2(_1586_),
    .Y(_1629_),
    .B1(_1334_));
 sg13g2_xnor2_1 _2477_ (.Y(_1630_),
    .A(_1462_),
    .B(_1629_));
 sg13g2_nand2_1 _2478_ (.Y(_1631_),
    .A(_1598_),
    .B(_1630_));
 sg13g2_a21oi_1 _2479_ (.A1(_1332_),
    .A2(_1333_),
    .Y(_1632_),
    .B1(net182));
 sg13g2_xor2_1 _2480_ (.B(_1632_),
    .A(_1467_),
    .X(_1633_));
 sg13g2_nor2_1 _2481_ (.A(_1597_),
    .B(_1633_),
    .Y(_1634_));
 sg13g2_nor2_1 _2482_ (.A(_1334_),
    .B(_1586_),
    .Y(_1635_));
 sg13g2_xnor2_1 _2483_ (.Y(_1636_),
    .A(_1463_),
    .B(_1635_));
 sg13g2_nor2_1 _2484_ (.A(net180),
    .B(_1636_),
    .Y(_1637_));
 sg13g2_nor2_2 _2485_ (.A(net180),
    .B(_1633_),
    .Y(_1638_));
 sg13g2_nor2b_1 _2486_ (.A(net180),
    .B_N(_1630_),
    .Y(_1639_));
 sg13g2_nor3_1 _2487_ (.A(_1597_),
    .B(_1636_),
    .C(_1638_),
    .Y(_1640_));
 sg13g2_a22oi_1 _2488_ (.Y(_1641_),
    .B1(_1639_),
    .B2(_1640_),
    .A2(_1637_),
    .A1(_1634_));
 sg13g2_or2_1 _2489_ (.X(_1642_),
    .B(_1641_),
    .A(_1631_));
 sg13g2_nor2_1 _2490_ (.A(net182),
    .B(net180),
    .Y(_1643_));
 sg13g2_a21oi_1 _2491_ (.A1(_1595_),
    .A2(_1596_),
    .Y(_1644_),
    .B1(net182));
 sg13g2_nor2_1 _2492_ (.A(_1602_),
    .B(_1636_),
    .Y(_1645_));
 sg13g2_xor2_1 _2493_ (.B(_1644_),
    .A(_1638_),
    .X(_1646_));
 sg13g2_a22oi_1 _2494_ (.Y(_1647_),
    .B1(_1645_),
    .B2(_1646_),
    .A2(_1643_),
    .A1(_1634_));
 sg13g2_xor2_1 _2495_ (.B(_1637_),
    .A(_1634_),
    .X(_1648_));
 sg13g2_nor2b_1 _2496_ (.A(_1647_),
    .B_N(_1648_),
    .Y(_1649_));
 sg13g2_nand2_1 _2497_ (.Y(_1650_),
    .A(_1603_),
    .B(_1630_));
 sg13g2_inv_1 _2498_ (.Y(_1651_),
    .A(_1650_));
 sg13g2_xnor2_1 _2499_ (.Y(_1652_),
    .A(_1647_),
    .B(_1648_));
 sg13g2_a21oi_1 _2500_ (.A1(_1651_),
    .A2(_1652_),
    .Y(_1653_),
    .B1(_1649_));
 sg13g2_xnor2_1 _2501_ (.Y(_1654_),
    .A(_1639_),
    .B(_1640_));
 sg13g2_nor2_1 _2502_ (.A(_1653_),
    .B(_1654_),
    .Y(_1655_));
 sg13g2_nor2_1 _2503_ (.A(net182),
    .B(_1602_),
    .Y(_1656_));
 sg13g2_nor2_1 _2504_ (.A(_1602_),
    .B(_1633_),
    .Y(_1657_));
 sg13g2_nor2_1 _2505_ (.A(net179),
    .B(_1636_),
    .Y(_1658_));
 sg13g2_xor2_1 _2506_ (.B(_1657_),
    .A(_1643_),
    .X(_1659_));
 sg13g2_a22oi_1 _2507_ (.Y(_1660_),
    .B1(_1658_),
    .B2(_1659_),
    .A2(_1656_),
    .A1(_1638_));
 sg13g2_xnor2_1 _2508_ (.Y(_1661_),
    .A(_1645_),
    .B(_1646_));
 sg13g2_nor2_1 _2509_ (.A(_1660_),
    .B(_1661_),
    .Y(_1662_));
 sg13g2_nor2b_1 _2510_ (.A(net179),
    .B_N(_1630_),
    .Y(_1663_));
 sg13g2_xor2_1 _2511_ (.B(_1661_),
    .A(_1660_),
    .X(_1664_));
 sg13g2_a21oi_1 _2512_ (.A1(_1663_),
    .A2(_1664_),
    .Y(_1665_),
    .B1(_1662_));
 sg13g2_xnor2_1 _2513_ (.Y(_1666_),
    .A(_1651_),
    .B(_1652_));
 sg13g2_nor2_1 _2514_ (.A(_1665_),
    .B(_1666_),
    .Y(_1667_));
 sg13g2_xor2_1 _2515_ (.B(_1659_),
    .A(_1658_),
    .X(_1668_));
 sg13g2_nor2_1 _2516_ (.A(net179),
    .B(_1633_),
    .Y(_1669_));
 sg13g2_and2_1 _2517_ (.A(_1656_),
    .B(_1669_),
    .X(_1670_));
 sg13g2_nand2_1 _2518_ (.Y(_1671_),
    .A(_1668_),
    .B(_1670_));
 sg13g2_xor2_1 _2519_ (.B(_1664_),
    .A(_1663_),
    .X(_1672_));
 sg13g2_nor2b_1 _2520_ (.A(_1671_),
    .B_N(_1672_),
    .Y(_1673_));
 sg13g2_xor2_1 _2521_ (.B(_1666_),
    .A(_1665_),
    .X(_1674_));
 sg13g2_a21o_1 _2522_ (.A2(_1674_),
    .A1(_1673_),
    .B1(_1667_),
    .X(_1675_));
 sg13g2_xor2_1 _2523_ (.B(_1654_),
    .A(_1653_),
    .X(_1676_));
 sg13g2_a21oi_1 _2524_ (.A1(_1675_),
    .A2(_1676_),
    .Y(_1677_),
    .B1(_1655_));
 sg13g2_and2_1 _2525_ (.A(_1631_),
    .B(_1641_),
    .X(_1678_));
 sg13g2_xor2_1 _2526_ (.B(_1641_),
    .A(_1631_),
    .X(_1679_));
 sg13g2_o21ai_1 _2527_ (.B1(_1642_),
    .Y(_1680_),
    .A1(_1677_),
    .A2(_1678_));
 sg13g2_xor2_1 _2528_ (.B(_1627_),
    .A(_1626_),
    .X(_1681_));
 sg13g2_a21oi_1 _2529_ (.A1(_1680_),
    .A2(_1681_),
    .Y(_1682_),
    .B1(_1628_));
 sg13g2_nor2_1 _2530_ (.A(_1618_),
    .B(_1682_),
    .Y(_1683_));
 sg13g2_nand2_1 _2531_ (.Y(_1684_),
    .A(_1618_),
    .B(_1682_));
 sg13g2_nand2b_1 _2532_ (.Y(_1685_),
    .B(_1684_),
    .A_N(_1683_));
 sg13g2_xnor2_1 _2533_ (.Y(_1686_),
    .A(_1574_),
    .B(_1575_));
 sg13g2_nor2_1 _2534_ (.A(_1581_),
    .B(_1686_),
    .Y(_1687_));
 sg13g2_xor2_1 _2535_ (.B(_1686_),
    .A(_1581_),
    .X(_1688_));
 sg13g2_a21oi_1 _2536_ (.A1(_1607_),
    .A2(_1688_),
    .Y(_1689_),
    .B1(_1687_));
 sg13g2_xnor2_1 _2537_ (.Y(_1690_),
    .A(_1624_),
    .B(_1625_));
 sg13g2_nor2_1 _2538_ (.A(_1689_),
    .B(_1690_),
    .Y(_1691_));
 sg13g2_xor2_1 _2539_ (.B(_1690_),
    .A(_1689_),
    .X(_1692_));
 sg13g2_xnor2_1 _2540_ (.Y(_1693_),
    .A(_1677_),
    .B(_1679_));
 sg13g2_a21oi_1 _2541_ (.A1(_1692_),
    .A2(_1693_),
    .Y(_1694_),
    .B1(_1691_));
 sg13g2_xnor2_1 _2542_ (.Y(_1695_),
    .A(_1680_),
    .B(_1681_));
 sg13g2_nor2_1 _2543_ (.A(_1694_),
    .B(_1695_),
    .Y(_1696_));
 sg13g2_xor2_1 _2544_ (.B(_1676_),
    .A(_1675_),
    .X(_1697_));
 sg13g2_xnor2_1 _2545_ (.Y(_1698_),
    .A(_1606_),
    .B(_1688_));
 sg13g2_nand2_1 _2546_ (.Y(_1699_),
    .A(_1697_),
    .B(_1698_));
 sg13g2_xnor2_1 _2547_ (.Y(_1700_),
    .A(_1692_),
    .B(_1693_));
 sg13g2_or2_1 _2548_ (.X(_1701_),
    .B(_1700_),
    .A(_1699_));
 sg13g2_xnor2_1 _2549_ (.Y(_1702_),
    .A(_1568_),
    .B(_1570_));
 sg13g2_nor2_1 _2550_ (.A(_1558_),
    .B(_1702_),
    .Y(_1703_));
 sg13g2_xor2_1 _2551_ (.B(_1702_),
    .A(_1558_),
    .X(_1704_));
 sg13g2_a21oi_1 _2552_ (.A1(_1590_),
    .A2(_1704_),
    .Y(_1705_),
    .B1(_1703_));
 sg13g2_o21ai_1 _2553_ (.B1(_1571_),
    .Y(_1706_),
    .A1(_1564_),
    .A2(_1572_));
 sg13g2_nor2b_2 _2554_ (.A(_1573_),
    .B_N(_1706_),
    .Y(_1707_));
 sg13g2_nor2b_1 _2555_ (.A(_1705_),
    .B_N(_1707_),
    .Y(_1708_));
 sg13g2_xnor2_1 _2556_ (.Y(_1709_),
    .A(_1673_),
    .B(_1674_));
 sg13g2_xnor2_1 _2557_ (.Y(_1710_),
    .A(_1705_),
    .B(_1707_));
 sg13g2_nor2b_1 _2558_ (.A(_1709_),
    .B_N(_1710_),
    .Y(_1711_));
 sg13g2_nor2_1 _2559_ (.A(_1708_),
    .B(_1711_),
    .Y(_1712_));
 sg13g2_xnor2_1 _2560_ (.Y(_1713_),
    .A(_1697_),
    .B(_1698_));
 sg13g2_nor2_1 _2561_ (.A(_1712_),
    .B(_1713_),
    .Y(_1714_));
 sg13g2_xnor2_1 _2562_ (.Y(_1715_),
    .A(_1709_),
    .B(_1710_));
 sg13g2_xnor2_1 _2563_ (.Y(_1716_),
    .A(_1554_),
    .B(_1567_));
 sg13g2_xnor2_1 _2564_ (.Y(_1717_),
    .A(_1668_),
    .B(_1670_));
 sg13g2_nor2_1 _2565_ (.A(_1716_),
    .B(_1717_),
    .Y(_1718_));
 sg13g2_xnor2_1 _2566_ (.Y(_1719_),
    .A(net179),
    .B(_1704_));
 sg13g2_nand2_1 _2567_ (.Y(_1720_),
    .A(_1718_),
    .B(_1719_));
 sg13g2_xnor2_1 _2568_ (.Y(_1721_),
    .A(_1671_),
    .B(_1672_));
 sg13g2_inv_1 _2569_ (.Y(_1722_),
    .A(_1721_));
 sg13g2_xnor2_1 _2570_ (.Y(_1723_),
    .A(_1718_),
    .B(_1719_));
 sg13g2_o21ai_1 _2571_ (.B1(_1720_),
    .Y(_1724_),
    .A1(_1722_),
    .A2(_1723_));
 sg13g2_nand2_1 _2572_ (.Y(_1725_),
    .A(_1715_),
    .B(_1724_));
 sg13g2_xnor2_1 _2573_ (.Y(_1726_),
    .A(_1715_),
    .B(_1724_));
 sg13g2_xnor2_1 _2574_ (.Y(_1727_),
    .A(_1716_),
    .B(_1717_));
 sg13g2_inv_1 _2575_ (.Y(_1728_),
    .A(_1727_));
 sg13g2_xor2_1 _2576_ (.B(_1669_),
    .A(_1656_),
    .X(_1729_));
 sg13g2_and2_1 _2577_ (.A(_1566_),
    .B(_1729_),
    .X(_1730_));
 sg13g2_nand2_1 _2578_ (.Y(_1731_),
    .A(_1728_),
    .B(_1730_));
 sg13g2_xnor2_1 _2579_ (.Y(_1732_),
    .A(_1722_),
    .B(_1723_));
 sg13g2_or2_1 _2580_ (.X(_1733_),
    .B(_1732_),
    .A(_1731_));
 sg13g2_o21ai_1 _2581_ (.B1(_1725_),
    .Y(_1734_),
    .A1(_1726_),
    .A2(_1733_));
 sg13g2_xor2_1 _2582_ (.B(_1713_),
    .A(_1712_),
    .X(_1735_));
 sg13g2_nand2_1 _2583_ (.Y(_1736_),
    .A(_1734_),
    .B(_1735_));
 sg13g2_a21oi_1 _2584_ (.A1(_1734_),
    .A2(_1735_),
    .Y(_1737_),
    .B1(_1714_));
 sg13g2_xnor2_1 _2585_ (.Y(_1738_),
    .A(_1699_),
    .B(_1700_));
 sg13g2_nor2_1 _2586_ (.A(_1737_),
    .B(_1738_),
    .Y(_1739_));
 sg13g2_o21ai_1 _2587_ (.B1(_1701_),
    .Y(_1740_),
    .A1(_1737_),
    .A2(_1738_));
 sg13g2_nand2_1 _2588_ (.Y(_1741_),
    .A(_1694_),
    .B(_1695_));
 sg13g2_nand2b_1 _2589_ (.Y(_1742_),
    .B(_1741_),
    .A_N(_1696_));
 sg13g2_a21o_1 _2590_ (.A2(_1741_),
    .A1(_1740_),
    .B1(_1696_),
    .X(_1743_));
 sg13g2_a21oi_1 _2591_ (.A1(_1684_),
    .A2(_1743_),
    .Y(_1744_),
    .B1(_1683_));
 sg13g2_o21ai_1 _2592_ (.B1(_1523_),
    .Y(_1745_),
    .A1(_1528_),
    .A2(_1547_));
 sg13g2_o21ai_1 _2593_ (.B1(_1598_),
    .Y(_1746_),
    .A1(net180),
    .A2(_1603_));
 sg13g2_nor2_1 _2594_ (.A(_1745_),
    .B(_1746_),
    .Y(_1747_));
 sg13g2_xnor2_1 _2595_ (.Y(_1748_),
    .A(_1745_),
    .B(_1746_));
 sg13g2_inv_1 _2596_ (.Y(_1749_),
    .A(_1748_));
 sg13g2_xnor2_1 _2597_ (.Y(_1750_),
    .A(_1614_),
    .B(_1748_));
 sg13g2_nand2_1 _2598_ (.Y(_1751_),
    .A(_1617_),
    .B(_1750_));
 sg13g2_xnor2_1 _2599_ (.Y(_1752_),
    .A(_1617_),
    .B(_1750_));
 sg13g2_xor2_1 _2600_ (.B(_1752_),
    .A(_1744_),
    .X(_1753_));
 sg13g2_xnor2_1 _2601_ (.Y(_1754_),
    .A(_1685_),
    .B(_1743_));
 sg13g2_nor2_1 _2602_ (.A(_1734_),
    .B(_1735_),
    .Y(_1755_));
 sg13g2_a21oi_1 _2603_ (.A1(_1701_),
    .A2(_1742_),
    .Y(_1756_),
    .B1(_1739_));
 sg13g2_a21oi_1 _2604_ (.A1(_1737_),
    .A2(_1738_),
    .Y(_1757_),
    .B1(_1755_));
 sg13g2_and3_1 _2605_ (.X(_1758_),
    .A(_1736_),
    .B(_1756_),
    .C(_1757_));
 sg13g2_xor2_1 _2606_ (.B(_1730_),
    .A(_1727_),
    .X(_1759_));
 sg13g2_nor3_1 _2607_ (.A(_1726_),
    .B(_1732_),
    .C(_1759_),
    .Y(_1760_));
 sg13g2_a21oi_1 _2608_ (.A1(_1758_),
    .A2(_1760_),
    .Y(_1761_),
    .B1(_1754_));
 sg13g2_nand2b_1 _2609_ (.Y(_1762_),
    .B(_1761_),
    .A_N(_1753_));
 sg13g2_o21ai_1 _2610_ (.B1(_1751_),
    .Y(_1763_),
    .A1(_1744_),
    .A2(_1752_));
 sg13g2_a21oi_1 _2611_ (.A1(_1614_),
    .A2(_1749_),
    .Y(_1764_),
    .B1(_1747_));
 sg13g2_xnor2_1 _2612_ (.Y(_1765_),
    .A(_1579_),
    .B(_1599_));
 sg13g2_xnor2_1 _2613_ (.Y(_1766_),
    .A(_1764_),
    .B(_1765_));
 sg13g2_nor2_1 _2614_ (.A(_1566_),
    .B(_1729_),
    .Y(_1767_));
 sg13g2_nor3_1 _2615_ (.A(_1585_),
    .B(net179),
    .C(_1767_),
    .Y(_1768_));
 sg13g2_nor3_1 _2616_ (.A(_1728_),
    .B(_1730_),
    .C(_1768_),
    .Y(_1769_));
 sg13g2_nor2_1 _2617_ (.A(_1732_),
    .B(_1769_),
    .Y(_1770_));
 sg13g2_mux2_1 _2618_ (.A0(_1733_),
    .A1(_1770_),
    .S(_1726_),
    .X(_1771_));
 sg13g2_a21o_1 _2619_ (.A2(_1771_),
    .A1(_1758_),
    .B1(_1754_),
    .X(_1772_));
 sg13g2_a221oi_1 _2620_ (.B2(_1772_),
    .C1(_1501_),
    .B1(_1753_),
    .A1(_1453_),
    .Y(_1773_),
    .A2(_1486_));
 sg13g2_xnor2_1 _2621_ (.Y(_1774_),
    .A(_1763_),
    .B(_1766_));
 sg13g2_and3_2 _2622_ (.X(_1775_),
    .A(_1762_),
    .B(_1773_),
    .C(_1774_));
 sg13g2_nand3_1 _2623_ (.B(_1773_),
    .C(_1774_),
    .A(_1762_),
    .Y(_1776_));
 sg13g2_nor2_1 _2624_ (.A(_1413_),
    .B(_1425_),
    .Y(_1777_));
 sg13g2_nor2_1 _2625_ (.A(_1406_),
    .B(_1479_),
    .Y(_1778_));
 sg13g2_o21ai_1 _2626_ (.B1(_1777_),
    .Y(_1779_),
    .A1(_1504_),
    .A2(_1778_));
 sg13g2_nor2_1 _2627_ (.A(_1452_),
    .B(_1779_),
    .Y(_1780_));
 sg13g2_nor4_1 _2628_ (.A(_1337_),
    .B(_1485_),
    .C(_1490_),
    .D(_1780_),
    .Y(_1781_));
 sg13g2_nand2_1 _2629_ (.Y(_1782_),
    .A(_1453_),
    .B(_1781_));
 sg13g2_or3_1 _2630_ (.A(_1460_),
    .B(_1462_),
    .C(_1468_),
    .X(_1783_));
 sg13g2_a21oi_1 _2631_ (.A1(_1593_),
    .A2(_1783_),
    .Y(_1784_),
    .B1(_1338_));
 sg13g2_nand2_1 _2632_ (.Y(_1785_),
    .A(_1334_),
    .B(_1784_));
 sg13g2_nand3_1 _2633_ (.B(_1487_),
    .C(_1785_),
    .A(_1483_),
    .Y(_1786_));
 sg13g2_nand3_1 _2634_ (.B(_1438_),
    .C(_1481_),
    .A(_1428_),
    .Y(_1787_));
 sg13g2_a22oi_1 _2635_ (.Y(_1788_),
    .B1(_1787_),
    .B2(_1450_),
    .A2(_1786_),
    .A1(_1782_));
 sg13g2_nand2_1 _2636_ (.Y(_1789_),
    .A(_1460_),
    .B(_1467_));
 sg13g2_nand3_1 _2637_ (.B(_1471_),
    .C(_1789_),
    .A(_1458_),
    .Y(_1790_));
 sg13g2_a21oi_1 _2638_ (.A1(_1489_),
    .A2(_1790_),
    .Y(_1791_),
    .B1(_1335_));
 sg13g2_o21ai_1 _2639_ (.B1(_1335_),
    .Y(_1792_),
    .A1(_1457_),
    .A2(_1783_));
 sg13g2_nor3_1 _2640_ (.A(_1337_),
    .B(_1339_),
    .C(_1792_),
    .Y(_1793_));
 sg13g2_a221oi_1 _2641_ (.B2(_1429_),
    .C1(_1438_),
    .B1(_1492_),
    .A1(_1444_),
    .Y(_1794_),
    .A2(_1446_));
 sg13g2_nor4_1 _2642_ (.A(_1494_),
    .B(_1791_),
    .C(_1793_),
    .D(_1794_),
    .Y(_1795_));
 sg13g2_a21o_1 _2643_ (.A2(_1777_),
    .A1(_1491_),
    .B1(_1429_),
    .X(_1796_));
 sg13g2_a21oi_1 _2644_ (.A1(_1472_),
    .A2(_1796_),
    .Y(_1797_),
    .B1(_1794_));
 sg13g2_nand2_1 _2645_ (.Y(_1798_),
    .A(_1452_),
    .B(_1797_));
 sg13g2_nand3_1 _2646_ (.B(_1462_),
    .C(_1468_),
    .A(_1460_),
    .Y(_1799_));
 sg13g2_nand3_1 _2647_ (.B(_1458_),
    .C(_1799_),
    .A(_1339_),
    .Y(_1800_));
 sg13g2_nand2_1 _2648_ (.Y(_1801_),
    .A(_1337_),
    .B(_1800_));
 sg13g2_nor4_1 _2649_ (.A(_1334_),
    .B(_1593_),
    .C(_1798_),
    .D(_1801_),
    .Y(_1802_));
 sg13g2_nor3_2 _2650_ (.A(_1788_),
    .B(_1795_),
    .C(_1802_),
    .Y(_1803_));
 sg13g2_inv_2 _2651_ (.Y(_1804_),
    .A(net175));
 sg13g2_nand2_2 _2652_ (.Y(_1805_),
    .A(net172),
    .B(net175));
 sg13g2_nor2b_1 _2653_ (.A(\sin_y_acc[23] ),
    .B_N(\cos_x_acc[23] ),
    .Y(_1806_));
 sg13g2_nand2b_1 _2654_ (.Y(_1807_),
    .B(\sin_y_acc[23] ),
    .A_N(\cos_x_acc[23] ));
 sg13g2_nand2b_2 _2655_ (.Y(_1808_),
    .B(_1807_),
    .A_N(_1806_));
 sg13g2_o21ai_1 _2656_ (.B1(_1332_),
    .Y(_1809_),
    .A1(\sin_y_acc[22] ),
    .A2(_1236_));
 sg13g2_xnor2_1 _2657_ (.Y(_1810_),
    .A(_1808_),
    .B(_1809_));
 sg13g2_xor2_1 _2658_ (.B(_1809_),
    .A(_1808_),
    .X(_1811_));
 sg13g2_a21oi_1 _2659_ (.A1(net247),
    .A2(\sin_x_acc[22] ),
    .Y(_1812_),
    .B1(_1443_));
 sg13g2_xor2_1 _2660_ (.B(\sin_x_acc[23] ),
    .A(\cos_y_acc[23] ),
    .X(_1813_));
 sg13g2_xnor2_1 _2661_ (.Y(_1814_),
    .A(_1812_),
    .B(_1813_));
 sg13g2_xnor2_1 _2662_ (.Y(_1815_),
    .A(_1811_),
    .B(_1814_));
 sg13g2_xnor2_1 _2663_ (.Y(_1816_),
    .A(_1810_),
    .B(_1814_));
 sg13g2_nand3_1 _2664_ (.B(net175),
    .C(net178),
    .A(net172),
    .Y(_1817_));
 sg13g2_a21oi_1 _2665_ (.A1(_1291_),
    .A2(_1301_),
    .Y(_1818_),
    .B1(_1305_));
 sg13g2_nor2b_1 _2666_ (.A(_1818_),
    .B_N(_1296_),
    .Y(_1819_));
 sg13g2_xnor2_1 _2667_ (.Y(_1820_),
    .A(_1296_),
    .B(_1818_));
 sg13g2_xnor2_1 _2668_ (.Y(_1821_),
    .A(\sin_x_acc[10] ),
    .B(_1820_));
 sg13g2_and2_1 _2669_ (.A(_1200_),
    .B(_1821_),
    .X(_1822_));
 sg13g2_a21o_1 _2670_ (.A2(_1820_),
    .A1(_1226_),
    .B1(_1822_),
    .X(_1823_));
 sg13g2_nor2_1 _2671_ (.A(_1295_),
    .B(_1819_),
    .Y(_1824_));
 sg13g2_xor2_1 _2672_ (.B(_1824_),
    .A(_1294_),
    .X(_1825_));
 sg13g2_nor2b_1 _2673_ (.A(_1377_),
    .B_N(_1382_),
    .Y(_1826_));
 sg13g2_xnor2_1 _2674_ (.Y(_1827_),
    .A(_1825_),
    .B(_1826_));
 sg13g2_nand2_1 _2675_ (.Y(_1828_),
    .A(_1823_),
    .B(_1827_));
 sg13g2_xnor2_1 _2676_ (.Y(_1829_),
    .A(\cos_y_acc[10] ),
    .B(_1821_));
 sg13g2_a21oi_1 _2677_ (.A1(_1291_),
    .A2(_1299_),
    .Y(_1830_),
    .B1(_1298_));
 sg13g2_xnor2_1 _2678_ (.Y(_1831_),
    .A(_1300_),
    .B(_1830_));
 sg13g2_a21oi_1 _2679_ (.A1(_1379_),
    .A2(_1831_),
    .Y(_1832_),
    .B1(_1385_));
 sg13g2_nor2b_1 _2680_ (.A(_1832_),
    .B_N(_1829_),
    .Y(_1833_));
 sg13g2_xor2_1 _2681_ (.B(_1832_),
    .A(_1829_),
    .X(_1834_));
 sg13g2_xor2_1 _2682_ (.B(_1299_),
    .A(_1291_),
    .X(_1835_));
 sg13g2_nor2b_1 _2683_ (.A(\sin_x_acc[8] ),
    .B_N(_1835_),
    .Y(_1836_));
 sg13g2_xnor2_1 _2684_ (.Y(_1837_),
    .A(\sin_x_acc[8] ),
    .B(_1835_));
 sg13g2_and2_1 _2685_ (.A(_1202_),
    .B(_1837_),
    .X(_1838_));
 sg13g2_xnor2_1 _2686_ (.Y(_1839_),
    .A(\cos_y_acc[9] ),
    .B(\sin_x_acc[9] ));
 sg13g2_xnor2_1 _2687_ (.Y(_1840_),
    .A(_1831_),
    .B(_1839_));
 sg13g2_or3_1 _2688_ (.A(_1836_),
    .B(_1838_),
    .C(_1840_),
    .X(_1841_));
 sg13g2_o21ai_1 _2689_ (.B1(_1840_),
    .Y(_1842_),
    .A1(_1836_),
    .A2(_1838_));
 sg13g2_xnor2_1 _2690_ (.Y(_1843_),
    .A(_1202_),
    .B(_1837_));
 sg13g2_xor2_1 _2691_ (.B(_1290_),
    .A(_1289_),
    .X(_1844_));
 sg13g2_xnor2_1 _2692_ (.Y(_1845_),
    .A(\sin_x_acc[7] ),
    .B(_1844_));
 sg13g2_and2_1 _2693_ (.A(_1203_),
    .B(_1845_),
    .X(_1846_));
 sg13g2_a21oi_1 _2694_ (.A1(_1225_),
    .A2(_1844_),
    .Y(_1847_),
    .B1(_1846_));
 sg13g2_nor2_1 _2695_ (.A(_1843_),
    .B(_1847_),
    .Y(_1848_));
 sg13g2_xnor2_1 _2696_ (.Y(_1849_),
    .A(_1270_),
    .B(_1288_));
 sg13g2_nand2b_1 _2697_ (.Y(_1850_),
    .B(_1849_),
    .A_N(\sin_x_acc[6] ));
 sg13g2_xnor2_1 _2698_ (.Y(_1851_),
    .A(\sin_x_acc[6] ),
    .B(_1849_));
 sg13g2_nand2b_1 _2699_ (.Y(_1852_),
    .B(_1851_),
    .A_N(\cos_y_acc[6] ));
 sg13g2_nand2_1 _2700_ (.Y(_1853_),
    .A(_1850_),
    .B(_1852_));
 sg13g2_xnor2_1 _2701_ (.Y(_1854_),
    .A(\cos_y_acc[7] ),
    .B(_1845_));
 sg13g2_nor2_1 _2702_ (.A(_1853_),
    .B(_1854_),
    .Y(_1855_));
 sg13g2_xor2_1 _2703_ (.B(_1283_),
    .A(_1281_),
    .X(_1856_));
 sg13g2_xnor2_1 _2704_ (.Y(_1857_),
    .A(\sin_x_acc[4] ),
    .B(_1856_));
 sg13g2_and2_1 _2705_ (.A(_1205_),
    .B(_1857_),
    .X(_1858_));
 sg13g2_a21oi_1 _2706_ (.A1(_1224_),
    .A2(_1856_),
    .Y(_1859_),
    .B1(_1858_));
 sg13g2_a21oi_1 _2707_ (.A1(_1281_),
    .A2(_1283_),
    .Y(_1860_),
    .B1(_1282_));
 sg13g2_xor2_1 _2708_ (.B(_1860_),
    .A(_1286_),
    .X(_1861_));
 sg13g2_nor2_1 _2709_ (.A(\sin_x_acc[5] ),
    .B(_1861_),
    .Y(_1862_));
 sg13g2_xor2_1 _2710_ (.B(_1861_),
    .A(\sin_x_acc[5] ),
    .X(_1863_));
 sg13g2_xnor2_1 _2711_ (.Y(_1864_),
    .A(_1204_),
    .B(_1863_));
 sg13g2_nor2_1 _2712_ (.A(_1859_),
    .B(_1864_),
    .Y(_1865_));
 sg13g2_xor2_1 _2713_ (.B(_1280_),
    .A(_1279_),
    .X(_1866_));
 sg13g2_xnor2_1 _2714_ (.Y(_1867_),
    .A(\sin_x_acc[3] ),
    .B(_1866_));
 sg13g2_and2_1 _2715_ (.A(_1206_),
    .B(_1867_),
    .X(_1868_));
 sg13g2_a21o_1 _2716_ (.A2(_1866_),
    .A1(_1213_),
    .B1(_1868_),
    .X(_1869_));
 sg13g2_xnor2_1 _2717_ (.Y(_1870_),
    .A(\cos_y_acc[4] ),
    .B(_1857_));
 sg13g2_nand2_1 _2718_ (.Y(_1871_),
    .A(_1869_),
    .B(_1870_));
 sg13g2_nor2_1 _2719_ (.A(_1869_),
    .B(_1870_),
    .Y(_1872_));
 sg13g2_xnor2_1 _2720_ (.Y(_1873_),
    .A(_1276_),
    .B(_1278_));
 sg13g2_nand2b_1 _2721_ (.Y(_1874_),
    .B(_1873_),
    .A_N(\sin_x_acc[2] ));
 sg13g2_xnor2_1 _2722_ (.Y(_1875_),
    .A(\sin_x_acc[2] ),
    .B(_1873_));
 sg13g2_nand2b_1 _2723_ (.Y(_1876_),
    .B(_1875_),
    .A_N(\cos_y_acc[2] ));
 sg13g2_and2_1 _2724_ (.A(_1874_),
    .B(_1876_),
    .X(_1877_));
 sg13g2_xnor2_1 _2725_ (.Y(_1878_),
    .A(_1206_),
    .B(_1867_));
 sg13g2_nor2_1 _2726_ (.A(_1877_),
    .B(_1878_),
    .Y(_1879_));
 sg13g2_nand2b_1 _2727_ (.Y(_1880_),
    .B(\cos_y_acc[2] ),
    .A_N(_1875_));
 sg13g2_xnor2_1 _2728_ (.Y(_1881_),
    .A(_1274_),
    .B(_1275_));
 sg13g2_nor2b_1 _2729_ (.A(\sin_y_acc[0] ),
    .B_N(\cos_x_acc[0] ),
    .Y(_1882_));
 sg13g2_o21ai_1 _2730_ (.B1(_1274_),
    .Y(_1883_),
    .A1(\cos_y_acc[0] ),
    .A2(\sin_x_acc[0] ));
 sg13g2_o21ai_1 _2731_ (.B1(_1359_),
    .Y(_1884_),
    .A1(_1882_),
    .A2(_1883_));
 sg13g2_nand2_1 _2732_ (.Y(_1885_),
    .A(_1881_),
    .B(_1884_));
 sg13g2_nand3_1 _2733_ (.B(_1881_),
    .C(_1884_),
    .A(_1358_),
    .Y(_1886_));
 sg13g2_nand3_1 _2734_ (.B(_1880_),
    .C(_1886_),
    .A(_1876_),
    .Y(_1887_));
 sg13g2_nor3_1 _2735_ (.A(_1358_),
    .B(_1881_),
    .C(_1884_),
    .Y(_1888_));
 sg13g2_a21oi_1 _2736_ (.A1(_1361_),
    .A2(_1885_),
    .Y(_1889_),
    .B1(_1888_));
 sg13g2_a22oi_1 _2737_ (.Y(_1890_),
    .B1(_1887_),
    .B2(_1889_),
    .A2(_1878_),
    .A1(_1877_));
 sg13g2_nor2_1 _2738_ (.A(_1879_),
    .B(_1890_),
    .Y(_1891_));
 sg13g2_o21ai_1 _2739_ (.B1(_1871_),
    .Y(_1892_),
    .A1(_1872_),
    .A2(_1891_));
 sg13g2_xor2_1 _2740_ (.B(_1851_),
    .A(\cos_y_acc[6] ),
    .X(_0147_));
 sg13g2_a21oi_1 _2741_ (.A1(_1204_),
    .A2(_1863_),
    .Y(_0148_),
    .B1(_1862_));
 sg13g2_a22oi_1 _2742_ (.Y(_0149_),
    .B1(_0147_),
    .B2(_0148_),
    .A2(_1864_),
    .A1(_1859_));
 sg13g2_o21ai_1 _2743_ (.B1(_0149_),
    .Y(_0150_),
    .A1(_1865_),
    .A2(_1892_));
 sg13g2_nor2_1 _2744_ (.A(_0147_),
    .B(_0148_),
    .Y(_0151_));
 sg13g2_a21oi_1 _2745_ (.A1(_1853_),
    .A2(_1854_),
    .Y(_0152_),
    .B1(_0151_));
 sg13g2_a221oi_1 _2746_ (.B2(_0152_),
    .C1(_1855_),
    .B1(_0150_),
    .A1(_1843_),
    .Y(_0153_),
    .A2(_1847_));
 sg13g2_nor2_1 _2747_ (.A(_1848_),
    .B(_0153_),
    .Y(_0154_));
 sg13g2_o21ai_1 _2748_ (.B1(_1841_),
    .Y(_0155_),
    .A1(_1848_),
    .A2(_0153_));
 sg13g2_nand2_1 _2749_ (.Y(_0156_),
    .A(_1842_),
    .B(_0155_));
 sg13g2_a21oi_1 _2750_ (.A1(_1842_),
    .A2(_0155_),
    .Y(_0157_),
    .B1(_1834_));
 sg13g2_nor2_1 _2751_ (.A(_1833_),
    .B(_0157_),
    .Y(_0158_));
 sg13g2_xor2_1 _2752_ (.B(_1827_),
    .A(_1823_),
    .X(_0159_));
 sg13g2_o21ai_1 _2753_ (.B1(_0159_),
    .Y(_0160_),
    .A1(_1833_),
    .A2(_0157_));
 sg13g2_nor2_1 _2754_ (.A(_1262_),
    .B(_1308_),
    .Y(_0161_));
 sg13g2_xor2_1 _2755_ (.B(_1308_),
    .A(_1262_),
    .X(_0162_));
 sg13g2_and2_1 _2756_ (.A(_1227_),
    .B(_0162_),
    .X(_0163_));
 sg13g2_xnor2_1 _2757_ (.Y(_0164_),
    .A(\sin_x_acc[12] ),
    .B(_0162_));
 sg13g2_and2_1 _2758_ (.A(_1198_),
    .B(_0164_),
    .X(_0165_));
 sg13g2_xnor2_1 _2759_ (.Y(_0166_),
    .A(\cos_y_acc[12] ),
    .B(_0164_));
 sg13g2_a21oi_1 _2760_ (.A1(_1382_),
    .A2(_1825_),
    .Y(_0167_),
    .B1(_1377_));
 sg13g2_and2_1 _2761_ (.A(_0166_),
    .B(_0167_),
    .X(_0168_));
 sg13g2_inv_1 _2762_ (.Y(_0169_),
    .A(_0168_));
 sg13g2_xnor2_1 _2763_ (.Y(_0170_),
    .A(_0166_),
    .B(_0167_));
 sg13g2_a21o_2 _2764_ (.A2(_0160_),
    .A1(_1828_),
    .B1(_0170_),
    .X(_0171_));
 sg13g2_nand3_1 _2765_ (.B(_0160_),
    .C(_0170_),
    .A(_1828_),
    .Y(_0172_));
 sg13g2_nand2_2 _2766_ (.Y(_0173_),
    .A(_0171_),
    .B(_0172_));
 sg13g2_xor2_1 _2767_ (.B(_0156_),
    .A(_1834_),
    .X(_0174_));
 sg13g2_xnor2_1 _2768_ (.Y(_0175_),
    .A(_0173_),
    .B(_0174_));
 sg13g2_nor2_1 _2769_ (.A(_1817_),
    .B(_0175_),
    .Y(_0176_));
 sg13g2_or4_1 _2770_ (.A(net173),
    .B(net174),
    .C(net176),
    .D(_0175_),
    .X(_0177_));
 sg13g2_xnor2_1 _2771_ (.Y(_0178_),
    .A(net251),
    .B(\hvsync_gen.hpos[1] ));
 sg13g2_xnor2_1 _2772_ (.Y(_0179_),
    .A(_1216_),
    .B(net245));
 sg13g2_nor2_1 _2773_ (.A(_0177_),
    .B(_0179_),
    .Y(_0180_));
 sg13g2_xnor2_1 _2774_ (.Y(_0181_),
    .A(_0158_),
    .B(_0159_));
 sg13g2_nand2_1 _2775_ (.Y(_0182_),
    .A(_0169_),
    .B(_0171_));
 sg13g2_nor2_1 _2776_ (.A(_1257_),
    .B(_0161_),
    .Y(_0183_));
 sg13g2_xnor2_1 _2777_ (.Y(_0184_),
    .A(_1263_),
    .B(_0183_));
 sg13g2_xnor2_1 _2778_ (.Y(_0185_),
    .A(_1355_),
    .B(_0184_));
 sg13g2_o21ai_1 _2779_ (.B1(_0185_),
    .Y(_0186_),
    .A1(_0163_),
    .A2(_0165_));
 sg13g2_inv_1 _2780_ (.Y(_0187_),
    .A(_0186_));
 sg13g2_nor3_1 _2781_ (.A(_0163_),
    .B(_0165_),
    .C(_0185_),
    .Y(_0188_));
 sg13g2_nor2_1 _2782_ (.A(_0187_),
    .B(_0188_),
    .Y(_0189_));
 sg13g2_xor2_1 _2783_ (.B(_0189_),
    .A(_0182_),
    .X(_0190_));
 sg13g2_xnor2_1 _2784_ (.Y(_0191_),
    .A(_0181_),
    .B(_0190_));
 sg13g2_nor4_2 _2785_ (.A(net173),
    .B(net174),
    .C(net176),
    .Y(_0192_),
    .D(_0191_));
 sg13g2_nand2_1 _2786_ (.Y(_0193_),
    .A(_0177_),
    .B(_0179_));
 sg13g2_xnor2_1 _2787_ (.Y(_0194_),
    .A(_0177_),
    .B(_0179_));
 sg13g2_a21oi_1 _2788_ (.A1(_0192_),
    .A2(_0193_),
    .Y(_0195_),
    .B1(_0180_));
 sg13g2_a21o_1 _2789_ (.A2(_0193_),
    .A1(_0192_),
    .B1(_0180_),
    .X(_0196_));
 sg13g2_xnor2_1 _2790_ (.Y(_0197_),
    .A(_1214_),
    .B(net182));
 sg13g2_nand2_1 _2791_ (.Y(_0198_),
    .A(_1197_),
    .B(_0197_));
 sg13g2_xnor2_1 _2792_ (.Y(_0199_),
    .A(\cos_y_acc[14] ),
    .B(_0197_));
 sg13g2_or2_1 _2793_ (.X(_0200_),
    .B(_0184_),
    .A(_1350_));
 sg13g2_nand2_1 _2794_ (.Y(_0201_),
    .A(_1347_),
    .B(_0200_));
 sg13g2_nand3_1 _2795_ (.B(_0199_),
    .C(_0200_),
    .A(_1347_),
    .Y(_0202_));
 sg13g2_xor2_1 _2796_ (.B(_0201_),
    .A(_0199_),
    .X(_0203_));
 sg13g2_inv_1 _2797_ (.Y(_0204_),
    .A(_0203_));
 sg13g2_a21oi_1 _2798_ (.A1(_0169_),
    .A2(_0171_),
    .Y(_0205_),
    .B1(_0188_));
 sg13g2_or2_1 _2799_ (.X(_0206_),
    .B(_0205_),
    .A(_0187_));
 sg13g2_o21ai_1 _2800_ (.B1(_0204_),
    .Y(_0207_),
    .A1(_0187_),
    .A2(_0205_));
 sg13g2_xnor2_1 _2801_ (.Y(_0208_),
    .A(_0203_),
    .B(_0206_));
 sg13g2_xnor2_1 _2802_ (.Y(_0209_),
    .A(_0173_),
    .B(_0208_));
 sg13g2_nor3_1 _2803_ (.A(net173),
    .B(net174),
    .C(_0209_),
    .Y(_0210_));
 sg13g2_nand3b_1 _2804_ (.B(net172),
    .C(net175),
    .Y(_0211_),
    .A_N(_0209_));
 sg13g2_nand2_2 _2805_ (.Y(_0212_),
    .A(net178),
    .B(_0211_));
 sg13g2_xnor2_1 _2806_ (.Y(_0213_),
    .A(net251),
    .B(\hvsync_gen.hpos[0] ));
 sg13g2_inv_4 _2807_ (.A(_0213_),
    .Y(_0214_));
 sg13g2_nand2_1 _2808_ (.Y(_0215_),
    .A(_0192_),
    .B(_0214_));
 sg13g2_xnor2_1 _2809_ (.Y(_0216_),
    .A(_0192_),
    .B(_0214_));
 sg13g2_xor2_1 _2810_ (.B(_0216_),
    .A(_0212_),
    .X(_0217_));
 sg13g2_xnor2_1 _2811_ (.Y(_0218_),
    .A(_0212_),
    .B(_0216_));
 sg13g2_nor4_1 _2812_ (.A(net173),
    .B(net174),
    .C(net176),
    .D(_0174_),
    .Y(_0219_));
 sg13g2_nor2b_1 _2813_ (.A(net245),
    .B_N(_0219_),
    .Y(_0220_));
 sg13g2_nand2_1 _2814_ (.Y(_0221_),
    .A(_1841_),
    .B(_1842_));
 sg13g2_xnor2_1 _2815_ (.Y(_0222_),
    .A(_0154_),
    .B(_0221_));
 sg13g2_xor2_1 _2816_ (.B(_0222_),
    .A(_0181_),
    .X(_0223_));
 sg13g2_nor2_1 _2817_ (.A(_1817_),
    .B(_0223_),
    .Y(_0224_));
 sg13g2_or2_1 _2818_ (.X(_0225_),
    .B(_0223_),
    .A(_1817_));
 sg13g2_o21ai_1 _2819_ (.B1(net245),
    .Y(_0226_),
    .A1(_1817_),
    .A2(_0174_));
 sg13g2_xnor2_1 _2820_ (.Y(_0227_),
    .A(net245),
    .B(_0219_));
 sg13g2_a21oi_1 _2821_ (.A1(_0224_),
    .A2(_0226_),
    .Y(_0228_),
    .B1(_0220_));
 sg13g2_a21o_1 _2822_ (.A2(_0226_),
    .A1(_0224_),
    .B1(_0220_),
    .X(_0229_));
 sg13g2_xnor2_1 _2823_ (.Y(_0230_),
    .A(_0192_),
    .B(_0194_));
 sg13g2_xor2_1 _2824_ (.B(_0194_),
    .A(_0192_),
    .X(_0231_));
 sg13g2_a22oi_1 _2825_ (.Y(_0232_),
    .B1(_0229_),
    .B2(_0230_),
    .A2(_0217_),
    .A1(_0196_));
 sg13g2_nor2_1 _2826_ (.A(_0196_),
    .B(_0217_),
    .Y(_0233_));
 sg13g2_o21ai_1 _2827_ (.B1(_0198_),
    .Y(_0234_),
    .A1(\sin_x_acc[14] ),
    .A2(net182));
 sg13g2_or2_1 _2828_ (.X(_0235_),
    .B(_1467_),
    .A(\sin_x_acc[15] ));
 sg13g2_xnor2_1 _2829_ (.Y(_0236_),
    .A(\sin_x_acc[15] ),
    .B(_1467_));
 sg13g2_xor2_1 _2830_ (.B(_0236_),
    .A(\cos_y_acc[15] ),
    .X(_0237_));
 sg13g2_xor2_1 _2831_ (.B(_0237_),
    .A(_0234_),
    .X(_0238_));
 sg13g2_inv_1 _2832_ (.Y(_0239_),
    .A(_0238_));
 sg13g2_a21oi_1 _2833_ (.A1(_0202_),
    .A2(_0207_),
    .Y(_0240_),
    .B1(_0239_));
 sg13g2_nand3_1 _2834_ (.B(_0207_),
    .C(_0239_),
    .A(_0202_),
    .Y(_0241_));
 sg13g2_nand2b_2 _2835_ (.Y(_0242_),
    .B(_0241_),
    .A_N(_0240_));
 sg13g2_xor2_1 _2836_ (.B(_0242_),
    .A(_0190_),
    .X(_0243_));
 sg13g2_nand3_1 _2837_ (.B(net175),
    .C(_0243_),
    .A(net172),
    .Y(_0244_));
 sg13g2_and2_1 _2838_ (.A(net178),
    .B(_0244_),
    .X(_0245_));
 sg13g2_xnor2_1 _2839_ (.Y(_0246_),
    .A(net251),
    .B(\hvsync_gen.hpos[2] ));
 sg13g2_xor2_1 _2840_ (.B(\hvsync_gen.hpos[2] ),
    .A(net251),
    .X(_0247_));
 sg13g2_a21oi_1 _2841_ (.A1(net178),
    .A2(_0244_),
    .Y(_0248_),
    .B1(_0247_));
 sg13g2_nand3_1 _2842_ (.B(_0244_),
    .C(_0247_),
    .A(net178),
    .Y(_0249_));
 sg13g2_o21ai_1 _2843_ (.B1(_0249_),
    .Y(_0250_),
    .A1(_0225_),
    .A2(_0248_));
 sg13g2_or2_1 _2844_ (.X(_0251_),
    .B(_0250_),
    .A(_0176_));
 sg13g2_xnor2_1 _2845_ (.Y(_0252_),
    .A(_0225_),
    .B(_0227_));
 sg13g2_a21o_1 _2846_ (.A2(_0250_),
    .A1(_0176_),
    .B1(_0252_),
    .X(_0253_));
 sg13g2_a22oi_1 _2847_ (.Y(_0254_),
    .B1(_0228_),
    .B2(_0231_),
    .A2(_0218_),
    .A1(_0195_));
 sg13g2_and4_1 _2848_ (.A(_0232_),
    .B(_0251_),
    .C(_0253_),
    .D(_0254_),
    .X(_0255_));
 sg13g2_o21ai_1 _2849_ (.B1(_0215_),
    .Y(_0256_),
    .A1(_0212_),
    .A2(_0216_));
 sg13g2_xnor2_1 _2850_ (.Y(_0257_),
    .A(_1215_),
    .B(_0213_));
 sg13g2_inv_2 _2851_ (.Y(_0258_),
    .A(_0257_));
 sg13g2_o21ai_1 _2852_ (.B1(_0257_),
    .Y(_0259_),
    .A1(net176),
    .A2(_0210_));
 sg13g2_nor3_1 _2853_ (.A(net177),
    .B(_0210_),
    .C(_0257_),
    .Y(_0260_));
 sg13g2_nand3_1 _2854_ (.B(_0211_),
    .C(_0258_),
    .A(_1815_),
    .Y(_0261_));
 sg13g2_a21o_1 _2855_ (.A2(_0261_),
    .A1(_0259_),
    .B1(_0245_),
    .X(_0262_));
 sg13g2_nand3b_1 _2856_ (.B(_0245_),
    .C(_0259_),
    .Y(_0263_),
    .A_N(_0260_));
 sg13g2_nand3_1 _2857_ (.B(_0262_),
    .C(_0263_),
    .A(_0256_),
    .Y(_0264_));
 sg13g2_o21ai_1 _2858_ (.B1(_0264_),
    .Y(_0265_),
    .A1(_0232_),
    .A2(_0233_));
 sg13g2_a21o_1 _2859_ (.A2(_0263_),
    .A1(_0262_),
    .B1(_0256_),
    .X(_0266_));
 sg13g2_o21ai_1 _2860_ (.B1(_0266_),
    .Y(_0267_),
    .A1(_0255_),
    .A2(_0265_));
 sg13g2_nand2_1 _2861_ (.Y(_0268_),
    .A(_0245_),
    .B(_0259_));
 sg13g2_o21ai_1 _2862_ (.B1(_0268_),
    .Y(_0269_),
    .A1(_0245_),
    .A2(_0260_));
 sg13g2_or2_1 _2863_ (.X(_0270_),
    .B(_0269_),
    .A(_0267_));
 sg13g2_nor2_1 _2864_ (.A(\hvsync_gen.hpos[8] ),
    .B(\hvsync_gen.hpos[7] ),
    .Y(_0271_));
 sg13g2_o21ai_1 _2865_ (.B1(\hvsync_gen.hpos[9] ),
    .Y(_0272_),
    .A1(\hvsync_gen.hpos[8] ),
    .A2(\hvsync_gen.hpos[7] ));
 sg13g2_nand2_1 _2866_ (.Y(_0273_),
    .A(net297),
    .B(net322));
 sg13g2_nand4_1 _2867_ (.B(\hvsync_gen.vpos[6] ),
    .C(\hvsync_gen.vpos[7] ),
    .A(\hvsync_gen.vpos[5] ),
    .Y(_0274_),
    .D(\hvsync_gen.vpos[8] ));
 sg13g2_nand3b_1 _2868_ (.B(_0272_),
    .C(_0274_),
    .Y(_0275_),
    .A_N(\hvsync_gen.vpos[9] ));
 sg13g2_a21oi_1 _2869_ (.A1(_0267_),
    .A2(_0269_),
    .Y(_0276_),
    .B1(_0275_));
 sg13g2_and2_1 _2870_ (.A(_0270_),
    .B(_0276_),
    .X(uo_out[6]));
 sg13g2_a21oi_2 _2871_ (.B1(_0275_),
    .Y(uo_out[2]),
    .A2(_0270_),
    .A1(_0268_));
 sg13g2_xnor2_1 _2872_ (.Y(_0277_),
    .A(\sin_x_acc[19] ),
    .B(_1457_));
 sg13g2_nor2_1 _2873_ (.A(\cos_y_acc[19] ),
    .B(_0277_),
    .Y(_0278_));
 sg13g2_a21oi_1 _2874_ (.A1(_1218_),
    .A2(_1458_),
    .Y(_0279_),
    .B1(_0278_));
 sg13g2_xnor2_1 _2875_ (.Y(_0280_),
    .A(\sin_x_acc[20] ),
    .B(_1339_));
 sg13g2_nand2b_1 _2876_ (.Y(_0281_),
    .B(_0280_),
    .A_N(net248));
 sg13g2_xnor2_1 _2877_ (.Y(_0282_),
    .A(net248),
    .B(_0280_));
 sg13g2_nand2b_1 _2878_ (.Y(_0283_),
    .B(_0282_),
    .A_N(_0279_));
 sg13g2_xnor2_1 _2879_ (.Y(_0284_),
    .A(_0279_),
    .B(_0282_));
 sg13g2_xnor2_1 _2880_ (.Y(_0285_),
    .A(\sin_x_acc[18] ),
    .B(_1459_));
 sg13g2_nor2b_1 _2881_ (.A(\cos_y_acc[18] ),
    .B_N(_0285_),
    .Y(_0286_));
 sg13g2_a21oi_1 _2882_ (.A1(_1219_),
    .A2(_1459_),
    .Y(_0287_),
    .B1(_0286_));
 sg13g2_xnor2_1 _2883_ (.Y(_0288_),
    .A(_1194_),
    .B(_0277_));
 sg13g2_nand2b_1 _2884_ (.Y(_0289_),
    .B(_0287_),
    .A_N(_0288_));
 sg13g2_nand2b_1 _2885_ (.Y(_0290_),
    .B(_0288_),
    .A_N(_0287_));
 sg13g2_nor2_1 _2886_ (.A(\sin_x_acc[17] ),
    .B(_1462_),
    .Y(_0291_));
 sg13g2_xnor2_1 _2887_ (.Y(_0292_),
    .A(_1220_),
    .B(_1462_));
 sg13g2_a21oi_1 _2888_ (.A1(_1195_),
    .A2(_0292_),
    .Y(_0293_),
    .B1(_0291_));
 sg13g2_xnor2_1 _2889_ (.Y(_0294_),
    .A(\cos_y_acc[18] ),
    .B(_0285_));
 sg13g2_nand2b_1 _2890_ (.Y(_0295_),
    .B(_0294_),
    .A_N(_0293_));
 sg13g2_xnor2_1 _2891_ (.Y(_0296_),
    .A(_0293_),
    .B(_0294_));
 sg13g2_nor2_1 _2892_ (.A(\sin_x_acc[16] ),
    .B(_1464_),
    .Y(_0297_));
 sg13g2_xnor2_1 _2893_ (.Y(_0298_),
    .A(\sin_x_acc[16] ),
    .B(_1463_));
 sg13g2_a21oi_1 _2894_ (.A1(_1196_),
    .A2(_0298_),
    .Y(_0299_),
    .B1(_0297_));
 sg13g2_xnor2_1 _2895_ (.Y(_0300_),
    .A(\cos_y_acc[17] ),
    .B(_0292_));
 sg13g2_nor2b_1 _2896_ (.A(_0299_),
    .B_N(_0300_),
    .Y(_0301_));
 sg13g2_o21ai_1 _2897_ (.B1(_0235_),
    .Y(_0302_),
    .A1(\cos_y_acc[15] ),
    .A2(_0236_));
 sg13g2_xnor2_1 _2898_ (.Y(_0303_),
    .A(\cos_y_acc[16] ),
    .B(_0298_));
 sg13g2_nand2_1 _2899_ (.Y(_0304_),
    .A(_0302_),
    .B(_0303_));
 sg13g2_a21o_1 _2900_ (.A2(_0237_),
    .A1(_0234_),
    .B1(_0240_),
    .X(_0305_));
 sg13g2_xnor2_1 _2901_ (.Y(_0306_),
    .A(_0302_),
    .B(_0303_));
 sg13g2_inv_1 _2902_ (.Y(_0307_),
    .A(_0306_));
 sg13g2_nand2_1 _2903_ (.Y(_0308_),
    .A(_0305_),
    .B(_0307_));
 sg13g2_xor2_1 _2904_ (.B(_0300_),
    .A(_0299_),
    .X(_0309_));
 sg13g2_a21oi_1 _2905_ (.A1(_0304_),
    .A2(_0308_),
    .Y(_0310_),
    .B1(_0309_));
 sg13g2_nor2_1 _2906_ (.A(_0301_),
    .B(_0310_),
    .Y(_0311_));
 sg13g2_o21ai_1 _2907_ (.B1(_0296_),
    .Y(_0312_),
    .A1(_0301_),
    .A2(_0310_));
 sg13g2_nand2_1 _2908_ (.Y(_0313_),
    .A(_0295_),
    .B(_0312_));
 sg13g2_nand3_1 _2909_ (.B(_0295_),
    .C(_0312_),
    .A(_0290_),
    .Y(_0314_));
 sg13g2_nand3_1 _2910_ (.B(_0289_),
    .C(_0314_),
    .A(_0284_),
    .Y(_0315_));
 sg13g2_o21ai_1 _2911_ (.B1(_0281_),
    .Y(_0316_),
    .A1(\sin_x_acc[20] ),
    .A2(_1340_));
 sg13g2_nor2_1 _2912_ (.A(\sin_x_acc[21] ),
    .B(_1338_),
    .Y(_0317_));
 sg13g2_xnor2_1 _2913_ (.Y(_0318_),
    .A(\sin_x_acc[21] ),
    .B(_1337_));
 sg13g2_xnor2_1 _2914_ (.Y(_0319_),
    .A(\cos_y_acc[21] ),
    .B(_0318_));
 sg13g2_and2_1 _2915_ (.A(_0316_),
    .B(_0319_),
    .X(_0320_));
 sg13g2_xor2_1 _2916_ (.B(_0319_),
    .A(_0316_),
    .X(_0321_));
 sg13g2_inv_1 _2917_ (.Y(_0322_),
    .A(_0321_));
 sg13g2_a21oi_1 _2918_ (.A1(_0283_),
    .A2(_0315_),
    .Y(_0323_),
    .B1(_0322_));
 sg13g2_nand3_1 _2919_ (.B(_0315_),
    .C(_0322_),
    .A(_0283_),
    .Y(_0324_));
 sg13g2_nand2b_2 _2920_ (.Y(_0325_),
    .B(_0324_),
    .A_N(_0323_));
 sg13g2_and2_1 _2921_ (.A(_0289_),
    .B(_0290_),
    .X(_0326_));
 sg13g2_xnor2_1 _2922_ (.Y(_0327_),
    .A(_0313_),
    .B(_0326_));
 sg13g2_o21ai_1 _2923_ (.B1(net178),
    .Y(_0328_),
    .A1(_0325_),
    .A2(_0327_));
 sg13g2_a21oi_1 _2924_ (.A1(_0325_),
    .A2(_0327_),
    .Y(_0329_),
    .B1(_0328_));
 sg13g2_inv_1 _2925_ (.Y(_0330_),
    .A(_0329_));
 sg13g2_nand3_1 _2926_ (.B(net175),
    .C(_0330_),
    .A(net172),
    .Y(_0331_));
 sg13g2_inv_1 _2927_ (.Y(_0332_),
    .A(_0331_));
 sg13g2_xnor2_1 _2928_ (.Y(_0333_),
    .A(_0296_),
    .B(_0311_));
 sg13g2_a21o_1 _2929_ (.A2(_0314_),
    .A1(_0289_),
    .B1(_0284_),
    .X(_0334_));
 sg13g2_nand2_1 _2930_ (.Y(_0335_),
    .A(_0315_),
    .B(_0334_));
 sg13g2_xnor2_1 _2931_ (.Y(_0336_),
    .A(_0333_),
    .B(_0335_));
 sg13g2_nand2_1 _2932_ (.Y(_0337_),
    .A(net178),
    .B(_0336_));
 sg13g2_nand3_1 _2933_ (.B(_1803_),
    .C(_0337_),
    .A(net172),
    .Y(_0338_));
 sg13g2_nor2_1 _2934_ (.A(_0258_),
    .B(_0338_),
    .Y(_0339_));
 sg13g2_nor2_1 _2935_ (.A(_0332_),
    .B(_0339_),
    .Y(_0340_));
 sg13g2_nand2_1 _2936_ (.Y(_0341_),
    .A(_0258_),
    .B(_0338_));
 sg13g2_a21oi_1 _2937_ (.A1(_0332_),
    .A2(_0341_),
    .Y(_0342_),
    .B1(_0340_));
 sg13g2_nand3_1 _2938_ (.B(_0308_),
    .C(_0309_),
    .A(_0304_),
    .Y(_0343_));
 sg13g2_nand2b_1 _2939_ (.Y(_0344_),
    .B(_0343_),
    .A_N(_0310_));
 sg13g2_xnor2_1 _2940_ (.Y(_0345_),
    .A(_0327_),
    .B(_0344_));
 sg13g2_nor2_1 _2941_ (.A(_1817_),
    .B(_0345_),
    .Y(_0346_));
 sg13g2_or4_1 _2942_ (.A(net173),
    .B(net174),
    .C(net176),
    .D(_0345_),
    .X(_0347_));
 sg13g2_xnor2_1 _2943_ (.Y(_0348_),
    .A(_0214_),
    .B(_0347_));
 sg13g2_nand2_1 _2944_ (.Y(_0349_),
    .A(_0338_),
    .B(_0348_));
 sg13g2_o21ai_1 _2945_ (.B1(_0349_),
    .Y(_0350_),
    .A1(_0213_),
    .A2(_0347_));
 sg13g2_inv_1 _2946_ (.Y(_0351_),
    .A(_0350_));
 sg13g2_xnor2_1 _2947_ (.Y(_0352_),
    .A(_0257_),
    .B(_0338_));
 sg13g2_xnor2_1 _2948_ (.Y(_0353_),
    .A(_0331_),
    .B(_0352_));
 sg13g2_inv_1 _2949_ (.Y(_0354_),
    .A(_0353_));
 sg13g2_xnor2_1 _2950_ (.Y(_0355_),
    .A(_0305_),
    .B(_0307_));
 sg13g2_xor2_1 _2951_ (.B(_0355_),
    .A(_0333_),
    .X(_0356_));
 sg13g2_or4_1 _2952_ (.A(net173),
    .B(net174),
    .C(net176),
    .D(_0356_),
    .X(_0357_));
 sg13g2_nor2_1 _2953_ (.A(_0179_),
    .B(_0357_),
    .Y(_0358_));
 sg13g2_xor2_1 _2954_ (.B(_0357_),
    .A(_0179_),
    .X(_0359_));
 sg13g2_a21oi_1 _2955_ (.A1(_0346_),
    .A2(_0359_),
    .Y(_0360_),
    .B1(_0358_));
 sg13g2_xnor2_1 _2956_ (.Y(_0361_),
    .A(_0338_),
    .B(_0348_));
 sg13g2_nor2_1 _2957_ (.A(_0360_),
    .B(_0361_),
    .Y(_0362_));
 sg13g2_nand2_1 _2958_ (.Y(_0363_),
    .A(_0247_),
    .B(_0331_));
 sg13g2_xnor2_1 _2959_ (.Y(_0364_),
    .A(_0242_),
    .B(_0344_));
 sg13g2_or4_1 _2960_ (.A(net173),
    .B(net174),
    .C(net176),
    .D(_0364_),
    .X(_0365_));
 sg13g2_a21o_1 _2961_ (.A2(_0330_),
    .A1(_0246_),
    .B1(_0365_),
    .X(_0366_));
 sg13g2_nand3_1 _2962_ (.B(_0363_),
    .C(_0366_),
    .A(_0357_),
    .Y(_0367_));
 sg13g2_xnor2_1 _2963_ (.Y(_0368_),
    .A(_0208_),
    .B(_0355_));
 sg13g2_nand4_1 _2964_ (.B(net175),
    .C(net178),
    .A(net172),
    .Y(_0369_),
    .D(_0368_));
 sg13g2_or2_1 _2965_ (.X(_0370_),
    .B(_0369_),
    .A(net245));
 sg13g2_xnor2_1 _2966_ (.Y(_0371_),
    .A(net245),
    .B(_0369_));
 sg13g2_or2_1 _2967_ (.X(_0372_),
    .B(_0371_),
    .A(_0365_));
 sg13g2_xnor2_1 _2968_ (.Y(_0373_),
    .A(_0346_),
    .B(_0359_));
 sg13g2_a21oi_1 _2969_ (.A1(_0370_),
    .A2(_0372_),
    .Y(_0374_),
    .B1(_0373_));
 sg13g2_and3_1 _2970_ (.X(_0375_),
    .A(_0370_),
    .B(_0372_),
    .C(_0373_));
 sg13g2_nand2_1 _2971_ (.Y(_0376_),
    .A(_0360_),
    .B(_0361_));
 sg13g2_xor2_1 _2972_ (.B(_0371_),
    .A(_0365_),
    .X(_0377_));
 sg13g2_a21oi_1 _2973_ (.A1(_0363_),
    .A2(_0366_),
    .Y(_0378_),
    .B1(_0357_));
 sg13g2_xnor2_1 _2974_ (.Y(_0379_),
    .A(_0360_),
    .B(_0361_));
 sg13g2_a21oi_1 _2975_ (.A1(_0367_),
    .A2(_0377_),
    .Y(_0380_),
    .B1(_0378_));
 sg13g2_or4_1 _2976_ (.A(_0374_),
    .B(_0375_),
    .C(_0379_),
    .D(_0380_),
    .X(_0381_));
 sg13g2_a221oi_1 _2977_ (.B2(_0376_),
    .C1(_0362_),
    .B1(_0374_),
    .A1(_0350_),
    .Y(_0382_),
    .A2(_0354_));
 sg13g2_a22oi_1 _2978_ (.Y(_0383_),
    .B1(_0381_),
    .B2(_0382_),
    .A2(_0353_),
    .A1(_0351_));
 sg13g2_nor2_1 _2979_ (.A(_0342_),
    .B(_0383_),
    .Y(_0384_));
 sg13g2_a21oi_1 _2980_ (.A1(_0342_),
    .A2(_0383_),
    .Y(_0385_),
    .B1(_0275_));
 sg13g2_nor2b_2 _2981_ (.A(_0384_),
    .B_N(_0385_),
    .Y(uo_out[5]));
 sg13g2_a21oi_1 _2982_ (.A1(_0342_),
    .A2(_0383_),
    .Y(_0386_),
    .B1(_0340_));
 sg13g2_nor2_2 _2983_ (.A(_0275_),
    .B(_0386_),
    .Y(uo_out[1]));
 sg13g2_xnor2_1 _2984_ (.Y(_0387_),
    .A(\sin_x_acc[23] ),
    .B(_1810_));
 sg13g2_nand2b_1 _2985_ (.Y(_0388_),
    .B(_0387_),
    .A_N(\cos_y_acc[23] ));
 sg13g2_o21ai_1 _2986_ (.B1(_0388_),
    .Y(_0389_),
    .A1(\sin_x_acc[23] ),
    .A2(_1811_));
 sg13g2_xnor2_1 _2987_ (.Y(_0390_),
    .A(\sin_y_acc[24] ),
    .B(\cos_x_acc[24] ));
 sg13g2_a21oi_1 _2988_ (.A1(_1807_),
    .A2(_1809_),
    .Y(_0391_),
    .B1(_1806_));
 sg13g2_nand2b_1 _2989_ (.Y(_0392_),
    .B(_0390_),
    .A_N(_0391_));
 sg13g2_xnor2_1 _2990_ (.Y(_0393_),
    .A(_0390_),
    .B(_0391_));
 sg13g2_xnor2_1 _2991_ (.Y(_0394_),
    .A(\sin_x_acc[24] ),
    .B(_0393_));
 sg13g2_nor2b_1 _2992_ (.A(\cos_y_acc[24] ),
    .B_N(_0394_),
    .Y(_0395_));
 sg13g2_xnor2_1 _2993_ (.Y(_0396_),
    .A(\cos_y_acc[24] ),
    .B(_0394_));
 sg13g2_and2_1 _2994_ (.A(_0389_),
    .B(_0396_),
    .X(_0397_));
 sg13g2_xnor2_1 _2995_ (.Y(_0398_),
    .A(\sin_x_acc[22] ),
    .B(_1334_));
 sg13g2_nand2b_1 _2996_ (.Y(_0399_),
    .B(_0398_),
    .A_N(net247));
 sg13g2_o21ai_1 _2997_ (.B1(_0399_),
    .Y(_0400_),
    .A1(\sin_x_acc[22] ),
    .A2(_1335_));
 sg13g2_xnor2_1 _2998_ (.Y(_0401_),
    .A(\cos_y_acc[23] ),
    .B(_0387_));
 sg13g2_a21oi_1 _2999_ (.A1(_1193_),
    .A2(_0318_),
    .Y(_0402_),
    .B1(_0317_));
 sg13g2_xnor2_1 _3000_ (.Y(_0403_),
    .A(net247),
    .B(_0398_));
 sg13g2_nand2b_1 _3001_ (.Y(_0404_),
    .B(_0403_),
    .A_N(_0402_));
 sg13g2_xnor2_1 _3002_ (.Y(_0405_),
    .A(_0402_),
    .B(_0403_));
 sg13g2_o21ai_1 _3003_ (.B1(_0405_),
    .Y(_0406_),
    .A1(_0320_),
    .A2(_0323_));
 sg13g2_xnor2_1 _3004_ (.Y(_0407_),
    .A(_0400_),
    .B(_0401_));
 sg13g2_a21oi_1 _3005_ (.A1(_0404_),
    .A2(_0406_),
    .Y(_0408_),
    .B1(_0407_));
 sg13g2_a21o_1 _3006_ (.A2(_0401_),
    .A1(_0400_),
    .B1(_0408_),
    .X(_0409_));
 sg13g2_xor2_1 _3007_ (.B(_0396_),
    .A(_0389_),
    .X(_0410_));
 sg13g2_a21oi_1 _3008_ (.A1(_0409_),
    .A2(_0410_),
    .Y(_0411_),
    .B1(_0397_));
 sg13g2_a21oi_1 _3009_ (.A1(_1223_),
    .A2(_0393_),
    .Y(_0412_),
    .B1(_0395_));
 sg13g2_inv_1 _3010_ (.Y(_0413_),
    .A(_0412_));
 sg13g2_nor2b_1 _3011_ (.A(\sin_y_acc[25] ),
    .B_N(\cos_x_acc[25] ),
    .Y(_0414_));
 sg13g2_nand2b_1 _3012_ (.Y(_0415_),
    .B(\sin_y_acc[25] ),
    .A_N(\cos_x_acc[25] ));
 sg13g2_nand2b_1 _3013_ (.Y(_0416_),
    .B(_0415_),
    .A_N(_0414_));
 sg13g2_o21ai_1 _3014_ (.B1(_0392_),
    .Y(_0417_),
    .A1(\sin_y_acc[24] ),
    .A2(_1221_));
 sg13g2_xnor2_1 _3015_ (.Y(_0418_),
    .A(_0416_),
    .B(_0417_));
 sg13g2_xnor2_1 _3016_ (.Y(_0419_),
    .A(\sin_x_acc[25] ),
    .B(_0418_));
 sg13g2_nor2b_1 _3017_ (.A(\cos_y_acc[25] ),
    .B_N(_0419_),
    .Y(_0420_));
 sg13g2_xnor2_1 _3018_ (.Y(_0421_),
    .A(\cos_y_acc[25] ),
    .B(_0419_));
 sg13g2_xnor2_1 _3019_ (.Y(_0422_),
    .A(_0412_),
    .B(_0421_));
 sg13g2_nor2b_1 _3020_ (.A(_0411_),
    .B_N(_0422_),
    .Y(_0423_));
 sg13g2_xnor2_1 _3021_ (.Y(_0424_),
    .A(_0411_),
    .B(_0422_));
 sg13g2_nand2_1 _3022_ (.Y(_0425_),
    .A(_1815_),
    .B(_0424_));
 sg13g2_nor2b_2 _3023_ (.A(_1805_),
    .B_N(_0425_),
    .Y(_0426_));
 sg13g2_nand3_1 _3024_ (.B(net175),
    .C(_0425_),
    .A(net172),
    .Y(_0427_));
 sg13g2_a21oi_1 _3025_ (.A1(_0413_),
    .A2(_0421_),
    .Y(_0428_),
    .B1(_0423_));
 sg13g2_xnor2_1 _3026_ (.Y(_0429_),
    .A(_0409_),
    .B(_0410_));
 sg13g2_a21o_1 _3027_ (.A2(_0418_),
    .A1(_1222_),
    .B1(_0420_),
    .X(_0430_));
 sg13g2_xor2_1 _3028_ (.B(\sin_x_acc[26] ),
    .A(\cos_x_acc[26] ),
    .X(_0431_));
 sg13g2_xor2_1 _3029_ (.B(\sin_y_acc[26] ),
    .A(\cos_y_acc[26] ),
    .X(_0432_));
 sg13g2_xnor2_1 _3030_ (.Y(_0433_),
    .A(_0431_),
    .B(_0432_));
 sg13g2_a21oi_1 _3031_ (.A1(_0415_),
    .A2(_0417_),
    .Y(_0434_),
    .B1(_0414_));
 sg13g2_xnor2_1 _3032_ (.Y(_0435_),
    .A(_0433_),
    .B(_0434_));
 sg13g2_xnor2_1 _3033_ (.Y(_0436_),
    .A(_0430_),
    .B(_0435_));
 sg13g2_xor2_1 _3034_ (.B(_0436_),
    .A(_0429_),
    .X(_0437_));
 sg13g2_xnor2_1 _3035_ (.Y(_0438_),
    .A(_0428_),
    .B(_0437_));
 sg13g2_a21oi_2 _3036_ (.B1(_1805_),
    .Y(_0439_),
    .A2(_0438_),
    .A1(_1815_));
 sg13g2_a21oi_1 _3037_ (.A1(_0257_),
    .A2(_0439_),
    .Y(_0440_),
    .B1(_0426_));
 sg13g2_o21ai_1 _3038_ (.B1(_0426_),
    .Y(_0441_),
    .A1(_0257_),
    .A2(_0439_));
 sg13g2_nor2b_1 _3039_ (.A(_0440_),
    .B_N(_0441_),
    .Y(_0442_));
 sg13g2_nand3_1 _3040_ (.B(_0406_),
    .C(_0407_),
    .A(_0404_),
    .Y(_0443_));
 sg13g2_nand2b_1 _3041_ (.Y(_0444_),
    .B(_0443_),
    .A_N(_0408_));
 sg13g2_xor2_1 _3042_ (.B(_0444_),
    .A(_0424_),
    .X(_0445_));
 sg13g2_nor4_2 _3043_ (.A(net173),
    .B(net174),
    .C(net177),
    .Y(_0446_),
    .D(_0445_));
 sg13g2_nand2_1 _3044_ (.Y(_0447_),
    .A(_0214_),
    .B(_0446_));
 sg13g2_xnor2_1 _3045_ (.Y(_0448_),
    .A(_0214_),
    .B(_0446_));
 sg13g2_o21ai_1 _3046_ (.B1(_0447_),
    .Y(_0449_),
    .A1(_0439_),
    .A2(_0448_));
 sg13g2_xnor2_1 _3047_ (.Y(_0450_),
    .A(_0258_),
    .B(_0439_));
 sg13g2_xnor2_1 _3048_ (.Y(_0451_),
    .A(_0426_),
    .B(_0450_));
 sg13g2_nor2_1 _3049_ (.A(_0449_),
    .B(_0451_),
    .Y(_0452_));
 sg13g2_or3_1 _3050_ (.A(_0320_),
    .B(_0323_),
    .C(_0405_),
    .X(_0453_));
 sg13g2_nand2_1 _3051_ (.Y(_0454_),
    .A(_0406_),
    .B(_0453_));
 sg13g2_xnor2_1 _3052_ (.Y(_0455_),
    .A(_0429_),
    .B(_0454_));
 sg13g2_nor4_2 _3053_ (.A(_1775_),
    .B(_1804_),
    .C(net177),
    .Y(_0456_),
    .D(_0455_));
 sg13g2_xnor2_1 _3054_ (.Y(_0457_),
    .A(_0325_),
    .B(_0444_));
 sg13g2_nor4_2 _3055_ (.A(_1775_),
    .B(_1804_),
    .C(net177),
    .Y(_0458_),
    .D(_0457_));
 sg13g2_nand2_1 _3056_ (.Y(_0459_),
    .A(_0246_),
    .B(_0425_));
 sg13g2_a22oi_1 _3057_ (.Y(_0460_),
    .B1(_0458_),
    .B2(_0459_),
    .A2(_0427_),
    .A1(_0247_));
 sg13g2_nor2b_1 _3058_ (.A(_0456_),
    .B_N(_0460_),
    .Y(_0461_));
 sg13g2_nor2b_1 _3059_ (.A(_0179_),
    .B_N(_0456_),
    .Y(_0462_));
 sg13g2_nand2b_1 _3060_ (.Y(_0463_),
    .B(_0179_),
    .A_N(_0456_));
 sg13g2_xnor2_1 _3061_ (.Y(_0464_),
    .A(_0179_),
    .B(_0456_));
 sg13g2_a21oi_1 _3062_ (.A1(_0446_),
    .A2(_0463_),
    .Y(_0465_),
    .B1(_0462_));
 sg13g2_a21o_1 _3063_ (.A2(_0463_),
    .A1(_0446_),
    .B1(_0462_),
    .X(_0466_));
 sg13g2_xor2_1 _3064_ (.B(_0448_),
    .A(_0439_),
    .X(_0467_));
 sg13g2_xnor2_1 _3065_ (.Y(_0468_),
    .A(_0439_),
    .B(_0448_));
 sg13g2_nor2_1 _3066_ (.A(_0465_),
    .B(_0468_),
    .Y(_0469_));
 sg13g2_a21oi_1 _3067_ (.A1(_0466_),
    .A2(_0467_),
    .Y(_0470_),
    .B1(_0461_));
 sg13g2_or2_1 _3068_ (.X(_0471_),
    .B(_0454_),
    .A(_0335_));
 sg13g2_a21oi_1 _3069_ (.A1(_0335_),
    .A2(_0454_),
    .Y(_0472_),
    .B1(net176));
 sg13g2_nand4_1 _3070_ (.B(_1803_),
    .C(_0471_),
    .A(_1776_),
    .Y(_0473_),
    .D(_0472_));
 sg13g2_nor2_1 _3071_ (.A(net245),
    .B(_0473_),
    .Y(_0474_));
 sg13g2_nand2_1 _3072_ (.Y(_0475_),
    .A(_0178_),
    .B(_0473_));
 sg13g2_xnor2_1 _3073_ (.Y(_0476_),
    .A(net245),
    .B(_0473_));
 sg13g2_xnor2_1 _3074_ (.Y(_0477_),
    .A(_0458_),
    .B(_0476_));
 sg13g2_nor2b_1 _3075_ (.A(_0460_),
    .B_N(_0456_),
    .Y(_0478_));
 sg13g2_or2_1 _3076_ (.X(_0479_),
    .B(_0478_),
    .A(_0477_));
 sg13g2_a21oi_1 _3077_ (.A1(_0458_),
    .A2(_0475_),
    .Y(_0480_),
    .B1(_0474_));
 sg13g2_xnor2_1 _3078_ (.Y(_0481_),
    .A(_0446_),
    .B(_0464_));
 sg13g2_nor2_1 _3079_ (.A(_0480_),
    .B(_0481_),
    .Y(_0482_));
 sg13g2_nand2_1 _3080_ (.Y(_0483_),
    .A(_0465_),
    .B(_0468_));
 sg13g2_xor2_1 _3081_ (.B(_0481_),
    .A(_0480_),
    .X(_0484_));
 sg13g2_nand4_1 _3082_ (.B(_0479_),
    .C(_0483_),
    .A(_0470_),
    .Y(_0485_),
    .D(_0484_));
 sg13g2_a221oi_1 _3083_ (.B2(_0483_),
    .C1(_0469_),
    .B1(_0482_),
    .A1(_0449_),
    .Y(_0486_),
    .A2(_0451_));
 sg13g2_a21oi_1 _3084_ (.A1(_0485_),
    .A2(_0486_),
    .Y(_0487_),
    .B1(_0452_));
 sg13g2_nor2_1 _3085_ (.A(_0442_),
    .B(_0487_),
    .Y(_0488_));
 sg13g2_a21oi_1 _3086_ (.A1(_0442_),
    .A2(_0487_),
    .Y(_0489_),
    .B1(_0275_));
 sg13g2_nor2b_2 _3087_ (.A(_0488_),
    .B_N(_0489_),
    .Y(uo_out[4]));
 sg13g2_a21oi_1 _3088_ (.A1(_0442_),
    .A2(_0487_),
    .Y(_0490_),
    .B1(_0440_));
 sg13g2_nor2_2 _3089_ (.A(_0275_),
    .B(_0490_),
    .Y(uo_out[0]));
 sg13g2_and2_1 _3090_ (.A(\hvsync_gen.vpos[2] ),
    .B(\hvsync_gen.vpos[3] ),
    .X(_0491_));
 sg13g2_nand3b_1 _3091_ (.B(\hvsync_gen.vpos[3] ),
    .C(net246),
    .Y(_0492_),
    .A_N(\hvsync_gen.vpos[9] ));
 sg13g2_nor4_1 _3092_ (.A(net271),
    .B(_0274_),
    .C(_0491_),
    .D(_0492_),
    .Y(_0001_));
 sg13g2_and3_1 _3093_ (.X(_0493_),
    .A(\hvsync_gen.hpos[4] ),
    .B(net302),
    .C(net329));
 sg13g2_nand3_1 _3094_ (.B(\hvsync_gen.hpos[7] ),
    .C(net292),
    .A(_1217_),
    .Y(_0494_));
 sg13g2_nor3_1 _3095_ (.A(\hvsync_gen.hpos[4] ),
    .B(\hvsync_gen.hpos[5] ),
    .C(\hvsync_gen.hpos[6] ),
    .Y(_0495_));
 sg13g2_nor3_1 _3096_ (.A(_0493_),
    .B(net293),
    .C(_0495_),
    .Y(_0000_));
 sg13g2_xnor2_1 _3097_ (.Y(_0496_),
    .A(net249),
    .B(net251));
 sg13g2_xor2_1 _3098_ (.B(net251),
    .A(net249),
    .X(_0497_));
 sg13g2_xor2_1 _3099_ (.B(\cos_addr[1] ),
    .A(net249),
    .X(_0498_));
 sg13g2_xnor2_1 _3100_ (.Y(_0499_),
    .A(net249),
    .B(\cos_addr[1] ));
 sg13g2_xnor2_1 _3101_ (.Y(_0500_),
    .A(net249),
    .B(\cos_addr[2] ));
 sg13g2_xor2_1 _3102_ (.B(\cos_addr[2] ),
    .A(net249),
    .X(_0501_));
 sg13g2_nor2_2 _3103_ (.A(net241),
    .B(net237),
    .Y(_0502_));
 sg13g2_o21ai_1 _3104_ (.B1(net244),
    .Y(_0503_),
    .A1(net241),
    .A2(net238));
 sg13g2_nand2_1 _3105_ (.Y(_0504_),
    .A(_0497_),
    .B(net240));
 sg13g2_nand2_1 _3106_ (.Y(_0505_),
    .A(net249),
    .B(\cos_addr[3] ));
 sg13g2_or2_1 _3107_ (.X(_0506_),
    .B(\cos_addr[3] ),
    .A(net249));
 sg13g2_xnor2_1 _3108_ (.Y(_0507_),
    .A(net250),
    .B(\cos_addr[3] ));
 sg13g2_xor2_1 _3109_ (.B(\cos_addr[3] ),
    .A(net250),
    .X(_0508_));
 sg13g2_xnor2_1 _3110_ (.Y(_0509_),
    .A(net250),
    .B(\cos_addr[4] ));
 sg13g2_xor2_1 _3111_ (.B(\cos_addr[4] ),
    .A(net250),
    .X(_0510_));
 sg13g2_nor2_2 _3112_ (.A(net230),
    .B(net223),
    .Y(_0511_));
 sg13g2_nand2_1 _3113_ (.Y(_0512_),
    .A(net232),
    .B(net227));
 sg13g2_a221oi_1 _3114_ (.B2(_0506_),
    .C1(net225),
    .B1(_0505_),
    .A1(net242),
    .Y(_0513_),
    .A2(net240));
 sg13g2_nor2_2 _3115_ (.A(_0507_),
    .B(net225),
    .Y(_0514_));
 sg13g2_mux2_1 _3116_ (.A0(_0514_),
    .A1(_0513_),
    .S(_0503_),
    .X(_0515_));
 sg13g2_nor2_1 _3117_ (.A(net230),
    .B(net228),
    .Y(_0516_));
 sg13g2_nor2_2 _3118_ (.A(net242),
    .B(net237),
    .Y(_0517_));
 sg13g2_nor2_1 _3119_ (.A(net241),
    .B(net235),
    .Y(_0518_));
 sg13g2_nand2_1 _3120_ (.Y(_0519_),
    .A(net239),
    .B(net237));
 sg13g2_nor2_1 _3121_ (.A(net240),
    .B(net236),
    .Y(_0520_));
 sg13g2_nor2_2 _3122_ (.A(net236),
    .B(net231),
    .Y(_0521_));
 sg13g2_nor2_2 _3123_ (.A(net242),
    .B(net229),
    .Y(_0522_));
 sg13g2_o21ai_1 _3124_ (.B1(net234),
    .Y(_0523_),
    .A1(net244),
    .A2(net238));
 sg13g2_nor3_1 _3125_ (.A(net228),
    .B(_0520_),
    .C(_0523_),
    .Y(_0524_));
 sg13g2_xor2_1 _3126_ (.B(\cos_addr[5] ),
    .A(net250),
    .X(_0525_));
 sg13g2_xnor2_1 _3127_ (.Y(_0526_),
    .A(net250),
    .B(\cos_addr[5] ));
 sg13g2_nor2_2 _3128_ (.A(net239),
    .B(net238),
    .Y(_0527_));
 sg13g2_nor2_1 _3129_ (.A(net244),
    .B(net239),
    .Y(_0528_));
 sg13g2_nor4_1 _3130_ (.A(net234),
    .B(net228),
    .C(_0527_),
    .D(net215),
    .Y(_0529_));
 sg13g2_or4_1 _3131_ (.A(_0515_),
    .B(_0524_),
    .C(net219),
    .D(_0529_),
    .X(_0530_));
 sg13g2_nor2_1 _3132_ (.A(net235),
    .B(net214),
    .Y(_0531_));
 sg13g2_o21ai_1 _3133_ (.B1(_0500_),
    .Y(_0532_),
    .A1(net244),
    .A2(net240));
 sg13g2_nor2_2 _3134_ (.A(net242),
    .B(net239),
    .Y(_0533_));
 sg13g2_nand2_1 _3135_ (.Y(_0534_),
    .A(net243),
    .B(net241));
 sg13g2_o21ai_1 _3136_ (.B1(net236),
    .Y(_0535_),
    .A1(net244),
    .A2(net241));
 sg13g2_xnor2_1 _3137_ (.Y(_0536_),
    .A(\cos_addr[1] ),
    .B(net251));
 sg13g2_nand2_1 _3138_ (.Y(_0537_),
    .A(net235),
    .B(net217));
 sg13g2_a21oi_1 _3139_ (.A1(_0532_),
    .A2(_0537_),
    .Y(_0538_),
    .B1(net231));
 sg13g2_mux2_1 _3140_ (.A0(_0496_),
    .A1(_0498_),
    .S(net238),
    .X(_0539_));
 sg13g2_a21oi_1 _3141_ (.A1(net243),
    .A2(net240),
    .Y(_0540_),
    .B1(net238));
 sg13g2_o21ai_1 _3142_ (.B1(net235),
    .Y(_0541_),
    .A1(net242),
    .A2(net241));
 sg13g2_nand2_1 _3143_ (.Y(_0542_),
    .A(net243),
    .B(net216));
 sg13g2_nor3_2 _3144_ (.A(net242),
    .B(_0498_),
    .C(_0500_),
    .Y(_0543_));
 sg13g2_a21oi_1 _3145_ (.A1(_0496_),
    .A2(net239),
    .Y(_0544_),
    .B1(net236));
 sg13g2_o21ai_1 _3146_ (.B1(net231),
    .Y(_0545_),
    .A1(_0543_),
    .A2(net213));
 sg13g2_nand2_1 _3147_ (.Y(_0546_),
    .A(_0507_),
    .B(_0539_));
 sg13g2_a21oi_1 _3148_ (.A1(_0545_),
    .A2(_0546_),
    .Y(_0547_),
    .B1(net225));
 sg13g2_o21ai_1 _3149_ (.B1(net225),
    .Y(_0548_),
    .A1(net234),
    .A2(_0539_));
 sg13g2_o21ai_1 _3150_ (.B1(net219),
    .Y(_0549_),
    .A1(_0538_),
    .A2(_0548_));
 sg13g2_o21ai_1 _3151_ (.B1(_0530_),
    .Y(_0550_),
    .A1(_0547_),
    .A2(_0549_));
 sg13g2_or2_1 _3152_ (.X(_0551_),
    .B(net187),
    .A(net318));
 sg13g2_nor3_1 _3153_ (.A(\hvsync_gen.hpos[2] ),
    .B(\hvsync_gen.hpos[9] ),
    .C(\hvsync_gen.hpos[3] ),
    .Y(_0552_));
 sg13g2_nor2_1 _3154_ (.A(net165),
    .B(net452),
    .Y(_0553_));
 sg13g2_and4_1 _3155_ (.A(_0271_),
    .B(_0495_),
    .C(_0552_),
    .D(_0553_),
    .X(_0554_));
 sg13g2_nand4_1 _3156_ (.B(_0495_),
    .C(_0552_),
    .A(_0271_),
    .Y(_0555_),
    .D(_0553_));
 sg13g2_nand2_2 _3157_ (.Y(_0556_),
    .A(net318),
    .B(net187));
 sg13g2_and3_1 _3158_ (.X(_0002_),
    .A(_0551_),
    .B(net203),
    .C(_0556_));
 sg13g2_o21ai_1 _3159_ (.B1(net231),
    .Y(_0557_),
    .A1(_0517_),
    .A2(net213));
 sg13g2_nand3_1 _3160_ (.B(net239),
    .C(net238),
    .A(net242),
    .Y(_0558_));
 sg13g2_nand3_1 _3161_ (.B(_0535_),
    .C(_0558_),
    .A(net234),
    .Y(_0559_));
 sg13g2_nand3_1 _3162_ (.B(_0557_),
    .C(_0559_),
    .A(net222),
    .Y(_0560_));
 sg13g2_nor2_1 _3163_ (.A(net235),
    .B(_0533_),
    .Y(_0561_));
 sg13g2_and2_1 _3164_ (.A(net238),
    .B(net217),
    .X(_0562_));
 sg13g2_nor2_1 _3165_ (.A(_0517_),
    .B(net217),
    .Y(_0563_));
 sg13g2_nor2_1 _3166_ (.A(net243),
    .B(_0520_),
    .Y(_0564_));
 sg13g2_nand2_1 _3167_ (.Y(_0565_),
    .A(_0532_),
    .B(_0541_));
 sg13g2_a221oi_1 _3168_ (.B2(_0514_),
    .C1(net220),
    .B1(_0565_),
    .A1(_0511_),
    .Y(_0566_),
    .A2(_0563_));
 sg13g2_nor2_1 _3169_ (.A(_0502_),
    .B(_0536_),
    .Y(_0567_));
 sg13g2_o21ai_1 _3170_ (.B1(net225),
    .Y(_0568_),
    .A1(_0538_),
    .A2(_0567_));
 sg13g2_nand2_1 _3171_ (.Y(_0569_),
    .A(net241),
    .B(net232));
 sg13g2_o21ai_1 _3172_ (.B1(net230),
    .Y(_0570_),
    .A1(_0517_),
    .A2(net217));
 sg13g2_a21oi_1 _3173_ (.A1(net241),
    .A2(net234),
    .Y(_0571_),
    .B1(net223));
 sg13g2_nand2_1 _3174_ (.Y(_0572_),
    .A(net226),
    .B(_0569_));
 sg13g2_a21oi_1 _3175_ (.A1(_0570_),
    .A2(_0571_),
    .Y(_0573_),
    .B1(net219));
 sg13g2_a22oi_1 _3176_ (.Y(_0574_),
    .B1(_0568_),
    .B2(_0573_),
    .A2(_0566_),
    .A1(_0560_));
 sg13g2_nand2_1 _3177_ (.Y(_0575_),
    .A(net489),
    .B(_0574_));
 sg13g2_xnor2_1 _3178_ (.Y(_0576_),
    .A(\cos_x_acc[1] ),
    .B(_0574_));
 sg13g2_o21ai_1 _3179_ (.B1(net203),
    .Y(_0577_),
    .A1(_0556_),
    .A2(_0576_));
 sg13g2_a21oi_1 _3180_ (.A1(_0556_),
    .A2(_0576_),
    .Y(_0003_),
    .B1(_0577_));
 sg13g2_nand2_2 _3181_ (.Y(_0578_),
    .A(net237),
    .B(net229));
 sg13g2_nor2_2 _3182_ (.A(net237),
    .B(net229),
    .Y(_0579_));
 sg13g2_nand2_2 _3183_ (.Y(_0580_),
    .A(net235),
    .B(net234));
 sg13g2_a21oi_1 _3184_ (.A1(_0578_),
    .A2(_0580_),
    .Y(_0581_),
    .B1(net243));
 sg13g2_nand2_1 _3185_ (.Y(_0582_),
    .A(_0504_),
    .B(net225));
 sg13g2_nor2_1 _3186_ (.A(_0581_),
    .B(_0582_),
    .Y(_0583_));
 sg13g2_nand2b_1 _3187_ (.Y(_0584_),
    .B(_0535_),
    .A_N(net213));
 sg13g2_nand2_1 _3188_ (.Y(_0585_),
    .A(net239),
    .B(net229));
 sg13g2_o21ai_1 _3189_ (.B1(net230),
    .Y(_0586_),
    .A1(_0518_),
    .A2(_0540_));
 sg13g2_mux2_1 _3190_ (.A0(net231),
    .A1(_0586_),
    .S(_0584_),
    .X(_0587_));
 sg13g2_a21oi_1 _3191_ (.A1(net228),
    .A2(_0587_),
    .Y(_0588_),
    .B1(_0583_));
 sg13g2_o21ai_1 _3192_ (.B1(_0503_),
    .Y(_0589_),
    .A1(_0504_),
    .A2(_0521_));
 sg13g2_o21ai_1 _3193_ (.B1(net233),
    .Y(_0590_),
    .A1(net237),
    .A2(_0534_));
 sg13g2_nor2_1 _3194_ (.A(net228),
    .B(net217),
    .Y(_0591_));
 sg13g2_a21oi_1 _3195_ (.A1(_0590_),
    .A2(_0591_),
    .Y(_0592_),
    .B1(net218));
 sg13g2_o21ai_1 _3196_ (.B1(_0592_),
    .Y(_0593_),
    .A1(_0572_),
    .A2(_0589_));
 sg13g2_o21ai_1 _3197_ (.B1(_0593_),
    .Y(_0594_),
    .A1(net220),
    .A2(_0588_));
 sg13g2_inv_1 _3198_ (.Y(_0595_),
    .A(_0594_));
 sg13g2_xor2_1 _3199_ (.B(_0594_),
    .A(\cos_x_acc[2] ),
    .X(_0596_));
 sg13g2_o21ai_1 _3200_ (.B1(_0575_),
    .Y(_0597_),
    .A1(_0556_),
    .A2(_0576_));
 sg13g2_nor2b_1 _3201_ (.A(_0597_),
    .B_N(_0596_),
    .Y(_0598_));
 sg13g2_nor2b_1 _3202_ (.A(_0596_),
    .B_N(_0597_),
    .Y(_0599_));
 sg13g2_nor3_1 _3203_ (.A(net211),
    .B(net490),
    .C(_0599_),
    .Y(_0004_));
 sg13g2_a21oi_2 _3204_ (.B1(net224),
    .Y(_0600_),
    .A2(_0533_),
    .A1(net233));
 sg13g2_nand3_1 _3205_ (.B(_0580_),
    .C(_0600_),
    .A(_0565_),
    .Y(_0601_));
 sg13g2_nor2_2 _3206_ (.A(net228),
    .B(_0521_),
    .Y(_0602_));
 sg13g2_o21ai_1 _3207_ (.B1(_0602_),
    .Y(_0603_),
    .A1(_0520_),
    .A2(net215));
 sg13g2_nor2_1 _3208_ (.A(_0511_),
    .B(net221),
    .Y(_0604_));
 sg13g2_a21oi_1 _3209_ (.A1(_0511_),
    .A2(_0543_),
    .Y(_0605_),
    .B1(net220));
 sg13g2_nand2_1 _3210_ (.Y(_0606_),
    .A(_0603_),
    .B(_0605_));
 sg13g2_nor2_1 _3211_ (.A(_0524_),
    .B(_0606_),
    .Y(_0607_));
 sg13g2_nand2_1 _3212_ (.Y(_0608_),
    .A(_0564_),
    .B(_0585_));
 sg13g2_a21oi_1 _3213_ (.A1(_0578_),
    .A2(_0608_),
    .Y(_0609_),
    .B1(net227));
 sg13g2_nor2_2 _3214_ (.A(net243),
    .B(net233),
    .Y(_0610_));
 sg13g2_nand2_1 _3215_ (.Y(_0611_),
    .A(net242),
    .B(net231));
 sg13g2_nor2_2 _3216_ (.A(net216),
    .B(_0527_),
    .Y(_0612_));
 sg13g2_a221oi_1 _3217_ (.B2(_0612_),
    .C1(net222),
    .B1(_0610_),
    .A1(net233),
    .Y(_0613_),
    .A2(_0527_));
 sg13g2_nor3_1 _3218_ (.A(net219),
    .B(_0609_),
    .C(_0613_),
    .Y(_0614_));
 sg13g2_a21oi_2 _3219_ (.B1(_0614_),
    .Y(_0615_),
    .A2(_0607_),
    .A1(_0601_));
 sg13g2_nand2b_1 _3220_ (.Y(_0616_),
    .B(net483),
    .A_N(_0615_));
 sg13g2_xnor2_1 _3221_ (.Y(_0617_),
    .A(net483),
    .B(_0615_));
 sg13g2_a21oi_1 _3222_ (.A1(net501),
    .A2(_0595_),
    .Y(_0618_),
    .B1(_0599_));
 sg13g2_nand2b_1 _3223_ (.Y(_0619_),
    .B(_0618_),
    .A_N(_0617_));
 sg13g2_nand2b_1 _3224_ (.Y(_0620_),
    .B(_0617_),
    .A_N(_0618_));
 sg13g2_and3_1 _3225_ (.X(_0005_),
    .A(net199),
    .B(_0619_),
    .C(_0620_));
 sg13g2_nor2_2 _3226_ (.A(net237),
    .B(net217),
    .Y(_0621_));
 sg13g2_a21oi_1 _3227_ (.A1(net230),
    .A2(net217),
    .Y(_0622_),
    .B1(net227));
 sg13g2_a21oi_1 _3228_ (.A1(net223),
    .A2(_0517_),
    .Y(_0623_),
    .B1(_0622_));
 sg13g2_nor2_1 _3229_ (.A(_0621_),
    .B(_0623_),
    .Y(_0624_));
 sg13g2_o21ai_1 _3230_ (.B1(net227),
    .Y(_0625_),
    .A1(net232),
    .A2(net216));
 sg13g2_or2_1 _3231_ (.X(_0626_),
    .B(net213),
    .A(_0502_));
 sg13g2_nor2b_1 _3232_ (.A(_0625_),
    .B_N(_0626_),
    .Y(_0627_));
 sg13g2_nor4_1 _3233_ (.A(net237),
    .B(net233),
    .C(net222),
    .D(_0534_),
    .Y(_0628_));
 sg13g2_nor4_1 _3234_ (.A(net220),
    .B(_0624_),
    .C(_0627_),
    .D(_0628_),
    .Y(_0629_));
 sg13g2_nor3_1 _3235_ (.A(net222),
    .B(net216),
    .C(net214),
    .Y(_0630_));
 sg13g2_o21ai_1 _3236_ (.B1(net220),
    .Y(_0631_),
    .A1(net226),
    .A2(_0535_));
 sg13g2_a21oi_1 _3237_ (.A1(_0611_),
    .A2(_0630_),
    .Y(_0632_),
    .B1(_0631_));
 sg13g2_nor2_2 _3238_ (.A(_0629_),
    .B(_0632_),
    .Y(_0633_));
 sg13g2_xnor2_1 _3239_ (.Y(_0634_),
    .A(_1228_),
    .B(_0633_));
 sg13g2_nand3_1 _3240_ (.B(_0620_),
    .C(_0634_),
    .A(_0616_),
    .Y(_0635_));
 sg13g2_a21o_1 _3241_ (.A2(_0620_),
    .A1(_0616_),
    .B1(_0634_),
    .X(_0636_));
 sg13g2_and3_1 _3242_ (.X(_0006_),
    .A(net199),
    .B(net484),
    .C(_0636_));
 sg13g2_o21ai_1 _3243_ (.B1(_0636_),
    .Y(_0637_),
    .A1(_1228_),
    .A2(_0633_));
 sg13g2_nor2_1 _3244_ (.A(net214),
    .B(_0579_),
    .Y(_0638_));
 sg13g2_o21ai_1 _3245_ (.B1(_0578_),
    .Y(_0639_),
    .A1(net214),
    .A2(_0579_));
 sg13g2_a221oi_1 _3246_ (.B2(_0542_),
    .C1(net226),
    .B1(_0639_),
    .A1(net214),
    .Y(_0640_),
    .A2(_0579_));
 sg13g2_nor2_1 _3247_ (.A(_0502_),
    .B(_0564_),
    .Y(_0641_));
 sg13g2_nand2_1 _3248_ (.Y(_0642_),
    .A(_0537_),
    .B(_0558_));
 sg13g2_inv_1 _3249_ (.Y(_0643_),
    .A(_0642_));
 sg13g2_a221oi_1 _3250_ (.B2(_0511_),
    .C1(_0640_),
    .B1(_0642_),
    .A1(_0514_),
    .Y(_0644_),
    .A2(_0641_));
 sg13g2_o21ai_1 _3251_ (.B1(net232),
    .Y(_0645_),
    .A1(_0517_),
    .A2(net213));
 sg13g2_o21ai_1 _3252_ (.B1(_0645_),
    .Y(_0646_),
    .A1(net232),
    .A2(_0541_));
 sg13g2_a221oi_1 _3253_ (.B2(net244),
    .C1(_0610_),
    .B1(_0521_),
    .A1(net240),
    .Y(_0647_),
    .A2(net235));
 sg13g2_a21oi_1 _3254_ (.A1(net227),
    .A2(_0647_),
    .Y(_0648_),
    .B1(net219));
 sg13g2_o21ai_1 _3255_ (.B1(_0648_),
    .Y(_0649_),
    .A1(net226),
    .A2(_0646_));
 sg13g2_o21ai_1 _3256_ (.B1(_0649_),
    .Y(_0650_),
    .A1(net220),
    .A2(_0644_));
 sg13g2_inv_1 _3257_ (.Y(_0651_),
    .A(_0650_));
 sg13g2_nand2b_1 _3258_ (.Y(_0652_),
    .B(_0650_),
    .A_N(net499));
 sg13g2_and2_1 _3259_ (.A(net457),
    .B(_0651_),
    .X(_0653_));
 sg13g2_xnor2_1 _3260_ (.Y(_0654_),
    .A(net457),
    .B(_0650_));
 sg13g2_o21ai_1 _3261_ (.B1(net199),
    .Y(_0655_),
    .A1(_0637_),
    .A2(_0654_));
 sg13g2_a21oi_1 _3262_ (.A1(_0637_),
    .A2(_0654_),
    .Y(_0007_),
    .B1(_0655_));
 sg13g2_a21oi_1 _3263_ (.A1(net235),
    .A2(net217),
    .Y(_0656_),
    .B1(net213));
 sg13g2_o21ai_1 _3264_ (.B1(_0611_),
    .Y(_0657_),
    .A1(net229),
    .A2(_0656_));
 sg13g2_nand3b_1 _3265_ (.B(_0557_),
    .C(_0580_),
    .Y(_0658_),
    .A_N(_0522_));
 sg13g2_a221oi_1 _3266_ (.B2(_0600_),
    .C1(net218),
    .B1(_0658_),
    .A1(net222),
    .Y(_0659_),
    .A2(_0657_));
 sg13g2_o21ai_1 _3267_ (.B1(_0535_),
    .Y(_0660_),
    .A1(_0522_),
    .A2(_0579_));
 sg13g2_nand2_1 _3268_ (.Y(_0661_),
    .A(net229),
    .B(_0564_));
 sg13g2_nand2_1 _3269_ (.Y(_0662_),
    .A(_0660_),
    .B(_0661_));
 sg13g2_a22oi_1 _3270_ (.Y(_0663_),
    .B1(_0662_),
    .B2(net222),
    .A2(_0531_),
    .A1(_0514_));
 sg13g2_a21o_2 _3271_ (.A2(_0663_),
    .A1(net218),
    .B1(_0659_),
    .X(_0664_));
 sg13g2_and2_1 _3272_ (.A(net496),
    .B(_0664_),
    .X(_0665_));
 sg13g2_xnor2_1 _3273_ (.Y(_0666_),
    .A(net496),
    .B(_0664_));
 sg13g2_a21oi_1 _3274_ (.A1(_0637_),
    .A2(_0652_),
    .Y(_0667_),
    .B1(_0653_));
 sg13g2_nor2_1 _3275_ (.A(_0666_),
    .B(_0667_),
    .Y(_0668_));
 sg13g2_a21oi_1 _3276_ (.A1(_0666_),
    .A2(_0667_),
    .Y(_0669_),
    .B1(net205));
 sg13g2_nor2b_1 _3277_ (.A(_0668_),
    .B_N(_0669_),
    .Y(_0008_));
 sg13g2_a21oi_1 _3278_ (.A1(net229),
    .A2(_0626_),
    .Y(_0670_),
    .B1(net226));
 sg13g2_o21ai_1 _3279_ (.B1(_0670_),
    .Y(_0671_),
    .A1(net216),
    .A2(_0590_));
 sg13g2_o21ai_1 _3280_ (.B1(net229),
    .Y(_0672_),
    .A1(net243),
    .A2(_0612_));
 sg13g2_nand3_1 _3281_ (.B(_0600_),
    .C(_0672_),
    .A(_0580_),
    .Y(_0673_));
 sg13g2_a21oi_1 _3282_ (.A1(_0671_),
    .A2(_0673_),
    .Y(_0674_),
    .B1(net220));
 sg13g2_o21ai_1 _3283_ (.B1(net233),
    .Y(_0675_),
    .A1(_0543_),
    .A2(_0544_));
 sg13g2_nand2_1 _3284_ (.Y(_0676_),
    .A(net222),
    .B(_0675_));
 sg13g2_o21ai_1 _3285_ (.B1(_0676_),
    .Y(_0677_),
    .A1(_0531_),
    .A2(_0572_));
 sg13g2_a22oi_1 _3286_ (.Y(_0678_),
    .B1(_0585_),
    .B2(_0677_),
    .A2(net216),
    .A1(net226));
 sg13g2_a21oi_2 _3287_ (.B1(_0674_),
    .Y(_0679_),
    .A2(_0678_),
    .A1(net220));
 sg13g2_nor2b_1 _3288_ (.A(_0679_),
    .B_N(net486),
    .Y(_0680_));
 sg13g2_xnor2_1 _3289_ (.Y(_0681_),
    .A(net486),
    .B(_0679_));
 sg13g2_nor2_1 _3290_ (.A(_0665_),
    .B(_0668_),
    .Y(_0682_));
 sg13g2_nor3_1 _3291_ (.A(_0665_),
    .B(_0668_),
    .C(_0681_),
    .Y(_0683_));
 sg13g2_nor2b_1 _3292_ (.A(_0682_),
    .B_N(_0681_),
    .Y(_0684_));
 sg13g2_nor3_1 _3293_ (.A(net205),
    .B(_0683_),
    .C(_0684_),
    .Y(_0009_));
 sg13g2_a21oi_1 _3294_ (.A1(_0507_),
    .A2(_0539_),
    .Y(_0685_),
    .B1(_0533_));
 sg13g2_o21ai_1 _3295_ (.B1(_0685_),
    .Y(_0686_),
    .A1(net243),
    .A2(_0612_));
 sg13g2_a22oi_1 _3296_ (.Y(_0687_),
    .B1(_0600_),
    .B2(_0686_),
    .A2(_0578_),
    .A1(net222));
 sg13g2_nor2_1 _3297_ (.A(net218),
    .B(_0687_),
    .Y(_0688_));
 sg13g2_o21ai_1 _3298_ (.B1(net232),
    .Y(_0689_),
    .A1(_0562_),
    .A2(_0621_));
 sg13g2_or2_1 _3299_ (.X(_0690_),
    .B(_0638_),
    .A(_0581_));
 sg13g2_a21oi_1 _3300_ (.A1(net230),
    .A2(net216),
    .Y(_0691_),
    .B1(net223));
 sg13g2_a22oi_1 _3301_ (.Y(_0692_),
    .B1(_0690_),
    .B2(_0691_),
    .A2(_0689_),
    .A1(_0670_));
 sg13g2_a21oi_2 _3302_ (.B1(_0688_),
    .Y(_0693_),
    .A2(_0692_),
    .A1(net218));
 sg13g2_xnor2_1 _3303_ (.Y(_0694_),
    .A(net470),
    .B(_0693_));
 sg13g2_or2_1 _3304_ (.X(_0695_),
    .B(_0684_),
    .A(_0680_));
 sg13g2_nor2b_1 _3305_ (.A(_0695_),
    .B_N(_0694_),
    .Y(_0696_));
 sg13g2_nor2b_1 _3306_ (.A(_0694_),
    .B_N(_0695_),
    .Y(_0697_));
 sg13g2_nor3_1 _3307_ (.A(net205),
    .B(_0696_),
    .C(_0697_),
    .Y(_0010_));
 sg13g2_a21o_1 _3308_ (.A2(_0693_),
    .A1(net470),
    .B1(_0697_),
    .X(_0698_));
 sg13g2_o21ai_1 _3309_ (.B1(_0571_),
    .Y(_0699_),
    .A1(_0561_),
    .A2(_0621_));
 sg13g2_o21ai_1 _3310_ (.B1(net223),
    .Y(_0700_),
    .A1(_0522_),
    .A2(_0610_));
 sg13g2_nand3_1 _3311_ (.B(_0699_),
    .C(_0700_),
    .A(net221),
    .Y(_0701_));
 sg13g2_a221oi_1 _3312_ (.B2(_0660_),
    .C1(net226),
    .B1(_0626_),
    .A1(net216),
    .Y(_0702_),
    .A2(_0522_));
 sg13g2_a22oi_1 _3313_ (.Y(_0703_),
    .B1(_0621_),
    .B2(_0511_),
    .A2(_0610_),
    .A1(net226));
 sg13g2_nand2_1 _3314_ (.Y(_0704_),
    .A(net218),
    .B(_0703_));
 sg13g2_o21ai_1 _3315_ (.B1(_0701_),
    .Y(_0705_),
    .A1(_0702_),
    .A2(_0704_));
 sg13g2_inv_2 _3316_ (.Y(_0706_),
    .A(_0705_));
 sg13g2_nor2_1 _3317_ (.A(_1229_),
    .B(_0706_),
    .Y(_0707_));
 sg13g2_nand2_1 _3318_ (.Y(_0708_),
    .A(_1229_),
    .B(_0706_));
 sg13g2_nor2b_1 _3319_ (.A(_0707_),
    .B_N(_0708_),
    .Y(_0709_));
 sg13g2_o21ai_1 _3320_ (.B1(net199),
    .Y(_0710_),
    .A1(_0698_),
    .A2(_0709_));
 sg13g2_a21oi_1 _3321_ (.A1(_0698_),
    .A2(_0709_),
    .Y(_0011_),
    .B1(_0710_));
 sg13g2_nand3_1 _3322_ (.B(_0570_),
    .C(_0689_),
    .A(net227),
    .Y(_0711_));
 sg13g2_a21oi_1 _3323_ (.A1(_0569_),
    .A2(_0622_),
    .Y(_0712_),
    .B1(net218));
 sg13g2_nand2_1 _3324_ (.Y(_0713_),
    .A(net232),
    .B(_0612_));
 sg13g2_a221oi_1 _3325_ (.B2(net244),
    .C1(net228),
    .B1(_0713_),
    .A1(_0521_),
    .Y(_0714_),
    .A2(net214));
 sg13g2_a221oi_1 _3326_ (.B2(_0579_),
    .C1(net223),
    .B1(net214),
    .A1(net239),
    .Y(_0715_),
    .A2(net230));
 sg13g2_nor3_1 _3327_ (.A(net221),
    .B(_0714_),
    .C(_0715_),
    .Y(_0716_));
 sg13g2_a21oi_2 _3328_ (.B1(_0716_),
    .Y(_0717_),
    .A2(_0712_),
    .A1(_0711_));
 sg13g2_inv_2 _3329_ (.Y(_0718_),
    .A(_0717_));
 sg13g2_xnor2_1 _3330_ (.Y(_0719_),
    .A(net448),
    .B(_0717_));
 sg13g2_o21ai_1 _3331_ (.B1(_0708_),
    .Y(_0720_),
    .A1(_0698_),
    .A2(_0707_));
 sg13g2_or2_1 _3332_ (.X(_0721_),
    .B(_0720_),
    .A(_0719_));
 sg13g2_nand2_1 _3333_ (.Y(_0722_),
    .A(net198),
    .B(_0721_));
 sg13g2_a21oi_1 _3334_ (.A1(_0719_),
    .A2(_0720_),
    .Y(_0012_),
    .B1(_0722_));
 sg13g2_o21ai_1 _3335_ (.B1(_0721_),
    .Y(_0723_),
    .A1(_1230_),
    .A2(_0718_));
 sg13g2_o21ai_1 _3336_ (.B1(net232),
    .Y(_0724_),
    .A1(net215),
    .A2(net213));
 sg13g2_o21ai_1 _3337_ (.B1(_0604_),
    .Y(_0725_),
    .A1(net223),
    .A2(_0612_));
 sg13g2_a21oi_1 _3338_ (.A1(_0622_),
    .A2(_0724_),
    .Y(_0726_),
    .B1(_0725_));
 sg13g2_a22oi_1 _3339_ (.Y(_0727_),
    .B1(_0535_),
    .B2(_0558_),
    .A2(_0533_),
    .A1(net233));
 sg13g2_a21oi_1 _3340_ (.A1(_0521_),
    .A2(_0533_),
    .Y(_0728_),
    .B1(_0727_));
 sg13g2_o21ai_1 _3341_ (.B1(net221),
    .Y(_0729_),
    .A1(_0512_),
    .A2(_0641_));
 sg13g2_a221oi_1 _3342_ (.B2(net223),
    .C1(_0729_),
    .B1(_0728_),
    .A1(_0514_),
    .Y(_0730_),
    .A2(_0643_));
 sg13g2_or2_1 _3343_ (.X(_0731_),
    .B(_0730_),
    .A(_0726_));
 sg13g2_inv_1 _3344_ (.Y(_0732_),
    .A(net183));
 sg13g2_nor2_1 _3345_ (.A(_1231_),
    .B(net183),
    .Y(_0733_));
 sg13g2_nand2_1 _3346_ (.Y(_0734_),
    .A(_1231_),
    .B(net183));
 sg13g2_nor2b_1 _3347_ (.A(_0733_),
    .B_N(_0734_),
    .Y(_0735_));
 sg13g2_o21ai_1 _3348_ (.B1(net200),
    .Y(_0736_),
    .A1(_0723_),
    .A2(_0735_));
 sg13g2_a21oi_1 _3349_ (.A1(_0723_),
    .A2(_0735_),
    .Y(_0013_),
    .B1(_0736_));
 sg13g2_o21ai_1 _3350_ (.B1(net219),
    .Y(_0737_),
    .A1(net224),
    .A2(_0527_));
 sg13g2_a21oi_1 _3351_ (.A1(_0545_),
    .A2(_0602_),
    .Y(_0738_),
    .B1(_0737_));
 sg13g2_o21ai_1 _3352_ (.B1(_0511_),
    .Y(_0739_),
    .A1(net214),
    .A2(net213));
 sg13g2_nand3_1 _3353_ (.B(_0532_),
    .C(_0541_),
    .A(_0516_),
    .Y(_0740_));
 sg13g2_nand3_1 _3354_ (.B(_0739_),
    .C(_0740_),
    .A(_0586_),
    .Y(_0741_));
 sg13g2_a22oi_1 _3355_ (.Y(_0742_),
    .B1(_0741_),
    .B2(net221),
    .A2(_0738_),
    .A1(_0512_));
 sg13g2_nand2_1 _3356_ (.Y(_0743_),
    .A(net450),
    .B(_0742_));
 sg13g2_xnor2_1 _3357_ (.Y(_0744_),
    .A(net450),
    .B(_0742_));
 sg13g2_o21ai_1 _3358_ (.B1(_0734_),
    .Y(_0745_),
    .A1(_0723_),
    .A2(_0733_));
 sg13g2_or2_1 _3359_ (.X(_0746_),
    .B(_0745_),
    .A(_0744_));
 sg13g2_nand2_1 _3360_ (.Y(_0747_),
    .A(net200),
    .B(_0746_));
 sg13g2_a21oi_1 _3361_ (.A1(_0744_),
    .A2(_0745_),
    .Y(_0014_),
    .B1(_0747_));
 sg13g2_nand2_1 _3362_ (.Y(_0748_),
    .A(_0743_),
    .B(_0746_));
 sg13g2_a21oi_1 _3363_ (.A1(net230),
    .A2(_0540_),
    .Y(_0749_),
    .B1(net221));
 sg13g2_o21ai_1 _3364_ (.B1(_0580_),
    .Y(_0750_),
    .A1(net234),
    .A2(_0519_));
 sg13g2_nor2_1 _3365_ (.A(net227),
    .B(_0543_),
    .Y(_0751_));
 sg13g2_a221oi_1 _3366_ (.B2(_0751_),
    .C1(net218),
    .B1(_0750_),
    .A1(_0580_),
    .Y(_0752_),
    .A2(_0691_));
 sg13g2_a21oi_2 _3367_ (.B1(_0752_),
    .Y(_0753_),
    .A2(_0749_),
    .A1(_0602_));
 sg13g2_inv_1 _3368_ (.Y(_0754_),
    .A(net186));
 sg13g2_xnor2_1 _3369_ (.Y(_0755_),
    .A(_1232_),
    .B(net186));
 sg13g2_o21ai_1 _3370_ (.B1(net200),
    .Y(_0756_),
    .A1(_0748_),
    .A2(_0755_));
 sg13g2_a21oi_1 _3371_ (.A1(_0748_),
    .A2(_0755_),
    .Y(_0015_),
    .B1(_0756_));
 sg13g2_a22oi_1 _3372_ (.Y(_0757_),
    .B1(_0541_),
    .B2(_0516_),
    .A2(_0519_),
    .A1(_0514_));
 sg13g2_nand2b_2 _3373_ (.Y(_0758_),
    .B(_0757_),
    .A_N(_0749_));
 sg13g2_nand2_1 _3374_ (.Y(_0759_),
    .A(net455),
    .B(_0758_));
 sg13g2_xnor2_1 _3375_ (.Y(_0760_),
    .A(net455),
    .B(_0758_));
 sg13g2_a21o_1 _3376_ (.A2(net186),
    .A1(\cos_x_acc[13] ),
    .B1(_0748_),
    .X(_0761_));
 sg13g2_o21ai_1 _3377_ (.B1(_0761_),
    .Y(_0762_),
    .A1(\cos_x_acc[13] ),
    .A2(net186));
 sg13g2_or2_1 _3378_ (.X(_0763_),
    .B(_0762_),
    .A(_0760_));
 sg13g2_nand2_1 _3379_ (.Y(_0764_),
    .A(net200),
    .B(_0763_));
 sg13g2_a21oi_1 _3380_ (.A1(_0760_),
    .A2(_0762_),
    .Y(_0016_),
    .B1(_0764_));
 sg13g2_nand2_1 _3381_ (.Y(_0765_),
    .A(_0759_),
    .B(_0763_));
 sg13g2_and2_1 _3382_ (.A(net221),
    .B(_0625_),
    .X(_0766_));
 sg13g2_nor2b_1 _3383_ (.A(net188),
    .B_N(net466),
    .Y(_0767_));
 sg13g2_nand2b_1 _3384_ (.Y(_0768_),
    .B(net188),
    .A_N(net466));
 sg13g2_nor2b_1 _3385_ (.A(_0767_),
    .B_N(_0768_),
    .Y(_0769_));
 sg13g2_o21ai_1 _3386_ (.B1(net201),
    .Y(_0770_),
    .A1(_0765_),
    .A2(_0769_));
 sg13g2_a21oi_1 _3387_ (.A1(_0765_),
    .A2(_0769_),
    .Y(_0017_),
    .B1(_0770_));
 sg13g2_o21ai_1 _3388_ (.B1(_0768_),
    .Y(_0771_),
    .A1(_0765_),
    .A2(_0767_));
 sg13g2_nand2b_1 _3389_ (.Y(_0772_),
    .B(_0771_),
    .A_N(net453));
 sg13g2_nand2b_1 _3390_ (.Y(_0773_),
    .B(net453),
    .A_N(_0771_));
 sg13g2_and3_1 _3391_ (.X(_0018_),
    .A(net200),
    .B(net454),
    .C(_0773_));
 sg13g2_or2_1 _3392_ (.X(_0774_),
    .B(_0773_),
    .A(_1233_));
 sg13g2_nand2_1 _3393_ (.Y(_0775_),
    .A(net200),
    .B(_0774_));
 sg13g2_a21oi_1 _3394_ (.A1(_1233_),
    .A2(_0773_),
    .Y(_0019_),
    .B1(_0775_));
 sg13g2_and2_1 _3395_ (.A(_1234_),
    .B(_0774_),
    .X(_0776_));
 sg13g2_nor2_1 _3396_ (.A(_1234_),
    .B(_0774_),
    .Y(_0777_));
 sg13g2_nor3_1 _3397_ (.A(net208),
    .B(_0776_),
    .C(_0777_),
    .Y(_0020_));
 sg13g2_nor3_2 _3398_ (.A(_1234_),
    .B(_1235_),
    .C(_0774_),
    .Y(_0778_));
 sg13g2_o21ai_1 _3399_ (.B1(net201),
    .Y(_0779_),
    .A1(net411),
    .A2(_0777_));
 sg13g2_nor2_1 _3400_ (.A(_0778_),
    .B(net412),
    .Y(_0021_));
 sg13g2_xnor2_1 _3401_ (.Y(_0780_),
    .A(net364),
    .B(_0778_));
 sg13g2_nor2_1 _3402_ (.A(net209),
    .B(net365),
    .Y(_0022_));
 sg13g2_a21oi_1 _3403_ (.A1(\cos_x_acc[20] ),
    .A2(_0778_),
    .Y(_0781_),
    .B1(net258));
 sg13g2_and3_2 _3404_ (.X(_0782_),
    .A(net364),
    .B(net258),
    .C(_0778_));
 sg13g2_nor3_1 _3405_ (.A(net209),
    .B(net259),
    .C(_0782_),
    .Y(_0023_));
 sg13g2_nor2_1 _3406_ (.A(net430),
    .B(_0782_),
    .Y(_0783_));
 sg13g2_and2_1 _3407_ (.A(net430),
    .B(_0782_),
    .X(_0784_));
 sg13g2_nor3_1 _3408_ (.A(net211),
    .B(_0783_),
    .C(_0784_),
    .Y(_0024_));
 sg13g2_o21ai_1 _3409_ (.B1(net204),
    .Y(_0785_),
    .A1(net168),
    .A2(_0784_));
 sg13g2_a21oi_1 _3410_ (.A1(net168),
    .A2(_0784_),
    .Y(_0025_),
    .B1(_0785_));
 sg13g2_a21oi_1 _3411_ (.A1(net168),
    .A2(_0784_),
    .Y(_0786_),
    .B1(net268));
 sg13g2_and4_1 _3412_ (.A(net268),
    .B(net168),
    .C(\cos_x_acc[22] ),
    .D(_0782_),
    .X(_0787_));
 sg13g2_nor3_1 _3413_ (.A(net211),
    .B(net269),
    .C(_0787_),
    .Y(_0026_));
 sg13g2_and2_1 _3414_ (.A(net390),
    .B(_0787_),
    .X(_0788_));
 sg13g2_o21ai_1 _3415_ (.B1(net204),
    .Y(_0789_),
    .A1(net390),
    .A2(_0787_));
 sg13g2_nor2_1 _3416_ (.A(_0788_),
    .B(net391),
    .Y(_0027_));
 sg13g2_a21oi_1 _3417_ (.A1(net400),
    .A2(_0788_),
    .Y(_0790_),
    .B1(net210));
 sg13g2_o21ai_1 _3418_ (.B1(_0790_),
    .Y(_0791_),
    .A1(net400),
    .A2(_0788_));
 sg13g2_inv_1 _3419_ (.Y(_0028_),
    .A(_0791_));
 sg13g2_and2_1 _3420_ (.A(net165),
    .B(net452),
    .X(_0792_));
 sg13g2_and2_1 _3421_ (.A(net377),
    .B(_0792_),
    .X(_0793_));
 sg13g2_and2_1 _3422_ (.A(net347),
    .B(_0793_),
    .X(_0794_));
 sg13g2_and2_1 _3423_ (.A(net394),
    .B(_0794_),
    .X(_0795_));
 sg13g2_nor3_1 _3424_ (.A(_1217_),
    .B(\hvsync_gen.hpos[7] ),
    .C(\hvsync_gen.hpos[6] ),
    .Y(_0796_));
 sg13g2_nand4_1 _3425_ (.B(_1242_),
    .C(_0795_),
    .A(net292),
    .Y(_0797_),
    .D(_0796_));
 sg13g2_and2_1 _3426_ (.A(net252),
    .B(_0797_),
    .X(_0798_));
 sg13g2_nand2_1 _3427_ (.Y(_0799_),
    .A(net252),
    .B(_0797_));
 sg13g2_nor2_1 _3428_ (.A(net165),
    .B(net185),
    .Y(_0029_));
 sg13g2_nor3_1 _3429_ (.A(_0553_),
    .B(_0792_),
    .C(net185),
    .Y(_0030_));
 sg13g2_nor2_1 _3430_ (.A(net377),
    .B(_0792_),
    .Y(_0800_));
 sg13g2_nor3_1 _3431_ (.A(_1248_),
    .B(_0793_),
    .C(net378),
    .Y(_0031_));
 sg13g2_o21ai_1 _3432_ (.B1(net254),
    .Y(_0801_),
    .A1(net347),
    .A2(_0793_));
 sg13g2_nor2_1 _3433_ (.A(_0794_),
    .B(net348),
    .Y(_0032_));
 sg13g2_o21ai_1 _3434_ (.B1(net254),
    .Y(_0802_),
    .A1(net394),
    .A2(_0794_));
 sg13g2_nor2_1 _3435_ (.A(_0795_),
    .B(_0802_),
    .Y(_0033_));
 sg13g2_and2_1 _3436_ (.A(net302),
    .B(_0795_),
    .X(_0803_));
 sg13g2_nor2_1 _3437_ (.A(net302),
    .B(_0795_),
    .Y(_0804_));
 sg13g2_nor3_1 _3438_ (.A(net185),
    .B(_0803_),
    .C(net303),
    .Y(_0034_));
 sg13g2_nor2_1 _3439_ (.A(net329),
    .B(_0803_),
    .Y(_0805_));
 sg13g2_and2_1 _3440_ (.A(_0493_),
    .B(_0794_),
    .X(_0806_));
 sg13g2_nor3_1 _3441_ (.A(net185),
    .B(net330),
    .C(_0806_),
    .Y(_0035_));
 sg13g2_xnor2_1 _3442_ (.Y(_0807_),
    .A(net392),
    .B(_0806_));
 sg13g2_nor2_1 _3443_ (.A(net185),
    .B(net393),
    .Y(_0036_));
 sg13g2_a21oi_1 _3444_ (.A1(\hvsync_gen.hpos[7] ),
    .A2(_0806_),
    .Y(_0808_),
    .B1(net273));
 sg13g2_and3_1 _3445_ (.X(_0809_),
    .A(net273),
    .B(net392),
    .C(_0806_));
 sg13g2_nor3_1 _3446_ (.A(net185),
    .B(net274),
    .C(_0809_),
    .Y(_0037_));
 sg13g2_a21oi_1 _3447_ (.A1(net292),
    .A2(_0809_),
    .Y(_0810_),
    .B1(net185));
 sg13g2_o21ai_1 _3448_ (.B1(_0810_),
    .Y(_0811_),
    .A1(net292),
    .A2(_0809_));
 sg13g2_inv_1 _3449_ (.Y(_0038_),
    .A(_0811_));
 sg13g2_nor3_1 _3450_ (.A(\bayer_j[0] ),
    .B(net246),
    .C(net305),
    .Y(_0812_));
 sg13g2_nor4_1 _3451_ (.A(\hvsync_gen.vpos[4] ),
    .B(\hvsync_gen.vpos[5] ),
    .C(\hvsync_gen.vpos[6] ),
    .D(net285),
    .Y(_0813_));
 sg13g2_nor3_1 _3452_ (.A(\hvsync_gen.vpos[9] ),
    .B(\hvsync_gen.vpos[2] ),
    .C(net332),
    .Y(_0814_));
 sg13g2_nand3_1 _3453_ (.B(_0813_),
    .C(_0814_),
    .A(_0812_),
    .Y(_0815_));
 sg13g2_nand2b_1 _3454_ (.Y(_0816_),
    .B(\y_prv[3] ),
    .A_N(\hvsync_gen.vpos[3] ));
 sg13g2_xnor2_1 _3455_ (.Y(_0817_),
    .A(\hvsync_gen.vpos[4] ),
    .B(\y_prv[4] ));
 sg13g2_nand2b_1 _3456_ (.Y(_0818_),
    .B(\hvsync_gen.vpos[5] ),
    .A_N(\y_prv[5] ));
 sg13g2_nand2b_1 _3457_ (.Y(_0819_),
    .B(\hvsync_gen.vpos[2] ),
    .A_N(\y_prv[2] ));
 sg13g2_xnor2_1 _3458_ (.Y(_0820_),
    .A(\hvsync_gen.vpos[9] ),
    .B(\y_prv[9] ));
 sg13g2_nand4_1 _3459_ (.B(_0818_),
    .C(_0819_),
    .A(_0817_),
    .Y(_0821_),
    .D(_0820_));
 sg13g2_a221oi_1 _3460_ (.B2(net322),
    .C1(_0821_),
    .B1(_1246_),
    .A1(_1215_),
    .Y(_0822_),
    .A2(net266));
 sg13g2_a22oi_1 _3461_ (.Y(_0823_),
    .B1(\y_prv[5] ),
    .B2(_1238_),
    .A2(_1243_),
    .A1(\bayer_j[0] ));
 sg13g2_o21ai_1 _3462_ (.B1(_0816_),
    .Y(_0824_),
    .A1(_1240_),
    .A2(\y_prv[7] ));
 sg13g2_a22oi_1 _3463_ (.Y(_0825_),
    .B1(_1247_),
    .B2(\hvsync_gen.vpos[8] ),
    .A2(_1244_),
    .A1(\bayer_j[1] ));
 sg13g2_a221oi_1 _3464_ (.B2(\hvsync_gen.vpos[3] ),
    .C1(_0824_),
    .B1(_1245_),
    .A1(_1237_),
    .Y(_0826_),
    .A2(\y_prv[2] ));
 sg13g2_a22oi_1 _3465_ (.Y(_0827_),
    .B1(\y_prv[8] ),
    .B2(_1241_),
    .A2(\y_prv[1] ),
    .A1(_1216_));
 sg13g2_nand4_1 _3466_ (.B(_0825_),
    .C(_0826_),
    .A(_0823_),
    .Y(_0828_),
    .D(_0827_));
 sg13g2_a221oi_1 _3467_ (.B2(_1240_),
    .C1(_0828_),
    .B1(net261),
    .A1(_1239_),
    .Y(_0829_),
    .A2(\y_prv[6] ));
 sg13g2_a21oi_1 _3468_ (.A1(_0822_),
    .A2(_0829_),
    .Y(_0830_),
    .B1(_0815_));
 sg13g2_nor2_1 _3469_ (.A(net251),
    .B(_0830_),
    .Y(_0831_));
 sg13g2_and2_1 _3470_ (.A(net467),
    .B(_0830_),
    .X(_0832_));
 sg13g2_nor3_1 _3471_ (.A(_1248_),
    .B(_0831_),
    .C(_0832_),
    .Y(_0039_));
 sg13g2_o21ai_1 _3472_ (.B1(net254),
    .Y(_0833_),
    .A1(net311),
    .A2(_0832_));
 sg13g2_a21oi_1 _3473_ (.A1(net311),
    .A2(_0832_),
    .Y(_0040_),
    .B1(_0833_));
 sg13g2_a21oi_1 _3474_ (.A1(\cos_addr[1] ),
    .A2(_0832_),
    .Y(_0834_),
    .B1(net282));
 sg13g2_and3_1 _3475_ (.X(_0835_),
    .A(net282),
    .B(net311),
    .C(_0832_));
 sg13g2_nor3_1 _3476_ (.A(_1248_),
    .B(net283),
    .C(_0835_),
    .Y(_0041_));
 sg13g2_and2_1 _3477_ (.A(net440),
    .B(_0835_),
    .X(_0836_));
 sg13g2_o21ai_1 _3478_ (.B1(net254),
    .Y(_0837_),
    .A1(net440),
    .A2(_0835_));
 sg13g2_nor2_1 _3479_ (.A(_0836_),
    .B(_0837_),
    .Y(_0042_));
 sg13g2_and2_1 _3480_ (.A(net402),
    .B(_0836_),
    .X(_0838_));
 sg13g2_o21ai_1 _3481_ (.B1(net254),
    .Y(_0839_),
    .A1(net402),
    .A2(_0836_));
 sg13g2_nor2_1 _3482_ (.A(_0838_),
    .B(net403),
    .Y(_0043_));
 sg13g2_and2_1 _3483_ (.A(net416),
    .B(_0838_),
    .X(_0840_));
 sg13g2_o21ai_1 _3484_ (.B1(net254),
    .Y(_0841_),
    .A1(net416),
    .A2(_0838_));
 sg13g2_nor2_1 _3485_ (.A(_0840_),
    .B(_0841_),
    .Y(_0044_));
 sg13g2_o21ai_1 _3486_ (.B1(net254),
    .Y(_0842_),
    .A1(net166),
    .A2(_0840_));
 sg13g2_a21oi_1 _3487_ (.A1(net166),
    .A2(_0840_),
    .Y(_0045_),
    .B1(_0842_));
 sg13g2_nor2_1 _3488_ (.A(net266),
    .B(net252),
    .Y(_0843_));
 sg13g2_a21oi_1 _3489_ (.A1(_1215_),
    .A2(net252),
    .Y(_0046_),
    .B1(_0843_));
 sg13g2_mux2_1 _3490_ (.A0(net313),
    .A1(\bayer_j[1] ),
    .S(net253),
    .X(_0047_));
 sg13g2_mux2_1 _3491_ (.A0(net315),
    .A1(net309),
    .S(net253),
    .X(_0048_));
 sg13g2_mux2_1 _3492_ (.A0(net320),
    .A1(\hvsync_gen.vpos[3] ),
    .S(net253),
    .X(_0049_));
 sg13g2_mux2_1 _3493_ (.A0(net291),
    .A1(net271),
    .S(net1),
    .X(_0050_));
 sg13g2_nor2_1 _3494_ (.A(net256),
    .B(net253),
    .Y(_0844_));
 sg13g2_a21oi_1 _3495_ (.A1(_1238_),
    .A2(net252),
    .Y(_0051_),
    .B1(_0844_));
 sg13g2_nand2_1 _3496_ (.Y(_0845_),
    .A(\hvsync_gen.vpos[6] ),
    .B(net252));
 sg13g2_o21ai_1 _3497_ (.B1(_0845_),
    .Y(_0052_),
    .A1(_1246_),
    .A2(net252));
 sg13g2_nor2_1 _3498_ (.A(net261),
    .B(net252),
    .Y(_0846_));
 sg13g2_a21oi_1 _3499_ (.A1(_1240_),
    .A2(net253),
    .Y(_0053_),
    .B1(_0846_));
 sg13g2_mux2_1 _3500_ (.A0(net308),
    .A1(net305),
    .S(net253),
    .X(_0054_));
 sg13g2_mux2_1 _3501_ (.A0(net316),
    .A1(\hvsync_gen.vpos[9] ),
    .S(net1),
    .X(_0055_));
 sg13g2_or2_1 _3502_ (.X(_0847_),
    .B(net187),
    .A(net370));
 sg13g2_nand2_1 _3503_ (.Y(_0848_),
    .A(net370),
    .B(net187));
 sg13g2_and3_1 _3504_ (.X(_0056_),
    .A(net203),
    .B(_0847_),
    .C(_0848_));
 sg13g2_nor2_2 _3505_ (.A(net187),
    .B(_0574_),
    .Y(_0849_));
 sg13g2_xor2_1 _3506_ (.B(_0574_),
    .A(net187),
    .X(_0850_));
 sg13g2_nand2_1 _3507_ (.Y(_0851_),
    .A(net478),
    .B(_0850_));
 sg13g2_xnor2_1 _3508_ (.Y(_0852_),
    .A(\sin_x_acc[1] ),
    .B(_0850_));
 sg13g2_or2_1 _3509_ (.X(_0853_),
    .B(_0852_),
    .A(_0848_));
 sg13g2_nand2_1 _3510_ (.Y(_0854_),
    .A(net203),
    .B(_0853_));
 sg13g2_a21oi_1 _3511_ (.A1(_0848_),
    .A2(_0852_),
    .Y(_0057_),
    .B1(_0854_));
 sg13g2_nand2_1 _3512_ (.Y(_0855_),
    .A(_0594_),
    .B(_0849_));
 sg13g2_xor2_1 _3513_ (.B(_0849_),
    .A(_0594_),
    .X(_0856_));
 sg13g2_xnor2_1 _3514_ (.Y(_0857_),
    .A(\sin_x_acc[2] ),
    .B(_0856_));
 sg13g2_and3_1 _3515_ (.X(_0858_),
    .A(_0851_),
    .B(_0853_),
    .C(_0857_));
 sg13g2_a21oi_1 _3516_ (.A1(_0851_),
    .A2(_0853_),
    .Y(_0859_),
    .B1(_0857_));
 sg13g2_nor3_1 _3517_ (.A(net211),
    .B(net479),
    .C(_0859_),
    .Y(_0058_));
 sg13g2_a21oi_1 _3518_ (.A1(\sin_x_acc[2] ),
    .A2(_0856_),
    .Y(_0860_),
    .B1(_0859_));
 sg13g2_nand3_1 _3519_ (.B(_0615_),
    .C(_0849_),
    .A(_0594_),
    .Y(_0861_));
 sg13g2_xnor2_1 _3520_ (.Y(_0862_),
    .A(_0615_),
    .B(_0855_));
 sg13g2_nand2_1 _3521_ (.Y(_0863_),
    .A(net476),
    .B(_0862_));
 sg13g2_xnor2_1 _3522_ (.Y(_0864_),
    .A(net476),
    .B(_0862_));
 sg13g2_o21ai_1 _3523_ (.B1(net203),
    .Y(_0865_),
    .A1(_0860_),
    .A2(_0864_));
 sg13g2_a21oi_1 _3524_ (.A1(_0860_),
    .A2(_0864_),
    .Y(_0059_),
    .B1(_0865_));
 sg13g2_o21ai_1 _3525_ (.B1(_0863_),
    .Y(_0866_),
    .A1(_0860_),
    .A2(_0864_));
 sg13g2_nand4_1 _3526_ (.B(_0615_),
    .C(_0633_),
    .A(_0594_),
    .Y(_0867_),
    .D(_0849_));
 sg13g2_xnor2_1 _3527_ (.Y(_0868_),
    .A(_0633_),
    .B(_0861_));
 sg13g2_xnor2_1 _3528_ (.Y(_0869_),
    .A(net495),
    .B(_0868_));
 sg13g2_nor2b_1 _3529_ (.A(_0866_),
    .B_N(_0869_),
    .Y(_0870_));
 sg13g2_nor2b_1 _3530_ (.A(_0869_),
    .B_N(_0866_),
    .Y(_0871_));
 sg13g2_nor3_1 _3531_ (.A(net207),
    .B(_0870_),
    .C(_0871_),
    .Y(_0060_));
 sg13g2_a21oi_1 _3532_ (.A1(\sin_x_acc[4] ),
    .A2(_0868_),
    .Y(_0872_),
    .B1(_0871_));
 sg13g2_xnor2_1 _3533_ (.Y(_0873_),
    .A(_0650_),
    .B(_0867_));
 sg13g2_nand2_1 _3534_ (.Y(_0874_),
    .A(net460),
    .B(_0873_));
 sg13g2_xnor2_1 _3535_ (.Y(_0875_),
    .A(net460),
    .B(_0873_));
 sg13g2_or2_1 _3536_ (.X(_0876_),
    .B(_0875_),
    .A(_0872_));
 sg13g2_nand2_1 _3537_ (.Y(_0877_),
    .A(net199),
    .B(_0876_));
 sg13g2_a21oi_1 _3538_ (.A1(_0872_),
    .A2(_0875_),
    .Y(_0061_),
    .B1(_0877_));
 sg13g2_o21ai_1 _3539_ (.B1(_0664_),
    .Y(_0878_),
    .A1(_0651_),
    .A2(_0867_));
 sg13g2_xnor2_1 _3540_ (.Y(_0879_),
    .A(net488),
    .B(_0878_));
 sg13g2_and3_1 _3541_ (.X(_0880_),
    .A(_0874_),
    .B(_0876_),
    .C(_0879_));
 sg13g2_a21oi_1 _3542_ (.A1(_0874_),
    .A2(_0876_),
    .Y(_0881_),
    .B1(_0879_));
 sg13g2_nor3_1 _3543_ (.A(net205),
    .B(_0880_),
    .C(_0881_),
    .Y(_0062_));
 sg13g2_xnor2_1 _3544_ (.Y(_0882_),
    .A(net498),
    .B(_0679_));
 sg13g2_a21oi_1 _3545_ (.A1(net488),
    .A2(_0878_),
    .Y(_0883_),
    .B1(_0881_));
 sg13g2_nor2_1 _3546_ (.A(_0882_),
    .B(_0883_),
    .Y(_0884_));
 sg13g2_a21oi_1 _3547_ (.A1(_0882_),
    .A2(_0883_),
    .Y(_0885_),
    .B1(net205));
 sg13g2_nor2b_1 _3548_ (.A(_0884_),
    .B_N(_0885_),
    .Y(_0063_));
 sg13g2_nor2b_1 _3549_ (.A(_0693_),
    .B_N(\sin_x_acc[8] ),
    .Y(_0886_));
 sg13g2_xnor2_1 _3550_ (.Y(_0887_),
    .A(net497),
    .B(_0693_));
 sg13g2_a21o_1 _3551_ (.A2(_0679_),
    .A1(net498),
    .B1(_0884_),
    .X(_0888_));
 sg13g2_or2_1 _3552_ (.X(_0889_),
    .B(_0888_),
    .A(_0887_));
 sg13g2_nand2_1 _3553_ (.Y(_0890_),
    .A(_0887_),
    .B(_0888_));
 sg13g2_and3_1 _3554_ (.X(_0064_),
    .A(net198),
    .B(_0889_),
    .C(_0890_));
 sg13g2_a21oi_1 _3555_ (.A1(_0887_),
    .A2(_0888_),
    .Y(_0891_),
    .B1(_0886_));
 sg13g2_nand2_1 _3556_ (.Y(_0892_),
    .A(net472),
    .B(_0706_));
 sg13g2_nor2_1 _3557_ (.A(net472),
    .B(_0706_),
    .Y(_0893_));
 sg13g2_xor2_1 _3558_ (.B(_0705_),
    .A(net472),
    .X(_0894_));
 sg13g2_o21ai_1 _3559_ (.B1(net198),
    .Y(_0895_),
    .A1(_0891_),
    .A2(_0894_));
 sg13g2_a21oi_1 _3560_ (.A1(_0891_),
    .A2(_0894_),
    .Y(_0065_),
    .B1(_0895_));
 sg13g2_xnor2_1 _3561_ (.Y(_0896_),
    .A(net493),
    .B(_0717_));
 sg13g2_a21oi_1 _3562_ (.A1(_0891_),
    .A2(_0892_),
    .Y(_0897_),
    .B1(_0893_));
 sg13g2_nor2_1 _3563_ (.A(_0896_),
    .B(_0897_),
    .Y(_0898_));
 sg13g2_and2_1 _3564_ (.A(_0896_),
    .B(_0897_),
    .X(_0899_));
 sg13g2_nor3_1 _3565_ (.A(net205),
    .B(_0898_),
    .C(_0899_),
    .Y(_0066_));
 sg13g2_a21o_1 _3566_ (.A2(_0718_),
    .A1(net493),
    .B1(_0899_),
    .X(_0900_));
 sg13g2_and2_1 _3567_ (.A(\sin_x_acc[11] ),
    .B(net183),
    .X(_0901_));
 sg13g2_or2_1 _3568_ (.X(_0902_),
    .B(net183),
    .A(\sin_x_acc[11] ));
 sg13g2_nor2b_1 _3569_ (.A(_0901_),
    .B_N(_0902_),
    .Y(_0903_));
 sg13g2_o21ai_1 _3570_ (.B1(net200),
    .Y(_0904_),
    .A1(_0900_),
    .A2(_0903_));
 sg13g2_a21oi_1 _3571_ (.A1(_0900_),
    .A2(_0903_),
    .Y(_0067_),
    .B1(_0904_));
 sg13g2_xnor2_1 _3572_ (.Y(_0905_),
    .A(_1227_),
    .B(_0742_));
 sg13g2_o21ai_1 _3573_ (.B1(_0902_),
    .Y(_0906_),
    .A1(_0900_),
    .A2(_0901_));
 sg13g2_or2_1 _3574_ (.X(_0907_),
    .B(_0906_),
    .A(_0905_));
 sg13g2_nand2_1 _3575_ (.Y(_0908_),
    .A(net201),
    .B(_0907_));
 sg13g2_a21oi_1 _3576_ (.A1(_0905_),
    .A2(_0906_),
    .Y(_0068_),
    .B1(_0908_));
 sg13g2_o21ai_1 _3577_ (.B1(_0907_),
    .Y(_0909_),
    .A1(_1227_),
    .A2(_0742_));
 sg13g2_nor2b_1 _3578_ (.A(net186),
    .B_N(net500),
    .Y(_0910_));
 sg13g2_nand2b_1 _3579_ (.Y(_0911_),
    .B(net186),
    .A_N(net500));
 sg13g2_nor2b_1 _3580_ (.A(_0910_),
    .B_N(_0911_),
    .Y(_0912_));
 sg13g2_o21ai_1 _3581_ (.B1(net201),
    .Y(_0913_),
    .A1(_0909_),
    .A2(_0912_));
 sg13g2_a21oi_1 _3582_ (.A1(_0909_),
    .A2(_0912_),
    .Y(_0069_),
    .B1(_0913_));
 sg13g2_xnor2_1 _3583_ (.Y(_0914_),
    .A(_1214_),
    .B(_0758_));
 sg13g2_o21ai_1 _3584_ (.B1(_0911_),
    .Y(_0915_),
    .A1(_0909_),
    .A2(_0910_));
 sg13g2_or2_1 _3585_ (.X(_0916_),
    .B(_0915_),
    .A(_0914_));
 sg13g2_nand2_1 _3586_ (.Y(_0917_),
    .A(net201),
    .B(_0916_));
 sg13g2_a21oi_1 _3587_ (.A1(_0914_),
    .A2(_0915_),
    .Y(_0070_),
    .B1(_0917_));
 sg13g2_o21ai_1 _3588_ (.B1(_0916_),
    .Y(_0918_),
    .A1(_1214_),
    .A2(_0758_));
 sg13g2_and2_1 _3589_ (.A(net502),
    .B(net188),
    .X(_0919_));
 sg13g2_or2_1 _3590_ (.X(_0920_),
    .B(net188),
    .A(net502));
 sg13g2_nor2b_1 _3591_ (.A(_0919_),
    .B_N(_0920_),
    .Y(_0921_));
 sg13g2_o21ai_1 _3592_ (.B1(net202),
    .Y(_0922_),
    .A1(_0918_),
    .A2(_0921_));
 sg13g2_a21oi_1 _3593_ (.A1(_0918_),
    .A2(_0921_),
    .Y(_0071_),
    .B1(_0922_));
 sg13g2_o21ai_1 _3594_ (.B1(_0920_),
    .Y(_0923_),
    .A1(_0918_),
    .A2(_0919_));
 sg13g2_nand2b_1 _3595_ (.Y(_0924_),
    .B(_0923_),
    .A_N(net465));
 sg13g2_nand2b_2 _3596_ (.Y(_0925_),
    .B(net465),
    .A_N(_0923_));
 sg13g2_and3_1 _3597_ (.X(_0072_),
    .A(net201),
    .B(_0924_),
    .C(_0925_));
 sg13g2_or2_1 _3598_ (.X(_0926_),
    .B(_0925_),
    .A(_1220_));
 sg13g2_nand2_1 _3599_ (.Y(_0927_),
    .A(net204),
    .B(_0926_));
 sg13g2_a21oi_1 _3600_ (.A1(_1220_),
    .A2(_0925_),
    .Y(_0073_),
    .B1(_0927_));
 sg13g2_and2_1 _3601_ (.A(_1219_),
    .B(_0926_),
    .X(_0928_));
 sg13g2_nor2_1 _3602_ (.A(_1219_),
    .B(_0926_),
    .Y(_0929_));
 sg13g2_nor3_1 _3603_ (.A(net210),
    .B(_0928_),
    .C(_0929_),
    .Y(_0074_));
 sg13g2_nor3_2 _3604_ (.A(_1218_),
    .B(_1219_),
    .C(_0926_),
    .Y(_0930_));
 sg13g2_o21ai_1 _3605_ (.B1(net204),
    .Y(_0931_),
    .A1(net436),
    .A2(_0929_));
 sg13g2_nor2_1 _3606_ (.A(_0930_),
    .B(net437),
    .Y(_0075_));
 sg13g2_xnor2_1 _3607_ (.Y(_0932_),
    .A(net441),
    .B(_0930_));
 sg13g2_nor2_1 _3608_ (.A(net210),
    .B(net442),
    .Y(_0076_));
 sg13g2_a21oi_1 _3609_ (.A1(\sin_x_acc[20] ),
    .A2(_0930_),
    .Y(_0933_),
    .B1(net326));
 sg13g2_and3_2 _3610_ (.X(_0934_),
    .A(net326),
    .B(\sin_x_acc[20] ),
    .C(_0930_));
 sg13g2_nor3_1 _3611_ (.A(net210),
    .B(net327),
    .C(_0934_),
    .Y(_0077_));
 sg13g2_xnor2_1 _3612_ (.Y(_0935_),
    .A(net428),
    .B(_0934_));
 sg13g2_nor2_1 _3613_ (.A(net210),
    .B(net429),
    .Y(_0078_));
 sg13g2_a21oi_1 _3614_ (.A1(\sin_x_acc[22] ),
    .A2(_0934_),
    .Y(_0936_),
    .B1(net299));
 sg13g2_and3_1 _3615_ (.X(_0937_),
    .A(net299),
    .B(\sin_x_acc[22] ),
    .C(_0934_));
 sg13g2_nor3_1 _3616_ (.A(net210),
    .B(net300),
    .C(_0937_),
    .Y(_0079_));
 sg13g2_nor2_1 _3617_ (.A(net356),
    .B(_0937_),
    .Y(_0938_));
 sg13g2_and2_1 _3618_ (.A(net356),
    .B(_0937_),
    .X(_0939_));
 sg13g2_nor3_1 _3619_ (.A(net210),
    .B(net357),
    .C(_0939_),
    .Y(_0080_));
 sg13g2_and2_1 _3620_ (.A(net421),
    .B(_0939_),
    .X(_0940_));
 sg13g2_o21ai_1 _3621_ (.B1(net204),
    .Y(_0941_),
    .A1(net421),
    .A2(_0939_));
 sg13g2_nor2_1 _3622_ (.A(_0940_),
    .B(_0941_),
    .Y(_0081_));
 sg13g2_nor2_1 _3623_ (.A(net288),
    .B(_0940_),
    .Y(_0942_));
 sg13g2_a21oi_1 _3624_ (.A1(net288),
    .A2(_0940_),
    .Y(_0943_),
    .B1(net210));
 sg13g2_nor2b_1 _3625_ (.A(net289),
    .B_N(_0943_),
    .Y(_0082_));
 sg13g2_nor2_1 _3626_ (.A(net204),
    .B(_0815_),
    .Y(_0944_));
 sg13g2_and2_1 _3627_ (.A(_0550_),
    .B(net211),
    .X(_0945_));
 sg13g2_xnor2_1 _3628_ (.Y(_0946_),
    .A(net388),
    .B(_0945_));
 sg13g2_nor2_1 _3629_ (.A(net197),
    .B(_0946_),
    .Y(_0083_));
 sg13g2_nand2_1 _3630_ (.Y(_0947_),
    .A(\sin_y_acc[0] ),
    .B(net187));
 sg13g2_nand2_1 _3631_ (.Y(_0948_),
    .A(net358),
    .B(_0850_));
 sg13g2_xnor2_1 _3632_ (.Y(_0949_),
    .A(net358),
    .B(_0850_));
 sg13g2_and2_1 _3633_ (.A(net211),
    .B(_0815_),
    .X(_0950_));
 sg13g2_o21ai_1 _3634_ (.B1(net192),
    .Y(_0951_),
    .A1(_0947_),
    .A2(_0949_));
 sg13g2_a21oi_1 _3635_ (.A1(_0947_),
    .A2(_0949_),
    .Y(_0952_),
    .B1(_0951_));
 sg13g2_a21o_1 _3636_ (.A2(net203),
    .A1(net358),
    .B1(_0952_),
    .X(_0084_));
 sg13g2_o21ai_1 _3637_ (.B1(_0948_),
    .Y(_0953_),
    .A1(_0947_),
    .A2(_0949_));
 sg13g2_nand2_1 _3638_ (.Y(_0954_),
    .A(\sin_y_acc[2] ),
    .B(_0856_));
 sg13g2_xnor2_1 _3639_ (.Y(_0955_),
    .A(net423),
    .B(_0856_));
 sg13g2_nand2b_1 _3640_ (.Y(_0956_),
    .B(_0953_),
    .A_N(_0955_));
 sg13g2_nand2b_1 _3641_ (.Y(_0957_),
    .B(_0955_),
    .A_N(_0953_));
 sg13g2_nand3_1 _3642_ (.B(_0956_),
    .C(_0957_),
    .A(net192),
    .Y(_0958_));
 sg13g2_o21ai_1 _3643_ (.B1(_0958_),
    .Y(_0085_),
    .A1(_1212_),
    .A2(net211));
 sg13g2_nand2_1 _3644_ (.Y(_0959_),
    .A(net278),
    .B(net203));
 sg13g2_nand2_1 _3645_ (.Y(_0960_),
    .A(_0954_),
    .B(_0956_));
 sg13g2_xnor2_1 _3646_ (.Y(_0961_),
    .A(net278),
    .B(_0862_));
 sg13g2_inv_1 _3647_ (.Y(_0962_),
    .A(_0961_));
 sg13g2_a21oi_1 _3648_ (.A1(_0954_),
    .A2(_0956_),
    .Y(_0963_),
    .B1(_0961_));
 sg13g2_o21ai_1 _3649_ (.B1(net192),
    .Y(_0964_),
    .A1(_0960_),
    .A2(_0962_));
 sg13g2_o21ai_1 _3650_ (.B1(_0959_),
    .Y(_0086_),
    .A1(_0963_),
    .A2(_0964_));
 sg13g2_nand2_1 _3651_ (.Y(_0965_),
    .A(net287),
    .B(net199));
 sg13g2_a21o_1 _3652_ (.A2(_0862_),
    .A1(net278),
    .B1(_0963_),
    .X(_0966_));
 sg13g2_xnor2_1 _3653_ (.Y(_0967_),
    .A(net287),
    .B(_0868_));
 sg13g2_inv_1 _3654_ (.Y(_0968_),
    .A(_0967_));
 sg13g2_and2_1 _3655_ (.A(_0966_),
    .B(_0968_),
    .X(_0969_));
 sg13g2_o21ai_1 _3656_ (.B1(net192),
    .Y(_0970_),
    .A1(_0966_),
    .A2(_0968_));
 sg13g2_o21ai_1 _3657_ (.B1(_0965_),
    .Y(_0087_),
    .A1(_0969_),
    .A2(_0970_));
 sg13g2_a21oi_1 _3658_ (.A1(net287),
    .A2(_0868_),
    .Y(_0971_),
    .B1(_0969_));
 sg13g2_nand2_1 _3659_ (.Y(_0972_),
    .A(\sin_y_acc[5] ),
    .B(_0873_));
 sg13g2_xnor2_1 _3660_ (.Y(_0973_),
    .A(net360),
    .B(_0873_));
 sg13g2_or2_1 _3661_ (.X(_0974_),
    .B(_0973_),
    .A(_0971_));
 sg13g2_nand2_1 _3662_ (.Y(_0975_),
    .A(net189),
    .B(_0974_));
 sg13g2_a21oi_1 _3663_ (.A1(_0971_),
    .A2(_0973_),
    .Y(_0976_),
    .B1(_0975_));
 sg13g2_a21o_1 _3664_ (.A2(net198),
    .A1(net360),
    .B1(_0976_),
    .X(_0088_));
 sg13g2_nand2_1 _3665_ (.Y(_0977_),
    .A(net295),
    .B(net198));
 sg13g2_xnor2_1 _3666_ (.Y(_0978_),
    .A(net295),
    .B(_0878_));
 sg13g2_a21oi_1 _3667_ (.A1(_0972_),
    .A2(_0974_),
    .Y(_0979_),
    .B1(_0978_));
 sg13g2_nand3_1 _3668_ (.B(_0974_),
    .C(_0978_),
    .A(_0972_),
    .Y(_0980_));
 sg13g2_nand2_1 _3669_ (.Y(_0981_),
    .A(net189),
    .B(_0980_));
 sg13g2_o21ai_1 _3670_ (.B1(_0977_),
    .Y(_0089_),
    .A1(_0979_),
    .A2(_0981_));
 sg13g2_xnor2_1 _3671_ (.Y(_0982_),
    .A(net369),
    .B(_0679_));
 sg13g2_a21oi_1 _3672_ (.A1(net295),
    .A2(_0878_),
    .Y(_0983_),
    .B1(_0979_));
 sg13g2_nor2_1 _3673_ (.A(_0982_),
    .B(_0983_),
    .Y(_0984_));
 sg13g2_o21ai_1 _3674_ (.B1(net189),
    .Y(_0985_),
    .A1(_0982_),
    .A2(_0983_));
 sg13g2_a21oi_1 _3675_ (.A1(_0982_),
    .A2(_0983_),
    .Y(_0986_),
    .B1(_0985_));
 sg13g2_a21o_1 _3676_ (.A2(net198),
    .A1(net369),
    .B1(_0986_),
    .X(_0090_));
 sg13g2_nor2b_1 _3677_ (.A(_0693_),
    .B_N(\sin_y_acc[8] ),
    .Y(_0987_));
 sg13g2_xnor2_1 _3678_ (.Y(_0988_),
    .A(net366),
    .B(_0693_));
 sg13g2_a21o_1 _3679_ (.A2(_0679_),
    .A1(\sin_y_acc[7] ),
    .B1(_0984_),
    .X(_0989_));
 sg13g2_o21ai_1 _3680_ (.B1(net189),
    .Y(_0990_),
    .A1(_0988_),
    .A2(_0989_));
 sg13g2_a21oi_1 _3681_ (.A1(_0988_),
    .A2(_0989_),
    .Y(_0991_),
    .B1(_0990_));
 sg13g2_a21o_1 _3682_ (.A2(net199),
    .A1(net366),
    .B1(_0991_),
    .X(_0091_));
 sg13g2_a21oi_1 _3683_ (.A1(_0988_),
    .A2(_0989_),
    .Y(_0992_),
    .B1(_0987_));
 sg13g2_xnor2_1 _3684_ (.Y(_0993_),
    .A(_1211_),
    .B(_0705_));
 sg13g2_o21ai_1 _3685_ (.B1(net189),
    .Y(_0994_),
    .A1(_0992_),
    .A2(_0993_));
 sg13g2_a21o_1 _3686_ (.A2(_0993_),
    .A1(_0992_),
    .B1(_0994_),
    .X(_0995_));
 sg13g2_o21ai_1 _3687_ (.B1(_0995_),
    .Y(_0092_),
    .A1(_1211_),
    .A2(net206));
 sg13g2_nand2_1 _3688_ (.Y(_0996_),
    .A(net280),
    .B(net198));
 sg13g2_xnor2_1 _3689_ (.Y(_0997_),
    .A(net280),
    .B(_0717_));
 sg13g2_a21oi_1 _3690_ (.A1(_1211_),
    .A2(_0705_),
    .Y(_0998_),
    .B1(_0992_));
 sg13g2_a21o_1 _3691_ (.A2(_0706_),
    .A1(\sin_y_acc[9] ),
    .B1(_0998_),
    .X(_0999_));
 sg13g2_and2_1 _3692_ (.A(_0997_),
    .B(_0999_),
    .X(_1000_));
 sg13g2_o21ai_1 _3693_ (.B1(net190),
    .Y(_1001_),
    .A1(_0997_),
    .A2(_0999_));
 sg13g2_o21ai_1 _3694_ (.B1(_0996_),
    .Y(_0093_),
    .A1(_1000_),
    .A2(_1001_));
 sg13g2_a21oi_1 _3695_ (.A1(net280),
    .A2(_0718_),
    .Y(_1002_),
    .B1(_1000_));
 sg13g2_nand2_1 _3696_ (.Y(_1003_),
    .A(\sin_y_acc[11] ),
    .B(net183));
 sg13g2_nor2_1 _3697_ (.A(net368),
    .B(net183),
    .Y(_1004_));
 sg13g2_xnor2_1 _3698_ (.Y(_1005_),
    .A(net368),
    .B(net183));
 sg13g2_o21ai_1 _3699_ (.B1(net190),
    .Y(_1006_),
    .A1(_1002_),
    .A2(_1005_));
 sg13g2_a21oi_1 _3700_ (.A1(_1002_),
    .A2(_1005_),
    .Y(_1007_),
    .B1(_1006_));
 sg13g2_a21o_1 _3701_ (.A2(net200),
    .A1(net368),
    .B1(_1007_),
    .X(_0094_));
 sg13g2_xnor2_1 _3702_ (.Y(_1008_),
    .A(net373),
    .B(_0742_));
 sg13g2_a21oi_1 _3703_ (.A1(_1002_),
    .A2(_1003_),
    .Y(_1009_),
    .B1(_1004_));
 sg13g2_nand2_1 _3704_ (.Y(_1010_),
    .A(_1008_),
    .B(_1009_));
 sg13g2_o21ai_1 _3705_ (.B1(net190),
    .Y(_1011_),
    .A1(_1008_),
    .A2(_1009_));
 sg13g2_nand2b_1 _3706_ (.Y(_1012_),
    .B(_1010_),
    .A_N(_1011_));
 sg13g2_o21ai_1 _3707_ (.B1(_1012_),
    .Y(_0095_),
    .A1(_1210_),
    .A2(net208));
 sg13g2_o21ai_1 _3708_ (.B1(_1010_),
    .Y(_1013_),
    .A1(_1210_),
    .A2(_0742_));
 sg13g2_xnor2_1 _3709_ (.Y(_1014_),
    .A(net446),
    .B(net186));
 sg13g2_o21ai_1 _3710_ (.B1(net190),
    .Y(_1015_),
    .A1(_1013_),
    .A2(_1014_));
 sg13g2_a21o_1 _3711_ (.A2(_1014_),
    .A1(_1013_),
    .B1(_1015_),
    .X(_1016_));
 sg13g2_o21ai_1 _3712_ (.B1(_1016_),
    .Y(_0096_),
    .A1(_1209_),
    .A2(net208));
 sg13g2_xnor2_1 _3713_ (.Y(_1017_),
    .A(_1208_),
    .B(_0758_));
 sg13g2_o21ai_1 _3714_ (.B1(_1013_),
    .Y(_1018_),
    .A1(net504),
    .A2(_0754_));
 sg13g2_o21ai_1 _3715_ (.B1(_1018_),
    .Y(_1019_),
    .A1(_1209_),
    .A2(net186));
 sg13g2_nand2b_1 _3716_ (.Y(_1020_),
    .B(_1019_),
    .A_N(_1017_));
 sg13g2_nand2b_1 _3717_ (.Y(_1021_),
    .B(_1017_),
    .A_N(_1019_));
 sg13g2_nand3_1 _3718_ (.B(_1020_),
    .C(_1021_),
    .A(net190),
    .Y(_1022_));
 sg13g2_o21ai_1 _3719_ (.B1(_1022_),
    .Y(_0097_),
    .A1(_1208_),
    .A2(net208));
 sg13g2_o21ai_1 _3720_ (.B1(_1020_),
    .Y(_1023_),
    .A1(_1208_),
    .A2(_0758_));
 sg13g2_or2_1 _3721_ (.X(_1024_),
    .B(net188),
    .A(net506));
 sg13g2_xnor2_1 _3722_ (.Y(_1025_),
    .A(net380),
    .B(net188));
 sg13g2_xnor2_1 _3723_ (.Y(_1026_),
    .A(_1023_),
    .B(_1025_));
 sg13g2_a22oi_1 _3724_ (.Y(_1027_),
    .B1(net190),
    .B2(_1026_),
    .A2(net201),
    .A1(net380));
 sg13g2_inv_1 _3725_ (.Y(_0098_),
    .A(_1027_));
 sg13g2_a21o_1 _3726_ (.A2(net188),
    .A1(net506),
    .B1(_1023_),
    .X(_1028_));
 sg13g2_and3_1 _3727_ (.X(_1029_),
    .A(net208),
    .B(_1024_),
    .C(_1028_));
 sg13g2_nor2_1 _3728_ (.A(net372),
    .B(_1029_),
    .Y(_1030_));
 sg13g2_and4_1 _3729_ (.A(net372),
    .B(net208),
    .C(_1024_),
    .D(_1028_),
    .X(_1031_));
 sg13g2_and2_1 _3730_ (.A(net372),
    .B(_1029_),
    .X(_1032_));
 sg13g2_nor3_1 _3731_ (.A(net194),
    .B(_1030_),
    .C(_1032_),
    .Y(_0099_));
 sg13g2_nor2_1 _3732_ (.A(net389),
    .B(_1031_),
    .Y(_1033_));
 sg13g2_and2_1 _3733_ (.A(net389),
    .B(_1032_),
    .X(_1034_));
 sg13g2_nor3_1 _3734_ (.A(net194),
    .B(_1033_),
    .C(_1034_),
    .Y(_0100_));
 sg13g2_nor2_1 _3735_ (.A(net415),
    .B(_1034_),
    .Y(_1035_));
 sg13g2_and2_1 _3736_ (.A(net415),
    .B(_1034_),
    .X(_1036_));
 sg13g2_nor3_1 _3737_ (.A(net194),
    .B(_1035_),
    .C(_1036_),
    .Y(_0101_));
 sg13g2_nor2_1 _3738_ (.A(net407),
    .B(_1036_),
    .Y(_1037_));
 sg13g2_and4_1 _3739_ (.A(net407),
    .B(\sin_y_acc[18] ),
    .C(net389),
    .D(_1031_),
    .X(_1038_));
 sg13g2_nor3_1 _3740_ (.A(net194),
    .B(net408),
    .C(_1038_),
    .Y(_0102_));
 sg13g2_nor2_1 _3741_ (.A(net383),
    .B(_1038_),
    .Y(_1039_));
 sg13g2_and3_1 _3742_ (.X(_1040_),
    .A(net383),
    .B(\sin_y_acc[19] ),
    .C(_1036_));
 sg13g2_nor3_1 _3743_ (.A(net194),
    .B(net384),
    .C(_1040_),
    .Y(_0103_));
 sg13g2_nor2_1 _3744_ (.A(net323),
    .B(_1040_),
    .Y(_1041_));
 sg13g2_and3_2 _3745_ (.X(_1042_),
    .A(net323),
    .B(\sin_y_acc[20] ),
    .C(_1038_));
 sg13g2_nor3_1 _3746_ (.A(net194),
    .B(net324),
    .C(_1042_),
    .Y(_0104_));
 sg13g2_nor2_1 _3747_ (.A(net345),
    .B(_1042_),
    .Y(_1043_));
 sg13g2_and2_1 _3748_ (.A(net345),
    .B(_1042_),
    .X(_1044_));
 sg13g2_nor3_1 _3749_ (.A(net197),
    .B(net346),
    .C(_1044_),
    .Y(_0105_));
 sg13g2_or2_1 _3750_ (.X(_1045_),
    .B(_1044_),
    .A(net445));
 sg13g2_a21oi_1 _3751_ (.A1(net445),
    .A2(_1044_),
    .Y(_1046_),
    .B1(net195));
 sg13g2_and2_1 _3752_ (.A(_1045_),
    .B(_1046_),
    .X(_0106_));
 sg13g2_a21oi_1 _3753_ (.A1(\sin_y_acc[23] ),
    .A2(_1044_),
    .Y(_1047_),
    .B1(net263));
 sg13g2_and3_2 _3754_ (.X(_1048_),
    .A(net263),
    .B(\sin_y_acc[23] ),
    .C(_1044_));
 sg13g2_nor3_1 _3755_ (.A(net196),
    .B(net264),
    .C(_1048_),
    .Y(_0107_));
 sg13g2_a21oi_1 _3756_ (.A1(net405),
    .A2(_1048_),
    .Y(_1049_),
    .B1(net195));
 sg13g2_o21ai_1 _3757_ (.B1(_1049_),
    .Y(_1050_),
    .A1(net405),
    .A2(_1048_));
 sg13g2_inv_1 _3758_ (.Y(_0108_),
    .A(net406));
 sg13g2_a21oi_1 _3759_ (.A1(\sin_y_acc[25] ),
    .A2(_1048_),
    .Y(_1051_),
    .B1(net170));
 sg13g2_and3_1 _3760_ (.X(_1052_),
    .A(net170),
    .B(\sin_y_acc[25] ),
    .C(_1048_));
 sg13g2_nor3_1 _3761_ (.A(net195),
    .B(net171),
    .C(_1052_),
    .Y(_0109_));
 sg13g2_xnor2_1 _3762_ (.Y(_1053_),
    .A(net398),
    .B(_0945_));
 sg13g2_nor2_1 _3763_ (.A(net197),
    .B(_1053_),
    .Y(_0110_));
 sg13g2_nand2_1 _3764_ (.Y(_1054_),
    .A(net398),
    .B(net187));
 sg13g2_nand2_1 _3765_ (.Y(_1055_),
    .A(\cos_y_acc[1] ),
    .B(_0574_));
 sg13g2_xor2_1 _3766_ (.B(_0574_),
    .A(net401),
    .X(_1056_));
 sg13g2_nand2b_1 _3767_ (.Y(_1057_),
    .B(_1056_),
    .A_N(_1054_));
 sg13g2_xnor2_1 _3768_ (.Y(_1058_),
    .A(_1054_),
    .B(_1056_));
 sg13g2_a22oi_1 _3769_ (.Y(_1059_),
    .B1(net192),
    .B2(_1058_),
    .A2(net204),
    .A1(net401));
 sg13g2_inv_1 _3770_ (.Y(_0111_),
    .A(_1059_));
 sg13g2_xor2_1 _3771_ (.B(_0594_),
    .A(net396),
    .X(_1060_));
 sg13g2_and2_1 _3772_ (.A(_1055_),
    .B(_1057_),
    .X(_1061_));
 sg13g2_nor2_1 _3773_ (.A(_1060_),
    .B(_1061_),
    .Y(_1062_));
 sg13g2_o21ai_1 _3774_ (.B1(net192),
    .Y(_1063_),
    .A1(_1060_),
    .A2(_1061_));
 sg13g2_a21oi_1 _3775_ (.A1(_1060_),
    .A2(_1061_),
    .Y(_1064_),
    .B1(_1063_));
 sg13g2_a21o_1 _3776_ (.A2(net203),
    .A1(net396),
    .B1(_1064_),
    .X(_0112_));
 sg13g2_nand2b_1 _3777_ (.Y(_1065_),
    .B(\cos_y_acc[3] ),
    .A_N(_0615_));
 sg13g2_xnor2_1 _3778_ (.Y(_1066_),
    .A(net399),
    .B(_0615_));
 sg13g2_a21oi_1 _3779_ (.A1(net396),
    .A2(_0595_),
    .Y(_1067_),
    .B1(_1062_));
 sg13g2_nand2b_1 _3780_ (.Y(_1068_),
    .B(_1066_),
    .A_N(_1067_));
 sg13g2_nand2b_1 _3781_ (.Y(_1069_),
    .B(_1067_),
    .A_N(_1066_));
 sg13g2_nand3_1 _3782_ (.B(_1068_),
    .C(_1069_),
    .A(net192),
    .Y(_1070_));
 sg13g2_o21ai_1 _3783_ (.B1(_1070_),
    .Y(_0113_),
    .A1(_1206_),
    .A2(net207));
 sg13g2_xnor2_1 _3784_ (.Y(_1071_),
    .A(net386),
    .B(_0633_));
 sg13g2_inv_1 _3785_ (.Y(_1072_),
    .A(_1071_));
 sg13g2_a21o_1 _3786_ (.A2(_1068_),
    .A1(_1065_),
    .B1(_1072_),
    .X(_1073_));
 sg13g2_nand3_1 _3787_ (.B(_1068_),
    .C(_1072_),
    .A(_1065_),
    .Y(_1074_));
 sg13g2_nand3_1 _3788_ (.B(_1073_),
    .C(_1074_),
    .A(net192),
    .Y(_1075_));
 sg13g2_o21ai_1 _3789_ (.B1(_1075_),
    .Y(_0114_),
    .A1(_1205_),
    .A2(net207));
 sg13g2_o21ai_1 _3790_ (.B1(_1073_),
    .Y(_1076_),
    .A1(_1205_),
    .A2(_0633_));
 sg13g2_nand2_1 _3791_ (.Y(_1077_),
    .A(_1204_),
    .B(_0650_));
 sg13g2_nor2_1 _3792_ (.A(_1204_),
    .B(_0650_),
    .Y(_1078_));
 sg13g2_xnor2_1 _3793_ (.Y(_1079_),
    .A(net410),
    .B(_0650_));
 sg13g2_o21ai_1 _3794_ (.B1(net191),
    .Y(_1080_),
    .A1(_1076_),
    .A2(_1079_));
 sg13g2_a21o_1 _3795_ (.A2(_1079_),
    .A1(_1076_),
    .B1(_1080_),
    .X(_1081_));
 sg13g2_o21ai_1 _3796_ (.B1(_1081_),
    .Y(_0115_),
    .A1(_1204_),
    .A2(net207));
 sg13g2_xnor2_1 _3797_ (.Y(_1082_),
    .A(net414),
    .B(_0664_));
 sg13g2_a21oi_1 _3798_ (.A1(_1076_),
    .A2(_1077_),
    .Y(_1083_),
    .B1(_1078_));
 sg13g2_nor2_1 _3799_ (.A(_1082_),
    .B(_1083_),
    .Y(_1084_));
 sg13g2_o21ai_1 _3800_ (.B1(net189),
    .Y(_1085_),
    .A1(_1082_),
    .A2(_1083_));
 sg13g2_a21oi_1 _3801_ (.A1(_1082_),
    .A2(_1083_),
    .Y(_1086_),
    .B1(_1085_));
 sg13g2_a21o_1 _3802_ (.A2(net198),
    .A1(net414),
    .B1(_1086_),
    .X(_0116_));
 sg13g2_xnor2_1 _3803_ (.Y(_1087_),
    .A(net434),
    .B(_0679_));
 sg13g2_a21o_1 _3804_ (.A2(_0664_),
    .A1(\cos_y_acc[6] ),
    .B1(_1084_),
    .X(_1088_));
 sg13g2_nand2_1 _3805_ (.Y(_1089_),
    .A(_1087_),
    .B(_1088_));
 sg13g2_o21ai_1 _3806_ (.B1(net189),
    .Y(_1090_),
    .A1(_1087_),
    .A2(_1088_));
 sg13g2_nand2b_1 _3807_ (.Y(_1091_),
    .B(_1089_),
    .A_N(_1090_));
 sg13g2_o21ai_1 _3808_ (.B1(_1091_),
    .Y(_0117_),
    .A1(_1203_),
    .A2(net205));
 sg13g2_nand2_1 _3809_ (.Y(_1092_),
    .A(\cos_y_acc[8] ),
    .B(_0693_));
 sg13g2_xnor2_1 _3810_ (.Y(_1093_),
    .A(net447),
    .B(_0693_));
 sg13g2_o21ai_1 _3811_ (.B1(_1089_),
    .Y(_1094_),
    .A1(_1203_),
    .A2(_0679_));
 sg13g2_nand2b_1 _3812_ (.Y(_1095_),
    .B(_1094_),
    .A_N(_1093_));
 sg13g2_nand2b_1 _3813_ (.Y(_1096_),
    .B(_1093_),
    .A_N(_1094_));
 sg13g2_nand3_1 _3814_ (.B(_1095_),
    .C(_1096_),
    .A(net189),
    .Y(_1097_));
 sg13g2_o21ai_1 _3815_ (.B1(_1097_),
    .Y(_0118_),
    .A1(_1202_),
    .A2(net205));
 sg13g2_nand2_1 _3816_ (.Y(_1098_),
    .A(_1092_),
    .B(_1095_));
 sg13g2_xnor2_1 _3817_ (.Y(_1099_),
    .A(_1201_),
    .B(_0705_));
 sg13g2_o21ai_1 _3818_ (.B1(net190),
    .Y(_1100_),
    .A1(_1098_),
    .A2(_1099_));
 sg13g2_a21o_1 _3819_ (.A2(_1099_),
    .A1(_1098_),
    .B1(_1100_),
    .X(_1101_));
 sg13g2_o21ai_1 _3820_ (.B1(_1101_),
    .Y(_0119_),
    .A1(_1201_),
    .A2(net206));
 sg13g2_xnor2_1 _3821_ (.Y(_1102_),
    .A(net432),
    .B(_0717_));
 sg13g2_a22oi_1 _3822_ (.Y(_1103_),
    .B1(_1092_),
    .B2(_1095_),
    .A2(_0706_),
    .A1(_1201_));
 sg13g2_a21oi_1 _3823_ (.A1(\cos_y_acc[9] ),
    .A2(_0705_),
    .Y(_1104_),
    .B1(_1103_));
 sg13g2_or2_1 _3824_ (.X(_1105_),
    .B(_1104_),
    .A(_1102_));
 sg13g2_nand2_1 _3825_ (.Y(_1106_),
    .A(_1102_),
    .B(_1104_));
 sg13g2_nand3_1 _3826_ (.B(_1105_),
    .C(_1106_),
    .A(net190),
    .Y(_1107_));
 sg13g2_o21ai_1 _3827_ (.B1(_1107_),
    .Y(_0120_),
    .A1(_1200_),
    .A2(net206));
 sg13g2_o21ai_1 _3828_ (.B1(_1105_),
    .Y(_1108_),
    .A1(_1200_),
    .A2(_0718_));
 sg13g2_xnor2_1 _3829_ (.Y(_1109_),
    .A(net425),
    .B(_0731_));
 sg13g2_o21ai_1 _3830_ (.B1(net191),
    .Y(_1110_),
    .A1(_1108_),
    .A2(_1109_));
 sg13g2_a21o_1 _3831_ (.A2(_1109_),
    .A1(_1108_),
    .B1(_1110_),
    .X(_1111_));
 sg13g2_o21ai_1 _3832_ (.B1(_1111_),
    .Y(_0121_),
    .A1(_1199_),
    .A2(net206));
 sg13g2_nand2_1 _3833_ (.Y(_1112_),
    .A(\cos_y_acc[12] ),
    .B(_0742_));
 sg13g2_xnor2_1 _3834_ (.Y(_1113_),
    .A(net426),
    .B(_0742_));
 sg13g2_o21ai_1 _3835_ (.B1(_1108_),
    .Y(_1114_),
    .A1(\cos_y_acc[11] ),
    .A2(_0732_));
 sg13g2_o21ai_1 _3836_ (.B1(_1114_),
    .Y(_1115_),
    .A1(_1199_),
    .A2(_0731_));
 sg13g2_nand2b_1 _3837_ (.Y(_1116_),
    .B(_1115_),
    .A_N(_1113_));
 sg13g2_nand2b_1 _3838_ (.Y(_1117_),
    .B(_1113_),
    .A_N(_1115_));
 sg13g2_nand3_1 _3839_ (.B(_1116_),
    .C(_1117_),
    .A(net193),
    .Y(_1118_));
 sg13g2_o21ai_1 _3840_ (.B1(_1118_),
    .Y(_0122_),
    .A1(_1198_),
    .A2(net208));
 sg13g2_nand2_1 _3841_ (.Y(_1119_),
    .A(net351),
    .B(net202));
 sg13g2_nand2_1 _3842_ (.Y(_1120_),
    .A(_1112_),
    .B(_1116_));
 sg13g2_nand2_1 _3843_ (.Y(_1121_),
    .A(net351),
    .B(_0753_));
 sg13g2_inv_1 _3844_ (.Y(_1122_),
    .A(_1121_));
 sg13g2_or2_1 _3845_ (.X(_1123_),
    .B(_0753_),
    .A(net351));
 sg13g2_nand3_1 _3846_ (.B(_1121_),
    .C(_1123_),
    .A(_1120_),
    .Y(_1124_));
 sg13g2_a21oi_1 _3847_ (.A1(_1121_),
    .A2(_1123_),
    .Y(_1125_),
    .B1(_1120_));
 sg13g2_nand2_1 _3848_ (.Y(_1126_),
    .A(net193),
    .B(_1124_));
 sg13g2_o21ai_1 _3849_ (.B1(_1119_),
    .Y(_0123_),
    .A1(_1125_),
    .A2(_1126_));
 sg13g2_nand2_1 _3850_ (.Y(_1127_),
    .A(net422),
    .B(_0758_));
 sg13g2_xnor2_1 _3851_ (.Y(_1128_),
    .A(_1197_),
    .B(_0758_));
 sg13g2_o21ai_1 _3852_ (.B1(_1123_),
    .Y(_1129_),
    .A1(_1120_),
    .A2(_1122_));
 sg13g2_nand2b_1 _3853_ (.Y(_1130_),
    .B(_1128_),
    .A_N(_1129_));
 sg13g2_nand2b_1 _3854_ (.Y(_1131_),
    .B(_1129_),
    .A_N(_1128_));
 sg13g2_nand3_1 _3855_ (.B(_1130_),
    .C(_1131_),
    .A(net193),
    .Y(_1132_));
 sg13g2_o21ai_1 _3856_ (.B1(_1132_),
    .Y(_0124_),
    .A1(_1197_),
    .A2(net208));
 sg13g2_nand2_1 _3857_ (.Y(_1133_),
    .A(_1127_),
    .B(_1130_));
 sg13g2_nor2b_1 _3858_ (.A(net188),
    .B_N(\cos_y_acc[15] ),
    .Y(_1134_));
 sg13g2_nand2b_1 _3859_ (.Y(_1135_),
    .B(_0766_),
    .A_N(\cos_y_acc[15] ));
 sg13g2_nor2b_1 _3860_ (.A(_1134_),
    .B_N(_1135_),
    .Y(_1136_));
 sg13g2_o21ai_1 _3861_ (.B1(net193),
    .Y(_1137_),
    .A1(_1133_),
    .A2(_1136_));
 sg13g2_a21oi_1 _3862_ (.A1(_1133_),
    .A2(_1136_),
    .Y(_1138_),
    .B1(_1137_));
 sg13g2_a21o_1 _3863_ (.A2(_0555_),
    .A1(net431),
    .B1(_1138_),
    .X(_0125_));
 sg13g2_or2_1 _3864_ (.X(_1139_),
    .B(_1134_),
    .A(_1133_));
 sg13g2_and3_1 _3865_ (.X(_1140_),
    .A(net209),
    .B(_1135_),
    .C(_1139_));
 sg13g2_nor2_1 _3866_ (.A(net420),
    .B(_1140_),
    .Y(_1141_));
 sg13g2_and4_1 _3867_ (.A(net420),
    .B(net209),
    .C(_1135_),
    .D(_1139_),
    .X(_1142_));
 sg13g2_nor3_1 _3868_ (.A(net194),
    .B(_1141_),
    .C(_1142_),
    .Y(_0126_));
 sg13g2_nor2_1 _3869_ (.A(net417),
    .B(_1142_),
    .Y(_1143_));
 sg13g2_and3_2 _3870_ (.X(_1144_),
    .A(net417),
    .B(net420),
    .C(_1140_));
 sg13g2_nor3_1 _3871_ (.A(net194),
    .B(net418),
    .C(_1144_),
    .Y(_0127_));
 sg13g2_xnor2_1 _3872_ (.Y(_1145_),
    .A(net439),
    .B(_1144_));
 sg13g2_nor2_1 _3873_ (.A(net196),
    .B(_1145_),
    .Y(_0128_));
 sg13g2_a21oi_1 _3874_ (.A1(\cos_y_acc[18] ),
    .A2(_1144_),
    .Y(_1146_),
    .B1(net336));
 sg13g2_and4_1 _3875_ (.A(net336),
    .B(net439),
    .C(net417),
    .D(_1142_),
    .X(_1147_));
 sg13g2_nor3_1 _3876_ (.A(net196),
    .B(net337),
    .C(_1147_),
    .Y(_0129_));
 sg13g2_nor2_1 _3877_ (.A(net248),
    .B(_1147_),
    .Y(_1148_));
 sg13g2_a21oi_1 _3878_ (.A1(net248),
    .A2(_1147_),
    .Y(_1149_),
    .B1(net196));
 sg13g2_nor2b_1 _3879_ (.A(_1148_),
    .B_N(_1149_),
    .Y(_0130_));
 sg13g2_a21oi_1 _3880_ (.A1(net248),
    .A2(_1147_),
    .Y(_1150_),
    .B1(net340));
 sg13g2_and3_2 _3881_ (.X(_1151_),
    .A(net340),
    .B(net463),
    .C(_1147_));
 sg13g2_nor3_1 _3882_ (.A(net196),
    .B(net341),
    .C(_1151_),
    .Y(_0131_));
 sg13g2_a21oi_1 _3883_ (.A1(net247),
    .A2(_1151_),
    .Y(_1152_),
    .B1(net195));
 sg13g2_o21ai_1 _3884_ (.B1(_1152_),
    .Y(_1153_),
    .A1(net247),
    .A2(_1151_));
 sg13g2_inv_1 _3885_ (.Y(_0132_),
    .A(_1153_));
 sg13g2_a21oi_1 _3886_ (.A1(net247),
    .A2(_1151_),
    .Y(_1154_),
    .B1(net361));
 sg13g2_and3_1 _3887_ (.X(_1155_),
    .A(net361),
    .B(net247),
    .C(_1151_));
 sg13g2_nor3_1 _3888_ (.A(net195),
    .B(net362),
    .C(_1155_),
    .Y(_0133_));
 sg13g2_nor2_1 _3889_ (.A(net353),
    .B(_1155_),
    .Y(_1156_));
 sg13g2_and4_1 _3890_ (.A(net353),
    .B(\cos_y_acc[23] ),
    .C(net503),
    .D(_1151_),
    .X(_1157_));
 sg13g2_nor3_1 _3891_ (.A(net195),
    .B(net354),
    .C(_1157_),
    .Y(_0134_));
 sg13g2_nor2_1 _3892_ (.A(net349),
    .B(_1157_),
    .Y(_1158_));
 sg13g2_and2_1 _3893_ (.A(net349),
    .B(_1157_),
    .X(_1159_));
 sg13g2_nor3_1 _3894_ (.A(net195),
    .B(net350),
    .C(_1159_),
    .Y(_0135_));
 sg13g2_a21oi_1 _3895_ (.A1(net395),
    .A2(_1159_),
    .Y(_1160_),
    .B1(net195));
 sg13g2_o21ai_1 _3896_ (.B1(_1160_),
    .Y(_1161_),
    .A1(net395),
    .A2(_1159_));
 sg13g2_inv_1 _3897_ (.Y(_0136_),
    .A(_1161_));
 sg13g2_nand4_1 _3898_ (.B(_0491_),
    .C(_0812_),
    .A(\hvsync_gen.vpos[9] ),
    .Y(_1162_),
    .D(_0813_));
 sg13g2_nand2_1 _3899_ (.Y(_1163_),
    .A(net253),
    .B(_1162_));
 sg13g2_or2_1 _3900_ (.X(_1164_),
    .B(_1163_),
    .A(_0797_));
 sg13g2_inv_1 _3901_ (.Y(_1165_),
    .A(net184));
 sg13g2_nor2_1 _3902_ (.A(_1215_),
    .B(_0798_),
    .Y(_1166_));
 sg13g2_a21oi_1 _3903_ (.A1(_1215_),
    .A2(net184),
    .Y(_0137_),
    .B1(_1166_));
 sg13g2_nand2_1 _3904_ (.Y(_1167_),
    .A(net246),
    .B(_0798_));
 sg13g2_xnor2_1 _3905_ (.Y(_1168_),
    .A(net343),
    .B(net246));
 sg13g2_o21ai_1 _3906_ (.B1(_1167_),
    .Y(_0138_),
    .A1(net184),
    .A2(_1168_));
 sg13g2_nand2_1 _3907_ (.Y(_1169_),
    .A(net309),
    .B(_0798_));
 sg13g2_a21oi_1 _3908_ (.A1(\bayer_j[0] ),
    .A2(net246),
    .Y(_1170_),
    .B1(net309));
 sg13g2_nand3_1 _3909_ (.B(net246),
    .C(net309),
    .A(\bayer_j[0] ),
    .Y(_1171_));
 sg13g2_nand2b_1 _3910_ (.Y(_1172_),
    .B(_1171_),
    .A_N(_1170_));
 sg13g2_o21ai_1 _3911_ (.B1(_1169_),
    .Y(_0139_),
    .A1(net184),
    .A2(_1172_));
 sg13g2_nand2_1 _3912_ (.Y(_1173_),
    .A(net332),
    .B(_0798_));
 sg13g2_nand3_1 _3913_ (.B(net246),
    .C(_0491_),
    .A(net343),
    .Y(_1174_));
 sg13g2_xor2_1 _3914_ (.B(_1171_),
    .A(net332),
    .X(_1175_));
 sg13g2_o21ai_1 _3915_ (.B1(_1173_),
    .Y(_0140_),
    .A1(net184),
    .A2(_1175_));
 sg13g2_nand2_1 _3916_ (.Y(_1176_),
    .A(net271),
    .B(_0798_));
 sg13g2_nand4_1 _3917_ (.B(net246),
    .C(net271),
    .A(net505),
    .Y(_1177_),
    .D(_0491_));
 sg13g2_xor2_1 _3918_ (.B(net344),
    .A(net271),
    .X(_1178_));
 sg13g2_o21ai_1 _3919_ (.B1(_1176_),
    .Y(_0141_),
    .A1(net184),
    .A2(_1178_));
 sg13g2_nand2_1 _3920_ (.Y(_1179_),
    .A(net297),
    .B(_0798_));
 sg13g2_xnor2_1 _3921_ (.Y(_1180_),
    .A(_1238_),
    .B(_1177_));
 sg13g2_o21ai_1 _3922_ (.B1(_1179_),
    .Y(_0142_),
    .A1(net184),
    .A2(_1180_));
 sg13g2_nand2_1 _3923_ (.Y(_1181_),
    .A(net322),
    .B(_0798_));
 sg13g2_o21ai_1 _3924_ (.B1(_1239_),
    .Y(_1182_),
    .A1(_1238_),
    .A2(_1177_));
 sg13g2_nor2_1 _3925_ (.A(_0273_),
    .B(_1177_),
    .Y(_1183_));
 sg13g2_o21ai_1 _3926_ (.B1(_1182_),
    .Y(_1184_),
    .A1(_0273_),
    .A2(_1177_));
 sg13g2_o21ai_1 _3927_ (.B1(_1181_),
    .Y(_0143_),
    .A1(net184),
    .A2(_1184_));
 sg13g2_nand2_1 _3928_ (.Y(_1185_),
    .A(net285),
    .B(_0798_));
 sg13g2_nor3_1 _3929_ (.A(_1240_),
    .B(_0273_),
    .C(_1177_),
    .Y(_1186_));
 sg13g2_xnor2_1 _3930_ (.Y(_1187_),
    .A(net285),
    .B(_1183_));
 sg13g2_o21ai_1 _3931_ (.B1(_1185_),
    .Y(_0144_),
    .A1(_1164_),
    .A2(_1187_));
 sg13g2_nand2_1 _3932_ (.Y(_1188_),
    .A(net305),
    .B(_1186_));
 sg13g2_nand2_1 _3933_ (.Y(_1189_),
    .A(_1165_),
    .B(_1188_));
 sg13g2_nand2_1 _3934_ (.Y(_1190_),
    .A(net185),
    .B(_1189_));
 sg13g2_a21oi_1 _3935_ (.A1(_1165_),
    .A2(_1186_),
    .Y(_1191_),
    .B1(net305));
 sg13g2_a21oi_1 _3936_ (.A1(_0799_),
    .A2(_1189_),
    .Y(_0145_),
    .B1(net306));
 sg13g2_nor3_1 _3937_ (.A(net424),
    .B(_1164_),
    .C(_1188_),
    .Y(_1192_));
 sg13g2_a21o_1 _3938_ (.A2(_1190_),
    .A1(net424),
    .B1(_1192_),
    .X(_0146_));
 sg13g2_dfrbpq_2 _3939_ (.RESET_B(net153),
    .D(_0002_),
    .Q(\cos_x_acc[0] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _3940_ (.RESET_B(net47),
    .D(net319),
    .Q(\cos_x_acc[1] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _3941_ (.RESET_B(net46),
    .D(net491),
    .Q(\cos_x_acc[2] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _3942_ (.RESET_B(net45),
    .D(_0005_),
    .Q(\cos_x_acc[3] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _3943_ (.RESET_B(net44),
    .D(net485),
    .Q(\cos_x_acc[4] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_2 _3944_ (.RESET_B(net43),
    .D(net458),
    .Q(\cos_x_acc[5] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 _3945_ (.RESET_B(net42),
    .D(_0008_),
    .Q(\cos_x_acc[6] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 _3946_ (.RESET_B(net41),
    .D(_0009_),
    .Q(\cos_x_acc[7] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 _3947_ (.RESET_B(net40),
    .D(_0010_),
    .Q(\cos_x_acc[8] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _3948_ (.RESET_B(net39),
    .D(net471),
    .Q(\cos_x_acc[9] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_2 _3949_ (.RESET_B(net38),
    .D(net449),
    .Q(\cos_x_acc[10] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _3950_ (.RESET_B(net37),
    .D(_0013_),
    .Q(\cos_x_acc[11] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_2 _3951_ (.RESET_B(net36),
    .D(net451),
    .Q(\cos_x_acc[12] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_2 _3952_ (.RESET_B(net35),
    .D(_0015_),
    .Q(\cos_x_acc[13] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_2 _3953_ (.RESET_B(net34),
    .D(net456),
    .Q(\cos_x_acc[14] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _3954_ (.RESET_B(net33),
    .D(_0017_),
    .Q(\cos_x_acc[15] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_2 _3955_ (.RESET_B(net32),
    .D(_0018_),
    .Q(\cos_x_acc[16] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _3956_ (.RESET_B(net31),
    .D(net376),
    .Q(\cos_x_acc[17] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _3957_ (.RESET_B(net30),
    .D(_0020_),
    .Q(\cos_x_acc[18] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_2 _3958_ (.RESET_B(net29),
    .D(net413),
    .Q(\cos_x_acc[19] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_2 _3959_ (.RESET_B(net28),
    .D(_0022_),
    .Q(\cos_x_acc[20] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _3960_ (.RESET_B(net27),
    .D(net260),
    .Q(\cos_x_acc[21] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _3961_ (.RESET_B(net26),
    .D(_0024_),
    .Q(\cos_x_acc[22] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 _3962_ (.RESET_B(net25),
    .D(net169),
    .Q(\cos_x_acc[23] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _3963_ (.RESET_B(net24),
    .D(net270),
    .Q(\cos_x_acc[24] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _3964_ (.RESET_B(net23),
    .D(_0027_),
    .Q(\cos_x_acc[25] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _3965_ (.RESET_B(net22),
    .D(_0028_),
    .Q(\cos_x_acc[26] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_2 _3966_ (.RESET_B(net21),
    .D(_0029_),
    .Q(\hvsync_gen.hpos[0] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _3967_ (.RESET_B(net20),
    .D(_0030_),
    .Q(\hvsync_gen.hpos[1] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _3968_ (.RESET_B(net19),
    .D(net379),
    .Q(\hvsync_gen.hpos[2] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _3969_ (.RESET_B(net18),
    .D(_0032_),
    .Q(\hvsync_gen.hpos[3] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _3970_ (.RESET_B(net163),
    .D(_0033_),
    .Q(\hvsync_gen.hpos[4] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 _3971_ (.RESET_B(net162),
    .D(net304),
    .Q(\hvsync_gen.hpos[5] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _3972_ (.RESET_B(net161),
    .D(net331),
    .Q(\hvsync_gen.hpos[6] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 _3973_ (.RESET_B(net160),
    .D(_0036_),
    .Q(\hvsync_gen.hpos[7] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 _3974_ (.RESET_B(net159),
    .D(net275),
    .Q(\hvsync_gen.hpos[8] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 _3975_ (.RESET_B(net158),
    .D(_0038_),
    .Q(\hvsync_gen.hpos[9] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _3976_ (.RESET_B(net157),
    .D(net468),
    .Q(\cos_addr[0] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 _3977_ (.RESET_B(net155),
    .D(net312),
    .Q(\cos_addr[1] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 _3978_ (.RESET_B(net152),
    .D(net284),
    .Q(\cos_addr[2] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _3979_ (.RESET_B(net150),
    .D(_0042_),
    .Q(\cos_addr[3] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 _3980_ (.RESET_B(net148),
    .D(net404),
    .Q(\cos_addr[4] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 _3981_ (.RESET_B(net146),
    .D(_0044_),
    .Q(\cos_addr[5] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 _3982_ (.RESET_B(net144),
    .D(net167),
    .Q(\cos_addr[6] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _3983_ (.RESET_B(net142),
    .D(net267),
    .Q(\y_prv[0] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _3984_ (.RESET_B(net141),
    .D(net314),
    .Q(\y_prv[1] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _3985_ (.RESET_B(net140),
    .D(_0048_),
    .Q(\y_prv[2] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _3986_ (.RESET_B(net139),
    .D(net321),
    .Q(\y_prv[3] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _3987_ (.RESET_B(net138),
    .D(_0050_),
    .Q(\y_prv[4] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _3988_ (.RESET_B(net137),
    .D(net257),
    .Q(\y_prv[5] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _3989_ (.RESET_B(net136),
    .D(net277),
    .Q(\y_prv[6] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _3990_ (.RESET_B(net135),
    .D(net262),
    .Q(\y_prv[7] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _3991_ (.RESET_B(net134),
    .D(_0054_),
    .Q(\y_prv[8] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _3992_ (.RESET_B(net133),
    .D(net317),
    .Q(\y_prv[9] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_2 _3993_ (.RESET_B(net132),
    .D(_0056_),
    .Q(\sin_x_acc[0] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _3994_ (.RESET_B(net131),
    .D(net371),
    .Q(\sin_x_acc[1] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _3995_ (.RESET_B(net130),
    .D(net480),
    .Q(\sin_x_acc[2] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _3996_ (.RESET_B(net129),
    .D(net477),
    .Q(\sin_x_acc[3] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 _3997_ (.RESET_B(net128),
    .D(_0060_),
    .Q(\sin_x_acc[4] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_2 _3998_ (.RESET_B(net127),
    .D(net461),
    .Q(\sin_x_acc[5] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 _3999_ (.RESET_B(net126),
    .D(_0062_),
    .Q(\sin_x_acc[6] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 _4000_ (.RESET_B(net125),
    .D(_0063_),
    .Q(\sin_x_acc[7] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_2 _4001_ (.RESET_B(net124),
    .D(_0064_),
    .Q(\sin_x_acc[8] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_2 _4002_ (.RESET_B(net123),
    .D(net473),
    .Q(\sin_x_acc[9] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_2 _4003_ (.RESET_B(net122),
    .D(_0066_),
    .Q(\sin_x_acc[10] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_2 _4004_ (.RESET_B(net121),
    .D(net494),
    .Q(\sin_x_acc[11] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_2 _4005_ (.RESET_B(net120),
    .D(net475),
    .Q(\sin_x_acc[12] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 _4006_ (.RESET_B(net119),
    .D(_0069_),
    .Q(\sin_x_acc[13] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_2 _4007_ (.RESET_B(net118),
    .D(net482),
    .Q(\sin_x_acc[14] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 _4008_ (.RESET_B(net117),
    .D(_0071_),
    .Q(\sin_x_acc[15] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 _4009_ (.RESET_B(net116),
    .D(_0072_),
    .Q(\sin_x_acc[16] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _4010_ (.RESET_B(net115),
    .D(net335),
    .Q(\sin_x_acc[17] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 _4011_ (.RESET_B(net114),
    .D(_0074_),
    .Q(\sin_x_acc[18] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 _4012_ (.RESET_B(net113),
    .D(net438),
    .Q(\sin_x_acc[19] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _4013_ (.RESET_B(net112),
    .D(_0076_),
    .Q(\sin_x_acc[20] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _4014_ (.RESET_B(net111),
    .D(net328),
    .Q(\sin_x_acc[21] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _4015_ (.RESET_B(net110),
    .D(_0078_),
    .Q(\sin_x_acc[22] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _4016_ (.RESET_B(net109),
    .D(net301),
    .Q(\sin_x_acc[23] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 _4017_ (.RESET_B(net108),
    .D(_0080_),
    .Q(\sin_x_acc[24] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 _4018_ (.RESET_B(net107),
    .D(_0081_),
    .Q(\sin_x_acc[25] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _4019_ (.RESET_B(net106),
    .D(net290),
    .Q(\sin_x_acc[26] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_2 _4020_ (.RESET_B(net105),
    .D(_0083_),
    .Q(\sin_y_acc[0] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 _4021_ (.RESET_B(net103),
    .D(net359),
    .Q(\sin_y_acc[1] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _4022_ (.RESET_B(net101),
    .D(_0085_),
    .Q(\sin_y_acc[2] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _4023_ (.RESET_B(net99),
    .D(net279),
    .Q(\sin_y_acc[3] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 _4024_ (.RESET_B(net97),
    .D(_0087_),
    .Q(\sin_y_acc[4] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 _4025_ (.RESET_B(net95),
    .D(_0088_),
    .Q(\sin_y_acc[5] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 _4026_ (.RESET_B(net93),
    .D(net296),
    .Q(\sin_y_acc[6] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_2 _4027_ (.RESET_B(net91),
    .D(_0090_),
    .Q(\sin_y_acc[7] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 _4028_ (.RESET_B(net89),
    .D(net367),
    .Q(\sin_y_acc[8] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 _4029_ (.RESET_B(net87),
    .D(net382),
    .Q(\sin_y_acc[9] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_2 _4030_ (.RESET_B(net85),
    .D(net281),
    .Q(\sin_y_acc[10] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_2 _4031_ (.RESET_B(net83),
    .D(_0094_),
    .Q(\sin_y_acc[11] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_2 _4032_ (.RESET_B(net81),
    .D(net374),
    .Q(\sin_y_acc[12] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_2 _4033_ (.RESET_B(net79),
    .D(_0096_),
    .Q(\sin_y_acc[13] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_2 _4034_ (.RESET_B(net77),
    .D(_0097_),
    .Q(\sin_y_acc[14] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_2 _4035_ (.RESET_B(net75),
    .D(_0098_),
    .Q(\sin_y_acc[15] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_2 _4036_ (.RESET_B(net73),
    .D(_0099_),
    .Q(\sin_y_acc[16] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _4037_ (.RESET_B(net71),
    .D(_0100_),
    .Q(\sin_y_acc[17] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _4038_ (.RESET_B(net69),
    .D(_0101_),
    .Q(\sin_y_acc[18] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _4039_ (.RESET_B(net67),
    .D(net409),
    .Q(\sin_y_acc[19] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _4040_ (.RESET_B(net65),
    .D(net385),
    .Q(\sin_y_acc[20] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_2 _4041_ (.RESET_B(net63),
    .D(net325),
    .Q(\sin_y_acc[21] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_2 _4042_ (.RESET_B(net61),
    .D(_0105_),
    .Q(\sin_y_acc[22] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _4043_ (.RESET_B(net59),
    .D(_0106_),
    .Q(\sin_y_acc[23] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _4044_ (.RESET_B(net57),
    .D(net265),
    .Q(\sin_y_acc[24] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _4045_ (.RESET_B(net55),
    .D(_0108_),
    .Q(\sin_y_acc[25] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _4046_ (.RESET_B(net53),
    .D(net255),
    .Q(\sin_y_acc[26] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _4047_ (.RESET_B(net51),
    .D(_0110_),
    .Q(\cos_y_acc[0] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _4048_ (.RESET_B(net49),
    .D(_0111_),
    .Q(\cos_y_acc[1] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _4049_ (.RESET_B(net156),
    .D(net397),
    .Q(\cos_y_acc[2] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_2 _4050_ (.RESET_B(net151),
    .D(_0113_),
    .Q(\cos_y_acc[3] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_2 _4051_ (.RESET_B(net147),
    .D(net387),
    .Q(\cos_y_acc[4] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_2 _4052_ (.RESET_B(net143),
    .D(_0115_),
    .Q(\cos_y_acc[5] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_2 _4053_ (.RESET_B(net102),
    .D(_0116_),
    .Q(\cos_y_acc[6] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 _4054_ (.RESET_B(net98),
    .D(net435),
    .Q(\cos_y_acc[7] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_2 _4055_ (.RESET_B(net94),
    .D(_0118_),
    .Q(\cos_y_acc[8] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_2 _4056_ (.RESET_B(net90),
    .D(net444),
    .Q(\cos_y_acc[9] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_2 _4057_ (.RESET_B(net86),
    .D(net433),
    .Q(\cos_y_acc[10] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_2 _4058_ (.RESET_B(net82),
    .D(_0121_),
    .Q(\cos_y_acc[11] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_2 _4059_ (.RESET_B(net78),
    .D(net427),
    .Q(\cos_y_acc[12] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 _4060_ (.RESET_B(net74),
    .D(net352),
    .Q(\cos_y_acc[13] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 _4061_ (.RESET_B(net70),
    .D(_0124_),
    .Q(\cos_y_acc[14] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 _4062_ (.RESET_B(net66),
    .D(_0125_),
    .Q(\cos_y_acc[15] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 _4063_ (.RESET_B(net62),
    .D(_0126_),
    .Q(\cos_y_acc[16] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 _4064_ (.RESET_B(net58),
    .D(net419),
    .Q(\cos_y_acc[17] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _4065_ (.RESET_B(net54),
    .D(_0128_),
    .Q(\cos_y_acc[18] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 _4066_ (.RESET_B(net50),
    .D(net338),
    .Q(\cos_y_acc[19] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _4067_ (.RESET_B(net154),
    .D(_0130_),
    .Q(\cos_y_acc[20] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _4068_ (.RESET_B(net145),
    .D(net342),
    .Q(\cos_y_acc[21] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _4069_ (.RESET_B(net100),
    .D(_0132_),
    .Q(\cos_y_acc[22] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _4070_ (.RESET_B(net92),
    .D(net363),
    .Q(\cos_y_acc[23] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _4071_ (.RESET_B(net84),
    .D(net355),
    .Q(\cos_y_acc[24] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _4072_ (.RESET_B(net76),
    .D(_0135_),
    .Q(\cos_y_acc[25] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _4073_ (.RESET_B(net164),
    .D(_0136_),
    .Q(\cos_y_acc[26] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _4074_ (.RESET_B(net68),
    .D(net294),
    .Q(hsync),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 _4075_ (.RESET_B(net60),
    .D(_0137_),
    .Q(\bayer_j[0] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_2 _4076_ (.RESET_B(net52),
    .D(_0138_),
    .Q(\bayer_j[1] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_2 _4077_ (.RESET_B(net149),
    .D(net310),
    .Q(\hvsync_gen.vpos[2] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 _4078_ (.RESET_B(net96),
    .D(net333),
    .Q(\hvsync_gen.vpos[3] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _4079_ (.RESET_B(net80),
    .D(_0141_),
    .Q(\hvsync_gen.vpos[4] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _4080_ (.RESET_B(net64),
    .D(net298),
    .Q(\hvsync_gen.vpos[5] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 _4081_ (.RESET_B(net48),
    .D(_0143_),
    .Q(\hvsync_gen.vpos[6] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _4082_ (.RESET_B(net88),
    .D(net286),
    .Q(\hvsync_gen.vpos[7] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_2 _4083_ (.RESET_B(net56),
    .D(net307),
    .Q(\hvsync_gen.vpos[8] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 _4084_ (.RESET_B(net104),
    .D(_0146_),
    .Q(\hvsync_gen.vpos[9] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _4085_ (.RESET_B(net72),
    .D(net272),
    .Q(\hvsync_gen.vsync ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_tiehi _3968__19 (.L_HI(net19));
 sg13g2_tiehi _3967__20 (.L_HI(net20));
 sg13g2_tiehi _3966__21 (.L_HI(net21));
 sg13g2_tiehi _3965__22 (.L_HI(net22));
 sg13g2_tiehi _3964__23 (.L_HI(net23));
 sg13g2_tiehi _3963__24 (.L_HI(net24));
 sg13g2_tiehi _3962__25 (.L_HI(net25));
 sg13g2_tiehi _3961__26 (.L_HI(net26));
 sg13g2_tiehi _3960__27 (.L_HI(net27));
 sg13g2_tiehi _3959__28 (.L_HI(net28));
 sg13g2_tiehi _3958__29 (.L_HI(net29));
 sg13g2_tiehi _3957__30 (.L_HI(net30));
 sg13g2_tiehi _3956__31 (.L_HI(net31));
 sg13g2_tiehi _3955__32 (.L_HI(net32));
 sg13g2_tiehi _3954__33 (.L_HI(net33));
 sg13g2_tiehi _3953__34 (.L_HI(net34));
 sg13g2_tiehi _3952__35 (.L_HI(net35));
 sg13g2_tiehi _3951__36 (.L_HI(net36));
 sg13g2_tiehi _3950__37 (.L_HI(net37));
 sg13g2_tiehi _3949__38 (.L_HI(net38));
 sg13g2_tiehi _3948__39 (.L_HI(net39));
 sg13g2_tiehi _3947__40 (.L_HI(net40));
 sg13g2_tiehi _3946__41 (.L_HI(net41));
 sg13g2_tiehi _3945__42 (.L_HI(net42));
 sg13g2_tiehi _3944__43 (.L_HI(net43));
 sg13g2_tiehi _3943__44 (.L_HI(net44));
 sg13g2_tiehi _3942__45 (.L_HI(net45));
 sg13g2_tiehi _3941__46 (.L_HI(net46));
 sg13g2_tiehi _3940__47 (.L_HI(net47));
 sg13g2_tiehi _4081__48 (.L_HI(net48));
 sg13g2_tiehi _4048__49 (.L_HI(net49));
 sg13g2_tiehi _4066__50 (.L_HI(net50));
 sg13g2_tiehi _4047__51 (.L_HI(net51));
 sg13g2_tiehi _4076__52 (.L_HI(net52));
 sg13g2_tiehi _4046__53 (.L_HI(net53));
 sg13g2_tiehi _4065__54 (.L_HI(net54));
 sg13g2_tiehi _4045__55 (.L_HI(net55));
 sg13g2_tiehi _4083__56 (.L_HI(net56));
 sg13g2_tiehi _4044__57 (.L_HI(net57));
 sg13g2_tiehi _4064__58 (.L_HI(net58));
 sg13g2_tiehi _4043__59 (.L_HI(net59));
 sg13g2_tiehi _4075__60 (.L_HI(net60));
 sg13g2_tiehi _4042__61 (.L_HI(net61));
 sg13g2_tiehi _4063__62 (.L_HI(net62));
 sg13g2_tiehi _4041__63 (.L_HI(net63));
 sg13g2_tiehi _4080__64 (.L_HI(net64));
 sg13g2_tiehi _4040__65 (.L_HI(net65));
 sg13g2_tiehi _4062__66 (.L_HI(net66));
 sg13g2_tiehi _4039__67 (.L_HI(net67));
 sg13g2_tiehi _4074__68 (.L_HI(net68));
 sg13g2_tiehi _4038__69 (.L_HI(net69));
 sg13g2_tiehi _4061__70 (.L_HI(net70));
 sg13g2_tiehi _4037__71 (.L_HI(net71));
 sg13g2_tiehi _4085__72 (.L_HI(net72));
 sg13g2_tiehi _4036__73 (.L_HI(net73));
 sg13g2_tiehi _4060__74 (.L_HI(net74));
 sg13g2_tiehi _4035__75 (.L_HI(net75));
 sg13g2_tiehi _4072__76 (.L_HI(net76));
 sg13g2_tiehi _4034__77 (.L_HI(net77));
 sg13g2_tiehi _4059__78 (.L_HI(net78));
 sg13g2_tiehi _4033__79 (.L_HI(net79));
 sg13g2_tiehi _4079__80 (.L_HI(net80));
 sg13g2_tiehi _4032__81 (.L_HI(net81));
 sg13g2_tiehi _4058__82 (.L_HI(net82));
 sg13g2_tiehi _4031__83 (.L_HI(net83));
 sg13g2_tiehi _4071__84 (.L_HI(net84));
 sg13g2_tiehi _4030__85 (.L_HI(net85));
 sg13g2_tiehi _4057__86 (.L_HI(net86));
 sg13g2_tiehi _4029__87 (.L_HI(net87));
 sg13g2_tiehi _4082__88 (.L_HI(net88));
 sg13g2_tiehi _4028__89 (.L_HI(net89));
 sg13g2_tiehi _4056__90 (.L_HI(net90));
 sg13g2_tiehi _4027__91 (.L_HI(net91));
 sg13g2_tiehi _4070__92 (.L_HI(net92));
 sg13g2_tiehi _4026__93 (.L_HI(net93));
 sg13g2_tiehi _4055__94 (.L_HI(net94));
 sg13g2_tiehi _4025__95 (.L_HI(net95));
 sg13g2_tiehi _4078__96 (.L_HI(net96));
 sg13g2_tiehi _4024__97 (.L_HI(net97));
 sg13g2_tiehi _4054__98 (.L_HI(net98));
 sg13g2_tiehi _4023__99 (.L_HI(net99));
 sg13g2_tiehi _4069__100 (.L_HI(net100));
 sg13g2_tiehi _4022__101 (.L_HI(net101));
 sg13g2_tiehi _4053__102 (.L_HI(net102));
 sg13g2_tiehi _4021__103 (.L_HI(net103));
 sg13g2_tiehi _4084__104 (.L_HI(net104));
 sg13g2_tiehi _4020__105 (.L_HI(net105));
 sg13g2_tiehi _4019__106 (.L_HI(net106));
 sg13g2_tiehi _4018__107 (.L_HI(net107));
 sg13g2_tiehi _4017__108 (.L_HI(net108));
 sg13g2_tiehi _4016__109 (.L_HI(net109));
 sg13g2_tiehi _4015__110 (.L_HI(net110));
 sg13g2_tiehi _4014__111 (.L_HI(net111));
 sg13g2_tiehi _4013__112 (.L_HI(net112));
 sg13g2_tiehi _4012__113 (.L_HI(net113));
 sg13g2_tiehi _4011__114 (.L_HI(net114));
 sg13g2_tiehi _4010__115 (.L_HI(net115));
 sg13g2_tiehi _4009__116 (.L_HI(net116));
 sg13g2_tiehi _4008__117 (.L_HI(net117));
 sg13g2_tiehi _4007__118 (.L_HI(net118));
 sg13g2_tiehi _4006__119 (.L_HI(net119));
 sg13g2_tiehi _4005__120 (.L_HI(net120));
 sg13g2_tiehi _4004__121 (.L_HI(net121));
 sg13g2_tiehi _4003__122 (.L_HI(net122));
 sg13g2_tiehi _4002__123 (.L_HI(net123));
 sg13g2_tiehi _4001__124 (.L_HI(net124));
 sg13g2_tiehi _4000__125 (.L_HI(net125));
 sg13g2_tiehi _3999__126 (.L_HI(net126));
 sg13g2_tiehi _3998__127 (.L_HI(net127));
 sg13g2_tiehi _3997__128 (.L_HI(net128));
 sg13g2_tiehi _3996__129 (.L_HI(net129));
 sg13g2_tiehi _3995__130 (.L_HI(net130));
 sg13g2_tiehi _3994__131 (.L_HI(net131));
 sg13g2_tiehi _3993__132 (.L_HI(net132));
 sg13g2_tiehi _3992__133 (.L_HI(net133));
 sg13g2_tiehi _3991__134 (.L_HI(net134));
 sg13g2_tiehi _3990__135 (.L_HI(net135));
 sg13g2_tiehi _3989__136 (.L_HI(net136));
 sg13g2_tiehi _3988__137 (.L_HI(net137));
 sg13g2_tiehi _3987__138 (.L_HI(net138));
 sg13g2_tiehi _3986__139 (.L_HI(net139));
 sg13g2_tiehi _3985__140 (.L_HI(net140));
 sg13g2_tiehi _3984__141 (.L_HI(net141));
 sg13g2_tiehi _3983__142 (.L_HI(net142));
 sg13g2_tiehi _4052__143 (.L_HI(net143));
 sg13g2_tiehi _3982__144 (.L_HI(net144));
 sg13g2_tiehi _4068__145 (.L_HI(net145));
 sg13g2_tiehi _3981__146 (.L_HI(net146));
 sg13g2_tiehi _4051__147 (.L_HI(net147));
 sg13g2_tiehi _3980__148 (.L_HI(net148));
 sg13g2_tiehi _4077__149 (.L_HI(net149));
 sg13g2_tiehi _3979__150 (.L_HI(net150));
 sg13g2_tiehi _4050__151 (.L_HI(net151));
 sg13g2_tiehi _3978__152 (.L_HI(net152));
 sg13g2_tiehi _3939__153 (.L_HI(net153));
 sg13g2_tiehi _4067__154 (.L_HI(net154));
 sg13g2_tiehi _3977__155 (.L_HI(net155));
 sg13g2_tiehi _4049__156 (.L_HI(net156));
 sg13g2_tiehi _3976__157 (.L_HI(net157));
 sg13g2_tiehi _3975__158 (.L_HI(net158));
 sg13g2_tiehi _3974__159 (.L_HI(net159));
 sg13g2_tiehi _3973__160 (.L_HI(net160));
 sg13g2_tiehi _3972__161 (.L_HI(net161));
 sg13g2_tiehi _3971__162 (.L_HI(net162));
 sg13g2_tiehi _3970__163 (.L_HI(net163));
 sg13g2_tiehi _4073__164 (.L_HI(net164));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_rejunity_vga_logo_3 (.L_LO(net3));
 sg13g2_tielo tt_um_rejunity_vga_logo_4 (.L_LO(net4));
 sg13g2_tielo tt_um_rejunity_vga_logo_5 (.L_LO(net5));
 sg13g2_tielo tt_um_rejunity_vga_logo_6 (.L_LO(net6));
 sg13g2_tielo tt_um_rejunity_vga_logo_7 (.L_LO(net7));
 sg13g2_tielo tt_um_rejunity_vga_logo_8 (.L_LO(net8));
 sg13g2_tielo tt_um_rejunity_vga_logo_9 (.L_LO(net9));
 sg13g2_tielo tt_um_rejunity_vga_logo_10 (.L_LO(net10));
 sg13g2_tielo tt_um_rejunity_vga_logo_11 (.L_LO(net11));
 sg13g2_tielo tt_um_rejunity_vga_logo_12 (.L_LO(net12));
 sg13g2_tielo tt_um_rejunity_vga_logo_13 (.L_LO(net13));
 sg13g2_tielo tt_um_rejunity_vga_logo_14 (.L_LO(net14));
 sg13g2_tielo tt_um_rejunity_vga_logo_15 (.L_LO(net15));
 sg13g2_tielo tt_um_rejunity_vga_logo_16 (.L_LO(net16));
 sg13g2_tielo tt_um_rejunity_vga_logo_17 (.L_LO(net17));
 sg13g2_tiehi _3969__18 (.L_HI(net18));
 sg13g2_buf_1 _4249_ (.A(\hvsync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _4250_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout172 (.A(_1776_),
    .X(net172));
 sg13g2_buf_8 fanout173 (.A(_1775_),
    .X(net173));
 sg13g2_buf_8 fanout174 (.A(_1804_),
    .X(net174));
 sg13g2_buf_8 fanout175 (.A(_1803_),
    .X(net175));
 sg13g2_buf_8 fanout176 (.A(_1816_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_1816_),
    .X(net177));
 sg13g2_buf_8 fanout178 (.A(_1815_),
    .X(net178));
 sg13g2_buf_8 fanout179 (.A(_1589_),
    .X(net179));
 sg13g2_buf_8 fanout180 (.A(_1592_),
    .X(net180));
 sg13g2_buf_8 fanout181 (.A(_1529_),
    .X(net181));
 sg13g2_buf_8 fanout182 (.A(_1585_),
    .X(net182));
 sg13g2_buf_8 fanout183 (.A(_0731_),
    .X(net183));
 sg13g2_buf_8 fanout184 (.A(_1164_),
    .X(net184));
 sg13g2_buf_8 fanout185 (.A(_0799_),
    .X(net185));
 sg13g2_buf_8 fanout186 (.A(_0753_),
    .X(net186));
 sg13g2_buf_8 fanout187 (.A(_0550_),
    .X(net187));
 sg13g2_buf_8 fanout188 (.A(_0766_),
    .X(net188));
 sg13g2_buf_8 fanout189 (.A(net191),
    .X(net189));
 sg13g2_buf_8 fanout190 (.A(net191),
    .X(net190));
 sg13g2_buf_8 fanout191 (.A(_0950_),
    .X(net191));
 sg13g2_buf_8 fanout192 (.A(_0950_),
    .X(net192));
 sg13g2_buf_1 fanout193 (.A(_0950_),
    .X(net193));
 sg13g2_buf_8 fanout194 (.A(net197),
    .X(net194));
 sg13g2_buf_8 fanout195 (.A(net196),
    .X(net195));
 sg13g2_buf_8 fanout196 (.A(net197),
    .X(net196));
 sg13g2_buf_8 fanout197 (.A(_0944_),
    .X(net197));
 sg13g2_buf_8 fanout198 (.A(net199),
    .X(net198));
 sg13g2_buf_8 fanout199 (.A(net202),
    .X(net199));
 sg13g2_buf_8 fanout200 (.A(net201),
    .X(net200));
 sg13g2_buf_8 fanout201 (.A(net202),
    .X(net201));
 sg13g2_buf_8 fanout202 (.A(_0555_),
    .X(net202));
 sg13g2_buf_8 fanout203 (.A(net204),
    .X(net203));
 sg13g2_buf_8 fanout204 (.A(_0555_),
    .X(net204));
 sg13g2_buf_8 fanout205 (.A(net207),
    .X(net205));
 sg13g2_buf_1 fanout206 (.A(net207),
    .X(net206));
 sg13g2_buf_8 fanout207 (.A(net212),
    .X(net207));
 sg13g2_buf_8 fanout208 (.A(net212),
    .X(net208));
 sg13g2_buf_1 fanout209 (.A(net212),
    .X(net209));
 sg13g2_buf_8 fanout210 (.A(net211),
    .X(net210));
 sg13g2_buf_8 fanout211 (.A(net212),
    .X(net211));
 sg13g2_buf_8 fanout212 (.A(_0554_),
    .X(net212));
 sg13g2_buf_8 fanout213 (.A(_0544_),
    .X(net213));
 sg13g2_buf_8 fanout214 (.A(net215),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_0528_),
    .X(net215));
 sg13g2_buf_8 fanout216 (.A(_0518_),
    .X(net216));
 sg13g2_buf_8 fanout217 (.A(_0536_),
    .X(net217));
 sg13g2_buf_8 fanout218 (.A(net219),
    .X(net218));
 sg13g2_buf_8 fanout219 (.A(_0526_),
    .X(net219));
 sg13g2_buf_8 fanout220 (.A(_0525_),
    .X(net220));
 sg13g2_buf_8 fanout221 (.A(_0525_),
    .X(net221));
 sg13g2_buf_8 fanout222 (.A(net224),
    .X(net222));
 sg13g2_buf_8 fanout223 (.A(net224),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(net225),
    .X(net224));
 sg13g2_buf_8 fanout225 (.A(_0510_),
    .X(net225));
 sg13g2_buf_8 fanout226 (.A(net227),
    .X(net226));
 sg13g2_buf_8 fanout227 (.A(net228),
    .X(net227));
 sg13g2_buf_8 fanout228 (.A(_0509_),
    .X(net228));
 sg13g2_buf_8 fanout229 (.A(net231),
    .X(net229));
 sg13g2_buf_8 fanout230 (.A(net231),
    .X(net230));
 sg13g2_buf_8 fanout231 (.A(_0508_),
    .X(net231));
 sg13g2_buf_8 fanout232 (.A(net233),
    .X(net232));
 sg13g2_buf_8 fanout233 (.A(net234),
    .X(net233));
 sg13g2_buf_8 fanout234 (.A(_0507_),
    .X(net234));
 sg13g2_buf_8 fanout235 (.A(_0501_),
    .X(net235));
 sg13g2_buf_1 fanout236 (.A(_0501_),
    .X(net236));
 sg13g2_buf_8 fanout237 (.A(net238),
    .X(net237));
 sg13g2_buf_8 fanout238 (.A(_0500_),
    .X(net238));
 sg13g2_buf_8 fanout239 (.A(net240),
    .X(net239));
 sg13g2_buf_8 fanout240 (.A(_0499_),
    .X(net240));
 sg13g2_buf_8 fanout241 (.A(_0498_),
    .X(net241));
 sg13g2_buf_8 fanout242 (.A(_0497_),
    .X(net242));
 sg13g2_buf_8 fanout243 (.A(net244),
    .X(net243));
 sg13g2_buf_8 fanout244 (.A(_0496_),
    .X(net244));
 sg13g2_buf_8 fanout245 (.A(_0178_),
    .X(net245));
 sg13g2_buf_8 fanout246 (.A(net459),
    .X(net246));
 sg13g2_buf_8 fanout247 (.A(net487),
    .X(net247));
 sg13g2_buf_8 fanout248 (.A(net463),
    .X(net248));
 sg13g2_buf_8 fanout249 (.A(net250),
    .X(net249));
 sg13g2_buf_8 fanout250 (.A(\cos_addr[6] ),
    .X(net250));
 sg13g2_buf_8 fanout251 (.A(net467),
    .X(net251));
 sg13g2_buf_8 fanout252 (.A(net253),
    .X(net252));
 sg13g2_buf_8 fanout253 (.A(net1),
    .X(net253));
 sg13g2_buf_8 fanout254 (.A(net1),
    .X(net254));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_tielo tt_um_rejunity_vga_logo_2 (.L_LO(net2));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_8 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_8 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_8 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_8 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_8 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_8 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_8 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_8 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_8 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_8 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_8 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_8 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_8 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_8 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_8 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_8 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_8 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_8 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_8 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_8 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_8 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_8 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_8 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_8 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_8 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_8 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_8 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_8 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_8 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_8 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_8 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\hvsync_gen.hpos[0] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold2 (.A(\cos_addr[6] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0045_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold4 (.A(\cos_x_acc[23] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0025_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold6 (.A(\sin_y_acc[26] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold7 (.A(_1051_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0109_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold9 (.A(\y_prv[5] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0051_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold11 (.A(\cos_x_acc[21] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0781_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0023_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold14 (.A(\y_prv[7] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0053_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold16 (.A(\sin_y_acc[24] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold17 (.A(_1047_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0107_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold19 (.A(\y_prv[0] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0046_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold21 (.A(\cos_x_acc[24] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0786_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0026_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold24 (.A(\hvsync_gen.vpos[4] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0001_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold26 (.A(\hvsync_gen.hpos[8] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0808_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0037_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold29 (.A(\y_prv[6] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0052_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold31 (.A(\sin_y_acc[3] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0086_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold33 (.A(\sin_y_acc[10] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0093_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold35 (.A(\cos_addr[2] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0834_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0041_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold38 (.A(\hvsync_gen.vpos[7] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0144_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold40 (.A(\sin_y_acc[4] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold41 (.A(\sin_x_acc[26] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0942_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0082_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold44 (.A(\y_prv[4] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold45 (.A(\hvsync_gen.hpos[9] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0494_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0000_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold48 (.A(\sin_y_acc[6] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0089_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold50 (.A(\hvsync_gen.vpos[5] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0142_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold52 (.A(\sin_x_acc[23] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0936_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0079_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold55 (.A(\hvsync_gen.hpos[5] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0804_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0034_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold58 (.A(\hvsync_gen.vpos[8] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold59 (.A(_1191_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0145_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold61 (.A(\y_prv[8] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold62 (.A(\hvsync_gen.vpos[2] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0139_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold64 (.A(\cos_addr[1] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0040_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold66 (.A(\y_prv[1] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0047_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold68 (.A(\y_prv[2] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold69 (.A(\y_prv[9] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0055_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold71 (.A(\cos_x_acc[0] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0003_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold73 (.A(\y_prv[3] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0049_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold75 (.A(\hvsync_gen.vpos[6] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold76 (.A(\sin_y_acc[21] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold77 (.A(_1041_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0104_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold79 (.A(\sin_x_acc[21] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0933_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0077_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold82 (.A(\hvsync_gen.hpos[6] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0805_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0035_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold85 (.A(\hvsync_gen.vpos[3] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0140_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold87 (.A(\sin_x_acc[17] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0073_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold89 (.A(\cos_y_acc[19] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold90 (.A(_1146_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0129_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold92 (.A(\sin_y_acc[14] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold93 (.A(\cos_y_acc[21] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold94 (.A(_1150_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0131_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold96 (.A(\bayer_j[0] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold97 (.A(_1174_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold98 (.A(\sin_y_acc[22] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold99 (.A(_1043_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold100 (.A(\hvsync_gen.hpos[3] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0801_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold102 (.A(\cos_y_acc[25] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold103 (.A(_1158_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold104 (.A(\cos_y_acc[13] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0123_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold106 (.A(\cos_y_acc[24] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold107 (.A(_1156_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0134_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold109 (.A(\sin_x_acc[24] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0938_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold111 (.A(\sin_y_acc[1] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0084_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold113 (.A(\sin_y_acc[5] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold114 (.A(\cos_y_acc[23] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold115 (.A(_1154_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0133_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold117 (.A(\cos_x_acc[20] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0780_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold119 (.A(\sin_y_acc[8] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0091_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold121 (.A(\sin_y_acc[11] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold122 (.A(\sin_y_acc[7] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold123 (.A(\sin_x_acc[0] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0057_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold125 (.A(\sin_y_acc[16] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold126 (.A(\sin_y_acc[12] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0095_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold128 (.A(\cos_x_acc[17] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0019_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold130 (.A(\hvsync_gen.hpos[2] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0800_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0031_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold133 (.A(\sin_y_acc[15] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold134 (.A(\sin_y_acc[9] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0092_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold136 (.A(\sin_y_acc[20] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold137 (.A(_1039_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0103_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold139 (.A(\cos_y_acc[4] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0114_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold141 (.A(\sin_y_acc[0] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold142 (.A(\sin_y_acc[17] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold143 (.A(\cos_x_acc[25] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0789_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold145 (.A(\hvsync_gen.hpos[7] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0807_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold147 (.A(\hvsync_gen.hpos[4] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold148 (.A(\cos_y_acc[26] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold149 (.A(\cos_y_acc[2] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0112_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold151 (.A(\cos_y_acc[0] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold152 (.A(\cos_y_acc[3] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold153 (.A(\cos_x_acc[26] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold154 (.A(\cos_y_acc[1] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold155 (.A(\cos_addr[4] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0839_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0043_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold158 (.A(\sin_y_acc[25] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold159 (.A(_1050_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold160 (.A(\sin_y_acc[19] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold161 (.A(_1037_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0102_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold163 (.A(\cos_y_acc[5] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold164 (.A(\cos_x_acc[19] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0779_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0021_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold167 (.A(\cos_y_acc[6] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold168 (.A(\sin_y_acc[18] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold169 (.A(\cos_addr[5] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold170 (.A(\cos_y_acc[17] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold171 (.A(_1143_),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0127_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold173 (.A(\cos_y_acc[16] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold174 (.A(\sin_x_acc[25] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold175 (.A(\cos_y_acc[14] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold176 (.A(\sin_y_acc[2] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold177 (.A(\hvsync_gen.vpos[9] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold178 (.A(\cos_y_acc[11] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold179 (.A(\cos_y_acc[12] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0122_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold181 (.A(\sin_x_acc[22] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0935_),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold183 (.A(\cos_x_acc[22] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold184 (.A(\cos_y_acc[15] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold185 (.A(\cos_y_acc[10] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0120_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold187 (.A(\cos_y_acc[7] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0117_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold189 (.A(\sin_x_acc[19] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0931_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0075_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold192 (.A(\cos_y_acc[18] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold193 (.A(\cos_addr[3] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold194 (.A(\sin_x_acc[20] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0932_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold196 (.A(\cos_y_acc[9] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0119_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold198 (.A(\sin_y_acc[23] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold199 (.A(\sin_y_acc[13] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold200 (.A(\cos_y_acc[8] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold201 (.A(\cos_x_acc[10] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0012_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold203 (.A(\cos_x_acc[12] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0014_),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold205 (.A(\hvsync_gen.hpos[1] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold206 (.A(\cos_x_acc[16] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0772_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold208 (.A(\cos_x_acc[14] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0016_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold210 (.A(\cos_x_acc[5] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0007_),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold212 (.A(\bayer_j[1] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold213 (.A(\sin_x_acc[5] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0061_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold215 (.A(\cos_x_acc[13] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold216 (.A(\cos_y_acc[20] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold217 (.A(\sin_x_acc[18] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold218 (.A(\sin_x_acc[16] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold219 (.A(\cos_x_acc[15] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold220 (.A(\cos_addr[0] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0039_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold222 (.A(\cos_x_acc[18] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold223 (.A(\cos_x_acc[8] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0011_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold225 (.A(\sin_x_acc[9] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0065_),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold227 (.A(\sin_x_acc[12] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0068_),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold229 (.A(\sin_x_acc[3] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0059_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold231 (.A(\sin_x_acc[1] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0858_),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0058_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold234 (.A(\sin_x_acc[14] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0070_),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold236 (.A(\cos_x_acc[3] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0635_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0006_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold239 (.A(\cos_x_acc[7] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold240 (.A(\cos_y_acc[22] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold241 (.A(\sin_x_acc[6] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold242 (.A(\cos_x_acc[1] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0598_),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0004_),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold245 (.A(\cos_x_acc[11] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold246 (.A(\sin_x_acc[10] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0067_),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold248 (.A(\sin_x_acc[4] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold249 (.A(\cos_x_acc[6] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold250 (.A(\sin_x_acc[8] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold251 (.A(\sin_x_acc[7] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold252 (.A(\cos_x_acc[5] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold253 (.A(\sin_x_acc[13] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold254 (.A(\cos_x_acc[2] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold255 (.A(\sin_x_acc[15] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold256 (.A(\cos_y_acc[22] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold257 (.A(\sin_y_acc[13] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold258 (.A(\bayer_j[0] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold259 (.A(\sin_y_acc[15] ),
    .X(net506));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_4 FILLER_13_224 ();
 sg13g2_fill_2 FILLER_13_228 ();
 sg13g2_fill_1 FILLER_13_234 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_163 ();
 sg13g2_decap_4 FILLER_14_170 ();
 sg13g2_decap_8 FILLER_14_187 ();
 sg13g2_decap_8 FILLER_14_194 ();
 sg13g2_decap_8 FILLER_14_201 ();
 sg13g2_decap_8 FILLER_14_208 ();
 sg13g2_decap_8 FILLER_14_215 ();
 sg13g2_fill_2 FILLER_14_222 ();
 sg13g2_fill_1 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_257 ();
 sg13g2_decap_8 FILLER_14_264 ();
 sg13g2_decap_8 FILLER_14_271 ();
 sg13g2_decap_8 FILLER_14_278 ();
 sg13g2_decap_8 FILLER_14_285 ();
 sg13g2_decap_8 FILLER_14_292 ();
 sg13g2_decap_8 FILLER_14_299 ();
 sg13g2_decap_8 FILLER_14_306 ();
 sg13g2_decap_8 FILLER_14_313 ();
 sg13g2_decap_8 FILLER_14_320 ();
 sg13g2_decap_8 FILLER_14_327 ();
 sg13g2_decap_8 FILLER_14_334 ();
 sg13g2_decap_8 FILLER_14_341 ();
 sg13g2_decap_8 FILLER_14_348 ();
 sg13g2_decap_8 FILLER_14_355 ();
 sg13g2_decap_8 FILLER_14_362 ();
 sg13g2_decap_8 FILLER_14_369 ();
 sg13g2_decap_8 FILLER_14_376 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_4 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_134 ();
 sg13g2_decap_4 FILLER_15_141 ();
 sg13g2_fill_1 FILLER_15_145 ();
 sg13g2_fill_1 FILLER_15_206 ();
 sg13g2_fill_2 FILLER_15_240 ();
 sg13g2_fill_1 FILLER_15_242 ();
 sg13g2_decap_8 FILLER_15_278 ();
 sg13g2_decap_8 FILLER_15_285 ();
 sg13g2_decap_8 FILLER_15_292 ();
 sg13g2_decap_8 FILLER_15_299 ();
 sg13g2_decap_8 FILLER_15_306 ();
 sg13g2_decap_8 FILLER_15_313 ();
 sg13g2_decap_8 FILLER_15_320 ();
 sg13g2_decap_8 FILLER_15_327 ();
 sg13g2_decap_8 FILLER_15_334 ();
 sg13g2_decap_8 FILLER_15_341 ();
 sg13g2_decap_8 FILLER_15_348 ();
 sg13g2_decap_8 FILLER_15_355 ();
 sg13g2_decap_8 FILLER_15_362 ();
 sg13g2_decap_8 FILLER_15_372 ();
 sg13g2_decap_8 FILLER_15_379 ();
 sg13g2_decap_8 FILLER_15_386 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_4 FILLER_16_119 ();
 sg13g2_fill_2 FILLER_16_123 ();
 sg13g2_fill_2 FILLER_16_153 ();
 sg13g2_fill_1 FILLER_16_155 ();
 sg13g2_decap_4 FILLER_16_184 ();
 sg13g2_fill_2 FILLER_16_188 ();
 sg13g2_fill_2 FILLER_16_248 ();
 sg13g2_fill_2 FILLER_16_268 ();
 sg13g2_decap_8 FILLER_16_274 ();
 sg13g2_decap_8 FILLER_16_281 ();
 sg13g2_decap_8 FILLER_16_288 ();
 sg13g2_decap_8 FILLER_16_295 ();
 sg13g2_decap_8 FILLER_16_302 ();
 sg13g2_decap_8 FILLER_16_309 ();
 sg13g2_decap_8 FILLER_16_316 ();
 sg13g2_decap_8 FILLER_16_323 ();
 sg13g2_decap_8 FILLER_16_330 ();
 sg13g2_decap_8 FILLER_16_337 ();
 sg13g2_decap_8 FILLER_16_344 ();
 sg13g2_decap_8 FILLER_16_351 ();
 sg13g2_decap_4 FILLER_16_358 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_decap_8 FILLER_16_388 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_4 FILLER_17_130 ();
 sg13g2_fill_1 FILLER_17_134 ();
 sg13g2_decap_8 FILLER_17_139 ();
 sg13g2_fill_1 FILLER_17_146 ();
 sg13g2_fill_1 FILLER_17_161 ();
 sg13g2_fill_1 FILLER_17_170 ();
 sg13g2_fill_2 FILLER_17_209 ();
 sg13g2_fill_1 FILLER_17_211 ();
 sg13g2_fill_2 FILLER_17_235 ();
 sg13g2_fill_1 FILLER_17_237 ();
 sg13g2_fill_1 FILLER_17_248 ();
 sg13g2_fill_2 FILLER_17_263 ();
 sg13g2_fill_1 FILLER_17_265 ();
 sg13g2_fill_2 FILLER_17_275 ();
 sg13g2_decap_8 FILLER_17_310 ();
 sg13g2_decap_8 FILLER_17_317 ();
 sg13g2_decap_8 FILLER_17_324 ();
 sg13g2_decap_8 FILLER_17_331 ();
 sg13g2_decap_4 FILLER_17_338 ();
 sg13g2_fill_2 FILLER_17_347 ();
 sg13g2_decap_8 FILLER_17_390 ();
 sg13g2_decap_8 FILLER_17_397 ();
 sg13g2_decap_4 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_fill_2 FILLER_18_84 ();
 sg13g2_fill_1 FILLER_18_86 ();
 sg13g2_decap_8 FILLER_18_108 ();
 sg13g2_fill_1 FILLER_18_115 ();
 sg13g2_fill_1 FILLER_18_167 ();
 sg13g2_decap_8 FILLER_18_172 ();
 sg13g2_decap_4 FILLER_18_179 ();
 sg13g2_fill_1 FILLER_18_194 ();
 sg13g2_fill_2 FILLER_18_200 ();
 sg13g2_decap_8 FILLER_18_237 ();
 sg13g2_decap_8 FILLER_18_244 ();
 sg13g2_fill_2 FILLER_18_251 ();
 sg13g2_fill_2 FILLER_18_262 ();
 sg13g2_fill_1 FILLER_18_264 ();
 sg13g2_fill_1 FILLER_18_302 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_fill_2 FILLER_18_329 ();
 sg13g2_fill_1 FILLER_18_331 ();
 sg13g2_fill_2 FILLER_18_352 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_4 FILLER_18_403 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_fill_2 FILLER_19_63 ();
 sg13g2_fill_1 FILLER_19_65 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_fill_2 FILLER_19_84 ();
 sg13g2_fill_1 FILLER_19_86 ();
 sg13g2_fill_2 FILLER_19_160 ();
 sg13g2_fill_1 FILLER_19_175 ();
 sg13g2_fill_2 FILLER_19_189 ();
 sg13g2_fill_1 FILLER_19_208 ();
 sg13g2_fill_2 FILLER_19_213 ();
 sg13g2_fill_1 FILLER_19_248 ();
 sg13g2_decap_4 FILLER_19_319 ();
 sg13g2_fill_2 FILLER_19_323 ();
 sg13g2_fill_2 FILLER_19_356 ();
 sg13g2_fill_1 FILLER_19_358 ();
 sg13g2_decap_8 FILLER_19_390 ();
 sg13g2_decap_8 FILLER_19_397 ();
 sg13g2_decap_4 FILLER_19_404 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_4 FILLER_20_56 ();
 sg13g2_fill_2 FILLER_20_88 ();
 sg13g2_fill_1 FILLER_20_208 ();
 sg13g2_fill_2 FILLER_20_241 ();
 sg13g2_fill_2 FILLER_20_290 ();
 sg13g2_fill_1 FILLER_20_292 ();
 sg13g2_fill_1 FILLER_20_324 ();
 sg13g2_fill_2 FILLER_20_337 ();
 sg13g2_fill_1 FILLER_20_339 ();
 sg13g2_decap_8 FILLER_20_345 ();
 sg13g2_decap_8 FILLER_20_352 ();
 sg13g2_fill_2 FILLER_20_359 ();
 sg13g2_fill_2 FILLER_20_369 ();
 sg13g2_fill_2 FILLER_20_375 ();
 sg13g2_fill_1 FILLER_20_377 ();
 sg13g2_decap_8 FILLER_20_386 ();
 sg13g2_fill_2 FILLER_20_393 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_4 FILLER_21_42 ();
 sg13g2_decap_4 FILLER_21_59 ();
 sg13g2_fill_2 FILLER_21_63 ();
 sg13g2_fill_2 FILLER_21_113 ();
 sg13g2_fill_1 FILLER_21_115 ();
 sg13g2_fill_2 FILLER_21_134 ();
 sg13g2_fill_2 FILLER_21_145 ();
 sg13g2_fill_2 FILLER_21_180 ();
 sg13g2_fill_2 FILLER_21_196 ();
 sg13g2_fill_2 FILLER_21_213 ();
 sg13g2_fill_2 FILLER_21_230 ();
 sg13g2_fill_2 FILLER_21_312 ();
 sg13g2_fill_1 FILLER_21_314 ();
 sg13g2_fill_2 FILLER_21_328 ();
 sg13g2_fill_1 FILLER_21_330 ();
 sg13g2_decap_8 FILLER_21_339 ();
 sg13g2_fill_2 FILLER_21_346 ();
 sg13g2_fill_1 FILLER_21_348 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_decap_4 FILLER_21_375 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_4 FILLER_22_49 ();
 sg13g2_fill_2 FILLER_22_53 ();
 sg13g2_fill_2 FILLER_22_88 ();
 sg13g2_fill_1 FILLER_22_99 ();
 sg13g2_decap_8 FILLER_22_120 ();
 sg13g2_decap_4 FILLER_22_127 ();
 sg13g2_fill_1 FILLER_22_131 ();
 sg13g2_fill_2 FILLER_22_135 ();
 sg13g2_decap_8 FILLER_22_150 ();
 sg13g2_decap_4 FILLER_22_157 ();
 sg13g2_fill_2 FILLER_22_187 ();
 sg13g2_fill_2 FILLER_22_225 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_4 FILLER_22_319 ();
 sg13g2_fill_2 FILLER_22_323 ();
 sg13g2_fill_1 FILLER_22_353 ();
 sg13g2_fill_2 FILLER_22_358 ();
 sg13g2_decap_8 FILLER_22_365 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_4 FILLER_23_42 ();
 sg13g2_fill_1 FILLER_23_46 ();
 sg13g2_decap_4 FILLER_23_104 ();
 sg13g2_fill_1 FILLER_23_121 ();
 sg13g2_fill_2 FILLER_23_144 ();
 sg13g2_fill_1 FILLER_23_146 ();
 sg13g2_decap_4 FILLER_23_151 ();
 sg13g2_fill_1 FILLER_23_155 ();
 sg13g2_decap_4 FILLER_23_174 ();
 sg13g2_fill_1 FILLER_23_178 ();
 sg13g2_decap_4 FILLER_23_183 ();
 sg13g2_fill_1 FILLER_23_216 ();
 sg13g2_fill_2 FILLER_23_230 ();
 sg13g2_fill_1 FILLER_23_232 ();
 sg13g2_fill_2 FILLER_23_254 ();
 sg13g2_decap_4 FILLER_23_319 ();
 sg13g2_fill_2 FILLER_23_381 ();
 sg13g2_fill_1 FILLER_23_383 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_fill_2 FILLER_24_35 ();
 sg13g2_fill_1 FILLER_24_37 ();
 sg13g2_fill_1 FILLER_24_127 ();
 sg13g2_fill_2 FILLER_24_149 ();
 sg13g2_fill_1 FILLER_24_211 ();
 sg13g2_decap_4 FILLER_24_221 ();
 sg13g2_fill_2 FILLER_24_247 ();
 sg13g2_fill_1 FILLER_24_249 ();
 sg13g2_fill_1 FILLER_24_327 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_fill_2 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_4 FILLER_24_385 ();
 sg13g2_fill_1 FILLER_24_389 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_fill_2 FILLER_25_28 ();
 sg13g2_fill_1 FILLER_25_30 ();
 sg13g2_fill_2 FILLER_25_64 ();
 sg13g2_fill_1 FILLER_25_66 ();
 sg13g2_decap_4 FILLER_25_88 ();
 sg13g2_fill_2 FILLER_25_92 ();
 sg13g2_fill_2 FILLER_25_104 ();
 sg13g2_decap_8 FILLER_25_145 ();
 sg13g2_decap_4 FILLER_25_152 ();
 sg13g2_fill_1 FILLER_25_156 ();
 sg13g2_decap_8 FILLER_25_171 ();
 sg13g2_decap_8 FILLER_25_178 ();
 sg13g2_fill_2 FILLER_25_185 ();
 sg13g2_fill_1 FILLER_25_187 ();
 sg13g2_fill_1 FILLER_25_197 ();
 sg13g2_fill_2 FILLER_25_215 ();
 sg13g2_fill_1 FILLER_25_217 ();
 sg13g2_fill_1 FILLER_25_237 ();
 sg13g2_fill_1 FILLER_25_243 ();
 sg13g2_fill_2 FILLER_25_309 ();
 sg13g2_fill_1 FILLER_25_311 ();
 sg13g2_fill_2 FILLER_25_332 ();
 sg13g2_fill_1 FILLER_25_334 ();
 sg13g2_fill_1 FILLER_25_346 ();
 sg13g2_decap_4 FILLER_25_350 ();
 sg13g2_fill_1 FILLER_25_354 ();
 sg13g2_fill_2 FILLER_25_360 ();
 sg13g2_fill_2 FILLER_25_367 ();
 sg13g2_fill_1 FILLER_25_369 ();
 sg13g2_decap_4 FILLER_25_378 ();
 sg13g2_fill_1 FILLER_25_382 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_fill_1 FILLER_26_35 ();
 sg13g2_fill_2 FILLER_26_53 ();
 sg13g2_fill_1 FILLER_26_59 ();
 sg13g2_decap_8 FILLER_26_69 ();
 sg13g2_fill_1 FILLER_26_76 ();
 sg13g2_decap_8 FILLER_26_90 ();
 sg13g2_decap_8 FILLER_26_97 ();
 sg13g2_decap_8 FILLER_26_104 ();
 sg13g2_fill_1 FILLER_26_127 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_176 ();
 sg13g2_decap_8 FILLER_26_183 ();
 sg13g2_decap_8 FILLER_26_190 ();
 sg13g2_decap_8 FILLER_26_197 ();
 sg13g2_fill_2 FILLER_26_204 ();
 sg13g2_fill_1 FILLER_26_206 ();
 sg13g2_decap_8 FILLER_26_246 ();
 sg13g2_fill_2 FILLER_26_253 ();
 sg13g2_fill_2 FILLER_26_259 ();
 sg13g2_fill_2 FILLER_26_265 ();
 sg13g2_fill_1 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_306 ();
 sg13g2_fill_2 FILLER_26_313 ();
 sg13g2_decap_8 FILLER_26_325 ();
 sg13g2_decap_8 FILLER_26_332 ();
 sg13g2_fill_1 FILLER_26_339 ();
 sg13g2_fill_2 FILLER_26_348 ();
 sg13g2_decap_4 FILLER_26_371 ();
 sg13g2_fill_1 FILLER_26_388 ();
 sg13g2_decap_8 FILLER_26_402 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_59 ();
 sg13g2_fill_1 FILLER_27_66 ();
 sg13g2_decap_8 FILLER_27_72 ();
 sg13g2_decap_8 FILLER_27_79 ();
 sg13g2_fill_1 FILLER_27_86 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_fill_2 FILLER_27_112 ();
 sg13g2_fill_1 FILLER_27_114 ();
 sg13g2_fill_2 FILLER_27_124 ();
 sg13g2_fill_1 FILLER_27_126 ();
 sg13g2_fill_2 FILLER_27_188 ();
 sg13g2_decap_8 FILLER_27_204 ();
 sg13g2_decap_4 FILLER_27_211 ();
 sg13g2_fill_1 FILLER_27_215 ();
 sg13g2_decap_4 FILLER_27_267 ();
 sg13g2_fill_1 FILLER_27_271 ();
 sg13g2_decap_4 FILLER_27_309 ();
 sg13g2_fill_2 FILLER_27_313 ();
 sg13g2_decap_8 FILLER_27_323 ();
 sg13g2_decap_8 FILLER_27_330 ();
 sg13g2_decap_8 FILLER_27_337 ();
 sg13g2_fill_1 FILLER_27_344 ();
 sg13g2_decap_8 FILLER_27_352 ();
 sg13g2_fill_1 FILLER_27_359 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_4 FILLER_27_385 ();
 sg13g2_fill_1 FILLER_27_393 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_fill_2 FILLER_28_21 ();
 sg13g2_fill_1 FILLER_28_23 ();
 sg13g2_decap_4 FILLER_28_52 ();
 sg13g2_fill_2 FILLER_28_61 ();
 sg13g2_fill_1 FILLER_28_127 ();
 sg13g2_fill_1 FILLER_28_146 ();
 sg13g2_fill_2 FILLER_28_160 ();
 sg13g2_decap_8 FILLER_28_218 ();
 sg13g2_fill_1 FILLER_28_225 ();
 sg13g2_decap_8 FILLER_28_230 ();
 sg13g2_decap_8 FILLER_28_237 ();
 sg13g2_fill_2 FILLER_28_244 ();
 sg13g2_fill_1 FILLER_28_282 ();
 sg13g2_decap_4 FILLER_28_334 ();
 sg13g2_fill_1 FILLER_28_338 ();
 sg13g2_fill_2 FILLER_28_357 ();
 sg13g2_fill_1 FILLER_28_359 ();
 sg13g2_decap_4 FILLER_28_364 ();
 sg13g2_fill_1 FILLER_28_368 ();
 sg13g2_fill_2 FILLER_28_381 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_4 FILLER_29_14 ();
 sg13g2_fill_2 FILLER_29_18 ();
 sg13g2_fill_2 FILLER_29_42 ();
 sg13g2_fill_1 FILLER_29_44 ();
 sg13g2_fill_2 FILLER_29_62 ();
 sg13g2_decap_4 FILLER_29_103 ();
 sg13g2_fill_2 FILLER_29_107 ();
 sg13g2_fill_1 FILLER_29_146 ();
 sg13g2_fill_1 FILLER_29_163 ();
 sg13g2_fill_2 FILLER_29_174 ();
 sg13g2_fill_1 FILLER_29_194 ();
 sg13g2_decap_8 FILLER_29_219 ();
 sg13g2_decap_8 FILLER_29_226 ();
 sg13g2_fill_2 FILLER_29_233 ();
 sg13g2_fill_2 FILLER_29_239 ();
 sg13g2_fill_2 FILLER_29_251 ();
 sg13g2_fill_1 FILLER_29_293 ();
 sg13g2_fill_1 FILLER_29_308 ();
 sg13g2_fill_1 FILLER_29_325 ();
 sg13g2_fill_1 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_29_368 ();
 sg13g2_decap_8 FILLER_29_375 ();
 sg13g2_decap_4 FILLER_29_382 ();
 sg13g2_fill_1 FILLER_29_386 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_fill_2 FILLER_30_28 ();
 sg13g2_fill_2 FILLER_30_52 ();
 sg13g2_fill_1 FILLER_30_54 ();
 sg13g2_fill_2 FILLER_30_63 ();
 sg13g2_fill_1 FILLER_30_65 ();
 sg13g2_decap_4 FILLER_30_87 ();
 sg13g2_fill_1 FILLER_30_98 ();
 sg13g2_fill_1 FILLER_30_126 ();
 sg13g2_decap_4 FILLER_30_174 ();
 sg13g2_fill_1 FILLER_30_178 ();
 sg13g2_fill_2 FILLER_30_228 ();
 sg13g2_fill_2 FILLER_30_258 ();
 sg13g2_fill_1 FILLER_30_260 ();
 sg13g2_decap_4 FILLER_30_292 ();
 sg13g2_fill_1 FILLER_30_296 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_decap_8 FILLER_30_328 ();
 sg13g2_fill_2 FILLER_30_335 ();
 sg13g2_fill_1 FILLER_30_350 ();
 sg13g2_fill_2 FILLER_30_358 ();
 sg13g2_fill_1 FILLER_30_360 ();
 sg13g2_fill_1 FILLER_30_366 ();
 sg13g2_decap_8 FILLER_30_380 ();
 sg13g2_fill_2 FILLER_30_387 ();
 sg13g2_fill_1 FILLER_30_389 ();
 sg13g2_fill_2 FILLER_30_395 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_fill_2 FILLER_31_43 ();
 sg13g2_decap_4 FILLER_31_54 ();
 sg13g2_fill_2 FILLER_31_58 ();
 sg13g2_fill_1 FILLER_31_64 ();
 sg13g2_fill_1 FILLER_31_69 ();
 sg13g2_fill_1 FILLER_31_83 ();
 sg13g2_decap_4 FILLER_31_107 ();
 sg13g2_fill_2 FILLER_31_156 ();
 sg13g2_fill_2 FILLER_31_166 ();
 sg13g2_fill_2 FILLER_31_205 ();
 sg13g2_fill_1 FILLER_31_207 ();
 sg13g2_fill_2 FILLER_31_246 ();
 sg13g2_fill_1 FILLER_31_269 ();
 sg13g2_fill_2 FILLER_31_279 ();
 sg13g2_fill_2 FILLER_31_288 ();
 sg13g2_fill_1 FILLER_31_290 ();
 sg13g2_decap_4 FILLER_31_313 ();
 sg13g2_decap_4 FILLER_31_336 ();
 sg13g2_fill_2 FILLER_31_340 ();
 sg13g2_fill_2 FILLER_31_350 ();
 sg13g2_fill_1 FILLER_31_352 ();
 sg13g2_fill_2 FILLER_31_371 ();
 sg13g2_fill_1 FILLER_31_373 ();
 sg13g2_decap_4 FILLER_31_386 ();
 sg13g2_fill_2 FILLER_31_390 ();
 sg13g2_decap_8 FILLER_31_396 ();
 sg13g2_decap_4 FILLER_31_403 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_14 ();
 sg13g2_fill_1 FILLER_32_53 ();
 sg13g2_fill_2 FILLER_32_100 ();
 sg13g2_fill_2 FILLER_32_115 ();
 sg13g2_fill_1 FILLER_32_117 ();
 sg13g2_fill_2 FILLER_32_122 ();
 sg13g2_fill_2 FILLER_32_134 ();
 sg13g2_decap_8 FILLER_32_172 ();
 sg13g2_fill_2 FILLER_32_179 ();
 sg13g2_fill_1 FILLER_32_181 ();
 sg13g2_decap_8 FILLER_32_186 ();
 sg13g2_fill_2 FILLER_32_197 ();
 sg13g2_fill_1 FILLER_32_199 ();
 sg13g2_fill_2 FILLER_32_244 ();
 sg13g2_fill_1 FILLER_32_246 ();
 sg13g2_fill_2 FILLER_32_306 ();
 sg13g2_fill_1 FILLER_32_308 ();
 sg13g2_decap_4 FILLER_32_346 ();
 sg13g2_fill_2 FILLER_32_350 ();
 sg13g2_fill_2 FILLER_32_360 ();
 sg13g2_fill_2 FILLER_32_385 ();
 sg13g2_fill_1 FILLER_32_387 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_25 ();
 sg13g2_fill_1 FILLER_33_39 ();
 sg13g2_decap_4 FILLER_33_49 ();
 sg13g2_fill_2 FILLER_33_63 ();
 sg13g2_fill_2 FILLER_33_72 ();
 sg13g2_fill_1 FILLER_33_74 ();
 sg13g2_fill_1 FILLER_33_112 ();
 sg13g2_fill_1 FILLER_33_137 ();
 sg13g2_fill_2 FILLER_33_151 ();
 sg13g2_fill_1 FILLER_33_153 ();
 sg13g2_fill_2 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_179 ();
 sg13g2_decap_8 FILLER_33_186 ();
 sg13g2_decap_8 FILLER_33_198 ();
 sg13g2_decap_8 FILLER_33_205 ();
 sg13g2_decap_4 FILLER_33_212 ();
 sg13g2_fill_2 FILLER_33_216 ();
 sg13g2_fill_1 FILLER_33_230 ();
 sg13g2_fill_1 FILLER_33_245 ();
 sg13g2_fill_2 FILLER_33_298 ();
 sg13g2_fill_1 FILLER_33_312 ();
 sg13g2_decap_4 FILLER_33_338 ();
 sg13g2_fill_1 FILLER_33_342 ();
 sg13g2_fill_2 FILLER_33_355 ();
 sg13g2_decap_8 FILLER_33_368 ();
 sg13g2_fill_2 FILLER_33_393 ();
 sg13g2_fill_1 FILLER_33_395 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_fill_1 FILLER_34_44 ();
 sg13g2_fill_1 FILLER_34_84 ();
 sg13g2_fill_1 FILLER_34_93 ();
 sg13g2_fill_1 FILLER_34_99 ();
 sg13g2_fill_2 FILLER_34_113 ();
 sg13g2_fill_1 FILLER_34_157 ();
 sg13g2_decap_4 FILLER_34_184 ();
 sg13g2_fill_2 FILLER_34_188 ();
 sg13g2_fill_1 FILLER_34_198 ();
 sg13g2_decap_4 FILLER_34_220 ();
 sg13g2_fill_1 FILLER_34_228 ();
 sg13g2_decap_4 FILLER_34_242 ();
 sg13g2_fill_2 FILLER_34_251 ();
 sg13g2_fill_1 FILLER_34_253 ();
 sg13g2_fill_2 FILLER_34_299 ();
 sg13g2_decap_4 FILLER_34_308 ();
 sg13g2_decap_8 FILLER_34_320 ();
 sg13g2_decap_8 FILLER_34_327 ();
 sg13g2_decap_8 FILLER_34_334 ();
 sg13g2_decap_8 FILLER_34_341 ();
 sg13g2_fill_1 FILLER_34_348 ();
 sg13g2_fill_1 FILLER_34_374 ();
 sg13g2_fill_2 FILLER_34_388 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_fill_2 FILLER_35_21 ();
 sg13g2_fill_1 FILLER_35_23 ();
 sg13g2_fill_2 FILLER_35_28 ();
 sg13g2_fill_1 FILLER_35_30 ();
 sg13g2_fill_2 FILLER_35_61 ();
 sg13g2_fill_1 FILLER_35_97 ();
 sg13g2_fill_2 FILLER_35_126 ();
 sg13g2_fill_2 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_fill_2 FILLER_35_182 ();
 sg13g2_fill_1 FILLER_35_184 ();
 sg13g2_fill_1 FILLER_35_193 ();
 sg13g2_fill_2 FILLER_35_261 ();
 sg13g2_fill_2 FILLER_35_267 ();
 sg13g2_decap_4 FILLER_35_286 ();
 sg13g2_decap_8 FILLER_35_307 ();
 sg13g2_decap_8 FILLER_35_314 ();
 sg13g2_fill_2 FILLER_35_325 ();
 sg13g2_decap_8 FILLER_35_336 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_fill_2 FILLER_35_350 ();
 sg13g2_fill_1 FILLER_35_352 ();
 sg13g2_fill_2 FILLER_35_374 ();
 sg13g2_fill_2 FILLER_35_380 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_4 FILLER_36_14 ();
 sg13g2_fill_1 FILLER_36_18 ();
 sg13g2_fill_2 FILLER_36_47 ();
 sg13g2_fill_1 FILLER_36_49 ();
 sg13g2_fill_1 FILLER_36_71 ();
 sg13g2_fill_2 FILLER_36_90 ();
 sg13g2_decap_8 FILLER_36_100 ();
 sg13g2_fill_1 FILLER_36_107 ();
 sg13g2_decap_4 FILLER_36_117 ();
 sg13g2_fill_1 FILLER_36_121 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_fill_1 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_150 ();
 sg13g2_decap_8 FILLER_36_157 ();
 sg13g2_fill_1 FILLER_36_164 ();
 sg13g2_decap_4 FILLER_36_198 ();
 sg13g2_fill_2 FILLER_36_207 ();
 sg13g2_fill_2 FILLER_36_270 ();
 sg13g2_fill_2 FILLER_36_290 ();
 sg13g2_fill_1 FILLER_36_292 ();
 sg13g2_decap_8 FILLER_36_340 ();
 sg13g2_fill_2 FILLER_36_347 ();
 sg13g2_decap_4 FILLER_36_354 ();
 sg13g2_fill_1 FILLER_36_358 ();
 sg13g2_decap_8 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_378 ();
 sg13g2_fill_2 FILLER_36_385 ();
 sg13g2_fill_2 FILLER_36_394 ();
 sg13g2_fill_1 FILLER_36_396 ();
 sg13g2_decap_8 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_fill_2 FILLER_37_21 ();
 sg13g2_fill_1 FILLER_37_23 ();
 sg13g2_fill_1 FILLER_37_46 ();
 sg13g2_fill_2 FILLER_37_54 ();
 sg13g2_fill_1 FILLER_37_56 ();
 sg13g2_fill_1 FILLER_37_80 ();
 sg13g2_decap_8 FILLER_37_129 ();
 sg13g2_decap_8 FILLER_37_136 ();
 sg13g2_decap_8 FILLER_37_143 ();
 sg13g2_decap_4 FILLER_37_177 ();
 sg13g2_fill_2 FILLER_37_194 ();
 sg13g2_fill_2 FILLER_37_207 ();
 sg13g2_fill_1 FILLER_37_209 ();
 sg13g2_decap_4 FILLER_37_213 ();
 sg13g2_fill_2 FILLER_37_217 ();
 sg13g2_fill_2 FILLER_37_228 ();
 sg13g2_fill_2 FILLER_37_242 ();
 sg13g2_fill_1 FILLER_37_260 ();
 sg13g2_decap_4 FILLER_37_283 ();
 sg13g2_fill_1 FILLER_37_287 ();
 sg13g2_fill_2 FILLER_37_316 ();
 sg13g2_fill_2 FILLER_37_345 ();
 sg13g2_fill_2 FILLER_37_362 ();
 sg13g2_fill_1 FILLER_37_364 ();
 sg13g2_decap_4 FILLER_37_386 ();
 sg13g2_fill_2 FILLER_37_390 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_4 FILLER_38_14 ();
 sg13g2_fill_2 FILLER_38_18 ();
 sg13g2_decap_4 FILLER_38_57 ();
 sg13g2_fill_2 FILLER_38_61 ();
 sg13g2_fill_2 FILLER_38_67 ();
 sg13g2_fill_1 FILLER_38_76 ();
 sg13g2_fill_2 FILLER_38_81 ();
 sg13g2_fill_2 FILLER_38_92 ();
 sg13g2_fill_2 FILLER_38_102 ();
 sg13g2_fill_2 FILLER_38_120 ();
 sg13g2_fill_2 FILLER_38_143 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_4 FILLER_38_168 ();
 sg13g2_fill_1 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_181 ();
 sg13g2_fill_2 FILLER_38_202 ();
 sg13g2_fill_1 FILLER_38_204 ();
 sg13g2_decap_4 FILLER_38_218 ();
 sg13g2_fill_1 FILLER_38_222 ();
 sg13g2_fill_2 FILLER_38_228 ();
 sg13g2_fill_1 FILLER_38_233 ();
 sg13g2_fill_1 FILLER_38_246 ();
 sg13g2_fill_1 FILLER_38_287 ();
 sg13g2_fill_1 FILLER_38_306 ();
 sg13g2_fill_2 FILLER_38_319 ();
 sg13g2_fill_1 FILLER_38_321 ();
 sg13g2_decap_4 FILLER_38_327 ();
 sg13g2_fill_1 FILLER_38_335 ();
 sg13g2_decap_8 FILLER_38_351 ();
 sg13g2_decap_8 FILLER_38_358 ();
 sg13g2_decap_8 FILLER_38_365 ();
 sg13g2_decap_4 FILLER_38_372 ();
 sg13g2_fill_1 FILLER_38_388 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_4 FILLER_39_7 ();
 sg13g2_fill_2 FILLER_39_11 ();
 sg13g2_fill_2 FILLER_39_26 ();
 sg13g2_fill_2 FILLER_39_36 ();
 sg13g2_fill_1 FILLER_39_52 ();
 sg13g2_decap_8 FILLER_39_85 ();
 sg13g2_fill_1 FILLER_39_92 ();
 sg13g2_decap_4 FILLER_39_106 ();
 sg13g2_fill_1 FILLER_39_146 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_decap_4 FILLER_39_182 ();
 sg13g2_fill_2 FILLER_39_194 ();
 sg13g2_fill_1 FILLER_39_196 ();
 sg13g2_decap_4 FILLER_39_205 ();
 sg13g2_fill_1 FILLER_39_209 ();
 sg13g2_fill_1 FILLER_39_218 ();
 sg13g2_decap_8 FILLER_39_239 ();
 sg13g2_decap_4 FILLER_39_246 ();
 sg13g2_fill_2 FILLER_39_250 ();
 sg13g2_fill_1 FILLER_39_264 ();
 sg13g2_decap_8 FILLER_39_299 ();
 sg13g2_decap_8 FILLER_39_311 ();
 sg13g2_fill_2 FILLER_39_318 ();
 sg13g2_fill_1 FILLER_39_320 ();
 sg13g2_fill_1 FILLER_39_329 ();
 sg13g2_fill_2 FILLER_39_345 ();
 sg13g2_decap_8 FILLER_39_352 ();
 sg13g2_decap_8 FILLER_39_359 ();
 sg13g2_fill_2 FILLER_39_366 ();
 sg13g2_fill_1 FILLER_39_376 ();
 sg13g2_fill_2 FILLER_39_394 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_7 ();
 sg13g2_fill_2 FILLER_40_46 ();
 sg13g2_fill_1 FILLER_40_48 ();
 sg13g2_fill_2 FILLER_40_66 ();
 sg13g2_decap_8 FILLER_40_94 ();
 sg13g2_decap_8 FILLER_40_101 ();
 sg13g2_decap_8 FILLER_40_108 ();
 sg13g2_fill_1 FILLER_40_119 ();
 sg13g2_decap_4 FILLER_40_123 ();
 sg13g2_fill_1 FILLER_40_127 ();
 sg13g2_fill_2 FILLER_40_132 ();
 sg13g2_fill_2 FILLER_40_175 ();
 sg13g2_fill_1 FILLER_40_177 ();
 sg13g2_fill_1 FILLER_40_199 ();
 sg13g2_decap_8 FILLER_40_209 ();
 sg13g2_decap_4 FILLER_40_216 ();
 sg13g2_fill_1 FILLER_40_220 ();
 sg13g2_decap_8 FILLER_40_238 ();
 sg13g2_decap_8 FILLER_40_245 ();
 sg13g2_fill_1 FILLER_40_252 ();
 sg13g2_fill_1 FILLER_40_265 ();
 sg13g2_fill_2 FILLER_40_280 ();
 sg13g2_decap_8 FILLER_40_295 ();
 sg13g2_decap_4 FILLER_40_302 ();
 sg13g2_decap_8 FILLER_40_310 ();
 sg13g2_fill_2 FILLER_40_317 ();
 sg13g2_fill_1 FILLER_40_319 ();
 sg13g2_fill_2 FILLER_40_340 ();
 sg13g2_fill_1 FILLER_40_356 ();
 sg13g2_fill_2 FILLER_40_378 ();
 sg13g2_fill_1 FILLER_40_380 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_fill_2 FILLER_41_21 ();
 sg13g2_fill_1 FILLER_41_23 ();
 sg13g2_decap_4 FILLER_41_29 ();
 sg13g2_fill_1 FILLER_41_33 ();
 sg13g2_decap_4 FILLER_41_55 ();
 sg13g2_fill_2 FILLER_41_59 ();
 sg13g2_fill_1 FILLER_41_65 ();
 sg13g2_fill_1 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_fill_1 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_fill_2 FILLER_41_147 ();
 sg13g2_fill_1 FILLER_41_177 ();
 sg13g2_decap_4 FILLER_41_211 ();
 sg13g2_fill_1 FILLER_41_215 ();
 sg13g2_decap_8 FILLER_41_241 ();
 sg13g2_fill_1 FILLER_41_248 ();
 sg13g2_fill_1 FILLER_41_306 ();
 sg13g2_decap_8 FILLER_41_320 ();
 sg13g2_fill_1 FILLER_41_357 ();
 sg13g2_decap_8 FILLER_41_379 ();
 sg13g2_decap_8 FILLER_41_402 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_fill_1 FILLER_42_28 ();
 sg13g2_decap_4 FILLER_42_33 ();
 sg13g2_fill_2 FILLER_42_37 ();
 sg13g2_decap_4 FILLER_42_49 ();
 sg13g2_fill_1 FILLER_42_53 ();
 sg13g2_fill_1 FILLER_42_80 ();
 sg13g2_decap_8 FILLER_42_114 ();
 sg13g2_fill_2 FILLER_42_121 ();
 sg13g2_fill_2 FILLER_42_127 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_fill_1 FILLER_42_158 ();
 sg13g2_fill_1 FILLER_42_167 ();
 sg13g2_fill_2 FILLER_42_182 ();
 sg13g2_fill_1 FILLER_42_184 ();
 sg13g2_decap_8 FILLER_42_198 ();
 sg13g2_fill_1 FILLER_42_247 ();
 sg13g2_fill_2 FILLER_42_264 ();
 sg13g2_fill_1 FILLER_42_295 ();
 sg13g2_decap_8 FILLER_42_324 ();
 sg13g2_decap_8 FILLER_42_331 ();
 sg13g2_decap_4 FILLER_42_338 ();
 sg13g2_fill_2 FILLER_42_346 ();
 sg13g2_fill_1 FILLER_42_357 ();
 sg13g2_fill_1 FILLER_42_362 ();
 sg13g2_fill_2 FILLER_42_376 ();
 sg13g2_fill_1 FILLER_42_378 ();
 sg13g2_decap_4 FILLER_42_387 ();
 sg13g2_fill_1 FILLER_42_391 ();
 sg13g2_decap_4 FILLER_42_404 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_fill_2 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_2 ();
 sg13g2_fill_1 FILLER_43_30 ();
 sg13g2_fill_2 FILLER_43_43 ();
 sg13g2_fill_1 FILLER_43_45 ();
 sg13g2_decap_8 FILLER_43_54 ();
 sg13g2_decap_4 FILLER_43_69 ();
 sg13g2_fill_1 FILLER_43_73 ();
 sg13g2_fill_1 FILLER_43_78 ();
 sg13g2_decap_4 FILLER_43_87 ();
 sg13g2_fill_2 FILLER_43_95 ();
 sg13g2_fill_1 FILLER_43_97 ();
 sg13g2_fill_2 FILLER_43_107 ();
 sg13g2_fill_1 FILLER_43_109 ();
 sg13g2_fill_2 FILLER_43_118 ();
 sg13g2_fill_2 FILLER_43_130 ();
 sg13g2_decap_8 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_158 ();
 sg13g2_decap_8 FILLER_43_165 ();
 sg13g2_fill_2 FILLER_43_172 ();
 sg13g2_fill_2 FILLER_43_219 ();
 sg13g2_fill_2 FILLER_43_263 ();
 sg13g2_fill_1 FILLER_43_273 ();
 sg13g2_fill_1 FILLER_43_282 ();
 sg13g2_decap_8 FILLER_43_328 ();
 sg13g2_decap_4 FILLER_43_335 ();
 sg13g2_fill_2 FILLER_43_339 ();
 sg13g2_decap_8 FILLER_43_364 ();
 sg13g2_decap_8 FILLER_43_383 ();
 sg13g2_decap_4 FILLER_43_390 ();
 sg13g2_fill_2 FILLER_43_394 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_2 ();
 sg13g2_fill_2 FILLER_44_16 ();
 sg13g2_fill_2 FILLER_44_28 ();
 sg13g2_fill_2 FILLER_44_47 ();
 sg13g2_decap_8 FILLER_44_92 ();
 sg13g2_fill_1 FILLER_44_99 ();
 sg13g2_fill_1 FILLER_44_132 ();
 sg13g2_fill_2 FILLER_44_139 ();
 sg13g2_fill_2 FILLER_44_149 ();
 sg13g2_fill_1 FILLER_44_151 ();
 sg13g2_decap_4 FILLER_44_162 ();
 sg13g2_fill_1 FILLER_44_193 ();
 sg13g2_fill_2 FILLER_44_230 ();
 sg13g2_fill_1 FILLER_44_232 ();
 sg13g2_fill_1 FILLER_44_250 ();
 sg13g2_decap_4 FILLER_44_307 ();
 sg13g2_fill_2 FILLER_44_311 ();
 sg13g2_decap_4 FILLER_44_325 ();
 sg13g2_fill_1 FILLER_44_329 ();
 sg13g2_decap_8 FILLER_44_334 ();
 sg13g2_fill_1 FILLER_44_341 ();
 sg13g2_decap_4 FILLER_44_369 ();
 sg13g2_fill_1 FILLER_44_373 ();
 sg13g2_decap_8 FILLER_44_389 ();
 sg13g2_decap_8 FILLER_44_396 ();
 sg13g2_decap_4 FILLER_44_403 ();
 sg13g2_fill_2 FILLER_44_407 ();
 sg13g2_fill_1 FILLER_45_0 ();
 sg13g2_decap_4 FILLER_45_68 ();
 sg13g2_fill_1 FILLER_45_72 ();
 sg13g2_decap_8 FILLER_45_101 ();
 sg13g2_fill_2 FILLER_45_127 ();
 sg13g2_fill_2 FILLER_45_145 ();
 sg13g2_fill_2 FILLER_45_192 ();
 sg13g2_fill_1 FILLER_45_194 ();
 sg13g2_decap_4 FILLER_45_210 ();
 sg13g2_fill_2 FILLER_45_214 ();
 sg13g2_fill_1 FILLER_45_244 ();
 sg13g2_decap_8 FILLER_45_254 ();
 sg13g2_decap_8 FILLER_45_261 ();
 sg13g2_decap_4 FILLER_45_268 ();
 sg13g2_decap_4 FILLER_45_291 ();
 sg13g2_decap_8 FILLER_45_300 ();
 sg13g2_decap_4 FILLER_45_307 ();
 sg13g2_fill_2 FILLER_45_323 ();
 sg13g2_fill_1 FILLER_45_340 ();
 sg13g2_fill_1 FILLER_45_346 ();
 sg13g2_fill_2 FILLER_45_366 ();
 sg13g2_fill_1 FILLER_45_377 ();
 sg13g2_decap_4 FILLER_45_382 ();
 sg13g2_fill_2 FILLER_45_391 ();
 sg13g2_fill_1 FILLER_45_393 ();
 sg13g2_decap_4 FILLER_45_404 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_4 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_4 ();
 sg13g2_fill_2 FILLER_46_16 ();
 sg13g2_fill_1 FILLER_46_18 ();
 sg13g2_fill_2 FILLER_46_35 ();
 sg13g2_fill_1 FILLER_46_37 ();
 sg13g2_decap_4 FILLER_46_84 ();
 sg13g2_fill_2 FILLER_46_108 ();
 sg13g2_fill_1 FILLER_46_110 ();
 sg13g2_fill_1 FILLER_46_133 ();
 sg13g2_fill_1 FILLER_46_144 ();
 sg13g2_decap_8 FILLER_46_165 ();
 sg13g2_fill_2 FILLER_46_172 ();
 sg13g2_decap_4 FILLER_46_215 ();
 sg13g2_fill_2 FILLER_46_219 ();
 sg13g2_decap_4 FILLER_46_225 ();
 sg13g2_fill_2 FILLER_46_229 ();
 sg13g2_decap_8 FILLER_46_236 ();
 sg13g2_decap_8 FILLER_46_243 ();
 sg13g2_decap_4 FILLER_46_250 ();
 sg13g2_fill_2 FILLER_46_254 ();
 sg13g2_decap_8 FILLER_46_281 ();
 sg13g2_fill_1 FILLER_46_296 ();
 sg13g2_fill_2 FILLER_46_305 ();
 sg13g2_fill_2 FILLER_46_348 ();
 sg13g2_fill_2 FILLER_46_358 ();
 sg13g2_fill_2 FILLER_46_373 ();
 sg13g2_fill_2 FILLER_46_407 ();
 sg13g2_fill_1 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_22 ();
 sg13g2_decap_4 FILLER_47_34 ();
 sg13g2_fill_1 FILLER_47_46 ();
 sg13g2_fill_2 FILLER_47_57 ();
 sg13g2_fill_1 FILLER_47_92 ();
 sg13g2_fill_1 FILLER_47_104 ();
 sg13g2_fill_2 FILLER_47_130 ();
 sg13g2_decap_4 FILLER_47_146 ();
 sg13g2_decap_4 FILLER_47_176 ();
 sg13g2_fill_1 FILLER_47_180 ();
 sg13g2_decap_8 FILLER_47_189 ();
 sg13g2_fill_2 FILLER_47_196 ();
 sg13g2_decap_8 FILLER_47_206 ();
 sg13g2_fill_1 FILLER_47_221 ();
 sg13g2_decap_4 FILLER_47_230 ();
 sg13g2_decap_8 FILLER_47_242 ();
 sg13g2_decap_4 FILLER_47_249 ();
 sg13g2_decap_4 FILLER_47_305 ();
 sg13g2_fill_2 FILLER_47_328 ();
 sg13g2_fill_1 FILLER_47_330 ();
 sg13g2_fill_2 FILLER_47_338 ();
 sg13g2_fill_2 FILLER_47_348 ();
 sg13g2_fill_1 FILLER_47_350 ();
 sg13g2_fill_2 FILLER_47_356 ();
 sg13g2_fill_1 FILLER_47_358 ();
 sg13g2_fill_1 FILLER_47_370 ();
 sg13g2_decap_8 FILLER_47_376 ();
 sg13g2_fill_2 FILLER_47_383 ();
 sg13g2_decap_4 FILLER_47_404 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_16 ();
 sg13g2_fill_2 FILLER_48_26 ();
 sg13g2_fill_1 FILLER_48_28 ();
 sg13g2_decap_4 FILLER_48_37 ();
 sg13g2_decap_8 FILLER_48_52 ();
 sg13g2_decap_4 FILLER_48_59 ();
 sg13g2_fill_1 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_83 ();
 sg13g2_decap_8 FILLER_48_90 ();
 sg13g2_decap_4 FILLER_48_97 ();
 sg13g2_decap_4 FILLER_48_116 ();
 sg13g2_fill_2 FILLER_48_120 ();
 sg13g2_decap_4 FILLER_48_137 ();
 sg13g2_fill_2 FILLER_48_141 ();
 sg13g2_fill_2 FILLER_48_148 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_fill_2 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_176 ();
 sg13g2_decap_4 FILLER_48_183 ();
 sg13g2_fill_2 FILLER_48_187 ();
 sg13g2_decap_8 FILLER_48_218 ();
 sg13g2_decap_8 FILLER_48_225 ();
 sg13g2_decap_8 FILLER_48_232 ();
 sg13g2_fill_2 FILLER_48_239 ();
 sg13g2_fill_1 FILLER_48_241 ();
 sg13g2_fill_2 FILLER_48_318 ();
 sg13g2_fill_1 FILLER_48_320 ();
 sg13g2_decap_8 FILLER_48_339 ();
 sg13g2_decap_8 FILLER_48_346 ();
 sg13g2_decap_4 FILLER_48_353 ();
 sg13g2_fill_2 FILLER_48_361 ();
 sg13g2_decap_8 FILLER_48_367 ();
 sg13g2_decap_8 FILLER_48_374 ();
 sg13g2_fill_1 FILLER_48_381 ();
 sg13g2_fill_2 FILLER_48_406 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_fill_1 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_29 ();
 sg13g2_fill_2 FILLER_49_39 ();
 sg13g2_fill_1 FILLER_49_41 ();
 sg13g2_decap_4 FILLER_49_50 ();
 sg13g2_fill_1 FILLER_49_54 ();
 sg13g2_fill_1 FILLER_49_73 ();
 sg13g2_decap_8 FILLER_49_93 ();
 sg13g2_decap_4 FILLER_49_100 ();
 sg13g2_fill_1 FILLER_49_104 ();
 sg13g2_fill_2 FILLER_49_130 ();
 sg13g2_fill_1 FILLER_49_132 ();
 sg13g2_fill_2 FILLER_49_146 ();
 sg13g2_decap_8 FILLER_49_160 ();
 sg13g2_fill_2 FILLER_49_193 ();
 sg13g2_fill_1 FILLER_49_195 ();
 sg13g2_decap_8 FILLER_49_214 ();
 sg13g2_fill_2 FILLER_49_221 ();
 sg13g2_decap_4 FILLER_49_231 ();
 sg13g2_fill_1 FILLER_49_248 ();
 sg13g2_decap_4 FILLER_49_257 ();
 sg13g2_decap_8 FILLER_49_265 ();
 sg13g2_fill_2 FILLER_49_272 ();
 sg13g2_fill_2 FILLER_49_286 ();
 sg13g2_fill_1 FILLER_49_293 ();
 sg13g2_fill_2 FILLER_49_304 ();
 sg13g2_fill_1 FILLER_49_306 ();
 sg13g2_decap_4 FILLER_49_334 ();
 sg13g2_fill_1 FILLER_49_338 ();
 sg13g2_decap_4 FILLER_49_343 ();
 sg13g2_fill_1 FILLER_49_347 ();
 sg13g2_decap_8 FILLER_49_356 ();
 sg13g2_decap_8 FILLER_49_363 ();
 sg13g2_decap_8 FILLER_49_370 ();
 sg13g2_fill_1 FILLER_49_377 ();
 sg13g2_fill_1 FILLER_49_392 ();
 sg13g2_decap_8 FILLER_49_398 ();
 sg13g2_decap_4 FILLER_49_405 ();
 sg13g2_decap_4 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_4 ();
 sg13g2_decap_4 FILLER_50_10 ();
 sg13g2_fill_1 FILLER_50_14 ();
 sg13g2_decap_4 FILLER_50_20 ();
 sg13g2_fill_1 FILLER_50_24 ();
 sg13g2_fill_2 FILLER_50_42 ();
 sg13g2_decap_4 FILLER_50_56 ();
 sg13g2_fill_2 FILLER_50_96 ();
 sg13g2_fill_1 FILLER_50_98 ();
 sg13g2_decap_8 FILLER_50_120 ();
 sg13g2_fill_2 FILLER_50_127 ();
 sg13g2_fill_1 FILLER_50_147 ();
 sg13g2_decap_8 FILLER_50_164 ();
 sg13g2_fill_1 FILLER_50_171 ();
 sg13g2_decap_4 FILLER_50_180 ();
 sg13g2_fill_1 FILLER_50_216 ();
 sg13g2_fill_1 FILLER_50_235 ();
 sg13g2_fill_1 FILLER_50_244 ();
 sg13g2_decap_8 FILLER_50_258 ();
 sg13g2_decap_8 FILLER_50_270 ();
 sg13g2_decap_4 FILLER_50_290 ();
 sg13g2_decap_4 FILLER_50_299 ();
 sg13g2_fill_1 FILLER_50_303 ();
 sg13g2_fill_1 FILLER_50_340 ();
 sg13g2_fill_2 FILLER_50_357 ();
 sg13g2_fill_2 FILLER_50_378 ();
 sg13g2_fill_1 FILLER_50_380 ();
 sg13g2_decap_8 FILLER_50_394 ();
 sg13g2_decap_8 FILLER_50_401 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_4 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_4 ();
 sg13g2_decap_4 FILLER_51_10 ();
 sg13g2_fill_2 FILLER_51_34 ();
 sg13g2_fill_1 FILLER_51_58 ();
 sg13g2_fill_2 FILLER_51_68 ();
 sg13g2_fill_1 FILLER_51_70 ();
 sg13g2_fill_1 FILLER_51_93 ();
 sg13g2_fill_1 FILLER_51_118 ();
 sg13g2_fill_1 FILLER_51_134 ();
 sg13g2_fill_2 FILLER_51_144 ();
 sg13g2_fill_2 FILLER_51_190 ();
 sg13g2_fill_1 FILLER_51_217 ();
 sg13g2_fill_1 FILLER_51_223 ();
 sg13g2_fill_1 FILLER_51_256 ();
 sg13g2_fill_1 FILLER_51_301 ();
 sg13g2_fill_2 FILLER_51_326 ();
 sg13g2_fill_2 FILLER_51_337 ();
 sg13g2_fill_2 FILLER_51_346 ();
 sg13g2_fill_1 FILLER_51_348 ();
 sg13g2_fill_2 FILLER_51_383 ();
 sg13g2_decap_8 FILLER_51_397 ();
 sg13g2_decap_4 FILLER_51_404 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_fill_1 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_32 ();
 sg13g2_decap_8 FILLER_52_72 ();
 sg13g2_decap_8 FILLER_52_79 ();
 sg13g2_decap_8 FILLER_52_86 ();
 sg13g2_fill_2 FILLER_52_93 ();
 sg13g2_fill_1 FILLER_52_95 ();
 sg13g2_decap_4 FILLER_52_124 ();
 sg13g2_fill_2 FILLER_52_128 ();
 sg13g2_fill_2 FILLER_52_135 ();
 sg13g2_fill_1 FILLER_52_164 ();
 sg13g2_decap_8 FILLER_52_179 ();
 sg13g2_fill_2 FILLER_52_186 ();
 sg13g2_fill_2 FILLER_52_195 ();
 sg13g2_fill_1 FILLER_52_197 ();
 sg13g2_fill_2 FILLER_52_210 ();
 sg13g2_fill_2 FILLER_52_217 ();
 sg13g2_fill_2 FILLER_52_224 ();
 sg13g2_fill_1 FILLER_52_226 ();
 sg13g2_decap_4 FILLER_52_231 ();
 sg13g2_fill_1 FILLER_52_235 ();
 sg13g2_fill_1 FILLER_52_264 ();
 sg13g2_decap_4 FILLER_52_275 ();
 sg13g2_fill_1 FILLER_52_279 ();
 sg13g2_decap_4 FILLER_52_295 ();
 sg13g2_fill_1 FILLER_52_299 ();
 sg13g2_fill_1 FILLER_52_305 ();
 sg13g2_fill_2 FILLER_52_311 ();
 sg13g2_fill_2 FILLER_52_342 ();
 sg13g2_fill_1 FILLER_52_344 ();
 sg13g2_fill_2 FILLER_52_350 ();
 sg13g2_fill_1 FILLER_52_352 ();
 sg13g2_decap_4 FILLER_52_364 ();
 sg13g2_fill_1 FILLER_52_368 ();
 sg13g2_fill_1 FILLER_52_375 ();
 sg13g2_fill_2 FILLER_52_381 ();
 sg13g2_decap_8 FILLER_52_388 ();
 sg13g2_decap_8 FILLER_52_395 ();
 sg13g2_decap_8 FILLER_52_402 ();
 sg13g2_decap_4 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_4 ();
 sg13g2_decap_8 FILLER_53_38 ();
 sg13g2_decap_8 FILLER_53_54 ();
 sg13g2_fill_2 FILLER_53_61 ();
 sg13g2_fill_1 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_75 ();
 sg13g2_decap_8 FILLER_53_82 ();
 sg13g2_decap_8 FILLER_53_89 ();
 sg13g2_fill_1 FILLER_53_96 ();
 sg13g2_fill_1 FILLER_53_110 ();
 sg13g2_decap_4 FILLER_53_116 ();
 sg13g2_fill_2 FILLER_53_120 ();
 sg13g2_fill_2 FILLER_53_131 ();
 sg13g2_fill_2 FILLER_53_138 ();
 sg13g2_fill_1 FILLER_53_140 ();
 sg13g2_decap_4 FILLER_53_147 ();
 sg13g2_fill_1 FILLER_53_151 ();
 sg13g2_fill_1 FILLER_53_171 ();
 sg13g2_decap_4 FILLER_53_185 ();
 sg13g2_decap_8 FILLER_53_202 ();
 sg13g2_decap_8 FILLER_53_209 ();
 sg13g2_decap_4 FILLER_53_221 ();
 sg13g2_fill_2 FILLER_53_225 ();
 sg13g2_decap_8 FILLER_53_243 ();
 sg13g2_decap_8 FILLER_53_254 ();
 sg13g2_fill_2 FILLER_53_261 ();
 sg13g2_fill_1 FILLER_53_263 ();
 sg13g2_decap_8 FILLER_53_268 ();
 sg13g2_decap_8 FILLER_53_275 ();
 sg13g2_fill_1 FILLER_53_282 ();
 sg13g2_decap_8 FILLER_53_288 ();
 sg13g2_fill_2 FILLER_53_295 ();
 sg13g2_fill_1 FILLER_53_297 ();
 sg13g2_decap_4 FILLER_53_319 ();
 sg13g2_fill_2 FILLER_53_328 ();
 sg13g2_fill_2 FILLER_53_344 ();
 sg13g2_fill_1 FILLER_53_346 ();
 sg13g2_decap_8 FILLER_53_367 ();
 sg13g2_decap_8 FILLER_53_374 ();
 sg13g2_decap_8 FILLER_53_381 ();
 sg13g2_decap_8 FILLER_53_388 ();
 sg13g2_decap_8 FILLER_53_395 ();
 sg13g2_decap_8 FILLER_53_402 ();
 sg13g2_fill_2 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_2 ();
 sg13g2_decap_8 FILLER_54_47 ();
 sg13g2_fill_2 FILLER_54_63 ();
 sg13g2_decap_4 FILLER_54_74 ();
 sg13g2_fill_2 FILLER_54_78 ();
 sg13g2_decap_8 FILLER_54_85 ();
 sg13g2_fill_1 FILLER_54_92 ();
 sg13g2_decap_4 FILLER_54_136 ();
 sg13g2_fill_1 FILLER_54_140 ();
 sg13g2_decap_4 FILLER_54_156 ();
 sg13g2_fill_2 FILLER_54_160 ();
 sg13g2_decap_4 FILLER_54_177 ();
 sg13g2_fill_2 FILLER_54_181 ();
 sg13g2_decap_8 FILLER_54_209 ();
 sg13g2_decap_8 FILLER_54_216 ();
 sg13g2_decap_8 FILLER_54_223 ();
 sg13g2_decap_8 FILLER_54_252 ();
 sg13g2_decap_8 FILLER_54_259 ();
 sg13g2_decap_4 FILLER_54_266 ();
 sg13g2_fill_1 FILLER_54_287 ();
 sg13g2_decap_8 FILLER_54_296 ();
 sg13g2_fill_1 FILLER_54_303 ();
 sg13g2_fill_1 FILLER_54_336 ();
 sg13g2_decap_8 FILLER_54_365 ();
 sg13g2_decap_8 FILLER_54_372 ();
 sg13g2_decap_8 FILLER_54_379 ();
 sg13g2_decap_8 FILLER_54_386 ();
 sg13g2_decap_8 FILLER_54_393 ();
 sg13g2_decap_8 FILLER_54_400 ();
 sg13g2_fill_2 FILLER_54_407 ();
 sg13g2_fill_1 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_38 ();
 sg13g2_fill_2 FILLER_55_48 ();
 sg13g2_fill_2 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_93 ();
 sg13g2_fill_1 FILLER_55_100 ();
 sg13g2_fill_2 FILLER_55_121 ();
 sg13g2_fill_2 FILLER_55_127 ();
 sg13g2_decap_8 FILLER_55_138 ();
 sg13g2_decap_8 FILLER_55_145 ();
 sg13g2_decap_8 FILLER_55_152 ();
 sg13g2_decap_8 FILLER_55_159 ();
 sg13g2_fill_1 FILLER_55_166 ();
 sg13g2_decap_4 FILLER_55_171 ();
 sg13g2_fill_1 FILLER_55_175 ();
 sg13g2_fill_2 FILLER_55_211 ();
 sg13g2_decap_8 FILLER_55_252 ();
 sg13g2_decap_4 FILLER_55_277 ();
 sg13g2_fill_1 FILLER_55_281 ();
 sg13g2_decap_4 FILLER_55_319 ();
 sg13g2_fill_1 FILLER_55_323 ();
 sg13g2_decap_8 FILLER_55_332 ();
 sg13g2_decap_4 FILLER_55_339 ();
 sg13g2_fill_2 FILLER_55_343 ();
 sg13g2_fill_2 FILLER_55_351 ();
 sg13g2_fill_1 FILLER_55_353 ();
 sg13g2_decap_8 FILLER_55_393 ();
 sg13g2_decap_8 FILLER_55_400 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_30 ();
 sg13g2_decap_8 FILLER_56_53 ();
 sg13g2_fill_2 FILLER_56_60 ();
 sg13g2_fill_2 FILLER_56_67 ();
 sg13g2_fill_1 FILLER_56_69 ();
 sg13g2_decap_4 FILLER_56_98 ();
 sg13g2_fill_2 FILLER_56_102 ();
 sg13g2_fill_2 FILLER_56_117 ();
 sg13g2_fill_2 FILLER_56_127 ();
 sg13g2_fill_1 FILLER_56_155 ();
 sg13g2_fill_2 FILLER_56_161 ();
 sg13g2_fill_1 FILLER_56_163 ();
 sg13g2_decap_8 FILLER_56_175 ();
 sg13g2_decap_4 FILLER_56_182 ();
 sg13g2_fill_2 FILLER_56_202 ();
 sg13g2_fill_1 FILLER_56_204 ();
 sg13g2_decap_4 FILLER_56_228 ();
 sg13g2_decap_4 FILLER_56_236 ();
 sg13g2_fill_2 FILLER_56_240 ();
 sg13g2_fill_1 FILLER_56_253 ();
 sg13g2_fill_1 FILLER_56_275 ();
 sg13g2_fill_2 FILLER_56_288 ();
 sg13g2_decap_4 FILLER_56_298 ();
 sg13g2_fill_1 FILLER_56_302 ();
 sg13g2_decap_4 FILLER_56_307 ();
 sg13g2_fill_1 FILLER_56_311 ();
 sg13g2_decap_8 FILLER_56_333 ();
 sg13g2_decap_4 FILLER_56_340 ();
 sg13g2_fill_2 FILLER_56_344 ();
 sg13g2_fill_2 FILLER_56_354 ();
 sg13g2_fill_1 FILLER_56_356 ();
 sg13g2_decap_8 FILLER_56_394 ();
 sg13g2_decap_8 FILLER_56_401 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_fill_1 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_29 ();
 sg13g2_fill_2 FILLER_57_44 ();
 sg13g2_fill_1 FILLER_57_46 ();
 sg13g2_decap_4 FILLER_57_59 ();
 sg13g2_fill_2 FILLER_57_63 ();
 sg13g2_fill_1 FILLER_57_82 ();
 sg13g2_fill_2 FILLER_57_97 ();
 sg13g2_fill_1 FILLER_57_99 ();
 sg13g2_decap_4 FILLER_57_143 ();
 sg13g2_fill_1 FILLER_57_162 ();
 sg13g2_decap_8 FILLER_57_176 ();
 sg13g2_decap_8 FILLER_57_183 ();
 sg13g2_fill_2 FILLER_57_202 ();
 sg13g2_fill_1 FILLER_57_209 ();
 sg13g2_decap_8 FILLER_57_248 ();
 sg13g2_fill_2 FILLER_57_255 ();
 sg13g2_decap_4 FILLER_57_340 ();
 sg13g2_fill_2 FILLER_57_344 ();
 sg13g2_decap_4 FILLER_57_404 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_decap_4 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_4 ();
 sg13g2_decap_4 FILLER_58_10 ();
 sg13g2_fill_2 FILLER_58_14 ();
 sg13g2_fill_1 FILLER_58_83 ();
 sg13g2_decap_4 FILLER_58_97 ();
 sg13g2_fill_1 FILLER_58_101 ();
 sg13g2_fill_2 FILLER_58_134 ();
 sg13g2_decap_8 FILLER_58_147 ();
 sg13g2_fill_1 FILLER_58_154 ();
 sg13g2_fill_1 FILLER_58_183 ();
 sg13g2_decap_4 FILLER_58_193 ();
 sg13g2_fill_1 FILLER_58_197 ();
 sg13g2_decap_4 FILLER_58_207 ();
 sg13g2_fill_2 FILLER_58_211 ();
 sg13g2_fill_2 FILLER_58_230 ();
 sg13g2_fill_1 FILLER_58_232 ();
 sg13g2_fill_2 FILLER_58_258 ();
 sg13g2_fill_1 FILLER_58_260 ();
 sg13g2_fill_2 FILLER_58_269 ();
 sg13g2_decap_8 FILLER_58_276 ();
 sg13g2_fill_1 FILLER_58_283 ();
 sg13g2_fill_2 FILLER_58_288 ();
 sg13g2_fill_1 FILLER_58_290 ();
 sg13g2_fill_2 FILLER_58_296 ();
 sg13g2_fill_1 FILLER_58_298 ();
 sg13g2_decap_4 FILLER_58_314 ();
 sg13g2_fill_1 FILLER_58_318 ();
 sg13g2_decap_8 FILLER_58_382 ();
 sg13g2_decap_8 FILLER_58_389 ();
 sg13g2_decap_8 FILLER_58_396 ();
 sg13g2_decap_4 FILLER_58_403 ();
 sg13g2_fill_2 FILLER_58_407 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_fill_1 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_62 ();
 sg13g2_fill_2 FILLER_59_69 ();
 sg13g2_fill_1 FILLER_59_71 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_4 FILLER_59_89 ();
 sg13g2_fill_1 FILLER_59_93 ();
 sg13g2_fill_1 FILLER_59_126 ();
 sg13g2_fill_2 FILLER_59_132 ();
 sg13g2_decap_4 FILLER_59_142 ();
 sg13g2_fill_2 FILLER_59_156 ();
 sg13g2_fill_2 FILLER_59_167 ();
 sg13g2_fill_1 FILLER_59_169 ();
 sg13g2_fill_1 FILLER_59_183 ();
 sg13g2_decap_8 FILLER_59_197 ();
 sg13g2_decap_8 FILLER_59_204 ();
 sg13g2_decap_4 FILLER_59_211 ();
 sg13g2_fill_2 FILLER_59_215 ();
 sg13g2_decap_8 FILLER_59_227 ();
 sg13g2_fill_2 FILLER_59_234 ();
 sg13g2_fill_1 FILLER_59_236 ();
 sg13g2_decap_8 FILLER_59_247 ();
 sg13g2_decap_8 FILLER_59_254 ();
 sg13g2_decap_4 FILLER_59_261 ();
 sg13g2_fill_2 FILLER_59_265 ();
 sg13g2_fill_2 FILLER_59_271 ();
 sg13g2_fill_1 FILLER_59_273 ();
 sg13g2_fill_2 FILLER_59_278 ();
 sg13g2_decap_8 FILLER_59_285 ();
 sg13g2_decap_8 FILLER_59_292 ();
 sg13g2_decap_8 FILLER_59_299 ();
 sg13g2_decap_8 FILLER_59_306 ();
 sg13g2_decap_4 FILLER_59_313 ();
 sg13g2_fill_2 FILLER_59_358 ();
 sg13g2_fill_1 FILLER_59_360 ();
 sg13g2_fill_2 FILLER_59_365 ();
 sg13g2_fill_1 FILLER_59_367 ();
 sg13g2_decap_8 FILLER_59_372 ();
 sg13g2_decap_8 FILLER_59_379 ();
 sg13g2_decap_8 FILLER_59_386 ();
 sg13g2_decap_8 FILLER_59_393 ();
 sg13g2_decap_8 FILLER_59_400 ();
 sg13g2_fill_2 FILLER_59_407 ();
 sg13g2_decap_4 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_4 ();
 sg13g2_decap_4 FILLER_60_18 ();
 sg13g2_fill_1 FILLER_60_22 ();
 sg13g2_decap_4 FILLER_60_55 ();
 sg13g2_fill_2 FILLER_60_73 ();
 sg13g2_fill_1 FILLER_60_75 ();
 sg13g2_fill_2 FILLER_60_95 ();
 sg13g2_fill_1 FILLER_60_97 ();
 sg13g2_fill_2 FILLER_60_128 ();
 sg13g2_fill_1 FILLER_60_130 ();
 sg13g2_decap_8 FILLER_60_145 ();
 sg13g2_fill_1 FILLER_60_196 ();
 sg13g2_decap_8 FILLER_60_211 ();
 sg13g2_decap_8 FILLER_60_218 ();
 sg13g2_decap_8 FILLER_60_225 ();
 sg13g2_fill_2 FILLER_60_232 ();
 sg13g2_fill_1 FILLER_60_234 ();
 sg13g2_decap_8 FILLER_60_239 ();
 sg13g2_fill_2 FILLER_60_246 ();
 sg13g2_fill_1 FILLER_60_248 ();
 sg13g2_decap_8 FILLER_60_254 ();
 sg13g2_fill_1 FILLER_60_274 ();
 sg13g2_fill_2 FILLER_60_295 ();
 sg13g2_fill_1 FILLER_60_297 ();
 sg13g2_fill_1 FILLER_60_338 ();
 sg13g2_fill_1 FILLER_60_352 ();
 sg13g2_decap_8 FILLER_60_390 ();
 sg13g2_decap_8 FILLER_60_397 ();
 sg13g2_decap_4 FILLER_60_404 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_fill_1 FILLER_61_0 ();
 sg13g2_decap_4 FILLER_61_46 ();
 sg13g2_fill_1 FILLER_61_122 ();
 sg13g2_fill_2 FILLER_61_133 ();
 sg13g2_fill_1 FILLER_61_135 ();
 sg13g2_decap_8 FILLER_61_154 ();
 sg13g2_fill_1 FILLER_61_161 ();
 sg13g2_decap_8 FILLER_61_175 ();
 sg13g2_decap_8 FILLER_61_182 ();
 sg13g2_fill_2 FILLER_61_189 ();
 sg13g2_fill_1 FILLER_61_191 ();
 sg13g2_decap_4 FILLER_61_213 ();
 sg13g2_fill_1 FILLER_61_217 ();
 sg13g2_fill_2 FILLER_61_222 ();
 sg13g2_decap_8 FILLER_61_232 ();
 sg13g2_fill_2 FILLER_61_239 ();
 sg13g2_decap_4 FILLER_61_294 ();
 sg13g2_fill_2 FILLER_61_322 ();
 sg13g2_decap_8 FILLER_61_398 ();
 sg13g2_decap_4 FILLER_61_405 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_4 FILLER_62_14 ();
 sg13g2_decap_4 FILLER_62_45 ();
 sg13g2_fill_2 FILLER_62_57 ();
 sg13g2_fill_1 FILLER_62_59 ();
 sg13g2_fill_2 FILLER_62_73 ();
 sg13g2_fill_1 FILLER_62_75 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_fill_1 FILLER_62_98 ();
 sg13g2_fill_1 FILLER_62_133 ();
 sg13g2_fill_1 FILLER_62_142 ();
 sg13g2_decap_8 FILLER_62_170 ();
 sg13g2_decap_8 FILLER_62_177 ();
 sg13g2_decap_4 FILLER_62_200 ();
 sg13g2_fill_1 FILLER_62_204 ();
 sg13g2_decap_4 FILLER_62_232 ();
 sg13g2_fill_2 FILLER_62_236 ();
 sg13g2_fill_1 FILLER_62_319 ();
 sg13g2_fill_2 FILLER_62_361 ();
 sg13g2_fill_1 FILLER_62_363 ();
 sg13g2_decap_8 FILLER_62_395 ();
 sg13g2_decap_8 FILLER_62_402 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_4 FILLER_63_47 ();
 sg13g2_fill_2 FILLER_63_61 ();
 sg13g2_fill_1 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_73 ();
 sg13g2_fill_1 FILLER_63_84 ();
 sg13g2_fill_2 FILLER_63_119 ();
 sg13g2_fill_1 FILLER_63_145 ();
 sg13g2_decap_8 FILLER_63_170 ();
 sg13g2_fill_2 FILLER_63_185 ();
 sg13g2_decap_4 FILLER_63_200 ();
 sg13g2_fill_2 FILLER_63_204 ();
 sg13g2_fill_2 FILLER_63_224 ();
 sg13g2_decap_4 FILLER_63_244 ();
 sg13g2_decap_4 FILLER_63_257 ();
 sg13g2_fill_2 FILLER_63_261 ();
 sg13g2_fill_2 FILLER_63_272 ();
 sg13g2_fill_1 FILLER_63_274 ();
 sg13g2_decap_8 FILLER_63_287 ();
 sg13g2_decap_4 FILLER_63_294 ();
 sg13g2_fill_2 FILLER_63_298 ();
 sg13g2_fill_2 FILLER_63_349 ();
 sg13g2_decap_8 FILLER_63_388 ();
 sg13g2_decap_8 FILLER_63_395 ();
 sg13g2_decap_8 FILLER_63_402 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_4 FILLER_64_25 ();
 sg13g2_decap_8 FILLER_64_62 ();
 sg13g2_fill_1 FILLER_64_69 ();
 sg13g2_fill_2 FILLER_64_100 ();
 sg13g2_fill_1 FILLER_64_102 ();
 sg13g2_decap_4 FILLER_64_116 ();
 sg13g2_fill_1 FILLER_64_120 ();
 sg13g2_fill_1 FILLER_64_142 ();
 sg13g2_fill_2 FILLER_64_156 ();
 sg13g2_fill_1 FILLER_64_158 ();
 sg13g2_decap_4 FILLER_64_199 ();
 sg13g2_fill_2 FILLER_64_203 ();
 sg13g2_decap_8 FILLER_64_260 ();
 sg13g2_fill_2 FILLER_64_267 ();
 sg13g2_decap_8 FILLER_64_278 ();
 sg13g2_decap_8 FILLER_64_285 ();
 sg13g2_decap_4 FILLER_64_292 ();
 sg13g2_fill_2 FILLER_64_330 ();
 sg13g2_fill_1 FILLER_64_362 ();
 sg13g2_decap_8 FILLER_64_386 ();
 sg13g2_decap_8 FILLER_64_393 ();
 sg13g2_decap_8 FILLER_64_400 ();
 sg13g2_fill_2 FILLER_64_407 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_107 ();
 sg13g2_decap_8 FILLER_65_114 ();
 sg13g2_fill_1 FILLER_65_121 ();
 sg13g2_decap_8 FILLER_65_135 ();
 sg13g2_fill_1 FILLER_65_142 ();
 sg13g2_fill_2 FILLER_65_249 ();
 sg13g2_decap_8 FILLER_65_260 ();
 sg13g2_decap_8 FILLER_65_267 ();
 sg13g2_decap_8 FILLER_65_274 ();
 sg13g2_decap_4 FILLER_65_281 ();
 sg13g2_fill_1 FILLER_65_285 ();
 sg13g2_fill_2 FILLER_65_319 ();
 sg13g2_fill_1 FILLER_65_356 ();
 sg13g2_decap_8 FILLER_65_390 ();
 sg13g2_decap_8 FILLER_65_397 ();
 sg13g2_decap_4 FILLER_65_404 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_4 FILLER_66_14 ();
 sg13g2_fill_2 FILLER_66_18 ();
 sg13g2_fill_2 FILLER_66_130 ();
 sg13g2_fill_1 FILLER_66_132 ();
 sg13g2_fill_1 FILLER_66_141 ();
 sg13g2_fill_2 FILLER_66_181 ();
 sg13g2_fill_1 FILLER_66_183 ();
 sg13g2_fill_1 FILLER_66_202 ();
 sg13g2_fill_1 FILLER_66_207 ();
 sg13g2_fill_2 FILLER_66_213 ();
 sg13g2_fill_1 FILLER_66_224 ();
 sg13g2_fill_2 FILLER_66_246 ();
 sg13g2_fill_1 FILLER_66_256 ();
 sg13g2_decap_4 FILLER_66_285 ();
 sg13g2_fill_2 FILLER_66_318 ();
 sg13g2_fill_1 FILLER_66_343 ();
 sg13g2_decap_8 FILLER_66_383 ();
 sg13g2_decap_8 FILLER_66_390 ();
 sg13g2_decap_8 FILLER_66_397 ();
 sg13g2_decap_4 FILLER_66_404 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_4 FILLER_67_21 ();
 sg13g2_fill_2 FILLER_67_25 ();
 sg13g2_decap_8 FILLER_67_31 ();
 sg13g2_decap_4 FILLER_67_38 ();
 sg13g2_fill_2 FILLER_67_164 ();
 sg13g2_fill_1 FILLER_67_197 ();
 sg13g2_fill_2 FILLER_67_278 ();
 sg13g2_fill_2 FILLER_67_293 ();
 sg13g2_decap_8 FILLER_67_382 ();
 sg13g2_decap_8 FILLER_67_389 ();
 sg13g2_decap_8 FILLER_67_396 ();
 sg13g2_decap_4 FILLER_67_403 ();
 sg13g2_fill_2 FILLER_67_407 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_4 FILLER_68_42 ();
 sg13g2_fill_2 FILLER_68_46 ();
 sg13g2_fill_2 FILLER_68_61 ();
 sg13g2_decap_8 FILLER_68_85 ();
 sg13g2_fill_1 FILLER_68_204 ();
 sg13g2_fill_2 FILLER_68_222 ();
 sg13g2_fill_2 FILLER_68_246 ();
 sg13g2_fill_1 FILLER_68_260 ();
 sg13g2_fill_2 FILLER_68_302 ();
 sg13g2_fill_1 FILLER_68_304 ();
 sg13g2_decap_4 FILLER_68_310 ();
 sg13g2_decap_8 FILLER_68_398 ();
 sg13g2_decap_4 FILLER_68_405 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_4 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_78 ();
 sg13g2_decap_8 FILLER_69_85 ();
 sg13g2_fill_2 FILLER_69_92 ();
 sg13g2_fill_1 FILLER_69_151 ();
 sg13g2_fill_1 FILLER_69_251 ();
 sg13g2_fill_1 FILLER_69_264 ();
 sg13g2_fill_2 FILLER_69_304 ();
 sg13g2_fill_1 FILLER_69_306 ();
 sg13g2_fill_2 FILLER_69_312 ();
 sg13g2_fill_2 FILLER_69_319 ();
 sg13g2_fill_1 FILLER_69_326 ();
 sg13g2_fill_1 FILLER_69_336 ();
 sg13g2_fill_1 FILLER_69_342 ();
 sg13g2_fill_2 FILLER_69_362 ();
 sg13g2_fill_2 FILLER_69_369 ();
 sg13g2_decap_8 FILLER_69_384 ();
 sg13g2_decap_8 FILLER_69_391 ();
 sg13g2_decap_8 FILLER_69_398 ();
 sg13g2_decap_4 FILLER_69_405 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_fill_2 FILLER_70_91 ();
 sg13g2_fill_1 FILLER_70_93 ();
 sg13g2_fill_2 FILLER_70_107 ();
 sg13g2_fill_1 FILLER_70_109 ();
 sg13g2_fill_2 FILLER_70_201 ();
 sg13g2_fill_2 FILLER_70_212 ();
 sg13g2_fill_1 FILLER_70_214 ();
 sg13g2_fill_2 FILLER_70_262 ();
 sg13g2_decap_4 FILLER_70_301 ();
 sg13g2_fill_1 FILLER_70_321 ();
 sg13g2_decap_4 FILLER_70_364 ();
 sg13g2_decap_8 FILLER_70_373 ();
 sg13g2_fill_1 FILLER_70_380 ();
 sg13g2_decap_8 FILLER_70_390 ();
 sg13g2_decap_8 FILLER_70_397 ();
 sg13g2_decap_4 FILLER_70_404 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_fill_1 FILLER_71_91 ();
 sg13g2_decap_4 FILLER_71_96 ();
 sg13g2_fill_1 FILLER_71_100 ();
 sg13g2_fill_1 FILLER_71_110 ();
 sg13g2_fill_2 FILLER_71_120 ();
 sg13g2_fill_1 FILLER_71_122 ();
 sg13g2_fill_1 FILLER_71_222 ();
 sg13g2_fill_1 FILLER_71_227 ();
 sg13g2_fill_1 FILLER_71_233 ();
 sg13g2_fill_1 FILLER_71_283 ();
 sg13g2_fill_2 FILLER_71_293 ();
 sg13g2_fill_1 FILLER_71_295 ();
 sg13g2_fill_1 FILLER_71_331 ();
 sg13g2_decap_8 FILLER_71_390 ();
 sg13g2_decap_8 FILLER_71_397 ();
 sg13g2_decap_4 FILLER_71_404 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_fill_2 FILLER_72_84 ();
 sg13g2_fill_2 FILLER_72_132 ();
 sg13g2_fill_2 FILLER_72_167 ();
 sg13g2_fill_2 FILLER_72_188 ();
 sg13g2_fill_1 FILLER_72_208 ();
 sg13g2_fill_2 FILLER_72_218 ();
 sg13g2_fill_2 FILLER_72_225 ();
 sg13g2_fill_2 FILLER_72_279 ();
 sg13g2_fill_1 FILLER_72_281 ();
 sg13g2_fill_1 FILLER_72_295 ();
 sg13g2_fill_1 FILLER_72_350 ();
 sg13g2_decap_8 FILLER_72_377 ();
 sg13g2_decap_8 FILLER_72_384 ();
 sg13g2_decap_8 FILLER_72_391 ();
 sg13g2_decap_8 FILLER_72_398 ();
 sg13g2_decap_4 FILLER_72_405 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_fill_1 FILLER_73_161 ();
 sg13g2_fill_2 FILLER_73_171 ();
 sg13g2_fill_2 FILLER_73_177 ();
 sg13g2_fill_2 FILLER_73_324 ();
 sg13g2_fill_2 FILLER_73_335 ();
 sg13g2_fill_1 FILLER_73_363 ();
 sg13g2_decap_8 FILLER_73_377 ();
 sg13g2_decap_8 FILLER_73_384 ();
 sg13g2_decap_8 FILLER_73_391 ();
 sg13g2_decap_8 FILLER_73_398 ();
 sg13g2_decap_4 FILLER_73_405 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_4 FILLER_74_84 ();
 sg13g2_fill_1 FILLER_74_88 ();
 sg13g2_fill_1 FILLER_74_145 ();
 sg13g2_fill_2 FILLER_74_153 ();
 sg13g2_fill_1 FILLER_74_189 ();
 sg13g2_fill_2 FILLER_74_199 ();
 sg13g2_fill_1 FILLER_74_236 ();
 sg13g2_fill_1 FILLER_74_265 ();
 sg13g2_fill_2 FILLER_74_317 ();
 sg13g2_fill_2 FILLER_74_342 ();
 sg13g2_fill_2 FILLER_74_360 ();
 sg13g2_decap_8 FILLER_74_389 ();
 sg13g2_decap_8 FILLER_74_396 ();
 sg13g2_decap_4 FILLER_74_403 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_fill_1 FILLER_75_98 ();
 sg13g2_fill_1 FILLER_75_103 ();
 sg13g2_fill_1 FILLER_75_117 ();
 sg13g2_fill_2 FILLER_75_136 ();
 sg13g2_fill_1 FILLER_75_156 ();
 sg13g2_fill_2 FILLER_75_189 ();
 sg13g2_fill_1 FILLER_75_198 ();
 sg13g2_fill_1 FILLER_75_204 ();
 sg13g2_fill_2 FILLER_75_218 ();
 sg13g2_fill_2 FILLER_75_238 ();
 sg13g2_fill_1 FILLER_75_240 ();
 sg13g2_fill_1 FILLER_75_309 ();
 sg13g2_fill_1 FILLER_75_324 ();
 sg13g2_fill_2 FILLER_75_338 ();
 sg13g2_fill_1 FILLER_75_349 ();
 sg13g2_decap_8 FILLER_75_393 ();
 sg13g2_decap_8 FILLER_75_400 ();
 sg13g2_fill_2 FILLER_75_407 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_4 FILLER_76_105 ();
 sg13g2_fill_1 FILLER_76_144 ();
 sg13g2_fill_2 FILLER_76_168 ();
 sg13g2_fill_2 FILLER_76_198 ();
 sg13g2_fill_1 FILLER_76_200 ();
 sg13g2_fill_2 FILLER_76_247 ();
 sg13g2_fill_1 FILLER_76_249 ();
 sg13g2_fill_1 FILLER_76_259 ();
 sg13g2_fill_1 FILLER_76_283 ();
 sg13g2_fill_2 FILLER_76_293 ();
 sg13g2_fill_1 FILLER_76_345 ();
 sg13g2_decap_8 FILLER_76_383 ();
 sg13g2_decap_8 FILLER_76_390 ();
 sg13g2_decap_8 FILLER_76_397 ();
 sg13g2_decap_4 FILLER_76_404 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_fill_2 FILLER_77_182 ();
 sg13g2_fill_1 FILLER_77_184 ();
 sg13g2_fill_1 FILLER_77_241 ();
 sg13g2_decap_8 FILLER_77_378 ();
 sg13g2_decap_8 FILLER_77_385 ();
 sg13g2_decap_8 FILLER_77_392 ();
 sg13g2_decap_8 FILLER_77_399 ();
 sg13g2_fill_2 FILLER_77_406 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_4 FILLER_78_105 ();
 sg13g2_fill_2 FILLER_78_109 ();
 sg13g2_fill_2 FILLER_78_141 ();
 sg13g2_fill_1 FILLER_78_156 ();
 sg13g2_fill_2 FILLER_78_213 ();
 sg13g2_fill_1 FILLER_78_238 ();
 sg13g2_fill_2 FILLER_78_334 ();
 sg13g2_decap_8 FILLER_78_368 ();
 sg13g2_decap_8 FILLER_78_375 ();
 sg13g2_decap_8 FILLER_78_382 ();
 sg13g2_decap_8 FILLER_78_389 ();
 sg13g2_decap_8 FILLER_78_396 ();
 sg13g2_decap_4 FILLER_78_403 ();
 sg13g2_fill_2 FILLER_78_407 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_fill_1 FILLER_79_112 ();
 sg13g2_fill_1 FILLER_79_158 ();
 sg13g2_fill_1 FILLER_79_263 ();
 sg13g2_fill_1 FILLER_79_319 ();
 sg13g2_decap_8 FILLER_79_360 ();
 sg13g2_decap_8 FILLER_79_367 ();
 sg13g2_decap_8 FILLER_79_374 ();
 sg13g2_decap_8 FILLER_79_381 ();
 sg13g2_decap_8 FILLER_79_388 ();
 sg13g2_decap_8 FILLER_79_395 ();
 sg13g2_decap_8 FILLER_79_402 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_fill_2 FILLER_80_92 ();
 sg13g2_decap_8 FILLER_80_221 ();
 sg13g2_fill_2 FILLER_80_228 ();
 sg13g2_fill_1 FILLER_80_230 ();
 sg13g2_fill_2 FILLER_80_243 ();
 sg13g2_fill_2 FILLER_80_250 ();
 sg13g2_fill_2 FILLER_80_262 ();
 sg13g2_fill_2 FILLER_80_289 ();
 sg13g2_decap_8 FILLER_80_352 ();
 sg13g2_decap_8 FILLER_80_359 ();
 sg13g2_decap_8 FILLER_80_366 ();
 sg13g2_fill_2 FILLER_80_373 ();
 sg13g2_fill_1 FILLER_80_375 ();
 sg13g2_decap_8 FILLER_80_381 ();
 sg13g2_decap_8 FILLER_80_388 ();
 sg13g2_decap_8 FILLER_80_395 ();
 sg13g2_decap_8 FILLER_80_402 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
endmodule
