module tt_um_LnL_SoC (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \P0.clkout ;
 wire \P0.countreg[0] ;
 wire \P0.countreg[1] ;
 wire \P0.countreg[2] ;
 wire \P0.uptime[0] ;
 wire \P0.uptime[1] ;
 wire \P0.uptime[2] ;
 wire \P0.uptimelat[0] ;
 wire \P0.uptimelat[1] ;
 wire \P0.uptimelat[2] ;
 wire \P0.uptimereg[0] ;
 wire \P0.uptimereg[1] ;
 wire \P0.uptimereg[2] ;
 wire \T0.clkout ;
 wire \T0.count[0] ;
 wire \T0.count[1] ;
 wire \T0.count[2] ;
 wire \T0.count[3] ;
 wire \T0.count[4] ;
 wire \T0.count[5] ;
 wire \T0.count[6] ;
 wire \T0.count[7] ;
 wire \T0.selreg[0] ;
 wire \T0.selreg[1] ;
 wire \T0.selreg[2] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire \addr_to_memio[0] ;
 wire \addr_to_memio[10] ;
 wire \addr_to_memio[11] ;
 wire \addr_to_memio[1] ;
 wire \addr_to_memio[2] ;
 wire \addr_to_memio[3] ;
 wire \addr_to_memio[4] ;
 wire \addr_to_memio[5] ;
 wire \addr_to_memio[6] ;
 wire \addr_to_memio[7] ;
 wire \addr_to_memio[8] ;
 wire \addr_to_memio[9] ;
 wire \boot_to_cpu[0] ;
 wire \boot_to_cpu[10] ;
 wire \boot_to_cpu[11] ;
 wire \boot_to_cpu[12] ;
 wire \boot_to_cpu[13] ;
 wire \boot_to_cpu[14] ;
 wire \boot_to_cpu[15] ;
 wire \boot_to_cpu[1] ;
 wire \boot_to_cpu[2] ;
 wire \boot_to_cpu[3] ;
 wire \boot_to_cpu[4] ;
 wire \boot_to_cpu[5] ;
 wire \boot_to_cpu[6] ;
 wire \boot_to_cpu[7] ;
 wire \boot_to_cpu[8] ;
 wire \boot_to_cpu[9] ;
 wire \cpu0.ac0 ;
 wire \cpu0.ac15 ;
 wire \cpu0.ac[0] ;
 wire \cpu0.ac[10] ;
 wire \cpu0.ac[11] ;
 wire \cpu0.ac[12] ;
 wire \cpu0.ac[13] ;
 wire \cpu0.ac[14] ;
 wire \cpu0.ac[15] ;
 wire \cpu0.ac[1] ;
 wire \cpu0.ac[2] ;
 wire \cpu0.ac[3] ;
 wire \cpu0.ac[4] ;
 wire \cpu0.ac[5] ;
 wire \cpu0.ac[6] ;
 wire \cpu0.ac[7] ;
 wire \cpu0.ac[8] ;
 wire \cpu0.ac[9] ;
 wire \cpu0.clk ;
 wire \cpu0.dataout[3] ;
 wire \cpu0.dataout[4] ;
 wire \cpu0.dataout[5] ;
 wire \cpu0.dataout[6] ;
 wire \cpu0.dataout[7] ;
 wire \cpu0.decode2.a[0] ;
 wire \cpu0.decode2.a[1] ;
 wire \cpu0.decode2.a[2] ;
 wire \cpu0.dr[0] ;
 wire \cpu0.dr[10] ;
 wire \cpu0.dr[11] ;
 wire \cpu0.dr[12] ;
 wire \cpu0.dr[13] ;
 wire \cpu0.dr[14] ;
 wire \cpu0.dr[15] ;
 wire \cpu0.dr[1] ;
 wire \cpu0.dr[2] ;
 wire \cpu0.dr[3] ;
 wire \cpu0.dr[4] ;
 wire \cpu0.dr[5] ;
 wire \cpu0.dr[6] ;
 wire \cpu0.dr[7] ;
 wire \cpu0.dr[8] ;
 wire \cpu0.dr[9] ;
 wire \cpu0.e ;
 wire \cpu0.en_out ;
 wire \cpu0.ir[0] ;
 wire \cpu0.ir[10] ;
 wire \cpu0.ir[11] ;
 wire \cpu0.ir[15] ;
 wire \cpu0.ir[1] ;
 wire \cpu0.ir[2] ;
 wire \cpu0.ir[3] ;
 wire \cpu0.ir[4] ;
 wire \cpu0.ir[5] ;
 wire \cpu0.ir[6] ;
 wire \cpu0.ir[7] ;
 wire \cpu0.ir[8] ;
 wire \cpu0.ir[9] ;
 wire \cpu0.pc[0] ;
 wire \cpu0.pc[10] ;
 wire \cpu0.pc[11] ;
 wire \cpu0.pc[1] ;
 wire \cpu0.pc[2] ;
 wire \cpu0.pc[3] ;
 wire \cpu0.pc[4] ;
 wire \cpu0.pc[5] ;
 wire \cpu0.pc[6] ;
 wire \cpu0.pc[7] ;
 wire \cpu0.pc[8] ;
 wire \cpu0.pc[9] ;
 wire \cpu0.rstT ;
 wire \cpu0.t[0] ;
 wire \cpu0.t[10] ;
 wire \cpu0.t[1] ;
 wire \cpu0.t[2] ;
 wire \cpu0.t[3] ;
 wire \cpu0.t[4] ;
 wire \cpu0.t[5] ;
 wire \cpu0.t[6] ;
 wire \cpu0.t[7] ;
 wire \cpu0.t[8] ;
 wire \cpu0.t[9] ;
 wire \mem0.dout_internal[0] ;
 wire \mem0.dout_internal[10] ;
 wire \mem0.dout_internal[11] ;
 wire \mem0.dout_internal[12] ;
 wire \mem0.dout_internal[13] ;
 wire \mem0.dout_internal[14] ;
 wire \mem0.dout_internal[15] ;
 wire \mem0.dout_internal[1] ;
 wire \mem0.dout_internal[2] ;
 wire \mem0.dout_internal[3] ;
 wire \mem0.dout_internal[4] ;
 wire \mem0.dout_internal[5] ;
 wire \mem0.dout_internal[6] ;
 wire \mem0.dout_internal[7] ;
 wire \mem0.dout_internal[8] ;
 wire \mem0.dout_internal[9] ;
 wire rst_n_i;
 wire \spi0.cntreg[0] ;
 wire \spi0.cntreg[1] ;
 wire \spi0.cntreg[2] ;
 wire \spi0.cntreg[3] ;
 wire \spi0.dataout[0] ;
 wire \spi0.dataout[1] ;
 wire \spi0.dataout[2] ;
 wire \spi0.dataout[3] ;
 wire \spi0.dataout[4] ;
 wire \spi0.dataout[5] ;
 wire \spi0.dataout[6] ;
 wire \spi0.dataout[7] ;
 wire \spi0.datareg[0] ;
 wire \spi0.datareg[1] ;
 wire \spi0.datareg[2] ;
 wire \spi0.datareg[3] ;
 wire \spi0.datareg[4] ;
 wire \spi0.datareg[5] ;
 wire \spi0.datareg[6] ;
 wire \spi0.datareg[7] ;
 wire \spi0.sclk ;
 wire \spi0.ssn_out ;
 wire \spi0.unload ;
 wire net14;
 wire net15;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire clk_regs;
 wire net16;
 wire net17;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_3_0__leaf_clk_regs;
 wire clknet_3_1__leaf_clk_regs;
 wire clknet_3_2__leaf_clk_regs;
 wire clknet_3_3__leaf_clk_regs;
 wire clknet_3_4__leaf_clk_regs;
 wire clknet_3_5__leaf_clk_regs;
 wire clknet_3_6__leaf_clk_regs;
 wire clknet_3_7__leaf_clk_regs;
 wire \clknet_0_cpu0.clk ;
 wire \clknet_4_0_0_cpu0.clk ;
 wire \clknet_4_1_0_cpu0.clk ;
 wire \clknet_4_2_0_cpu0.clk ;
 wire \clknet_4_3_0_cpu0.clk ;
 wire \clknet_4_4_0_cpu0.clk ;
 wire \clknet_4_5_0_cpu0.clk ;
 wire \clknet_4_6_0_cpu0.clk ;
 wire \clknet_4_7_0_cpu0.clk ;
 wire \clknet_4_8_0_cpu0.clk ;
 wire \clknet_4_9_0_cpu0.clk ;
 wire \clknet_4_10_0_cpu0.clk ;
 wire \clknet_4_11_0_cpu0.clk ;
 wire \clknet_4_12_0_cpu0.clk ;
 wire \clknet_4_13_0_cpu0.clk ;
 wire \clknet_4_14_0_cpu0.clk ;
 wire \clknet_4_15_0_cpu0.clk ;
 wire delaynet_0_clk;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;

 sg13g2_inv_1 _0848_ (.Y(_0009_),
    .A(net39));
 sg13g2_inv_2 _0849_ (.Y(_0233_),
    .A(net160));
 sg13g2_inv_1 _0850_ (.Y(_0234_),
    .A(net152));
 sg13g2_inv_2 _0851_ (.Y(_0235_),
    .A(net298));
 sg13g2_inv_2 _0852_ (.Y(_0236_),
    .A(net137));
 sg13g2_inv_1 _0853_ (.Y(_0237_),
    .A(net78));
 sg13g2_inv_2 _0854_ (.Y(_0238_),
    .A(net217));
 sg13g2_inv_1 _0855_ (.Y(_0239_),
    .A(net317));
 sg13g2_inv_1 _0856_ (.Y(_0240_),
    .A(net153));
 sg13g2_inv_1 _0857_ (.Y(_0241_),
    .A(net316));
 sg13g2_inv_1 _0858_ (.Y(_0242_),
    .A(net146));
 sg13g2_inv_1 _0859_ (.Y(_0243_),
    .A(net315));
 sg13g2_inv_2 _0860_ (.Y(_0244_),
    .A(net150));
 sg13g2_inv_2 _0861_ (.Y(_0245_),
    .A(net179));
 sg13g2_inv_1 _0862_ (.Y(_0246_),
    .A(net92));
 sg13g2_inv_1 _0863_ (.Y(_0247_),
    .A(net344));
 sg13g2_inv_2 _0864_ (.Y(_0248_),
    .A(net97));
 sg13g2_inv_1 _0865_ (.Y(_0249_),
    .A(net299));
 sg13g2_inv_2 _0866_ (.Y(_0250_),
    .A(net135));
 sg13g2_inv_1 _0867_ (.Y(_0251_),
    .A(net87));
 sg13g2_inv_1 _0868_ (.Y(_0252_),
    .A(net333));
 sg13g2_inv_1 _0869_ (.Y(_0253_),
    .A(net331));
 sg13g2_inv_1 _0870_ (.Y(_0254_),
    .A(net332));
 sg13g2_inv_1 _0871_ (.Y(_0255_),
    .A(net327));
 sg13g2_inv_1 _0872_ (.Y(_0256_),
    .A(net329));
 sg13g2_inv_2 _0873_ (.Y(_0257_),
    .A(net325));
 sg13g2_inv_1 _0874_ (.Y(_0258_),
    .A(net326));
 sg13g2_inv_2 _0875_ (.Y(_0259_),
    .A(net166));
 sg13g2_inv_2 _0876_ (.Y(_0260_),
    .A(net181));
 sg13g2_inv_1 _0877_ (.Y(_0261_),
    .A(net350));
 sg13g2_inv_1 _0878_ (.Y(_0262_),
    .A(net351));
 sg13g2_inv_2 _0879_ (.Y(_0263_),
    .A(net162));
 sg13g2_inv_1 _0880_ (.Y(_0264_),
    .A(net349));
 sg13g2_inv_2 _0881_ (.Y(_0265_),
    .A(net184));
 sg13g2_inv_1 _0882_ (.Y(_0266_),
    .A(net182));
 sg13g2_inv_1 _0883_ (.Y(_0267_),
    .A(net118));
 sg13g2_inv_1 _0884_ (.Y(_0268_),
    .A(net86));
 sg13g2_inv_2 _0885_ (.Y(_0269_),
    .A(net69));
 sg13g2_inv_4 _0886_ (.A(net313),
    .Y(_0270_));
 sg13g2_inv_1 _0887_ (.Y(_0271_),
    .A(net107));
 sg13g2_inv_1 _0888_ (.Y(_0272_),
    .A(net77));
 sg13g2_inv_1 _0889_ (.Y(_0273_),
    .A(net104));
 sg13g2_inv_1 _0890_ (.Y(_0274_),
    .A(net121));
 sg13g2_inv_1 _0891_ (.Y(_0275_),
    .A(net123));
 sg13g2_inv_1 _0892_ (.Y(_0276_),
    .A(\cpu0.pc[0] ));
 sg13g2_inv_4 _0893_ (.A(net158),
    .Y(_0277_));
 sg13g2_inv_2 _0894_ (.Y(_0278_),
    .A(net155));
 sg13g2_inv_1 _0895_ (.Y(_0279_),
    .A(net164));
 sg13g2_inv_2 _0896_ (.Y(_0280_),
    .A(\addr_to_memio[3] ));
 sg13g2_inv_2 _0897_ (.Y(_0281_),
    .A(net126));
 sg13g2_inv_1 _0898_ (.Y(_0282_),
    .A(\cpu0.pc[5] ));
 sg13g2_inv_1 _0899_ (.Y(_0283_),
    .A(net98));
 sg13g2_inv_1 _0900_ (.Y(_0284_),
    .A(net131));
 sg13g2_inv_1 _0901_ (.Y(_0285_),
    .A(net90));
 sg13g2_inv_1 _0902_ (.Y(_0286_),
    .A(\T0.count[3] ));
 sg13g2_inv_1 _0903_ (.Y(_0012_),
    .A(net42));
 sg13g2_nand2_1 _0904_ (.Y(_0287_),
    .A(\cpu0.decode2.a[0] ),
    .B(\cpu0.decode2.a[1] ));
 sg13g2_nor2_2 _0905_ (.A(net298),
    .B(_0287_),
    .Y(_0288_));
 sg13g2_and2_1 _0906_ (.A(\cpu0.t[6] ),
    .B(net297),
    .X(_0289_));
 sg13g2_a21oi_2 _0907_ (.B1(net293),
    .Y(_0290_),
    .A2(net338),
    .A1(net296));
 sg13g2_nand2b_2 _0908_ (.Y(_0816_),
    .B(net291),
    .A_N(_0290_));
 sg13g2_nand2_1 _0909_ (.Y(_0291_),
    .A(_0234_),
    .B(\cpu0.decode2.a[2] ));
 sg13g2_nor2b_2 _0910_ (.A(\cpu0.decode2.a[0] ),
    .B_N(\cpu0.decode2.a[1] ),
    .Y(_0292_));
 sg13g2_and2_1 _0911_ (.A(net298),
    .B(_0292_),
    .X(_0293_));
 sg13g2_nand2_2 _0912_ (.Y(_0294_),
    .A(net298),
    .B(_0292_));
 sg13g2_nor2b_2 _0913_ (.A(net297),
    .B_N(\cpu0.t[7] ),
    .Y(_0295_));
 sg13g2_o21ai_1 _0914_ (.B1(net290),
    .Y(_0808_),
    .A1(net293),
    .A2(net292));
 sg13g2_nand2_2 _0915_ (.Y(_0296_),
    .A(\cpu0.decode2.a[0] ),
    .B(_0236_));
 sg13g2_nor2_2 _0916_ (.A(_0235_),
    .B(_0296_),
    .Y(_0297_));
 sg13g2_inv_1 _0917_ (.Y(_0298_),
    .A(net285));
 sg13g2_nand2_2 _0918_ (.Y(_0825_),
    .A(net337),
    .B(_0297_));
 sg13g2_and3_1 _0919_ (.X(_0299_),
    .A(\cpu0.decode2.a[0] ),
    .B(\cpu0.decode2.a[2] ),
    .C(\cpu0.decode2.a[1] ));
 sg13g2_nand3_1 _0920_ (.B(\cpu0.decode2.a[2] ),
    .C(\cpu0.decode2.a[1] ),
    .A(\cpu0.decode2.a[0] ),
    .Y(_0300_));
 sg13g2_nor2_2 _0921_ (.A(net296),
    .B(net294),
    .Y(_0301_));
 sg13g2_nand2_1 _0922_ (.Y(_0302_),
    .A(net342),
    .B(_0299_));
 sg13g2_nor2_1 _0923_ (.A(net296),
    .B(_0302_),
    .Y(_0303_));
 sg13g2_and2_1 _0924_ (.A(\cpu0.ir[10] ),
    .B(_0303_),
    .X(\cpu0.en_out ));
 sg13g2_nor3_1 _0925_ (.A(\P0.uptimereg[1] ),
    .B(\P0.uptimereg[0] ),
    .C(\P0.uptimereg[2] ),
    .Y(_0304_));
 sg13g2_inv_1 _0926_ (.Y(\P0.clkout ),
    .A(_0304_));
 sg13g2_nor2_1 _0927_ (.A(\spi0.cntreg[1] ),
    .B(net112),
    .Y(_0305_));
 sg13g2_nor4_1 _0928_ (.A(net59),
    .B(\spi0.cntreg[2] ),
    .C(net116),
    .D(net112),
    .Y(\spi0.ssn_out ));
 sg13g2_nand2_1 _0929_ (.Y(_0306_),
    .A(net297),
    .B(net54));
 sg13g2_o21ai_1 _0930_ (.B1(_0816_),
    .Y(_0307_),
    .A1(_0294_),
    .A2(_0306_));
 sg13g2_o21ai_1 _0931_ (.B1(net290),
    .Y(_0308_),
    .A1(\cpu0.t[6] ),
    .A2(\cpu0.t[7] ));
 sg13g2_a21oi_1 _0932_ (.A1(_0825_),
    .A2(_0308_),
    .Y(_0309_),
    .B1(net297));
 sg13g2_or2_1 _0933_ (.X(_0310_),
    .B(_0309_),
    .A(_0307_));
 sg13g2_inv_1 _0934_ (.Y(_0311_),
    .A(_0310_));
 sg13g2_or2_1 _0935_ (.X(_0312_),
    .B(\addr_to_memio[7] ),
    .A(\addr_to_memio[8] ));
 sg13g2_nor4_2 _0936_ (.A(\addr_to_memio[10] ),
    .B(\addr_to_memio[9] ),
    .C(\addr_to_memio[11] ),
    .Y(_0313_),
    .D(_0312_));
 sg13g2_a21oi_1 _0937_ (.A1(net297),
    .A2(_0236_),
    .Y(_0314_),
    .B1(_0292_));
 sg13g2_nand3_1 _0938_ (.B(_0296_),
    .C(_0314_),
    .A(net298),
    .Y(_0315_));
 sg13g2_nand2b_1 _0939_ (.Y(_0316_),
    .B(_0308_),
    .A_N(\cpu0.t[1] ));
 sg13g2_a221oi_1 _0940_ (.B2(net338),
    .C1(_0316_),
    .B1(_0315_),
    .A1(net293),
    .Y(_0317_),
    .A2(_0300_));
 sg13g2_nor2_2 _0941_ (.A(_0313_),
    .B(_0317_),
    .Y(_0318_));
 sg13g2_or2_1 _0942_ (.X(_0319_),
    .B(_0317_),
    .A(_0313_));
 sg13g2_nand2_2 _0943_ (.Y(_0320_),
    .A(_0310_),
    .B(net276));
 sg13g2_nor2b_1 _0944_ (.A(net12),
    .B_N(net11),
    .Y(_0321_));
 sg13g2_mux2_1 _0945_ (.A0(\P0.uptime[0] ),
    .A1(_0321_),
    .S(net267),
    .X(_0001_));
 sg13g2_mux2_1 _0946_ (.A0(\P0.uptime[1] ),
    .A1(net106),
    .S(net267),
    .X(_0002_));
 sg13g2_mux2_1 _0947_ (.A0(\P0.uptime[2] ),
    .A1(net80),
    .S(net267),
    .X(_0003_));
 sg13g2_mux2_1 _0948_ (.A0(\cpu0.dataout[3] ),
    .A1(net96),
    .S(net267),
    .X(_0004_));
 sg13g2_mux2_1 _0949_ (.A0(\cpu0.dataout[4] ),
    .A1(net79),
    .S(net267),
    .X(_0005_));
 sg13g2_mux2_1 _0950_ (.A0(\cpu0.dataout[5] ),
    .A1(net100),
    .S(net267),
    .X(_0006_));
 sg13g2_mux2_1 _0951_ (.A0(\cpu0.dataout[6] ),
    .A1(net83),
    .S(net267),
    .X(_0007_));
 sg13g2_mux2_1 _0952_ (.A0(\cpu0.dataout[7] ),
    .A1(net91),
    .S(_0320_),
    .X(_0008_));
 sg13g2_nor2_2 _0953_ (.A(\addr_to_memio[2] ),
    .B(\addr_to_memio[3] ),
    .Y(_0322_));
 sg13g2_and2_1 _0954_ (.A(net323),
    .B(net322),
    .X(_0323_));
 sg13g2_nand2_1 _0955_ (.Y(_0324_),
    .A(net323),
    .B(net322));
 sg13g2_nor2_1 _0956_ (.A(net320),
    .B(_0324_),
    .Y(_0325_));
 sg13g2_and2_1 _0957_ (.A(_0322_),
    .B(_0325_),
    .X(_0326_));
 sg13g2_nor2_1 _0958_ (.A(net323),
    .B(net322),
    .Y(_0327_));
 sg13g2_nor2_2 _0959_ (.A(net323),
    .B(net321),
    .Y(_0328_));
 sg13g2_nor3_1 _0960_ (.A(net323),
    .B(net322),
    .C(net321),
    .Y(_0329_));
 sg13g2_nor2b_2 _0961_ (.A(net322),
    .B_N(net323),
    .Y(_0330_));
 sg13g2_and2_1 _0962_ (.A(net321),
    .B(_0322_),
    .X(_0331_));
 sg13g2_a221oi_1 _0963_ (.B2(_0331_),
    .C1(_0326_),
    .B1(_0330_),
    .A1(\addr_to_memio[3] ),
    .Y(_0332_),
    .A2(_0329_));
 sg13g2_nor2_2 _0964_ (.A(_0278_),
    .B(_0280_),
    .Y(_0333_));
 sg13g2_nand2_1 _0965_ (.Y(_0334_),
    .A(_0328_),
    .B(_0333_));
 sg13g2_nor2_1 _0966_ (.A(net324),
    .B(_0277_),
    .Y(_0335_));
 sg13g2_nand2b_1 _0967_ (.Y(_0336_),
    .B(net322),
    .A_N(net323));
 sg13g2_nor2_2 _0968_ (.A(\addr_to_memio[2] ),
    .B(_0280_),
    .Y(_0337_));
 sg13g2_nand2_1 _0969_ (.Y(_0338_),
    .A(_0330_),
    .B(_0337_));
 sg13g2_a22oi_1 _0970_ (.Y(_0339_),
    .B1(_0337_),
    .B2(_0330_),
    .A2(_0335_),
    .A1(_0333_));
 sg13g2_or2_1 _0971_ (.X(_0340_),
    .B(_0339_),
    .A(net320));
 sg13g2_and2_1 _0972_ (.A(_0332_),
    .B(_0340_),
    .X(_0341_));
 sg13g2_nand2_1 _0973_ (.Y(_0342_),
    .A(net320),
    .B(_0333_));
 sg13g2_inv_1 _0974_ (.Y(_0343_),
    .A(_0342_));
 sg13g2_nor2_1 _0975_ (.A(net322),
    .B(_0342_),
    .Y(_0344_));
 sg13g2_nand2_1 _0976_ (.Y(_0345_),
    .A(_0330_),
    .B(_0333_));
 sg13g2_nor2_1 _0977_ (.A(_0278_),
    .B(\addr_to_memio[3] ),
    .Y(_0346_));
 sg13g2_nor3_2 _0978_ (.A(_0277_),
    .B(_0278_),
    .C(\addr_to_memio[3] ),
    .Y(_0347_));
 sg13g2_a22oi_1 _0979_ (.Y(_0348_),
    .B1(_0347_),
    .B2(net324),
    .A2(_0333_),
    .A1(_0330_));
 sg13g2_or2_1 _0980_ (.X(_0349_),
    .B(_0348_),
    .A(net320));
 sg13g2_nand3b_1 _0981_ (.B(_0349_),
    .C(_0341_),
    .Y(\mem0.dout_internal[0] ),
    .A_N(_0344_));
 sg13g2_nand2_1 _0982_ (.Y(_0350_),
    .A(net320),
    .B(_0337_));
 sg13g2_nor2_1 _0983_ (.A(_0324_),
    .B(_0350_),
    .Y(_0351_));
 sg13g2_nand3_1 _0984_ (.B(net321),
    .C(_0323_),
    .A(\addr_to_memio[3] ),
    .Y(_0352_));
 sg13g2_nand2_1 _0985_ (.Y(\mem0.dout_internal[1] ),
    .A(_0341_),
    .B(_0352_));
 sg13g2_a21oi_1 _0986_ (.A1(net322),
    .A2(_0343_),
    .Y(_0353_),
    .B1(_0351_));
 sg13g2_nor2_1 _0987_ (.A(net320),
    .B(_0336_),
    .Y(_0354_));
 sg13g2_nand2_1 _0988_ (.Y(_0355_),
    .A(_0337_),
    .B(_0354_));
 sg13g2_nand3_1 _0989_ (.B(_0353_),
    .C(_0355_),
    .A(_0332_),
    .Y(\mem0.dout_internal[2] ));
 sg13g2_nand2b_1 _0990_ (.Y(_0356_),
    .B(_0331_),
    .A_N(net323));
 sg13g2_nand2b_1 _0991_ (.Y(_0357_),
    .B(_0277_),
    .A_N(_0356_));
 sg13g2_nand3_1 _0992_ (.B(_0353_),
    .C(_0357_),
    .A(_0340_),
    .Y(\mem0.dout_internal[3] ));
 sg13g2_nand2_1 _0993_ (.Y(_0358_),
    .A(_0330_),
    .B(_0346_));
 sg13g2_nor2_1 _0994_ (.A(net320),
    .B(_0358_),
    .Y(_0359_));
 sg13g2_inv_1 _0995_ (.Y(_0360_),
    .A(_0359_));
 sg13g2_a21oi_1 _0996_ (.A1(_0328_),
    .A2(_0347_),
    .Y(_0361_),
    .B1(_0359_));
 sg13g2_nand3_1 _0997_ (.B(_0353_),
    .C(_0361_),
    .A(_0349_),
    .Y(\mem0.dout_internal[4] ));
 sg13g2_nand2_1 _0998_ (.Y(_0362_),
    .A(net320),
    .B(_0347_));
 sg13g2_nand2_1 _0999_ (.Y(_0363_),
    .A(_0325_),
    .B(_0337_));
 sg13g2_nand2_1 _1000_ (.Y(\mem0.dout_internal[5] ),
    .A(_0362_),
    .B(_0363_));
 sg13g2_a21o_1 _1001_ (.A2(_0358_),
    .A1(_0338_),
    .B1(_0281_),
    .X(_0364_));
 sg13g2_o21ai_1 _1002_ (.B1(_0364_),
    .Y(\mem0.dout_internal[6] ),
    .A1(_0336_),
    .A2(_0350_));
 sg13g2_nand2_1 _1003_ (.Y(_0365_),
    .A(_0327_),
    .B(_0343_));
 sg13g2_nand2_1 _1004_ (.Y(_0366_),
    .A(_0331_),
    .B(_0335_));
 sg13g2_nand4_1 _1005_ (.B(_0363_),
    .C(_0365_),
    .A(_0360_),
    .Y(\mem0.dout_internal[7] ),
    .D(_0366_));
 sg13g2_nand3_1 _1006_ (.B(_0327_),
    .C(_0337_),
    .A(net321),
    .Y(_0367_));
 sg13g2_inv_1 _1007_ (.Y(\mem0.dout_internal[8] ),
    .A(_0367_));
 sg13g2_nand2_1 _1008_ (.Y(_0368_),
    .A(_0325_),
    .B(_0333_));
 sg13g2_nand2_2 _1009_ (.Y(_0369_),
    .A(_0322_),
    .B(_0328_));
 sg13g2_o21ai_1 _1010_ (.B1(_0368_),
    .Y(\mem0.dout_internal[9] ),
    .A1(\addr_to_memio[1] ),
    .A2(_0369_));
 sg13g2_nand2_1 _1011_ (.Y(_0370_),
    .A(_0327_),
    .B(_0346_));
 sg13g2_nand2_1 _1012_ (.Y(_0371_),
    .A(_0323_),
    .B(_0331_));
 sg13g2_nand2_1 _1013_ (.Y(\mem0.dout_internal[10] ),
    .A(_0370_),
    .B(_0371_));
 sg13g2_nor2_1 _1014_ (.A(_0277_),
    .B(_0369_),
    .Y(\mem0.dout_internal[11] ));
 sg13g2_nand4_1 _1015_ (.B(_0368_),
    .C(_0370_),
    .A(_0356_),
    .Y(_0372_),
    .D(_0371_));
 sg13g2_nand3_1 _1016_ (.B(_0362_),
    .C(_0367_),
    .A(_0355_),
    .Y(_0373_));
 sg13g2_nor3_1 _1017_ (.A(\mem0.dout_internal[6] ),
    .B(_0372_),
    .C(_0373_),
    .Y(_0374_));
 sg13g2_and2_1 _1018_ (.A(_0361_),
    .B(_0369_),
    .X(_0375_));
 sg13g2_o21ai_1 _1019_ (.B1(_0345_),
    .Y(_0376_),
    .A1(_0277_),
    .A2(_0334_));
 sg13g2_nor3_1 _1020_ (.A(_0326_),
    .B(_0351_),
    .C(_0376_),
    .Y(_0377_));
 sg13g2_nand3_1 _1021_ (.B(_0375_),
    .C(_0377_),
    .A(_0374_),
    .Y(\mem0.dout_internal[12] ));
 sg13g2_a221oi_1 _1022_ (.B2(_0329_),
    .C1(_0344_),
    .B1(_0337_),
    .A1(_0328_),
    .Y(_0378_),
    .A2(_0333_));
 sg13g2_nand3_1 _1023_ (.B(_0375_),
    .C(_0378_),
    .A(_0374_),
    .Y(\mem0.dout_internal[13] ));
 sg13g2_nand3_1 _1024_ (.B(net321),
    .C(_0347_),
    .A(net324),
    .Y(_0379_));
 sg13g2_nand3_1 _1025_ (.B(_0322_),
    .C(_0330_),
    .A(_0281_),
    .Y(_0380_));
 sg13g2_nand3_1 _1026_ (.B(_0379_),
    .C(_0380_),
    .A(_0367_),
    .Y(_0381_));
 sg13g2_o21ai_1 _1027_ (.B1(_0354_),
    .Y(_0382_),
    .A1(_0337_),
    .A2(_0346_));
 sg13g2_nand4_1 _1028_ (.B(_0364_),
    .C(_0369_),
    .A(_0352_),
    .Y(_0383_),
    .D(_0382_));
 sg13g2_or4_1 _1029_ (.A(_0344_),
    .B(_0372_),
    .C(_0381_),
    .D(_0383_),
    .X(\mem0.dout_internal[14] ));
 sg13g2_nand2_1 _1030_ (.Y(_0384_),
    .A(_0345_),
    .B(_0370_));
 sg13g2_a22oi_1 _1031_ (.Y(_0385_),
    .B1(_0384_),
    .B2(_0281_),
    .A2(_0343_),
    .A1(_0323_));
 sg13g2_nand4_1 _1032_ (.B(_0369_),
    .C(_0371_),
    .A(_0334_),
    .Y(\mem0.dout_internal[15] ),
    .D(_0385_));
 sg13g2_mux2_1 _1033_ (.A0(\T0.count[4] ),
    .A1(\T0.count[5] ),
    .S(\T0.selreg[0] ),
    .X(_0386_));
 sg13g2_nor2b_1 _1034_ (.A(\T0.selreg[0] ),
    .B_N(\T0.count[6] ),
    .Y(_0387_));
 sg13g2_a21oi_1 _1035_ (.A1(\T0.selreg[0] ),
    .A2(\T0.count[7] ),
    .Y(_0388_),
    .B1(_0387_));
 sg13g2_o21ai_1 _1036_ (.B1(\T0.selreg[2] ),
    .Y(_0389_),
    .A1(\T0.selreg[1] ),
    .A2(_0386_));
 sg13g2_a21oi_1 _1037_ (.A1(\T0.selreg[1] ),
    .A2(_0388_),
    .Y(_0390_),
    .B1(_0389_));
 sg13g2_a21oi_1 _1038_ (.A1(\T0.selreg[0] ),
    .A2(\T0.count[1] ),
    .Y(_0391_),
    .B1(\T0.selreg[1] ));
 sg13g2_o21ai_1 _1039_ (.B1(_0391_),
    .Y(_0392_),
    .A1(\T0.selreg[0] ),
    .A2(_0012_));
 sg13g2_nor2b_1 _1040_ (.A(\T0.selreg[0] ),
    .B_N(\T0.count[2] ),
    .Y(_0393_));
 sg13g2_a21oi_1 _1041_ (.A1(\T0.selreg[0] ),
    .A2(\T0.count[3] ),
    .Y(_0394_),
    .B1(_0393_));
 sg13g2_a21oi_1 _1042_ (.A1(\T0.selreg[1] ),
    .A2(_0394_),
    .Y(_0395_),
    .B1(\T0.selreg[2] ));
 sg13g2_a21o_1 _1043_ (.A2(_0395_),
    .A1(_0392_),
    .B1(_0390_),
    .X(\T0.clkout ));
 sg13g2_nor2_2 _1044_ (.A(net311),
    .B(net306),
    .Y(_0396_));
 sg13g2_nor2_1 _1045_ (.A(_0300_),
    .B(_0396_),
    .Y(_0397_));
 sg13g2_a21o_1 _1046_ (.A2(net291),
    .A1(net296),
    .B1(_0397_),
    .X(_0398_));
 sg13g2_nor2_1 _1047_ (.A(\cpu0.decode2.a[1] ),
    .B(_0291_),
    .Y(_0399_));
 sg13g2_or2_1 _1048_ (.X(_0400_),
    .B(_0399_),
    .A(net291));
 sg13g2_nand2_1 _1049_ (.Y(_0401_),
    .A(net187),
    .B(net290));
 sg13g2_nand3_1 _1050_ (.B(_0299_),
    .C(_0396_),
    .A(net338),
    .Y(_0402_));
 sg13g2_a21o_1 _1051_ (.A2(\cpu0.t[9] ),
    .A1(_0235_),
    .B1(net292),
    .X(_0403_));
 sg13g2_nand3_1 _1052_ (.B(_0291_),
    .C(_0403_),
    .A(_0287_),
    .Y(_0404_));
 sg13g2_nand4_1 _1053_ (.B(_0401_),
    .C(_0402_),
    .A(net363),
    .Y(_0405_),
    .D(_0404_));
 sg13g2_a221oi_1 _1054_ (.B2(net72),
    .C1(_0405_),
    .B1(_0400_),
    .A1(net78),
    .Y(_0406_),
    .A2(_0398_));
 sg13g2_inv_1 _1055_ (.Y(\cpu0.rstT ),
    .A(net278));
 sg13g2_nor2_2 _1056_ (.A(\cpu0.ir[15] ),
    .B(_0302_),
    .Y(_0407_));
 sg13g2_a21o_1 _1057_ (.A2(_0407_),
    .A1(\cpu0.ir[0] ),
    .B1(clknet_1_0__leaf_clk),
    .X(\cpu0.clk ));
 sg13g2_nand2_1 _1058_ (.Y(_0408_),
    .A(_0283_),
    .B(_0313_));
 sg13g2_nor4_1 _1059_ (.A(\addr_to_memio[6] ),
    .B(_0310_),
    .C(_0317_),
    .D(_0408_),
    .Y(_0000_));
 sg13g2_nor2b_1 _1060_ (.A(\spi0.ssn_out ),
    .B_N(clknet_1_1__leaf_clk),
    .Y(\spi0.sclk ));
 sg13g2_nand2_1 _1061_ (.Y(_0409_),
    .A(net39),
    .B(net43));
 sg13g2_xor2_1 _1062_ (.B(net43),
    .A(net39),
    .X(_0010_));
 sg13g2_xnor2_1 _1063_ (.Y(_0011_),
    .A(net56),
    .B(_0409_));
 sg13g2_xor2_1 _1064_ (.B(net42),
    .A(net44),
    .X(_0013_));
 sg13g2_nand3_1 _1065_ (.B(net44),
    .C(net42),
    .A(net172),
    .Y(_0410_));
 sg13g2_a21o_1 _1066_ (.A2(net42),
    .A1(net44),
    .B1(net172),
    .X(_0411_));
 sg13g2_and2_1 _1067_ (.A(_0410_),
    .B(_0411_),
    .X(_0014_));
 sg13g2_nor2_1 _1068_ (.A(_0286_),
    .B(_0410_),
    .Y(_0412_));
 sg13g2_xnor2_1 _1069_ (.Y(_0015_),
    .A(net67),
    .B(_0410_));
 sg13g2_and2_1 _1070_ (.A(net52),
    .B(_0412_),
    .X(_0413_));
 sg13g2_xor2_1 _1071_ (.B(_0412_),
    .A(net52),
    .X(_0016_));
 sg13g2_xor2_1 _1072_ (.B(_0413_),
    .A(net57),
    .X(_0017_));
 sg13g2_nand3_1 _1073_ (.B(net57),
    .C(_0413_),
    .A(net177),
    .Y(_0414_));
 sg13g2_a21o_1 _1074_ (.A2(_0413_),
    .A1(net57),
    .B1(net177),
    .X(_0415_));
 sg13g2_and2_1 _1075_ (.A(_0414_),
    .B(_0415_),
    .X(_0018_));
 sg13g2_xnor2_1 _1076_ (.Y(_0019_),
    .A(net45),
    .B(_0414_));
 sg13g2_nor2_2 _1077_ (.A(_0310_),
    .B(net275),
    .Y(\spi0.unload ));
 sg13g2_nor2_2 _1078_ (.A(net338),
    .B(net342),
    .Y(_0416_));
 sg13g2_inv_1 _1079_ (.Y(_0417_),
    .A(_0416_));
 sg13g2_nand2_1 _1080_ (.Y(_0418_),
    .A(net88),
    .B(net296));
 sg13g2_a21oi_1 _1081_ (.A1(\cpu0.t[6] ),
    .A2(_0233_),
    .Y(_0419_),
    .B1(net54));
 sg13g2_nand2b_1 _1082_ (.Y(_0420_),
    .B(_0416_),
    .A_N(_0419_));
 sg13g2_a21oi_1 _1083_ (.A1(\cpu0.decode2.a[0] ),
    .A2(\cpu0.decode2.a[1] ),
    .Y(_0421_),
    .B1(net298));
 sg13g2_nor2_2 _1084_ (.A(net294),
    .B(net77),
    .Y(_0422_));
 sg13g2_nand2_2 _1085_ (.Y(_0423_),
    .A(net342),
    .B(_0272_));
 sg13g2_nand2_2 _1086_ (.Y(_0424_),
    .A(net296),
    .B(_0422_));
 sg13g2_nor4_1 _1087_ (.A(net299),
    .B(net311),
    .C(\cpu0.ir[5] ),
    .D(net310),
    .Y(_0425_));
 sg13g2_nor2_1 _1088_ (.A(_0300_),
    .B(_0424_),
    .Y(_0426_));
 sg13g2_a22oi_1 _1089_ (.Y(_0427_),
    .B1(_0425_),
    .B2(_0426_),
    .A2(_0420_),
    .A1(_0302_));
 sg13g2_o21ai_1 _1090_ (.B1(_0427_),
    .Y(_0428_),
    .A1(_0417_),
    .A2(_0421_));
 sg13g2_or2_1 _1091_ (.X(_0429_),
    .B(_0428_),
    .A(_0303_));
 sg13g2_and2_1 _1092_ (.A(net318),
    .B(net333),
    .X(_0430_));
 sg13g2_nand2_1 _1093_ (.Y(_0431_),
    .A(net318),
    .B(net333));
 sg13g2_and2_1 _1094_ (.A(net319),
    .B(net336),
    .X(_0432_));
 sg13g2_or2_1 _1095_ (.X(_0433_),
    .B(net333),
    .A(net318));
 sg13g2_nand3_1 _1096_ (.B(_0432_),
    .C(_0433_),
    .A(_0431_),
    .Y(_0434_));
 sg13g2_a21oi_1 _1097_ (.A1(_0432_),
    .A2(_0433_),
    .Y(_0435_),
    .B1(_0430_));
 sg13g2_nand2_1 _1098_ (.Y(_0436_),
    .A(\cpu0.dr[2] ),
    .B(net332));
 sg13g2_xnor2_1 _1099_ (.Y(_0437_),
    .A(\cpu0.dr[2] ),
    .B(net332));
 sg13g2_or2_1 _1100_ (.X(_0438_),
    .B(_0437_),
    .A(_0435_));
 sg13g2_nand2_1 _1101_ (.Y(_0439_),
    .A(\cpu0.dr[3] ),
    .B(net331));
 sg13g2_and2_1 _1102_ (.A(_0436_),
    .B(_0439_),
    .X(_0440_));
 sg13g2_o21ai_1 _1103_ (.B1(_0440_),
    .Y(_0441_),
    .A1(_0435_),
    .A2(_0437_));
 sg13g2_nand2_1 _1104_ (.Y(_0442_),
    .A(_0238_),
    .B(_0253_));
 sg13g2_and2_1 _1105_ (.A(_0441_),
    .B(_0442_),
    .X(_0443_));
 sg13g2_nand2_1 _1106_ (.Y(_0444_),
    .A(net316),
    .B(net325));
 sg13g2_xnor2_1 _1107_ (.Y(_0445_),
    .A(net316),
    .B(net325));
 sg13g2_and2_1 _1108_ (.A(\cpu0.dr[6] ),
    .B(net326),
    .X(_0446_));
 sg13g2_or2_1 _1109_ (.X(_0447_),
    .B(net326),
    .A(\cpu0.dr[6] ));
 sg13g2_xnor2_1 _1110_ (.Y(_0448_),
    .A(\cpu0.dr[6] ),
    .B(net326));
 sg13g2_or2_1 _1111_ (.X(_0449_),
    .B(_0448_),
    .A(_0445_));
 sg13g2_nand2_1 _1112_ (.Y(_0450_),
    .A(net317),
    .B(net327));
 sg13g2_nor2_1 _1113_ (.A(net317),
    .B(net327),
    .Y(_0451_));
 sg13g2_xnor2_1 _1114_ (.Y(_0452_),
    .A(net317),
    .B(net327));
 sg13g2_and2_1 _1115_ (.A(\cpu0.dr[4] ),
    .B(net329),
    .X(_0453_));
 sg13g2_nor2_1 _1116_ (.A(\cpu0.dr[4] ),
    .B(net329),
    .Y(_0454_));
 sg13g2_nor2_1 _1117_ (.A(_0453_),
    .B(_0454_),
    .Y(_0455_));
 sg13g2_nor4_1 _1118_ (.A(_0449_),
    .B(_0452_),
    .C(_0453_),
    .D(_0454_),
    .Y(_0456_));
 sg13g2_and3_1 _1119_ (.X(_0457_),
    .A(_0441_),
    .B(_0442_),
    .C(_0456_));
 sg13g2_nand3_1 _1120_ (.B(_0442_),
    .C(_0456_),
    .A(_0441_),
    .Y(_0458_));
 sg13g2_o21ai_1 _1121_ (.B1(_0446_),
    .Y(_0459_),
    .A1(\cpu0.dr[7] ),
    .A2(net325));
 sg13g2_nand2_1 _1122_ (.Y(_0460_),
    .A(_0444_),
    .B(_0459_));
 sg13g2_a21oi_1 _1123_ (.A1(net317),
    .A2(net327),
    .Y(_0461_),
    .B1(_0453_));
 sg13g2_nor3_1 _1124_ (.A(_0449_),
    .B(_0451_),
    .C(_0461_),
    .Y(_0462_));
 sg13g2_nor2_1 _1125_ (.A(_0460_),
    .B(_0462_),
    .Y(_0463_));
 sg13g2_or2_1 _1126_ (.X(_0464_),
    .B(_0462_),
    .A(_0460_));
 sg13g2_nand2_1 _1127_ (.Y(_0465_),
    .A(net315),
    .B(\cpu0.ac[8] ));
 sg13g2_xor2_1 _1128_ (.B(\cpu0.ac[8] ),
    .A(net315),
    .X(_0466_));
 sg13g2_inv_1 _1129_ (.Y(_0467_),
    .A(_0466_));
 sg13g2_nand3_1 _1130_ (.B(_0463_),
    .C(_0467_),
    .A(_0458_),
    .Y(_0468_));
 sg13g2_a21oi_1 _1131_ (.A1(_0458_),
    .A2(_0463_),
    .Y(_0469_),
    .B1(_0467_));
 sg13g2_nor2_2 _1132_ (.A(net298),
    .B(_0296_),
    .Y(_0470_));
 sg13g2_nand2b_2 _1133_ (.Y(_0471_),
    .B(_0235_),
    .A_N(_0296_));
 sg13g2_nor2_1 _1134_ (.A(_0469_),
    .B(net281),
    .Y(_0472_));
 sg13g2_and2_1 _1135_ (.A(_0235_),
    .B(_0292_),
    .X(_0473_));
 sg13g2_nand2_2 _1136_ (.Y(_0474_),
    .A(_0235_),
    .B(_0292_));
 sg13g2_nor2_1 _1137_ (.A(_0465_),
    .B(net284),
    .Y(_0475_));
 sg13g2_a21oi_1 _1138_ (.A1(_0468_),
    .A2(_0472_),
    .Y(_0476_),
    .B1(_0475_));
 sg13g2_o21ai_1 _1139_ (.B1(net294),
    .Y(_0477_),
    .A1(net315),
    .A2(_0474_));
 sg13g2_a21oi_1 _1140_ (.A1(_0474_),
    .A2(_0476_),
    .Y(_0478_),
    .B1(_0477_));
 sg13g2_nand2_1 _1141_ (.Y(_0479_),
    .A(net334),
    .B(net335));
 sg13g2_and4_1 _1142_ (.A(net334),
    .B(net336),
    .C(net331),
    .D(net332),
    .X(_0480_));
 sg13g2_and2_1 _1143_ (.A(net329),
    .B(_0480_),
    .X(_0481_));
 sg13g2_nand4_1 _1144_ (.B(net329),
    .C(net326),
    .A(net327),
    .Y(_0482_),
    .D(_0480_));
 sg13g2_nor2_1 _1145_ (.A(_0257_),
    .B(_0482_),
    .Y(_0483_));
 sg13g2_xnor2_1 _1146_ (.Y(_0484_),
    .A(_0260_),
    .B(_0483_));
 sg13g2_a21oi_1 _1147_ (.A1(_0257_),
    .A2(net312),
    .Y(_0485_),
    .B1(net307));
 sg13g2_o21ai_1 _1148_ (.B1(_0485_),
    .Y(_0486_),
    .A1(net312),
    .A2(_0484_));
 sg13g2_a21oi_1 _1149_ (.A1(net166),
    .A2(net307),
    .Y(_0487_),
    .B1(net302));
 sg13g2_a221oi_1 _1150_ (.B2(_0487_),
    .C1(_0423_),
    .B1(_0486_),
    .A1(net302),
    .Y(_0488_),
    .A2(net181));
 sg13g2_nor3_1 _1151_ (.A(net263),
    .B(_0478_),
    .C(_0488_),
    .Y(_0489_));
 sg13g2_a21oi_1 _1152_ (.A1(_0260_),
    .A2(net263),
    .Y(_0020_),
    .B1(_0489_));
 sg13g2_nand2_1 _1153_ (.Y(_0490_),
    .A(\cpu0.dr[9] ),
    .B(\cpu0.ac[9] ));
 sg13g2_nor2_1 _1154_ (.A(\cpu0.dr[9] ),
    .B(\cpu0.ac[9] ),
    .Y(_0491_));
 sg13g2_nand2_1 _1155_ (.Y(_0492_),
    .A(_0242_),
    .B(_0259_));
 sg13g2_o21ai_1 _1156_ (.B1(_0490_),
    .Y(_0493_),
    .A1(_0465_),
    .A2(_0491_));
 sg13g2_a21oi_1 _1157_ (.A1(_0469_),
    .A2(_0492_),
    .Y(_0494_),
    .B1(_0493_));
 sg13g2_nand2_1 _1158_ (.Y(_0495_),
    .A(net284),
    .B(_0494_));
 sg13g2_a22oi_1 _1159_ (.Y(_0496_),
    .B1(_0490_),
    .B2(_0492_),
    .A2(\cpu0.ac[8] ),
    .A1(\cpu0.dr[8] ));
 sg13g2_a22oi_1 _1160_ (.Y(_0497_),
    .B1(_0496_),
    .B2(_0472_),
    .A2(_0495_),
    .A1(_0490_));
 sg13g2_a21oi_1 _1161_ (.A1(_0242_),
    .A2(net288),
    .Y(_0498_),
    .B1(net343));
 sg13g2_o21ai_1 _1162_ (.B1(_0498_),
    .Y(_0499_),
    .A1(net288),
    .A2(_0497_));
 sg13g2_nor4_2 _1163_ (.A(_0257_),
    .B(_0259_),
    .C(_0260_),
    .Y(_0500_),
    .D(_0482_));
 sg13g2_a21oi_1 _1164_ (.A1(\cpu0.ac[8] ),
    .A2(_0483_),
    .Y(_0501_),
    .B1(\cpu0.ac[9] ));
 sg13g2_o21ai_1 _1165_ (.B1(_0270_),
    .Y(_0502_),
    .A1(_0500_),
    .A2(_0501_));
 sg13g2_a21oi_1 _1166_ (.A1(_0260_),
    .A2(net312),
    .Y(_0503_),
    .B1(net307));
 sg13g2_a221oi_1 _1167_ (.B2(_0503_),
    .C1(net302),
    .B1(_0502_),
    .A1(net351),
    .Y(_0504_),
    .A2(net308));
 sg13g2_a21oi_1 _1168_ (.A1(net302),
    .A2(net166),
    .Y(_0505_),
    .B1(_0504_));
 sg13g2_a21oi_1 _1169_ (.A1(_0422_),
    .A2(_0505_),
    .Y(_0506_),
    .B1(net263));
 sg13g2_a22oi_1 _1170_ (.Y(_0021_),
    .B1(_0499_),
    .B2(_0506_),
    .A2(_0429_),
    .A1(_0259_));
 sg13g2_nand2_1 _1171_ (.Y(_0507_),
    .A(\cpu0.dr[10] ),
    .B(net351));
 sg13g2_xnor2_1 _1172_ (.Y(_0508_),
    .A(\cpu0.dr[10] ),
    .B(net351));
 sg13g2_xnor2_1 _1173_ (.Y(_0509_),
    .A(_0494_),
    .B(_0508_));
 sg13g2_nand2_1 _1174_ (.Y(_0510_),
    .A(net281),
    .B(_0507_));
 sg13g2_a21oi_1 _1175_ (.A1(net284),
    .A2(_0509_),
    .Y(_0511_),
    .B1(net288));
 sg13g2_a22oi_1 _1176_ (.Y(_0512_),
    .B1(_0510_),
    .B2(_0511_),
    .A2(net288),
    .A1(net143));
 sg13g2_or2_1 _1177_ (.X(_0513_),
    .B(_0512_),
    .A(net343));
 sg13g2_nand2_1 _1178_ (.Y(_0514_),
    .A(net351),
    .B(_0500_));
 sg13g2_xnor2_1 _1179_ (.Y(_0515_),
    .A(net351),
    .B(_0500_));
 sg13g2_mux2_1 _1180_ (.A0(_0259_),
    .A1(_0515_),
    .S(_0270_),
    .X(_0516_));
 sg13g2_a21oi_1 _1181_ (.A1(net350),
    .A2(net308),
    .Y(_0517_),
    .B1(net303));
 sg13g2_o21ai_1 _1182_ (.B1(_0517_),
    .Y(_0518_),
    .A1(net308),
    .A2(_0516_));
 sg13g2_a21oi_1 _1183_ (.A1(net303),
    .A2(net197),
    .Y(_0519_),
    .B1(_0423_));
 sg13g2_a21oi_1 _1184_ (.A1(_0518_),
    .A2(_0519_),
    .Y(_0520_),
    .B1(net263));
 sg13g2_a22oi_1 _1185_ (.Y(_0022_),
    .B1(_0513_),
    .B2(_0520_),
    .A2(net263),
    .A1(_0262_));
 sg13g2_a21oi_1 _1186_ (.A1(net150),
    .A2(net350),
    .Y(_0521_),
    .B1(net284));
 sg13g2_xor2_1 _1187_ (.B(net350),
    .A(\cpu0.dr[11] ),
    .X(_0522_));
 sg13g2_o21ai_1 _1188_ (.B1(_0507_),
    .Y(_0523_),
    .A1(_0494_),
    .A2(_0508_));
 sg13g2_xnor2_1 _1189_ (.Y(_0524_),
    .A(_0522_),
    .B(_0523_));
 sg13g2_a21oi_1 _1190_ (.A1(_0470_),
    .A2(_0524_),
    .Y(_0525_),
    .B1(_0521_));
 sg13g2_a21oi_1 _1191_ (.A1(_0244_),
    .A2(net287),
    .Y(_0526_),
    .B1(net343));
 sg13g2_o21ai_1 _1192_ (.B1(_0526_),
    .Y(_0527_),
    .A1(net288),
    .A2(_0525_));
 sg13g2_xnor2_1 _1193_ (.Y(_0528_),
    .A(net350),
    .B(_0514_));
 sg13g2_a21oi_1 _1194_ (.A1(_0262_),
    .A2(net313),
    .Y(_0529_),
    .B1(net308));
 sg13g2_o21ai_1 _1195_ (.B1(_0529_),
    .Y(_0530_),
    .A1(net313),
    .A2(_0528_));
 sg13g2_a21oi_1 _1196_ (.A1(net349),
    .A2(net308),
    .Y(_0531_),
    .B1(net303));
 sg13g2_a22oi_1 _1197_ (.Y(_0532_),
    .B1(_0530_),
    .B2(_0531_),
    .A2(net202),
    .A1(net303));
 sg13g2_a21oi_1 _1198_ (.A1(_0422_),
    .A2(_0532_),
    .Y(_0533_),
    .B1(net263));
 sg13g2_a22oi_1 _1199_ (.Y(_0023_),
    .B1(_0527_),
    .B2(_0533_),
    .A2(net263),
    .A1(_0261_));
 sg13g2_nand4_1 _1200_ (.B(net351),
    .C(net349),
    .A(\cpu0.ac[11] ),
    .Y(_0534_),
    .D(_0500_));
 sg13g2_o21ai_1 _1201_ (.B1(_0264_),
    .Y(_0535_),
    .A1(_0261_),
    .A2(_0514_));
 sg13g2_a21o_1 _1202_ (.A2(_0535_),
    .A1(_0534_),
    .B1(net313),
    .X(_0536_));
 sg13g2_o21ai_1 _1203_ (.B1(_0536_),
    .Y(_0537_),
    .A1(net350),
    .A2(_0270_));
 sg13g2_a21oi_1 _1204_ (.A1(net162),
    .A2(net305),
    .Y(_0538_),
    .B1(net299));
 sg13g2_o21ai_1 _1205_ (.B1(_0538_),
    .Y(_0539_),
    .A1(net305),
    .A2(_0537_));
 sg13g2_a21oi_1 _1206_ (.A1(net300),
    .A2(net196),
    .Y(_0540_),
    .B1(_0423_));
 sg13g2_nor2b_1 _1207_ (.A(_0508_),
    .B_N(_0522_),
    .Y(_0541_));
 sg13g2_and4_1 _1208_ (.A(_0466_),
    .B(_0490_),
    .C(_0492_),
    .D(_0541_),
    .X(_0542_));
 sg13g2_o21ai_1 _1209_ (.B1(_0542_),
    .Y(_0543_),
    .A1(_0457_),
    .A2(_0464_));
 sg13g2_a21oi_1 _1210_ (.A1(_0244_),
    .A2(_0261_),
    .Y(_0544_),
    .B1(_0507_));
 sg13g2_a221oi_1 _1211_ (.B2(_0541_),
    .C1(_0544_),
    .B1(_0493_),
    .A1(\cpu0.dr[11] ),
    .Y(_0545_),
    .A2(net350));
 sg13g2_nand2_1 _1212_ (.Y(_0546_),
    .A(\cpu0.dr[12] ),
    .B(net349));
 sg13g2_xnor2_1 _1213_ (.Y(_0547_),
    .A(\cpu0.dr[12] ),
    .B(net349));
 sg13g2_a21oi_1 _1214_ (.A1(_0543_),
    .A2(_0545_),
    .Y(_0548_),
    .B1(_0547_));
 sg13g2_and3_1 _1215_ (.X(_0549_),
    .A(_0543_),
    .B(_0545_),
    .C(_0547_));
 sg13g2_o21ai_1 _1216_ (.B1(_0470_),
    .Y(_0550_),
    .A1(_0548_),
    .A2(_0549_));
 sg13g2_o21ai_1 _1217_ (.B1(net133),
    .Y(_0551_),
    .A1(net349),
    .A2(net287));
 sg13g2_a21oi_1 _1218_ (.A1(_0471_),
    .A2(_0551_),
    .Y(_0552_),
    .B1(net343));
 sg13g2_a221oi_1 _1219_ (.B2(_0552_),
    .C1(net264),
    .B1(_0550_),
    .A1(_0539_),
    .Y(_0553_),
    .A2(_0540_));
 sg13g2_a21oi_1 _1220_ (.A1(_0264_),
    .A2(net263),
    .Y(_0024_),
    .B1(_0553_));
 sg13g2_nand2_1 _1221_ (.Y(_0554_),
    .A(_0263_),
    .B(_0534_));
 sg13g2_nor2_1 _1222_ (.A(_0263_),
    .B(_0534_),
    .Y(_0555_));
 sg13g2_nor2_1 _1223_ (.A(net311),
    .B(_0555_),
    .Y(_0556_));
 sg13g2_a22oi_1 _1224_ (.Y(_0557_),
    .B1(_0554_),
    .B2(_0556_),
    .A2(net311),
    .A1(net349));
 sg13g2_a21oi_1 _1225_ (.A1(\cpu0.ac[14] ),
    .A2(net306),
    .Y(_0558_),
    .B1(net299));
 sg13g2_o21ai_1 _1226_ (.B1(_0558_),
    .Y(_0559_),
    .A1(net306),
    .A2(_0557_));
 sg13g2_a21oi_1 _1227_ (.A1(net299),
    .A2(net162),
    .Y(_0560_),
    .B1(_0423_));
 sg13g2_nor2_1 _1228_ (.A(_0245_),
    .B(_0263_),
    .Y(_0561_));
 sg13g2_xnor2_1 _1229_ (.Y(_0562_),
    .A(\cpu0.dr[13] ),
    .B(\cpu0.ac[13] ));
 sg13g2_a21oi_1 _1230_ (.A1(\cpu0.dr[12] ),
    .A2(net349),
    .Y(_0563_),
    .B1(_0548_));
 sg13g2_xnor2_1 _1231_ (.Y(_0564_),
    .A(_0562_),
    .B(_0563_));
 sg13g2_a21oi_1 _1232_ (.A1(net282),
    .A2(_0561_),
    .Y(_0565_),
    .B1(net287));
 sg13g2_o21ai_1 _1233_ (.B1(_0565_),
    .Y(_0566_),
    .A1(net282),
    .A2(_0564_));
 sg13g2_a21oi_1 _1234_ (.A1(_0245_),
    .A2(net287),
    .Y(_0567_),
    .B1(net343));
 sg13g2_a221oi_1 _1235_ (.B2(_0567_),
    .C1(net264),
    .B1(_0566_),
    .A1(_0559_),
    .Y(_0568_),
    .A2(_0560_));
 sg13g2_a21oi_1 _1236_ (.A1(_0263_),
    .A2(net264),
    .Y(_0025_),
    .B1(_0568_));
 sg13g2_xnor2_1 _1237_ (.Y(_0569_),
    .A(_0266_),
    .B(_0555_));
 sg13g2_a21oi_1 _1238_ (.A1(_0263_),
    .A2(net311),
    .Y(_0570_),
    .B1(net306));
 sg13g2_o21ai_1 _1239_ (.B1(_0570_),
    .Y(_0571_),
    .A1(net311),
    .A2(_0569_));
 sg13g2_a21oi_1 _1240_ (.A1(\cpu0.ac[15] ),
    .A2(net305),
    .Y(_0572_),
    .B1(net300));
 sg13g2_a221oi_1 _1241_ (.B2(_0572_),
    .C1(_0423_),
    .B1(_0571_),
    .A1(net300),
    .Y(_0573_),
    .A2(net182));
 sg13g2_nand2_1 _1242_ (.Y(_0574_),
    .A(\cpu0.dr[14] ),
    .B(\cpu0.ac[14] ));
 sg13g2_xnor2_1 _1243_ (.Y(_0575_),
    .A(\cpu0.dr[14] ),
    .B(\cpu0.ac[14] ));
 sg13g2_or2_1 _1244_ (.X(_0576_),
    .B(_0562_),
    .A(_0547_));
 sg13g2_a21o_1 _1245_ (.A2(_0545_),
    .A1(_0543_),
    .B1(_0576_),
    .X(_0577_));
 sg13g2_a21oi_1 _1246_ (.A1(_0245_),
    .A2(_0263_),
    .Y(_0578_),
    .B1(_0546_));
 sg13g2_nor2_1 _1247_ (.A(_0561_),
    .B(_0578_),
    .Y(_0579_));
 sg13g2_a21o_1 _1248_ (.A2(_0579_),
    .A1(_0577_),
    .B1(_0575_),
    .X(_0580_));
 sg13g2_nand3_1 _1249_ (.B(_0577_),
    .C(_0579_),
    .A(_0575_),
    .Y(_0581_));
 sg13g2_a21oi_1 _1250_ (.A1(_0580_),
    .A2(_0581_),
    .Y(_0582_),
    .B1(net282));
 sg13g2_a21oi_1 _1251_ (.A1(net282),
    .A2(_0574_),
    .Y(_0583_),
    .B1(net287));
 sg13g2_nand2b_1 _1252_ (.Y(_0584_),
    .B(_0583_),
    .A_N(_0582_));
 sg13g2_nand2_1 _1253_ (.Y(_0585_),
    .A(\cpu0.dr[14] ),
    .B(net287));
 sg13g2_a21o_1 _1254_ (.A2(_0585_),
    .A1(_0584_),
    .B1(net342),
    .X(_0586_));
 sg13g2_nor2_1 _1255_ (.A(net264),
    .B(_0573_),
    .Y(_0587_));
 sg13g2_a22oi_1 _1256_ (.Y(_0026_),
    .B1(_0586_),
    .B2(_0587_),
    .A2(net264),
    .A1(_0266_));
 sg13g2_nor2_1 _1257_ (.A(_0246_),
    .B(_0265_),
    .Y(_0588_));
 sg13g2_xnor2_1 _1258_ (.Y(_0589_),
    .A(net92),
    .B(\cpu0.ac[15] ));
 sg13g2_a21oi_1 _1259_ (.A1(_0574_),
    .A2(_0580_),
    .Y(_0590_),
    .B1(_0589_));
 sg13g2_and3_1 _1260_ (.X(_0591_),
    .A(_0574_),
    .B(_0580_),
    .C(_0589_));
 sg13g2_nor3_1 _1261_ (.A(net282),
    .B(_0590_),
    .C(_0591_),
    .Y(_0592_));
 sg13g2_a21o_1 _1262_ (.A2(_0588_),
    .A1(net282),
    .B1(net287),
    .X(_0593_));
 sg13g2_a21oi_1 _1263_ (.A1(_0246_),
    .A2(net287),
    .Y(_0594_),
    .B1(net342));
 sg13g2_o21ai_1 _1264_ (.B1(_0594_),
    .Y(_0595_),
    .A1(_0592_),
    .A2(_0593_));
 sg13g2_nor2_1 _1265_ (.A(_0266_),
    .B(_0556_),
    .Y(_0596_));
 sg13g2_nor2_1 _1266_ (.A(_0265_),
    .B(net311),
    .Y(_0597_));
 sg13g2_xnor2_1 _1267_ (.Y(_0598_),
    .A(_0596_),
    .B(_0597_));
 sg13g2_a21oi_1 _1268_ (.A1(net135),
    .A2(net305),
    .Y(_0599_),
    .B1(net300));
 sg13g2_o21ai_1 _1269_ (.B1(_0599_),
    .Y(_0600_),
    .A1(net305),
    .A2(_0598_));
 sg13g2_a21oi_1 _1270_ (.A1(net300),
    .A2(net184),
    .Y(_0601_),
    .B1(_0423_));
 sg13g2_a21oi_1 _1271_ (.A1(_0600_),
    .A2(_0601_),
    .Y(_0602_),
    .B1(net264));
 sg13g2_a22oi_1 _1272_ (.Y(_0027_),
    .B1(_0595_),
    .B2(_0602_),
    .A2(net264),
    .A1(_0265_));
 sg13g2_and2_1 _1273_ (.A(net348),
    .B(net278),
    .X(_0028_));
 sg13g2_and2_1 _1274_ (.A(net40),
    .B(_0406_),
    .X(_0029_));
 sg13g2_and2_1 _1275_ (.A(net50),
    .B(net278),
    .X(_0030_));
 sg13g2_nor2_1 _1276_ (.A(net294),
    .B(\cpu0.rstT ),
    .Y(_0031_));
 sg13g2_and2_1 _1277_ (.A(net338),
    .B(net278),
    .X(_0032_));
 sg13g2_nor2_1 _1278_ (.A(_0237_),
    .B(\cpu0.rstT ),
    .Y(_0033_));
 sg13g2_and2_1 _1279_ (.A(net88),
    .B(net278),
    .X(_0034_));
 sg13g2_and2_1 _1280_ (.A(net72),
    .B(net278),
    .X(_0035_));
 sg13g2_and2_1 _1281_ (.A(net54),
    .B(net278),
    .X(_0036_));
 sg13g2_and2_1 _1282_ (.A(net74),
    .B(net278),
    .X(_0037_));
 sg13g2_and2_1 _1283_ (.A(net340),
    .B(net310),
    .X(_0603_));
 sg13g2_nand2_1 _1284_ (.Y(_0604_),
    .A(net305),
    .B(_0407_));
 sg13g2_mux2_1 _1285_ (.A0(net335),
    .A1(net94),
    .S(_0604_),
    .X(_0038_));
 sg13g2_nand2_1 _1286_ (.Y(_0605_),
    .A(net10),
    .B(\cpu0.ir[11] ));
 sg13g2_a21o_1 _1287_ (.A2(_0605_),
    .A1(_0301_),
    .B1(_0428_),
    .X(_0606_));
 sg13g2_nand2_1 _1288_ (.Y(_0607_),
    .A(net335),
    .B(net262));
 sg13g2_a21oi_1 _1289_ (.A1(net335),
    .A2(net283),
    .Y(_0608_),
    .B1(net319));
 sg13g2_nand3_1 _1290_ (.B(net335),
    .C(net283),
    .A(\cpu0.dr[0] ),
    .Y(_0609_));
 sg13g2_o21ai_1 _1291_ (.B1(_0609_),
    .Y(_0610_),
    .A1(net335),
    .A2(net283));
 sg13g2_a21oi_1 _1292_ (.A1(_0474_),
    .A2(_0610_),
    .Y(_0611_),
    .B1(_0608_));
 sg13g2_nand2_1 _1293_ (.Y(_0612_),
    .A(net333),
    .B(net306));
 sg13g2_o21ai_1 _1294_ (.B1(_0612_),
    .Y(_0613_),
    .A1(_0250_),
    .A2(net306));
 sg13g2_nor3_1 _1295_ (.A(net299),
    .B(_0396_),
    .C(_0613_),
    .Y(_0614_));
 sg13g2_o21ai_1 _1296_ (.B1(net335),
    .Y(_0615_),
    .A1(net299),
    .A2(_0396_));
 sg13g2_nand3_1 _1297_ (.B(_0272_),
    .C(_0615_),
    .A(net296),
    .Y(_0616_));
 sg13g2_a21oi_1 _1298_ (.A1(net297),
    .A2(net2),
    .Y(_0617_),
    .B1(net294));
 sg13g2_o21ai_1 _1299_ (.B1(_0617_),
    .Y(_0618_),
    .A1(_0614_),
    .A2(_0616_));
 sg13g2_o21ai_1 _1300_ (.B1(_0618_),
    .Y(_0619_),
    .A1(net343),
    .A2(_0611_));
 sg13g2_o21ai_1 _1301_ (.B1(_0607_),
    .Y(_0039_),
    .A1(net262),
    .A2(_0619_));
 sg13g2_a21oi_1 _1302_ (.A1(net3),
    .A2(_0301_),
    .Y(_0620_),
    .B1(net260));
 sg13g2_a21oi_1 _1303_ (.A1(_0431_),
    .A2(_0433_),
    .Y(_0621_),
    .B1(_0432_));
 sg13g2_nand2_1 _1304_ (.Y(_0622_),
    .A(_0434_),
    .B(net283));
 sg13g2_a22oi_1 _1305_ (.Y(_0623_),
    .B1(net286),
    .B2(net199),
    .A2(net281),
    .A1(_0430_));
 sg13g2_o21ai_1 _1306_ (.B1(_0623_),
    .Y(_0624_),
    .A1(_0621_),
    .A2(_0622_));
 sg13g2_a21oi_1 _1307_ (.A1(net334),
    .A2(net336),
    .Y(_0625_),
    .B1(net314));
 sg13g2_or2_1 _1308_ (.X(_0626_),
    .B(net336),
    .A(net333));
 sg13g2_a22oi_1 _1309_ (.Y(_0627_),
    .B1(_0625_),
    .B2(_0626_),
    .A2(net314),
    .A1(net336));
 sg13g2_a21oi_1 _1310_ (.A1(net332),
    .A2(net309),
    .Y(_0628_),
    .B1(net304));
 sg13g2_o21ai_1 _1311_ (.B1(_0628_),
    .Y(_0629_),
    .A1(net309),
    .A2(_0627_));
 sg13g2_a21oi_1 _1312_ (.A1(net304),
    .A2(net334),
    .Y(_0630_),
    .B1(_0424_));
 sg13g2_a22oi_1 _1313_ (.Y(_0631_),
    .B1(_0629_),
    .B2(_0630_),
    .A2(_0624_),
    .A1(net294));
 sg13g2_a22oi_1 _1314_ (.Y(_0040_),
    .B1(_0620_),
    .B2(_0631_),
    .A2(net260),
    .A1(_0252_));
 sg13g2_a21oi_1 _1315_ (.A1(_0435_),
    .A2(_0437_),
    .Y(_0632_),
    .B1(net281));
 sg13g2_nand2_1 _1316_ (.Y(_0633_),
    .A(_0438_),
    .B(_0632_));
 sg13g2_nor2_1 _1317_ (.A(_0436_),
    .B(net284),
    .Y(_0634_));
 sg13g2_nor2_1 _1318_ (.A(net286),
    .B(_0634_),
    .Y(_0635_));
 sg13g2_o21ai_1 _1319_ (.B1(net294),
    .Y(_0636_),
    .A1(net188),
    .A2(_0474_));
 sg13g2_a21oi_1 _1320_ (.A1(_0633_),
    .A2(_0635_),
    .Y(_0637_),
    .B1(_0636_));
 sg13g2_xnor2_1 _1321_ (.Y(_0638_),
    .A(net332),
    .B(_0479_));
 sg13g2_a21oi_1 _1322_ (.A1(_0252_),
    .A2(net314),
    .Y(_0639_),
    .B1(net310));
 sg13g2_o21ai_1 _1323_ (.B1(_0639_),
    .Y(_0640_),
    .A1(net314),
    .A2(_0638_));
 sg13g2_a21oi_1 _1324_ (.A1(net331),
    .A2(net310),
    .Y(_0641_),
    .B1(net304));
 sg13g2_a221oi_1 _1325_ (.B2(_0641_),
    .C1(_0424_),
    .B1(_0640_),
    .A1(net304),
    .Y(_0642_),
    .A2(net207));
 sg13g2_nand2_1 _1326_ (.Y(_0643_),
    .A(net4),
    .B(_0301_));
 sg13g2_nor3_1 _1327_ (.A(net260),
    .B(_0637_),
    .C(_0642_),
    .Y(_0644_));
 sg13g2_a22oi_1 _1328_ (.Y(_0041_),
    .B1(_0643_),
    .B2(_0644_),
    .A2(net260),
    .A1(_0254_));
 sg13g2_o21ai_1 _1329_ (.B1(_0439_),
    .Y(_0645_),
    .A1(_0443_),
    .A2(net281));
 sg13g2_nand2_1 _1330_ (.Y(_0646_),
    .A(_0440_),
    .B(_0442_));
 sg13g2_nand4_1 _1331_ (.B(_0438_),
    .C(net283),
    .A(_0436_),
    .Y(_0647_),
    .D(_0646_));
 sg13g2_a21oi_1 _1332_ (.A1(_0645_),
    .A2(_0647_),
    .Y(_0648_),
    .B1(net289));
 sg13g2_o21ai_1 _1333_ (.B1(net295),
    .Y(_0649_),
    .A1(net218),
    .A2(_0474_));
 sg13g2_nor2_1 _1334_ (.A(_0648_),
    .B(_0649_),
    .Y(_0650_));
 sg13g2_nand2_1 _1335_ (.Y(_0651_),
    .A(\cpu0.ac[3] ),
    .B(_0270_));
 sg13g2_o21ai_1 _1336_ (.B1(_0651_),
    .Y(_0652_),
    .A1(_0254_),
    .A2(_0625_));
 sg13g2_a21oi_1 _1337_ (.A1(_0270_),
    .A2(_0480_),
    .Y(_0653_),
    .B1(net309));
 sg13g2_nand2_1 _1338_ (.Y(_0654_),
    .A(_0652_),
    .B(_0653_));
 sg13g2_a21oi_1 _1339_ (.A1(net330),
    .A2(net309),
    .Y(_0655_),
    .B1(net304));
 sg13g2_a221oi_1 _1340_ (.B2(_0655_),
    .C1(_0424_),
    .B1(_0654_),
    .A1(net304),
    .Y(_0656_),
    .A2(net331));
 sg13g2_nand2_1 _1341_ (.Y(_0657_),
    .A(net5),
    .B(_0301_));
 sg13g2_nor3_1 _1342_ (.A(net260),
    .B(_0650_),
    .C(_0656_),
    .Y(_0658_));
 sg13g2_a22oi_1 _1343_ (.Y(_0042_),
    .B1(_0657_),
    .B2(net219),
    .A2(net260),
    .A1(_0253_));
 sg13g2_a22oi_1 _1344_ (.Y(_0659_),
    .B1(net286),
    .B2(net153),
    .A2(net281),
    .A1(_0453_));
 sg13g2_a21oi_1 _1345_ (.A1(_0443_),
    .A2(_0455_),
    .Y(_0660_),
    .B1(net281));
 sg13g2_o21ai_1 _1346_ (.B1(_0660_),
    .Y(_0661_),
    .A1(_0443_),
    .A2(_0455_));
 sg13g2_a21o_1 _1347_ (.A2(_0661_),
    .A1(_0659_),
    .B1(net344),
    .X(_0662_));
 sg13g2_nor2_1 _1348_ (.A(net329),
    .B(_0480_),
    .Y(_0663_));
 sg13g2_nor3_1 _1349_ (.A(net314),
    .B(_0481_),
    .C(_0663_),
    .Y(_0664_));
 sg13g2_a21oi_1 _1350_ (.A1(net331),
    .A2(net314),
    .Y(_0665_),
    .B1(_0664_));
 sg13g2_a21oi_1 _1351_ (.A1(net328),
    .A2(net309),
    .Y(_0666_),
    .B1(net301));
 sg13g2_o21ai_1 _1352_ (.B1(_0666_),
    .Y(_0667_),
    .A1(net309),
    .A2(_0665_));
 sg13g2_a21oi_1 _1353_ (.A1(net301),
    .A2(net330),
    .Y(_0668_),
    .B1(_0424_));
 sg13g2_a221oi_1 _1354_ (.B2(_0668_),
    .C1(net261),
    .B1(_0667_),
    .A1(net6),
    .Y(_0669_),
    .A2(_0301_));
 sg13g2_a22oi_1 _1355_ (.Y(_0043_),
    .B1(_0662_),
    .B2(_0669_),
    .A2(net260),
    .A1(_0256_));
 sg13g2_a21oi_1 _1356_ (.A1(_0443_),
    .A2(_0455_),
    .Y(_0670_),
    .B1(_0453_));
 sg13g2_o21ai_1 _1357_ (.B1(net283),
    .Y(_0671_),
    .A1(_0451_),
    .A2(_0670_));
 sg13g2_and2_1 _1358_ (.A(net283),
    .B(_0670_),
    .X(_0672_));
 sg13g2_a22oi_1 _1359_ (.Y(_0673_),
    .B1(_0672_),
    .B2(_0452_),
    .A2(_0671_),
    .A1(_0450_));
 sg13g2_a21oi_1 _1360_ (.A1(_0239_),
    .A2(net286),
    .Y(_0674_),
    .B1(net344));
 sg13g2_o21ai_1 _1361_ (.B1(_0674_),
    .Y(_0675_),
    .A1(net286),
    .A2(_0673_));
 sg13g2_or2_1 _1362_ (.X(_0676_),
    .B(_0481_),
    .A(net328));
 sg13g2_a21oi_1 _1363_ (.A1(net328),
    .A2(_0481_),
    .Y(_0677_),
    .B1(net312));
 sg13g2_a22oi_1 _1364_ (.Y(_0678_),
    .B1(_0676_),
    .B2(_0677_),
    .A2(net312),
    .A1(net330));
 sg13g2_a21oi_1 _1365_ (.A1(net326),
    .A2(net307),
    .Y(_0679_),
    .B1(net301));
 sg13g2_o21ai_1 _1366_ (.B1(_0679_),
    .Y(_0680_),
    .A1(net309),
    .A2(_0678_));
 sg13g2_a21oi_1 _1367_ (.A1(net301),
    .A2(net328),
    .Y(_0681_),
    .B1(_0424_));
 sg13g2_a221oi_1 _1368_ (.B2(_0681_),
    .C1(net261),
    .B1(_0680_),
    .A1(net7),
    .Y(_0682_),
    .A2(_0301_));
 sg13g2_a22oi_1 _1369_ (.Y(_0044_),
    .B1(_0675_),
    .B2(_0682_),
    .A2(net261),
    .A1(_0255_));
 sg13g2_o21ai_1 _1370_ (.B1(_0450_),
    .Y(_0683_),
    .A1(_0451_),
    .A2(_0670_));
 sg13g2_xor2_1 _1371_ (.B(_0683_),
    .A(_0448_),
    .X(_0684_));
 sg13g2_o21ai_1 _1372_ (.B1(_0474_),
    .Y(_0685_),
    .A1(_0446_),
    .A2(net283));
 sg13g2_a21oi_1 _1373_ (.A1(net284),
    .A2(_0684_),
    .Y(_0686_),
    .B1(_0685_));
 sg13g2_a21oi_1 _1374_ (.A1(net174),
    .A2(net286),
    .Y(_0687_),
    .B1(_0686_));
 sg13g2_or2_1 _1375_ (.X(_0688_),
    .B(_0687_),
    .A(net344));
 sg13g2_a21o_1 _1376_ (.A2(_0481_),
    .A1(net328),
    .B1(\cpu0.ac[6] ),
    .X(_0689_));
 sg13g2_and2_1 _1377_ (.A(_0482_),
    .B(_0689_),
    .X(_0690_));
 sg13g2_a21oi_1 _1378_ (.A1(_0255_),
    .A2(net312),
    .Y(_0691_),
    .B1(net307));
 sg13g2_o21ai_1 _1379_ (.B1(_0691_),
    .Y(_0692_),
    .A1(net312),
    .A2(_0690_));
 sg13g2_a21oi_1 _1380_ (.A1(net325),
    .A2(net307),
    .Y(_0693_),
    .B1(net301));
 sg13g2_nand2_1 _1381_ (.Y(_0694_),
    .A(_0692_),
    .B(_0693_));
 sg13g2_a21oi_1 _1382_ (.A1(net301),
    .A2(net210),
    .Y(_0695_),
    .B1(_0424_));
 sg13g2_a221oi_1 _1383_ (.B2(_0695_),
    .C1(net261),
    .B1(_0694_),
    .A1(net8),
    .Y(_0696_),
    .A2(_0301_));
 sg13g2_a22oi_1 _1384_ (.Y(_0045_),
    .B1(_0688_),
    .B2(_0696_),
    .A2(net261),
    .A1(_0258_));
 sg13g2_and2_1 _1385_ (.A(_0444_),
    .B(net281),
    .X(_0697_));
 sg13g2_a21oi_1 _1386_ (.A1(_0447_),
    .A2(_0683_),
    .Y(_0698_),
    .B1(_0446_));
 sg13g2_xnor2_1 _1387_ (.Y(_0699_),
    .A(_0445_),
    .B(_0698_));
 sg13g2_a21oi_1 _1388_ (.A1(net284),
    .A2(_0699_),
    .Y(_0700_),
    .B1(_0697_));
 sg13g2_a21oi_1 _1389_ (.A1(_0241_),
    .A2(net286),
    .Y(_0701_),
    .B1(net343));
 sg13g2_o21ai_1 _1390_ (.B1(_0701_),
    .Y(_0702_),
    .A1(net286),
    .A2(_0700_));
 sg13g2_xnor2_1 _1391_ (.Y(_0703_),
    .A(net325),
    .B(_0482_));
 sg13g2_a21oi_1 _1392_ (.A1(_0258_),
    .A2(net313),
    .Y(_0704_),
    .B1(net307));
 sg13g2_o21ai_1 _1393_ (.B1(_0704_),
    .Y(_0705_),
    .A1(net312),
    .A2(_0703_));
 sg13g2_a21oi_1 _1394_ (.A1(\cpu0.ac[8] ),
    .A2(net307),
    .Y(_0706_),
    .B1(net301));
 sg13g2_nand2_1 _1395_ (.Y(_0707_),
    .A(_0705_),
    .B(_0706_));
 sg13g2_a21oi_1 _1396_ (.A1(net301),
    .A2(net214),
    .Y(_0708_),
    .B1(_0424_));
 sg13g2_a221oi_1 _1397_ (.B2(_0708_),
    .C1(net261),
    .B1(_0707_),
    .A1(net9),
    .Y(_0709_),
    .A2(_0301_));
 sg13g2_a22oi_1 _1398_ (.Y(_0046_),
    .B1(_0702_),
    .B2(_0709_),
    .A2(net260),
    .A1(_0257_));
 sg13g2_a21o_1 _1399_ (.A2(_0402_),
    .A1(net294),
    .B1(_0407_),
    .X(_0710_));
 sg13g2_o21ai_1 _1400_ (.B1(_0416_),
    .Y(_0711_),
    .A1(_0419_),
    .A2(net282));
 sg13g2_nand2b_2 _1401_ (.Y(_0712_),
    .B(net342),
    .A_N(\cpu0.ir[10] ));
 sg13g2_nand3b_1 _1402_ (.B(_0248_),
    .C(_0299_),
    .Y(_0713_),
    .A_N(_0712_));
 sg13g2_o21ai_1 _1403_ (.B1(net338),
    .Y(_0714_),
    .A1(\cpu0.ir[15] ),
    .A2(_0300_));
 sg13g2_nand4_1 _1404_ (.B(_0711_),
    .C(_0713_),
    .A(_0710_),
    .Y(_0715_),
    .D(_0714_));
 sg13g2_o21ai_1 _1405_ (.B1(_0416_),
    .Y(_0716_),
    .A1(_0588_),
    .A2(_0590_));
 sg13g2_nor2_1 _1406_ (.A(net135),
    .B(_0712_),
    .Y(_0717_));
 sg13g2_nor2b_1 _1407_ (.A(net94),
    .B_N(net305),
    .Y(_0718_));
 sg13g2_o21ai_1 _1408_ (.B1(net338),
    .Y(_0719_),
    .A1(net305),
    .A2(net62));
 sg13g2_nor3_1 _1409_ (.A(net342),
    .B(_0718_),
    .C(_0719_),
    .Y(_0720_));
 sg13g2_nor3_1 _1410_ (.A(_0715_),
    .B(_0717_),
    .C(_0720_),
    .Y(_0721_));
 sg13g2_a22oi_1 _1411_ (.Y(_0047_),
    .B1(_0716_),
    .B2(_0721_),
    .A2(_0715_),
    .A1(_0250_));
 sg13g2_mux2_1 _1412_ (.A0(\boot_to_cpu[0] ),
    .A1(\spi0.dataout[0] ),
    .S(net276),
    .X(_0722_));
 sg13g2_nand2_1 _1413_ (.Y(_0723_),
    .A(net295),
    .B(_0722_));
 sg13g2_nor3_1 _1414_ (.A(net296),
    .B(_0237_),
    .C(_0307_),
    .Y(_0724_));
 sg13g2_nor3_1 _1415_ (.A(net347),
    .B(net340),
    .C(_0724_),
    .Y(_0725_));
 sg13g2_a21oi_1 _1416_ (.A1(net339),
    .A2(\cpu0.ir[0] ),
    .Y(_0726_),
    .B1(net345));
 sg13g2_a221oi_1 _1417_ (.B2(_0726_),
    .C1(net271),
    .B1(_0723_),
    .A1(net345),
    .Y(_0727_),
    .A2(_0276_));
 sg13g2_a21o_1 _1418_ (.A2(net270),
    .A1(net108),
    .B1(_0727_),
    .X(_0048_));
 sg13g2_mux2_1 _1419_ (.A0(\boot_to_cpu[1] ),
    .A1(\spi0.dataout[1] ),
    .S(net276),
    .X(_0728_));
 sg13g2_a21oi_1 _1420_ (.A1(net339),
    .A2(_0251_),
    .Y(_0729_),
    .B1(net346));
 sg13g2_o21ai_1 _1421_ (.B1(_0729_),
    .Y(_0730_),
    .A1(net339),
    .A2(_0728_));
 sg13g2_a21oi_1 _1422_ (.A1(net345),
    .A2(\cpu0.pc[1] ),
    .Y(_0731_),
    .B1(net270));
 sg13g2_a22oi_1 _1423_ (.Y(_0049_),
    .B1(_0730_),
    .B2(_0731_),
    .A2(net270),
    .A1(_0277_));
 sg13g2_mux2_1 _1424_ (.A0(\boot_to_cpu[2] ),
    .A1(\spi0.dataout[2] ),
    .S(net276),
    .X(_0732_));
 sg13g2_inv_1 _1425_ (.Y(_0733_),
    .A(_0732_));
 sg13g2_a21oi_1 _1426_ (.A1(net340),
    .A2(_0267_),
    .Y(_0734_),
    .B1(net346));
 sg13g2_o21ai_1 _1427_ (.B1(_0734_),
    .Y(_0735_),
    .A1(net340),
    .A2(_0732_));
 sg13g2_a21oi_1 _1428_ (.A1(net345),
    .A2(net168),
    .Y(_0736_),
    .B1(net270));
 sg13g2_a22oi_1 _1429_ (.Y(_0050_),
    .B1(_0735_),
    .B2(_0736_),
    .A2(net270),
    .A1(_0278_));
 sg13g2_mux2_1 _1430_ (.A0(\boot_to_cpu[3] ),
    .A1(\spi0.dataout[3] ),
    .S(net276),
    .X(_0737_));
 sg13g2_a21oi_1 _1431_ (.A1(net339),
    .A2(_0268_),
    .Y(_0738_),
    .B1(net346));
 sg13g2_o21ai_1 _1432_ (.B1(_0738_),
    .Y(_0739_),
    .A1(net339),
    .A2(_0737_));
 sg13g2_a21oi_1 _1433_ (.A1(net345),
    .A2(net164),
    .Y(_0740_),
    .B1(net270));
 sg13g2_a22oi_1 _1434_ (.Y(_0051_),
    .B1(_0739_),
    .B2(_0740_),
    .A2(net270),
    .A1(_0280_));
 sg13g2_mux2_1 _1435_ (.A0(\boot_to_cpu[4] ),
    .A1(\spi0.dataout[4] ),
    .S(net276),
    .X(_0741_));
 sg13g2_a21oi_1 _1436_ (.A1(net339),
    .A2(_0269_),
    .Y(_0742_),
    .B1(net345));
 sg13g2_o21ai_1 _1437_ (.B1(_0742_),
    .Y(_0743_),
    .A1(net339),
    .A2(_0741_));
 sg13g2_a21oi_1 _1438_ (.A1(net345),
    .A2(net138),
    .Y(_0744_),
    .B1(net271));
 sg13g2_a22oi_1 _1439_ (.Y(_0052_),
    .B1(_0743_),
    .B2(net139),
    .A2(net270),
    .A1(_0281_));
 sg13g2_mux2_1 _1440_ (.A0(\boot_to_cpu[5] ),
    .A1(\spi0.dataout[5] ),
    .S(_0318_),
    .X(_0745_));
 sg13g2_a21oi_1 _1441_ (.A1(net340),
    .A2(_0271_),
    .Y(_0746_),
    .B1(net346));
 sg13g2_o21ai_1 _1442_ (.B1(_0746_),
    .Y(_0747_),
    .A1(net339),
    .A2(_0745_));
 sg13g2_a21oi_1 _1443_ (.A1(net345),
    .A2(net142),
    .Y(_0748_),
    .B1(net271));
 sg13g2_a22oi_1 _1444_ (.Y(_0053_),
    .B1(_0747_),
    .B2(_0748_),
    .A2(net271),
    .A1(_0283_));
 sg13g2_mux2_1 _1445_ (.A0(\boot_to_cpu[6] ),
    .A1(\spi0.dataout[6] ),
    .S(net276),
    .X(_0749_));
 sg13g2_nand2_1 _1446_ (.Y(_0750_),
    .A(net295),
    .B(_0749_));
 sg13g2_a21oi_1 _1447_ (.A1(net342),
    .A2(net311),
    .Y(_0751_),
    .B1(net348));
 sg13g2_a221oi_1 _1448_ (.B2(_0751_),
    .C1(net272),
    .B1(_0750_),
    .A1(net346),
    .Y(_0752_),
    .A2(_0284_));
 sg13g2_a21o_1 _1449_ (.A2(net272),
    .A1(net90),
    .B1(net132),
    .X(_0054_));
 sg13g2_mux2_1 _1450_ (.A0(\boot_to_cpu[7] ),
    .A1(\spi0.dataout[7] ),
    .S(net276),
    .X(_0753_));
 sg13g2_nand2_1 _1451_ (.Y(_0754_),
    .A(net347),
    .B(\cpu0.pc[7] ));
 sg13g2_a21oi_1 _1452_ (.A1(net295),
    .A2(_0753_),
    .Y(_0755_),
    .B1(_0603_));
 sg13g2_o21ai_1 _1453_ (.B1(_0754_),
    .Y(_0756_),
    .A1(net347),
    .A2(_0755_));
 sg13g2_mux2_1 _1454_ (.A0(_0756_),
    .A1(net119),
    .S(net272),
    .X(_0055_));
 sg13g2_and2_1 _1455_ (.A(\boot_to_cpu[8] ),
    .B(net275),
    .X(_0757_));
 sg13g2_a21oi_1 _1456_ (.A1(net340),
    .A2(_0248_),
    .Y(_0758_),
    .B1(net348));
 sg13g2_o21ai_1 _1457_ (.B1(_0758_),
    .Y(_0759_),
    .A1(net340),
    .A2(_0757_));
 sg13g2_a21oi_1 _1458_ (.A1(net347),
    .A2(\cpu0.pc[8] ),
    .Y(_0760_),
    .B1(net272));
 sg13g2_a22oi_1 _1459_ (.Y(_0056_),
    .B1(_0759_),
    .B2(_0760_),
    .A2(net272),
    .A1(_0273_));
 sg13g2_and2_1 _1460_ (.A(\boot_to_cpu[9] ),
    .B(net274),
    .X(_0761_));
 sg13g2_a21oi_1 _1461_ (.A1(net341),
    .A2(_0249_),
    .Y(_0762_),
    .B1(net347));
 sg13g2_o21ai_1 _1462_ (.B1(_0762_),
    .Y(_0763_),
    .A1(net341),
    .A2(_0761_));
 sg13g2_a21oi_1 _1463_ (.A1(net348),
    .A2(net81),
    .Y(_0764_),
    .B1(net272));
 sg13g2_a22oi_1 _1464_ (.Y(_0057_),
    .B1(_0763_),
    .B2(_0764_),
    .A2(net273),
    .A1(_0274_));
 sg13g2_and2_1 _1465_ (.A(\boot_to_cpu[10] ),
    .B(net274),
    .X(_0765_));
 sg13g2_o21ai_1 _1466_ (.B1(_0712_),
    .Y(_0766_),
    .A1(net341),
    .A2(_0765_));
 sg13g2_nor2_1 _1467_ (.A(net347),
    .B(_0766_),
    .Y(_0767_));
 sg13g2_a21oi_1 _1468_ (.A1(net347),
    .A2(\cpu0.pc[10] ),
    .Y(_0768_),
    .B1(_0767_));
 sg13g2_nand2_1 _1469_ (.Y(_0769_),
    .A(net84),
    .B(net272));
 sg13g2_o21ai_1 _1470_ (.B1(_0769_),
    .Y(_0058_),
    .A1(net272),
    .A2(_0768_));
 sg13g2_nand2_1 _1471_ (.Y(_0770_),
    .A(\boot_to_cpu[11] ),
    .B(net274));
 sg13g2_a21oi_1 _1472_ (.A1(\boot_to_cpu[11] ),
    .A2(net274),
    .Y(_0771_),
    .B1(net341));
 sg13g2_or3_1 _1473_ (.A(net348),
    .B(_0422_),
    .C(_0771_),
    .X(_0772_));
 sg13g2_a21oi_1 _1474_ (.A1(net347),
    .A2(net101),
    .Y(_0773_),
    .B1(net273));
 sg13g2_a22oi_1 _1475_ (.Y(_0059_),
    .B1(_0772_),
    .B2(_0773_),
    .A2(net273),
    .A1(_0275_));
 sg13g2_nand2_1 _1476_ (.Y(_0774_),
    .A(\cpu0.ir[6] ),
    .B(_0407_));
 sg13g2_nand2_1 _1477_ (.Y(_0775_),
    .A(net62),
    .B(_0774_));
 sg13g2_o21ai_1 _1478_ (.B1(net63),
    .Y(_0060_),
    .A1(_0265_),
    .A2(_0774_));
 sg13g2_a22oi_1 _1479_ (.Y(_0776_),
    .B1(\cpu0.t[5] ),
    .B2(_0298_),
    .A2(\cpu0.t[7] ),
    .A1(net297));
 sg13g2_nor2_1 _1480_ (.A(_0310_),
    .B(_0776_),
    .Y(_0777_));
 sg13g2_or2_1 _1481_ (.X(_0778_),
    .B(_0776_),
    .A(_0310_));
 sg13g2_a21oi_2 _1482_ (.B1(_0294_),
    .Y(_0779_),
    .A2(_0418_),
    .A1(_0306_));
 sg13g2_nor2_2 _1483_ (.A(net257),
    .B(net280),
    .Y(_0780_));
 sg13g2_nand2b_1 _1484_ (.Y(_0781_),
    .B(_0780_),
    .A_N(net319));
 sg13g2_o21ai_1 _1485_ (.B1(_0781_),
    .Y(_0782_),
    .A1(_0722_),
    .A2(_0778_));
 sg13g2_a21oi_1 _1486_ (.A1(net319),
    .A2(net280),
    .Y(_0061_),
    .B1(_0782_));
 sg13g2_nand2_1 _1487_ (.Y(_0783_),
    .A(_0728_),
    .B(net257));
 sg13g2_a21oi_1 _1488_ (.A1(net319),
    .A2(net280),
    .Y(_0784_),
    .B1(net318));
 sg13g2_nand3_1 _1489_ (.B(net319),
    .C(net280),
    .A(net318),
    .Y(_0785_));
 sg13g2_nand2_1 _1490_ (.Y(_0786_),
    .A(_0778_),
    .B(_0785_));
 sg13g2_o21ai_1 _1491_ (.B1(_0783_),
    .Y(_0062_),
    .A1(_0784_),
    .A2(_0786_));
 sg13g2_nand3_1 _1492_ (.B(net319),
    .C(net188),
    .A(net318),
    .Y(_0787_));
 sg13g2_nand2b_1 _1493_ (.Y(_0788_),
    .B(net280),
    .A_N(_0787_));
 sg13g2_o21ai_1 _1494_ (.B1(_0788_),
    .Y(_0789_),
    .A1(net188),
    .A2(_0786_));
 sg13g2_a21oi_1 _1495_ (.A1(_0733_),
    .A2(net257),
    .Y(_0063_),
    .B1(_0789_));
 sg13g2_o21ai_1 _1496_ (.B1(_0238_),
    .Y(_0790_),
    .A1(_0780_),
    .A2(_0787_));
 sg13g2_nor2_1 _1497_ (.A(_0238_),
    .B(_0787_),
    .Y(_0791_));
 sg13g2_a21oi_1 _1498_ (.A1(net280),
    .A2(_0791_),
    .Y(_0792_),
    .B1(net257));
 sg13g2_a22oi_1 _1499_ (.Y(_0793_),
    .B1(_0790_),
    .B2(_0792_),
    .A2(net257),
    .A1(_0737_));
 sg13g2_inv_1 _1500_ (.Y(_0064_),
    .A(_0793_));
 sg13g2_nor3_1 _1501_ (.A(_0238_),
    .B(_0240_),
    .C(_0787_),
    .Y(_0794_));
 sg13g2_a21oi_1 _1502_ (.A1(net280),
    .A2(_0794_),
    .Y(_0795_),
    .B1(net257));
 sg13g2_a21oi_1 _1503_ (.A1(_0741_),
    .A2(net257),
    .Y(_0796_),
    .B1(_0795_));
 sg13g2_a21oi_1 _1504_ (.A1(_0240_),
    .A2(_0792_),
    .Y(_0065_),
    .B1(_0796_));
 sg13g2_nand2_1 _1505_ (.Y(_0797_),
    .A(_0745_),
    .B(net257));
 sg13g2_nand3_1 _1506_ (.B(net280),
    .C(_0794_),
    .A(net317),
    .Y(_0798_));
 sg13g2_nand2_1 _1507_ (.Y(_0799_),
    .A(_0778_),
    .B(_0798_));
 sg13g2_a22oi_1 _1508_ (.Y(_0066_),
    .B1(_0797_),
    .B2(_0799_),
    .A2(_0795_),
    .A1(_0239_));
 sg13g2_nand3_1 _1509_ (.B(\cpu0.dr[6] ),
    .C(_0794_),
    .A(net317),
    .Y(_0800_));
 sg13g2_inv_1 _1510_ (.Y(_0801_),
    .A(_0800_));
 sg13g2_a21oi_2 _1511_ (.B1(net258),
    .Y(_0802_),
    .A2(_0801_),
    .A1(_0779_));
 sg13g2_a21oi_1 _1512_ (.A1(_0749_),
    .A2(net259),
    .Y(_0803_),
    .B1(_0802_));
 sg13g2_nor2_1 _1513_ (.A(net174),
    .B(_0799_),
    .Y(_0804_));
 sg13g2_nor2_1 _1514_ (.A(_0803_),
    .B(net175),
    .Y(_0067_));
 sg13g2_a21o_1 _1515_ (.A2(_0778_),
    .A1(_0241_),
    .B1(_0802_),
    .X(_0805_));
 sg13g2_a21oi_1 _1516_ (.A1(_0753_),
    .A2(net258),
    .Y(_0806_),
    .B1(_0805_));
 sg13g2_a21oi_1 _1517_ (.A1(_0241_),
    .A2(_0802_),
    .Y(_0068_),
    .B1(_0806_));
 sg13g2_nand2_1 _1518_ (.Y(_0807_),
    .A(_0757_),
    .B(net259));
 sg13g2_a21oi_1 _1519_ (.A1(net316),
    .A2(net315),
    .Y(_0118_),
    .B1(net258));
 sg13g2_nor2_1 _1520_ (.A(_0802_),
    .B(_0118_),
    .Y(_0119_));
 sg13g2_a22oi_1 _1521_ (.Y(_0069_),
    .B1(_0807_),
    .B2(_0119_),
    .A2(_0805_),
    .A1(_0243_));
 sg13g2_nand2_1 _1522_ (.Y(_0120_),
    .A(_0761_),
    .B(net258));
 sg13g2_nand3_1 _1523_ (.B(net146),
    .C(net315),
    .A(net316),
    .Y(_0121_));
 sg13g2_a21oi_1 _1524_ (.A1(_0778_),
    .A2(_0121_),
    .Y(_0122_),
    .B1(_0802_));
 sg13g2_nor2_1 _1525_ (.A(net146),
    .B(_0119_),
    .Y(_0123_));
 sg13g2_a21oi_1 _1526_ (.A1(_0120_),
    .A2(_0122_),
    .Y(_0070_),
    .B1(net147));
 sg13g2_nand2_1 _1527_ (.Y(_0124_),
    .A(_0765_),
    .B(net258));
 sg13g2_nand4_1 _1528_ (.B(net146),
    .C(net315),
    .A(net316),
    .Y(_0125_),
    .D(net143));
 sg13g2_a21oi_1 _1529_ (.A1(_0778_),
    .A2(_0125_),
    .Y(_0126_),
    .B1(_0802_));
 sg13g2_nor2_1 _1530_ (.A(net143),
    .B(_0122_),
    .Y(_0127_));
 sg13g2_a21oi_1 _1531_ (.A1(_0124_),
    .A2(_0126_),
    .Y(_0071_),
    .B1(net144));
 sg13g2_nor2_1 _1532_ (.A(net150),
    .B(_0126_),
    .Y(_0128_));
 sg13g2_nor3_1 _1533_ (.A(_0244_),
    .B(_0800_),
    .C(_0125_),
    .Y(_0129_));
 sg13g2_a221oi_1 _1534_ (.B2(_0129_),
    .C1(_0128_),
    .B1(_0779_),
    .A1(_0770_),
    .Y(_0072_),
    .A2(net258));
 sg13g2_a21oi_1 _1535_ (.A1(net133),
    .A2(_0129_),
    .Y(_0130_),
    .B1(net258));
 sg13g2_or2_1 _1536_ (.X(_0131_),
    .B(_0130_),
    .A(_0780_));
 sg13g2_nand2_1 _1537_ (.Y(_0132_),
    .A(net133),
    .B(_0131_));
 sg13g2_and2_1 _1538_ (.A(\boot_to_cpu[12] ),
    .B(net275),
    .X(_0133_));
 sg13g2_a22oi_1 _1539_ (.Y(_0134_),
    .B1(_0133_),
    .B2(net258),
    .A2(_0130_),
    .A1(_0129_));
 sg13g2_o21ai_1 _1540_ (.B1(_0132_),
    .Y(_0073_),
    .A1(_0780_),
    .A2(_0134_));
 sg13g2_nand2_1 _1541_ (.Y(_0135_),
    .A(\boot_to_cpu[13] ),
    .B(net274));
 sg13g2_and4_1 _1542_ (.A(net179),
    .B(net133),
    .C(_0779_),
    .D(_0129_),
    .X(_0136_));
 sg13g2_a221oi_1 _1543_ (.B2(net259),
    .C1(_0136_),
    .B1(_0135_),
    .A1(_0245_),
    .Y(_0074_),
    .A2(_0131_));
 sg13g2_nand2_1 _1544_ (.Y(_0137_),
    .A(\cpu0.dr[14] ),
    .B(_0136_));
 sg13g2_a21oi_1 _1545_ (.A1(net193),
    .A2(_0136_),
    .Y(_0138_),
    .B1(net259));
 sg13g2_o21ai_1 _1546_ (.B1(_0138_),
    .Y(_0139_),
    .A1(net193),
    .A2(_0136_));
 sg13g2_nand2_1 _1547_ (.Y(_0140_),
    .A(\boot_to_cpu[14] ),
    .B(net274));
 sg13g2_o21ai_1 _1548_ (.B1(_0139_),
    .Y(_0075_),
    .A1(_0778_),
    .A2(_0140_));
 sg13g2_and2_1 _1549_ (.A(\boot_to_cpu[15] ),
    .B(net274),
    .X(_0141_));
 sg13g2_a22oi_1 _1550_ (.Y(_0142_),
    .B1(_0141_),
    .B2(net259),
    .A2(_0138_),
    .A1(net92));
 sg13g2_o21ai_1 _1551_ (.B1(_0142_),
    .Y(_0076_),
    .A1(net92),
    .A2(_0137_));
 sg13g2_nand2_1 _1552_ (.Y(_0143_),
    .A(\addr_to_memio[5] ),
    .B(_0313_));
 sg13g2_nor3_2 _1553_ (.A(\addr_to_memio[6] ),
    .B(_0317_),
    .C(_0143_),
    .Y(_0144_));
 sg13g2_mux2_1 _1554_ (.A0(net176),
    .A1(\P0.uptime[0] ),
    .S(_0144_),
    .X(_0077_));
 sg13g2_mux2_1 _1555_ (.A0(net141),
    .A1(\P0.uptime[1] ),
    .S(_0144_),
    .X(_0078_));
 sg13g2_mux2_1 _1556_ (.A0(net115),
    .A1(\P0.uptime[2] ),
    .S(_0144_),
    .X(_0079_));
 sg13g2_nand2_2 _1557_ (.Y(_0145_),
    .A(net50),
    .B(_0311_));
 sg13g2_mux2_1 _1558_ (.A0(_0722_),
    .A1(net130),
    .S(net253),
    .X(_0080_));
 sg13g2_nor2_1 _1559_ (.A(_0728_),
    .B(net252),
    .Y(_0146_));
 sg13g2_a21oi_1 _1560_ (.A1(_0251_),
    .A2(net252),
    .Y(_0081_),
    .B1(_0146_));
 sg13g2_nor2_1 _1561_ (.A(_0732_),
    .B(net253),
    .Y(_0147_));
 sg13g2_a21oi_1 _1562_ (.A1(_0267_),
    .A2(net253),
    .Y(_0082_),
    .B1(_0147_));
 sg13g2_nor2_1 _1563_ (.A(_0737_),
    .B(net252),
    .Y(_0148_));
 sg13g2_a21oi_1 _1564_ (.A1(_0268_),
    .A2(net252),
    .Y(_0083_),
    .B1(_0148_));
 sg13g2_nor2_1 _1565_ (.A(_0741_),
    .B(net252),
    .Y(_0149_));
 sg13g2_a21oi_1 _1566_ (.A1(_0269_),
    .A2(net252),
    .Y(_0084_),
    .B1(_0149_));
 sg13g2_nor2_1 _1567_ (.A(_0745_),
    .B(net252),
    .Y(_0150_));
 sg13g2_a21oi_1 _1568_ (.A1(_0271_),
    .A2(net253),
    .Y(_0085_),
    .B1(_0150_));
 sg13g2_nor2_1 _1569_ (.A(_0749_),
    .B(net256),
    .Y(_0151_));
 sg13g2_a21oi_1 _1570_ (.A1(_0270_),
    .A2(net256),
    .Y(_0086_),
    .B1(_0151_));
 sg13g2_mux2_1 _1571_ (.A0(_0753_),
    .A1(net310),
    .S(net253),
    .X(_0087_));
 sg13g2_nor2_1 _1572_ (.A(_0757_),
    .B(net252),
    .Y(_0152_));
 sg13g2_a21oi_1 _1573_ (.A1(_0248_),
    .A2(net254),
    .Y(_0088_),
    .B1(_0152_));
 sg13g2_nor2_1 _1574_ (.A(_0761_),
    .B(net254),
    .Y(_0153_));
 sg13g2_a21oi_1 _1575_ (.A1(_0249_),
    .A2(net254),
    .Y(_0089_),
    .B1(_0153_));
 sg13g2_mux2_1 _1576_ (.A0(_0765_),
    .A1(net129),
    .S(net254),
    .X(_0090_));
 sg13g2_nand2_1 _1577_ (.Y(_0154_),
    .A(net77),
    .B(net256));
 sg13g2_o21ai_1 _1578_ (.B1(_0154_),
    .Y(_0091_),
    .A1(_0770_),
    .A2(net256));
 sg13g2_nor2_1 _1579_ (.A(_0133_),
    .B(net255),
    .Y(_0155_));
 sg13g2_a21oi_1 _1580_ (.A1(_0234_),
    .A2(net255),
    .Y(_0092_),
    .B1(_0155_));
 sg13g2_a21oi_1 _1581_ (.A1(\boot_to_cpu[13] ),
    .A2(net274),
    .Y(_0156_),
    .B1(net254));
 sg13g2_a21oi_1 _1582_ (.A1(_0236_),
    .A2(net254),
    .Y(_0093_),
    .B1(_0156_));
 sg13g2_nand2_1 _1583_ (.Y(_0157_),
    .A(net298),
    .B(net255));
 sg13g2_o21ai_1 _1584_ (.B1(_0157_),
    .Y(_0094_),
    .A1(_0140_),
    .A2(net254));
 sg13g2_nor2_1 _1585_ (.A(_0141_),
    .B(net255),
    .Y(_0158_));
 sg13g2_a21oi_1 _1586_ (.A1(_0233_),
    .A2(net254),
    .Y(_0095_),
    .B1(_0158_));
 sg13g2_a22oi_1 _1587_ (.Y(_0159_),
    .B1(\cpu0.ac[15] ),
    .B2(\cpu0.ir[3] ),
    .A2(\cpu0.ir[1] ),
    .A1(_0250_));
 sg13g2_or4_1 _1588_ (.A(\cpu0.ac[3] ),
    .B(\cpu0.ac[2] ),
    .C(net328),
    .D(net330),
    .X(_0160_));
 sg13g2_nor4_1 _1589_ (.A(net350),
    .B(net351),
    .C(\cpu0.ac[13] ),
    .D(\cpu0.ac[12] ),
    .Y(_0161_));
 sg13g2_nor2_1 _1590_ (.A(\cpu0.ac[15] ),
    .B(\cpu0.ac[14] ),
    .Y(_0162_));
 sg13g2_o21ai_1 _1591_ (.B1(_0159_),
    .Y(_0163_),
    .A1(\cpu0.ac[15] ),
    .A2(_0269_));
 sg13g2_nor4_1 _1592_ (.A(\cpu0.ac[7] ),
    .B(\cpu0.ac[6] ),
    .C(\cpu0.ac[9] ),
    .D(\cpu0.ac[8] ),
    .Y(_0164_));
 sg13g2_nand4_1 _1593_ (.B(_0161_),
    .C(_0162_),
    .A(\cpu0.ir[2] ),
    .Y(_0165_),
    .D(_0164_));
 sg13g2_nor3_1 _1594_ (.A(_0626_),
    .B(_0160_),
    .C(_0165_),
    .Y(_0166_));
 sg13g2_o21ai_1 _1595_ (.B1(_0407_),
    .Y(_0167_),
    .A1(_0163_),
    .A2(_0166_));
 sg13g2_a21oi_1 _1596_ (.A1(net297),
    .A2(\cpu0.t[9] ),
    .Y(_0168_),
    .B1(net292));
 sg13g2_nor2_1 _1597_ (.A(_0294_),
    .B(_0168_),
    .Y(_0169_));
 sg13g2_nor4_1 _1598_ (.A(\cpu0.dr[5] ),
    .B(\cpu0.dr[4] ),
    .C(net316),
    .D(\cpu0.dr[6] ),
    .Y(_0170_));
 sg13g2_nor4_1 _1599_ (.A(net318),
    .B(\cpu0.dr[0] ),
    .C(\cpu0.dr[3] ),
    .D(\cpu0.dr[2] ),
    .Y(_0171_));
 sg13g2_nor4_1 _1600_ (.A(\cpu0.dr[13] ),
    .B(\cpu0.dr[12] ),
    .C(\cpu0.dr[15] ),
    .D(\cpu0.dr[14] ),
    .Y(_0172_));
 sg13g2_nor4_1 _1601_ (.A(\cpu0.dr[9] ),
    .B(net315),
    .C(\cpu0.dr[11] ),
    .D(\cpu0.dr[10] ),
    .Y(_0173_));
 sg13g2_and4_1 _1602_ (.A(_0170_),
    .B(_0171_),
    .C(_0172_),
    .D(_0173_),
    .X(_0174_));
 sg13g2_a221oi_1 _1603_ (.B2(_0174_),
    .C1(net348),
    .B1(_0169_),
    .A1(\cpu0.t[6] ),
    .Y(_0175_),
    .A2(_0297_));
 sg13g2_a22oi_1 _1604_ (.Y(_0176_),
    .B1(net10),
    .B2(net299),
    .A2(\cpu0.ir[8] ),
    .A1(\cpu0.ir[10] ));
 sg13g2_nand2b_1 _1605_ (.Y(_0177_),
    .B(_0303_),
    .A_N(_0176_));
 sg13g2_nand3_1 _1606_ (.B(_0175_),
    .C(_0177_),
    .A(_0167_),
    .Y(_0178_));
 sg13g2_inv_4 _1607_ (.A(net277),
    .Y(_0179_));
 sg13g2_or2_1 _1608_ (.X(_0180_),
    .B(net293),
    .A(net338));
 sg13g2_a22oi_1 _1609_ (.Y(_0181_),
    .B1(_0399_),
    .B2(_0180_),
    .A2(_0297_),
    .A1(net78));
 sg13g2_nor2b_2 _1610_ (.A(net277),
    .B_N(_0181_),
    .Y(_0182_));
 sg13g2_inv_1 _1611_ (.Y(_0183_),
    .A(_0182_));
 sg13g2_nor2_1 _1612_ (.A(net277),
    .B(_0181_),
    .Y(_0184_));
 sg13g2_nor2_1 _1613_ (.A(net161),
    .B(_0179_),
    .Y(_0185_));
 sg13g2_a221oi_1 _1614_ (.B2(net108),
    .C1(_0185_),
    .B1(net268),
    .A1(net161),
    .Y(_0186_),
    .A2(_0182_));
 sg13g2_inv_1 _1615_ (.Y(_0096_),
    .A(_0186_));
 sg13g2_xnor2_1 _1616_ (.Y(_0187_),
    .A(net161),
    .B(net171));
 sg13g2_a22oi_1 _1617_ (.Y(_0188_),
    .B1(net268),
    .B2(net158),
    .A2(_0182_),
    .A1(net171));
 sg13g2_o21ai_1 _1618_ (.B1(_0188_),
    .Y(_0097_),
    .A1(_0179_),
    .A2(_0187_));
 sg13g2_nand3_1 _1619_ (.B(\cpu0.pc[1] ),
    .C(net168),
    .A(net161),
    .Y(_0189_));
 sg13g2_a21o_1 _1620_ (.A2(\cpu0.pc[1] ),
    .A1(\cpu0.pc[0] ),
    .B1(\cpu0.pc[2] ),
    .X(_0190_));
 sg13g2_nand2_1 _1621_ (.Y(_0191_),
    .A(_0189_),
    .B(_0190_));
 sg13g2_a22oi_1 _1622_ (.Y(_0192_),
    .B1(net268),
    .B2(net155),
    .A2(_0182_),
    .A1(\cpu0.pc[2] ));
 sg13g2_o21ai_1 _1623_ (.B1(net156),
    .Y(_0098_),
    .A1(_0179_),
    .A2(_0191_));
 sg13g2_nor2_1 _1624_ (.A(_0279_),
    .B(_0189_),
    .Y(_0193_));
 sg13g2_xnor2_1 _1625_ (.Y(_0194_),
    .A(_0279_),
    .B(_0189_));
 sg13g2_a22oi_1 _1626_ (.Y(_0195_),
    .B1(net268),
    .B2(net169),
    .A2(_0182_),
    .A1(net164));
 sg13g2_o21ai_1 _1627_ (.B1(_0195_),
    .Y(_0099_),
    .A1(_0179_),
    .A2(_0194_));
 sg13g2_and2_1 _1628_ (.A(\cpu0.pc[4] ),
    .B(_0193_),
    .X(_0196_));
 sg13g2_xnor2_1 _1629_ (.Y(_0197_),
    .A(\cpu0.pc[4] ),
    .B(_0193_));
 sg13g2_a22oi_1 _1630_ (.Y(_0198_),
    .B1(net268),
    .B2(net126),
    .A2(_0182_),
    .A1(\cpu0.pc[4] ));
 sg13g2_o21ai_1 _1631_ (.B1(net127),
    .Y(_0100_),
    .A1(_0179_),
    .A2(_0197_));
 sg13g2_nand2_1 _1632_ (.Y(_0199_),
    .A(net98),
    .B(_0179_));
 sg13g2_and2_1 _1633_ (.A(net142),
    .B(_0196_),
    .X(_0200_));
 sg13g2_a21oi_1 _1634_ (.A1(net277),
    .A2(_0200_),
    .Y(_0201_),
    .B1(net268));
 sg13g2_o21ai_1 _1635_ (.B1(_0201_),
    .Y(_0202_),
    .A1(\cpu0.pc[5] ),
    .A2(_0196_));
 sg13g2_a22oi_1 _1636_ (.Y(_0101_),
    .B1(_0199_),
    .B2(_0202_),
    .A2(_0182_),
    .A1(_0282_));
 sg13g2_and3_1 _1637_ (.X(_0203_),
    .A(net131),
    .B(net277),
    .C(_0200_));
 sg13g2_a221oi_1 _1638_ (.B2(_0284_),
    .C1(_0203_),
    .B1(_0201_),
    .A1(_0285_),
    .Y(_0102_),
    .A2(net268));
 sg13g2_nor3_1 _1639_ (.A(net178),
    .B(net268),
    .C(_0203_),
    .Y(_0204_));
 sg13g2_nor3_1 _1640_ (.A(net119),
    .B(net277),
    .C(_0181_),
    .Y(_0205_));
 sg13g2_and4_1 _1641_ (.A(net131),
    .B(net178),
    .C(net277),
    .D(_0200_),
    .X(_0206_));
 sg13g2_nor3_1 _1642_ (.A(_0204_),
    .B(_0205_),
    .C(_0206_),
    .Y(_0103_));
 sg13g2_nor3_1 _1643_ (.A(net180),
    .B(net269),
    .C(_0206_),
    .Y(_0207_));
 sg13g2_nor3_1 _1644_ (.A(net104),
    .B(net277),
    .C(_0181_),
    .Y(_0208_));
 sg13g2_and2_1 _1645_ (.A(net180),
    .B(_0206_),
    .X(_0209_));
 sg13g2_nor3_1 _1646_ (.A(_0207_),
    .B(_0208_),
    .C(_0209_),
    .Y(_0104_));
 sg13g2_nor3_1 _1647_ (.A(net81),
    .B(net269),
    .C(_0209_),
    .Y(_0210_));
 sg13g2_nand2_1 _1648_ (.Y(_0211_),
    .A(net81),
    .B(_0209_));
 sg13g2_a221oi_1 _1649_ (.B2(net81),
    .C1(_0210_),
    .B1(_0209_),
    .A1(_0274_),
    .Y(_0105_),
    .A2(net269));
 sg13g2_nand3_1 _1650_ (.B(net110),
    .C(_0209_),
    .A(net81),
    .Y(_0212_));
 sg13g2_nand2b_1 _1651_ (.Y(_0213_),
    .B(_0212_),
    .A_N(net269));
 sg13g2_nand2_1 _1652_ (.Y(_0214_),
    .A(net84),
    .B(_0179_));
 sg13g2_nor2_1 _1653_ (.A(net110),
    .B(net269),
    .Y(_0215_));
 sg13g2_a22oi_1 _1654_ (.Y(_0106_),
    .B1(_0215_),
    .B2(_0211_),
    .A2(_0214_),
    .A1(_0213_));
 sg13g2_nand4_1 _1655_ (.B(\cpu0.pc[10] ),
    .C(net101),
    .A(net81),
    .Y(_0216_),
    .D(_0209_));
 sg13g2_o21ai_1 _1656_ (.B1(_0216_),
    .Y(_0217_),
    .A1(\addr_to_memio[11] ),
    .A2(_0178_));
 sg13g2_nor2_1 _1657_ (.A(net101),
    .B(_0213_),
    .Y(_0218_));
 sg13g2_a21oi_1 _1658_ (.A1(_0183_),
    .A2(_0217_),
    .Y(_0107_),
    .B1(net102));
 sg13g2_nand2b_1 _1659_ (.Y(_0219_),
    .B(net361),
    .A_N(net112));
 sg13g2_a21oi_1 _1660_ (.A1(net117),
    .A2(net267),
    .Y(_0108_),
    .B1(_0219_));
 sg13g2_nand2_1 _1661_ (.Y(_0220_),
    .A(net59),
    .B(net112));
 sg13g2_nand2_1 _1662_ (.Y(_0221_),
    .A(net361),
    .B(_0220_));
 sg13g2_and2_1 _1663_ (.A(net116),
    .B(net112),
    .X(_0222_));
 sg13g2_nor3_1 _1664_ (.A(net113),
    .B(_0221_),
    .C(_0222_),
    .Y(_0109_));
 sg13g2_xnor2_1 _1665_ (.Y(_0223_),
    .A(net125),
    .B(_0222_));
 sg13g2_nor2_1 _1666_ (.A(_0221_),
    .B(_0223_),
    .Y(_0110_));
 sg13g2_a21oi_1 _1667_ (.A1(\spi0.cntreg[2] ),
    .A2(_0222_),
    .Y(_0224_),
    .B1(net59));
 sg13g2_nor2_1 _1668_ (.A(_0221_),
    .B(net60),
    .Y(_0111_));
 sg13g2_nand3b_1 _1669_ (.B(_0313_),
    .C(\addr_to_memio[6] ),
    .Y(_0225_),
    .A_N(_0317_));
 sg13g2_mux2_1 _1670_ (.A0(\P0.uptime[0] ),
    .A1(net47),
    .S(_0225_),
    .X(_0112_));
 sg13g2_mux2_1 _1671_ (.A0(\P0.uptime[1] ),
    .A1(net70),
    .S(_0225_),
    .X(_0113_));
 sg13g2_mux2_1 _1672_ (.A0(\P0.uptime[2] ),
    .A1(net65),
    .S(_0225_),
    .X(_0114_));
 sg13g2_nor3_2 _1673_ (.A(net39),
    .B(net43),
    .C(net56),
    .Y(_0226_));
 sg13g2_or2_1 _1674_ (.X(_0227_),
    .B(_0226_),
    .A(_0304_));
 sg13g2_nand2_1 _1675_ (.Y(_0228_),
    .A(net47),
    .B(_0226_));
 sg13g2_o21ai_1 _1676_ (.B1(net48),
    .Y(_0115_),
    .A1(\P0.uptimereg[0] ),
    .A2(_0227_));
 sg13g2_xor2_1 _1677_ (.B(\P0.uptimereg[0] ),
    .A(\P0.uptimereg[1] ),
    .X(_0229_));
 sg13g2_nand2_1 _1678_ (.Y(_0230_),
    .A(net70),
    .B(_0226_));
 sg13g2_o21ai_1 _1679_ (.B1(_0230_),
    .Y(_0116_),
    .A1(_0227_),
    .A2(_0229_));
 sg13g2_nand2_1 _1680_ (.Y(_0231_),
    .A(net65),
    .B(_0226_));
 sg13g2_o21ai_1 _1681_ (.B1(\P0.uptimereg[2] ),
    .Y(_0232_),
    .A1(\P0.uptimereg[1] ),
    .A2(\P0.uptimereg[0] ));
 sg13g2_o21ai_1 _1682_ (.B1(_0231_),
    .Y(_0117_),
    .A1(_0226_),
    .A2(_0232_));
 sg13g2_o21ai_1 _1683_ (.B1(net290),
    .Y(_0809_),
    .A1(net293),
    .A2(net292));
 sg13g2_o21ai_1 _1684_ (.B1(net290),
    .Y(_0810_),
    .A1(net293),
    .A2(net292));
 sg13g2_o21ai_1 _1685_ (.B1(net290),
    .Y(_0811_),
    .A1(net293),
    .A2(net292));
 sg13g2_o21ai_1 _1686_ (.B1(net290),
    .Y(_0812_),
    .A1(net293),
    .A2(net292));
 sg13g2_o21ai_1 _1687_ (.B1(net290),
    .Y(_0813_),
    .A1(_0289_),
    .A2(net292));
 sg13g2_o21ai_1 _1688_ (.B1(_0293_),
    .Y(_0814_),
    .A1(_0289_),
    .A2(_0295_));
 sg13g2_o21ai_1 _1689_ (.B1(_0293_),
    .Y(_0815_),
    .A1(_0289_),
    .A2(_0295_));
 sg13g2_nand2b_2 _1690_ (.Y(_0817_),
    .B(net291),
    .A_N(_0290_));
 sg13g2_nand2b_2 _1691_ (.Y(_0818_),
    .B(net291),
    .A_N(_0290_));
 sg13g2_nand2b_2 _1692_ (.Y(_0819_),
    .B(net291),
    .A_N(_0290_));
 sg13g2_nand2b_2 _1693_ (.Y(_0820_),
    .B(net291),
    .A_N(_0290_));
 sg13g2_nand2b_2 _1694_ (.Y(_0821_),
    .B(net291),
    .A_N(_0290_));
 sg13g2_nand2b_2 _1695_ (.Y(_0822_),
    .B(_0288_),
    .A_N(_0290_));
 sg13g2_nand2b_2 _1696_ (.Y(_0823_),
    .B(_0288_),
    .A_N(_0290_));
 sg13g2_nand2_2 _1697_ (.Y(_0826_),
    .A(net337),
    .B(net285));
 sg13g2_nand2_2 _1698_ (.Y(_0827_),
    .A(net337),
    .B(net285));
 sg13g2_nand2_2 _1699_ (.Y(_0828_),
    .A(net337),
    .B(net285));
 sg13g2_nand2_2 _1700_ (.Y(_0829_),
    .A(net337),
    .B(net285));
 sg13g2_nand2_2 _1701_ (.Y(_0830_),
    .A(net337),
    .B(net285));
 sg13g2_nand2_2 _1702_ (.Y(_0831_),
    .A(net337),
    .B(net285));
 sg13g2_nand2_2 _1703_ (.Y(_0824_),
    .A(net337),
    .B(net285));
 sg13g2_dfrbpq_1 _1704_ (.RESET_B(net1),
    .D(net17),
    .Q(rst_n_i),
    .CLK(clknet_3_7__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1705_ (.RESET_B(net366),
    .D(_0020_),
    .Q(\cpu0.ac[8] ),
    .CLK(\clknet_4_14_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1706_ (.RESET_B(net366),
    .D(net167),
    .Q(\cpu0.ac[9] ),
    .CLK(\clknet_4_14_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1707_ (.RESET_B(net366),
    .D(net198),
    .Q(\cpu0.ac[10] ),
    .CLK(\clknet_4_14_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1708_ (.RESET_B(net366),
    .D(net203),
    .Q(\cpu0.ac[11] ),
    .CLK(\clknet_4_14_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1709_ (.RESET_B(net366),
    .D(_0024_),
    .Q(\cpu0.ac[12] ),
    .CLK(\clknet_4_14_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1710_ (.RESET_B(net366),
    .D(net163),
    .Q(\cpu0.ac[13] ),
    .CLK(\clknet_4_11_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1711_ (.RESET_B(net363),
    .D(net183),
    .Q(\cpu0.ac[14] ),
    .CLK(\clknet_4_11_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1712_ (.RESET_B(net363),
    .D(_0027_),
    .Q(\cpu0.ac[15] ),
    .CLK(\clknet_4_11_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1713_ (.RESET_B(net28),
    .D(\cpu0.rstT ),
    .Q(\cpu0.t[0] ),
    .CLK(\clknet_4_6_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1714_ (.RESET_B(net27),
    .D(_0028_),
    .Q(\cpu0.t[1] ),
    .CLK(\clknet_4_9_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1715_ (.RESET_B(net26),
    .D(net41),
    .Q(\cpu0.t[2] ),
    .CLK(\clknet_4_8_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1716_ (.RESET_B(net25),
    .D(net51),
    .Q(\cpu0.t[3] ),
    .CLK(\clknet_4_8_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1717_ (.RESET_B(net24),
    .D(_0031_),
    .Q(\cpu0.t[4] ),
    .CLK(\clknet_4_10_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1718_ (.RESET_B(net23),
    .D(net186),
    .Q(\cpu0.t[5] ),
    .CLK(\clknet_4_9_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1719_ (.RESET_B(net22),
    .D(_0033_),
    .Q(\cpu0.t[6] ),
    .CLK(\clknet_4_8_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1720_ (.RESET_B(net21),
    .D(net89),
    .Q(\cpu0.t[7] ),
    .CLK(\clknet_4_8_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1721_ (.RESET_B(net20),
    .D(net73),
    .Q(\cpu0.t[8] ),
    .CLK(\clknet_4_8_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1722_ (.RESET_B(net19),
    .D(net55),
    .Q(\cpu0.t[9] ),
    .CLK(\clknet_4_10_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1723_ (.RESET_B(net18),
    .D(net75),
    .Q(\cpu0.t[10] ),
    .CLK(\clknet_4_8_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1724_ (.RESET_B(net363),
    .D(net95),
    .Q(\cpu0.ac0 ),
    .CLK(\clknet_4_10_0_cpu0.clk ));
 sg13g2_dlhq_1 _1725_ (.D(net336),
    .GATE(net279),
    .Q(uo_out[0]));
 sg13g2_dlhq_1 _1726_ (.D(net333),
    .GATE(net279),
    .Q(uo_out[1]));
 sg13g2_dlhq_1 _1727_ (.D(net332),
    .GATE(net279),
    .Q(uo_out[2]));
 sg13g2_dlhq_1 _1728_ (.D(net331),
    .GATE(net279),
    .Q(uo_out[3]));
 sg13g2_dlhq_1 _1729_ (.D(net329),
    .GATE(\cpu0.en_out ),
    .Q(uo_out[4]));
 sg13g2_dlhq_1 _1730_ (.D(net327),
    .GATE(net279),
    .Q(uo_out[5]));
 sg13g2_dlhq_1 _1731_ (.D(net326),
    .GATE(net279),
    .Q(uo_out[6]));
 sg13g2_dlhq_1 _1732_ (.D(net325),
    .GATE(net279),
    .Q(uo_out[7]));
 sg13g2_dfrbpq_1 _1733_ (.RESET_B(net363),
    .D(_0039_),
    .Q(\cpu0.ac[0] ),
    .CLK(\clknet_4_12_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1734_ (.RESET_B(net365),
    .D(net213),
    .Q(\cpu0.ac[1] ),
    .CLK(\clknet_4_13_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1735_ (.RESET_B(net367),
    .D(_0041_),
    .Q(\cpu0.ac[2] ),
    .CLK(\clknet_4_15_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1736_ (.RESET_B(net365),
    .D(_0042_),
    .Q(\cpu0.ac[3] ),
    .CLK(\clknet_4_13_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1737_ (.RESET_B(net368),
    .D(net192),
    .Q(\cpu0.ac[4] ),
    .CLK(\clknet_4_15_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1738_ (.RESET_B(net367),
    .D(net205),
    .Q(\cpu0.ac[5] ),
    .CLK(\clknet_4_15_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1739_ (.RESET_B(net367),
    .D(net211),
    .Q(\cpu0.ac[6] ),
    .CLK(\clknet_4_15_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1740_ (.RESET_B(net367),
    .D(net215),
    .Q(\cpu0.ac[7] ),
    .CLK(\clknet_4_15_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1741_ (.RESET_B(net364),
    .D(net136),
    .Q(\cpu0.e ),
    .CLK(\clknet_4_11_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1742_ (.RESET_B(net352),
    .D(net109),
    .Q(\addr_to_memio[0] ),
    .CLK(\clknet_4_1_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1743_ (.RESET_B(net355),
    .D(net159),
    .Q(\addr_to_memio[1] ),
    .CLK(\clknet_4_1_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1744_ (.RESET_B(net352),
    .D(_0050_),
    .Q(\addr_to_memio[2] ),
    .CLK(\clknet_4_1_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1745_ (.RESET_B(net352),
    .D(net165),
    .Q(\addr_to_memio[3] ),
    .CLK(\clknet_4_1_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1746_ (.RESET_B(net352),
    .D(net140),
    .Q(\addr_to_memio[4] ),
    .CLK(\clknet_4_1_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1747_ (.RESET_B(net353),
    .D(_0053_),
    .Q(\addr_to_memio[5] ),
    .CLK(\clknet_4_2_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1748_ (.RESET_B(net355),
    .D(_0054_),
    .Q(\addr_to_memio[6] ),
    .CLK(\clknet_4_0_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1749_ (.RESET_B(net353),
    .D(net120),
    .Q(\addr_to_memio[7] ),
    .CLK(\clknet_4_3_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1750_ (.RESET_B(net362),
    .D(net105),
    .Q(\addr_to_memio[8] ),
    .CLK(\clknet_4_6_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1751_ (.RESET_B(net362),
    .D(net122),
    .Q(\addr_to_memio[9] ),
    .CLK(\clknet_4_6_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1752_ (.RESET_B(net353),
    .D(net85),
    .Q(\addr_to_memio[10] ),
    .CLK(\clknet_4_2_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1753_ (.RESET_B(net353),
    .D(net124),
    .Q(\addr_to_memio[11] ),
    .CLK(\clknet_4_3_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1754_ (.RESET_B(net363),
    .D(net64),
    .Q(\cpu0.ac15 ),
    .CLK(\clknet_4_10_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1755_ (.RESET_B(net360),
    .D(_0061_),
    .Q(\cpu0.dr[0] ),
    .CLK(\clknet_4_4_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1756_ (.RESET_B(net360),
    .D(_0062_),
    .Q(\cpu0.dr[1] ),
    .CLK(\clknet_4_4_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1757_ (.RESET_B(net360),
    .D(_0063_),
    .Q(\cpu0.dr[2] ),
    .CLK(\clknet_4_5_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1758_ (.RESET_B(net360),
    .D(_0064_),
    .Q(\cpu0.dr[3] ),
    .CLK(\clknet_4_5_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1759_ (.RESET_B(net360),
    .D(net154),
    .Q(\cpu0.dr[4] ),
    .CLK(\clknet_4_5_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1760_ (.RESET_B(net359),
    .D(_0066_),
    .Q(\cpu0.dr[5] ),
    .CLK(\clknet_4_5_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1761_ (.RESET_B(net359),
    .D(_0067_),
    .Q(\cpu0.dr[6] ),
    .CLK(\clknet_4_5_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1762_ (.RESET_B(net365),
    .D(_0068_),
    .Q(\cpu0.dr[7] ),
    .CLK(\clknet_4_13_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1763_ (.RESET_B(net365),
    .D(net201),
    .Q(\cpu0.dr[8] ),
    .CLK(\clknet_4_13_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1764_ (.RESET_B(net365),
    .D(net148),
    .Q(\cpu0.dr[9] ),
    .CLK(\clknet_4_13_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1765_ (.RESET_B(net365),
    .D(net145),
    .Q(\cpu0.dr[10] ),
    .CLK(\clknet_4_12_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1766_ (.RESET_B(net365),
    .D(net151),
    .Q(\cpu0.dr[11] ),
    .CLK(\clknet_4_12_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1767_ (.RESET_B(net365),
    .D(net134),
    .Q(\cpu0.dr[12] ),
    .CLK(\clknet_4_12_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1768_ (.RESET_B(net366),
    .D(_0074_),
    .Q(\cpu0.dr[13] ),
    .CLK(\clknet_4_12_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1769_ (.RESET_B(net362),
    .D(_0075_),
    .Q(\cpu0.dr[14] ),
    .CLK(\clknet_4_4_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1770_ (.RESET_B(net364),
    .D(net93),
    .Q(\cpu0.dr[15] ),
    .CLK(\clknet_4_7_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1771_ (.RESET_B(net357),
    .D(_0077_),
    .Q(\T0.selreg[0] ),
    .CLK(clknet_3_3__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1772_ (.RESET_B(net356),
    .D(_0078_),
    .Q(\T0.selreg[1] ),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1773_ (.RESET_B(net356),
    .D(_0079_),
    .Q(\T0.selreg[2] ),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1774_ (.RESET_B(net354),
    .D(_0080_),
    .Q(\cpu0.ir[0] ),
    .CLK(\clknet_4_4_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1775_ (.RESET_B(net354),
    .D(_0081_),
    .Q(\cpu0.ir[1] ),
    .CLK(\clknet_4_3_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1776_ (.RESET_B(net360),
    .D(_0082_),
    .Q(\cpu0.ir[2] ),
    .CLK(\clknet_4_4_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1777_ (.RESET_B(net354),
    .D(_0083_),
    .Q(\cpu0.ir[3] ),
    .CLK(\clknet_4_7_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1778_ (.RESET_B(net354),
    .D(_0084_),
    .Q(\cpu0.ir[4] ),
    .CLK(\clknet_4_3_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1779_ (.RESET_B(net355),
    .D(_0085_),
    .Q(\cpu0.ir[5] ),
    .CLK(\clknet_4_7_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1780_ (.RESET_B(net366),
    .D(_0086_),
    .Q(\cpu0.ir[6] ),
    .CLK(\clknet_4_12_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1781_ (.RESET_B(net354),
    .D(_0087_),
    .Q(\cpu0.ir[7] ),
    .CLK(\clknet_4_4_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1782_ (.RESET_B(net364),
    .D(_0088_),
    .Q(\cpu0.ir[8] ),
    .CLK(\clknet_4_7_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1783_ (.RESET_B(net363),
    .D(_0089_),
    .Q(\cpu0.ir[9] ),
    .CLK(\clknet_4_10_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1784_ (.RESET_B(net362),
    .D(_0090_),
    .Q(\cpu0.ir[10] ),
    .CLK(\clknet_4_7_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1785_ (.RESET_B(net362),
    .D(_0091_),
    .Q(\cpu0.ir[11] ),
    .CLK(\clknet_4_11_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1786_ (.RESET_B(net362),
    .D(_0092_),
    .Q(\cpu0.decode2.a[0] ),
    .CLK(\clknet_4_9_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1787_ (.RESET_B(net364),
    .D(_0093_),
    .Q(\cpu0.decode2.a[1] ),
    .CLK(\clknet_4_9_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1788_ (.RESET_B(net362),
    .D(_0094_),
    .Q(\cpu0.decode2.a[2] ),
    .CLK(\clknet_4_9_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1789_ (.RESET_B(net363),
    .D(_0095_),
    .Q(\cpu0.ir[15] ),
    .CLK(\clknet_4_10_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1790_ (.RESET_B(net352),
    .D(_0096_),
    .Q(\cpu0.pc[0] ),
    .CLK(\clknet_4_0_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1791_ (.RESET_B(net352),
    .D(_0097_),
    .Q(\cpu0.pc[1] ),
    .CLK(\clknet_4_0_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1792_ (.RESET_B(net355),
    .D(net157),
    .Q(\cpu0.pc[2] ),
    .CLK(\clknet_4_0_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1793_ (.RESET_B(net352),
    .D(net170),
    .Q(\cpu0.pc[3] ),
    .CLK(\clknet_4_0_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1794_ (.RESET_B(net352),
    .D(net128),
    .Q(\cpu0.pc[4] ),
    .CLK(\clknet_4_2_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1795_ (.RESET_B(net353),
    .D(net99),
    .Q(\cpu0.pc[5] ),
    .CLK(\clknet_4_2_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1796_ (.RESET_B(net353),
    .D(_0102_),
    .Q(\cpu0.pc[6] ),
    .CLK(\clknet_4_0_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1797_ (.RESET_B(net353),
    .D(_0103_),
    .Q(\cpu0.pc[7] ),
    .CLK(\clknet_4_2_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1798_ (.RESET_B(net354),
    .D(_0104_),
    .Q(\cpu0.pc[8] ),
    .CLK(\clknet_4_6_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1799_ (.RESET_B(net362),
    .D(net82),
    .Q(\cpu0.pc[9] ),
    .CLK(\clknet_4_6_0_cpu0.clk ));
 sg13g2_dfrbpq_2 _1800_ (.RESET_B(net354),
    .D(net111),
    .Q(\cpu0.pc[10] ),
    .CLK(\clknet_4_3_0_cpu0.clk ));
 sg13g2_dfrbpq_1 _1801_ (.RESET_B(net353),
    .D(net103),
    .Q(\cpu0.pc[11] ),
    .CLK(\clknet_4_2_0_cpu0.clk ));
 sg13g2_dlhq_1 _1802_ (.D(\mem0.dout_internal[0] ),
    .GATE(net266),
    .Q(\boot_to_cpu[0] ));
 sg13g2_dlhq_1 _1803_ (.D(\mem0.dout_internal[1] ),
    .GATE(net266),
    .Q(\boot_to_cpu[1] ));
 sg13g2_dlhq_1 _1804_ (.D(\mem0.dout_internal[2] ),
    .GATE(net266),
    .Q(\boot_to_cpu[2] ));
 sg13g2_dlhq_1 _1805_ (.D(\mem0.dout_internal[3] ),
    .GATE(net266),
    .Q(\boot_to_cpu[3] ));
 sg13g2_dlhq_1 _1806_ (.D(\mem0.dout_internal[4] ),
    .GATE(net266),
    .Q(\boot_to_cpu[4] ));
 sg13g2_dlhq_1 _1807_ (.D(\mem0.dout_internal[5] ),
    .GATE(_0000_),
    .Q(\boot_to_cpu[5] ));
 sg13g2_dlhq_1 _1808_ (.D(\mem0.dout_internal[6] ),
    .GATE(net266),
    .Q(\boot_to_cpu[6] ));
 sg13g2_dlhq_1 _1809_ (.D(\mem0.dout_internal[7] ),
    .GATE(net266),
    .Q(\boot_to_cpu[7] ));
 sg13g2_dlhq_1 _1810_ (.D(\mem0.dout_internal[8] ),
    .GATE(net265),
    .Q(\boot_to_cpu[8] ));
 sg13g2_dlhq_1 _1811_ (.D(\mem0.dout_internal[9] ),
    .GATE(net265),
    .Q(\boot_to_cpu[9] ));
 sg13g2_dlhq_1 _1812_ (.D(\mem0.dout_internal[10] ),
    .GATE(net265),
    .Q(\boot_to_cpu[10] ));
 sg13g2_dlhq_1 _1813_ (.D(\mem0.dout_internal[11] ),
    .GATE(net265),
    .Q(\boot_to_cpu[11] ));
 sg13g2_dlhq_1 _1814_ (.D(\mem0.dout_internal[12] ),
    .GATE(net265),
    .Q(\boot_to_cpu[12] ));
 sg13g2_dlhq_1 _1815_ (.D(\mem0.dout_internal[13] ),
    .GATE(net265),
    .Q(\boot_to_cpu[13] ));
 sg13g2_dlhq_1 _1816_ (.D(\mem0.dout_internal[14] ),
    .GATE(net265),
    .Q(\boot_to_cpu[14] ));
 sg13g2_dlhq_1 _1817_ (.D(\mem0.dout_internal[15] ),
    .GATE(net265),
    .Q(\boot_to_cpu[15] ));
 sg13g2_dfrbpq_2 _1818_ (.RESET_B(net31),
    .D(_0108_),
    .Q(\spi0.cntreg[0] ),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1819_ (.RESET_B(net30),
    .D(net114),
    .Q(\spi0.cntreg[1] ),
    .CLK(clknet_3_7__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1820_ (.RESET_B(net29),
    .D(_0110_),
    .Q(\spi0.cntreg[2] ),
    .CLK(clknet_3_7__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1821_ (.RESET_B(net32),
    .D(net61),
    .Q(\spi0.cntreg[3] ),
    .CLK(clknet_3_7__leaf_clk_regs));
 sg13g2_dlhq_1 _1822_ (.D(\spi0.datareg[0] ),
    .GATE(\spi0.unload ),
    .Q(\spi0.dataout[0] ));
 sg13g2_dlhq_1 _1823_ (.D(\spi0.datareg[1] ),
    .GATE(\spi0.unload ),
    .Q(\spi0.dataout[1] ));
 sg13g2_dlhq_1 _1824_ (.D(\spi0.datareg[2] ),
    .GATE(\spi0.unload ),
    .Q(\spi0.dataout[2] ));
 sg13g2_dlhq_1 _1825_ (.D(\spi0.datareg[3] ),
    .GATE(\spi0.unload ),
    .Q(\spi0.dataout[3] ));
 sg13g2_dlhq_1 _1826_ (.D(\spi0.datareg[4] ),
    .GATE(\spi0.unload ),
    .Q(\spi0.dataout[4] ));
 sg13g2_dlhq_1 _1827_ (.D(\spi0.datareg[5] ),
    .GATE(\spi0.unload ),
    .Q(\spi0.dataout[5] ));
 sg13g2_dlhq_1 _1828_ (.D(\spi0.datareg[6] ),
    .GATE(\spi0.unload ),
    .Q(\spi0.dataout[6] ));
 sg13g2_dlhq_1 _1829_ (.D(\spi0.datareg[7] ),
    .GATE(\spi0.unload ),
    .Q(\spi0.dataout[7] ));
 sg13g2_dfrbpq_1 _1830_ (.RESET_B(net359),
    .D(_0001_),
    .Q(\spi0.datareg[0] ),
    .CLK(clknet_3_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1831_ (.RESET_B(net358),
    .D(_0002_),
    .Q(\spi0.datareg[1] ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1832_ (.RESET_B(net358),
    .D(_0003_),
    .Q(\spi0.datareg[2] ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1833_ (.RESET_B(net358),
    .D(_0004_),
    .Q(\spi0.datareg[3] ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1834_ (.RESET_B(net358),
    .D(_0005_),
    .Q(\spi0.datareg[4] ),
    .CLK(clknet_3_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1835_ (.RESET_B(net358),
    .D(_0006_),
    .Q(\spi0.datareg[5] ),
    .CLK(clknet_3_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1836_ (.RESET_B(net358),
    .D(_0007_),
    .Q(\spi0.datareg[6] ),
    .CLK(clknet_3_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1837_ (.RESET_B(net360),
    .D(_0008_),
    .Q(\spi0.datareg[7] ),
    .CLK(clknet_3_1__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1838_ (.RESET_B(net357),
    .D(_0012_),
    .Q(\T0.count[0] ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1839_ (.RESET_B(net357),
    .D(_0013_),
    .Q(\T0.count[1] ),
    .CLK(clknet_3_5__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1840_ (.RESET_B(net356),
    .D(_0014_),
    .Q(\T0.count[2] ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1841_ (.RESET_B(net356),
    .D(net68),
    .Q(\T0.count[3] ),
    .CLK(clknet_3_5__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1842_ (.RESET_B(net357),
    .D(net53),
    .Q(\T0.count[4] ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1843_ (.RESET_B(net357),
    .D(net58),
    .Q(\T0.count[5] ),
    .CLK(clknet_3_5__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1844_ (.RESET_B(net357),
    .D(_0018_),
    .Q(\T0.count[6] ),
    .CLK(clknet_3_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1845_ (.RESET_B(net356),
    .D(net46),
    .Q(\T0.count[7] ),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1846_ (.RESET_B(net359),
    .D(_0112_),
    .Q(\P0.uptimelat[0] ),
    .CLK(clknet_3_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1847_ (.RESET_B(net359),
    .D(_0113_),
    .Q(\P0.uptimelat[1] ),
    .CLK(clknet_3_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1848_ (.RESET_B(net357),
    .D(_0114_),
    .Q(\P0.uptimelat[2] ),
    .CLK(clknet_3_5__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1849_ (.RESET_B(net356),
    .D(_0009_),
    .Q(\P0.countreg[0] ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1850_ (.RESET_B(net356),
    .D(_0010_),
    .Q(\P0.countreg[1] ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1851_ (.RESET_B(net356),
    .D(_0011_),
    .Q(\P0.countreg[2] ),
    .CLK(clknet_3_2__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1852_ (.RESET_B(net359),
    .D(net49),
    .Q(\P0.uptimereg[0] ),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1853_ (.RESET_B(net359),
    .D(net71),
    .Q(\P0.uptimereg[1] ),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1854_ (.RESET_B(net359),
    .D(net66),
    .Q(\P0.uptimereg[2] ),
    .CLK(clknet_3_6__leaf_clk_regs));
 sg13g2_tiehi _1723__18 (.L_HI(net18));
 sg13g2_tiehi _1722__19 (.L_HI(net19));
 sg13g2_tiehi _1721__20 (.L_HI(net20));
 sg13g2_tiehi _1720__21 (.L_HI(net21));
 sg13g2_tiehi _1719__22 (.L_HI(net22));
 sg13g2_tiehi _1718__23 (.L_HI(net23));
 sg13g2_tiehi _1717__24 (.L_HI(net24));
 sg13g2_tiehi _1716__25 (.L_HI(net25));
 sg13g2_tiehi _1715__26 (.L_HI(net26));
 sg13g2_tiehi _1714__27 (.L_HI(net27));
 sg13g2_tiehi _1713__28 (.L_HI(net28));
 sg13g2_tiehi _1820__29 (.L_HI(net29));
 sg13g2_tiehi _1819__30 (.L_HI(net30));
 sg13g2_tiehi _1818__31 (.L_HI(net31));
 sg13g2_tiehi _1821__32 (.L_HI(net32));
 sg13g2_tiehi tt_um_LnL_SoC_33 (.L_HI(net33));
 sg13g2_tiehi tt_um_LnL_SoC_34 (.L_HI(net34));
 sg13g2_tiehi tt_um_LnL_SoC_35 (.L_HI(net35));
 sg13g2_tiehi tt_um_LnL_SoC_36 (.L_HI(net36));
 sg13g2_tiehi tt_um_LnL_SoC_37 (.L_HI(net37));
 sg13g2_tiehi tt_um_LnL_SoC_38 (.L_HI(net38));
 sg13g2_buf_8 clkbuf_regs_0_clk (.A(clk),
    .X(delaynet_0_clk));
 sg13g2_tielo tt_um_LnL_SoC_14 (.L_LO(net14));
 sg13g2_tielo tt_um_LnL_SoC_15 (.L_LO(net15));
 sg13g2_tielo tt_um_LnL_SoC_16 (.L_LO(net16));
 sg13g2_tiehi _1704__17 (.L_HI(net17));
 sg13g2_buf_1 _1881_ (.A(\P0.clkout ),
    .X(uio_out[2]));
 sg13g2_buf_1 _1882_ (.A(\T0.clkout ),
    .X(uio_out[3]));
 sg13g2_buf_1 _1883_ (.A(\spi0.ssn_out ),
    .X(uio_out[4]));
 sg13g2_buf_1 _1884_ (.A(\spi0.datareg[7] ),
    .X(uio_out[5]));
 sg13g2_buf_1 _1885_ (.A(\spi0.sclk ),
    .X(uio_out[6]));
 sg13g2_buf_1 _1886_ (.A(net279),
    .X(uio_out[7]));
 sg13g2_ebufn_8 _1887_ (.Z(\P0.uptime[0] ),
    .A(net319),
    .TE_B(_0808_));
 sg13g2_ebufn_8 _1888_ (.Z(\P0.uptime[1] ),
    .A(net318),
    .TE_B(_0809_));
 sg13g2_ebufn_8 _1889_ (.Z(\P0.uptime[2] ),
    .A(\cpu0.dr[2] ),
    .TE_B(_0810_));
 sg13g2_ebufn_8 _1890_ (.Z(\cpu0.dataout[3] ),
    .A(\cpu0.dr[3] ),
    .TE_B(_0811_));
 sg13g2_ebufn_8 _1891_ (.Z(\cpu0.dataout[4] ),
    .A(\cpu0.dr[4] ),
    .TE_B(_0812_));
 sg13g2_ebufn_8 _1892_ (.Z(\cpu0.dataout[5] ),
    .A(net317),
    .TE_B(_0813_));
 sg13g2_ebufn_8 _1893_ (.Z(\cpu0.dataout[6] ),
    .A(\cpu0.dr[6] ),
    .TE_B(_0814_));
 sg13g2_ebufn_8 _1894_ (.Z(\cpu0.dataout[7] ),
    .A(net316),
    .TE_B(_0815_));
 sg13g2_ebufn_8 _1895_ (.Z(\P0.uptime[0] ),
    .A(net335),
    .TE_B(_0816_));
 sg13g2_ebufn_8 _1896_ (.Z(\P0.uptime[1] ),
    .A(net333),
    .TE_B(_0817_));
 sg13g2_ebufn_8 _1897_ (.Z(\P0.uptime[2] ),
    .A(net332),
    .TE_B(_0818_));
 sg13g2_ebufn_8 _1898_ (.Z(\cpu0.dataout[3] ),
    .A(net331),
    .TE_B(_0819_));
 sg13g2_ebufn_8 _1899_ (.Z(\cpu0.dataout[4] ),
    .A(net329),
    .TE_B(_0820_));
 sg13g2_ebufn_8 _1900_ (.Z(\cpu0.dataout[5] ),
    .A(net327),
    .TE_B(_0821_));
 sg13g2_ebufn_8 _1901_ (.Z(\cpu0.dataout[6] ),
    .A(net326),
    .TE_B(_0822_));
 sg13g2_ebufn_8 _1902_ (.Z(\cpu0.dataout[7] ),
    .A(net325),
    .TE_B(_0823_));
 sg13g2_ebufn_8 _1903_ (.Z(\P0.uptime[0] ),
    .A(\cpu0.pc[0] ),
    .TE_B(_0824_));
 sg13g2_ebufn_8 _1904_ (.Z(\P0.uptime[1] ),
    .A(\cpu0.pc[1] ),
    .TE_B(_0825_));
 sg13g2_ebufn_8 _1905_ (.Z(\P0.uptime[2] ),
    .A(\cpu0.pc[2] ),
    .TE_B(_0826_));
 sg13g2_ebufn_8 _1906_ (.Z(\cpu0.dataout[3] ),
    .A(\cpu0.pc[3] ),
    .TE_B(_0827_));
 sg13g2_ebufn_8 _1907_ (.Z(\cpu0.dataout[4] ),
    .A(\cpu0.pc[4] ),
    .TE_B(_0828_));
 sg13g2_ebufn_8 _1908_ (.Z(\cpu0.dataout[5] ),
    .A(\cpu0.pc[5] ),
    .TE_B(_0829_));
 sg13g2_ebufn_8 _1909_ (.Z(\cpu0.dataout[6] ),
    .A(\cpu0.pc[6] ),
    .TE_B(_0830_));
 sg13g2_ebufn_8 _1910_ (.Z(\cpu0.dataout[7] ),
    .A(\cpu0.pc[7] ),
    .TE_B(_0831_));
 sg13g2_buf_2 fanout252 (.A(net253),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_0145_),
    .X(net253));
 sg13g2_buf_8 fanout254 (.A(net256),
    .X(net254));
 sg13g2_buf_1 fanout255 (.A(net256),
    .X(net255));
 sg13g2_buf_8 fanout256 (.A(_0145_),
    .X(net256));
 sg13g2_buf_8 fanout257 (.A(net259),
    .X(net257));
 sg13g2_buf_8 fanout258 (.A(net259),
    .X(net258));
 sg13g2_buf_8 fanout259 (.A(_0777_),
    .X(net259));
 sg13g2_buf_8 fanout260 (.A(net262),
    .X(net260));
 sg13g2_buf_1 fanout261 (.A(net262),
    .X(net261));
 sg13g2_buf_1 fanout262 (.A(_0606_),
    .X(net262));
 sg13g2_buf_8 fanout263 (.A(net264),
    .X(net263));
 sg13g2_buf_8 fanout264 (.A(_0429_),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(net266),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_0000_),
    .X(net266));
 sg13g2_buf_8 fanout267 (.A(_0320_),
    .X(net267));
 sg13g2_buf_8 fanout268 (.A(_0184_),
    .X(net268));
 sg13g2_buf_1 fanout269 (.A(_0184_),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(net271),
    .X(net270));
 sg13g2_buf_1 fanout271 (.A(net273),
    .X(net271));
 sg13g2_buf_8 fanout272 (.A(net273),
    .X(net272));
 sg13g2_buf_1 fanout273 (.A(_0725_),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(net275),
    .X(net274));
 sg13g2_buf_1 fanout275 (.A(_0319_),
    .X(net275));
 sg13g2_buf_8 fanout276 (.A(_0318_),
    .X(net276));
 sg13g2_buf_8 fanout277 (.A(_0178_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_0406_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(\cpu0.en_out ),
    .X(net279));
 sg13g2_buf_8 fanout280 (.A(_0779_),
    .X(net280));
 sg13g2_buf_8 fanout281 (.A(net282),
    .X(net281));
 sg13g2_buf_8 fanout282 (.A(_0471_),
    .X(net282));
 sg13g2_buf_8 fanout283 (.A(net284),
    .X(net283));
 sg13g2_buf_8 fanout284 (.A(_0470_),
    .X(net284));
 sg13g2_buf_8 fanout285 (.A(_0297_),
    .X(net285));
 sg13g2_buf_8 fanout286 (.A(net289),
    .X(net286));
 sg13g2_buf_8 fanout287 (.A(net289),
    .X(net287));
 sg13g2_buf_1 fanout288 (.A(net289),
    .X(net288));
 sg13g2_buf_8 fanout289 (.A(_0473_),
    .X(net289));
 sg13g2_buf_8 fanout290 (.A(_0293_),
    .X(net290));
 sg13g2_buf_8 fanout291 (.A(_0288_),
    .X(net291));
 sg13g2_buf_8 fanout292 (.A(_0295_),
    .X(net292));
 sg13g2_buf_8 fanout293 (.A(_0289_),
    .X(net293));
 sg13g2_buf_8 fanout294 (.A(net295),
    .X(net294));
 sg13g2_buf_8 fanout295 (.A(_0247_),
    .X(net295));
 sg13g2_buf_8 fanout296 (.A(_0233_),
    .X(net296));
 sg13g2_buf_8 fanout297 (.A(\cpu0.ir[15] ),
    .X(net297));
 sg13g2_buf_8 fanout298 (.A(net190),
    .X(net298));
 sg13g2_buf_8 fanout299 (.A(net216),
    .X(net299));
 sg13g2_buf_1 fanout300 (.A(net221),
    .X(net300));
 sg13g2_buf_8 fanout301 (.A(net303),
    .X(net301));
 sg13g2_buf_1 fanout302 (.A(net303),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(net304),
    .X(net303));
 sg13g2_buf_8 fanout304 (.A(net220),
    .X(net304));
 sg13g2_buf_8 fanout305 (.A(net306),
    .X(net305));
 sg13g2_buf_8 fanout306 (.A(net310),
    .X(net306));
 sg13g2_buf_8 fanout307 (.A(net308),
    .X(net307));
 sg13g2_buf_8 fanout308 (.A(net309),
    .X(net308));
 sg13g2_buf_8 fanout309 (.A(net310),
    .X(net309));
 sg13g2_buf_8 fanout310 (.A(net195),
    .X(net310));
 sg13g2_buf_8 fanout311 (.A(\cpu0.ir[6] ),
    .X(net311));
 sg13g2_buf_8 fanout312 (.A(net313),
    .X(net312));
 sg13g2_buf_8 fanout313 (.A(net314),
    .X(net313));
 sg13g2_buf_8 fanout314 (.A(net194),
    .X(net314));
 sg13g2_buf_8 fanout315 (.A(net200),
    .X(net315));
 sg13g2_buf_8 fanout316 (.A(net206),
    .X(net316));
 sg13g2_buf_8 fanout317 (.A(net208),
    .X(net317));
 sg13g2_buf_8 fanout318 (.A(net199),
    .X(net318));
 sg13g2_buf_8 fanout319 (.A(net173),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(net321),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(\addr_to_memio[4] ),
    .X(net321));
 sg13g2_buf_8 fanout322 (.A(\addr_to_memio[1] ),
    .X(net322));
 sg13g2_buf_8 fanout323 (.A(net324),
    .X(net323));
 sg13g2_buf_1 fanout324 (.A(\addr_to_memio[0] ),
    .X(net324));
 sg13g2_buf_8 fanout325 (.A(net214),
    .X(net325));
 sg13g2_buf_8 fanout326 (.A(net210),
    .X(net326));
 sg13g2_buf_8 fanout327 (.A(net204),
    .X(net327));
 sg13g2_buf_1 fanout328 (.A(\cpu0.ac[5] ),
    .X(net328));
 sg13g2_buf_8 fanout329 (.A(net191),
    .X(net329));
 sg13g2_buf_1 fanout330 (.A(\cpu0.ac[4] ),
    .X(net330));
 sg13g2_buf_8 fanout331 (.A(net209),
    .X(net331));
 sg13g2_buf_8 fanout332 (.A(net207),
    .X(net332));
 sg13g2_buf_8 fanout333 (.A(net212),
    .X(net333));
 sg13g2_buf_1 fanout334 (.A(net212),
    .X(net334));
 sg13g2_buf_8 fanout335 (.A(net189),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(\cpu0.ac[0] ),
    .X(net336));
 sg13g2_buf_8 fanout337 (.A(\cpu0.t[4] ),
    .X(net337));
 sg13g2_buf_8 fanout338 (.A(net185),
    .X(net338));
 sg13g2_buf_8 fanout339 (.A(net340),
    .X(net339));
 sg13g2_buf_8 fanout340 (.A(net344),
    .X(net340));
 sg13g2_buf_1 fanout341 (.A(net344),
    .X(net341));
 sg13g2_buf_8 fanout342 (.A(net343),
    .X(net342));
 sg13g2_buf_8 fanout343 (.A(net344),
    .X(net343));
 sg13g2_buf_8 fanout344 (.A(\cpu0.t[3] ),
    .X(net344));
 sg13g2_buf_8 fanout345 (.A(net149),
    .X(net345));
 sg13g2_buf_1 fanout346 (.A(net149),
    .X(net346));
 sg13g2_buf_8 fanout347 (.A(net348),
    .X(net347));
 sg13g2_buf_8 fanout348 (.A(net149),
    .X(net348));
 sg13g2_buf_8 fanout349 (.A(net196),
    .X(net349));
 sg13g2_buf_8 fanout350 (.A(net202),
    .X(net350));
 sg13g2_buf_8 fanout351 (.A(net197),
    .X(net351));
 sg13g2_buf_8 fanout352 (.A(net355),
    .X(net352));
 sg13g2_buf_8 fanout353 (.A(net354),
    .X(net353));
 sg13g2_buf_8 fanout354 (.A(net355),
    .X(net354));
 sg13g2_buf_8 fanout355 (.A(net369),
    .X(net355));
 sg13g2_buf_8 fanout356 (.A(net357),
    .X(net356));
 sg13g2_buf_8 fanout357 (.A(net358),
    .X(net357));
 sg13g2_buf_8 fanout358 (.A(net361),
    .X(net358));
 sg13g2_buf_8 fanout359 (.A(net360),
    .X(net359));
 sg13g2_buf_8 fanout360 (.A(net361),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(net369),
    .X(net361));
 sg13g2_buf_8 fanout362 (.A(net364),
    .X(net362));
 sg13g2_buf_8 fanout363 (.A(net364),
    .X(net363));
 sg13g2_buf_8 fanout364 (.A(net369),
    .X(net364));
 sg13g2_buf_8 fanout365 (.A(net368),
    .X(net365));
 sg13g2_buf_8 fanout366 (.A(net368),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(net368),
    .X(net367));
 sg13g2_buf_8 fanout368 (.A(net369),
    .X(net368));
 sg13g2_buf_8 fanout369 (.A(net76),
    .X(net369));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[0]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[1]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[2]),
    .X(net12));
 sg13g2_tielo tt_um_LnL_SoC_13 (.L_LO(net13));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_1_1__leaf_clk));
 sg13g2_buf_8 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_8 clkbuf_3_0__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_0__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_1__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_1__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_2__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_2__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_3__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_3__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_4__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_4__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_5__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_5__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_6__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_6__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_3_7__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_7__leaf_clk_regs));
 sg13g2_inv_1 clkload1 (.A(clknet_3_1__leaf_clk_regs));
 sg13g2_inv_1 clkload2 (.A(clknet_3_2__leaf_clk_regs));
 sg13g2_inv_1 clkload3 (.A(clknet_3_3__leaf_clk_regs));
 sg13g2_inv_1 clkload4 (.A(clknet_3_4__leaf_clk_regs));
 sg13g2_inv_1 clkload5 (.A(clknet_3_5__leaf_clk_regs));
 sg13g2_inv_1 clkload6 (.A(clknet_3_6__leaf_clk_regs));
 sg13g2_inv_1 clkload7 (.A(clknet_3_7__leaf_clk_regs));
 sg13g2_buf_8 \clkbuf_0_cpu0.clk  (.A(\cpu0.clk ),
    .X(\clknet_0_cpu0.clk ));
 sg13g2_buf_8 \clkbuf_4_0_0_cpu0.clk  (.A(\clknet_0_cpu0.clk ),
    .X(\clknet_4_0_0_cpu0.clk ));
 sg13g2_buf_8 \clkbuf_4_1_0_cpu0.clk  (.A(\clknet_0_cpu0.clk ),
    .X(\clknet_4_1_0_cpu0.clk ));
 sg13g2_buf_8 \clkbuf_4_2_0_cpu0.clk  (.A(\clknet_0_cpu0.clk ),
    .X(\clknet_4_2_0_cpu0.clk ));
 sg13g2_buf_8 \clkbuf_4_3_0_cpu0.clk  (.A(\clknet_0_cpu0.clk ),
    .X(\clknet_4_3_0_cpu0.clk ));
 sg13g2_buf_8 \clkbuf_4_4_0_cpu0.clk  (.A(\clknet_0_cpu0.clk ),
    .X(\clknet_4_4_0_cpu0.clk ));
 sg13g2_buf_8 \clkbuf_4_5_0_cpu0.clk  (.A(\clknet_0_cpu0.clk ),
    .X(\clknet_4_5_0_cpu0.clk ));
 sg13g2_buf_8 \clkbuf_4_6_0_cpu0.clk  (.A(\clknet_0_cpu0.clk ),
    .X(\clknet_4_6_0_cpu0.clk ));
 sg13g2_buf_8 \clkbuf_4_7_0_cpu0.clk  (.A(\clknet_0_cpu0.clk ),
    .X(\clknet_4_7_0_cpu0.clk ));
 sg13g2_buf_8 \clkbuf_4_8_0_cpu0.clk  (.A(\clknet_0_cpu0.clk ),
    .X(\clknet_4_8_0_cpu0.clk ));
 sg13g2_buf_8 \clkbuf_4_9_0_cpu0.clk  (.A(\clknet_0_cpu0.clk ),
    .X(\clknet_4_9_0_cpu0.clk ));
 sg13g2_buf_8 \clkbuf_4_10_0_cpu0.clk  (.A(\clknet_0_cpu0.clk ),
    .X(\clknet_4_10_0_cpu0.clk ));
 sg13g2_buf_8 \clkbuf_4_11_0_cpu0.clk  (.A(\clknet_0_cpu0.clk ),
    .X(\clknet_4_11_0_cpu0.clk ));
 sg13g2_buf_8 \clkbuf_4_12_0_cpu0.clk  (.A(\clknet_0_cpu0.clk ),
    .X(\clknet_4_12_0_cpu0.clk ));
 sg13g2_buf_8 \clkbuf_4_13_0_cpu0.clk  (.A(\clknet_0_cpu0.clk ),
    .X(\clknet_4_13_0_cpu0.clk ));
 sg13g2_buf_8 \clkbuf_4_14_0_cpu0.clk  (.A(\clknet_0_cpu0.clk ),
    .X(\clknet_4_14_0_cpu0.clk ));
 sg13g2_buf_8 \clkbuf_4_15_0_cpu0.clk  (.A(\clknet_0_cpu0.clk ),
    .X(\clknet_4_15_0_cpu0.clk ));
 sg13g2_inv_1 clkload8 (.A(\clknet_4_1_0_cpu0.clk ));
 sg13g2_buf_1 clkload9 (.A(\clknet_4_2_0_cpu0.clk ));
 sg13g2_inv_1 clkload10 (.A(\clknet_4_3_0_cpu0.clk ));
 sg13g2_buf_1 clkload11 (.A(\clknet_4_4_0_cpu0.clk ));
 sg13g2_inv_1 clkload12 (.A(\clknet_4_5_0_cpu0.clk ));
 sg13g2_inv_1 clkload13 (.A(\clknet_4_6_0_cpu0.clk ));
 sg13g2_inv_1 clkload14 (.A(\clknet_4_7_0_cpu0.clk ));
 sg13g2_buf_1 clkload15 (.A(\clknet_4_8_0_cpu0.clk ));
 sg13g2_inv_1 clkload16 (.A(\clknet_4_9_0_cpu0.clk ));
 sg13g2_buf_1 clkload17 (.A(\clknet_4_10_0_cpu0.clk ));
 sg13g2_inv_1 clkload18 (.A(\clknet_4_11_0_cpu0.clk ));
 sg13g2_buf_1 clkload19 (.A(\clknet_4_12_0_cpu0.clk ));
 sg13g2_inv_1 clkload20 (.A(\clknet_4_13_0_cpu0.clk ));
 sg13g2_inv_1 clkload21 (.A(\clknet_4_14_0_cpu0.clk ));
 sg13g2_inv_1 clkload22 (.A(\clknet_4_15_0_cpu0.clk ));
 sg13g2_buf_8 delaybuf_0_clk (.A(delaynet_0_clk),
    .X(clk_regs));
 sg13g2_dlygate4sd3_1 hold1 (.A(\P0.countreg[0] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold2 (.A(\cpu0.t[1] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0029_),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold4 (.A(\T0.count[0] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold5 (.A(\P0.countreg[1] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold6 (.A(\T0.count[1] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold7 (.A(\T0.count[7] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0019_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold9 (.A(\P0.uptimelat[0] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0228_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0115_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold12 (.A(\cpu0.t[2] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0030_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold14 (.A(\T0.count[4] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0016_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold16 (.A(\cpu0.t[8] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0036_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold18 (.A(\P0.countreg[2] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold19 (.A(\T0.count[5] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0017_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold21 (.A(\spi0.cntreg[3] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0224_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0111_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold24 (.A(\cpu0.ac15 ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0775_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0060_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold27 (.A(\P0.uptimelat[2] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0117_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold29 (.A(\T0.count[3] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0015_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold31 (.A(\cpu0.ir[4] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold32 (.A(\P0.uptimelat[1] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0116_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold34 (.A(\cpu0.t[7] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0035_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold36 (.A(\cpu0.t[9] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0037_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold38 (.A(rst_n_i),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold39 (.A(\cpu0.ir[11] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold40 (.A(\cpu0.t[5] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold41 (.A(\spi0.datareg[3] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold42 (.A(\spi0.datareg[1] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold43 (.A(\cpu0.pc[9] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0105_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold45 (.A(\spi0.datareg[5] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold46 (.A(\addr_to_memio[10] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0058_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold48 (.A(\cpu0.ir[3] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold49 (.A(\cpu0.ir[1] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold50 (.A(\cpu0.t[6] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0034_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold52 (.A(\addr_to_memio[6] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold53 (.A(\spi0.datareg[6] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold54 (.A(\cpu0.dr[15] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0076_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold56 (.A(\cpu0.ac0 ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0038_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold58 (.A(\spi0.datareg[2] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold59 (.A(\cpu0.ir[8] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold60 (.A(\addr_to_memio[5] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0101_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold62 (.A(\spi0.datareg[4] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold63 (.A(\cpu0.pc[11] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0218_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0107_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold66 (.A(\addr_to_memio[8] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0056_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold68 (.A(\spi0.datareg[0] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold69 (.A(\cpu0.ir[5] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold70 (.A(\addr_to_memio[0] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0048_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold72 (.A(\cpu0.pc[10] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0106_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold74 (.A(\spi0.cntreg[0] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0305_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0109_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold77 (.A(\T0.selreg[2] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold78 (.A(\spi0.cntreg[1] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold79 (.A(\spi0.ssn_out ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold80 (.A(\cpu0.ir[2] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold81 (.A(\addr_to_memio[7] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0055_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold83 (.A(\addr_to_memio[9] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0057_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold85 (.A(\addr_to_memio[11] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0059_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold87 (.A(\spi0.cntreg[2] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold88 (.A(\addr_to_memio[4] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0198_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0100_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold91 (.A(\cpu0.ir[10] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold92 (.A(\cpu0.ir[0] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold93 (.A(\cpu0.pc[6] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0752_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold95 (.A(\cpu0.dr[12] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0073_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold97 (.A(\cpu0.e ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0047_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold99 (.A(\cpu0.decode2.a[1] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold100 (.A(\cpu0.pc[4] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0744_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0052_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold103 (.A(\T0.selreg[1] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold104 (.A(\cpu0.pc[5] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold105 (.A(\cpu0.dr[10] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0127_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0071_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold108 (.A(\cpu0.dr[9] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0123_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0070_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold111 (.A(\cpu0.t[0] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold112 (.A(\cpu0.dr[11] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0072_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold114 (.A(\cpu0.decode2.a[0] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold115 (.A(\cpu0.dr[4] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0065_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold117 (.A(\addr_to_memio[2] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0192_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0098_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold120 (.A(\addr_to_memio[1] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0049_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold122 (.A(\cpu0.ir[15] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold123 (.A(\cpu0.pc[0] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold124 (.A(\cpu0.ac[13] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0025_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold126 (.A(\cpu0.pc[3] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0051_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold128 (.A(\cpu0.ac[9] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0021_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold130 (.A(\cpu0.pc[2] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold131 (.A(\addr_to_memio[3] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0099_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold133 (.A(\cpu0.pc[1] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold134 (.A(\T0.count[2] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold135 (.A(\cpu0.dr[0] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold136 (.A(\cpu0.dr[6] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0804_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold138 (.A(\T0.selreg[0] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold139 (.A(\T0.count[6] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold140 (.A(\cpu0.pc[7] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold141 (.A(\cpu0.dr[13] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold142 (.A(\cpu0.pc[8] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold143 (.A(\cpu0.ac[8] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold144 (.A(\cpu0.ac[14] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0026_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold146 (.A(\cpu0.ac[15] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold147 (.A(\cpu0.t[4] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0032_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold149 (.A(\cpu0.t[10] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold150 (.A(\cpu0.dr[2] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold151 (.A(\cpu0.ac[0] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold152 (.A(\cpu0.decode2.a[2] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold153 (.A(\cpu0.ac[4] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0043_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold155 (.A(\cpu0.dr[14] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold156 (.A(\cpu0.ir[6] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold157 (.A(\cpu0.ir[7] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold158 (.A(\cpu0.ac[12] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold159 (.A(\cpu0.ac[10] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0022_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold161 (.A(\cpu0.dr[1] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold162 (.A(\cpu0.dr[8] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0069_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold164 (.A(\cpu0.ac[11] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0023_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold166 (.A(\cpu0.ac[5] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0044_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold168 (.A(\cpu0.dr[7] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold169 (.A(\cpu0.ac[2] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold170 (.A(\cpu0.dr[5] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold171 (.A(\cpu0.ac[3] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold172 (.A(\cpu0.ac[6] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0045_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold174 (.A(\cpu0.ac[1] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0040_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold176 (.A(\cpu0.ac[7] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0046_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold178 (.A(\cpu0.ir[9] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold179 (.A(\cpu0.dr[3] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold180 (.A(\cpu0.dr[3] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0658_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold182 (.A(\cpu0.ir[9] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold183 (.A(\cpu0.ir[9] ),
    .X(net221));
 sg13g2_antennanp ANTENNA_1 (.A(ui_in[4]));
 sg13g2_antennanp ANTENNA_2 (.A(ui_in[5]));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_fill_2 FILLER_3_140 ();
 sg13g2_decap_4 FILLER_3_154 ();
 sg13g2_fill_2 FILLER_3_158 ();
 sg13g2_decap_8 FILLER_3_169 ();
 sg13g2_decap_8 FILLER_3_176 ();
 sg13g2_decap_8 FILLER_3_183 ();
 sg13g2_decap_8 FILLER_3_190 ();
 sg13g2_decap_8 FILLER_3_197 ();
 sg13g2_decap_8 FILLER_3_204 ();
 sg13g2_decap_8 FILLER_3_211 ();
 sg13g2_decap_8 FILLER_3_218 ();
 sg13g2_decap_8 FILLER_3_225 ();
 sg13g2_decap_8 FILLER_3_232 ();
 sg13g2_decap_8 FILLER_3_239 ();
 sg13g2_decap_8 FILLER_3_246 ();
 sg13g2_decap_8 FILLER_3_253 ();
 sg13g2_decap_8 FILLER_3_260 ();
 sg13g2_decap_8 FILLER_3_267 ();
 sg13g2_decap_8 FILLER_3_274 ();
 sg13g2_decap_8 FILLER_3_281 ();
 sg13g2_decap_8 FILLER_3_288 ();
 sg13g2_decap_8 FILLER_3_295 ();
 sg13g2_decap_8 FILLER_3_302 ();
 sg13g2_decap_8 FILLER_3_309 ();
 sg13g2_decap_8 FILLER_3_316 ();
 sg13g2_decap_8 FILLER_3_323 ();
 sg13g2_decap_8 FILLER_3_330 ();
 sg13g2_decap_8 FILLER_3_337 ();
 sg13g2_decap_8 FILLER_3_344 ();
 sg13g2_decap_8 FILLER_3_351 ();
 sg13g2_decap_8 FILLER_3_358 ();
 sg13g2_decap_8 FILLER_3_365 ();
 sg13g2_decap_8 FILLER_3_372 ();
 sg13g2_decap_8 FILLER_3_379 ();
 sg13g2_decap_8 FILLER_3_386 ();
 sg13g2_decap_8 FILLER_3_393 ();
 sg13g2_decap_8 FILLER_3_400 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_4 FILLER_4_119 ();
 sg13g2_fill_2 FILLER_4_123 ();
 sg13g2_decap_4 FILLER_4_129 ();
 sg13g2_fill_1 FILLER_4_133 ();
 sg13g2_fill_2 FILLER_4_143 ();
 sg13g2_fill_2 FILLER_4_155 ();
 sg13g2_fill_1 FILLER_4_157 ();
 sg13g2_fill_2 FILLER_4_163 ();
 sg13g2_decap_8 FILLER_4_184 ();
 sg13g2_decap_8 FILLER_4_191 ();
 sg13g2_decap_8 FILLER_4_198 ();
 sg13g2_decap_8 FILLER_4_205 ();
 sg13g2_decap_8 FILLER_4_212 ();
 sg13g2_decap_8 FILLER_4_219 ();
 sg13g2_decap_8 FILLER_4_226 ();
 sg13g2_decap_8 FILLER_4_233 ();
 sg13g2_decap_8 FILLER_4_240 ();
 sg13g2_decap_8 FILLER_4_247 ();
 sg13g2_decap_8 FILLER_4_254 ();
 sg13g2_decap_8 FILLER_4_261 ();
 sg13g2_decap_8 FILLER_4_268 ();
 sg13g2_decap_8 FILLER_4_275 ();
 sg13g2_decap_8 FILLER_4_282 ();
 sg13g2_decap_8 FILLER_4_289 ();
 sg13g2_decap_8 FILLER_4_296 ();
 sg13g2_decap_8 FILLER_4_303 ();
 sg13g2_decap_8 FILLER_4_310 ();
 sg13g2_decap_8 FILLER_4_317 ();
 sg13g2_decap_8 FILLER_4_324 ();
 sg13g2_decap_8 FILLER_4_331 ();
 sg13g2_decap_8 FILLER_4_338 ();
 sg13g2_decap_8 FILLER_4_345 ();
 sg13g2_decap_8 FILLER_4_352 ();
 sg13g2_decap_8 FILLER_4_359 ();
 sg13g2_decap_8 FILLER_4_366 ();
 sg13g2_decap_8 FILLER_4_373 ();
 sg13g2_decap_8 FILLER_4_380 ();
 sg13g2_decap_8 FILLER_4_387 ();
 sg13g2_decap_8 FILLER_4_394 ();
 sg13g2_decap_8 FILLER_4_401 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_4 FILLER_5_105 ();
 sg13g2_fill_2 FILLER_5_109 ();
 sg13g2_fill_1 FILLER_5_116 ();
 sg13g2_fill_1 FILLER_5_160 ();
 sg13g2_fill_1 FILLER_5_166 ();
 sg13g2_fill_2 FILLER_5_186 ();
 sg13g2_decap_8 FILLER_5_201 ();
 sg13g2_decap_8 FILLER_5_208 ();
 sg13g2_decap_8 FILLER_5_215 ();
 sg13g2_decap_8 FILLER_5_222 ();
 sg13g2_decap_8 FILLER_5_229 ();
 sg13g2_decap_8 FILLER_5_236 ();
 sg13g2_decap_4 FILLER_5_243 ();
 sg13g2_fill_1 FILLER_5_247 ();
 sg13g2_decap_4 FILLER_5_262 ();
 sg13g2_fill_1 FILLER_5_266 ();
 sg13g2_decap_4 FILLER_5_271 ();
 sg13g2_fill_2 FILLER_5_275 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_4 FILLER_6_28 ();
 sg13g2_fill_1 FILLER_6_32 ();
 sg13g2_decap_8 FILLER_6_44 ();
 sg13g2_decap_8 FILLER_6_51 ();
 sg13g2_decap_8 FILLER_6_58 ();
 sg13g2_decap_8 FILLER_6_65 ();
 sg13g2_decap_8 FILLER_6_72 ();
 sg13g2_decap_4 FILLER_6_79 ();
 sg13g2_fill_1 FILLER_6_83 ();
 sg13g2_fill_2 FILLER_6_99 ();
 sg13g2_decap_8 FILLER_6_209 ();
 sg13g2_decap_4 FILLER_6_216 ();
 sg13g2_fill_1 FILLER_6_220 ();
 sg13g2_fill_1 FILLER_6_239 ();
 sg13g2_fill_1 FILLER_6_272 ();
 sg13g2_decap_8 FILLER_6_299 ();
 sg13g2_decap_8 FILLER_6_306 ();
 sg13g2_decap_8 FILLER_6_313 ();
 sg13g2_decap_8 FILLER_6_320 ();
 sg13g2_decap_8 FILLER_6_327 ();
 sg13g2_decap_8 FILLER_6_334 ();
 sg13g2_decap_8 FILLER_6_341 ();
 sg13g2_decap_8 FILLER_6_348 ();
 sg13g2_decap_8 FILLER_6_355 ();
 sg13g2_decap_8 FILLER_6_362 ();
 sg13g2_decap_8 FILLER_6_369 ();
 sg13g2_decap_8 FILLER_6_376 ();
 sg13g2_decap_8 FILLER_6_383 ();
 sg13g2_decap_8 FILLER_6_390 ();
 sg13g2_decap_8 FILLER_6_397 ();
 sg13g2_decap_4 FILLER_6_404 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_4 FILLER_7_21 ();
 sg13g2_fill_1 FILLER_7_25 ();
 sg13g2_decap_8 FILLER_7_50 ();
 sg13g2_decap_8 FILLER_7_57 ();
 sg13g2_decap_8 FILLER_7_64 ();
 sg13g2_decap_4 FILLER_7_71 ();
 sg13g2_fill_1 FILLER_7_156 ();
 sg13g2_fill_2 FILLER_7_223 ();
 sg13g2_fill_1 FILLER_7_225 ();
 sg13g2_fill_2 FILLER_7_259 ();
 sg13g2_fill_1 FILLER_7_261 ();
 sg13g2_decap_8 FILLER_7_311 ();
 sg13g2_decap_8 FILLER_7_318 ();
 sg13g2_decap_8 FILLER_7_325 ();
 sg13g2_decap_8 FILLER_7_332 ();
 sg13g2_decap_8 FILLER_7_339 ();
 sg13g2_decap_8 FILLER_7_346 ();
 sg13g2_decap_8 FILLER_7_353 ();
 sg13g2_decap_8 FILLER_7_360 ();
 sg13g2_decap_8 FILLER_7_367 ();
 sg13g2_decap_8 FILLER_7_374 ();
 sg13g2_decap_8 FILLER_7_381 ();
 sg13g2_decap_8 FILLER_7_388 ();
 sg13g2_decap_8 FILLER_7_395 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_fill_1 FILLER_8_14 ();
 sg13g2_fill_2 FILLER_8_92 ();
 sg13g2_fill_1 FILLER_8_114 ();
 sg13g2_fill_2 FILLER_8_173 ();
 sg13g2_fill_1 FILLER_8_188 ();
 sg13g2_decap_4 FILLER_8_225 ();
 sg13g2_fill_2 FILLER_8_229 ();
 sg13g2_fill_1 FILLER_8_286 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_fill_2 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_335 ();
 sg13g2_decap_4 FILLER_8_342 ();
 sg13g2_fill_1 FILLER_8_346 ();
 sg13g2_decap_8 FILLER_8_351 ();
 sg13g2_decap_8 FILLER_8_358 ();
 sg13g2_decap_8 FILLER_8_365 ();
 sg13g2_decap_8 FILLER_8_372 ();
 sg13g2_decap_8 FILLER_8_379 ();
 sg13g2_decap_8 FILLER_8_386 ();
 sg13g2_decap_8 FILLER_8_393 ();
 sg13g2_decap_8 FILLER_8_400 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_61 ();
 sg13g2_fill_1 FILLER_9_63 ();
 sg13g2_fill_2 FILLER_9_173 ();
 sg13g2_fill_2 FILLER_9_284 ();
 sg13g2_fill_1 FILLER_9_330 ();
 sg13g2_fill_2 FILLER_9_344 ();
 sg13g2_fill_2 FILLER_9_350 ();
 sg13g2_fill_2 FILLER_9_356 ();
 sg13g2_fill_1 FILLER_9_358 ();
 sg13g2_decap_4 FILLER_9_367 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_fill_1 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_4 FILLER_9_403 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_7 ();
 sg13g2_fill_1 FILLER_10_11 ();
 sg13g2_fill_2 FILLER_10_235 ();
 sg13g2_fill_1 FILLER_10_270 ();
 sg13g2_fill_2 FILLER_10_331 ();
 sg13g2_fill_1 FILLER_10_350 ();
 sg13g2_fill_2 FILLER_10_359 ();
 sg13g2_fill_1 FILLER_10_361 ();
 sg13g2_decap_8 FILLER_10_394 ();
 sg13g2_decap_8 FILLER_10_401 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_fill_1 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_29 ();
 sg13g2_fill_1 FILLER_11_31 ();
 sg13g2_fill_1 FILLER_11_50 ();
 sg13g2_fill_1 FILLER_11_71 ();
 sg13g2_fill_2 FILLER_11_81 ();
 sg13g2_fill_1 FILLER_11_89 ();
 sg13g2_fill_2 FILLER_11_202 ();
 sg13g2_fill_1 FILLER_11_204 ();
 sg13g2_fill_2 FILLER_11_222 ();
 sg13g2_fill_1 FILLER_11_241 ();
 sg13g2_fill_1 FILLER_11_260 ();
 sg13g2_fill_2 FILLER_11_306 ();
 sg13g2_fill_1 FILLER_11_321 ();
 sg13g2_fill_2 FILLER_11_363 ();
 sg13g2_fill_1 FILLER_11_365 ();
 sg13g2_fill_2 FILLER_11_385 ();
 sg13g2_fill_1 FILLER_11_403 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_2 ();
 sg13g2_fill_1 FILLER_12_26 ();
 sg13g2_fill_1 FILLER_12_69 ();
 sg13g2_fill_1 FILLER_12_149 ();
 sg13g2_fill_2 FILLER_12_193 ();
 sg13g2_fill_1 FILLER_12_225 ();
 sg13g2_fill_2 FILLER_12_256 ();
 sg13g2_fill_2 FILLER_12_271 ();
 sg13g2_fill_1 FILLER_12_304 ();
 sg13g2_fill_1 FILLER_12_318 ();
 sg13g2_fill_2 FILLER_12_388 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_fill_2 FILLER_13_27 ();
 sg13g2_fill_1 FILLER_13_87 ();
 sg13g2_fill_1 FILLER_13_224 ();
 sg13g2_fill_2 FILLER_13_313 ();
 sg13g2_fill_1 FILLER_13_320 ();
 sg13g2_fill_1 FILLER_13_326 ();
 sg13g2_fill_1 FILLER_13_390 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_fill_1 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_112 ();
 sg13g2_fill_1 FILLER_14_127 ();
 sg13g2_fill_1 FILLER_14_134 ();
 sg13g2_fill_2 FILLER_14_186 ();
 sg13g2_fill_1 FILLER_14_188 ();
 sg13g2_fill_2 FILLER_14_216 ();
 sg13g2_fill_2 FILLER_14_230 ();
 sg13g2_fill_1 FILLER_14_258 ();
 sg13g2_fill_1 FILLER_14_271 ();
 sg13g2_fill_2 FILLER_14_296 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_25 ();
 sg13g2_fill_1 FILLER_15_221 ();
 sg13g2_fill_1 FILLER_15_235 ();
 sg13g2_fill_2 FILLER_15_297 ();
 sg13g2_fill_1 FILLER_15_315 ();
 sg13g2_fill_2 FILLER_15_379 ();
 sg13g2_fill_1 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_29 ();
 sg13g2_fill_1 FILLER_16_31 ();
 sg13g2_fill_1 FILLER_16_65 ();
 sg13g2_fill_2 FILLER_16_124 ();
 sg13g2_fill_2 FILLER_16_194 ();
 sg13g2_fill_1 FILLER_16_196 ();
 sg13g2_fill_1 FILLER_16_207 ();
 sg13g2_fill_2 FILLER_16_240 ();
 sg13g2_fill_1 FILLER_16_262 ();
 sg13g2_fill_2 FILLER_16_289 ();
 sg13g2_fill_1 FILLER_16_306 ();
 sg13g2_fill_1 FILLER_16_312 ();
 sg13g2_fill_2 FILLER_16_335 ();
 sg13g2_fill_1 FILLER_16_362 ();
 sg13g2_fill_1 FILLER_16_382 ();
 sg13g2_fill_1 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_36 ();
 sg13g2_fill_1 FILLER_17_38 ();
 sg13g2_fill_1 FILLER_17_78 ();
 sg13g2_fill_2 FILLER_17_111 ();
 sg13g2_fill_2 FILLER_17_229 ();
 sg13g2_fill_1 FILLER_17_268 ();
 sg13g2_fill_1 FILLER_17_303 ();
 sg13g2_fill_2 FILLER_17_345 ();
 sg13g2_fill_1 FILLER_17_347 ();
 sg13g2_fill_2 FILLER_17_364 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_fill_1 FILLER_18_30 ();
 sg13g2_fill_2 FILLER_18_58 ();
 sg13g2_fill_2 FILLER_18_96 ();
 sg13g2_fill_2 FILLER_18_136 ();
 sg13g2_fill_2 FILLER_18_226 ();
 sg13g2_fill_1 FILLER_18_228 ();
 sg13g2_fill_2 FILLER_18_242 ();
 sg13g2_fill_2 FILLER_18_281 ();
 sg13g2_fill_2 FILLER_18_291 ();
 sg13g2_fill_1 FILLER_18_302 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_26 ();
 sg13g2_fill_2 FILLER_19_39 ();
 sg13g2_fill_2 FILLER_19_60 ();
 sg13g2_fill_1 FILLER_19_62 ();
 sg13g2_fill_1 FILLER_19_98 ();
 sg13g2_fill_1 FILLER_19_124 ();
 sg13g2_fill_2 FILLER_19_139 ();
 sg13g2_fill_1 FILLER_19_255 ();
 sg13g2_fill_1 FILLER_19_313 ();
 sg13g2_fill_1 FILLER_19_318 ();
 sg13g2_fill_1 FILLER_19_336 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_7 ();
 sg13g2_fill_2 FILLER_20_15 ();
 sg13g2_fill_1 FILLER_20_17 ();
 sg13g2_fill_2 FILLER_20_28 ();
 sg13g2_fill_1 FILLER_20_30 ();
 sg13g2_fill_2 FILLER_20_39 ();
 sg13g2_fill_2 FILLER_20_61 ();
 sg13g2_decap_8 FILLER_20_78 ();
 sg13g2_fill_1 FILLER_20_85 ();
 sg13g2_decap_8 FILLER_20_128 ();
 sg13g2_fill_1 FILLER_20_135 ();
 sg13g2_fill_1 FILLER_20_176 ();
 sg13g2_fill_2 FILLER_20_218 ();
 sg13g2_fill_1 FILLER_20_234 ();
 sg13g2_fill_2 FILLER_20_240 ();
 sg13g2_fill_1 FILLER_20_242 ();
 sg13g2_fill_2 FILLER_20_271 ();
 sg13g2_fill_1 FILLER_20_311 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_2 ();
 sg13g2_fill_2 FILLER_21_30 ();
 sg13g2_fill_2 FILLER_21_51 ();
 sg13g2_decap_4 FILLER_21_69 ();
 sg13g2_fill_2 FILLER_21_83 ();
 sg13g2_fill_1 FILLER_21_85 ();
 sg13g2_decap_4 FILLER_21_107 ();
 sg13g2_fill_2 FILLER_21_111 ();
 sg13g2_decap_8 FILLER_21_117 ();
 sg13g2_fill_1 FILLER_21_150 ();
 sg13g2_fill_1 FILLER_21_176 ();
 sg13g2_fill_1 FILLER_21_221 ();
 sg13g2_fill_1 FILLER_21_274 ();
 sg13g2_fill_1 FILLER_21_292 ();
 sg13g2_fill_1 FILLER_21_357 ();
 sg13g2_fill_2 FILLER_21_369 ();
 sg13g2_fill_2 FILLER_21_393 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_7 ();
 sg13g2_fill_2 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_78 ();
 sg13g2_decap_4 FILLER_22_85 ();
 sg13g2_fill_2 FILLER_22_89 ();
 sg13g2_fill_2 FILLER_22_101 ();
 sg13g2_fill_1 FILLER_22_158 ();
 sg13g2_fill_2 FILLER_22_194 ();
 sg13g2_fill_2 FILLER_22_314 ();
 sg13g2_fill_1 FILLER_22_316 ();
 sg13g2_fill_1 FILLER_22_322 ();
 sg13g2_fill_2 FILLER_22_364 ();
 sg13g2_fill_2 FILLER_22_379 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_24 ();
 sg13g2_fill_1 FILLER_23_41 ();
 sg13g2_fill_2 FILLER_23_47 ();
 sg13g2_fill_2 FILLER_23_70 ();
 sg13g2_fill_2 FILLER_23_106 ();
 sg13g2_fill_1 FILLER_23_108 ();
 sg13g2_fill_2 FILLER_23_119 ();
 sg13g2_fill_1 FILLER_23_131 ();
 sg13g2_fill_1 FILLER_23_137 ();
 sg13g2_fill_2 FILLER_23_142 ();
 sg13g2_fill_2 FILLER_23_239 ();
 sg13g2_fill_2 FILLER_23_274 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_4 ();
 sg13g2_decap_8 FILLER_24_64 ();
 sg13g2_decap_8 FILLER_24_71 ();
 sg13g2_fill_1 FILLER_24_98 ();
 sg13g2_fill_2 FILLER_24_256 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_fill_2 FILLER_25_21 ();
 sg13g2_fill_2 FILLER_25_95 ();
 sg13g2_fill_1 FILLER_25_136 ();
 sg13g2_fill_2 FILLER_25_145 ();
 sg13g2_fill_2 FILLER_25_184 ();
 sg13g2_fill_1 FILLER_25_232 ();
 sg13g2_fill_2 FILLER_25_244 ();
 sg13g2_fill_2 FILLER_25_292 ();
 sg13g2_fill_1 FILLER_25_294 ();
 sg13g2_fill_2 FILLER_25_326 ();
 sg13g2_fill_2 FILLER_25_356 ();
 sg13g2_fill_2 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_4 FILLER_26_14 ();
 sg13g2_fill_1 FILLER_26_18 ();
 sg13g2_fill_2 FILLER_26_64 ();
 sg13g2_decap_4 FILLER_26_74 ();
 sg13g2_fill_2 FILLER_26_113 ();
 sg13g2_fill_1 FILLER_26_195 ();
 sg13g2_fill_2 FILLER_26_214 ();
 sg13g2_fill_1 FILLER_26_329 ();
 sg13g2_fill_2 FILLER_26_351 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_12 ();
 sg13g2_fill_1 FILLER_27_14 ();
 sg13g2_fill_1 FILLER_27_91 ();
 sg13g2_fill_2 FILLER_27_131 ();
 sg13g2_fill_1 FILLER_27_236 ();
 sg13g2_fill_1 FILLER_27_283 ();
 sg13g2_fill_2 FILLER_27_297 ();
 sg13g2_fill_2 FILLER_27_354 ();
 sg13g2_fill_2 FILLER_28_72 ();
 sg13g2_fill_2 FILLER_28_206 ();
 sg13g2_fill_2 FILLER_28_294 ();
 sg13g2_fill_1 FILLER_28_296 ();
 sg13g2_fill_1 FILLER_28_369 ();
 sg13g2_fill_2 FILLER_28_398 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_86 ();
 sg13g2_fill_1 FILLER_29_189 ();
 sg13g2_fill_1 FILLER_29_200 ();
 sg13g2_fill_1 FILLER_29_223 ();
 sg13g2_fill_1 FILLER_29_251 ();
 sg13g2_fill_2 FILLER_29_295 ();
 sg13g2_fill_1 FILLER_29_297 ();
 sg13g2_fill_2 FILLER_29_305 ();
 sg13g2_fill_1 FILLER_29_332 ();
 sg13g2_fill_2 FILLER_29_395 ();
 sg13g2_fill_1 FILLER_29_397 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_112 ();
 sg13g2_fill_2 FILLER_30_203 ();
 sg13g2_fill_1 FILLER_30_205 ();
 sg13g2_fill_1 FILLER_30_245 ();
 sg13g2_fill_1 FILLER_30_256 ();
 sg13g2_fill_1 FILLER_30_331 ();
 sg13g2_fill_1 FILLER_30_383 ();
 sg13g2_fill_1 FILLER_31_133 ();
 sg13g2_fill_1 FILLER_31_167 ();
 sg13g2_fill_2 FILLER_31_200 ();
 sg13g2_fill_1 FILLER_31_202 ();
 sg13g2_fill_2 FILLER_31_225 ();
 sg13g2_fill_2 FILLER_31_296 ();
 sg13g2_fill_2 FILLER_31_309 ();
 sg13g2_fill_2 FILLER_31_324 ();
 sg13g2_fill_1 FILLER_31_344 ();
 sg13g2_fill_2 FILLER_31_351 ();
 sg13g2_fill_1 FILLER_31_353 ();
 sg13g2_fill_1 FILLER_31_359 ();
 sg13g2_fill_2 FILLER_31_375 ();
 sg13g2_fill_1 FILLER_32_53 ();
 sg13g2_fill_2 FILLER_32_190 ();
 sg13g2_fill_1 FILLER_32_250 ();
 sg13g2_fill_2 FILLER_32_264 ();
 sg13g2_fill_1 FILLER_32_266 ();
 sg13g2_fill_1 FILLER_32_312 ();
 sg13g2_fill_2 FILLER_32_358 ();
 sg13g2_fill_1 FILLER_32_360 ();
 sg13g2_fill_1 FILLER_32_380 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_96 ();
 sg13g2_fill_1 FILLER_33_165 ();
 sg13g2_fill_2 FILLER_33_318 ();
 sg13g2_fill_1 FILLER_33_350 ();
 sg13g2_fill_2 FILLER_33_378 ();
 sg13g2_fill_1 FILLER_33_386 ();
 sg13g2_fill_1 FILLER_34_125 ();
 sg13g2_fill_2 FILLER_34_172 ();
 sg13g2_fill_1 FILLER_34_220 ();
 sg13g2_fill_2 FILLER_34_286 ();
 sg13g2_fill_1 FILLER_34_325 ();
 sg13g2_fill_2 FILLER_34_345 ();
 sg13g2_fill_1 FILLER_35_53 ();
 sg13g2_fill_1 FILLER_35_64 ();
 sg13g2_fill_1 FILLER_35_131 ();
 sg13g2_fill_1 FILLER_35_234 ();
 sg13g2_fill_2 FILLER_35_331 ();
 sg13g2_fill_2 FILLER_35_398 ();
 sg13g2_fill_1 FILLER_36_54 ();
 sg13g2_fill_1 FILLER_36_90 ();
 sg13g2_fill_1 FILLER_36_119 ();
 sg13g2_fill_1 FILLER_36_161 ();
 sg13g2_fill_1 FILLER_36_182 ();
 sg13g2_fill_2 FILLER_36_231 ();
 sg13g2_fill_1 FILLER_36_233 ();
 sg13g2_fill_1 FILLER_36_314 ();
 sg13g2_fill_2 FILLER_36_346 ();
 sg13g2_fill_1 FILLER_36_362 ();
 sg13g2_fill_2 FILLER_37_131 ();
 sg13g2_fill_1 FILLER_37_138 ();
 sg13g2_fill_1 FILLER_37_332 ();
 sg13g2_fill_1 FILLER_37_385 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_fill_2 FILLER_38_176 ();
 sg13g2_fill_1 FILLER_38_192 ();
 sg13g2_fill_1 FILLER_38_271 ();
 sg13g2_fill_1 FILLER_38_312 ();
 sg13g2_fill_1 FILLER_38_369 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net13;
 assign uio_oe[1] = net14;
 assign uio_oe[2] = net33;
 assign uio_oe[3] = net34;
 assign uio_oe[4] = net35;
 assign uio_oe[5] = net36;
 assign uio_oe[6] = net37;
 assign uio_oe[7] = net38;
 assign uio_out[0] = net15;
 assign uio_out[1] = net16;
endmodule
