module tt_um_coastalwhite_canright_sbox (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire clknet_0_clk;
 wire \data_i[0] ;
 wire \data_i[1] ;
 wire \data_i[2] ;
 wire \data_i[3] ;
 wire \data_i[4] ;
 wire \data_i[5] ;
 wire \data_i[6] ;
 wire \data_i[7] ;
 wire \key[0] ;
 wire \key[1] ;
 wire \key[2] ;
 wire \key[3] ;
 wire \key[4] ;
 wire \key[5] ;
 wire \key[6] ;
 wire \key[7] ;
 wire \mask_i[0] ;
 wire \mask_i[1] ;
 wire \mask_i[2] ;
 wire \mask_i[3] ;
 wire \mask_i[4] ;
 wire \mask_i[5] ;
 wire \mask_i[6] ;
 wire \mask_i[7] ;
 wire \prd_i[0] ;
 wire \prd_i[10] ;
 wire \prd_i[11] ;
 wire \prd_i[12] ;
 wire \prd_i[13] ;
 wire \prd_i[14] ;
 wire \prd_i[15] ;
 wire \prd_i[16] ;
 wire \prd_i[17] ;
 wire \prd_i[1] ;
 wire \prd_i[2] ;
 wire \prd_i[3] ;
 wire \prd_i[4] ;
 wire \prd_i[5] ;
 wire \prd_i[6] ;
 wire \prd_i[7] ;
 wire \prd_i[8] ;
 wire \prd_i[9] ;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;

 sg13g2_inv_1 _0949_ (.Y(_0057_),
    .A(net113));
 sg13g2_inv_2 _0950_ (.Y(_0058_),
    .A(net8));
 sg13g2_inv_2 _0951_ (.Y(_0059_),
    .A(net7));
 sg13g2_inv_2 _0952_ (.Y(_0060_),
    .A(net6));
 sg13g2_inv_4 _0953_ (.A(net5),
    .Y(_0061_));
 sg13g2_inv_4 _0954_ (.A(net4),
    .Y(_0062_));
 sg13g2_inv_2 _0955_ (.Y(_0063_),
    .A(net3));
 sg13g2_inv_4 _0956_ (.A(net2),
    .Y(_0064_));
 sg13g2_inv_4 _0957_ (.A(net1),
    .Y(_0065_));
 sg13g2_inv_4 _0958_ (.A(net97),
    .Y(_0066_));
 sg13g2_inv_2 _0959_ (.Y(_0067_),
    .A(net93));
 sg13g2_nand2b_2 _0960_ (.Y(_0068_),
    .B(net9),
    .A_N(net10));
 sg13g2_nor3_2 _0961_ (.A(net11),
    .B(net12),
    .C(_0068_),
    .Y(_0069_));
 sg13g2_o21ai_1 _0962_ (.B1(net95),
    .Y(_0070_),
    .A1(net145),
    .A2(net82));
 sg13g2_a21oi_1 _0963_ (.A1(_0065_),
    .A2(net82),
    .Y(_0000_),
    .B1(_0070_));
 sg13g2_o21ai_1 _0964_ (.B1(net95),
    .Y(_0071_),
    .A1(net160),
    .A2(net82));
 sg13g2_a21oi_1 _0965_ (.A1(_0064_),
    .A2(net82),
    .Y(_0001_),
    .B1(_0071_));
 sg13g2_o21ai_1 _0966_ (.B1(net95),
    .Y(_0072_),
    .A1(net163),
    .A2(net82));
 sg13g2_a21oi_1 _0967_ (.A1(_0063_),
    .A2(net82),
    .Y(_0002_),
    .B1(_0072_));
 sg13g2_o21ai_1 _0968_ (.B1(net96),
    .Y(_0073_),
    .A1(net146),
    .A2(net83));
 sg13g2_a21oi_1 _0969_ (.A1(_0062_),
    .A2(net83),
    .Y(_0003_),
    .B1(_0073_));
 sg13g2_o21ai_1 _0970_ (.B1(net95),
    .Y(_0074_),
    .A1(net144),
    .A2(_0069_));
 sg13g2_a21oi_1 _0971_ (.A1(_0061_),
    .A2(net83),
    .Y(_0004_),
    .B1(_0074_));
 sg13g2_o21ai_1 _0972_ (.B1(net95),
    .Y(_0075_),
    .A1(net141),
    .A2(net82));
 sg13g2_a21oi_1 _0973_ (.A1(_0060_),
    .A2(net82),
    .Y(_0005_),
    .B1(_0075_));
 sg13g2_o21ai_1 _0974_ (.B1(net96),
    .Y(_0076_),
    .A1(net158),
    .A2(net83));
 sg13g2_a21oi_1 _0975_ (.A1(_0059_),
    .A2(net83),
    .Y(_0006_),
    .B1(_0076_));
 sg13g2_o21ai_1 _0976_ (.B1(net97),
    .Y(_0077_),
    .A1(net154),
    .A2(net83));
 sg13g2_a21oi_1 _0977_ (.A1(_0058_),
    .A2(net83),
    .Y(_0007_),
    .B1(_0077_));
 sg13g2_nand2b_2 _0978_ (.Y(_0078_),
    .B(net10),
    .A_N(net9));
 sg13g2_nor3_2 _0979_ (.A(net11),
    .B(net12),
    .C(_0078_),
    .Y(_0079_));
 sg13g2_o21ai_1 _0980_ (.B1(net95),
    .Y(_0080_),
    .A1(net147),
    .A2(net80));
 sg13g2_a21oi_1 _0981_ (.A1(_0065_),
    .A2(net80),
    .Y(_0008_),
    .B1(_0080_));
 sg13g2_o21ai_1 _0982_ (.B1(net95),
    .Y(_0081_),
    .A1(net161),
    .A2(net80));
 sg13g2_a21oi_1 _0983_ (.A1(_0064_),
    .A2(net80),
    .Y(_0009_),
    .B1(_0081_));
 sg13g2_o21ai_1 _0984_ (.B1(net95),
    .Y(_0082_),
    .A1(net162),
    .A2(net80));
 sg13g2_a21oi_1 _0985_ (.A1(_0063_),
    .A2(net80),
    .Y(_0010_),
    .B1(_0082_));
 sg13g2_o21ai_1 _0986_ (.B1(net96),
    .Y(_0083_),
    .A1(net143),
    .A2(net81));
 sg13g2_a21oi_1 _0987_ (.A1(_0062_),
    .A2(net81),
    .Y(_0011_),
    .B1(_0083_));
 sg13g2_o21ai_1 _0988_ (.B1(net96),
    .Y(_0084_),
    .A1(net156),
    .A2(_0079_));
 sg13g2_a21oi_1 _0989_ (.A1(_0061_),
    .A2(net81),
    .Y(_0012_),
    .B1(_0084_));
 sg13g2_o21ai_1 _0990_ (.B1(net96),
    .Y(_0085_),
    .A1(net150),
    .A2(net80));
 sg13g2_a21oi_1 _0991_ (.A1(_0060_),
    .A2(net80),
    .Y(_0013_),
    .B1(_0085_));
 sg13g2_o21ai_1 _0992_ (.B1(net97),
    .Y(_0086_),
    .A1(net153),
    .A2(net81));
 sg13g2_a21oi_1 _0993_ (.A1(_0059_),
    .A2(net81),
    .Y(_0014_),
    .B1(_0086_));
 sg13g2_o21ai_1 _0994_ (.B1(net97),
    .Y(_0087_),
    .A1(net155),
    .A2(net81));
 sg13g2_a21oi_1 _0995_ (.A1(_0058_),
    .A2(net81),
    .Y(_0015_),
    .B1(_0087_));
 sg13g2_nand2b_2 _0996_ (.Y(_0088_),
    .B(net12),
    .A_N(net11));
 sg13g2_a21oi_1 _0997_ (.A1(net10),
    .A2(net9),
    .Y(_0089_),
    .B1(net84));
 sg13g2_a21o_2 _0998_ (.A2(net9),
    .A1(net10),
    .B1(net84),
    .X(_0090_));
 sg13g2_nor2_2 _0999_ (.A(net10),
    .B(net9),
    .Y(_0091_));
 sg13g2_nor2_2 _1000_ (.A(net79),
    .B(_0091_),
    .Y(_0092_));
 sg13g2_nand2b_2 _1001_ (.Y(_0093_),
    .B(_0089_),
    .A_N(_0091_));
 sg13g2_xor2_1 _1002_ (.B(\data_i[6] ),
    .A(\key[6] ),
    .X(_0094_));
 sg13g2_xnor2_1 _1003_ (.Y(_0095_),
    .A(\key[5] ),
    .B(\data_i[5] ));
 sg13g2_xnor2_1 _1004_ (.Y(_0096_),
    .A(_0094_),
    .B(_0095_));
 sg13g2_nand2_2 _1005_ (.Y(_0097_),
    .A(net85),
    .B(_0096_));
 sg13g2_xor2_1 _1006_ (.B(\data_i[7] ),
    .A(\key[7] ),
    .X(_0098_));
 sg13g2_nand2_2 _1007_ (.Y(_0099_),
    .A(net85),
    .B(_0098_));
 sg13g2_xor2_1 _1008_ (.B(_0099_),
    .A(_0097_),
    .X(_0100_));
 sg13g2_xnor2_1 _1009_ (.Y(_0101_),
    .A(\key[4] ),
    .B(\data_i[4] ));
 sg13g2_xnor2_1 _1010_ (.Y(_0102_),
    .A(_0096_),
    .B(_0101_));
 sg13g2_nand2_2 _1011_ (.Y(_0103_),
    .A(net85),
    .B(_0102_));
 sg13g2_xor2_1 _1012_ (.B(_0103_),
    .A(_0100_),
    .X(_0104_));
 sg13g2_xor2_1 _1013_ (.B(\data_i[2] ),
    .A(\key[2] ),
    .X(_0105_));
 sg13g2_xnor2_1 _1014_ (.Y(_0106_),
    .A(\key[2] ),
    .B(\data_i[2] ));
 sg13g2_xnor2_1 _1015_ (.Y(_0107_),
    .A(_0094_),
    .B(_0106_));
 sg13g2_nand2_1 _1016_ (.Y(_0108_),
    .A(net85),
    .B(_0107_));
 sg13g2_xor2_1 _1017_ (.B(\data_i[0] ),
    .A(\key[0] ),
    .X(_0109_));
 sg13g2_nand2_2 _1018_ (.Y(_0110_),
    .A(net85),
    .B(_0109_));
 sg13g2_xor2_1 _1019_ (.B(\data_i[1] ),
    .A(\key[1] ),
    .X(_0111_));
 sg13g2_xnor2_1 _1020_ (.Y(_0112_),
    .A(\key[1] ),
    .B(\data_i[1] ));
 sg13g2_nand2_2 _1021_ (.Y(_0113_),
    .A(net85),
    .B(_0111_));
 sg13g2_mux2_1 _1022_ (.A0(_0111_),
    .A1(_0113_),
    .S(_0110_),
    .X(_0114_));
 sg13g2_xor2_1 _1023_ (.B(\data_i[3] ),
    .A(\key[3] ),
    .X(_0115_));
 sg13g2_nand2_1 _1024_ (.Y(_0116_),
    .A(net85),
    .B(_0115_));
 sg13g2_xor2_1 _1025_ (.B(_0116_),
    .A(_0114_),
    .X(_0117_));
 sg13g2_xnor2_1 _1026_ (.Y(_0118_),
    .A(_0108_),
    .B(_0117_));
 sg13g2_xor2_1 _1027_ (.B(_0110_),
    .A(_0097_),
    .X(_0119_));
 sg13g2_xor2_1 _1028_ (.B(_0119_),
    .A(_0099_),
    .X(_0120_));
 sg13g2_nor2b_2 _1029_ (.A(_0118_),
    .B_N(_0120_),
    .Y(_0121_));
 sg13g2_xnor2_1 _1030_ (.Y(_0122_),
    .A(_0118_),
    .B(_0120_));
 sg13g2_xnor2_1 _1031_ (.Y(_0123_),
    .A(_0097_),
    .B(_0114_));
 sg13g2_xnor2_1 _1032_ (.Y(_0124_),
    .A(_0120_),
    .B(_0123_));
 sg13g2_xnor2_1 _1033_ (.Y(_0125_),
    .A(_0118_),
    .B(_0119_));
 sg13g2_nor2_1 _1034_ (.A(_0124_),
    .B(_0125_),
    .Y(_0126_));
 sg13g2_nor3_1 _1035_ (.A(_0121_),
    .B(_0124_),
    .C(_0125_),
    .Y(_0127_));
 sg13g2_a21oi_1 _1036_ (.A1(net85),
    .A2(_0111_),
    .Y(_0128_),
    .B1(_0121_));
 sg13g2_o21ai_1 _1037_ (.B1(_0128_),
    .Y(_0129_),
    .A1(_0119_),
    .A2(_0126_));
 sg13g2_o21ai_1 _1038_ (.B1(_0129_),
    .Y(_0130_),
    .A1(_0113_),
    .A2(_0127_));
 sg13g2_xor2_1 _1039_ (.B(_0130_),
    .A(_0122_),
    .X(_0131_));
 sg13g2_xor2_1 _1040_ (.B(_0118_),
    .A(_0110_),
    .X(_0132_));
 sg13g2_nor2_1 _1041_ (.A(_0104_),
    .B(_0132_),
    .Y(_0133_));
 sg13g2_xnor2_1 _1042_ (.Y(_0134_),
    .A(_0104_),
    .B(_0117_));
 sg13g2_xnor2_1 _1043_ (.Y(_0135_),
    .A(_0119_),
    .B(_0134_));
 sg13g2_xnor2_1 _1044_ (.Y(_0136_),
    .A(_0132_),
    .B(_0135_));
 sg13g2_nand2_1 _1045_ (.Y(_0137_),
    .A(net13),
    .B(_0105_));
 sg13g2_xor2_1 _1046_ (.B(_0137_),
    .A(_0114_),
    .X(_0138_));
 sg13g2_xnor2_1 _1047_ (.Y(_0139_),
    .A(_0100_),
    .B(_0138_));
 sg13g2_inv_2 _1048_ (.Y(_0140_),
    .A(_0139_));
 sg13g2_xor2_1 _1049_ (.B(_0137_),
    .A(_0099_),
    .X(_0141_));
 sg13g2_xor2_1 _1050_ (.B(_0141_),
    .A(_0104_),
    .X(_0142_));
 sg13g2_nor2_1 _1051_ (.A(_0136_),
    .B(_0142_),
    .Y(_0143_));
 sg13g2_xnor2_1 _1052_ (.Y(_0144_),
    .A(_0133_),
    .B(_0143_));
 sg13g2_xnor2_1 _1053_ (.Y(_0145_),
    .A(_0131_),
    .B(_0144_));
 sg13g2_nor2b_1 _1054_ (.A(_0135_),
    .B_N(_0141_),
    .Y(_0146_));
 sg13g2_xnor2_1 _1055_ (.Y(_0147_),
    .A(_0133_),
    .B(_0146_));
 sg13g2_nor2_1 _1056_ (.A(_0134_),
    .B(_0140_),
    .Y(_0148_));
 sg13g2_xnor2_1 _1057_ (.Y(_0149_),
    .A(_0134_),
    .B(_0140_));
 sg13g2_xnor2_1 _1058_ (.Y(_0150_),
    .A(_0113_),
    .B(_0149_));
 sg13g2_nor2_1 _1059_ (.A(_0102_),
    .B(_0110_),
    .Y(_0151_));
 sg13g2_xor2_1 _1060_ (.B(_0110_),
    .A(_0103_),
    .X(_0152_));
 sg13g2_xnor2_1 _1061_ (.Y(_0153_),
    .A(_0139_),
    .B(_0152_));
 sg13g2_xnor2_1 _1062_ (.Y(_0154_),
    .A(_0110_),
    .B(_0134_));
 sg13g2_a21oi_1 _1063_ (.A1(_0153_),
    .A2(_0154_),
    .Y(_0155_),
    .B1(_0151_));
 sg13g2_a21oi_1 _1064_ (.A1(_0148_),
    .A2(_0151_),
    .Y(_0156_),
    .B1(_0155_));
 sg13g2_xnor2_1 _1065_ (.Y(_0157_),
    .A(_0147_),
    .B(_0156_));
 sg13g2_xnor2_1 _1066_ (.Y(_0158_),
    .A(_0150_),
    .B(_0157_));
 sg13g2_nand2b_1 _1067_ (.Y(_0159_),
    .B(_0158_),
    .A_N(_0145_));
 sg13g2_xnor2_1 _1068_ (.Y(_0160_),
    .A(_0121_),
    .B(_0126_));
 sg13g2_xnor2_1 _1069_ (.Y(_0161_),
    .A(_0147_),
    .B(_0160_));
 sg13g2_and3_1 _1070_ (.X(_0162_),
    .A(_0103_),
    .B(_0110_),
    .C(_0140_));
 sg13g2_a22oi_1 _1071_ (.Y(_0163_),
    .B1(_0153_),
    .B2(_0154_),
    .A2(_0140_),
    .A1(_0134_));
 sg13g2_a21oi_1 _1072_ (.A1(_0134_),
    .A2(_0162_),
    .Y(_0164_),
    .B1(_0163_));
 sg13g2_xor2_1 _1073_ (.B(_0122_),
    .A(_0103_),
    .X(_0165_));
 sg13g2_xnor2_1 _1074_ (.Y(_0166_),
    .A(_0164_),
    .B(_0165_));
 sg13g2_xnor2_1 _1075_ (.Y(_0167_),
    .A(_0144_),
    .B(_0166_));
 sg13g2_inv_1 _1076_ (.Y(_0168_),
    .A(_0167_));
 sg13g2_nand2_1 _1077_ (.Y(_0169_),
    .A(_0145_),
    .B(_0167_));
 sg13g2_nor2_1 _1078_ (.A(_0158_),
    .B(_0161_),
    .Y(_0170_));
 sg13g2_xor2_1 _1079_ (.B(_0170_),
    .A(_0169_),
    .X(_0171_));
 sg13g2_and2_1 _1080_ (.A(_0145_),
    .B(_0171_),
    .X(_0172_));
 sg13g2_inv_1 _1081_ (.Y(_0173_),
    .A(_0172_));
 sg13g2_a21o_2 _1082_ (.A2(_0161_),
    .A1(_0159_),
    .B1(_0172_),
    .X(_0174_));
 sg13g2_and2_1 _1083_ (.A(_0158_),
    .B(_0167_),
    .X(_0175_));
 sg13g2_nor2_1 _1084_ (.A(_0158_),
    .B(_0167_),
    .Y(_0176_));
 sg13g2_nor2_1 _1085_ (.A(_0175_),
    .B(_0176_),
    .Y(_0177_));
 sg13g2_nand2_1 _1086_ (.Y(_0178_),
    .A(_0171_),
    .B(_0177_));
 sg13g2_a21oi_1 _1087_ (.A1(_0158_),
    .A2(_0161_),
    .Y(_0179_),
    .B1(_0178_));
 sg13g2_nor2_1 _1088_ (.A(_0175_),
    .B(_0179_),
    .Y(_0180_));
 sg13g2_xnor2_1 _1089_ (.Y(_0181_),
    .A(_0174_),
    .B(_0180_));
 sg13g2_nand2b_1 _1090_ (.Y(_0182_),
    .B(_0181_),
    .A_N(_0104_));
 sg13g2_a21oi_1 _1091_ (.A1(_0159_),
    .A2(_0178_),
    .Y(_0183_),
    .B1(_0168_));
 sg13g2_nor2_2 _1092_ (.A(_0176_),
    .B(_0183_),
    .Y(_0184_));
 sg13g2_nor2_1 _1093_ (.A(_0145_),
    .B(_0161_),
    .Y(_0185_));
 sg13g2_nor2_2 _1094_ (.A(_0172_),
    .B(_0185_),
    .Y(_0186_));
 sg13g2_xnor2_1 _1095_ (.Y(_0187_),
    .A(_0184_),
    .B(_0186_));
 sg13g2_xor2_1 _1096_ (.B(_0187_),
    .A(_0181_),
    .X(_0188_));
 sg13g2_nor2_1 _1097_ (.A(_0142_),
    .B(_0188_),
    .Y(_0189_));
 sg13g2_xnor2_1 _1098_ (.Y(_0190_),
    .A(_0182_),
    .B(_0189_));
 sg13g2_nor2_1 _1099_ (.A(_0180_),
    .B(_0183_),
    .Y(_0191_));
 sg13g2_nor2_1 _1100_ (.A(_0176_),
    .B(_0191_),
    .Y(_0192_));
 sg13g2_nand2b_1 _1101_ (.Y(_0193_),
    .B(_0192_),
    .A_N(_0124_));
 sg13g2_nand2b_1 _1102_ (.Y(_0194_),
    .B(_0184_),
    .A_N(_0123_));
 sg13g2_xnor2_1 _1103_ (.Y(_0195_),
    .A(_0193_),
    .B(_0194_));
 sg13g2_xnor2_1 _1104_ (.Y(_0196_),
    .A(_0190_),
    .B(_0195_));
 sg13g2_nor2b_1 _1105_ (.A(_0110_),
    .B_N(_0174_),
    .Y(_0197_));
 sg13g2_o21ai_1 _1106_ (.B1(_0173_),
    .Y(_0198_),
    .A1(_0174_),
    .A2(_0185_));
 sg13g2_nand2_1 _1107_ (.Y(_0199_),
    .A(_0154_),
    .B(_0198_));
 sg13g2_xnor2_1 _1108_ (.Y(_0200_),
    .A(_0197_),
    .B(_0199_));
 sg13g2_nand2b_1 _1109_ (.Y(_0201_),
    .B(_0192_),
    .A_N(_0125_));
 sg13g2_o21ai_1 _1110_ (.B1(_0118_),
    .Y(_0202_),
    .A1(_0175_),
    .A2(_0179_));
 sg13g2_xor2_1 _1111_ (.B(_0202_),
    .A(_0201_),
    .X(_0203_));
 sg13g2_xor2_1 _1112_ (.B(_0203_),
    .A(_0200_),
    .X(_0204_));
 sg13g2_xor2_1 _1113_ (.B(_0204_),
    .A(_0196_),
    .X(_0205_));
 sg13g2_o21ai_1 _1114_ (.B1(_0093_),
    .Y(_0206_),
    .A1(net78),
    .A2(_0205_));
 sg13g2_nor2_2 _1115_ (.A(_0068_),
    .B(net84),
    .Y(_0207_));
 sg13g2_or2_1 _1116_ (.X(_0208_),
    .B(net84),
    .A(_0068_));
 sg13g2_and2_1 _1117_ (.A(net87),
    .B(_0109_),
    .X(_0209_));
 sg13g2_nand2_2 _1118_ (.Y(_0210_),
    .A(net86),
    .B(_0109_));
 sg13g2_and2_1 _1119_ (.A(net90),
    .B(_0094_),
    .X(_0211_));
 sg13g2_nand3_1 _1120_ (.B(_0109_),
    .C(_0112_),
    .A(net93),
    .Y(_0212_));
 sg13g2_nand2_1 _1121_ (.Y(_0213_),
    .A(net93),
    .B(_0111_));
 sg13g2_nor3_1 _1122_ (.A(_0067_),
    .B(_0109_),
    .C(_0112_),
    .Y(_0214_));
 sg13g2_nand3b_1 _1123_ (.B(_0111_),
    .C(net90),
    .Y(_0215_),
    .A_N(_0109_));
 sg13g2_nand2_2 _1124_ (.Y(_0216_),
    .A(_0212_),
    .B(_0215_));
 sg13g2_nor3_1 _1125_ (.A(_0067_),
    .B(_0106_),
    .C(_0115_),
    .Y(_0217_));
 sg13g2_nand3b_1 _1126_ (.B(_0105_),
    .C(net93),
    .Y(_0218_),
    .A_N(_0115_));
 sg13g2_and2_1 _1127_ (.A(net90),
    .B(_0115_),
    .X(_0219_));
 sg13g2_nand3_1 _1128_ (.B(_0106_),
    .C(_0115_),
    .A(net93),
    .Y(_0220_));
 sg13g2_a221oi_1 _1129_ (.B2(_0106_),
    .C1(_0217_),
    .B1(_0219_),
    .A1(_0212_),
    .Y(_0221_),
    .A2(_0215_));
 sg13g2_a221oi_1 _1130_ (.B2(_0220_),
    .C1(_0214_),
    .B1(_0218_),
    .A1(_0112_),
    .Y(_0222_),
    .A2(net70));
 sg13g2_or3_1 _1131_ (.A(_0211_),
    .B(_0221_),
    .C(_0222_),
    .X(_0223_));
 sg13g2_o21ai_1 _1132_ (.B1(_0211_),
    .Y(_0224_),
    .A1(_0221_),
    .A2(_0222_));
 sg13g2_nand2_2 _1133_ (.Y(_0225_),
    .A(_0223_),
    .B(_0224_));
 sg13g2_xnor2_1 _1134_ (.Y(_0226_),
    .A(net70),
    .B(_0225_));
 sg13g2_inv_1 _1135_ (.Y(_0227_),
    .A(_0226_));
 sg13g2_nand2b_2 _1136_ (.Y(_0228_),
    .B(net70),
    .A_N(_0102_));
 sg13g2_nand2_1 _1137_ (.Y(_0229_),
    .A(net87),
    .B(_0102_));
 sg13g2_nand3_1 _1138_ (.B(_0102_),
    .C(_0210_),
    .A(net86),
    .Y(_0230_));
 sg13g2_nand2_2 _1139_ (.Y(_0231_),
    .A(_0228_),
    .B(_0230_));
 sg13g2_inv_1 _1140_ (.Y(_0232_),
    .A(_0231_));
 sg13g2_nand2_1 _1141_ (.Y(_0233_),
    .A(net87),
    .B(_0096_));
 sg13g2_and2_1 _1142_ (.A(_0096_),
    .B(net70),
    .X(_0234_));
 sg13g2_nand2_1 _1143_ (.Y(_0235_),
    .A(_0096_),
    .B(net70));
 sg13g2_a21oi_1 _1144_ (.A1(net86),
    .A2(_0096_),
    .Y(_0236_),
    .B1(net70));
 sg13g2_a21o_2 _1145_ (.A2(_0096_),
    .A1(net87),
    .B1(_0209_),
    .X(_0237_));
 sg13g2_nand2_2 _1146_ (.Y(_0238_),
    .A(_0235_),
    .B(_0237_));
 sg13g2_nor2_1 _1147_ (.A(_0234_),
    .B(_0236_),
    .Y(_0239_));
 sg13g2_and2_1 _1148_ (.A(net86),
    .B(_0098_),
    .X(_0240_));
 sg13g2_nand2_1 _1149_ (.Y(_0241_),
    .A(net86),
    .B(_0098_));
 sg13g2_o21ai_1 _1150_ (.B1(_0240_),
    .Y(_0242_),
    .A1(_0234_),
    .A2(_0236_));
 sg13g2_nand3_1 _1151_ (.B(_0237_),
    .C(_0241_),
    .A(_0235_),
    .Y(_0243_));
 sg13g2_nand3_1 _1152_ (.B(_0237_),
    .C(_0240_),
    .A(_0235_),
    .Y(_0244_));
 sg13g2_o21ai_1 _1153_ (.B1(_0241_),
    .Y(_0245_),
    .A1(_0234_),
    .A2(_0236_));
 sg13g2_nand2_2 _1154_ (.Y(_0246_),
    .A(_0244_),
    .B(_0245_));
 sg13g2_and4_1 _1155_ (.A(_0228_),
    .B(_0230_),
    .C(_0244_),
    .D(_0245_),
    .X(_0247_));
 sg13g2_a22oi_1 _1156_ (.Y(_0248_),
    .B1(_0244_),
    .B2(_0245_),
    .A2(_0230_),
    .A1(_0228_));
 sg13g2_and4_1 _1157_ (.A(_0228_),
    .B(_0230_),
    .C(_0242_),
    .D(_0243_),
    .X(_0249_));
 sg13g2_a22oi_1 _1158_ (.Y(_0250_),
    .B1(_0242_),
    .B2(_0243_),
    .A2(_0230_),
    .A1(_0228_));
 sg13g2_nor2_2 _1159_ (.A(_0249_),
    .B(_0250_),
    .Y(_0251_));
 sg13g2_and2_1 _1160_ (.A(_0226_),
    .B(_0251_),
    .X(_0252_));
 sg13g2_nand3b_1 _1161_ (.B(_0105_),
    .C(net86),
    .Y(_0253_),
    .A_N(_0098_));
 sg13g2_o21ai_1 _1162_ (.B1(_0253_),
    .Y(_0254_),
    .A1(_0105_),
    .A2(_0241_));
 sg13g2_nor3_1 _1163_ (.A(_0249_),
    .B(_0250_),
    .C(net69),
    .Y(_0255_));
 sg13g2_or3_1 _1164_ (.A(_0249_),
    .B(_0250_),
    .C(net69),
    .X(_0256_));
 sg13g2_o21ai_1 _1165_ (.B1(net69),
    .Y(_0257_),
    .A1(_0249_),
    .A2(_0250_));
 sg13g2_nand2_1 _1166_ (.Y(_0258_),
    .A(_0256_),
    .B(_0257_));
 sg13g2_xnor2_1 _1167_ (.Y(_0259_),
    .A(_0216_),
    .B(_0219_));
 sg13g2_inv_1 _1168_ (.Y(_0260_),
    .A(_0259_));
 sg13g2_nor3_1 _1169_ (.A(_0247_),
    .B(_0248_),
    .C(_0260_),
    .Y(_0261_));
 sg13g2_o21ai_1 _1170_ (.B1(_0259_),
    .Y(_0262_),
    .A1(_0249_),
    .A2(_0250_));
 sg13g2_nor3_1 _1171_ (.A(_0249_),
    .B(_0250_),
    .C(_0259_),
    .Y(_0263_));
 sg13g2_o21ai_1 _1172_ (.B1(_0260_),
    .Y(_0264_),
    .A1(_0247_),
    .A2(_0248_));
 sg13g2_nand2_2 _1173_ (.Y(_0265_),
    .A(_0262_),
    .B(_0264_));
 sg13g2_nor3_2 _1174_ (.A(_0239_),
    .B(_0261_),
    .C(_0263_),
    .Y(_0266_));
 sg13g2_nand3_1 _1175_ (.B(_0262_),
    .C(_0264_),
    .A(_0238_),
    .Y(_0267_));
 sg13g2_a21oi_2 _1176_ (.B1(_0238_),
    .Y(_0268_),
    .A2(_0264_),
    .A1(_0262_));
 sg13g2_o21ai_1 _1177_ (.B1(_0239_),
    .Y(_0269_),
    .A1(_0261_),
    .A2(_0263_));
 sg13g2_nor2_1 _1178_ (.A(_0266_),
    .B(_0268_),
    .Y(_0270_));
 sg13g2_nor3_1 _1179_ (.A(_0227_),
    .B(_0266_),
    .C(_0268_),
    .Y(_0271_));
 sg13g2_nand3_1 _1180_ (.B(_0267_),
    .C(_0269_),
    .A(_0226_),
    .Y(_0272_));
 sg13g2_o21ai_1 _1181_ (.B1(_0227_),
    .Y(_0273_),
    .A1(_0266_),
    .A2(_0268_));
 sg13g2_nand2_1 _1182_ (.Y(_0274_),
    .A(_0272_),
    .B(_0273_));
 sg13g2_a22oi_1 _1183_ (.Y(_0275_),
    .B1(_0272_),
    .B2(_0273_),
    .A2(_0257_),
    .A1(_0256_));
 sg13g2_nand2_1 _1184_ (.Y(_0276_),
    .A(_0255_),
    .B(_0271_));
 sg13g2_o21ai_1 _1185_ (.B1(_0276_),
    .Y(_0277_),
    .A1(_0252_),
    .A2(_0275_));
 sg13g2_and2_1 _1186_ (.A(net92),
    .B(\mask_i[7] ),
    .X(_0278_));
 sg13g2_nand3b_1 _1187_ (.B(\mask_i[7] ),
    .C(net92),
    .Y(_0279_),
    .A_N(\mask_i[4] ));
 sg13g2_and2_1 _1188_ (.A(net92),
    .B(\mask_i[4] ),
    .X(_0280_));
 sg13g2_nand2_1 _1189_ (.Y(_0281_),
    .A(net92),
    .B(\mask_i[4] ));
 sg13g2_o21ai_1 _1190_ (.B1(_0279_),
    .Y(_0282_),
    .A1(\mask_i[7] ),
    .A2(_0281_));
 sg13g2_nand2_1 _1191_ (.Y(_0283_),
    .A(_0226_),
    .B(_0282_));
 sg13g2_nand2_2 _1192_ (.Y(_0284_),
    .A(net92),
    .B(\mask_i[0] ));
 sg13g2_inv_2 _1193_ (.Y(_0285_),
    .A(_0284_));
 sg13g2_nand2_2 _1194_ (.Y(_0286_),
    .A(net92),
    .B(\mask_i[1] ));
 sg13g2_nand3b_1 _1195_ (.B(\mask_i[1] ),
    .C(net92),
    .Y(_0287_),
    .A_N(\mask_i[0] ));
 sg13g2_o21ai_1 _1196_ (.B1(_0287_),
    .Y(_0288_),
    .A1(\mask_i[1] ),
    .A2(_0284_));
 sg13g2_xnor2_1 _1197_ (.Y(_0289_),
    .A(\mask_i[6] ),
    .B(\mask_i[5] ));
 sg13g2_or2_1 _1198_ (.X(_0290_),
    .B(_0289_),
    .A(_0067_));
 sg13g2_xor2_1 _1199_ (.B(_0290_),
    .A(_0288_),
    .X(_0291_));
 sg13g2_nand2_1 _1200_ (.Y(_0292_),
    .A(net93),
    .B(\mask_i[2] ));
 sg13g2_xor2_1 _1201_ (.B(_0292_),
    .A(_0288_),
    .X(_0293_));
 sg13g2_nor3_1 _1202_ (.A(_0067_),
    .B(\mask_i[7] ),
    .C(_0289_),
    .Y(_0294_));
 sg13g2_a21oi_1 _1203_ (.A1(_0278_),
    .A2(_0289_),
    .Y(_0295_),
    .B1(_0294_));
 sg13g2_xnor2_1 _1204_ (.Y(_0296_),
    .A(_0293_),
    .B(_0295_));
 sg13g2_xnor2_1 _1205_ (.Y(_0297_),
    .A(_0291_),
    .B(net68));
 sg13g2_and2_1 _1206_ (.A(_0282_),
    .B(_0297_),
    .X(_0298_));
 sg13g2_xor2_1 _1207_ (.B(_0297_),
    .A(_0282_),
    .X(_0299_));
 sg13g2_xnor2_1 _1208_ (.Y(_0300_),
    .A(_0282_),
    .B(_0297_));
 sg13g2_a21o_1 _1209_ (.A2(_0273_),
    .A1(_0272_),
    .B1(_0299_),
    .X(_0301_));
 sg13g2_a22oi_1 _1210_ (.Y(_0302_),
    .B1(_0301_),
    .B2(_0283_),
    .A2(_0298_),
    .A1(_0271_));
 sg13g2_xnor2_1 _1211_ (.Y(_0303_),
    .A(_0277_),
    .B(_0302_));
 sg13g2_nand3_1 _1212_ (.B(_0224_),
    .C(_0238_),
    .A(_0223_),
    .Y(_0304_));
 sg13g2_a21o_1 _1213_ (.A2(_0224_),
    .A1(_0223_),
    .B1(_0238_),
    .X(_0305_));
 sg13g2_nand2_1 _1214_ (.Y(_0306_),
    .A(_0304_),
    .B(_0305_));
 sg13g2_xnor2_1 _1215_ (.Y(_0307_),
    .A(_0284_),
    .B(_0295_));
 sg13g2_inv_1 _1216_ (.Y(_0308_),
    .A(_0307_));
 sg13g2_xor2_1 _1217_ (.B(_0307_),
    .A(_0291_),
    .X(_0309_));
 sg13g2_nand2_1 _1218_ (.Y(_0310_),
    .A(_0306_),
    .B(_0309_));
 sg13g2_xnor2_1 _1219_ (.Y(_0311_),
    .A(\mask_i[6] ),
    .B(\mask_i[3] ));
 sg13g2_nor2_1 _1220_ (.A(_0067_),
    .B(_0311_),
    .Y(_0312_));
 sg13g2_xnor2_1 _1221_ (.Y(_0313_),
    .A(_0293_),
    .B(_0312_));
 sg13g2_nor2_1 _1222_ (.A(_0308_),
    .B(_0313_),
    .Y(_0314_));
 sg13g2_nor2_1 _1223_ (.A(\mask_i[0] ),
    .B(_0290_),
    .Y(_0315_));
 sg13g2_a21oi_2 _1224_ (.B1(_0315_),
    .Y(_0316_),
    .A2(_0289_),
    .A1(_0285_));
 sg13g2_a22oi_1 _1225_ (.Y(_0317_),
    .B1(_0316_),
    .B2(_0308_),
    .A2(_0313_),
    .A1(_0291_));
 sg13g2_nand4_1 _1226_ (.B(_0308_),
    .C(_0313_),
    .A(_0291_),
    .Y(_0318_),
    .D(_0316_));
 sg13g2_nor2b_1 _1227_ (.A(_0317_),
    .B_N(_0318_),
    .Y(_0319_));
 sg13g2_inv_1 _1228_ (.Y(_0320_),
    .A(_0319_));
 sg13g2_nor2_1 _1229_ (.A(_0314_),
    .B(_0319_),
    .Y(_0321_));
 sg13g2_nor2_1 _1230_ (.A(_0238_),
    .B(_0291_),
    .Y(_0322_));
 sg13g2_nand2_2 _1231_ (.Y(_0323_),
    .A(net91),
    .B(\prd_i[11] ));
 sg13g2_nand2b_1 _1232_ (.Y(_0324_),
    .B(_0112_),
    .A_N(_0323_));
 sg13g2_o21ai_1 _1233_ (.B1(_0324_),
    .Y(_0325_),
    .A1(\prd_i[11] ),
    .A2(_0213_));
 sg13g2_xor2_1 _1234_ (.B(_0325_),
    .A(_0322_),
    .X(_0326_));
 sg13g2_xor2_1 _1235_ (.B(_0321_),
    .A(_0310_),
    .X(_0327_));
 sg13g2_xnor2_1 _1236_ (.Y(_0328_),
    .A(_0326_),
    .B(_0327_));
 sg13g2_xor2_1 _1237_ (.B(_0233_),
    .A(_0216_),
    .X(_0329_));
 sg13g2_xnor2_1 _1238_ (.Y(_0330_),
    .A(_0216_),
    .B(_0233_));
 sg13g2_nor2_1 _1239_ (.A(_0238_),
    .B(_0329_),
    .Y(_0331_));
 sg13g2_nand3_1 _1240_ (.B(_0245_),
    .C(_0329_),
    .A(_0244_),
    .Y(_0332_));
 sg13g2_nand3_1 _1241_ (.B(_0243_),
    .C(_0330_),
    .A(_0242_),
    .Y(_0333_));
 sg13g2_nand2_2 _1242_ (.Y(_0334_),
    .A(_0332_),
    .B(_0333_));
 sg13g2_a22oi_1 _1243_ (.Y(_0335_),
    .B1(_0332_),
    .B2(_0333_),
    .A2(_0305_),
    .A1(_0304_));
 sg13g2_nand2_1 _1244_ (.Y(_0336_),
    .A(_0225_),
    .B(_0246_));
 sg13g2_mux2_1 _1245_ (.A0(_0335_),
    .A1(_0336_),
    .S(_0331_),
    .X(_0337_));
 sg13g2_xor2_1 _1246_ (.B(_0313_),
    .A(_0307_),
    .X(_0338_));
 sg13g2_xor2_1 _1247_ (.B(_0338_),
    .A(_0286_),
    .X(_0339_));
 sg13g2_xnor2_1 _1248_ (.Y(_0340_),
    .A(_0337_),
    .B(_0339_));
 sg13g2_xnor2_1 _1249_ (.Y(_0341_),
    .A(_0284_),
    .B(_0313_));
 sg13g2_nand2_1 _1250_ (.Y(_0342_),
    .A(_0282_),
    .B(net66));
 sg13g2_nand2_1 _1251_ (.Y(_0343_),
    .A(net92),
    .B(\mask_i[3] ));
 sg13g2_xnor2_1 _1252_ (.Y(_0344_),
    .A(_0282_),
    .B(_0288_));
 sg13g2_xnor2_1 _1253_ (.Y(_0345_),
    .A(_0343_),
    .B(_0344_));
 sg13g2_xor2_1 _1254_ (.B(net67),
    .A(_0316_),
    .X(_0346_));
 sg13g2_nor2b_2 _1255_ (.A(_0346_),
    .B_N(net66),
    .Y(_0347_));
 sg13g2_xnor2_1 _1256_ (.Y(_0348_),
    .A(net66),
    .B(_0346_));
 sg13g2_xor2_1 _1257_ (.B(_0346_),
    .A(net66),
    .X(_0349_));
 sg13g2_o21ai_1 _1258_ (.B1(_0342_),
    .Y(_0350_),
    .A1(_0299_),
    .A2(_0348_));
 sg13g2_nand2_2 _1259_ (.Y(_0351_),
    .A(_0298_),
    .B(_0347_));
 sg13g2_and2_1 _1260_ (.A(_0350_),
    .B(_0351_),
    .X(_0352_));
 sg13g2_nor2_1 _1261_ (.A(_0225_),
    .B(_0246_),
    .Y(_0353_));
 sg13g2_xnor2_1 _1262_ (.Y(_0354_),
    .A(_0225_),
    .B(_0246_));
 sg13g2_inv_1 _1263_ (.Y(_0355_),
    .A(_0354_));
 sg13g2_nand3_1 _1264_ (.B(_0351_),
    .C(_0355_),
    .A(_0350_),
    .Y(_0356_));
 sg13g2_a21o_1 _1265_ (.A2(_0351_),
    .A1(_0350_),
    .B1(_0355_),
    .X(_0357_));
 sg13g2_and3_1 _1266_ (.X(_0358_),
    .A(_0340_),
    .B(_0356_),
    .C(_0357_));
 sg13g2_a21oi_1 _1267_ (.A1(_0356_),
    .A2(_0357_),
    .Y(_0359_),
    .B1(_0340_));
 sg13g2_and2_1 _1268_ (.A(_0251_),
    .B(net66),
    .X(_0360_));
 sg13g2_a21oi_1 _1269_ (.A1(_0256_),
    .A2(_0257_),
    .Y(_0361_),
    .B1(_0348_));
 sg13g2_nand2_1 _1270_ (.Y(_0362_),
    .A(_0255_),
    .B(_0347_));
 sg13g2_o21ai_1 _1271_ (.B1(_0362_),
    .Y(_0363_),
    .A1(_0360_),
    .A2(_0361_));
 sg13g2_xnor2_1 _1272_ (.Y(_0364_),
    .A(_0313_),
    .B(_0316_));
 sg13g2_and2_1 _1273_ (.A(_0334_),
    .B(_0364_),
    .X(_0365_));
 sg13g2_nor2_1 _1274_ (.A(_0316_),
    .B(_0329_),
    .Y(_0366_));
 sg13g2_xnor2_1 _1275_ (.Y(_0367_),
    .A(_0365_),
    .B(_0366_));
 sg13g2_xnor2_1 _1276_ (.Y(_0368_),
    .A(_0363_),
    .B(_0367_));
 sg13g2_or3_1 _1277_ (.A(_0358_),
    .B(_0359_),
    .C(_0368_),
    .X(_0369_));
 sg13g2_o21ai_1 _1278_ (.B1(_0368_),
    .Y(_0370_),
    .A1(_0358_),
    .A2(_0359_));
 sg13g2_nand3_1 _1279_ (.B(_0369_),
    .C(_0370_),
    .A(_0328_),
    .Y(_0371_));
 sg13g2_a21o_1 _1280_ (.A2(_0370_),
    .A1(_0369_),
    .B1(_0328_),
    .X(_0372_));
 sg13g2_nand3_1 _1281_ (.B(_0371_),
    .C(_0372_),
    .A(_0303_),
    .Y(_0373_));
 sg13g2_a21o_2 _1282_ (.A2(_0372_),
    .A1(_0371_),
    .B1(_0303_),
    .X(_0374_));
 sg13g2_and2_1 _1283_ (.A(_0373_),
    .B(_0374_),
    .X(_0375_));
 sg13g2_nand2_1 _1284_ (.Y(_0376_),
    .A(_0373_),
    .B(_0374_));
 sg13g2_nor2b_1 _1285_ (.A(_0297_),
    .B_N(_0346_),
    .Y(_0377_));
 sg13g2_xnor2_1 _1286_ (.Y(_0378_),
    .A(_0342_),
    .B(_0377_));
 sg13g2_nand2_2 _1287_ (.Y(_0379_),
    .A(net91),
    .B(\prd_i[10] ));
 sg13g2_xnor2_1 _1288_ (.Y(_0380_),
    .A(_0354_),
    .B(_0379_));
 sg13g2_xnor2_1 _1289_ (.Y(_0381_),
    .A(_0378_),
    .B(_0380_));
 sg13g2_a21oi_1 _1290_ (.A1(_0267_),
    .A2(_0269_),
    .Y(_0382_),
    .B1(_0297_));
 sg13g2_xnor2_1 _1291_ (.Y(_0383_),
    .A(_0283_),
    .B(_0382_));
 sg13g2_o21ai_1 _1292_ (.B1(net69),
    .Y(_0384_),
    .A1(_0266_),
    .A2(_0268_));
 sg13g2_xor2_1 _1293_ (.B(_0384_),
    .A(_0252_),
    .X(_0385_));
 sg13g2_o21ai_1 _1294_ (.B1(_0320_),
    .Y(_0386_),
    .A1(_0291_),
    .A2(_0316_));
 sg13g2_xnor2_1 _1295_ (.Y(_0387_),
    .A(_0381_),
    .B(_0385_));
 sg13g2_xor2_1 _1296_ (.B(_0386_),
    .A(_0383_),
    .X(_0388_));
 sg13g2_xnor2_1 _1297_ (.Y(_0389_),
    .A(_0387_),
    .B(_0388_));
 sg13g2_or2_1 _1298_ (.X(_0390_),
    .B(_0332_),
    .A(_0304_));
 sg13g2_o21ai_1 _1299_ (.B1(_0390_),
    .Y(_0391_),
    .A1(_0335_),
    .A2(_0353_));
 sg13g2_nor2_1 _1300_ (.A(_0225_),
    .B(_0307_),
    .Y(_0392_));
 sg13g2_xnor2_1 _1301_ (.Y(_0393_),
    .A(_0310_),
    .B(_0392_));
 sg13g2_xnor2_1 _1302_ (.Y(_0394_),
    .A(_0391_),
    .B(_0393_));
 sg13g2_nand2_1 _1303_ (.Y(_0395_),
    .A(net69),
    .B(_0346_));
 sg13g2_xor2_1 _1304_ (.B(_0395_),
    .A(_0360_),
    .X(_0396_));
 sg13g2_nand3_1 _1305_ (.B(_0245_),
    .C(_0313_),
    .A(_0244_),
    .Y(_0397_));
 sg13g2_xnor2_1 _1306_ (.Y(_0398_),
    .A(_0365_),
    .B(_0397_));
 sg13g2_xnor2_1 _1307_ (.Y(_0399_),
    .A(_0396_),
    .B(_0398_));
 sg13g2_xnor2_1 _1308_ (.Y(_0400_),
    .A(_0394_),
    .B(_0399_));
 sg13g2_xnor2_1 _1309_ (.Y(_0401_),
    .A(_0389_),
    .B(_0400_));
 sg13g2_xor2_1 _1310_ (.B(_0400_),
    .A(_0389_),
    .X(_0402_));
 sg13g2_a21oi_1 _1311_ (.A1(_0373_),
    .A2(_0374_),
    .Y(_0403_),
    .B1(_0401_));
 sg13g2_nand3_1 _1312_ (.B(_0374_),
    .C(_0401_),
    .A(_0373_),
    .Y(_0404_));
 sg13g2_nor2b_1 _1313_ (.A(_0403_),
    .B_N(_0404_),
    .Y(_0405_));
 sg13g2_or2_1 _1314_ (.X(_0406_),
    .B(_0323_),
    .A(\prd_i[10] ));
 sg13g2_o21ai_1 _1315_ (.B1(_0406_),
    .Y(_0407_),
    .A1(\prd_i[11] ),
    .A2(_0379_));
 sg13g2_nand2_2 _1316_ (.Y(_0408_),
    .A(net91),
    .B(\prd_i[12] ));
 sg13g2_or2_1 _1317_ (.X(_0409_),
    .B(_0408_),
    .A(\prd_i[13] ));
 sg13g2_nand2_2 _1318_ (.Y(_0410_),
    .A(net91),
    .B(\prd_i[13] ));
 sg13g2_o21ai_1 _1319_ (.B1(_0409_),
    .Y(_0411_),
    .A1(\prd_i[12] ),
    .A2(_0410_));
 sg13g2_nor2_1 _1320_ (.A(\mask_i[4] ),
    .B(_0290_),
    .Y(_0412_));
 sg13g2_a21oi_2 _1321_ (.B1(_0412_),
    .Y(_0413_),
    .A2(_0289_),
    .A1(_0280_));
 sg13g2_nand2_1 _1322_ (.Y(_0414_),
    .A(_0285_),
    .B(_0413_));
 sg13g2_nor2_1 _1323_ (.A(_0285_),
    .B(net67),
    .Y(_0415_));
 sg13g2_nand2_1 _1324_ (.Y(_0416_),
    .A(_0285_),
    .B(net67));
 sg13g2_nand2b_2 _1325_ (.Y(_0417_),
    .B(_0416_),
    .A_N(_0415_));
 sg13g2_xnor2_1 _1326_ (.Y(_0418_),
    .A(_0284_),
    .B(_0413_));
 sg13g2_xnor2_1 _1327_ (.Y(_0419_),
    .A(net68),
    .B(_0418_));
 sg13g2_xor2_1 _1328_ (.B(_0418_),
    .A(net68),
    .X(_0420_));
 sg13g2_and2_1 _1329_ (.A(_0417_),
    .B(_0420_),
    .X(_0421_));
 sg13g2_a21oi_1 _1330_ (.A1(_0296_),
    .A2(net67),
    .Y(_0422_),
    .B1(_0414_));
 sg13g2_a21o_1 _1331_ (.A2(_0421_),
    .A1(_0414_),
    .B1(_0422_),
    .X(_0423_));
 sg13g2_xnor2_1 _1332_ (.Y(_0424_),
    .A(net69),
    .B(_0330_));
 sg13g2_xnor2_1 _1333_ (.Y(_0425_),
    .A(_0254_),
    .B(_0329_));
 sg13g2_nand2_1 _1334_ (.Y(_0426_),
    .A(_0231_),
    .B(_0424_));
 sg13g2_nor2_1 _1335_ (.A(_0231_),
    .B(_0424_),
    .Y(_0427_));
 sg13g2_xnor2_1 _1336_ (.Y(_0428_),
    .A(_0231_),
    .B(_0425_));
 sg13g2_xnor2_1 _1337_ (.Y(_0429_),
    .A(_0231_),
    .B(_0424_));
 sg13g2_nand2_1 _1338_ (.Y(_0430_),
    .A(_0417_),
    .B(_0429_));
 sg13g2_o21ai_1 _1339_ (.B1(_0430_),
    .Y(_0431_),
    .A1(_0232_),
    .A2(_0284_));
 sg13g2_o21ai_1 _1340_ (.B1(_0431_),
    .Y(_0432_),
    .A1(_0416_),
    .A2(_0426_));
 sg13g2_xor2_1 _1341_ (.B(_0423_),
    .A(_0385_),
    .X(_0433_));
 sg13g2_xor2_1 _1342_ (.B(_0432_),
    .A(_0383_),
    .X(_0434_));
 sg13g2_xnor2_1 _1343_ (.Y(_0435_),
    .A(_0433_),
    .B(_0434_));
 sg13g2_nor2_1 _1344_ (.A(_0265_),
    .B(_0424_),
    .Y(_0436_));
 sg13g2_nand2_1 _1345_ (.Y(_0437_),
    .A(_0265_),
    .B(_0424_));
 sg13g2_nand2b_1 _1346_ (.Y(_0438_),
    .B(_0437_),
    .A_N(_0436_));
 sg13g2_nor2_1 _1347_ (.A(_0210_),
    .B(_0418_),
    .Y(_0439_));
 sg13g2_xnor2_1 _1348_ (.Y(_0440_),
    .A(_0396_),
    .B(_0439_));
 sg13g2_xnor2_1 _1349_ (.Y(_0441_),
    .A(_0438_),
    .B(_0440_));
 sg13g2_nand3_1 _1350_ (.B(_0262_),
    .C(_0264_),
    .A(_0210_),
    .Y(_0442_));
 sg13g2_o21ai_1 _1351_ (.B1(net70),
    .Y(_0443_),
    .A1(_0261_),
    .A2(_0263_));
 sg13g2_and2_1 _1352_ (.A(_0442_),
    .B(_0443_),
    .X(_0444_));
 sg13g2_nor2_1 _1353_ (.A(_0419_),
    .B(_0444_),
    .Y(_0445_));
 sg13g2_nor2_1 _1354_ (.A(net68),
    .B(net67),
    .Y(_0446_));
 sg13g2_xor2_1 _1355_ (.B(_0345_),
    .A(_0296_),
    .X(_0447_));
 sg13g2_nand2b_1 _1356_ (.Y(_0448_),
    .B(_0112_),
    .A_N(_0408_));
 sg13g2_o21ai_1 _1357_ (.B1(_0448_),
    .Y(_0449_),
    .A1(\prd_i[12] ),
    .A2(_0213_));
 sg13g2_xnor2_1 _1358_ (.Y(_0450_),
    .A(_0447_),
    .B(_0449_));
 sg13g2_xnor2_1 _1359_ (.Y(_0451_),
    .A(_0378_),
    .B(_0450_));
 sg13g2_xnor2_1 _1360_ (.Y(_0452_),
    .A(_0286_),
    .B(_0451_));
 sg13g2_xnor2_1 _1361_ (.Y(_0453_),
    .A(_0445_),
    .B(_0452_));
 sg13g2_xnor2_1 _1362_ (.Y(_0454_),
    .A(_0441_),
    .B(_0453_));
 sg13g2_a21oi_1 _1363_ (.A1(_0442_),
    .A2(_0443_),
    .Y(_0455_),
    .B1(_0428_));
 sg13g2_mux2_1 _1364_ (.A0(_0437_),
    .A1(_0455_),
    .S(_0228_),
    .X(_0456_));
 sg13g2_xnor2_1 _1365_ (.Y(_0457_),
    .A(_0435_),
    .B(_0456_));
 sg13g2_xnor2_1 _1366_ (.Y(_0458_),
    .A(_0454_),
    .B(_0457_));
 sg13g2_nor2_1 _1367_ (.A(_0265_),
    .B(net68),
    .Y(_0459_));
 sg13g2_xnor2_1 _1368_ (.Y(_0460_),
    .A(_0445_),
    .B(_0459_));
 sg13g2_nand2b_1 _1369_ (.Y(_0461_),
    .B(_0425_),
    .A_N(net67));
 sg13g2_a22oi_1 _1370_ (.Y(_0462_),
    .B1(_0430_),
    .B2(_0461_),
    .A2(_0427_),
    .A1(_0415_));
 sg13g2_xnor2_1 _1371_ (.Y(_0463_),
    .A(_0460_),
    .B(_0462_));
 sg13g2_nand4_1 _1372_ (.B(_0262_),
    .C(_0264_),
    .A(_0210_),
    .Y(_0464_),
    .D(_0427_));
 sg13g2_o21ai_1 _1373_ (.B1(_0464_),
    .Y(_0465_),
    .A1(_0436_),
    .A2(_0455_));
 sg13g2_xnor2_1 _1374_ (.Y(_0466_),
    .A(_0363_),
    .B(_0465_));
 sg13g2_xor2_1 _1375_ (.B(_0413_),
    .A(_0410_),
    .X(_0467_));
 sg13g2_xnor2_1 _1376_ (.Y(_0468_),
    .A(_0229_),
    .B(_0338_));
 sg13g2_xnor2_1 _1377_ (.Y(_0469_),
    .A(_0354_),
    .B(_0467_));
 sg13g2_xnor2_1 _1378_ (.Y(_0470_),
    .A(_0468_),
    .B(_0469_));
 sg13g2_nand3b_1 _1379_ (.B(_0415_),
    .C(_0418_),
    .Y(_0471_),
    .A_N(net68));
 sg13g2_o21ai_1 _1380_ (.B1(_0471_),
    .Y(_0472_),
    .A1(_0421_),
    .A2(_0446_));
 sg13g2_xnor2_1 _1381_ (.Y(_0473_),
    .A(_0352_),
    .B(_0472_));
 sg13g2_xnor2_1 _1382_ (.Y(_0474_),
    .A(_0470_),
    .B(_0473_));
 sg13g2_xnor2_1 _1383_ (.Y(_0475_),
    .A(_0466_),
    .B(_0474_));
 sg13g2_xnor2_1 _1384_ (.Y(_0476_),
    .A(_0303_),
    .B(_0475_));
 sg13g2_xnor2_1 _1385_ (.Y(_0477_),
    .A(_0463_),
    .B(_0476_));
 sg13g2_xor2_1 _1386_ (.B(_0477_),
    .A(_0458_),
    .X(_0478_));
 sg13g2_xor2_1 _1387_ (.B(_0478_),
    .A(_0411_),
    .X(_0479_));
 sg13g2_nand2_1 _1388_ (.Y(_0480_),
    .A(_0407_),
    .B(_0479_));
 sg13g2_xnor2_1 _1389_ (.Y(_0481_),
    .A(\prd_i[12] ),
    .B(_0458_));
 sg13g2_nor2b_1 _1390_ (.A(_0379_),
    .B_N(_0481_),
    .Y(_0482_));
 sg13g2_xnor2_1 _1391_ (.Y(_0483_),
    .A(_0480_),
    .B(_0482_));
 sg13g2_nand2_1 _1392_ (.Y(_0484_),
    .A(_0402_),
    .B(_0408_));
 sg13g2_nand2_2 _1393_ (.Y(_0485_),
    .A(net91),
    .B(\prd_i[8] ));
 sg13g2_mux2_1 _1394_ (.A0(\prd_i[12] ),
    .A1(_0408_),
    .S(_0379_),
    .X(_0486_));
 sg13g2_nand3_1 _1395_ (.B(\prd_i[13] ),
    .C(\prd_i[11] ),
    .A(net91),
    .Y(_0487_));
 sg13g2_nand2_1 _1396_ (.Y(_0488_),
    .A(_0323_),
    .B(_0410_));
 sg13g2_nand2_1 _1397_ (.Y(_0489_),
    .A(_0487_),
    .B(_0488_));
 sg13g2_xnor2_1 _1398_ (.Y(_0490_),
    .A(_0486_),
    .B(_0489_));
 sg13g2_xnor2_1 _1399_ (.Y(_0491_),
    .A(_0485_),
    .B(_0490_));
 sg13g2_xnor2_1 _1400_ (.Y(_0492_),
    .A(_0458_),
    .B(_0491_));
 sg13g2_xnor2_1 _1401_ (.Y(_0493_),
    .A(_0484_),
    .B(_0492_));
 sg13g2_nand3b_1 _1402_ (.B(_0404_),
    .C(_0411_),
    .Y(_0494_),
    .A_N(_0403_));
 sg13g2_and2_1 _1403_ (.A(_0375_),
    .B(_0477_),
    .X(_0495_));
 sg13g2_nor2_1 _1404_ (.A(_0375_),
    .B(_0477_),
    .Y(_0496_));
 sg13g2_xnor2_1 _1405_ (.Y(_0497_),
    .A(_0376_),
    .B(_0477_));
 sg13g2_xnor2_1 _1406_ (.Y(_0498_),
    .A(_0494_),
    .B(_0497_));
 sg13g2_xnor2_1 _1407_ (.Y(_0499_),
    .A(_0493_),
    .B(_0498_));
 sg13g2_nor2_1 _1408_ (.A(_0401_),
    .B(_0458_),
    .Y(_0500_));
 sg13g2_nand2_1 _1409_ (.Y(_0501_),
    .A(_0405_),
    .B(_0478_));
 sg13g2_mux2_1 _1410_ (.A0(_0501_),
    .A1(_0495_),
    .S(_0500_),
    .X(_0502_));
 sg13g2_xor2_1 _1411_ (.B(_0502_),
    .A(_0499_),
    .X(_0503_));
 sg13g2_xnor2_1 _1412_ (.Y(_0504_),
    .A(_0483_),
    .B(_0503_));
 sg13g2_nand2_1 _1413_ (.Y(_0505_),
    .A(net91),
    .B(\prd_i[9] ));
 sg13g2_xor2_1 _1414_ (.B(_0505_),
    .A(_0489_),
    .X(_0506_));
 sg13g2_nand2_1 _1415_ (.Y(_0507_),
    .A(_0407_),
    .B(_0478_));
 sg13g2_xnor2_1 _1416_ (.Y(_0508_),
    .A(_0497_),
    .B(_0506_));
 sg13g2_xor2_1 _1417_ (.B(_0507_),
    .A(_0494_),
    .X(_0509_));
 sg13g2_xnor2_1 _1418_ (.Y(_0510_),
    .A(_0508_),
    .B(_0509_));
 sg13g2_and2_1 _1419_ (.A(_0401_),
    .B(_0458_),
    .X(_0511_));
 sg13g2_mux2_1 _1420_ (.A0(_0501_),
    .A1(_0511_),
    .S(_0496_),
    .X(_0512_));
 sg13g2_nor2_1 _1421_ (.A(_0323_),
    .B(_0477_),
    .Y(_0513_));
 sg13g2_nand2_1 _1422_ (.Y(_0514_),
    .A(_0407_),
    .B(_0411_));
 sg13g2_xor2_1 _1423_ (.B(_0514_),
    .A(_0487_),
    .X(_0515_));
 sg13g2_nor2_1 _1424_ (.A(_0375_),
    .B(_0410_),
    .Y(_0516_));
 sg13g2_xnor2_1 _1425_ (.Y(_0517_),
    .A(_0515_),
    .B(_0516_));
 sg13g2_xnor2_1 _1426_ (.Y(_0518_),
    .A(_0513_),
    .B(_0517_));
 sg13g2_xnor2_1 _1427_ (.Y(_0519_),
    .A(_0512_),
    .B(_0518_));
 sg13g2_xnor2_1 _1428_ (.Y(_0520_),
    .A(_0510_),
    .B(_0519_));
 sg13g2_xnor2_1 _1429_ (.Y(_0521_),
    .A(_0504_),
    .B(_0520_));
 sg13g2_nand2_1 _1430_ (.Y(_0522_),
    .A(_0405_),
    .B(_0521_));
 sg13g2_nor2_1 _1431_ (.A(_0401_),
    .B(_0520_),
    .Y(_0523_));
 sg13g2_nand2_2 _1432_ (.Y(_0524_),
    .A(net86),
    .B(\prd_i[16] ));
 sg13g2_or2_1 _1433_ (.X(_0525_),
    .B(_0485_),
    .A(\prd_i[9] ));
 sg13g2_o21ai_1 _1434_ (.B1(_0525_),
    .Y(_0526_),
    .A1(\prd_i[8] ),
    .A2(_0505_));
 sg13g2_nand2_1 _1435_ (.Y(_0527_),
    .A(_0405_),
    .B(_0526_));
 sg13g2_xnor2_1 _1436_ (.Y(_0528_),
    .A(_0524_),
    .B(_0527_));
 sg13g2_xnor2_1 _1437_ (.Y(_0529_),
    .A(_0523_),
    .B(_0528_));
 sg13g2_xnor2_1 _1438_ (.Y(_0530_),
    .A(_0522_),
    .B(_0529_));
 sg13g2_nand2_1 _1439_ (.Y(_0531_),
    .A(_0407_),
    .B(_0521_));
 sg13g2_nor2_1 _1440_ (.A(_0379_),
    .B(_0520_),
    .Y(_0532_));
 sg13g2_nand2_1 _1441_ (.Y(_0533_),
    .A(_0407_),
    .B(_0526_));
 sg13g2_xnor2_1 _1442_ (.Y(_0534_),
    .A(\prd_i[10] ),
    .B(_0402_));
 sg13g2_nor2_1 _1443_ (.A(_0505_),
    .B(_0534_),
    .Y(_0535_));
 sg13g2_xor2_1 _1444_ (.B(_0535_),
    .A(_0533_),
    .X(_0536_));
 sg13g2_xnor2_1 _1445_ (.Y(_0537_),
    .A(_0532_),
    .B(_0536_));
 sg13g2_xnor2_1 _1446_ (.Y(_0538_),
    .A(_0531_),
    .B(_0537_));
 sg13g2_xnor2_1 _1447_ (.Y(_0539_),
    .A(_0530_),
    .B(_0538_));
 sg13g2_nand2_1 _1448_ (.Y(_0540_),
    .A(_0376_),
    .B(_0504_));
 sg13g2_nor2_1 _1449_ (.A(_0375_),
    .B(_0485_),
    .Y(_0541_));
 sg13g2_nand2_2 _1450_ (.Y(_0542_),
    .A(net87),
    .B(\prd_i[17] ));
 sg13g2_xnor2_1 _1451_ (.Y(_0543_),
    .A(_0541_),
    .B(_0542_));
 sg13g2_xnor2_1 _1452_ (.Y(_0544_),
    .A(_0527_),
    .B(_0543_));
 sg13g2_xnor2_1 _1453_ (.Y(_0545_),
    .A(_0540_),
    .B(_0544_));
 sg13g2_or2_1 _1454_ (.X(_0546_),
    .B(_0533_),
    .A(_0521_));
 sg13g2_nand3_1 _1455_ (.B(_0521_),
    .C(_0533_),
    .A(_0407_),
    .Y(_0547_));
 sg13g2_xnor2_1 _1456_ (.Y(_0548_),
    .A(\prd_i[8] ),
    .B(_0504_));
 sg13g2_or2_1 _1457_ (.X(_0549_),
    .B(_0548_),
    .A(_0323_));
 sg13g2_a21oi_1 _1458_ (.A1(_0546_),
    .A2(_0547_),
    .Y(_0550_),
    .B1(_0549_));
 sg13g2_and3_1 _1459_ (.X(_0551_),
    .A(_0546_),
    .B(_0547_),
    .C(_0549_));
 sg13g2_xnor2_1 _1460_ (.Y(_0552_),
    .A(_0522_),
    .B(_0545_));
 sg13g2_o21ai_1 _1461_ (.B1(_0552_),
    .Y(_0553_),
    .A1(_0550_),
    .A2(_0551_));
 sg13g2_or3_1 _1462_ (.A(_0550_),
    .B(_0551_),
    .C(_0552_),
    .X(_0554_));
 sg13g2_and2_1 _1463_ (.A(_0553_),
    .B(_0554_),
    .X(_0555_));
 sg13g2_or2_1 _1464_ (.X(_0556_),
    .B(_0555_),
    .A(_0539_));
 sg13g2_nand2_1 _1465_ (.Y(_0557_),
    .A(_0539_),
    .B(_0555_));
 sg13g2_xnor2_1 _1466_ (.Y(_0558_),
    .A(_0417_),
    .B(_0444_));
 sg13g2_nand3_1 _1467_ (.B(_0557_),
    .C(_0558_),
    .A(_0556_),
    .Y(_0559_));
 sg13g2_or2_1 _1468_ (.X(_0560_),
    .B(_0542_),
    .A(\prd_i[16] ));
 sg13g2_or2_1 _1469_ (.X(_0561_),
    .B(_0524_),
    .A(\prd_i[17] ));
 sg13g2_and2_1 _1470_ (.A(_0560_),
    .B(_0561_),
    .X(_0562_));
 sg13g2_nand2_1 _1471_ (.Y(_0563_),
    .A(_0560_),
    .B(_0561_));
 sg13g2_nand2_1 _1472_ (.Y(_0564_),
    .A(_0417_),
    .B(_0563_));
 sg13g2_nand3_1 _1473_ (.B(\prd_i[16] ),
    .C(\mask_i[0] ),
    .A(net86),
    .Y(_0565_));
 sg13g2_xnor2_1 _1474_ (.Y(_0566_),
    .A(_0564_),
    .B(_0565_));
 sg13g2_nand2_2 _1475_ (.Y(_0567_),
    .A(net87),
    .B(\prd_i[14] ));
 sg13g2_or2_1 _1476_ (.X(_0568_),
    .B(_0524_),
    .A(\prd_i[14] ));
 sg13g2_o21ai_1 _1477_ (.B1(_0568_),
    .Y(_0569_),
    .A1(\prd_i[16] ),
    .A2(_0567_));
 sg13g2_nand2_1 _1478_ (.Y(_0570_),
    .A(_0341_),
    .B(_0569_));
 sg13g2_nand2_2 _1479_ (.Y(_0571_),
    .A(net87),
    .B(\prd_i[15] ));
 sg13g2_or2_1 _1480_ (.X(_0572_),
    .B(_0571_),
    .A(\prd_i[17] ));
 sg13g2_o21ai_1 _1481_ (.B1(_0572_),
    .Y(_0573_),
    .A1(\prd_i[15] ),
    .A2(_0542_));
 sg13g2_nand2_1 _1482_ (.Y(_0574_),
    .A(_0346_),
    .B(_0573_));
 sg13g2_xor2_1 _1483_ (.B(_0574_),
    .A(_0570_),
    .X(_0575_));
 sg13g2_xnor2_1 _1484_ (.Y(_0576_),
    .A(_0566_),
    .B(_0575_));
 sg13g2_nand2_1 _1485_ (.Y(_0577_),
    .A(_0226_),
    .B(_0569_));
 sg13g2_nor2b_1 _1486_ (.A(_0270_),
    .B_N(_0573_),
    .Y(_0578_));
 sg13g2_xnor2_1 _1487_ (.Y(_0579_),
    .A(_0577_),
    .B(_0578_));
 sg13g2_nor2_1 _1488_ (.A(_0444_),
    .B(_0562_),
    .Y(_0580_));
 sg13g2_nand2_1 _1489_ (.Y(_0581_),
    .A(\prd_i[16] ),
    .B(net70));
 sg13g2_nand2_2 _1490_ (.Y(_0582_),
    .A(net88),
    .B(\prd_i[4] ));
 sg13g2_inv_1 _1491_ (.Y(_0583_),
    .A(_0582_));
 sg13g2_or2_1 _1492_ (.X(_0584_),
    .B(_0582_),
    .A(\prd_i[6] ));
 sg13g2_nand2_2 _1493_ (.Y(_0585_),
    .A(net88),
    .B(\prd_i[6] ));
 sg13g2_o21ai_1 _1494_ (.B1(_0584_),
    .Y(_0586_),
    .A1(\prd_i[4] ),
    .A2(_0585_));
 sg13g2_nand2_1 _1495_ (.Y(_0587_),
    .A(net119),
    .B(net89));
 sg13g2_or2_1 _1496_ (.X(_0588_),
    .B(_0587_),
    .A(\prd_i[1] ));
 sg13g2_nand2_1 _1497_ (.Y(_0589_),
    .A(net88),
    .B(\prd_i[1] ));
 sg13g2_o21ai_1 _1498_ (.B1(_0588_),
    .Y(_0590_),
    .A1(\prd_i[0] ),
    .A2(_0589_));
 sg13g2_xor2_1 _1499_ (.B(_0590_),
    .A(_0586_),
    .X(_0591_));
 sg13g2_xor2_1 _1500_ (.B(_0591_),
    .A(_0581_),
    .X(_0592_));
 sg13g2_xnor2_1 _1501_ (.Y(_0593_),
    .A(_0580_),
    .B(_0592_));
 sg13g2_xnor2_1 _1502_ (.Y(_0594_),
    .A(_0579_),
    .B(_0593_));
 sg13g2_nor2_1 _1503_ (.A(_0284_),
    .B(_0539_),
    .Y(_0595_));
 sg13g2_nor2_1 _1504_ (.A(_0210_),
    .B(_0539_),
    .Y(_0596_));
 sg13g2_xnor2_1 _1505_ (.Y(_0597_),
    .A(_0576_),
    .B(_0595_));
 sg13g2_xnor2_1 _1506_ (.Y(_0598_),
    .A(_0594_),
    .B(_0596_));
 sg13g2_xnor2_1 _1507_ (.Y(_0599_),
    .A(_0559_),
    .B(_0598_));
 sg13g2_xnor2_1 _1508_ (.Y(_0600_),
    .A(_0597_),
    .B(_0599_));
 sg13g2_nand2_1 _1509_ (.Y(_0601_),
    .A(_0479_),
    .B(_0521_));
 sg13g2_nor2_1 _1510_ (.A(_0458_),
    .B(_0520_),
    .Y(_0602_));
 sg13g2_nand2_1 _1511_ (.Y(_0603_),
    .A(_0479_),
    .B(_0526_));
 sg13g2_nand3_1 _1512_ (.B(\prd_i[9] ),
    .C(_0481_),
    .A(net91),
    .Y(_0604_));
 sg13g2_xor2_1 _1513_ (.B(_0604_),
    .A(_0603_),
    .X(_0605_));
 sg13g2_nor2_1 _1514_ (.A(_0408_),
    .B(_0520_),
    .Y(_0606_));
 sg13g2_xor2_1 _1515_ (.B(_0602_),
    .A(_0567_),
    .X(_0607_));
 sg13g2_xnor2_1 _1516_ (.Y(_0608_),
    .A(_0605_),
    .B(_0606_));
 sg13g2_xnor2_1 _1517_ (.Y(_0609_),
    .A(_0607_),
    .B(_0608_));
 sg13g2_xnor2_1 _1518_ (.Y(_0610_),
    .A(_0601_),
    .B(_0609_));
 sg13g2_nor2_1 _1519_ (.A(_0410_),
    .B(_0548_),
    .Y(_0611_));
 sg13g2_nor2_1 _1520_ (.A(_0477_),
    .B(_0485_),
    .Y(_0612_));
 sg13g2_xnor2_1 _1521_ (.Y(_0613_),
    .A(_0571_),
    .B(_0612_));
 sg13g2_xor2_1 _1522_ (.B(_0613_),
    .A(_0603_),
    .X(_0614_));
 sg13g2_xnor2_1 _1523_ (.Y(_0615_),
    .A(_0611_),
    .B(_0614_));
 sg13g2_nor2b_1 _1524_ (.A(_0477_),
    .B_N(_0504_),
    .Y(_0616_));
 sg13g2_xnor2_1 _1525_ (.Y(_0617_),
    .A(_0601_),
    .B(_0616_));
 sg13g2_xor2_1 _1526_ (.B(_0617_),
    .A(_0615_),
    .X(_0618_));
 sg13g2_xnor2_1 _1527_ (.Y(_0619_),
    .A(_0615_),
    .B(_0617_));
 sg13g2_nand2b_1 _1528_ (.Y(_0620_),
    .B(_0619_),
    .A_N(net65));
 sg13g2_xnor2_1 _1529_ (.Y(_0621_),
    .A(net65),
    .B(_0618_));
 sg13g2_xor2_1 _1530_ (.B(_0364_),
    .A(_0306_),
    .X(_0622_));
 sg13g2_nand2_2 _1531_ (.Y(_0623_),
    .A(_0621_),
    .B(_0622_));
 sg13g2_xor2_1 _1532_ (.B(net65),
    .A(_0567_),
    .X(_0624_));
 sg13g2_nand2_1 _1533_ (.Y(_0625_),
    .A(_0313_),
    .B(_0624_));
 sg13g2_or2_1 _1534_ (.X(_0626_),
    .B(_0571_),
    .A(\prd_i[14] ));
 sg13g2_o21ai_1 _1535_ (.B1(_0626_),
    .Y(_0627_),
    .A1(\prd_i[15] ),
    .A2(_0567_));
 sg13g2_and2_1 _1536_ (.A(_0622_),
    .B(_0627_),
    .X(_0628_));
 sg13g2_nor2_1 _1537_ (.A(_0225_),
    .B(_0567_),
    .Y(_0629_));
 sg13g2_nand3b_1 _1538_ (.B(net88),
    .C(\prd_i[3] ),
    .Y(_0630_),
    .A_N(\prd_i[0] ));
 sg13g2_o21ai_1 _1539_ (.B1(_0630_),
    .Y(_0631_),
    .A1(\prd_i[3] ),
    .A2(_0587_));
 sg13g2_xor2_1 _1540_ (.B(_0631_),
    .A(_0585_),
    .X(_0632_));
 sg13g2_mux2_1 _1541_ (.A0(\prd_i[1] ),
    .A1(_0589_),
    .S(_0632_),
    .X(_0633_));
 sg13g2_xnor2_1 _1542_ (.Y(_0634_),
    .A(_0629_),
    .B(_0633_));
 sg13g2_xnor2_1 _1543_ (.Y(_0635_),
    .A(_0575_),
    .B(_0634_));
 sg13g2_xnor2_1 _1544_ (.Y(_0636_),
    .A(_0628_),
    .B(_0635_));
 sg13g2_xnor2_1 _1545_ (.Y(_0637_),
    .A(_0579_),
    .B(_0636_));
 sg13g2_nor2_1 _1546_ (.A(_0225_),
    .B(net65),
    .Y(_0638_));
 sg13g2_xnor2_1 _1547_ (.Y(_0639_),
    .A(_0637_),
    .B(_0638_));
 sg13g2_xnor2_1 _1548_ (.Y(_0640_),
    .A(_0625_),
    .B(_0639_));
 sg13g2_xnor2_1 _1549_ (.Y(_0641_),
    .A(_0623_),
    .B(_0640_));
 sg13g2_xnor2_1 _1550_ (.Y(_0642_),
    .A(_0539_),
    .B(net65));
 sg13g2_xor2_1 _1551_ (.B(net65),
    .A(_0539_),
    .X(_0643_));
 sg13g2_nand2_1 _1552_ (.Y(_0644_),
    .A(_0226_),
    .B(_0643_));
 sg13g2_a21o_2 _1553_ (.A2(_0554_),
    .A1(_0553_),
    .B1(_0619_),
    .X(_0645_));
 sg13g2_nand3_1 _1554_ (.B(_0554_),
    .C(_0619_),
    .A(_0553_),
    .Y(_0646_));
 sg13g2_nand2_1 _1555_ (.Y(_0647_),
    .A(_0645_),
    .B(_0646_));
 sg13g2_nand2_1 _1556_ (.Y(_0648_),
    .A(net66),
    .B(_0643_));
 sg13g2_nand3_1 _1557_ (.B(net66),
    .C(_0643_),
    .A(_0227_),
    .Y(_0649_));
 sg13g2_o21ai_1 _1558_ (.B1(_0649_),
    .Y(_0650_),
    .A1(net66),
    .A2(_0644_));
 sg13g2_xor2_1 _1559_ (.B(_0346_),
    .A(_0270_),
    .X(_0651_));
 sg13g2_nor2_1 _1560_ (.A(_0647_),
    .B(_0651_),
    .Y(_0652_));
 sg13g2_xor2_1 _1561_ (.B(_0652_),
    .A(_0650_),
    .X(_0653_));
 sg13g2_xnor2_1 _1562_ (.Y(_0654_),
    .A(_0600_),
    .B(_0653_));
 sg13g2_xor2_1 _1563_ (.B(_0653_),
    .A(_0641_),
    .X(_0655_));
 sg13g2_xnor2_1 _1564_ (.Y(_0656_),
    .A(_0600_),
    .B(_0641_));
 sg13g2_a21oi_2 _1565_ (.B1(_0642_),
    .Y(_0657_),
    .A2(_0646_),
    .A1(_0645_));
 sg13g2_nand2_1 _1566_ (.Y(_0658_),
    .A(_0251_),
    .B(_0643_));
 sg13g2_and3_2 _1567_ (.X(_0659_),
    .A(_0642_),
    .B(_0645_),
    .C(_0646_));
 sg13g2_o21ai_1 _1568_ (.B1(_0258_),
    .Y(_0660_),
    .A1(_0657_),
    .A2(_0659_));
 sg13g2_a22oi_1 _1569_ (.Y(_0661_),
    .B1(_0658_),
    .B2(_0660_),
    .A2(_0657_),
    .A1(_0255_));
 sg13g2_nand2_1 _1570_ (.Y(_0662_),
    .A(_0282_),
    .B(_0643_));
 sg13g2_o21ai_1 _1571_ (.B1(_0300_),
    .Y(_0663_),
    .A1(_0657_),
    .A2(_0659_));
 sg13g2_a22oi_1 _1572_ (.Y(_0664_),
    .B1(_0662_),
    .B2(_0663_),
    .A2(_0657_),
    .A1(_0298_));
 sg13g2_xnor2_1 _1573_ (.Y(_0665_),
    .A(_0661_),
    .B(_0664_));
 sg13g2_nand2_1 _1574_ (.Y(_0666_),
    .A(_0309_),
    .B(_0621_));
 sg13g2_nor2_1 _1575_ (.A(_0291_),
    .B(_0619_),
    .Y(_0667_));
 sg13g2_and2_1 _1576_ (.A(_0251_),
    .B(_0569_),
    .X(_0668_));
 sg13g2_xor2_1 _1577_ (.B(_0573_),
    .A(_0569_),
    .X(_0669_));
 sg13g2_nand2_1 _1578_ (.Y(_0670_),
    .A(_0258_),
    .B(_0669_));
 sg13g2_xor2_1 _1579_ (.B(_0670_),
    .A(_0668_),
    .X(_0671_));
 sg13g2_nand2_1 _1580_ (.Y(_0672_),
    .A(_0334_),
    .B(_0627_));
 sg13g2_nor2_1 _1581_ (.A(_0329_),
    .B(_0571_),
    .Y(_0673_));
 sg13g2_xnor2_1 _1582_ (.Y(_0674_),
    .A(_0672_),
    .B(_0673_));
 sg13g2_xnor2_1 _1583_ (.Y(_0675_),
    .A(_0671_),
    .B(_0674_));
 sg13g2_xnor2_1 _1584_ (.Y(_0676_),
    .A(_0667_),
    .B(_0675_));
 sg13g2_nor2_1 _1585_ (.A(_0291_),
    .B(_0571_),
    .Y(_0677_));
 sg13g2_nand2_1 _1586_ (.Y(_0678_),
    .A(_0309_),
    .B(_0627_));
 sg13g2_xnor2_1 _1587_ (.Y(_0679_),
    .A(_0582_),
    .B(_0631_));
 sg13g2_xnor2_1 _1588_ (.Y(_0680_),
    .A(_0678_),
    .B(_0679_));
 sg13g2_xnor2_1 _1589_ (.Y(_0681_),
    .A(_0677_),
    .B(_0680_));
 sg13g2_nor2b_1 _1590_ (.A(_0333_),
    .B_N(net65),
    .Y(_0682_));
 sg13g2_a22oi_1 _1591_ (.Y(_0683_),
    .B1(_0621_),
    .B2(_0334_),
    .A2(_0618_),
    .A1(_0330_));
 sg13g2_a21oi_1 _1592_ (.A1(_0618_),
    .A2(_0682_),
    .Y(_0684_),
    .B1(_0683_));
 sg13g2_nand2_1 _1593_ (.Y(_0685_),
    .A(_0282_),
    .B(_0569_));
 sg13g2_nand2_1 _1594_ (.Y(_0686_),
    .A(_0300_),
    .B(_0669_));
 sg13g2_xor2_1 _1595_ (.B(_0686_),
    .A(_0685_),
    .X(_0687_));
 sg13g2_xnor2_1 _1596_ (.Y(_0688_),
    .A(_0666_),
    .B(_0676_));
 sg13g2_xnor2_1 _1597_ (.Y(_0689_),
    .A(_0684_),
    .B(_0688_));
 sg13g2_xnor2_1 _1598_ (.Y(_0690_),
    .A(_0681_),
    .B(_0687_));
 sg13g2_xnor2_1 _1599_ (.Y(_0691_),
    .A(_0689_),
    .B(_0690_));
 sg13g2_xnor2_1 _1600_ (.Y(_0692_),
    .A(_0665_),
    .B(_0691_));
 sg13g2_xnor2_1 _1601_ (.Y(_0693_),
    .A(_0656_),
    .B(_0692_));
 sg13g2_nor2_2 _1602_ (.A(_0078_),
    .B(net84),
    .Y(_0694_));
 sg13g2_nor3_1 _1603_ (.A(_0078_),
    .B(net84),
    .C(_0587_),
    .Y(_0695_));
 sg13g2_a21oi_1 _1604_ (.A1(_0207_),
    .A2(_0693_),
    .Y(_0696_),
    .B1(_0695_));
 sg13g2_nand2_1 _1605_ (.Y(_0697_),
    .A(_0092_),
    .B(_0696_));
 sg13g2_a22oi_1 _1606_ (.Y(_0698_),
    .B1(_0206_),
    .B2(_0697_),
    .A2(net79),
    .A1(net138));
 sg13g2_nor2_1 _1607_ (.A(_0066_),
    .B(_0698_),
    .Y(_0016_));
 sg13g2_nand2b_2 _1608_ (.Y(_0699_),
    .B(_0181_),
    .A_N(_0132_));
 sg13g2_nor2_1 _1609_ (.A(_0135_),
    .B(_0187_),
    .Y(_0700_));
 sg13g2_xnor2_1 _1610_ (.Y(_0701_),
    .A(_0699_),
    .B(_0700_));
 sg13g2_xnor2_1 _1611_ (.Y(_0702_),
    .A(_0203_),
    .B(_0701_));
 sg13g2_o21ai_1 _1612_ (.B1(_0699_),
    .Y(_0703_),
    .A1(_0136_),
    .A2(_0188_));
 sg13g2_nand2_1 _1613_ (.Y(_0704_),
    .A(_0135_),
    .B(_0187_));
 sg13g2_o21ai_1 _1614_ (.B1(_0703_),
    .Y(_0705_),
    .A1(_0699_),
    .A2(_0704_));
 sg13g2_nand2_1 _1615_ (.Y(_0706_),
    .A(_0119_),
    .B(_0184_));
 sg13g2_xnor2_1 _1616_ (.Y(_0707_),
    .A(_0201_),
    .B(_0706_));
 sg13g2_xnor2_1 _1617_ (.Y(_0708_),
    .A(_0705_),
    .B(_0707_));
 sg13g2_xnor2_1 _1618_ (.Y(_0709_),
    .A(_0702_),
    .B(_0708_));
 sg13g2_xnor2_1 _1619_ (.Y(_0710_),
    .A(_0196_),
    .B(_0709_));
 sg13g2_o21ai_1 _1620_ (.B1(_0093_),
    .Y(_0711_),
    .A1(net78),
    .A2(_0710_));
 sg13g2_o21ai_1 _1621_ (.B1(_0274_),
    .Y(_0712_),
    .A1(_0657_),
    .A2(_0659_));
 sg13g2_a22oi_1 _1622_ (.Y(_0713_),
    .B1(_0712_),
    .B2(_0644_),
    .A2(_0657_),
    .A1(_0271_));
 sg13g2_o21ai_1 _1623_ (.B1(_0349_),
    .Y(_0714_),
    .A1(_0657_),
    .A2(_0659_));
 sg13g2_a22oi_1 _1624_ (.Y(_0715_),
    .B1(_0714_),
    .B2(_0648_),
    .A2(_0657_),
    .A1(_0347_));
 sg13g2_xnor2_1 _1625_ (.Y(_0716_),
    .A(_0713_),
    .B(_0715_));
 sg13g2_nand2_1 _1626_ (.Y(_0717_),
    .A(_0349_),
    .B(_0669_));
 sg13g2_xor2_1 _1627_ (.B(_0717_),
    .A(_0570_),
    .X(_0718_));
 sg13g2_nand2_1 _1628_ (.Y(_0719_),
    .A(_0274_),
    .B(_0669_));
 sg13g2_xor2_1 _1629_ (.B(_0719_),
    .A(_0577_),
    .X(_0720_));
 sg13g2_xnor2_1 _1630_ (.Y(_0721_),
    .A(_0718_),
    .B(_0720_));
 sg13g2_xnor2_1 _1631_ (.Y(_0722_),
    .A(_0238_),
    .B(_0316_));
 sg13g2_nor2_1 _1632_ (.A(_0571_),
    .B(_0722_),
    .Y(_0723_));
 sg13g2_xnor2_1 _1633_ (.Y(_0724_),
    .A(_0586_),
    .B(_0628_));
 sg13g2_xnor2_1 _1634_ (.Y(_0725_),
    .A(_0723_),
    .B(_0724_));
 sg13g2_xnor2_1 _1635_ (.Y(_0726_),
    .A(_0721_),
    .B(_0725_));
 sg13g2_nor2_1 _1636_ (.A(_0619_),
    .B(_0722_),
    .Y(_0727_));
 sg13g2_xnor2_1 _1637_ (.Y(_0728_),
    .A(_0726_),
    .B(_0727_));
 sg13g2_xnor2_1 _1638_ (.Y(_0729_),
    .A(_0623_),
    .B(_0728_));
 sg13g2_xnor2_1 _1639_ (.Y(_0730_),
    .A(_0716_),
    .B(_0729_));
 sg13g2_xnor2_1 _1640_ (.Y(_0731_),
    .A(_0655_),
    .B(_0730_));
 sg13g2_a21oi_1 _1641_ (.A1(_0692_),
    .A2(_0731_),
    .Y(_0732_),
    .B1(_0208_));
 sg13g2_o21ai_1 _1642_ (.B1(_0732_),
    .Y(_0733_),
    .A1(_0692_),
    .A2(_0731_));
 sg13g2_nand2b_1 _1643_ (.Y(_0734_),
    .B(_0694_),
    .A_N(_0589_));
 sg13g2_nand3_1 _1644_ (.B(_0733_),
    .C(_0734_),
    .A(_0092_),
    .Y(_0735_));
 sg13g2_a22oi_1 _1645_ (.Y(_0736_),
    .B1(_0711_),
    .B2(_0735_),
    .A2(net79),
    .A1(net137));
 sg13g2_nor2_1 _1646_ (.A(_0066_),
    .B(_0736_),
    .Y(_0017_));
 sg13g2_nand3_1 _1647_ (.B(_0556_),
    .C(_0557_),
    .A(_0420_),
    .Y(_0737_));
 sg13g2_nand4_1 _1648_ (.B(_0429_),
    .C(_0556_),
    .A(_0419_),
    .Y(_0738_),
    .D(_0557_));
 sg13g2_o21ai_1 _1649_ (.B1(_0738_),
    .Y(_0739_),
    .A1(_0429_),
    .A2(_0737_));
 sg13g2_xnor2_1 _1650_ (.Y(_0740_),
    .A(net68),
    .B(_0424_));
 sg13g2_nor2_1 _1651_ (.A(_0555_),
    .B(_0740_),
    .Y(_0741_));
 sg13g2_nand2_1 _1652_ (.Y(_0742_),
    .A(_0420_),
    .B(_0563_));
 sg13g2_nor2_1 _1653_ (.A(net68),
    .B(_0542_),
    .Y(_0743_));
 sg13g2_xor2_1 _1654_ (.B(_0743_),
    .A(_0742_),
    .X(_0744_));
 sg13g2_nor2_1 _1655_ (.A(_0424_),
    .B(_0542_),
    .Y(_0745_));
 sg13g2_nand2_1 _1656_ (.Y(_0746_),
    .A(net88),
    .B(\prd_i[7] ));
 sg13g2_or2_1 _1657_ (.X(_0747_),
    .B(_0746_),
    .A(\prd_i[4] ));
 sg13g2_o21ai_1 _1658_ (.B1(_0747_),
    .Y(_0748_),
    .A1(\prd_i[7] ),
    .A2(_0582_));
 sg13g2_xor2_1 _1659_ (.B(_0748_),
    .A(_0745_),
    .X(_0749_));
 sg13g2_nor2_1 _1660_ (.A(_0428_),
    .B(_0562_),
    .Y(_0750_));
 sg13g2_xnor2_1 _1661_ (.Y(_0751_),
    .A(_0749_),
    .B(_0750_));
 sg13g2_xnor2_1 _1662_ (.Y(_0752_),
    .A(_0687_),
    .B(_0751_));
 sg13g2_xnor2_1 _1663_ (.Y(_0753_),
    .A(_0585_),
    .B(_0671_));
 sg13g2_xnor2_1 _1664_ (.Y(_0754_),
    .A(_0752_),
    .B(_0753_));
 sg13g2_xnor2_1 _1665_ (.Y(_0755_),
    .A(_0744_),
    .B(_0754_));
 sg13g2_xnor2_1 _1666_ (.Y(_0756_),
    .A(_0741_),
    .B(_0755_));
 sg13g2_xnor2_1 _1667_ (.Y(_0757_),
    .A(_0739_),
    .B(_0756_));
 sg13g2_xnor2_1 _1668_ (.Y(_0758_),
    .A(_0665_),
    .B(_0757_));
 sg13g2_nand3_1 _1669_ (.B(_0645_),
    .C(_0646_),
    .A(net69),
    .Y(_0759_));
 sg13g2_xor2_1 _1670_ (.B(_0759_),
    .A(_0658_),
    .X(_0760_));
 sg13g2_or2_1 _1671_ (.X(_0761_),
    .B(_0678_),
    .A(_0621_));
 sg13g2_o21ai_1 _1672_ (.B1(_0761_),
    .Y(_0762_),
    .A1(_0627_),
    .A2(_0666_));
 sg13g2_nor2_1 _1673_ (.A(_0307_),
    .B(_0567_),
    .Y(_0763_));
 sg13g2_xor2_1 _1674_ (.B(_0763_),
    .A(_0591_),
    .X(_0764_));
 sg13g2_xnor2_1 _1675_ (.Y(_0765_),
    .A(_0762_),
    .B(_0764_));
 sg13g2_xnor2_1 _1676_ (.Y(_0766_),
    .A(_0760_),
    .B(_0765_));
 sg13g2_nor2_1 _1677_ (.A(_0297_),
    .B(_0647_),
    .Y(_0767_));
 sg13g2_xor2_1 _1678_ (.B(_0767_),
    .A(_0662_),
    .X(_0768_));
 sg13g2_nor2_1 _1679_ (.A(_0246_),
    .B(net65),
    .Y(_0769_));
 sg13g2_a21o_1 _1680_ (.A2(_0621_),
    .A1(_0334_),
    .B1(_0769_),
    .X(_0770_));
 sg13g2_o21ai_1 _1681_ (.B1(_0770_),
    .Y(_0771_),
    .A1(_0332_),
    .A2(_0620_));
 sg13g2_nor2_1 _1682_ (.A(_0307_),
    .B(_0610_),
    .Y(_0772_));
 sg13g2_nand2_1 _1683_ (.Y(_0773_),
    .A(net69),
    .B(_0573_));
 sg13g2_nor2b_1 _1684_ (.A(_0297_),
    .B_N(_0573_),
    .Y(_0774_));
 sg13g2_xnor2_1 _1685_ (.Y(_0775_),
    .A(_0685_),
    .B(_0774_));
 sg13g2_xnor2_1 _1686_ (.Y(_0776_),
    .A(_0668_),
    .B(_0775_));
 sg13g2_xnor2_1 _1687_ (.Y(_0777_),
    .A(_0773_),
    .B(_0776_));
 sg13g2_nor2_1 _1688_ (.A(_0246_),
    .B(_0567_),
    .Y(_0778_));
 sg13g2_nand2_2 _1689_ (.Y(_0779_),
    .A(net89),
    .B(net122));
 sg13g2_xor2_1 _1690_ (.B(_0779_),
    .A(_0672_),
    .X(_0780_));
 sg13g2_xnor2_1 _1691_ (.Y(_0781_),
    .A(_0778_),
    .B(_0780_));
 sg13g2_xnor2_1 _1692_ (.Y(_0782_),
    .A(_0777_),
    .B(_0781_));
 sg13g2_xnor2_1 _1693_ (.Y(_0783_),
    .A(_0772_),
    .B(_0782_));
 sg13g2_xnor2_1 _1694_ (.Y(_0784_),
    .A(_0771_),
    .B(_0783_));
 sg13g2_xnor2_1 _1695_ (.Y(_0785_),
    .A(_0768_),
    .B(_0784_));
 sg13g2_xor2_1 _1696_ (.B(_0785_),
    .A(_0766_),
    .X(_0786_));
 sg13g2_nor2_1 _1697_ (.A(_0418_),
    .B(_0539_),
    .Y(_0787_));
 sg13g2_nor2_1 _1698_ (.A(_0232_),
    .B(_0539_),
    .Y(_0788_));
 sg13g2_xor2_1 _1699_ (.B(_0750_),
    .A(_0742_),
    .X(_0789_));
 sg13g2_xor2_1 _1700_ (.B(_0418_),
    .A(_0231_),
    .X(_0790_));
 sg13g2_nor2_1 _1701_ (.A(_0524_),
    .B(_0790_),
    .Y(_0791_));
 sg13g2_nand3b_1 _1702_ (.B(\prd_i[2] ),
    .C(net89),
    .Y(_0792_),
    .A_N(\prd_i[5] ));
 sg13g2_o21ai_1 _1703_ (.B1(_0792_),
    .Y(_0793_),
    .A1(\prd_i[2] ),
    .A2(_0779_));
 sg13g2_mux2_1 _1704_ (.A0(_0746_),
    .A1(\prd_i[7] ),
    .S(_0793_),
    .X(_0794_));
 sg13g2_xnor2_1 _1705_ (.Y(_0795_),
    .A(_0791_),
    .B(_0794_));
 sg13g2_xnor2_1 _1706_ (.Y(_0796_),
    .A(_0789_),
    .B(_0795_));
 sg13g2_xnor2_1 _1707_ (.Y(_0797_),
    .A(_0777_),
    .B(_0796_));
 sg13g2_xnor2_1 _1708_ (.Y(_0798_),
    .A(_0788_),
    .B(_0797_));
 sg13g2_xnor2_1 _1709_ (.Y(_0799_),
    .A(_0787_),
    .B(_0798_));
 sg13g2_xnor2_1 _1710_ (.Y(_0800_),
    .A(_0739_),
    .B(_0799_));
 sg13g2_xnor2_1 _1711_ (.Y(_0801_),
    .A(_0760_),
    .B(_0768_));
 sg13g2_xnor2_1 _1712_ (.Y(_0802_),
    .A(_0800_),
    .B(_0801_));
 sg13g2_xnor2_1 _1713_ (.Y(_0803_),
    .A(_0786_),
    .B(_0802_));
 sg13g2_xnor2_1 _1714_ (.Y(_0804_),
    .A(_0758_),
    .B(_0803_));
 sg13g2_xor2_1 _1715_ (.B(_0730_),
    .A(_0654_),
    .X(_0805_));
 sg13g2_xnor2_1 _1716_ (.Y(_0806_),
    .A(_0804_),
    .B(_0805_));
 sg13g2_nand3_1 _1717_ (.B(net128),
    .C(_0694_),
    .A(net88),
    .Y(_0807_));
 sg13g2_and2_1 _1718_ (.A(_0092_),
    .B(_0807_),
    .X(_0808_));
 sg13g2_o21ai_1 _1719_ (.B1(_0808_),
    .Y(_0809_),
    .A1(_0208_),
    .A2(_0806_));
 sg13g2_nand2_1 _1720_ (.Y(_0810_),
    .A(_0153_),
    .B(_0198_));
 sg13g2_nand2_1 _1721_ (.Y(_0811_),
    .A(_0140_),
    .B(_0186_));
 sg13g2_xnor2_1 _1722_ (.Y(_0812_),
    .A(_0810_),
    .B(_0811_));
 sg13g2_xnor2_1 _1723_ (.Y(_0813_),
    .A(_0190_),
    .B(_0812_));
 sg13g2_xnor2_1 _1724_ (.Y(_0814_),
    .A(_0708_),
    .B(_0813_));
 sg13g2_nor2_1 _1725_ (.A(_0120_),
    .B(_0180_),
    .Y(_0815_));
 sg13g2_xnor2_1 _1726_ (.Y(_0816_),
    .A(_0193_),
    .B(_0815_));
 sg13g2_nand2_1 _1727_ (.Y(_0817_),
    .A(_0152_),
    .B(_0174_));
 sg13g2_xnor2_1 _1728_ (.Y(_0818_),
    .A(_0810_),
    .B(_0817_));
 sg13g2_xnor2_1 _1729_ (.Y(_0819_),
    .A(_0816_),
    .B(_0818_));
 sg13g2_xnor2_1 _1730_ (.Y(_0820_),
    .A(_0200_),
    .B(_0701_));
 sg13g2_xnor2_1 _1731_ (.Y(_0821_),
    .A(_0819_),
    .B(_0820_));
 sg13g2_xnor2_1 _1732_ (.Y(_0822_),
    .A(_0814_),
    .B(_0821_));
 sg13g2_o21ai_1 _1733_ (.B1(_0093_),
    .Y(_0823_),
    .A1(net78),
    .A2(_0822_));
 sg13g2_a22oi_1 _1734_ (.Y(_0824_),
    .B1(_0809_),
    .B2(_0823_),
    .A2(net79),
    .A1(net157));
 sg13g2_nor2_1 _1735_ (.A(_0066_),
    .B(_0824_),
    .Y(_0018_));
 sg13g2_nand2_1 _1736_ (.Y(_0825_),
    .A(net115),
    .B(net79));
 sg13g2_nand2_1 _1737_ (.Y(_0826_),
    .A(_0134_),
    .B(_0186_));
 sg13g2_xnor2_1 _1738_ (.Y(_0827_),
    .A(_0199_),
    .B(_0826_));
 sg13g2_xnor2_1 _1739_ (.Y(_0828_),
    .A(_0705_),
    .B(_0827_));
 sg13g2_xor2_1 _1740_ (.B(_0828_),
    .A(_0814_),
    .X(_0829_));
 sg13g2_xor2_1 _1741_ (.B(_0829_),
    .A(_0204_),
    .X(_0830_));
 sg13g2_o21ai_1 _1742_ (.B1(_0093_),
    .Y(_0831_),
    .A1(net78),
    .A2(_0830_));
 sg13g2_nor2_1 _1743_ (.A(_0265_),
    .B(_0555_),
    .Y(_0832_));
 sg13g2_xor2_1 _1744_ (.B(_0748_),
    .A(_0564_),
    .X(_0833_));
 sg13g2_xnor2_1 _1745_ (.Y(_0834_),
    .A(_0265_),
    .B(net67));
 sg13g2_nor2_1 _1746_ (.A(_0542_),
    .B(_0834_),
    .Y(_0835_));
 sg13g2_xnor2_1 _1747_ (.Y(_0836_),
    .A(_0833_),
    .B(_0835_));
 sg13g2_xnor2_1 _1748_ (.Y(_0837_),
    .A(_0580_),
    .B(_0836_));
 sg13g2_xnor2_1 _1749_ (.Y(_0838_),
    .A(_0721_),
    .B(_0837_));
 sg13g2_nor2_1 _1750_ (.A(net67),
    .B(_0555_),
    .Y(_0839_));
 sg13g2_xnor2_1 _1751_ (.Y(_0840_),
    .A(_0838_),
    .B(_0839_));
 sg13g2_xnor2_1 _1752_ (.Y(_0841_),
    .A(_0559_),
    .B(_0840_));
 sg13g2_xnor2_1 _1753_ (.Y(_0842_),
    .A(_0832_),
    .B(_0841_));
 sg13g2_xnor2_1 _1754_ (.Y(_0843_),
    .A(_0716_),
    .B(_0842_));
 sg13g2_xor2_1 _1755_ (.B(_0758_),
    .A(_0730_),
    .X(_0844_));
 sg13g2_xor2_1 _1756_ (.B(_0844_),
    .A(_0843_),
    .X(_0845_));
 sg13g2_xor2_1 _1757_ (.B(_0845_),
    .A(_0656_),
    .X(_0846_));
 sg13g2_nand3_1 _1758_ (.B(\prd_i[3] ),
    .C(_0694_),
    .A(net88),
    .Y(_0847_));
 sg13g2_o21ai_1 _1759_ (.B1(_0847_),
    .Y(_0848_),
    .A1(_0208_),
    .A2(_0846_));
 sg13g2_o21ai_1 _1760_ (.B1(_0831_),
    .Y(_0849_),
    .A1(_0093_),
    .A2(_0848_));
 sg13g2_a21oi_1 _1761_ (.A1(_0825_),
    .A2(_0849_),
    .Y(_0019_),
    .B1(_0066_));
 sg13g2_a22oi_1 _1762_ (.Y(_0850_),
    .B1(_0845_),
    .B2(_0207_),
    .A2(_0694_),
    .A1(_0583_));
 sg13g2_a22oi_1 _1763_ (.Y(_0851_),
    .B1(_0850_),
    .B2(_0092_),
    .A2(_0829_),
    .A1(_0091_));
 sg13g2_o21ai_1 _1764_ (.B1(net97),
    .Y(_0852_),
    .A1(net79),
    .A2(_0851_));
 sg13g2_a21oi_1 _1765_ (.A1(_0057_),
    .A2(net79),
    .Y(_0020_),
    .B1(_0852_));
 sg13g2_xor2_1 _1766_ (.B(_0786_),
    .A(_0654_),
    .X(_0853_));
 sg13g2_nor2b_1 _1767_ (.A(_0187_),
    .B_N(_0141_),
    .Y(_0854_));
 sg13g2_xnor2_1 _1768_ (.Y(_0855_),
    .A(_0182_),
    .B(_0854_));
 sg13g2_xnor2_1 _1769_ (.Y(_0856_),
    .A(_0816_),
    .B(_0855_));
 sg13g2_nor2b_1 _1770_ (.A(_0088_),
    .B_N(_0091_),
    .Y(_0857_));
 sg13g2_xnor2_1 _1771_ (.Y(_0858_),
    .A(_0820_),
    .B(_0856_));
 sg13g2_nor3_1 _1772_ (.A(_0078_),
    .B(net84),
    .C(_0779_),
    .Y(_0859_));
 sg13g2_a21oi_1 _1773_ (.A1(_0207_),
    .A2(_0853_),
    .Y(_0860_),
    .B1(_0859_));
 sg13g2_a22oi_1 _1774_ (.Y(_0861_),
    .B1(_0857_),
    .B2(_0858_),
    .A2(net78),
    .A1(net164));
 sg13g2_a21oi_1 _1775_ (.A1(_0860_),
    .A2(_0861_),
    .Y(_0021_),
    .B1(_0066_));
 sg13g2_xor2_1 _1776_ (.B(_0843_),
    .A(_0758_),
    .X(_0862_));
 sg13g2_nor3_1 _1777_ (.A(_0078_),
    .B(net84),
    .C(_0585_),
    .Y(_0863_));
 sg13g2_a21oi_1 _1778_ (.A1(_0207_),
    .A2(_0862_),
    .Y(_0864_),
    .B1(_0863_));
 sg13g2_nand2_1 _1779_ (.Y(_0865_),
    .A(_0092_),
    .B(_0864_));
 sg13g2_xnor2_1 _1780_ (.Y(_0866_),
    .A(_0813_),
    .B(_0828_));
 sg13g2_o21ai_1 _1781_ (.B1(_0093_),
    .Y(_0867_),
    .A1(net78),
    .A2(_0866_));
 sg13g2_a22oi_1 _1782_ (.Y(_0868_),
    .B1(_0865_),
    .B2(_0867_),
    .A2(net78),
    .A1(net151));
 sg13g2_nor2_1 _1783_ (.A(_0066_),
    .B(net152),
    .Y(_0022_));
 sg13g2_nand3_1 _1784_ (.B(net136),
    .C(_0694_),
    .A(net88),
    .Y(_0869_));
 sg13g2_and2_1 _1785_ (.A(_0092_),
    .B(_0869_),
    .X(_0870_));
 sg13g2_o21ai_1 _1786_ (.B1(_0870_),
    .Y(_0871_),
    .A1(_0208_),
    .A2(_0844_));
 sg13g2_a21o_1 _1787_ (.A2(_0814_),
    .A1(_0089_),
    .B1(_0092_),
    .X(_0872_));
 sg13g2_a22oi_1 _1788_ (.Y(_0873_),
    .B1(_0871_),
    .B2(_0872_),
    .A2(net78),
    .A1(net142));
 sg13g2_nor2_1 _1789_ (.A(_0066_),
    .B(_0873_),
    .Y(_0023_));
 sg13g2_nand3_1 _1790_ (.B(net9),
    .C(net97),
    .A(net10),
    .Y(_0874_));
 sg13g2_nor3_2 _1791_ (.A(net11),
    .B(net12),
    .C(_0874_),
    .Y(_0875_));
 sg13g2_nor2_1 _1792_ (.A(net149),
    .B(net77),
    .Y(_0876_));
 sg13g2_a21oi_1 _1793_ (.A1(_0065_),
    .A2(net77),
    .Y(_0024_),
    .B1(_0876_));
 sg13g2_nor2_1 _1794_ (.A(net124),
    .B(net77),
    .Y(_0877_));
 sg13g2_a21oi_1 _1795_ (.A1(_0064_),
    .A2(net77),
    .Y(_0025_),
    .B1(_0877_));
 sg13g2_nor2_1 _1796_ (.A(net114),
    .B(net76),
    .Y(_0878_));
 sg13g2_a21oi_1 _1797_ (.A1(_0063_),
    .A2(net76),
    .Y(_0026_),
    .B1(_0878_));
 sg13g2_nor2_1 _1798_ (.A(net118),
    .B(net76),
    .Y(_0879_));
 sg13g2_a21oi_1 _1799_ (.A1(_0062_),
    .A2(net76),
    .Y(_0027_),
    .B1(_0879_));
 sg13g2_nor2_1 _1800_ (.A(net123),
    .B(net77),
    .Y(_0880_));
 sg13g2_a21oi_1 _1801_ (.A1(_0061_),
    .A2(net77),
    .Y(_0028_),
    .B1(_0880_));
 sg13g2_nor2_1 _1802_ (.A(net117),
    .B(_0875_),
    .Y(_0881_));
 sg13g2_a21oi_1 _1803_ (.A1(_0060_),
    .A2(net77),
    .Y(_0029_),
    .B1(_0881_));
 sg13g2_nor2_1 _1804_ (.A(net125),
    .B(net76),
    .Y(_0882_));
 sg13g2_a21oi_1 _1805_ (.A1(_0059_),
    .A2(net76),
    .Y(_0030_),
    .B1(_0882_));
 sg13g2_nor2_1 _1806_ (.A(net129),
    .B(net76),
    .Y(_0883_));
 sg13g2_a21oi_1 _1807_ (.A1(_0058_),
    .A2(net76),
    .Y(_0031_),
    .B1(_0883_));
 sg13g2_nand3b_1 _1808_ (.B(net97),
    .C(net11),
    .Y(_0884_),
    .A_N(net12));
 sg13g2_nor2_2 _1809_ (.A(_0078_),
    .B(_0884_),
    .Y(_0885_));
 sg13g2_nor2_1 _1810_ (.A(net148),
    .B(_0885_),
    .Y(_0886_));
 sg13g2_a21oi_1 _1811_ (.A1(_0065_),
    .A2(_0885_),
    .Y(_0032_),
    .B1(_0886_));
 sg13g2_nor2_1 _1812_ (.A(net133),
    .B(_0885_),
    .Y(_0887_));
 sg13g2_a21oi_1 _1813_ (.A1(_0064_),
    .A2(_0885_),
    .Y(_0033_),
    .B1(_0887_));
 sg13g2_nor2_1 _1814_ (.A(_0068_),
    .B(_0884_),
    .Y(_0888_));
 sg13g2_nor2_1 _1815_ (.A(net134),
    .B(net73),
    .Y(_0889_));
 sg13g2_a21oi_1 _1816_ (.A1(_0065_),
    .A2(net73),
    .Y(_0034_),
    .B1(_0889_));
 sg13g2_nor2_1 _1817_ (.A(net121),
    .B(net73),
    .Y(_0890_));
 sg13g2_a21oi_1 _1818_ (.A1(_0064_),
    .A2(net73),
    .Y(_0035_),
    .B1(_0890_));
 sg13g2_nor2_1 _1819_ (.A(net140),
    .B(net74),
    .Y(_0891_));
 sg13g2_a21oi_1 _1820_ (.A1(_0063_),
    .A2(net73),
    .Y(_0036_),
    .B1(_0891_));
 sg13g2_nor2_1 _1821_ (.A(net139),
    .B(net74),
    .Y(_0892_));
 sg13g2_a21oi_1 _1822_ (.A1(_0062_),
    .A2(net73),
    .Y(_0037_),
    .B1(_0892_));
 sg13g2_nor2_1 _1823_ (.A(net159),
    .B(net73),
    .Y(_0893_));
 sg13g2_a21oi_1 _1824_ (.A1(_0061_),
    .A2(net73),
    .Y(_0038_),
    .B1(_0893_));
 sg13g2_nor2_1 _1825_ (.A(net130),
    .B(net74),
    .Y(_0894_));
 sg13g2_a21oi_1 _1826_ (.A1(_0060_),
    .A2(net74),
    .Y(_0039_),
    .B1(_0894_));
 sg13g2_nor2_1 _1827_ (.A(net132),
    .B(net75),
    .Y(_0895_));
 sg13g2_a21oi_1 _1828_ (.A1(_0059_),
    .A2(net75),
    .Y(_0040_),
    .B1(_0895_));
 sg13g2_nor2_1 _1829_ (.A(net135),
    .B(net75),
    .Y(_0896_));
 sg13g2_a21oi_1 _1830_ (.A1(_0058_),
    .A2(net75),
    .Y(_0041_),
    .B1(_0896_));
 sg13g2_nor3_2 _1831_ (.A(net10),
    .B(net9),
    .C(_0884_),
    .Y(_0897_));
 sg13g2_nor2_1 _1832_ (.A(net119),
    .B(net71),
    .Y(_0898_));
 sg13g2_a21oi_1 _1833_ (.A1(_0065_),
    .A2(net71),
    .Y(_0042_),
    .B1(_0898_));
 sg13g2_nor2_1 _1834_ (.A(net120),
    .B(net71),
    .Y(_0050_));
 sg13g2_a21oi_1 _1835_ (.A1(_0064_),
    .A2(net71),
    .Y(_0043_),
    .B1(_0050_));
 sg13g2_nor2_1 _1836_ (.A(net128),
    .B(net72),
    .Y(_0051_));
 sg13g2_a21oi_1 _1837_ (.A1(_0063_),
    .A2(net72),
    .Y(_0044_),
    .B1(_0051_));
 sg13g2_nor2_1 _1838_ (.A(net127),
    .B(net72),
    .Y(_0052_));
 sg13g2_a21oi_1 _1839_ (.A1(_0062_),
    .A2(net72),
    .Y(_0045_),
    .B1(_0052_));
 sg13g2_nor2_1 _1840_ (.A(net131),
    .B(net72),
    .Y(_0053_));
 sg13g2_a21oi_1 _1841_ (.A1(_0061_),
    .A2(net72),
    .Y(_0046_),
    .B1(_0053_));
 sg13g2_nor2_1 _1842_ (.A(net122),
    .B(net72),
    .Y(_0054_));
 sg13g2_a21oi_1 _1843_ (.A1(_0060_),
    .A2(net72),
    .Y(_0047_),
    .B1(_0054_));
 sg13g2_nor2_1 _1844_ (.A(net126),
    .B(net71),
    .Y(_0055_));
 sg13g2_a21oi_1 _1845_ (.A1(_0059_),
    .A2(net71),
    .Y(_0048_),
    .B1(_0055_));
 sg13g2_nor2_1 _1846_ (.A(net136),
    .B(net71),
    .Y(_0056_));
 sg13g2_a21oi_1 _1847_ (.A1(_0058_),
    .A2(net71),
    .Y(_0049_),
    .B1(_0056_));
 sg13g2_dfrbpq_1 _1848_ (.RESET_B(net53),
    .D(_0000_),
    .Q(\data_i[0] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_2 _1849_ (.RESET_B(net48),
    .D(_0001_),
    .Q(\data_i[1] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_2 _1850_ (.RESET_B(net46),
    .D(_0002_),
    .Q(\data_i[2] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_1 _1851_ (.RESET_B(net44),
    .D(_0003_),
    .Q(\data_i[3] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _1852_ (.RESET_B(net42),
    .D(_0004_),
    .Q(\data_i[4] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_1 _1853_ (.RESET_B(net40),
    .D(_0005_),
    .Q(\data_i[5] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _1854_ (.RESET_B(net38),
    .D(_0006_),
    .Q(\data_i[6] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_1 _1855_ (.RESET_B(net36),
    .D(_0007_),
    .Q(\data_i[7] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_1 _1856_ (.RESET_B(net34),
    .D(_0008_),
    .Q(\key[0] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_2 _1857_ (.RESET_B(net32),
    .D(_0009_),
    .Q(\key[1] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_2 _1858_ (.RESET_B(net30),
    .D(_0010_),
    .Q(\key[2] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_1 _1859_ (.RESET_B(net111),
    .D(_0011_),
    .Q(\key[3] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _1860_ (.RESET_B(net109),
    .D(_0012_),
    .Q(\key[4] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _1861_ (.RESET_B(net107),
    .D(_0013_),
    .Q(\key[5] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_1 _1862_ (.RESET_B(net105),
    .D(_0014_),
    .Q(\key[6] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _1863_ (.RESET_B(net103),
    .D(_0015_),
    .Q(\key[7] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_2 _1864_ (.RESET_B(net101),
    .D(_0016_),
    .Q(uo_out[0]),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _1865_ (.RESET_B(net99),
    .D(_0017_),
    .Q(uo_out[1]),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _1866_ (.RESET_B(net64),
    .D(_0018_),
    .Q(uo_out[2]),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _1867_ (.RESET_B(net62),
    .D(net116),
    .Q(uo_out[3]),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _1868_ (.RESET_B(net60),
    .D(_0020_),
    .Q(uo_out[4]),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_2 _1869_ (.RESET_B(net58),
    .D(_0021_),
    .Q(uo_out[5]),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _1870_ (.RESET_B(net56),
    .D(_0022_),
    .Q(uo_out[6]),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _1871_ (.RESET_B(net54),
    .D(_0023_),
    .Q(uo_out[7]),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _1872_ (.RESET_B(net52),
    .D(_0024_),
    .Q(\mask_i[0] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _1873_ (.RESET_B(net51),
    .D(_0025_),
    .Q(\mask_i[1] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_1 _1874_ (.RESET_B(net50),
    .D(_0026_),
    .Q(\mask_i[2] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _1875_ (.RESET_B(net49),
    .D(_0027_),
    .Q(\mask_i[3] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _1876_ (.RESET_B(net47),
    .D(_0028_),
    .Q(\mask_i[4] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_1 _1877_ (.RESET_B(net45),
    .D(_0029_),
    .Q(\mask_i[5] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _1878_ (.RESET_B(net43),
    .D(_0030_),
    .Q(\mask_i[6] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_2 _1879_ (.RESET_B(net41),
    .D(_0031_),
    .Q(\mask_i[7] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _1880_ (.RESET_B(net39),
    .D(_0032_),
    .Q(\prd_i[16] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _1881_ (.RESET_B(net37),
    .D(_0033_),
    .Q(\prd_i[17] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_2 _1882_ (.RESET_B(net35),
    .D(_0034_),
    .Q(\prd_i[8] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _1883_ (.RESET_B(net33),
    .D(_0035_),
    .Q(\prd_i[9] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_2 _1884_ (.RESET_B(net31),
    .D(_0036_),
    .Q(\prd_i[10] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_2 _1885_ (.RESET_B(net112),
    .D(_0037_),
    .Q(\prd_i[11] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_2 _1886_ (.RESET_B(net110),
    .D(_0038_),
    .Q(\prd_i[12] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_2 _1887_ (.RESET_B(net108),
    .D(_0039_),
    .Q(\prd_i[13] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_2 _1888_ (.RESET_B(net106),
    .D(_0040_),
    .Q(\prd_i[14] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _1889_ (.RESET_B(net104),
    .D(_0041_),
    .Q(\prd_i[15] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _1890_ (.RESET_B(net102),
    .D(_0042_),
    .Q(\prd_i[0] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _1891_ (.RESET_B(net100),
    .D(_0043_),
    .Q(\prd_i[1] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _1892_ (.RESET_B(net98),
    .D(_0044_),
    .Q(\prd_i[2] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_2 _1893_ (.RESET_B(net63),
    .D(_0045_),
    .Q(\prd_i[3] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_2 _1894_ (.RESET_B(net61),
    .D(_0046_),
    .Q(\prd_i[4] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_2 _1895_ (.RESET_B(net59),
    .D(_0047_),
    .Q(\prd_i[5] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _1896_ (.RESET_B(net57),
    .D(_0048_),
    .Q(\prd_i[6] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _1897_ (.RESET_B(net55),
    .D(_0049_),
    .Q(\prd_i[7] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_tiehi _1884__31 (.L_HI(net31));
 sg13g2_tiehi _1857__32 (.L_HI(net32));
 sg13g2_tiehi _1883__33 (.L_HI(net33));
 sg13g2_tiehi _1856__34 (.L_HI(net34));
 sg13g2_tiehi _1882__35 (.L_HI(net35));
 sg13g2_tiehi _1855__36 (.L_HI(net36));
 sg13g2_tiehi _1881__37 (.L_HI(net37));
 sg13g2_tiehi _1854__38 (.L_HI(net38));
 sg13g2_tiehi _1880__39 (.L_HI(net39));
 sg13g2_tiehi _1853__40 (.L_HI(net40));
 sg13g2_tiehi _1879__41 (.L_HI(net41));
 sg13g2_tiehi _1852__42 (.L_HI(net42));
 sg13g2_tiehi _1878__43 (.L_HI(net43));
 sg13g2_tiehi _1851__44 (.L_HI(net44));
 sg13g2_tiehi _1877__45 (.L_HI(net45));
 sg13g2_tiehi _1850__46 (.L_HI(net46));
 sg13g2_tiehi _1876__47 (.L_HI(net47));
 sg13g2_tiehi _1849__48 (.L_HI(net48));
 sg13g2_tiehi _1875__49 (.L_HI(net49));
 sg13g2_tiehi _1874__50 (.L_HI(net50));
 sg13g2_tiehi _1873__51 (.L_HI(net51));
 sg13g2_tiehi _1872__52 (.L_HI(net52));
 sg13g2_tiehi _1848__53 (.L_HI(net53));
 sg13g2_tiehi _1871__54 (.L_HI(net54));
 sg13g2_tiehi _1897__55 (.L_HI(net55));
 sg13g2_tiehi _1870__56 (.L_HI(net56));
 sg13g2_tiehi _1896__57 (.L_HI(net57));
 sg13g2_tiehi _1869__58 (.L_HI(net58));
 sg13g2_tiehi _1895__59 (.L_HI(net59));
 sg13g2_tiehi _1868__60 (.L_HI(net60));
 sg13g2_tiehi _1894__61 (.L_HI(net61));
 sg13g2_tiehi _1867__62 (.L_HI(net62));
 sg13g2_tiehi _1893__63 (.L_HI(net63));
 sg13g2_tiehi _1866__64 (.L_HI(net64));
 sg13g2_tiehi _1892__65 (.L_HI(net98));
 sg13g2_tiehi _1865__66 (.L_HI(net99));
 sg13g2_tiehi _1891__67 (.L_HI(net100));
 sg13g2_tiehi _1864__68 (.L_HI(net101));
 sg13g2_tiehi _1890__69 (.L_HI(net102));
 sg13g2_tiehi _1863__70 (.L_HI(net103));
 sg13g2_tiehi _1889__71 (.L_HI(net104));
 sg13g2_tiehi _1862__72 (.L_HI(net105));
 sg13g2_tiehi _1888__73 (.L_HI(net106));
 sg13g2_tiehi _1861__74 (.L_HI(net107));
 sg13g2_tiehi _1887__75 (.L_HI(net108));
 sg13g2_tiehi _1860__76 (.L_HI(net109));
 sg13g2_tiehi _1886__77 (.L_HI(net110));
 sg13g2_tiehi _1859__78 (.L_HI(net111));
 sg13g2_tiehi _1885__79 (.L_HI(net112));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_coastalwhite_canright_sbox_15 (.L_LO(net15));
 sg13g2_tielo tt_um_coastalwhite_canright_sbox_16 (.L_LO(net16));
 sg13g2_tielo tt_um_coastalwhite_canright_sbox_17 (.L_LO(net17));
 sg13g2_tielo tt_um_coastalwhite_canright_sbox_18 (.L_LO(net18));
 sg13g2_tielo tt_um_coastalwhite_canright_sbox_19 (.L_LO(net19));
 sg13g2_tielo tt_um_coastalwhite_canright_sbox_20 (.L_LO(net20));
 sg13g2_tielo tt_um_coastalwhite_canright_sbox_21 (.L_LO(net21));
 sg13g2_tielo tt_um_coastalwhite_canright_sbox_22 (.L_LO(net22));
 sg13g2_tielo tt_um_coastalwhite_canright_sbox_23 (.L_LO(net23));
 sg13g2_tielo tt_um_coastalwhite_canright_sbox_24 (.L_LO(net24));
 sg13g2_tielo tt_um_coastalwhite_canright_sbox_25 (.L_LO(net25));
 sg13g2_tielo tt_um_coastalwhite_canright_sbox_26 (.L_LO(net26));
 sg13g2_tielo tt_um_coastalwhite_canright_sbox_27 (.L_LO(net27));
 sg13g2_tielo tt_um_coastalwhite_canright_sbox_28 (.L_LO(net28));
 sg13g2_tielo tt_um_coastalwhite_canright_sbox_29 (.L_LO(net29));
 sg13g2_tiehi _1858__30 (.L_HI(net30));
 sg13g2_buf_8 fanout65 (.A(_0610_),
    .X(net65));
 sg13g2_buf_8 fanout66 (.A(_0341_),
    .X(net66));
 sg13g2_buf_8 fanout67 (.A(_0345_),
    .X(net67));
 sg13g2_buf_8 fanout68 (.A(_0296_),
    .X(net68));
 sg13g2_buf_8 fanout69 (.A(_0254_),
    .X(net69));
 sg13g2_buf_8 fanout70 (.A(_0209_),
    .X(net70));
 sg13g2_buf_8 fanout71 (.A(_0897_),
    .X(net71));
 sg13g2_buf_8 fanout72 (.A(_0897_),
    .X(net72));
 sg13g2_buf_8 fanout73 (.A(net75),
    .X(net73));
 sg13g2_buf_1 fanout74 (.A(net75),
    .X(net74));
 sg13g2_buf_8 fanout75 (.A(_0888_),
    .X(net75));
 sg13g2_buf_8 fanout76 (.A(net77),
    .X(net76));
 sg13g2_buf_8 fanout77 (.A(_0875_),
    .X(net77));
 sg13g2_buf_8 fanout78 (.A(_0090_),
    .X(net78));
 sg13g2_buf_8 fanout79 (.A(_0090_),
    .X(net79));
 sg13g2_buf_8 fanout80 (.A(net81),
    .X(net80));
 sg13g2_buf_8 fanout81 (.A(_0079_),
    .X(net81));
 sg13g2_buf_8 fanout82 (.A(net83),
    .X(net82));
 sg13g2_buf_8 fanout83 (.A(_0069_),
    .X(net83));
 sg13g2_buf_8 fanout84 (.A(_0088_),
    .X(net84));
 sg13g2_buf_8 fanout85 (.A(net13),
    .X(net85));
 sg13g2_buf_8 fanout86 (.A(net94),
    .X(net86));
 sg13g2_buf_8 fanout87 (.A(net94),
    .X(net87));
 sg13g2_buf_8 fanout88 (.A(net89),
    .X(net88));
 sg13g2_buf_1 fanout89 (.A(net90),
    .X(net89));
 sg13g2_buf_1 fanout90 (.A(net94),
    .X(net90));
 sg13g2_buf_8 fanout91 (.A(net93),
    .X(net91));
 sg13g2_buf_8 fanout92 (.A(net93),
    .X(net92));
 sg13g2_buf_8 fanout93 (.A(net94),
    .X(net93));
 sg13g2_buf_8 fanout94 (.A(uio_in[6]),
    .X(net94));
 sg13g2_buf_8 fanout95 (.A(net96),
    .X(net95));
 sg13g2_buf_8 fanout96 (.A(net97),
    .X(net96));
 sg13g2_buf_8 fanout97 (.A(rst_n),
    .X(net97));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_2 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[7]),
    .X(net13));
 sg13g2_tielo tt_um_coastalwhite_canright_sbox_14 (.L_LO(net14));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_2__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_3_4__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_3_5__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_3_6__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(uo_out[4]),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold2 (.A(\mask_i[2] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold3 (.A(uo_out[3]),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0019_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold5 (.A(\mask_i[5] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold6 (.A(\mask_i[3] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold7 (.A(\prd_i[0] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold8 (.A(\prd_i[1] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold9 (.A(\prd_i[9] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold10 (.A(\prd_i[5] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold11 (.A(\mask_i[4] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold12 (.A(\mask_i[1] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold13 (.A(\mask_i[6] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold14 (.A(\prd_i[6] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold15 (.A(\prd_i[3] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold16 (.A(\prd_i[2] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold17 (.A(\mask_i[7] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold18 (.A(\prd_i[13] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold19 (.A(\prd_i[4] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold20 (.A(\prd_i[14] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold21 (.A(\prd_i[17] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold22 (.A(\prd_i[8] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold23 (.A(\prd_i[15] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold24 (.A(\prd_i[7] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold25 (.A(uo_out[1]),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold26 (.A(uo_out[0]),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold27 (.A(\prd_i[11] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold28 (.A(\prd_i[10] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold29 (.A(\data_i[5] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold30 (.A(uo_out[7]),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold31 (.A(\key[3] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold32 (.A(\data_i[4] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold33 (.A(\data_i[0] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold34 (.A(\data_i[3] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold35 (.A(\key[0] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold36 (.A(\prd_i[16] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold37 (.A(\mask_i[0] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold38 (.A(\key[5] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold39 (.A(uo_out[6]),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0868_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold41 (.A(\key[6] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold42 (.A(\data_i[7] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold43 (.A(\key[7] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold44 (.A(\key[4] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold45 (.A(uo_out[2]),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold46 (.A(\data_i[6] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold47 (.A(\prd_i[12] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold48 (.A(\data_i[1] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold49 (.A(\key[1] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold50 (.A(\key[2] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold51 (.A(\data_i[2] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold52 (.A(uo_out[5]),
    .X(net164));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_fill_2 FILLER_7_98 ();
 sg13g2_fill_1 FILLER_7_100 ();
 sg13g2_decap_8 FILLER_7_106 ();
 sg13g2_decap_8 FILLER_7_113 ();
 sg13g2_fill_2 FILLER_7_120 ();
 sg13g2_fill_1 FILLER_7_122 ();
 sg13g2_decap_8 FILLER_7_128 ();
 sg13g2_decap_8 FILLER_7_135 ();
 sg13g2_decap_8 FILLER_7_142 ();
 sg13g2_fill_1 FILLER_7_149 ();
 sg13g2_fill_1 FILLER_7_159 ();
 sg13g2_decap_4 FILLER_7_168 ();
 sg13g2_fill_1 FILLER_7_172 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_4 FILLER_7_224 ();
 sg13g2_fill_2 FILLER_7_228 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_4 FILLER_7_252 ();
 sg13g2_fill_1 FILLER_7_256 ();
 sg13g2_decap_8 FILLER_7_269 ();
 sg13g2_fill_1 FILLER_7_276 ();
 sg13g2_fill_2 FILLER_7_285 ();
 sg13g2_fill_1 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_293 ();
 sg13g2_decap_8 FILLER_7_300 ();
 sg13g2_decap_8 FILLER_7_307 ();
 sg13g2_decap_8 FILLER_7_318 ();
 sg13g2_decap_8 FILLER_7_325 ();
 sg13g2_decap_4 FILLER_7_332 ();
 sg13g2_fill_2 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_347 ();
 sg13g2_decap_8 FILLER_7_354 ();
 sg13g2_decap_8 FILLER_7_361 ();
 sg13g2_decap_8 FILLER_7_368 ();
 sg13g2_decap_8 FILLER_7_375 ();
 sg13g2_decap_8 FILLER_7_382 ();
 sg13g2_decap_8 FILLER_7_389 ();
 sg13g2_decap_8 FILLER_7_396 ();
 sg13g2_decap_4 FILLER_7_403 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_4 FILLER_8_63 ();
 sg13g2_fill_2 FILLER_8_67 ();
 sg13g2_fill_1 FILLER_8_77 ();
 sg13g2_decap_4 FILLER_8_84 ();
 sg13g2_fill_2 FILLER_8_88 ();
 sg13g2_fill_1 FILLER_8_103 ();
 sg13g2_decap_8 FILLER_8_113 ();
 sg13g2_decap_8 FILLER_8_136 ();
 sg13g2_fill_2 FILLER_8_143 ();
 sg13g2_decap_4 FILLER_8_168 ();
 sg13g2_fill_2 FILLER_8_188 ();
 sg13g2_fill_1 FILLER_8_190 ();
 sg13g2_decap_8 FILLER_8_215 ();
 sg13g2_fill_1 FILLER_8_222 ();
 sg13g2_decap_8 FILLER_8_239 ();
 sg13g2_decap_4 FILLER_8_246 ();
 sg13g2_decap_4 FILLER_8_272 ();
 sg13g2_fill_1 FILLER_8_276 ();
 sg13g2_decap_4 FILLER_8_305 ();
 sg13g2_decap_8 FILLER_8_324 ();
 sg13g2_fill_2 FILLER_8_331 ();
 sg13g2_fill_1 FILLER_8_333 ();
 sg13g2_decap_8 FILLER_8_353 ();
 sg13g2_decap_8 FILLER_8_360 ();
 sg13g2_decap_4 FILLER_8_367 ();
 sg13g2_fill_1 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_380 ();
 sg13g2_decap_4 FILLER_8_387 ();
 sg13g2_fill_2 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_401 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_4 FILLER_9_49 ();
 sg13g2_fill_1 FILLER_9_53 ();
 sg13g2_decap_8 FILLER_9_61 ();
 sg13g2_fill_2 FILLER_9_68 ();
 sg13g2_fill_1 FILLER_9_70 ();
 sg13g2_fill_2 FILLER_9_76 ();
 sg13g2_decap_8 FILLER_9_90 ();
 sg13g2_fill_1 FILLER_9_97 ();
 sg13g2_decap_4 FILLER_9_103 ();
 sg13g2_fill_2 FILLER_9_107 ();
 sg13g2_decap_4 FILLER_9_113 ();
 sg13g2_fill_1 FILLER_9_117 ();
 sg13g2_decap_4 FILLER_9_123 ();
 sg13g2_fill_2 FILLER_9_127 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_4 FILLER_9_140 ();
 sg13g2_fill_2 FILLER_9_149 ();
 sg13g2_fill_1 FILLER_9_151 ();
 sg13g2_decap_4 FILLER_9_156 ();
 sg13g2_decap_8 FILLER_9_164 ();
 sg13g2_decap_8 FILLER_9_171 ();
 sg13g2_decap_8 FILLER_9_178 ();
 sg13g2_decap_8 FILLER_9_185 ();
 sg13g2_fill_1 FILLER_9_192 ();
 sg13g2_fill_1 FILLER_9_209 ();
 sg13g2_decap_4 FILLER_9_218 ();
 sg13g2_fill_2 FILLER_9_222 ();
 sg13g2_decap_4 FILLER_9_245 ();
 sg13g2_fill_2 FILLER_9_249 ();
 sg13g2_decap_8 FILLER_9_264 ();
 sg13g2_fill_2 FILLER_9_271 ();
 sg13g2_fill_1 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_282 ();
 sg13g2_decap_8 FILLER_9_289 ();
 sg13g2_fill_2 FILLER_9_296 ();
 sg13g2_decap_8 FILLER_9_306 ();
 sg13g2_fill_2 FILLER_9_313 ();
 sg13g2_fill_1 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_331 ();
 sg13g2_fill_1 FILLER_9_338 ();
 sg13g2_fill_2 FILLER_9_353 ();
 sg13g2_decap_4 FILLER_9_403 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_fill_2 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_61 ();
 sg13g2_decap_4 FILLER_10_68 ();
 sg13g2_fill_1 FILLER_10_79 ();
 sg13g2_fill_1 FILLER_10_109 ();
 sg13g2_fill_1 FILLER_10_123 ();
 sg13g2_fill_2 FILLER_10_143 ();
 sg13g2_fill_1 FILLER_10_145 ();
 sg13g2_decap_4 FILLER_10_165 ();
 sg13g2_fill_2 FILLER_10_169 ();
 sg13g2_fill_1 FILLER_10_186 ();
 sg13g2_decap_4 FILLER_10_196 ();
 sg13g2_fill_1 FILLER_10_200 ();
 sg13g2_fill_1 FILLER_10_209 ();
 sg13g2_fill_1 FILLER_10_229 ();
 sg13g2_decap_8 FILLER_10_240 ();
 sg13g2_fill_2 FILLER_10_247 ();
 sg13g2_fill_1 FILLER_10_249 ();
 sg13g2_fill_1 FILLER_10_258 ();
 sg13g2_decap_8 FILLER_10_267 ();
 sg13g2_fill_2 FILLER_10_298 ();
 sg13g2_fill_2 FILLER_10_312 ();
 sg13g2_fill_1 FILLER_10_314 ();
 sg13g2_fill_2 FILLER_10_332 ();
 sg13g2_decap_8 FILLER_10_342 ();
 sg13g2_decap_8 FILLER_10_349 ();
 sg13g2_fill_1 FILLER_10_356 ();
 sg13g2_decap_8 FILLER_10_365 ();
 sg13g2_decap_8 FILLER_10_380 ();
 sg13g2_decap_4 FILLER_10_387 ();
 sg13g2_fill_2 FILLER_10_391 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_fill_2 FILLER_11_49 ();
 sg13g2_fill_1 FILLER_11_51 ();
 sg13g2_decap_4 FILLER_11_70 ();
 sg13g2_fill_1 FILLER_11_84 ();
 sg13g2_fill_1 FILLER_11_89 ();
 sg13g2_decap_8 FILLER_11_102 ();
 sg13g2_decap_8 FILLER_11_109 ();
 sg13g2_decap_8 FILLER_11_116 ();
 sg13g2_fill_2 FILLER_11_128 ();
 sg13g2_fill_1 FILLER_11_130 ();
 sg13g2_decap_8 FILLER_11_136 ();
 sg13g2_decap_4 FILLER_11_143 ();
 sg13g2_fill_1 FILLER_11_147 ();
 sg13g2_fill_2 FILLER_11_153 ();
 sg13g2_fill_1 FILLER_11_155 ();
 sg13g2_decap_4 FILLER_11_164 ();
 sg13g2_fill_2 FILLER_11_168 ();
 sg13g2_fill_1 FILLER_11_182 ();
 sg13g2_decap_4 FILLER_11_188 ();
 sg13g2_fill_2 FILLER_11_192 ();
 sg13g2_fill_2 FILLER_11_202 ();
 sg13g2_fill_1 FILLER_11_204 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_4 FILLER_11_217 ();
 sg13g2_fill_2 FILLER_11_221 ();
 sg13g2_fill_2 FILLER_11_243 ();
 sg13g2_fill_1 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_262 ();
 sg13g2_fill_2 FILLER_11_269 ();
 sg13g2_fill_1 FILLER_11_271 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_4 FILLER_11_308 ();
 sg13g2_fill_1 FILLER_11_328 ();
 sg13g2_fill_2 FILLER_11_333 ();
 sg13g2_fill_1 FILLER_11_335 ();
 sg13g2_fill_2 FILLER_11_364 ();
 sg13g2_fill_1 FILLER_11_366 ();
 sg13g2_decap_8 FILLER_11_379 ();
 sg13g2_fill_2 FILLER_11_386 ();
 sg13g2_fill_1 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_4 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_66 ();
 sg13g2_decap_8 FILLER_12_73 ();
 sg13g2_fill_2 FILLER_12_80 ();
 sg13g2_fill_2 FILLER_12_88 ();
 sg13g2_fill_1 FILLER_12_90 ();
 sg13g2_decap_8 FILLER_12_102 ();
 sg13g2_decap_8 FILLER_12_109 ();
 sg13g2_fill_1 FILLER_12_125 ();
 sg13g2_decap_4 FILLER_12_131 ();
 sg13g2_decap_8 FILLER_12_148 ();
 sg13g2_fill_2 FILLER_12_155 ();
 sg13g2_fill_1 FILLER_12_157 ();
 sg13g2_decap_8 FILLER_12_164 ();
 sg13g2_fill_2 FILLER_12_179 ();
 sg13g2_decap_8 FILLER_12_184 ();
 sg13g2_fill_2 FILLER_12_191 ();
 sg13g2_decap_8 FILLER_12_214 ();
 sg13g2_decap_4 FILLER_12_221 ();
 sg13g2_decap_8 FILLER_12_237 ();
 sg13g2_decap_4 FILLER_12_244 ();
 sg13g2_decap_8 FILLER_12_260 ();
 sg13g2_decap_4 FILLER_12_267 ();
 sg13g2_fill_1 FILLER_12_271 ();
 sg13g2_decap_8 FILLER_12_312 ();
 sg13g2_decap_8 FILLER_12_319 ();
 sg13g2_decap_8 FILLER_12_326 ();
 sg13g2_decap_4 FILLER_12_333 ();
 sg13g2_decap_8 FILLER_12_341 ();
 sg13g2_fill_1 FILLER_12_348 ();
 sg13g2_decap_8 FILLER_12_353 ();
 sg13g2_decap_8 FILLER_12_360 ();
 sg13g2_fill_1 FILLER_12_367 ();
 sg13g2_fill_2 FILLER_12_389 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_fill_2 FILLER_13_65 ();
 sg13g2_fill_1 FILLER_13_97 ();
 sg13g2_decap_8 FILLER_13_110 ();
 sg13g2_fill_2 FILLER_13_117 ();
 sg13g2_decap_8 FILLER_13_124 ();
 sg13g2_decap_8 FILLER_13_131 ();
 sg13g2_fill_2 FILLER_13_138 ();
 sg13g2_fill_1 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_171 ();
 sg13g2_decap_8 FILLER_13_178 ();
 sg13g2_fill_2 FILLER_13_185 ();
 sg13g2_fill_2 FILLER_13_195 ();
 sg13g2_fill_2 FILLER_13_202 ();
 sg13g2_decap_8 FILLER_13_212 ();
 sg13g2_decap_8 FILLER_13_219 ();
 sg13g2_fill_1 FILLER_13_226 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_fill_2 FILLER_13_245 ();
 sg13g2_fill_1 FILLER_13_269 ();
 sg13g2_decap_8 FILLER_13_286 ();
 sg13g2_decap_8 FILLER_13_293 ();
 sg13g2_fill_1 FILLER_13_300 ();
 sg13g2_decap_4 FILLER_13_309 ();
 sg13g2_fill_2 FILLER_13_321 ();
 sg13g2_fill_1 FILLER_13_323 ();
 sg13g2_fill_1 FILLER_13_336 ();
 sg13g2_fill_1 FILLER_13_349 ();
 sg13g2_decap_4 FILLER_13_362 ();
 sg13g2_decap_8 FILLER_13_379 ();
 sg13g2_decap_4 FILLER_13_386 ();
 sg13g2_decap_8 FILLER_13_400 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_fill_2 FILLER_14_42 ();
 sg13g2_fill_1 FILLER_14_44 ();
 sg13g2_fill_1 FILLER_14_53 ();
 sg13g2_decap_4 FILLER_14_67 ();
 sg13g2_fill_2 FILLER_14_71 ();
 sg13g2_decap_8 FILLER_14_78 ();
 sg13g2_fill_2 FILLER_14_85 ();
 sg13g2_fill_2 FILLER_14_103 ();
 sg13g2_fill_1 FILLER_14_105 ();
 sg13g2_decap_4 FILLER_14_111 ();
 sg13g2_fill_2 FILLER_14_115 ();
 sg13g2_fill_1 FILLER_14_125 ();
 sg13g2_decap_8 FILLER_14_134 ();
 sg13g2_decap_8 FILLER_14_141 ();
 sg13g2_decap_8 FILLER_14_148 ();
 sg13g2_fill_1 FILLER_14_155 ();
 sg13g2_fill_1 FILLER_14_162 ();
 sg13g2_fill_2 FILLER_14_178 ();
 sg13g2_fill_1 FILLER_14_180 ();
 sg13g2_decap_8 FILLER_14_185 ();
 sg13g2_fill_1 FILLER_14_192 ();
 sg13g2_fill_2 FILLER_14_230 ();
 sg13g2_fill_1 FILLER_14_232 ();
 sg13g2_decap_4 FILLER_14_243 ();
 sg13g2_fill_1 FILLER_14_247 ();
 sg13g2_decap_8 FILLER_14_257 ();
 sg13g2_fill_2 FILLER_14_264 ();
 sg13g2_fill_2 FILLER_14_278 ();
 sg13g2_fill_1 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_289 ();
 sg13g2_decap_4 FILLER_14_296 ();
 sg13g2_fill_1 FILLER_14_300 ();
 sg13g2_fill_1 FILLER_14_313 ();
 sg13g2_decap_8 FILLER_14_319 ();
 sg13g2_decap_4 FILLER_14_326 ();
 sg13g2_fill_2 FILLER_14_330 ();
 sg13g2_decap_4 FILLER_14_342 ();
 sg13g2_fill_1 FILLER_14_346 ();
 sg13g2_fill_2 FILLER_14_351 ();
 sg13g2_decap_8 FILLER_14_361 ();
 sg13g2_decap_8 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_14_380 ();
 sg13g2_fill_2 FILLER_14_387 ();
 sg13g2_fill_1 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_fill_1 FILLER_15_42 ();
 sg13g2_fill_2 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_82 ();
 sg13g2_decap_8 FILLER_15_93 ();
 sg13g2_fill_2 FILLER_15_100 ();
 sg13g2_fill_1 FILLER_15_102 ();
 sg13g2_decap_4 FILLER_15_111 ();
 sg13g2_fill_2 FILLER_15_158 ();
 sg13g2_fill_2 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_186 ();
 sg13g2_decap_4 FILLER_15_193 ();
 sg13g2_decap_8 FILLER_15_201 ();
 sg13g2_decap_8 FILLER_15_208 ();
 sg13g2_decap_4 FILLER_15_215 ();
 sg13g2_fill_1 FILLER_15_219 ();
 sg13g2_fill_1 FILLER_15_225 ();
 sg13g2_decap_4 FILLER_15_236 ();
 sg13g2_fill_1 FILLER_15_240 ();
 sg13g2_decap_8 FILLER_15_262 ();
 sg13g2_decap_4 FILLER_15_269 ();
 sg13g2_fill_2 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_299 ();
 sg13g2_fill_2 FILLER_15_306 ();
 sg13g2_fill_1 FILLER_15_308 ();
 sg13g2_fill_1 FILLER_15_324 ();
 sg13g2_decap_4 FILLER_15_341 ();
 sg13g2_decap_8 FILLER_15_354 ();
 sg13g2_fill_2 FILLER_15_361 ();
 sg13g2_decap_4 FILLER_15_367 ();
 sg13g2_fill_1 FILLER_15_376 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_fill_2 FILLER_16_35 ();
 sg13g2_fill_1 FILLER_16_37 ();
 sg13g2_decap_8 FILLER_16_58 ();
 sg13g2_decap_4 FILLER_16_65 ();
 sg13g2_fill_1 FILLER_16_69 ();
 sg13g2_decap_4 FILLER_16_78 ();
 sg13g2_fill_2 FILLER_16_82 ();
 sg13g2_decap_4 FILLER_16_88 ();
 sg13g2_fill_2 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_fill_2 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_132 ();
 sg13g2_fill_1 FILLER_16_139 ();
 sg13g2_decap_8 FILLER_16_153 ();
 sg13g2_decap_8 FILLER_16_160 ();
 sg13g2_decap_8 FILLER_16_167 ();
 sg13g2_fill_2 FILLER_16_178 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_fill_2 FILLER_16_210 ();
 sg13g2_fill_1 FILLER_16_212 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_4 FILLER_16_224 ();
 sg13g2_fill_1 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_271 ();
 sg13g2_decap_8 FILLER_16_290 ();
 sg13g2_decap_4 FILLER_16_297 ();
 sg13g2_fill_2 FILLER_16_317 ();
 sg13g2_fill_1 FILLER_16_319 ();
 sg13g2_decap_4 FILLER_16_333 ();
 sg13g2_fill_2 FILLER_16_341 ();
 sg13g2_fill_2 FILLER_16_355 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_4 FILLER_17_35 ();
 sg13g2_fill_1 FILLER_17_39 ();
 sg13g2_decap_4 FILLER_17_60 ();
 sg13g2_fill_2 FILLER_17_64 ();
 sg13g2_decap_8 FILLER_17_103 ();
 sg13g2_decap_8 FILLER_17_110 ();
 sg13g2_decap_4 FILLER_17_117 ();
 sg13g2_fill_2 FILLER_17_129 ();
 sg13g2_fill_1 FILLER_17_131 ();
 sg13g2_decap_8 FILLER_17_136 ();
 sg13g2_fill_2 FILLER_17_143 ();
 sg13g2_fill_2 FILLER_17_157 ();
 sg13g2_fill_2 FILLER_17_171 ();
 sg13g2_fill_1 FILLER_17_173 ();
 sg13g2_fill_2 FILLER_17_182 ();
 sg13g2_decap_4 FILLER_17_192 ();
 sg13g2_fill_2 FILLER_17_204 ();
 sg13g2_decap_8 FILLER_17_234 ();
 sg13g2_decap_4 FILLER_17_241 ();
 sg13g2_decap_8 FILLER_17_260 ();
 sg13g2_decap_4 FILLER_17_267 ();
 sg13g2_decap_4 FILLER_17_275 ();
 sg13g2_decap_4 FILLER_17_295 ();
 sg13g2_fill_2 FILLER_17_299 ();
 sg13g2_decap_8 FILLER_17_309 ();
 sg13g2_fill_2 FILLER_17_316 ();
 sg13g2_decap_8 FILLER_17_326 ();
 sg13g2_fill_2 FILLER_17_333 ();
 sg13g2_fill_1 FILLER_17_335 ();
 sg13g2_decap_8 FILLER_17_352 ();
 sg13g2_decap_4 FILLER_17_359 ();
 sg13g2_fill_1 FILLER_17_363 ();
 sg13g2_decap_8 FILLER_17_374 ();
 sg13g2_decap_8 FILLER_17_387 ();
 sg13g2_fill_1 FILLER_17_394 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_4 FILLER_18_42 ();
 sg13g2_fill_1 FILLER_18_46 ();
 sg13g2_decap_8 FILLER_18_59 ();
 sg13g2_decap_8 FILLER_18_82 ();
 sg13g2_fill_2 FILLER_18_89 ();
 sg13g2_fill_1 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_108 ();
 sg13g2_decap_4 FILLER_18_115 ();
 sg13g2_decap_8 FILLER_18_135 ();
 sg13g2_decap_8 FILLER_18_158 ();
 sg13g2_decap_4 FILLER_18_165 ();
 sg13g2_fill_1 FILLER_18_169 ();
 sg13g2_decap_4 FILLER_18_178 ();
 sg13g2_fill_2 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_188 ();
 sg13g2_decap_8 FILLER_18_195 ();
 sg13g2_fill_1 FILLER_18_202 ();
 sg13g2_decap_8 FILLER_18_208 ();
 sg13g2_fill_2 FILLER_18_215 ();
 sg13g2_fill_2 FILLER_18_242 ();
 sg13g2_decap_4 FILLER_18_250 ();
 sg13g2_decap_8 FILLER_18_268 ();
 sg13g2_decap_8 FILLER_18_275 ();
 sg13g2_decap_8 FILLER_18_282 ();
 sg13g2_fill_1 FILLER_18_289 ();
 sg13g2_decap_8 FILLER_18_311 ();
 sg13g2_fill_1 FILLER_18_318 ();
 sg13g2_decap_8 FILLER_18_327 ();
 sg13g2_decap_8 FILLER_18_334 ();
 sg13g2_decap_8 FILLER_18_341 ();
 sg13g2_decap_8 FILLER_18_348 ();
 sg13g2_fill_2 FILLER_18_355 ();
 sg13g2_fill_1 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_4 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_62 ();
 sg13g2_fill_2 FILLER_19_69 ();
 sg13g2_fill_1 FILLER_19_71 ();
 sg13g2_decap_4 FILLER_19_104 ();
 sg13g2_fill_2 FILLER_19_108 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_4 FILLER_19_156 ();
 sg13g2_fill_1 FILLER_19_180 ();
 sg13g2_decap_4 FILLER_19_212 ();
 sg13g2_fill_2 FILLER_19_216 ();
 sg13g2_decap_4 FILLER_19_237 ();
 sg13g2_fill_2 FILLER_19_241 ();
 sg13g2_fill_1 FILLER_19_249 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_fill_2 FILLER_19_284 ();
 sg13g2_fill_2 FILLER_19_304 ();
 sg13g2_fill_1 FILLER_19_318 ();
 sg13g2_decap_4 FILLER_19_360 ();
 sg13g2_fill_2 FILLER_19_368 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_4 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_58 ();
 sg13g2_fill_2 FILLER_20_65 ();
 sg13g2_decap_8 FILLER_20_75 ();
 sg13g2_decap_8 FILLER_20_82 ();
 sg13g2_decap_8 FILLER_20_89 ();
 sg13g2_decap_8 FILLER_20_100 ();
 sg13g2_fill_2 FILLER_20_107 ();
 sg13g2_fill_1 FILLER_20_117 ();
 sg13g2_decap_8 FILLER_20_134 ();
 sg13g2_fill_2 FILLER_20_141 ();
 sg13g2_decap_8 FILLER_20_151 ();
 sg13g2_fill_2 FILLER_20_158 ();
 sg13g2_fill_1 FILLER_20_160 ();
 sg13g2_decap_8 FILLER_20_177 ();
 sg13g2_decap_4 FILLER_20_184 ();
 sg13g2_fill_1 FILLER_20_188 ();
 sg13g2_decap_8 FILLER_20_194 ();
 sg13g2_decap_8 FILLER_20_206 ();
 sg13g2_fill_2 FILLER_20_213 ();
 sg13g2_fill_1 FILLER_20_215 ();
 sg13g2_fill_2 FILLER_20_220 ();
 sg13g2_fill_1 FILLER_20_222 ();
 sg13g2_decap_8 FILLER_20_228 ();
 sg13g2_decap_4 FILLER_20_235 ();
 sg13g2_fill_2 FILLER_20_239 ();
 sg13g2_fill_1 FILLER_20_253 ();
 sg13g2_fill_2 FILLER_20_258 ();
 sg13g2_fill_1 FILLER_20_260 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_fill_1 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_299 ();
 sg13g2_fill_2 FILLER_20_306 ();
 sg13g2_decap_8 FILLER_20_320 ();
 sg13g2_fill_1 FILLER_20_327 ();
 sg13g2_fill_2 FILLER_20_337 ();
 sg13g2_fill_1 FILLER_20_339 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_4 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_54 ();
 sg13g2_fill_2 FILLER_21_61 ();
 sg13g2_fill_2 FILLER_21_79 ();
 sg13g2_fill_1 FILLER_21_81 ();
 sg13g2_fill_2 FILLER_21_90 ();
 sg13g2_decap_8 FILLER_21_104 ();
 sg13g2_decap_4 FILLER_21_111 ();
 sg13g2_fill_1 FILLER_21_123 ();
 sg13g2_fill_1 FILLER_21_128 ();
 sg13g2_fill_2 FILLER_21_141 ();
 sg13g2_decap_8 FILLER_21_151 ();
 sg13g2_decap_4 FILLER_21_158 ();
 sg13g2_fill_1 FILLER_21_162 ();
 sg13g2_decap_8 FILLER_21_171 ();
 sg13g2_decap_8 FILLER_21_178 ();
 sg13g2_fill_2 FILLER_21_185 ();
 sg13g2_fill_2 FILLER_21_211 ();
 sg13g2_fill_1 FILLER_21_213 ();
 sg13g2_fill_1 FILLER_21_224 ();
 sg13g2_fill_2 FILLER_21_254 ();
 sg13g2_fill_2 FILLER_21_262 ();
 sg13g2_fill_2 FILLER_21_277 ();
 sg13g2_fill_1 FILLER_21_279 ();
 sg13g2_decap_4 FILLER_21_301 ();
 sg13g2_fill_2 FILLER_21_329 ();
 sg13g2_fill_1 FILLER_21_331 ();
 sg13g2_fill_2 FILLER_21_340 ();
 sg13g2_fill_1 FILLER_21_342 ();
 sg13g2_fill_2 FILLER_21_352 ();
 sg13g2_fill_1 FILLER_21_358 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_decap_8 FILLER_21_375 ();
 sg13g2_fill_2 FILLER_21_382 ();
 sg13g2_fill_1 FILLER_21_384 ();
 sg13g2_decap_8 FILLER_21_398 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_4 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_54 ();
 sg13g2_decap_8 FILLER_22_61 ();
 sg13g2_fill_1 FILLER_22_68 ();
 sg13g2_fill_1 FILLER_22_73 ();
 sg13g2_decap_8 FILLER_22_79 ();
 sg13g2_fill_2 FILLER_22_86 ();
 sg13g2_fill_1 FILLER_22_88 ();
 sg13g2_decap_8 FILLER_22_109 ();
 sg13g2_fill_2 FILLER_22_116 ();
 sg13g2_fill_2 FILLER_22_126 ();
 sg13g2_fill_1 FILLER_22_128 ();
 sg13g2_decap_4 FILLER_22_153 ();
 sg13g2_fill_2 FILLER_22_157 ();
 sg13g2_decap_4 FILLER_22_179 ();
 sg13g2_fill_1 FILLER_22_183 ();
 sg13g2_decap_8 FILLER_22_200 ();
 sg13g2_fill_2 FILLER_22_207 ();
 sg13g2_decap_8 FILLER_22_220 ();
 sg13g2_decap_8 FILLER_22_227 ();
 sg13g2_decap_4 FILLER_22_234 ();
 sg13g2_fill_2 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_253 ();
 sg13g2_decap_8 FILLER_22_260 ();
 sg13g2_fill_2 FILLER_22_280 ();
 sg13g2_fill_1 FILLER_22_282 ();
 sg13g2_decap_8 FILLER_22_306 ();
 sg13g2_fill_1 FILLER_22_313 ();
 sg13g2_decap_8 FILLER_22_319 ();
 sg13g2_decap_4 FILLER_22_326 ();
 sg13g2_fill_1 FILLER_22_330 ();
 sg13g2_decap_4 FILLER_22_364 ();
 sg13g2_fill_1 FILLER_22_368 ();
 sg13g2_fill_2 FILLER_22_378 ();
 sg13g2_fill_1 FILLER_22_380 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_29 ();
 sg13g2_decap_8 FILLER_23_36 ();
 sg13g2_decap_8 FILLER_23_86 ();
 sg13g2_decap_4 FILLER_23_93 ();
 sg13g2_fill_2 FILLER_23_97 ();
 sg13g2_decap_8 FILLER_23_107 ();
 sg13g2_decap_4 FILLER_23_114 ();
 sg13g2_fill_2 FILLER_23_118 ();
 sg13g2_fill_2 FILLER_23_128 ();
 sg13g2_fill_1 FILLER_23_130 ();
 sg13g2_decap_8 FILLER_23_139 ();
 sg13g2_decap_8 FILLER_23_146 ();
 sg13g2_decap_8 FILLER_23_153 ();
 sg13g2_fill_2 FILLER_23_160 ();
 sg13g2_fill_1 FILLER_23_162 ();
 sg13g2_decap_8 FILLER_23_171 ();
 sg13g2_decap_4 FILLER_23_178 ();
 sg13g2_fill_1 FILLER_23_182 ();
 sg13g2_decap_4 FILLER_23_187 ();
 sg13g2_decap_8 FILLER_23_195 ();
 sg13g2_decap_8 FILLER_23_202 ();
 sg13g2_fill_2 FILLER_23_209 ();
 sg13g2_decap_8 FILLER_23_220 ();
 sg13g2_decap_4 FILLER_23_239 ();
 sg13g2_fill_1 FILLER_23_243 ();
 sg13g2_fill_2 FILLER_23_250 ();
 sg13g2_decap_4 FILLER_23_264 ();
 sg13g2_fill_2 FILLER_23_268 ();
 sg13g2_decap_8 FILLER_23_275 ();
 sg13g2_decap_8 FILLER_23_282 ();
 sg13g2_fill_2 FILLER_23_289 ();
 sg13g2_decap_8 FILLER_23_299 ();
 sg13g2_decap_4 FILLER_23_306 ();
 sg13g2_decap_4 FILLER_23_322 ();
 sg13g2_fill_2 FILLER_23_326 ();
 sg13g2_fill_1 FILLER_23_337 ();
 sg13g2_fill_2 FILLER_23_349 ();
 sg13g2_fill_2 FILLER_23_360 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_4 ();
 sg13g2_fill_1 FILLER_24_13 ();
 sg13g2_decap_8 FILLER_24_31 ();
 sg13g2_decap_4 FILLER_24_38 ();
 sg13g2_fill_1 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_51 ();
 sg13g2_decap_8 FILLER_24_58 ();
 sg13g2_fill_2 FILLER_24_65 ();
 sg13g2_fill_1 FILLER_24_67 ();
 sg13g2_fill_2 FILLER_24_72 ();
 sg13g2_fill_1 FILLER_24_82 ();
 sg13g2_decap_8 FILLER_24_87 ();
 sg13g2_decap_8 FILLER_24_94 ();
 sg13g2_decap_4 FILLER_24_101 ();
 sg13g2_fill_2 FILLER_24_105 ();
 sg13g2_fill_2 FILLER_24_123 ();
 sg13g2_fill_1 FILLER_24_125 ();
 sg13g2_decap_4 FILLER_24_134 ();
 sg13g2_fill_1 FILLER_24_154 ();
 sg13g2_fill_2 FILLER_24_171 ();
 sg13g2_fill_1 FILLER_24_173 ();
 sg13g2_decap_4 FILLER_24_198 ();
 sg13g2_fill_1 FILLER_24_202 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_fill_2 FILLER_24_231 ();
 sg13g2_fill_1 FILLER_24_238 ();
 sg13g2_decap_4 FILLER_24_259 ();
 sg13g2_fill_1 FILLER_24_263 ();
 sg13g2_decap_4 FILLER_24_284 ();
 sg13g2_fill_2 FILLER_24_288 ();
 sg13g2_fill_1 FILLER_24_294 ();
 sg13g2_fill_2 FILLER_24_307 ();
 sg13g2_fill_1 FILLER_24_309 ();
 sg13g2_fill_2 FILLER_24_360 ();
 sg13g2_fill_1 FILLER_24_375 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_4 ();
 sg13g2_fill_2 FILLER_25_14 ();
 sg13g2_fill_1 FILLER_25_16 ();
 sg13g2_fill_2 FILLER_25_34 ();
 sg13g2_fill_1 FILLER_25_45 ();
 sg13g2_decap_4 FILLER_25_54 ();
 sg13g2_fill_2 FILLER_25_74 ();
 sg13g2_decap_4 FILLER_25_92 ();
 sg13g2_decap_4 FILLER_25_112 ();
 sg13g2_decap_4 FILLER_25_132 ();
 sg13g2_fill_1 FILLER_25_136 ();
 sg13g2_decap_8 FILLER_25_145 ();
 sg13g2_decap_4 FILLER_25_152 ();
 sg13g2_fill_2 FILLER_25_156 ();
 sg13g2_decap_4 FILLER_25_174 ();
 sg13g2_fill_1 FILLER_25_178 ();
 sg13g2_decap_4 FILLER_25_187 ();
 sg13g2_decap_8 FILLER_25_195 ();
 sg13g2_decap_8 FILLER_25_202 ();
 sg13g2_decap_4 FILLER_25_209 ();
 sg13g2_fill_1 FILLER_25_213 ();
 sg13g2_fill_2 FILLER_25_218 ();
 sg13g2_fill_1 FILLER_25_225 ();
 sg13g2_decap_8 FILLER_25_230 ();
 sg13g2_decap_8 FILLER_25_237 ();
 sg13g2_decap_4 FILLER_25_244 ();
 sg13g2_fill_1 FILLER_25_248 ();
 sg13g2_decap_4 FILLER_25_253 ();
 sg13g2_fill_1 FILLER_25_257 ();
 sg13g2_fill_2 FILLER_25_262 ();
 sg13g2_fill_1 FILLER_25_264 ();
 sg13g2_decap_4 FILLER_25_279 ();
 sg13g2_fill_1 FILLER_25_283 ();
 sg13g2_fill_2 FILLER_25_317 ();
 sg13g2_fill_1 FILLER_25_319 ();
 sg13g2_fill_2 FILLER_25_328 ();
 sg13g2_fill_2 FILLER_25_335 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_9 ();
 sg13g2_decap_8 FILLER_26_31 ();
 sg13g2_fill_1 FILLER_26_38 ();
 sg13g2_fill_1 FILLER_26_44 ();
 sg13g2_fill_2 FILLER_26_52 ();
 sg13g2_fill_1 FILLER_26_54 ();
 sg13g2_decap_8 FILLER_26_65 ();
 sg13g2_decap_8 FILLER_26_72 ();
 sg13g2_decap_4 FILLER_26_83 ();
 sg13g2_fill_2 FILLER_26_87 ();
 sg13g2_decap_8 FILLER_26_113 ();
 sg13g2_decap_4 FILLER_26_120 ();
 sg13g2_decap_8 FILLER_26_148 ();
 sg13g2_decap_8 FILLER_26_155 ();
 sg13g2_fill_2 FILLER_26_162 ();
 sg13g2_fill_1 FILLER_26_164 ();
 sg13g2_fill_1 FILLER_26_173 ();
 sg13g2_decap_8 FILLER_26_179 ();
 sg13g2_fill_1 FILLER_26_214 ();
 sg13g2_decap_4 FILLER_26_285 ();
 sg13g2_fill_2 FILLER_26_289 ();
 sg13g2_decap_4 FILLER_26_299 ();
 sg13g2_fill_2 FILLER_26_303 ();
 sg13g2_fill_2 FILLER_26_314 ();
 sg13g2_decap_8 FILLER_26_324 ();
 sg13g2_fill_2 FILLER_26_331 ();
 sg13g2_decap_4 FILLER_26_363 ();
 sg13g2_decap_4 FILLER_26_371 ();
 sg13g2_fill_2 FILLER_26_384 ();
 sg13g2_fill_1 FILLER_26_386 ();
 sg13g2_fill_2 FILLER_26_391 ();
 sg13g2_fill_1 FILLER_26_393 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_4 ();
 sg13g2_fill_2 FILLER_27_15 ();
 sg13g2_decap_8 FILLER_27_25 ();
 sg13g2_decap_4 FILLER_27_32 ();
 sg13g2_fill_2 FILLER_27_36 ();
 sg13g2_decap_4 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_86 ();
 sg13g2_fill_1 FILLER_27_93 ();
 sg13g2_decap_4 FILLER_27_110 ();
 sg13g2_decap_8 FILLER_27_132 ();
 sg13g2_fill_2 FILLER_27_139 ();
 sg13g2_fill_1 FILLER_27_141 ();
 sg13g2_decap_4 FILLER_27_158 ();
 sg13g2_decap_8 FILLER_27_185 ();
 sg13g2_decap_4 FILLER_27_192 ();
 sg13g2_fill_2 FILLER_27_210 ();
 sg13g2_fill_1 FILLER_27_212 ();
 sg13g2_fill_1 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_222 ();
 sg13g2_decap_4 FILLER_27_229 ();
 sg13g2_decap_4 FILLER_27_242 ();
 sg13g2_fill_2 FILLER_27_246 ();
 sg13g2_fill_1 FILLER_27_253 ();
 sg13g2_fill_2 FILLER_27_272 ();
 sg13g2_fill_1 FILLER_27_274 ();
 sg13g2_fill_2 FILLER_27_284 ();
 sg13g2_fill_1 FILLER_27_286 ();
 sg13g2_decap_4 FILLER_27_320 ();
 sg13g2_fill_1 FILLER_27_324 ();
 sg13g2_decap_4 FILLER_27_369 ();
 sg13g2_fill_1 FILLER_27_373 ();
 sg13g2_fill_2 FILLER_27_378 ();
 sg13g2_fill_1 FILLER_27_380 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_12 ();
 sg13g2_fill_1 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_34 ();
 sg13g2_decap_8 FILLER_28_41 ();
 sg13g2_decap_8 FILLER_28_48 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_fill_2 FILLER_28_77 ();
 sg13g2_fill_1 FILLER_28_79 ();
 sg13g2_decap_8 FILLER_28_88 ();
 sg13g2_fill_1 FILLER_28_95 ();
 sg13g2_decap_8 FILLER_28_104 ();
 sg13g2_decap_8 FILLER_28_111 ();
 sg13g2_decap_8 FILLER_28_134 ();
 sg13g2_decap_4 FILLER_28_141 ();
 sg13g2_fill_1 FILLER_28_145 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_fill_2 FILLER_28_168 ();
 sg13g2_fill_1 FILLER_28_170 ();
 sg13g2_decap_4 FILLER_28_186 ();
 sg13g2_fill_2 FILLER_28_190 ();
 sg13g2_fill_2 FILLER_28_219 ();
 sg13g2_fill_1 FILLER_28_221 ();
 sg13g2_decap_4 FILLER_28_290 ();
 sg13g2_decap_4 FILLER_28_302 ();
 sg13g2_fill_2 FILLER_28_306 ();
 sg13g2_decap_8 FILLER_28_321 ();
 sg13g2_decap_4 FILLER_28_328 ();
 sg13g2_fill_1 FILLER_28_341 ();
 sg13g2_decap_4 FILLER_28_360 ();
 sg13g2_decap_4 FILLER_28_372 ();
 sg13g2_fill_2 FILLER_28_376 ();
 sg13g2_decap_4 FILLER_28_389 ();
 sg13g2_decap_8 FILLER_28_402 ();
 sg13g2_fill_2 FILLER_29_16 ();
 sg13g2_fill_1 FILLER_29_18 ();
 sg13g2_decap_8 FILLER_29_23 ();
 sg13g2_fill_2 FILLER_29_30 ();
 sg13g2_fill_2 FILLER_29_40 ();
 sg13g2_fill_1 FILLER_29_42 ();
 sg13g2_decap_4 FILLER_29_47 ();
 sg13g2_fill_1 FILLER_29_51 ();
 sg13g2_decap_4 FILLER_29_70 ();
 sg13g2_fill_1 FILLER_29_74 ();
 sg13g2_fill_2 FILLER_29_80 ();
 sg13g2_fill_2 FILLER_29_86 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_fill_2 FILLER_29_119 ();
 sg13g2_fill_1 FILLER_29_121 ();
 sg13g2_fill_2 FILLER_29_141 ();
 sg13g2_fill_1 FILLER_29_164 ();
 sg13g2_fill_2 FILLER_29_173 ();
 sg13g2_fill_2 FILLER_29_181 ();
 sg13g2_decap_4 FILLER_29_193 ();
 sg13g2_fill_1 FILLER_29_197 ();
 sg13g2_decap_8 FILLER_29_202 ();
 sg13g2_decap_8 FILLER_29_209 ();
 sg13g2_decap_4 FILLER_29_216 ();
 sg13g2_fill_2 FILLER_29_233 ();
 sg13g2_decap_8 FILLER_29_244 ();
 sg13g2_fill_1 FILLER_29_256 ();
 sg13g2_fill_2 FILLER_29_270 ();
 sg13g2_decap_8 FILLER_29_288 ();
 sg13g2_fill_2 FILLER_29_295 ();
 sg13g2_fill_1 FILLER_29_297 ();
 sg13g2_decap_8 FILLER_29_335 ();
 sg13g2_fill_1 FILLER_29_342 ();
 sg13g2_fill_1 FILLER_29_347 ();
 sg13g2_decap_8 FILLER_29_353 ();
 sg13g2_decap_4 FILLER_29_360 ();
 sg13g2_fill_2 FILLER_29_372 ();
 sg13g2_fill_1 FILLER_29_374 ();
 sg13g2_fill_1 FILLER_29_380 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_4 FILLER_30_29 ();
 sg13g2_fill_1 FILLER_30_33 ();
 sg13g2_fill_2 FILLER_30_42 ();
 sg13g2_fill_1 FILLER_30_44 ();
 sg13g2_fill_2 FILLER_30_53 ();
 sg13g2_decap_4 FILLER_30_72 ();
 sg13g2_decap_4 FILLER_30_92 ();
 sg13g2_fill_2 FILLER_30_96 ();
 sg13g2_decap_8 FILLER_30_106 ();
 sg13g2_decap_8 FILLER_30_113 ();
 sg13g2_decap_4 FILLER_30_120 ();
 sg13g2_fill_1 FILLER_30_124 ();
 sg13g2_fill_1 FILLER_30_131 ();
 sg13g2_decap_8 FILLER_30_137 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_fill_2 FILLER_30_161 ();
 sg13g2_fill_2 FILLER_30_169 ();
 sg13g2_fill_1 FILLER_30_171 ();
 sg13g2_decap_8 FILLER_30_177 ();
 sg13g2_decap_4 FILLER_30_184 ();
 sg13g2_fill_2 FILLER_30_218 ();
 sg13g2_fill_1 FILLER_30_220 ();
 sg13g2_fill_1 FILLER_30_249 ();
 sg13g2_decap_4 FILLER_30_278 ();
 sg13g2_fill_2 FILLER_30_282 ();
 sg13g2_decap_4 FILLER_30_293 ();
 sg13g2_decap_4 FILLER_30_306 ();
 sg13g2_fill_2 FILLER_30_310 ();
 sg13g2_fill_1 FILLER_30_338 ();
 sg13g2_fill_1 FILLER_30_371 ();
 sg13g2_decap_4 FILLER_30_382 ();
 sg13g2_fill_1 FILLER_30_386 ();
 sg13g2_fill_1 FILLER_30_391 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_14 ();
 sg13g2_decap_4 FILLER_31_31 ();
 sg13g2_fill_2 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_41 ();
 sg13g2_fill_2 FILLER_31_48 ();
 sg13g2_fill_2 FILLER_31_58 ();
 sg13g2_decap_8 FILLER_31_76 ();
 sg13g2_decap_8 FILLER_31_83 ();
 sg13g2_fill_2 FILLER_31_90 ();
 sg13g2_decap_8 FILLER_31_100 ();
 sg13g2_fill_1 FILLER_31_107 ();
 sg13g2_fill_2 FILLER_31_136 ();
 sg13g2_fill_1 FILLER_31_138 ();
 sg13g2_fill_1 FILLER_31_195 ();
 sg13g2_decap_8 FILLER_31_205 ();
 sg13g2_decap_8 FILLER_31_212 ();
 sg13g2_fill_2 FILLER_31_232 ();
 sg13g2_fill_2 FILLER_31_243 ();
 sg13g2_fill_1 FILLER_31_253 ();
 sg13g2_decap_4 FILLER_31_276 ();
 sg13g2_fill_2 FILLER_31_280 ();
 sg13g2_fill_2 FILLER_31_310 ();
 sg13g2_fill_1 FILLER_31_345 ();
 sg13g2_decap_4 FILLER_31_371 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_4 ();
 sg13g2_fill_1 FILLER_32_13 ();
 sg13g2_decap_4 FILLER_32_28 ();
 sg13g2_fill_1 FILLER_32_32 ();
 sg13g2_decap_8 FILLER_32_47 ();
 sg13g2_decap_4 FILLER_32_54 ();
 sg13g2_fill_1 FILLER_32_58 ();
 sg13g2_decap_8 FILLER_32_67 ();
 sg13g2_fill_2 FILLER_32_74 ();
 sg13g2_fill_1 FILLER_32_76 ();
 sg13g2_decap_8 FILLER_32_93 ();
 sg13g2_decap_8 FILLER_32_100 ();
 sg13g2_decap_8 FILLER_32_107 ();
 sg13g2_decap_4 FILLER_32_118 ();
 sg13g2_fill_2 FILLER_32_122 ();
 sg13g2_fill_2 FILLER_32_144 ();
 sg13g2_fill_1 FILLER_32_146 ();
 sg13g2_decap_4 FILLER_32_160 ();
 sg13g2_decap_4 FILLER_32_175 ();
 sg13g2_fill_1 FILLER_32_179 ();
 sg13g2_fill_1 FILLER_32_183 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_fill_2 FILLER_32_210 ();
 sg13g2_fill_1 FILLER_32_220 ();
 sg13g2_decap_4 FILLER_32_227 ();
 sg13g2_fill_1 FILLER_32_244 ();
 sg13g2_fill_1 FILLER_32_258 ();
 sg13g2_fill_1 FILLER_32_291 ();
 sg13g2_decap_4 FILLER_32_301 ();
 sg13g2_fill_2 FILLER_32_305 ();
 sg13g2_decap_4 FILLER_32_320 ();
 sg13g2_fill_2 FILLER_32_324 ();
 sg13g2_fill_1 FILLER_32_340 ();
 sg13g2_fill_1 FILLER_32_344 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_4 FILLER_33_14 ();
 sg13g2_fill_2 FILLER_33_18 ();
 sg13g2_fill_2 FILLER_33_28 ();
 sg13g2_decap_4 FILLER_33_46 ();
 sg13g2_fill_2 FILLER_33_50 ();
 sg13g2_fill_1 FILLER_33_60 ();
 sg13g2_decap_4 FILLER_33_85 ();
 sg13g2_fill_2 FILLER_33_89 ();
 sg13g2_decap_8 FILLER_33_153 ();
 sg13g2_decap_4 FILLER_33_160 ();
 sg13g2_fill_2 FILLER_33_164 ();
 sg13g2_fill_2 FILLER_33_172 ();
 sg13g2_fill_1 FILLER_33_174 ();
 sg13g2_decap_4 FILLER_33_193 ();
 sg13g2_fill_1 FILLER_33_210 ();
 sg13g2_decap_4 FILLER_33_228 ();
 sg13g2_fill_1 FILLER_33_232 ();
 sg13g2_fill_2 FILLER_33_249 ();
 sg13g2_decap_4 FILLER_33_260 ();
 sg13g2_fill_1 FILLER_33_268 ();
 sg13g2_fill_2 FILLER_33_278 ();
 sg13g2_fill_2 FILLER_33_321 ();
 sg13g2_fill_2 FILLER_33_360 ();
 sg13g2_fill_2 FILLER_33_372 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_4 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_92 ();
 sg13g2_decap_4 FILLER_34_99 ();
 sg13g2_fill_1 FILLER_34_103 ();
 sg13g2_decap_4 FILLER_34_124 ();
 sg13g2_fill_2 FILLER_34_128 ();
 sg13g2_fill_1 FILLER_34_173 ();
 sg13g2_decap_8 FILLER_34_200 ();
 sg13g2_decap_8 FILLER_34_207 ();
 sg13g2_fill_2 FILLER_34_214 ();
 sg13g2_decap_4 FILLER_34_221 ();
 sg13g2_fill_1 FILLER_34_225 ();
 sg13g2_fill_1 FILLER_34_243 ();
 sg13g2_decap_8 FILLER_34_269 ();
 sg13g2_decap_4 FILLER_34_281 ();
 sg13g2_fill_1 FILLER_34_285 ();
 sg13g2_fill_2 FILLER_34_299 ();
 sg13g2_fill_1 FILLER_34_323 ();
 sg13g2_fill_2 FILLER_34_338 ();
 sg13g2_fill_1 FILLER_34_340 ();
 sg13g2_fill_1 FILLER_34_354 ();
 sg13g2_fill_2 FILLER_34_363 ();
 sg13g2_fill_2 FILLER_34_392 ();
 sg13g2_fill_1 FILLER_34_394 ();
 sg13g2_decap_4 FILLER_34_404 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_fill_1 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_101 ();
 sg13g2_decap_8 FILLER_35_108 ();
 sg13g2_fill_2 FILLER_35_115 ();
 sg13g2_decap_4 FILLER_35_121 ();
 sg13g2_fill_1 FILLER_35_125 ();
 sg13g2_fill_1 FILLER_35_146 ();
 sg13g2_fill_2 FILLER_35_153 ();
 sg13g2_fill_2 FILLER_35_170 ();
 sg13g2_fill_1 FILLER_35_172 ();
 sg13g2_fill_2 FILLER_35_183 ();
 sg13g2_fill_1 FILLER_35_185 ();
 sg13g2_decap_4 FILLER_35_218 ();
 sg13g2_fill_1 FILLER_35_249 ();
 sg13g2_fill_2 FILLER_35_267 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_fill_2 FILLER_36_139 ();
 sg13g2_fill_1 FILLER_36_150 ();
 sg13g2_fill_2 FILLER_36_166 ();
 sg13g2_fill_1 FILLER_36_209 ();
 sg13g2_decap_8 FILLER_36_239 ();
 sg13g2_fill_2 FILLER_36_246 ();
 sg13g2_fill_1 FILLER_36_248 ();
 sg13g2_fill_2 FILLER_36_254 ();
 sg13g2_fill_2 FILLER_36_264 ();
 sg13g2_decap_4 FILLER_36_270 ();
 sg13g2_fill_2 FILLER_36_274 ();
 sg13g2_fill_1 FILLER_36_286 ();
 sg13g2_fill_2 FILLER_36_291 ();
 sg13g2_fill_2 FILLER_36_302 ();
 sg13g2_fill_1 FILLER_36_304 ();
 sg13g2_fill_2 FILLER_36_330 ();
 sg13g2_fill_1 FILLER_36_332 ();
 sg13g2_fill_1 FILLER_36_365 ();
 sg13g2_fill_2 FILLER_36_372 ();
 sg13g2_fill_2 FILLER_36_379 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_4 FILLER_37_119 ();
 sg13g2_fill_2 FILLER_37_123 ();
 sg13g2_fill_1 FILLER_37_152 ();
 sg13g2_fill_2 FILLER_37_203 ();
 sg13g2_fill_1 FILLER_37_205 ();
 sg13g2_fill_2 FILLER_37_265 ();
 sg13g2_fill_1 FILLER_37_298 ();
 sg13g2_fill_2 FILLER_37_326 ();
 sg13g2_fill_1 FILLER_37_328 ();
 sg13g2_fill_1 FILLER_37_334 ();
 sg13g2_fill_2 FILLER_37_344 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_fill_1 FILLER_38_124 ();
 sg13g2_fill_2 FILLER_38_141 ();
 sg13g2_fill_1 FILLER_38_143 ();
 sg13g2_fill_1 FILLER_38_148 ();
 sg13g2_fill_2 FILLER_38_157 ();
 sg13g2_fill_1 FILLER_38_159 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_fill_1 FILLER_38_180 ();
 sg13g2_fill_1 FILLER_38_190 ();
 sg13g2_decap_4 FILLER_38_195 ();
 sg13g2_fill_2 FILLER_38_199 ();
 sg13g2_fill_1 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_decap_4 FILLER_38_222 ();
 sg13g2_fill_1 FILLER_38_226 ();
 sg13g2_fill_1 FILLER_38_236 ();
 sg13g2_decap_4 FILLER_38_241 ();
 sg13g2_fill_2 FILLER_38_245 ();
 sg13g2_decap_4 FILLER_38_256 ();
 sg13g2_fill_2 FILLER_38_269 ();
 sg13g2_fill_1 FILLER_38_271 ();
 sg13g2_fill_2 FILLER_38_319 ();
 sg13g2_fill_1 FILLER_38_321 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net14;
 assign uio_oe[1] = net15;
 assign uio_oe[2] = net16;
 assign uio_oe[3] = net17;
 assign uio_oe[4] = net18;
 assign uio_oe[5] = net19;
 assign uio_oe[6] = net20;
 assign uio_oe[7] = net21;
 assign uio_out[0] = net22;
 assign uio_out[1] = net23;
 assign uio_out[2] = net24;
 assign uio_out[3] = net25;
 assign uio_out[4] = net26;
 assign uio_out[5] = net27;
 assign uio_out[6] = net28;
 assign uio_out[7] = net29;
endmodule
