module tt_um_MichaelBell_photo_frame (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire clk_regs;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire \addr_in[0] ;
 wire \addr_in[10] ;
 wire \addr_in[11] ;
 wire \addr_in[12] ;
 wire \addr_in[13] ;
 wire \addr_in[14] ;
 wire \addr_in[15] ;
 wire \addr_in[16] ;
 wire \addr_in[17] ;
 wire \addr_in[18] ;
 wire \addr_in[19] ;
 wire \addr_in[1] ;
 wire \addr_in[20] ;
 wire \addr_in[21] ;
 wire \addr_in[22] ;
 wire \addr_in[23] ;
 wire \addr_in[2] ;
 wire \addr_in[3] ;
 wire \addr_in[4] ;
 wire \addr_in[5] ;
 wire \addr_in[6] ;
 wire \addr_in[7] ;
 wire \addr_in[8] ;
 wire \addr_in[9] ;
 wire hsync;
 wire hsync_r;
 wire \i_display.cfg[0] ;
 wire \i_display.cfg[10] ;
 wire \i_display.cfg[11] ;
 wire \i_display.cfg[12] ;
 wire \i_display.cfg[13] ;
 wire \i_display.cfg[14] ;
 wire \i_display.cfg[15] ;
 wire \i_display.cfg[16] ;
 wire \i_display.cfg[17] ;
 wire \i_display.cfg[18] ;
 wire \i_display.cfg[19] ;
 wire \i_display.cfg[1] ;
 wire \i_display.cfg[20] ;
 wire \i_display.cfg[21] ;
 wire \i_display.cfg[22] ;
 wire \i_display.cfg[23] ;
 wire \i_display.cfg[24] ;
 wire \i_display.cfg[25] ;
 wire \i_display.cfg[26] ;
 wire \i_display.cfg[27] ;
 wire \i_display.cfg[28] ;
 wire \i_display.cfg[29] ;
 wire \i_display.cfg[2] ;
 wire \i_display.cfg[30] ;
 wire \i_display.cfg[31] ;
 wire \i_display.cfg[32] ;
 wire \i_display.cfg[33] ;
 wire \i_display.cfg[34] ;
 wire \i_display.cfg[35] ;
 wire \i_display.cfg[36] ;
 wire \i_display.cfg[37] ;
 wire \i_display.cfg[38] ;
 wire \i_display.cfg[39] ;
 wire \i_display.cfg[3] ;
 wire \i_display.cfg[40] ;
 wire \i_display.cfg[41] ;
 wire \i_display.cfg[42] ;
 wire \i_display.cfg[43] ;
 wire \i_display.cfg[44] ;
 wire \i_display.cfg[45] ;
 wire \i_display.cfg[46] ;
 wire \i_display.cfg[47] ;
 wire \i_display.cfg[48] ;
 wire \i_display.cfg[49] ;
 wire \i_display.cfg[4] ;
 wire \i_display.cfg[50] ;
 wire \i_display.cfg[51] ;
 wire \i_display.cfg[52] ;
 wire \i_display.cfg[53] ;
 wire \i_display.cfg[54] ;
 wire \i_display.cfg[55] ;
 wire \i_display.cfg[56] ;
 wire \i_display.cfg[57] ;
 wire \i_display.cfg[58] ;
 wire \i_display.cfg[59] ;
 wire \i_display.cfg[5] ;
 wire \i_display.cfg[60] ;
 wire \i_display.cfg[61] ;
 wire \i_display.cfg[62] ;
 wire \i_display.cfg[63] ;
 wire \i_display.cfg[64] ;
 wire \i_display.cfg[65] ;
 wire \i_display.cfg[66] ;
 wire \i_display.cfg[67] ;
 wire \i_display.cfg[68] ;
 wire \i_display.cfg[69] ;
 wire \i_display.cfg[6] ;
 wire \i_display.cfg[70] ;
 wire \i_display.cfg[71] ;
 wire \i_display.cfg[72] ;
 wire \i_display.cfg[73] ;
 wire \i_display.cfg[74] ;
 wire \i_display.cfg[7] ;
 wire \i_display.cfg[8] ;
 wire \i_display.cfg[9] ;
 wire \i_display.cfg_clk_sync[0] ;
 wire \i_display.cfg_clk_sync[1] ;
 wire \i_display.cfg_clk_sync[2] ;
 wire \i_display.cfg_data_sync[0] ;
 wire \i_display.cfg_data_sync[1] ;
 wire \i_display.h_count[0] ;
 wire \i_display.h_count[10] ;
 wire \i_display.h_count[1] ;
 wire \i_display.h_count[2] ;
 wire \i_display.h_count[3] ;
 wire \i_display.h_count[4] ;
 wire \i_display.h_count[5] ;
 wire \i_display.h_count[6] ;
 wire \i_display.h_count[7] ;
 wire \i_display.h_count[8] ;
 wire \i_display.h_count[9] ;
 wire \i_display.h_state[0] ;
 wire \i_display.h_state[1] ;
 wire \i_display.v_count[0] ;
 wire \i_display.v_count[10] ;
 wire \i_display.v_count[1] ;
 wire \i_display.v_count[2] ;
 wire \i_display.v_count[3] ;
 wire \i_display.v_count[4] ;
 wire \i_display.v_count[5] ;
 wire \i_display.v_count[6] ;
 wire \i_display.v_count[7] ;
 wire \i_display.v_count[8] ;
 wire \i_display.v_count[9] ;
 wire \i_display.v_state[0] ;
 wire \i_display.v_state[1] ;
 wire \i_display.vsync ;
 wire \i_qpsi.addr[0] ;
 wire \i_qpsi.addr[10] ;
 wire \i_qpsi.addr[11] ;
 wire \i_qpsi.addr[12] ;
 wire \i_qpsi.addr[13] ;
 wire \i_qpsi.addr[14] ;
 wire \i_qpsi.addr[15] ;
 wire \i_qpsi.addr[16] ;
 wire \i_qpsi.addr[17] ;
 wire \i_qpsi.addr[18] ;
 wire \i_qpsi.addr[19] ;
 wire \i_qpsi.addr[1] ;
 wire \i_qpsi.addr[20] ;
 wire \i_qpsi.addr[21] ;
 wire \i_qpsi.addr[22] ;
 wire \i_qpsi.addr[23] ;
 wire \i_qpsi.addr[2] ;
 wire \i_qpsi.addr[3] ;
 wire \i_qpsi.addr[4] ;
 wire \i_qpsi.addr[5] ;
 wire \i_qpsi.addr[6] ;
 wire \i_qpsi.addr[7] ;
 wire \i_qpsi.addr[8] ;
 wire \i_qpsi.addr[9] ;
 wire \i_qpsi.bits_remaining[0] ;
 wire \i_qpsi.bits_remaining[1] ;
 wire \i_qpsi.bits_remaining[2] ;
 wire \i_qpsi.data[0] ;
 wire \i_qpsi.data[1] ;
 wire \i_qpsi.data[2] ;
 wire \i_qpsi.data[3] ;
 wire \i_qpsi.data[4] ;
 wire \i_qpsi.data[5] ;
 wire \i_qpsi.data[6] ;
 wire \i_qpsi.data[7] ;
 wire \i_qpsi.fsm_state[0] ;
 wire \i_qpsi.fsm_state[1] ;
 wire \i_qpsi.fsm_state[2] ;
 wire \i_qpsi.spi_clk ;
 wire \i_qpsi.spi_clk_n ;
 wire \i_qpsi.spi_data_in[0] ;
 wire \i_qpsi.spi_data_in[1] ;
 wire \i_qpsi.spi_data_oe[0] ;
 wire \i_qpsi.spi_miso_buf[0] ;
 wire \i_qpsi.spi_miso_buf[10] ;
 wire \i_qpsi.spi_miso_buf[11] ;
 wire \i_qpsi.spi_miso_buf[1] ;
 wire \i_qpsi.spi_miso_buf[2] ;
 wire \i_qpsi.spi_miso_buf[3] ;
 wire \i_qpsi.spi_miso_buf[4] ;
 wire \i_qpsi.spi_miso_buf[5] ;
 wire \i_qpsi.spi_miso_buf[6] ;
 wire \i_qpsi.spi_miso_buf[7] ;
 wire \i_qpsi.spi_miso_buf[8] ;
 wire \i_qpsi.spi_miso_buf[9] ;
 wire \i_qpsi.spi_select ;
 wire \i_qpsi.valid ;
 wire net15;
 wire net16;
 wire net266;
 wire net267;
 wire vsync_r;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire clknet_5_0__leaf_clk_regs;
 wire clknet_5_1__leaf_clk_regs;
 wire clknet_5_2__leaf_clk_regs;
 wire clknet_5_3__leaf_clk_regs;
 wire clknet_5_4__leaf_clk_regs;
 wire clknet_5_5__leaf_clk_regs;
 wire clknet_5_6__leaf_clk_regs;
 wire clknet_5_7__leaf_clk_regs;
 wire clknet_5_8__leaf_clk_regs;
 wire clknet_5_9__leaf_clk_regs;
 wire clknet_5_10__leaf_clk_regs;
 wire clknet_5_11__leaf_clk_regs;
 wire clknet_5_12__leaf_clk_regs;
 wire clknet_5_13__leaf_clk_regs;
 wire clknet_5_14__leaf_clk_regs;
 wire clknet_5_15__leaf_clk_regs;
 wire clknet_5_16__leaf_clk_regs;
 wire clknet_5_17__leaf_clk_regs;
 wire clknet_5_18__leaf_clk_regs;
 wire clknet_5_19__leaf_clk_regs;
 wire clknet_5_20__leaf_clk_regs;
 wire clknet_5_21__leaf_clk_regs;
 wire clknet_5_22__leaf_clk_regs;
 wire clknet_5_23__leaf_clk_regs;
 wire clknet_5_24__leaf_clk_regs;
 wire clknet_5_25__leaf_clk_regs;
 wire clknet_5_26__leaf_clk_regs;
 wire clknet_5_27__leaf_clk_regs;
 wire clknet_5_28__leaf_clk_regs;
 wire clknet_5_29__leaf_clk_regs;
 wire clknet_5_30__leaf_clk_regs;
 wire clknet_5_31__leaf_clk_regs;
 wire delaynet_0_clk;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;

 sg13g2_inv_1 _0791_ (.Y(_0173_),
    .A(net556));
 sg13g2_inv_1 _0792_ (.Y(_0174_),
    .A(net360));
 sg13g2_inv_1 _0793_ (.Y(_0175_),
    .A(net376));
 sg13g2_inv_1 _0794_ (.Y(_0176_),
    .A(net461));
 sg13g2_inv_1 _0795_ (.Y(_0177_),
    .A(net397));
 sg13g2_inv_1 _0796_ (.Y(_0178_),
    .A(net472));
 sg13g2_inv_1 _0797_ (.Y(_0179_),
    .A(net380));
 sg13g2_inv_2 _0798_ (.Y(_0180_),
    .A(net337));
 sg13g2_inv_2 _0799_ (.Y(_0181_),
    .A(net410));
 sg13g2_inv_2 _0800_ (.Y(_0182_),
    .A(net7));
 sg13g2_inv_1 _0801_ (.Y(_0183_),
    .A(net402));
 sg13g2_inv_1 _0802_ (.Y(_0184_),
    .A(\i_display.cfg[4] ));
 sg13g2_inv_1 _0803_ (.Y(_0185_),
    .A(net348));
 sg13g2_inv_1 _0804_ (.Y(_0186_),
    .A(net354));
 sg13g2_buf_8 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_nor2_1 _0806_ (.A(net508),
    .B(net556),
    .Y(_0187_));
 sg13g2_nand2b_2 _0807_ (.Y(_0188_),
    .B(_0187_),
    .A_N(net474));
 sg13g2_inv_2 _0808_ (.Y(\i_qpsi.spi_select ),
    .A(_0188_));
 sg13g2_nand2_1 _0809_ (.Y(_0189_),
    .A(net474),
    .B(_0187_));
 sg13g2_inv_1 _0810_ (.Y(_0190_),
    .A(net140));
 sg13g2_nor3_2 _0811_ (.A(net443),
    .B(\i_qpsi.bits_remaining[1] ),
    .C(net545),
    .Y(_0191_));
 sg13g2_or3_1 _0812_ (.A(net443),
    .B(net557),
    .C(net545),
    .X(_0192_));
 sg13g2_nor2_1 _0813_ (.A(net140),
    .B(_0192_),
    .Y(_0009_));
 sg13g2_and2_1 _0814_ (.A(net1),
    .B(net4),
    .X(_0193_));
 sg13g2_nand2_1 _0815_ (.Y(_0194_),
    .A(net172),
    .B(net4));
 sg13g2_nor3_1 _0816_ (.A(\i_display.h_count[1] ),
    .B(\i_display.h_count[0] ),
    .C(\i_display.h_count[2] ),
    .Y(_0195_));
 sg13g2_nand2b_2 _0817_ (.Y(_0196_),
    .B(_0195_),
    .A_N(net394));
 sg13g2_nor3_1 _0818_ (.A(\i_display.h_count[4] ),
    .B(\i_display.h_count[5] ),
    .C(_0196_),
    .Y(_0197_));
 sg13g2_nor3_1 _0819_ (.A(\i_display.h_count[7] ),
    .B(\i_display.h_count[6] ),
    .C(\i_display.h_count[8] ),
    .Y(_0198_));
 sg13g2_nand2b_1 _0820_ (.Y(_0199_),
    .B(_0197_),
    .A_N(net515));
 sg13g2_and2_1 _0821_ (.A(_0197_),
    .B(_0198_),
    .X(_0200_));
 sg13g2_nor2b_1 _0822_ (.A(\i_display.h_count[9] ),
    .B_N(_0200_),
    .Y(_0201_));
 sg13g2_nand2b_1 _0823_ (.Y(_0202_),
    .B(_0200_),
    .A_N(\i_display.h_count[9] ));
 sg13g2_nor2_2 _0824_ (.A(\i_display.h_count[10] ),
    .B(\i_display.h_count[9] ),
    .Y(_0203_));
 sg13g2_nor2_1 _0825_ (.A(\i_display.h_count[10] ),
    .B(_0202_),
    .Y(_0204_));
 sg13g2_nand2_2 _0826_ (.Y(_0205_),
    .A(_0200_),
    .B(_0203_));
 sg13g2_nor2_1 _0827_ (.A(net159),
    .B(net160),
    .Y(_0206_));
 sg13g2_nor2b_2 _0828_ (.A(net160),
    .B_N(net159),
    .Y(_0207_));
 sg13g2_nor2b_2 _0829_ (.A(net159),
    .B_N(net160),
    .Y(_0208_));
 sg13g2_and2_1 _0830_ (.A(\i_display.h_state[1] ),
    .B(\i_display.h_state[0] ),
    .X(_0209_));
 sg13g2_mux4_1 _0831_ (.S0(\i_display.h_state[0] ),
    .A0(\i_display.cfg[47] ),
    .A1(net325),
    .A2(net461),
    .A3(\i_display.cfg[56] ),
    .S1(\i_display.h_state[1] ),
    .X(_0210_));
 sg13g2_o21ai_1 _0832_ (.B1(_0193_),
    .Y(_0211_),
    .A1(\i_display.h_count[0] ),
    .A2(net129));
 sg13g2_a21oi_1 _0833_ (.A1(net129),
    .A2(_0210_),
    .Y(_0212_),
    .B1(_0211_));
 sg13g2_a21oi_1 _0834_ (.A1(_0176_),
    .A2(net165),
    .Y(_0000_),
    .B1(_0212_));
 sg13g2_a22oi_1 _0835_ (.Y(_0213_),
    .B1(_0208_),
    .B2(net435),
    .A2(net157),
    .A1(net467));
 sg13g2_a22oi_1 _0836_ (.Y(_0214_),
    .B1(_0209_),
    .B2(net495),
    .A2(_0207_),
    .A1(net346));
 sg13g2_nand3_1 _0837_ (.B(_0213_),
    .C(_0214_),
    .A(net130),
    .Y(_0215_));
 sg13g2_xor2_1 _0838_ (.B(\i_display.h_count[0] ),
    .A(net503),
    .X(_0216_));
 sg13g2_nor2_1 _0839_ (.A(net166),
    .B(net504),
    .Y(_0217_));
 sg13g2_a22oi_1 _0840_ (.Y(_0218_),
    .B1(_0215_),
    .B2(_0217_),
    .A2(net166),
    .A1(net346));
 sg13g2_inv_1 _0841_ (.Y(_0001_),
    .A(_0218_));
 sg13g2_o21ai_1 _0842_ (.B1(\i_display.h_count[2] ),
    .Y(_0219_),
    .A1(\i_display.h_count[1] ),
    .A2(\i_display.h_count[0] ));
 sg13g2_nor2b_1 _0843_ (.A(_0195_),
    .B_N(_0219_),
    .Y(_0220_));
 sg13g2_a22oi_1 _0844_ (.Y(_0221_),
    .B1(_0209_),
    .B2(net491),
    .A2(_0208_),
    .A1(\i_display.cfg[40] ));
 sg13g2_a21oi_1 _0845_ (.A1(net397),
    .A2(_0207_),
    .Y(_0222_),
    .B1(net157));
 sg13g2_a221oi_1 _0846_ (.B2(_0222_),
    .C1(_0205_),
    .B1(net492),
    .A1(_0178_),
    .Y(_0223_),
    .A2(net157));
 sg13g2_o21ai_1 _0847_ (.B1(net168),
    .Y(_0224_),
    .A1(net130),
    .A2(_0220_));
 sg13g2_nor2_1 _0848_ (.A(net493),
    .B(_0224_),
    .Y(_0225_));
 sg13g2_a21oi_1 _0849_ (.A1(_0177_),
    .A2(net167),
    .Y(_0002_),
    .B1(net494));
 sg13g2_nor2_1 _0850_ (.A(net343),
    .B(net168),
    .Y(_0226_));
 sg13g2_mux4_1 _0851_ (.S0(net160),
    .A0(\i_display.cfg[50] ),
    .A1(\i_display.cfg[41] ),
    .A2(\i_display.cfg[32] ),
    .A3(\i_display.cfg[59] ),
    .S1(net159),
    .X(_0227_));
 sg13g2_nand2b_1 _0852_ (.Y(_0228_),
    .B(net394),
    .A_N(_0195_));
 sg13g2_a21oi_1 _0853_ (.A1(_0196_),
    .A2(_0228_),
    .Y(_0229_),
    .B1(net129));
 sg13g2_a21oi_1 _0854_ (.A1(net129),
    .A2(_0227_),
    .Y(_0230_),
    .B1(net395));
 sg13g2_a21oi_1 _0855_ (.A1(net169),
    .A2(net396),
    .Y(_0003_),
    .B1(_0226_));
 sg13g2_nand2_1 _0856_ (.Y(_0231_),
    .A(net356),
    .B(net167));
 sg13g2_xor2_1 _0857_ (.B(_0196_),
    .A(\i_display.h_count[4] ),
    .X(_0232_));
 sg13g2_mux4_1 _0858_ (.S0(net160),
    .A0(\i_display.cfg[51] ),
    .A1(\i_display.cfg[42] ),
    .A2(\i_display.cfg[33] ),
    .A3(\i_display.cfg[60] ),
    .S1(net159),
    .X(_0233_));
 sg13g2_o21ai_1 _0859_ (.B1(net169),
    .Y(_0234_),
    .A1(_0205_),
    .A2(_0233_));
 sg13g2_o21ai_1 _0860_ (.B1(_0231_),
    .Y(_0004_),
    .A1(_0232_),
    .A2(_0234_));
 sg13g2_nor2_1 _0861_ (.A(net389),
    .B(net168),
    .Y(_0235_));
 sg13g2_a22oi_1 _0862_ (.Y(_0236_),
    .B1(_0209_),
    .B2(\i_display.cfg[61] ),
    .A2(_0208_),
    .A1(\i_display.cfg[43] ));
 sg13g2_inv_1 _0863_ (.Y(_0237_),
    .A(_0236_));
 sg13g2_a221oi_1 _0864_ (.B2(net389),
    .C1(_0237_),
    .B1(_0207_),
    .A1(\i_display.cfg[52] ),
    .Y(_0238_),
    .A2(net156));
 sg13g2_o21ai_1 _0865_ (.B1(\i_display.h_count[5] ),
    .Y(_0239_),
    .A1(\i_display.h_count[4] ),
    .A2(_0196_));
 sg13g2_nor2b_1 _0866_ (.A(_0197_),
    .B_N(_0239_),
    .Y(_0240_));
 sg13g2_mux2_1 _0867_ (.A0(_0238_),
    .A1(_0240_),
    .S(_0205_),
    .X(_0241_));
 sg13g2_a21oi_1 _0868_ (.A1(net168),
    .A2(_0241_),
    .Y(_0005_),
    .B1(_0235_));
 sg13g2_a21oi_1 _0869_ (.A1(net499),
    .A2(_0209_),
    .Y(_0242_),
    .B1(net156));
 sg13g2_a22oi_1 _0870_ (.Y(_0243_),
    .B1(_0208_),
    .B2(net448),
    .A2(_0207_),
    .A1(net380));
 sg13g2_a22oi_1 _0871_ (.Y(_0244_),
    .B1(_0242_),
    .B2(_0243_),
    .A2(net156),
    .A1(_0180_));
 sg13g2_nand2b_1 _0872_ (.Y(_0245_),
    .B(net515),
    .A_N(_0197_));
 sg13g2_a21o_1 _0873_ (.A2(_0245_),
    .A1(_0199_),
    .B1(net129),
    .X(_0246_));
 sg13g2_a21oi_1 _0874_ (.A1(net129),
    .A2(_0244_),
    .Y(_0247_),
    .B1(net167));
 sg13g2_a22oi_1 _0875_ (.Y(_0006_),
    .B1(_0246_),
    .B2(_0247_),
    .A2(net167),
    .A1(_0179_));
 sg13g2_nor2_1 _0876_ (.A(net378),
    .B(net168),
    .Y(_0248_));
 sg13g2_xnor2_1 _0877_ (.Y(_0249_),
    .A(net446),
    .B(_0199_));
 sg13g2_a22oi_1 _0878_ (.Y(_0250_),
    .B1(_0208_),
    .B2(\i_display.cfg[45] ),
    .A2(_0207_),
    .A1(net378));
 sg13g2_a22oi_1 _0879_ (.Y(_0251_),
    .B1(_0209_),
    .B2(\i_display.cfg[63] ),
    .A2(net156),
    .A1(net345));
 sg13g2_a21oi_1 _0880_ (.A1(_0250_),
    .A2(_0251_),
    .Y(_0252_),
    .B1(_0205_));
 sg13g2_a21oi_1 _0881_ (.A1(_0205_),
    .A2(_0249_),
    .Y(_0253_),
    .B1(_0252_));
 sg13g2_a21oi_1 _0882_ (.A1(net168),
    .A2(net447),
    .Y(_0007_),
    .B1(_0248_));
 sg13g2_mux4_1 _0883_ (.S0(net160),
    .A0(\i_display.cfg[55] ),
    .A1(\i_display.cfg[46] ),
    .A2(net410),
    .A3(\i_display.cfg[64] ),
    .S1(net159),
    .X(_0254_));
 sg13g2_o21ai_1 _0884_ (.B1(\i_display.h_count[8] ),
    .Y(_0255_),
    .A1(\i_display.h_count[7] ),
    .A2(_0199_));
 sg13g2_nand2b_1 _0885_ (.Y(_0256_),
    .B(_0200_),
    .A_N(_0203_));
 sg13g2_nand3_1 _0886_ (.B(_0255_),
    .C(_0256_),
    .A(net168),
    .Y(_0257_));
 sg13g2_a21oi_1 _0887_ (.A1(net129),
    .A2(_0254_),
    .Y(_0258_),
    .B1(_0257_));
 sg13g2_a21oi_1 _0888_ (.A1(_0181_),
    .A2(net167),
    .Y(_0008_),
    .B1(_0258_));
 sg13g2_mux2_1 _0889_ (.A0(net9),
    .A1(net10),
    .S(net171),
    .X(\i_qpsi.spi_data_in[0] ));
 sg13g2_mux2_1 _0890_ (.A0(net10),
    .A1(net11),
    .S(net171),
    .X(\i_qpsi.spi_data_in[1] ));
 sg13g2_nor2b_1 _0891_ (.A(net474),
    .B_N(\i_qpsi.fsm_state[1] ),
    .Y(_0259_));
 sg13g2_and2_1 _0892_ (.A(_0173_),
    .B(_0259_),
    .X(_0260_));
 sg13g2_nor3_1 _0893_ (.A(\i_qpsi.fsm_state[2] ),
    .B(\i_qpsi.fsm_state[1] ),
    .C(_0173_),
    .Y(_0261_));
 sg13g2_o21ai_1 _0894_ (.B1(\i_qpsi.bits_remaining[2] ),
    .Y(_0262_),
    .A1(\i_qpsi.bits_remaining[1] ),
    .A2(\i_qpsi.bits_remaining[0] ));
 sg13g2_nor2b_1 _0895_ (.A(\i_qpsi.bits_remaining[1] ),
    .B_N(\i_qpsi.bits_remaining[0] ),
    .Y(_0263_));
 sg13g2_o21ai_1 _0896_ (.B1(_0262_),
    .Y(_0264_),
    .A1(\i_qpsi.bits_remaining[2] ),
    .A2(_0263_));
 sg13g2_a22oi_1 _0897_ (.Y(_0265_),
    .B1(_0261_),
    .B2(_0264_),
    .A2(net135),
    .A1(\i_qpsi.addr[20] ));
 sg13g2_mux2_1 _0898_ (.A0(\i_qpsi.spi_clk ),
    .A1(\i_qpsi.spi_clk_n ),
    .S(net5),
    .X(_0266_));
 sg13g2_nand2_1 _0899_ (.Y(_0267_),
    .A(net171),
    .B(_0266_));
 sg13g2_o21ai_1 _0900_ (.B1(_0267_),
    .Y(uio_out[1]),
    .A1(net170),
    .A2(_0265_));
 sg13g2_nand2_1 _0901_ (.Y(_0268_),
    .A(\i_qpsi.addr[21] ),
    .B(net135));
 sg13g2_a21oi_1 _0902_ (.A1(\i_qpsi.addr[21] ),
    .A2(net135),
    .Y(_0269_),
    .B1(net170));
 sg13g2_a21oi_1 _0903_ (.A1(net170),
    .A2(_0265_),
    .Y(uio_out[2]),
    .B1(_0269_));
 sg13g2_nor2_1 _0904_ (.A(net170),
    .B(_0266_),
    .Y(_0270_));
 sg13g2_a21oi_1 _0905_ (.A1(net170),
    .A2(_0268_),
    .Y(uio_out[3]),
    .B1(_0270_));
 sg13g2_o21ai_1 _0906_ (.B1(net172),
    .Y(_0271_),
    .A1(\i_qpsi.spi_data_oe[0] ),
    .A2(net170));
 sg13g2_inv_2 _0907_ (.Y(uio_oe[1]),
    .A(_0271_));
 sg13g2_and3_2 _0908_ (.X(uio_oe[2]),
    .A(\i_qpsi.spi_data_oe[0] ),
    .B(net172),
    .C(net170));
 sg13g2_nor2b_2 _0909_ (.A(net170),
    .B_N(net172),
    .Y(uio_oe[3]));
 sg13g2_and2_1 _0910_ (.A(\i_qpsi.addr[22] ),
    .B(net137),
    .X(uio_out[4]));
 sg13g2_and2_1 _0911_ (.A(\i_qpsi.addr[23] ),
    .B(net137),
    .X(uio_out[5]));
 sg13g2_nor2b_1 _0912_ (.A(net162),
    .B_N(net161),
    .Y(_0272_));
 sg13g2_xor2_1 _0913_ (.B(_0272_),
    .A(net317),
    .X(\i_display.vsync ));
 sg13g2_xor2_1 _0914_ (.B(_0207_),
    .A(net281),
    .X(hsync));
 sg13g2_nor3_1 _0915_ (.A(net532),
    .B(\i_display.v_count[0] ),
    .C(net513),
    .Y(_0273_));
 sg13g2_nor2b_1 _0916_ (.A(\i_display.v_count[3] ),
    .B_N(_0273_),
    .Y(_0274_));
 sg13g2_nor2b_1 _0917_ (.A(net418),
    .B_N(_0274_),
    .Y(_0275_));
 sg13g2_nand2b_1 _0918_ (.Y(_0276_),
    .B(_0275_),
    .A_N(net560));
 sg13g2_nand3_1 _0919_ (.B(net160),
    .C(net130),
    .A(net159),
    .Y(_0277_));
 sg13g2_or2_1 _0920_ (.X(_0278_),
    .B(_0277_),
    .A(_0276_));
 sg13g2_nand2_2 _0921_ (.Y(_0279_),
    .A(net130),
    .B(_0209_));
 sg13g2_nor2_1 _0922_ (.A(net398),
    .B(\i_display.v_count[9] ),
    .Y(_0280_));
 sg13g2_nor3_1 _0923_ (.A(net549),
    .B(net371),
    .C(net473),
    .Y(_0281_));
 sg13g2_nand2_1 _0924_ (.Y(_0282_),
    .A(_0280_),
    .B(_0281_));
 sg13g2_or2_1 _0925_ (.X(_0283_),
    .B(_0282_),
    .A(_0276_));
 sg13g2_and2_1 _0926_ (.A(net161),
    .B(net162),
    .X(_0284_));
 sg13g2_a21oi_1 _0927_ (.A1(net466),
    .A2(_0284_),
    .Y(_0285_),
    .B1(net131));
 sg13g2_nor3_1 _0928_ (.A(net473),
    .B(_0278_),
    .C(_0285_),
    .Y(_0286_));
 sg13g2_a21oi_1 _0929_ (.A1(net473),
    .A2(_0278_),
    .Y(_0287_),
    .B1(_0286_));
 sg13g2_nor2_1 _0930_ (.A(net165),
    .B(_0287_),
    .Y(_0011_));
 sg13g2_o21ai_1 _0931_ (.B1(net371),
    .Y(_0288_),
    .A1(\i_display.v_count[6] ),
    .A2(_0278_));
 sg13g2_a21oi_1 _0932_ (.A1(\i_display.cfg[25] ),
    .A2(_0284_),
    .Y(_0289_),
    .B1(net131));
 sg13g2_nor4_1 _0933_ (.A(net371),
    .B(net473),
    .C(_0276_),
    .D(_0279_),
    .Y(_0290_));
 sg13g2_nand2b_1 _0934_ (.Y(_0291_),
    .B(_0290_),
    .A_N(_0289_));
 sg13g2_a21oi_1 _0935_ (.A1(net372),
    .A2(_0291_),
    .Y(_0012_),
    .B1(net165));
 sg13g2_nor2b_1 _0936_ (.A(_0290_),
    .B_N(net549),
    .Y(_0292_));
 sg13g2_nor2b_1 _0937_ (.A(net549),
    .B_N(_0290_),
    .Y(_0293_));
 sg13g2_nor2_1 _0938_ (.A(_0278_),
    .B(_0282_),
    .Y(_0294_));
 sg13g2_and2_1 _0939_ (.A(_0284_),
    .B(_0294_),
    .X(_0295_));
 sg13g2_nand2b_1 _0940_ (.Y(_0296_),
    .B(_0293_),
    .A_N(net553));
 sg13g2_a221oi_1 _0941_ (.B2(net429),
    .C1(net550),
    .B1(_0295_),
    .A1(net131),
    .Y(_0297_),
    .A2(_0293_));
 sg13g2_nor2_1 _0942_ (.A(net165),
    .B(_0297_),
    .Y(_0013_));
 sg13g2_nand2b_1 _0943_ (.Y(_0298_),
    .B(net553),
    .A_N(_0293_));
 sg13g2_a21oi_1 _0944_ (.A1(net454),
    .A2(_0284_),
    .Y(_0299_),
    .B1(net398));
 sg13g2_o21ai_1 _0945_ (.B1(_0298_),
    .Y(_0300_),
    .A1(_0296_),
    .A2(_0299_));
 sg13g2_and2_1 _0946_ (.A(net169),
    .B(_0300_),
    .X(_0014_));
 sg13g2_a22oi_1 _0947_ (.Y(_0301_),
    .B1(_0296_),
    .B2(net398),
    .A2(_0295_),
    .A1(net384));
 sg13g2_nor2_1 _0948_ (.A(net165),
    .B(net399),
    .Y(_0015_));
 sg13g2_nand2_2 _0949_ (.Y(_0302_),
    .A(net169),
    .B(_0279_));
 sg13g2_nor2_2 _0950_ (.A(net165),
    .B(_0279_),
    .Y(_0303_));
 sg13g2_nor2_2 _0951_ (.A(net161),
    .B(net162),
    .Y(_0304_));
 sg13g2_nor2b_1 _0952_ (.A(net161),
    .B_N(net162),
    .Y(_0305_));
 sg13g2_or2_1 _0953_ (.X(_0306_),
    .B(_0304_),
    .A(\i_display.cfg[18] ));
 sg13g2_mux4_1 _0954_ (.S0(net162),
    .A0(\i_display.cfg[12] ),
    .A1(\i_display.cfg[6] ),
    .A2(\i_display.cfg[0] ),
    .A3(\i_display.cfg[18] ),
    .S1(net161),
    .X(_0307_));
 sg13g2_nor2_1 _0955_ (.A(net132),
    .B(_0307_),
    .Y(_0308_));
 sg13g2_o21ai_1 _0956_ (.B1(_0303_),
    .Y(_0309_),
    .A1(\i_display.v_count[0] ),
    .A2(_0308_));
 sg13g2_o21ai_1 _0957_ (.B1(_0309_),
    .Y(_0310_),
    .A1(\i_display.v_count[0] ),
    .A2(_0302_));
 sg13g2_a21oi_1 _0958_ (.A1(_0183_),
    .A2(net166),
    .Y(_0016_),
    .B1(_0310_));
 sg13g2_nand2b_1 _0959_ (.Y(_0311_),
    .B(net165),
    .A_N(net339));
 sg13g2_o21ai_1 _0960_ (.B1(_0311_),
    .Y(_0312_),
    .A1(net532),
    .A2(_0302_));
 sg13g2_xnor2_1 _0961_ (.Y(_0313_),
    .A(net532),
    .B(\i_display.v_count[0] ));
 sg13g2_mux4_1 _0962_ (.S0(net162),
    .A0(\i_display.cfg[13] ),
    .A1(\i_display.cfg[7] ),
    .A2(\i_display.cfg[1] ),
    .A3(\i_display.cfg[19] ),
    .S1(net161),
    .X(_0314_));
 sg13g2_nor2b_1 _0963_ (.A(net131),
    .B_N(_0314_),
    .Y(_0315_));
 sg13g2_a21oi_1 _0964_ (.A1(net131),
    .A2(_0313_),
    .Y(_0316_),
    .B1(_0315_));
 sg13g2_a21oi_1 _0965_ (.A1(_0303_),
    .A2(_0316_),
    .Y(_0017_),
    .B1(_0312_));
 sg13g2_nand2b_1 _0966_ (.Y(_0317_),
    .B(net165),
    .A_N(net483));
 sg13g2_o21ai_1 _0967_ (.B1(_0317_),
    .Y(_0318_),
    .A1(net513),
    .A2(_0302_));
 sg13g2_o21ai_1 _0968_ (.B1(net513),
    .Y(_0319_),
    .A1(\i_display.v_count[1] ),
    .A2(\i_display.v_count[0] ));
 sg13g2_nand2b_1 _0969_ (.Y(_0320_),
    .B(_0319_),
    .A_N(_0273_));
 sg13g2_mux4_1 _0970_ (.S0(net162),
    .A0(\i_display.cfg[14] ),
    .A1(\i_display.cfg[8] ),
    .A2(\i_display.cfg[2] ),
    .A3(\i_display.cfg[20] ),
    .S1(net161),
    .X(_0321_));
 sg13g2_nor2b_1 _0971_ (.A(net131),
    .B_N(_0321_),
    .Y(_0322_));
 sg13g2_a21oi_1 _0972_ (.A1(net131),
    .A2(_0320_),
    .Y(_0323_),
    .B1(_0322_));
 sg13g2_a21oi_1 _0973_ (.A1(_0303_),
    .A2(_0323_),
    .Y(_0018_),
    .B1(_0318_));
 sg13g2_xor2_1 _0974_ (.B(_0273_),
    .A(net543),
    .X(_0324_));
 sg13g2_mux4_1 _0975_ (.S0(net162),
    .A0(\i_display.cfg[15] ),
    .A1(\i_display.cfg[9] ),
    .A2(\i_display.cfg[3] ),
    .A3(\i_display.cfg[21] ),
    .S1(net528),
    .X(_0325_));
 sg13g2_o21ai_1 _0976_ (.B1(_0324_),
    .Y(_0326_),
    .A1(net132),
    .A2(_0325_));
 sg13g2_nand2b_1 _0977_ (.Y(_0327_),
    .B(net166),
    .A_N(net400));
 sg13g2_o21ai_1 _0978_ (.B1(_0327_),
    .Y(_0328_),
    .A1(net543),
    .A2(_0302_));
 sg13g2_a21oi_1 _0979_ (.A1(_0303_),
    .A2(_0326_),
    .Y(_0019_),
    .B1(_0328_));
 sg13g2_nor2_1 _0980_ (.A(net418),
    .B(_0302_),
    .Y(_0329_));
 sg13g2_xor2_1 _0981_ (.B(_0274_),
    .A(net418),
    .X(_0330_));
 sg13g2_mux4_1 _0982_ (.S0(\i_display.v_state[0] ),
    .A0(\i_display.cfg[16] ),
    .A1(\i_display.cfg[10] ),
    .A2(\i_display.cfg[4] ),
    .A3(\i_display.cfg[22] ),
    .S1(\i_display.v_state[1] ),
    .X(_0331_));
 sg13g2_o21ai_1 _0983_ (.B1(_0330_),
    .Y(_0332_),
    .A1(net132),
    .A2(_0331_));
 sg13g2_a221oi_1 _0984_ (.B2(_0332_),
    .C1(_0329_),
    .B1(_0303_),
    .A1(_0184_),
    .Y(_0020_),
    .A2(net166));
 sg13g2_a22oi_1 _0985_ (.Y(_0333_),
    .B1(_0305_),
    .B2(net425),
    .A2(_0272_),
    .A1(net366));
 sg13g2_a22oi_1 _0986_ (.Y(_0334_),
    .B1(_0304_),
    .B2(net431),
    .A2(_0284_),
    .A1(net428));
 sg13g2_nand2_1 _0987_ (.Y(_0335_),
    .A(_0333_),
    .B(_0334_));
 sg13g2_xor2_1 _0988_ (.B(_0275_),
    .A(net522),
    .X(_0336_));
 sg13g2_o21ai_1 _0989_ (.B1(_0336_),
    .Y(_0337_),
    .A1(net131),
    .A2(_0335_));
 sg13g2_nand2b_1 _0990_ (.Y(_0338_),
    .B(net166),
    .A_N(net366));
 sg13g2_o21ai_1 _0991_ (.B1(_0338_),
    .Y(_0339_),
    .A1(net522),
    .A2(_0302_));
 sg13g2_a21oi_1 _0992_ (.A1(_0303_),
    .A2(_0337_),
    .Y(_0021_),
    .B1(_0339_));
 sg13g2_nand2_2 _0993_ (.Y(_0340_),
    .A(net157),
    .B(_0304_));
 sg13g2_nor2b_1 _0994_ (.A(net163),
    .B_N(net368),
    .Y(_0341_));
 sg13g2_a21oi_1 _0995_ (.A1(net163),
    .A2(net283),
    .Y(_0342_),
    .B1(net369));
 sg13g2_nor2_1 _0996_ (.A(_0340_),
    .B(net370),
    .Y(_0022_));
 sg13g2_nor2b_1 _0997_ (.A(net164),
    .B_N(net422),
    .Y(_0343_));
 sg13g2_a21oi_1 _0998_ (.A1(net164),
    .A2(net313),
    .Y(_0344_),
    .B1(net423));
 sg13g2_nor2_1 _0999_ (.A(_0340_),
    .B(net424),
    .Y(_0023_));
 sg13g2_nor2b_1 _1000_ (.A(net163),
    .B_N(net412),
    .Y(_0345_));
 sg13g2_a21oi_1 _1001_ (.A1(net164),
    .A2(net330),
    .Y(_0346_),
    .B1(net413));
 sg13g2_nor2_1 _1002_ (.A(_0340_),
    .B(net414),
    .Y(_0024_));
 sg13g2_nor2b_1 _1003_ (.A(net163),
    .B_N(net391),
    .Y(_0347_));
 sg13g2_a21oi_1 _1004_ (.A1(net163),
    .A2(net303),
    .Y(_0348_),
    .B1(net392));
 sg13g2_nor2_1 _1005_ (.A(_0340_),
    .B(net393),
    .Y(_0025_));
 sg13g2_nor2b_1 _1006_ (.A(net163),
    .B_N(net404),
    .Y(_0349_));
 sg13g2_a21oi_1 _1007_ (.A1(net163),
    .A2(net376),
    .Y(_0350_),
    .B1(net405));
 sg13g2_nor2_1 _1008_ (.A(_0340_),
    .B(net406),
    .Y(_0026_));
 sg13g2_nor2b_1 _1009_ (.A(net163),
    .B_N(uo_out[0]),
    .Y(_0351_));
 sg13g2_a21oi_1 _1010_ (.A1(net360),
    .A2(net164),
    .Y(_0352_),
    .B1(_0351_));
 sg13g2_nor2_1 _1011_ (.A(_0340_),
    .B(net361),
    .Y(_0027_));
 sg13g2_xnor2_1 _1012_ (.Y(_0353_),
    .A(\i_display.h_count[1] ),
    .B(\i_display.cfg[70] ));
 sg13g2_xnor2_1 _1013_ (.Y(_0354_),
    .A(\i_display.cfg[74] ),
    .B(\i_display.h_count[5] ));
 sg13g2_xnor2_1 _1014_ (.Y(_0355_),
    .A(\i_display.cfg[69] ),
    .B(\i_display.h_count[0] ));
 sg13g2_xor2_1 _1015_ (.B(\i_display.h_count[3] ),
    .A(\i_display.cfg[72] ),
    .X(_0356_));
 sg13g2_nor2b_1 _1016_ (.A(\i_display.h_count[2] ),
    .B_N(\i_display.cfg[71] ),
    .Y(_0357_));
 sg13g2_o21ai_1 _1017_ (.B1(_0198_),
    .Y(_0358_),
    .A1(_0284_),
    .A2(_0304_));
 sg13g2_nand2b_1 _1018_ (.Y(_0359_),
    .B(\i_display.cfg[73] ),
    .A_N(\i_display.h_count[4] ));
 sg13g2_nand2b_1 _1019_ (.Y(_0360_),
    .B(\i_display.h_count[4] ),
    .A_N(\i_display.cfg[73] ));
 sg13g2_nand2b_1 _1020_ (.Y(_0361_),
    .B(\i_display.h_count[2] ),
    .A_N(\i_display.cfg[71] ));
 sg13g2_nand4_1 _1021_ (.B(_0359_),
    .C(_0360_),
    .A(_0203_),
    .Y(_0362_),
    .D(_0361_));
 sg13g2_nor4_1 _1022_ (.A(_0356_),
    .B(_0357_),
    .C(_0358_),
    .D(_0362_),
    .Y(_0363_));
 sg13g2_nand4_1 _1023_ (.B(_0354_),
    .C(_0355_),
    .A(_0353_),
    .Y(_0364_),
    .D(_0363_));
 sg13g2_a21o_2 _1024_ (.A2(net132),
    .A1(net161),
    .B1(_0364_),
    .X(_0365_));
 sg13g2_nor2_1 _1025_ (.A(_0188_),
    .B(_0365_),
    .Y(_0366_));
 sg13g2_nor2b_1 _1026_ (.A(net133),
    .B_N(\i_qpsi.addr[4] ),
    .Y(_0367_));
 sg13g2_a21oi_1 _1027_ (.A1(net329),
    .A2(net133),
    .Y(_0368_),
    .B1(_0367_));
 sg13g2_nand2_1 _1028_ (.Y(_0369_),
    .A(net364),
    .B(net124));
 sg13g2_o21ai_1 _1029_ (.B1(_0369_),
    .Y(_0028_),
    .A1(net124),
    .A2(_0368_));
 sg13g2_nor2_2 _1030_ (.A(net133),
    .B(net124),
    .Y(_0370_));
 sg13g2_nand2_1 _1031_ (.Y(_0371_),
    .A(net291),
    .B(_0370_));
 sg13g2_a22oi_1 _1032_ (.Y(_0372_),
    .B1(net124),
    .B2(\addr_in[5] ),
    .A2(net133),
    .A1(\i_qpsi.addr[1] ));
 sg13g2_nand2_1 _1033_ (.Y(_0029_),
    .A(_0371_),
    .B(_0372_));
 sg13g2_nand2_1 _1034_ (.Y(_0373_),
    .A(net289),
    .B(net119));
 sg13g2_a22oi_1 _1035_ (.Y(_0374_),
    .B1(net125),
    .B2(\addr_in[6] ),
    .A2(net134),
    .A1(\i_qpsi.addr[2] ));
 sg13g2_nand2_1 _1036_ (.Y(_0030_),
    .A(_0373_),
    .B(_0374_));
 sg13g2_nand2_1 _1037_ (.Y(_0375_),
    .A(net307),
    .B(net119));
 sg13g2_a22oi_1 _1038_ (.Y(_0376_),
    .B1(net125),
    .B2(\addr_in[7] ),
    .A2(net134),
    .A1(\i_qpsi.addr[3] ));
 sg13g2_nand2_1 _1039_ (.Y(_0031_),
    .A(_0375_),
    .B(_0376_));
 sg13g2_nor2b_1 _1040_ (.A(net137),
    .B_N(\i_qpsi.addr[8] ),
    .Y(_0377_));
 sg13g2_a21oi_1 _1041_ (.A1(\i_qpsi.addr[4] ),
    .A2(net133),
    .Y(_0378_),
    .B1(_0377_));
 sg13g2_nand2_1 _1042_ (.Y(_0379_),
    .A(net362),
    .B(net124));
 sg13g2_o21ai_1 _1043_ (.B1(_0379_),
    .Y(_0032_),
    .A1(net128),
    .A2(_0378_));
 sg13g2_nand2_1 _1044_ (.Y(_0380_),
    .A(net299),
    .B(_0370_));
 sg13g2_a22oi_1 _1045_ (.Y(_0381_),
    .B1(net124),
    .B2(\addr_in[9] ),
    .A2(net133),
    .A1(net291));
 sg13g2_nand2_1 _1046_ (.Y(_0033_),
    .A(_0380_),
    .B(_0381_));
 sg13g2_nand2_1 _1047_ (.Y(_0382_),
    .A(net295),
    .B(net119));
 sg13g2_a22oi_1 _1048_ (.Y(_0383_),
    .B1(net125),
    .B2(\addr_in[10] ),
    .A2(net134),
    .A1(net289));
 sg13g2_nand2_1 _1049_ (.Y(_0034_),
    .A(_0382_),
    .B(_0383_));
 sg13g2_nand2_1 _1050_ (.Y(_0384_),
    .A(net311),
    .B(net119));
 sg13g2_a22oi_1 _1051_ (.Y(_0385_),
    .B1(net125),
    .B2(\addr_in[11] ),
    .A2(net134),
    .A1(net307));
 sg13g2_nand2_1 _1052_ (.Y(_0035_),
    .A(_0384_),
    .B(_0385_));
 sg13g2_nand2_1 _1053_ (.Y(_0386_),
    .A(net315),
    .B(net120));
 sg13g2_a22oi_1 _1054_ (.Y(_0387_),
    .B1(net128),
    .B2(\addr_in[12] ),
    .A2(net133),
    .A1(\i_qpsi.addr[8] ));
 sg13g2_nand2_1 _1055_ (.Y(_0036_),
    .A(_0386_),
    .B(_0387_));
 sg13g2_nand2_1 _1056_ (.Y(_0388_),
    .A(net285),
    .B(net120));
 sg13g2_a22oi_1 _1057_ (.Y(_0389_),
    .B1(net125),
    .B2(\addr_in[13] ),
    .A2(net134),
    .A1(\i_qpsi.addr[9] ));
 sg13g2_nand2_1 _1058_ (.Y(_0037_),
    .A(_0388_),
    .B(_0389_));
 sg13g2_nand2_1 _1059_ (.Y(_0390_),
    .A(net321),
    .B(net119));
 sg13g2_a22oi_1 _1060_ (.Y(_0391_),
    .B1(net125),
    .B2(\addr_in[14] ),
    .A2(net134),
    .A1(net295));
 sg13g2_nand2_1 _1061_ (.Y(_0038_),
    .A(_0390_),
    .B(_0391_));
 sg13g2_nand2_1 _1062_ (.Y(_0392_),
    .A(net305),
    .B(net119));
 sg13g2_a22oi_1 _1063_ (.Y(_0393_),
    .B1(net126),
    .B2(\addr_in[15] ),
    .A2(net134),
    .A1(\i_qpsi.addr[11] ));
 sg13g2_nand2_1 _1064_ (.Y(_0039_),
    .A(_0392_),
    .B(_0393_));
 sg13g2_nand2_1 _1065_ (.Y(_0394_),
    .A(net297),
    .B(net120));
 sg13g2_a22oi_1 _1066_ (.Y(_0395_),
    .B1(net127),
    .B2(\addr_in[16] ),
    .A2(net133),
    .A1(\i_qpsi.addr[12] ));
 sg13g2_nand2_1 _1067_ (.Y(_0040_),
    .A(_0394_),
    .B(_0395_));
 sg13g2_nand2_1 _1068_ (.Y(_0396_),
    .A(net279),
    .B(net120));
 sg13g2_a22oi_1 _1069_ (.Y(_0397_),
    .B1(net126),
    .B2(\addr_in[17] ),
    .A2(net136),
    .A1(\i_qpsi.addr[13] ));
 sg13g2_nand2_1 _1070_ (.Y(_0041_),
    .A(_0396_),
    .B(_0397_));
 sg13g2_nand2_1 _1071_ (.Y(_0398_),
    .A(net287),
    .B(net120));
 sg13g2_a22oi_1 _1072_ (.Y(_0399_),
    .B1(net126),
    .B2(\addr_in[18] ),
    .A2(net136),
    .A1(\i_qpsi.addr[14] ));
 sg13g2_nand2_1 _1073_ (.Y(_0042_),
    .A(_0398_),
    .B(_0399_));
 sg13g2_nand2_1 _1074_ (.Y(_0400_),
    .A(net309),
    .B(net120));
 sg13g2_a22oi_1 _1075_ (.Y(_0401_),
    .B1(net126),
    .B2(\addr_in[19] ),
    .A2(net136),
    .A1(net305));
 sg13g2_nand2_1 _1076_ (.Y(_0043_),
    .A(_0400_),
    .B(_0401_));
 sg13g2_nor2b_1 _1077_ (.A(net135),
    .B_N(\i_qpsi.addr[20] ),
    .Y(_0402_));
 sg13g2_a21oi_1 _1078_ (.A1(net297),
    .A2(net135),
    .Y(_0403_),
    .B1(_0402_));
 sg13g2_nand2_1 _1079_ (.Y(_0404_),
    .A(net374),
    .B(net127));
 sg13g2_o21ai_1 _1080_ (.B1(_0404_),
    .Y(_0044_),
    .A1(net127),
    .A2(_0403_));
 sg13g2_nor2b_1 _1081_ (.A(net137),
    .B_N(net353),
    .Y(_0405_));
 sg13g2_a21oi_1 _1082_ (.A1(net279),
    .A2(net135),
    .Y(_0406_),
    .B1(_0405_));
 sg13g2_nand2_1 _1083_ (.Y(_0407_),
    .A(net350),
    .B(net126));
 sg13g2_o21ai_1 _1084_ (.B1(_0407_),
    .Y(_0045_),
    .A1(net126),
    .A2(_0406_));
 sg13g2_nor2b_1 _1085_ (.A(net136),
    .B_N(\i_qpsi.addr[22] ),
    .Y(_0408_));
 sg13g2_a21oi_1 _1086_ (.A1(net287),
    .A2(net136),
    .Y(_0409_),
    .B1(_0408_));
 sg13g2_nand2_1 _1087_ (.Y(_0410_),
    .A(net323),
    .B(net126));
 sg13g2_o21ai_1 _1088_ (.B1(_0410_),
    .Y(_0046_),
    .A1(net126),
    .A2(_0409_));
 sg13g2_nor2b_1 _1089_ (.A(net136),
    .B_N(\i_qpsi.addr[23] ),
    .Y(_0411_));
 sg13g2_a21oi_1 _1090_ (.A1(net309),
    .A2(net136),
    .Y(_0412_),
    .B1(_0411_));
 sg13g2_nand2_1 _1091_ (.Y(_0413_),
    .A(net319),
    .B(net127));
 sg13g2_o21ai_1 _1092_ (.B1(_0413_),
    .Y(_0047_),
    .A1(net127),
    .A2(_0412_));
 sg13g2_mux2_1 _1093_ (.A0(\i_display.cfg[57] ),
    .A1(\i_display.h_count[1] ),
    .S(net158),
    .X(_0414_));
 sg13g2_mux2_1 _1094_ (.A0(\i_display.cfg[58] ),
    .A1(\i_display.h_count[2] ),
    .S(net158),
    .X(_0415_));
 sg13g2_mux2_1 _1095_ (.A0(\i_display.cfg[64] ),
    .A1(\i_display.h_count[8] ),
    .S(net156),
    .X(_0416_));
 sg13g2_mux2_1 _1096_ (.A0(\i_display.cfg[63] ),
    .A1(\i_display.h_count[7] ),
    .S(net157),
    .X(_0417_));
 sg13g2_mux2_1 _1097_ (.A0(\i_display.cfg[62] ),
    .A1(\i_display.h_count[6] ),
    .S(net157),
    .X(_0418_));
 sg13g2_mux2_1 _1098_ (.A0(\i_display.cfg[61] ),
    .A1(\i_display.h_count[5] ),
    .S(net157),
    .X(_0419_));
 sg13g2_mux2_1 _1099_ (.A0(\i_display.cfg[60] ),
    .A1(\i_display.h_count[4] ),
    .S(net156),
    .X(_0420_));
 sg13g2_mux2_1 _1100_ (.A0(\i_display.cfg[65] ),
    .A1(\i_display.h_count[9] ),
    .S(net156),
    .X(_0421_));
 sg13g2_mux2_1 _1101_ (.A0(\i_display.cfg[56] ),
    .A1(\i_display.h_count[0] ),
    .S(net158),
    .X(_0422_));
 sg13g2_mux2_1 _1102_ (.A0(\i_display.cfg[59] ),
    .A1(\i_display.h_count[3] ),
    .S(net158),
    .X(_0423_));
 sg13g2_mux2_1 _1103_ (.A0(\i_display.cfg[66] ),
    .A1(\i_display.h_count[10] ),
    .S(net156),
    .X(_0424_));
 sg13g2_nor3_1 _1104_ (.A(_0419_),
    .B(_0421_),
    .C(_0423_),
    .Y(_0425_));
 sg13g2_nor4_1 _1105_ (.A(_0415_),
    .B(_0417_),
    .C(_0422_),
    .D(_0424_),
    .Y(_0426_));
 sg13g2_nor4_1 _1106_ (.A(_0414_),
    .B(_0416_),
    .C(_0418_),
    .D(_0420_),
    .Y(_0427_));
 sg13g2_nand3_1 _1107_ (.B(_0426_),
    .C(_0427_),
    .A(_0425_),
    .Y(_0428_));
 sg13g2_nand2_2 _1108_ (.Y(_0429_),
    .A(net172),
    .B(_0428_));
 sg13g2_xor2_1 _1109_ (.B(\i_qpsi.spi_select ),
    .A(net518),
    .X(_0430_));
 sg13g2_nor2_1 _1110_ (.A(_0429_),
    .B(net519),
    .Y(_0048_));
 sg13g2_nor3_1 _1111_ (.A(_0173_),
    .B(\i_qpsi.spi_clk ),
    .C(_0191_),
    .Y(_0431_));
 sg13g2_nor2_1 _1112_ (.A(_0187_),
    .B(_0192_),
    .Y(_0432_));
 sg13g2_a221oi_1 _1113_ (.B2(net474),
    .C1(_0431_),
    .B1(_0432_),
    .A1(\i_qpsi.spi_select ),
    .Y(_0433_),
    .A2(_0365_));
 sg13g2_nor2_1 _1114_ (.A(net545),
    .B(_0433_),
    .Y(_0434_));
 sg13g2_or2_1 _1115_ (.X(_0435_),
    .B(_0261_),
    .A(net135));
 sg13g2_and2_1 _1116_ (.A(\i_qpsi.fsm_state[0] ),
    .B(_0259_),
    .X(_0436_));
 sg13g2_a21o_1 _1117_ (.A2(_0436_),
    .A1(net6),
    .B1(_0435_),
    .X(_0437_));
 sg13g2_a22oi_1 _1118_ (.Y(_0438_),
    .B1(_0191_),
    .B2(_0437_),
    .A2(_0188_),
    .A1(net545));
 sg13g2_nor2b_1 _1119_ (.A(_0438_),
    .B_N(_0433_),
    .Y(_0439_));
 sg13g2_nor3_1 _1120_ (.A(_0429_),
    .B(_0434_),
    .C(_0439_),
    .Y(_0049_));
 sg13g2_and2_1 _1121_ (.A(net6),
    .B(net7),
    .X(_0440_));
 sg13g2_xor2_1 _1122_ (.B(net7),
    .A(net6),
    .X(_0441_));
 sg13g2_a21oi_1 _1123_ (.A1(_0436_),
    .A2(_0441_),
    .Y(_0442_),
    .B1(_0435_));
 sg13g2_nor2_1 _1124_ (.A(\i_qpsi.spi_select ),
    .B(_0192_),
    .Y(_0443_));
 sg13g2_xnor2_1 _1125_ (.Y(_0444_),
    .A(\i_qpsi.bits_remaining[1] ),
    .B(\i_qpsi.bits_remaining[0] ));
 sg13g2_a21oi_1 _1126_ (.A1(_0192_),
    .A2(_0444_),
    .Y(_0445_),
    .B1(\i_qpsi.spi_select ));
 sg13g2_o21ai_1 _1127_ (.B1(_0445_),
    .Y(_0446_),
    .A1(_0192_),
    .A2(_0442_));
 sg13g2_mux2_1 _1128_ (.A0(net557),
    .A1(_0446_),
    .S(_0433_),
    .X(_0447_));
 sg13g2_nor2b_1 _1129_ (.A(_0429_),
    .B_N(_0447_),
    .Y(_0050_));
 sg13g2_nor2_1 _1130_ (.A(net443),
    .B(_0433_),
    .Y(_0448_));
 sg13g2_a21oi_1 _1131_ (.A1(_0436_),
    .A2(_0440_),
    .Y(_0449_),
    .B1(_0435_));
 sg13g2_o21ai_1 _1132_ (.B1(_0262_),
    .Y(_0450_),
    .A1(_0192_),
    .A2(_0449_));
 sg13g2_nor2_1 _1133_ (.A(\i_qpsi.spi_select ),
    .B(_0450_),
    .Y(_0451_));
 sg13g2_a21oi_1 _1134_ (.A1(_0433_),
    .A2(_0451_),
    .Y(_0452_),
    .B1(_0429_));
 sg13g2_nor2b_1 _1135_ (.A(net444),
    .B_N(_0452_),
    .Y(_0051_));
 sg13g2_nor2_1 _1136_ (.A(_0173_),
    .B(_0192_),
    .Y(_0453_));
 sg13g2_nor3_1 _1137_ (.A(net556),
    .B(net127),
    .C(_0443_),
    .Y(_0454_));
 sg13g2_nor4_1 _1138_ (.A(_0190_),
    .B(_0429_),
    .C(_0453_),
    .D(_0454_),
    .Y(_0052_));
 sg13g2_nand2_1 _1139_ (.Y(_0455_),
    .A(\i_qpsi.fsm_state[1] ),
    .B(_0453_));
 sg13g2_xnor2_1 _1140_ (.Y(_0456_),
    .A(net508),
    .B(_0453_));
 sg13g2_nor2_1 _1141_ (.A(_0429_),
    .B(net509),
    .Y(_0053_));
 sg13g2_a22oi_1 _1142_ (.Y(_0457_),
    .B1(_0455_),
    .B2(net474),
    .A2(_0436_),
    .A1(_0191_));
 sg13g2_nor2_1 _1143_ (.A(_0429_),
    .B(net475),
    .Y(_0054_));
 sg13g2_a21oi_1 _1144_ (.A1(_0182_),
    .A2(net271),
    .Y(_0458_),
    .B1(net138));
 sg13g2_nor2_2 _1145_ (.A(net6),
    .B(_0182_),
    .Y(_0459_));
 sg13g2_a22oi_1 _1146_ (.Y(_0460_),
    .B1(_0459_),
    .B2(net270),
    .A2(_0440_),
    .A1(\i_qpsi.spi_miso_buf[8] ));
 sg13g2_a22oi_1 _1147_ (.Y(_0055_),
    .B1(_0458_),
    .B2(_0460_),
    .A2(net138),
    .A1(_0185_));
 sg13g2_a21oi_1 _1148_ (.A1(_0182_),
    .A2(net275),
    .Y(_0461_),
    .B1(net140));
 sg13g2_a22oi_1 _1149_ (.Y(_0462_),
    .B1(_0459_),
    .B2(net276),
    .A2(_0440_),
    .A1(\i_qpsi.spi_miso_buf[9] ));
 sg13g2_a22oi_1 _1150_ (.Y(_0056_),
    .B1(_0461_),
    .B2(_0462_),
    .A2(net138),
    .A1(_0175_));
 sg13g2_a21oi_1 _1151_ (.A1(_0182_),
    .A2(net272),
    .Y(_0463_),
    .B1(net138));
 sg13g2_a22oi_1 _1152_ (.Y(_0464_),
    .B1(_0459_),
    .B2(net273),
    .A2(_0440_),
    .A1(net381));
 sg13g2_a22oi_1 _1153_ (.Y(_0057_),
    .B1(_0463_),
    .B2(_0464_),
    .A2(net139),
    .A1(_0174_));
 sg13g2_a21oi_1 _1154_ (.A1(_0182_),
    .A2(net274),
    .Y(_0465_),
    .B1(net138));
 sg13g2_a22oi_1 _1155_ (.Y(_0466_),
    .B1(_0459_),
    .B2(net277),
    .A2(_0440_),
    .A1(\i_qpsi.spi_miso_buf[11] ));
 sg13g2_a22oi_1 _1156_ (.Y(_0058_),
    .B1(_0465_),
    .B2(_0466_),
    .A2(net138),
    .A1(_0186_));
 sg13g2_nand2_1 _1157_ (.Y(_0467_),
    .A(net330),
    .B(net138));
 sg13g2_o21ai_1 _1158_ (.B1(_0467_),
    .Y(_0059_),
    .A1(_0185_),
    .A2(net138));
 sg13g2_nand2_1 _1159_ (.Y(_0468_),
    .A(net303),
    .B(net139));
 sg13g2_o21ai_1 _1160_ (.B1(_0468_),
    .Y(_0060_),
    .A1(_0175_),
    .A2(net139));
 sg13g2_nand2_1 _1161_ (.Y(_0469_),
    .A(net283),
    .B(net139));
 sg13g2_o21ai_1 _1162_ (.B1(_0469_),
    .Y(_0061_),
    .A1(_0174_),
    .A2(net139));
 sg13g2_nand2_1 _1163_ (.Y(_0470_),
    .A(net313),
    .B(net139));
 sg13g2_o21ai_1 _1164_ (.B1(_0470_),
    .Y(_0062_),
    .A1(_0186_),
    .A2(net139));
 sg13g2_nand2b_2 _1165_ (.Y(_0471_),
    .B(net278),
    .A_N(\i_display.cfg_clk_sync[2] ));
 sg13g2_nor2_1 _1166_ (.A(net442),
    .B(net153),
    .Y(_0472_));
 sg13g2_a21oi_1 _1167_ (.A1(_0183_),
    .A2(net151),
    .Y(_0063_),
    .B1(_0472_));
 sg13g2_nand2_1 _1168_ (.Y(_0473_),
    .A(net339),
    .B(net151));
 sg13g2_o21ai_1 _1169_ (.B1(_0473_),
    .Y(_0064_),
    .A1(_0183_),
    .A2(net151));
 sg13g2_mux2_1 _1170_ (.A0(net339),
    .A1(net483),
    .S(net153),
    .X(_0065_));
 sg13g2_mux2_1 _1171_ (.A0(net483),
    .A1(net400),
    .S(net153),
    .X(_0066_));
 sg13g2_nor2_1 _1172_ (.A(net400),
    .B(net154),
    .Y(_0474_));
 sg13g2_a21oi_1 _1173_ (.A1(_0184_),
    .A2(net154),
    .Y(_0067_),
    .B1(_0474_));
 sg13g2_nand2_1 _1174_ (.Y(_0475_),
    .A(net366),
    .B(net154));
 sg13g2_o21ai_1 _1175_ (.B1(_0475_),
    .Y(_0068_),
    .A1(_0184_),
    .A2(net154));
 sg13g2_mux2_1 _1176_ (.A0(net366),
    .A1(net441),
    .S(net152),
    .X(_0069_));
 sg13g2_mux2_1 _1177_ (.A0(net441),
    .A1(net440),
    .S(net151),
    .X(_0070_));
 sg13g2_mux2_1 _1178_ (.A0(net440),
    .A1(net433),
    .S(net153),
    .X(_0071_));
 sg13g2_mux2_1 _1179_ (.A0(net433),
    .A1(\i_display.cfg[9] ),
    .S(net153),
    .X(_0072_));
 sg13g2_mux2_1 _1180_ (.A0(net501),
    .A1(net458),
    .S(net155),
    .X(_0073_));
 sg13g2_mux2_1 _1181_ (.A0(net458),
    .A1(net425),
    .S(net151),
    .X(_0074_));
 sg13g2_mux2_1 _1182_ (.A0(net425),
    .A1(net408),
    .S(net151),
    .X(_0075_));
 sg13g2_mux2_1 _1183_ (.A0(net408),
    .A1(\i_display.cfg[13] ),
    .S(net151),
    .X(_0076_));
 sg13g2_mux2_1 _1184_ (.A0(net436),
    .A1(net426),
    .S(net153),
    .X(_0077_));
 sg13g2_mux2_1 _1185_ (.A0(net426),
    .A1(\i_display.cfg[15] ),
    .S(net153),
    .X(_0078_));
 sg13g2_mux2_1 _1186_ (.A0(\i_display.cfg[15] ),
    .A1(net469),
    .S(net154),
    .X(_0079_));
 sg13g2_mux2_1 _1187_ (.A0(\i_display.cfg[16] ),
    .A1(net431),
    .S(net152),
    .X(_0080_));
 sg13g2_mux2_1 _1188_ (.A0(net431),
    .A1(net490),
    .S(net152),
    .X(_0081_));
 sg13g2_mux2_1 _1189_ (.A0(\i_display.cfg[18] ),
    .A1(net452),
    .S(net151),
    .X(_0082_));
 sg13g2_mux2_1 _1190_ (.A0(net452),
    .A1(net464),
    .S(net153),
    .X(_0083_));
 sg13g2_mux2_1 _1191_ (.A0(net464),
    .A1(\i_display.cfg[21] ),
    .S(net155),
    .X(_0084_));
 sg13g2_mux2_1 _1192_ (.A0(\i_display.cfg[21] ),
    .A1(net416),
    .S(net154),
    .X(_0085_));
 sg13g2_mux2_1 _1193_ (.A0(net416),
    .A1(net428),
    .S(net154),
    .X(_0086_));
 sg13g2_mux2_1 _1194_ (.A0(net428),
    .A1(net466),
    .S(net150),
    .X(_0087_));
 sg13g2_mux2_1 _1195_ (.A0(\i_display.cfg[24] ),
    .A1(net455),
    .S(net150),
    .X(_0088_));
 sg13g2_mux2_1 _1196_ (.A0(net455),
    .A1(net429),
    .S(net150),
    .X(_0089_));
 sg13g2_mux2_1 _1197_ (.A0(net429),
    .A1(\i_display.cfg[27] ),
    .S(net150),
    .X(_0090_));
 sg13g2_mux2_1 _1198_ (.A0(net454),
    .A1(net384),
    .S(net150),
    .X(_0091_));
 sg13g2_nor2_1 _1199_ (.A(net384),
    .B(net150),
    .Y(_0476_));
 sg13g2_a21oi_1 _1200_ (.A1(_0176_),
    .A2(net150),
    .Y(_0092_),
    .B1(_0476_));
 sg13g2_nand2_1 _1201_ (.Y(_0477_),
    .A(net346),
    .B(net148));
 sg13g2_o21ai_1 _1202_ (.B1(_0477_),
    .Y(_0093_),
    .A1(_0176_),
    .A2(net149));
 sg13g2_nor2_1 _1203_ (.A(net346),
    .B(net148),
    .Y(_0478_));
 sg13g2_a21oi_1 _1204_ (.A1(_0177_),
    .A2(net148),
    .Y(_0094_),
    .B1(_0478_));
 sg13g2_nand2_1 _1205_ (.Y(_0479_),
    .A(net343),
    .B(net145));
 sg13g2_o21ai_1 _1206_ (.B1(_0479_),
    .Y(_0095_),
    .A1(_0177_),
    .A2(net145));
 sg13g2_mux2_1 _1207_ (.A0(net343),
    .A1(net356),
    .S(net145),
    .X(_0096_));
 sg13g2_mux2_1 _1208_ (.A0(net356),
    .A1(net389),
    .S(net141),
    .X(_0097_));
 sg13g2_nor2_1 _1209_ (.A(net389),
    .B(net141),
    .Y(_0480_));
 sg13g2_a21oi_1 _1210_ (.A1(_0179_),
    .A2(net142),
    .Y(_0098_),
    .B1(_0480_));
 sg13g2_nand2_1 _1211_ (.Y(_0481_),
    .A(net378),
    .B(net142));
 sg13g2_o21ai_1 _1212_ (.B1(_0481_),
    .Y(_0099_),
    .A1(_0179_),
    .A2(net142));
 sg13g2_nor2_1 _1213_ (.A(net378),
    .B(net143),
    .Y(_0482_));
 sg13g2_a21oi_1 _1214_ (.A1(_0181_),
    .A2(net143),
    .Y(_0100_),
    .B1(_0482_));
 sg13g2_nand2_1 _1215_ (.Y(_0483_),
    .A(net325),
    .B(net148));
 sg13g2_o21ai_1 _1216_ (.B1(_0483_),
    .Y(_0101_),
    .A1(_0181_),
    .A2(net148));
 sg13g2_mux2_1 _1217_ (.A0(net325),
    .A1(net435),
    .S(net148),
    .X(_0102_));
 sg13g2_mux2_1 _1218_ (.A0(net435),
    .A1(net498),
    .S(net149),
    .X(_0103_));
 sg13g2_mux2_1 _1219_ (.A0(\i_display.cfg[40] ),
    .A1(net496),
    .S(net145),
    .X(_0104_));
 sg13g2_mux2_1 _1220_ (.A0(\i_display.cfg[41] ),
    .A1(net481),
    .S(net145),
    .X(_0105_));
 sg13g2_mux2_1 _1221_ (.A0(net481),
    .A1(net489),
    .S(net141),
    .X(_0106_));
 sg13g2_mux2_1 _1222_ (.A0(\i_display.cfg[43] ),
    .A1(net448),
    .S(net141),
    .X(_0107_));
 sg13g2_mux2_1 _1223_ (.A0(net448),
    .A1(net463),
    .S(net141),
    .X(_0108_));
 sg13g2_mux2_1 _1224_ (.A0(net463),
    .A1(net471),
    .S(net143),
    .X(_0109_));
 sg13g2_mux2_1 _1225_ (.A0(net471),
    .A1(net480),
    .S(net146),
    .X(_0110_));
 sg13g2_mux2_1 _1226_ (.A0(\i_display.cfg[47] ),
    .A1(net467),
    .S(net148),
    .X(_0111_));
 sg13g2_mux2_1 _1227_ (.A0(net467),
    .A1(net472),
    .S(net148),
    .X(_0112_));
 sg13g2_mux2_1 _1228_ (.A0(\i_display.cfg[49] ),
    .A1(net459),
    .S(net146),
    .X(_0113_));
 sg13g2_mux2_1 _1229_ (.A0(net459),
    .A1(net438),
    .S(net143),
    .X(_0114_));
 sg13g2_mux2_1 _1230_ (.A0(net438),
    .A1(\i_display.cfg[52] ),
    .S(net141),
    .X(_0115_));
 sg13g2_nor2_1 _1231_ (.A(\i_display.cfg[52] ),
    .B(net141),
    .Y(_0484_));
 sg13g2_a21oi_1 _1232_ (.A1(_0180_),
    .A2(net141),
    .Y(_0116_),
    .B1(_0484_));
 sg13g2_nand2_1 _1233_ (.Y(_0485_),
    .A(net345),
    .B(net142));
 sg13g2_o21ai_1 _1234_ (.B1(_0485_),
    .Y(_0117_),
    .A1(_0180_),
    .A2(net142));
 sg13g2_mux2_1 _1235_ (.A0(net345),
    .A1(net437),
    .S(net142),
    .X(_0118_));
 sg13g2_mux2_1 _1236_ (.A0(net437),
    .A1(net502),
    .S(net145),
    .X(_0119_));
 sg13g2_mux2_1 _1237_ (.A0(net502),
    .A1(net495),
    .S(net149),
    .X(_0120_));
 sg13g2_mux2_1 _1238_ (.A0(net495),
    .A1(net491),
    .S(net146),
    .X(_0121_));
 sg13g2_mux2_1 _1239_ (.A0(net491),
    .A1(net487),
    .S(net145),
    .X(_0122_));
 sg13g2_mux2_1 _1240_ (.A0(net487),
    .A1(\i_display.cfg[60] ),
    .S(net145),
    .X(_0123_));
 sg13g2_mux2_1 _1241_ (.A0(\i_display.cfg[60] ),
    .A1(net520),
    .S(net144),
    .X(_0124_));
 sg13g2_mux2_1 _1242_ (.A0(\i_display.cfg[61] ),
    .A1(net499),
    .S(net144),
    .X(_0125_));
 sg13g2_mux2_1 _1243_ (.A0(\i_display.cfg[62] ),
    .A1(net485),
    .S(net144),
    .X(_0126_));
 sg13g2_mux2_1 _1244_ (.A0(net485),
    .A1(net484),
    .S(net144),
    .X(_0127_));
 sg13g2_mux2_1 _1245_ (.A0(net484),
    .A1(net386),
    .S(net144),
    .X(_0128_));
 sg13g2_mux2_1 _1246_ (.A0(net386),
    .A1(net358),
    .S(net147),
    .X(_0129_));
 sg13g2_mux2_1 _1247_ (.A0(net358),
    .A1(net317),
    .S(net147),
    .X(_0130_));
 sg13g2_mux2_1 _1248_ (.A0(net317),
    .A1(net281),
    .S(net147),
    .X(_0131_));
 sg13g2_mux2_1 _1249_ (.A0(net281),
    .A1(net457),
    .S(net147),
    .X(_0132_));
 sg13g2_mux2_1 _1250_ (.A0(net457),
    .A1(net450),
    .S(net152),
    .X(_0133_));
 sg13g2_mux2_1 _1251_ (.A0(net450),
    .A1(\i_display.cfg[71] ),
    .S(net149),
    .X(_0134_));
 sg13g2_mux2_1 _1252_ (.A0(net507),
    .A1(net478),
    .S(net149),
    .X(_0135_));
 sg13g2_mux2_1 _1253_ (.A0(net478),
    .A1(\i_display.cfg[73] ),
    .S(net146),
    .X(_0136_));
 sg13g2_mux2_1 _1254_ (.A0(\i_display.cfg[73] ),
    .A1(net420),
    .S(net146),
    .X(_0137_));
 sg13g2_nand2_1 _1255_ (.Y(_0486_),
    .A(_0191_),
    .B(net135));
 sg13g2_a21oi_1 _1256_ (.A1(net382),
    .A2(_0486_),
    .Y(_0487_),
    .B1(net127));
 sg13g2_nor2_1 _1257_ (.A(_0429_),
    .B(net383),
    .Y(_0138_));
 sg13g2_a22oi_1 _1258_ (.Y(_0488_),
    .B1(net120),
    .B2(net329),
    .A2(net124),
    .A1(net293));
 sg13g2_inv_1 _1259_ (.Y(_0139_),
    .A(_0488_));
 sg13g2_a22oi_1 _1260_ (.Y(_0489_),
    .B1(_0370_),
    .B2(net341),
    .A2(net124),
    .A1(\addr_in[1] ));
 sg13g2_inv_1 _1261_ (.Y(_0140_),
    .A(net342));
 sg13g2_a22oi_1 _1262_ (.Y(_0490_),
    .B1(net119),
    .B2(net327),
    .A2(net125),
    .A1(\addr_in[2] ));
 sg13g2_inv_1 _1263_ (.Y(_0141_),
    .A(net328));
 sg13g2_a22oi_1 _1264_ (.Y(_0491_),
    .B1(net119),
    .B2(net335),
    .A2(net125),
    .A1(\addr_in[3] ));
 sg13g2_inv_1 _1265_ (.Y(_0142_),
    .A(net336));
 sg13g2_nor3_1 _1266_ (.A(_0205_),
    .B(net132),
    .C(_0340_),
    .Y(_0492_));
 sg13g2_nand2b_2 _1267_ (.Y(_0493_),
    .B(net1),
    .A_N(_0492_));
 sg13g2_inv_1 _1268_ (.Y(_0494_),
    .A(_0493_));
 sg13g2_nand2b_1 _1269_ (.Y(_0495_),
    .B(_0304_),
    .A_N(\i_display.v_count[0] ));
 sg13g2_a21oi_1 _1270_ (.A1(_0306_),
    .A2(_0495_),
    .Y(_0496_),
    .B1(_0365_));
 sg13g2_a21o_1 _1271_ (.A2(_0495_),
    .A1(_0306_),
    .B1(_0365_),
    .X(_0497_));
 sg13g2_nand2_1 _1272_ (.Y(_0498_),
    .A(\addr_in[1] ),
    .B(_0415_));
 sg13g2_nor2_1 _1273_ (.A(net293),
    .B(_0414_),
    .Y(_0499_));
 sg13g2_nor2_1 _1274_ (.A(\addr_in[1] ),
    .B(_0415_),
    .Y(_0500_));
 sg13g2_xor2_1 _1275_ (.B(_0415_),
    .A(net517),
    .X(_0501_));
 sg13g2_o21ai_1 _1276_ (.B1(_0498_),
    .Y(_0502_),
    .A1(_0499_),
    .A2(_0500_));
 sg13g2_nor2_1 _1277_ (.A(\addr_in[3] ),
    .B(_0420_),
    .Y(_0503_));
 sg13g2_xor2_1 _1278_ (.B(_0420_),
    .A(net540),
    .X(_0504_));
 sg13g2_and2_1 _1279_ (.A(net542),
    .B(_0423_),
    .X(_0505_));
 sg13g2_xor2_1 _1280_ (.B(_0423_),
    .A(\addr_in[2] ),
    .X(_0506_));
 sg13g2_and2_1 _1281_ (.A(_0504_),
    .B(_0506_),
    .X(_0507_));
 sg13g2_nor2b_1 _1282_ (.A(_0503_),
    .B_N(_0505_),
    .Y(_0508_));
 sg13g2_a221oi_1 _1283_ (.B2(_0507_),
    .C1(_0508_),
    .B1(_0502_),
    .A1(net540),
    .Y(_0509_),
    .A2(_0420_));
 sg13g2_nor2_1 _1284_ (.A(\addr_in[7] ),
    .B(_0416_),
    .Y(_0510_));
 sg13g2_xor2_1 _1285_ (.B(_0416_),
    .A(net537),
    .X(_0511_));
 sg13g2_nand2_1 _1286_ (.Y(_0512_),
    .A(net534),
    .B(_0417_));
 sg13g2_xor2_1 _1287_ (.B(_0417_),
    .A(net534),
    .X(_0513_));
 sg13g2_and2_1 _1288_ (.A(_0511_),
    .B(_0513_),
    .X(_0514_));
 sg13g2_nand2_1 _1289_ (.Y(_0515_),
    .A(\addr_in[5] ),
    .B(_0418_));
 sg13g2_nor2_1 _1290_ (.A(\addr_in[5] ),
    .B(_0418_),
    .Y(_0516_));
 sg13g2_xor2_1 _1291_ (.B(_0418_),
    .A(net547),
    .X(_0517_));
 sg13g2_nand2_1 _1292_ (.Y(_0518_),
    .A(net364),
    .B(_0419_));
 sg13g2_xor2_1 _1293_ (.B(_0419_),
    .A(net364),
    .X(_0519_));
 sg13g2_nand3_1 _1294_ (.B(_0517_),
    .C(_0519_),
    .A(_0514_),
    .Y(_0520_));
 sg13g2_o21ai_1 _1295_ (.B1(_0515_),
    .Y(_0521_),
    .A1(_0516_),
    .A2(_0518_));
 sg13g2_nor2_1 _1296_ (.A(_0510_),
    .B(_0512_),
    .Y(_0522_));
 sg13g2_a221oi_1 _1297_ (.B2(_0521_),
    .C1(_0522_),
    .B1(_0514_),
    .A1(\addr_in[7] ),
    .Y(_0523_),
    .A2(_0416_));
 sg13g2_o21ai_1 _1298_ (.B1(net538),
    .Y(_0524_),
    .A1(_0509_),
    .A2(_0520_));
 sg13g2_nand2_1 _1299_ (.Y(_0525_),
    .A(\addr_in[9] ),
    .B(_0424_));
 sg13g2_nor2_1 _1300_ (.A(\addr_in[9] ),
    .B(_0424_),
    .Y(_0526_));
 sg13g2_xor2_1 _1301_ (.B(_0424_),
    .A(net548),
    .X(_0527_));
 sg13g2_nand2_1 _1302_ (.Y(_0528_),
    .A(net362),
    .B(_0421_));
 sg13g2_xor2_1 _1303_ (.B(_0421_),
    .A(net362),
    .X(_0529_));
 sg13g2_and2_1 _1304_ (.A(_0527_),
    .B(_0529_),
    .X(_0530_));
 sg13g2_o21ai_1 _1305_ (.B1(_0525_),
    .Y(_0531_),
    .A1(_0526_),
    .A2(_0528_));
 sg13g2_a21o_1 _1306_ (.A2(_0530_),
    .A1(_0524_),
    .B1(_0531_),
    .X(_0532_));
 sg13g2_and2_1 _1307_ (.A(net122),
    .B(_0532_),
    .X(_0533_));
 sg13g2_and2_1 _1308_ (.A(net539),
    .B(_0533_),
    .X(_0534_));
 sg13g2_and4_1 _1309_ (.A(net510),
    .B(\addr_in[10] ),
    .C(net122),
    .D(_0532_),
    .X(_0535_));
 sg13g2_and3_1 _1310_ (.X(_0536_),
    .A(net332),
    .B(net301),
    .C(net526));
 sg13g2_and2_1 _1311_ (.A(_0535_),
    .B(_0536_),
    .X(_0537_));
 sg13g2_nand2_1 _1312_ (.Y(_0538_),
    .A(net536),
    .B(_0537_));
 sg13g2_and4_1 _1313_ (.A(net476),
    .B(net536),
    .C(_0535_),
    .D(_0536_),
    .X(_0539_));
 sg13g2_and3_1 _1314_ (.X(_0540_),
    .A(net524),
    .B(net530),
    .C(_0539_));
 sg13g2_and4_1 _1315_ (.A(net505),
    .B(\addr_in[18] ),
    .C(\addr_in[17] ),
    .D(_0539_),
    .X(_0541_));
 sg13g2_and3_1 _1316_ (.X(_0542_),
    .A(net350),
    .B(net374),
    .C(_0541_));
 sg13g2_nand4_1 _1317_ (.B(net350),
    .C(net374),
    .A(net323),
    .Y(_0543_),
    .D(net525));
 sg13g2_xnor2_1 _1318_ (.Y(_0544_),
    .A(net319),
    .B(_0543_));
 sg13g2_mux2_1 _1319_ (.A0(net8),
    .A1(_0544_),
    .S(net118),
    .X(_0143_));
 sg13g2_nor2_1 _1320_ (.A(_0414_),
    .B(_0497_),
    .Y(_0545_));
 sg13g2_o21ai_1 _1321_ (.B1(net117),
    .Y(_0546_),
    .A1(net293),
    .A2(_0545_));
 sg13g2_a21oi_1 _1322_ (.A1(net293),
    .A2(_0545_),
    .Y(_0144_),
    .B1(_0546_));
 sg13g2_nor2_1 _1323_ (.A(net517),
    .B(net123),
    .Y(_0547_));
 sg13g2_xnor2_1 _1324_ (.Y(_0548_),
    .A(_0499_),
    .B(_0501_));
 sg13g2_nor2_1 _1325_ (.A(_0497_),
    .B(_0548_),
    .Y(_0549_));
 sg13g2_nor3_1 _1326_ (.A(_0493_),
    .B(_0547_),
    .C(_0549_),
    .Y(_0145_));
 sg13g2_xnor2_1 _1327_ (.Y(_0550_),
    .A(_0502_),
    .B(_0506_));
 sg13g2_nand2_1 _1328_ (.Y(_0551_),
    .A(net121),
    .B(_0550_));
 sg13g2_o21ai_1 _1329_ (.B1(_0551_),
    .Y(_0552_),
    .A1(net542),
    .A2(net121));
 sg13g2_nor2_1 _1330_ (.A(_0493_),
    .B(_0552_),
    .Y(_0146_));
 sg13g2_a21oi_1 _1331_ (.A1(_0502_),
    .A2(_0506_),
    .Y(_0553_),
    .B1(_0505_));
 sg13g2_xor2_1 _1332_ (.B(_0553_),
    .A(_0504_),
    .X(_0554_));
 sg13g2_o21ai_1 _1333_ (.B1(net116),
    .Y(_0555_),
    .A1(net540),
    .A2(net121));
 sg13g2_a21oi_1 _1334_ (.A1(net121),
    .A2(_0554_),
    .Y(_0147_),
    .B1(_0555_));
 sg13g2_nand2b_1 _1335_ (.Y(_0556_),
    .B(_0519_),
    .A_N(_0509_));
 sg13g2_xor2_1 _1336_ (.B(_0519_),
    .A(net541),
    .X(_0557_));
 sg13g2_o21ai_1 _1337_ (.B1(net117),
    .Y(_0558_),
    .A1(net364),
    .A2(net123));
 sg13g2_a21oi_1 _1338_ (.A1(net123),
    .A2(_0557_),
    .Y(_0148_),
    .B1(_0558_));
 sg13g2_and2_1 _1339_ (.A(_0518_),
    .B(_0556_),
    .X(_0559_));
 sg13g2_xor2_1 _1340_ (.B(_0559_),
    .A(_0517_),
    .X(_0560_));
 sg13g2_o21ai_1 _1341_ (.B1(net116),
    .Y(_0561_),
    .A1(net547),
    .A2(net122));
 sg13g2_a21oi_1 _1342_ (.A1(net122),
    .A2(_0560_),
    .Y(_0149_),
    .B1(_0561_));
 sg13g2_a21oi_1 _1343_ (.A1(_0515_),
    .A2(_0559_),
    .Y(_0562_),
    .B1(_0516_));
 sg13g2_nand2_1 _1344_ (.Y(_0563_),
    .A(_0513_),
    .B(_0562_));
 sg13g2_xnor2_1 _1345_ (.Y(_0564_),
    .A(_0513_),
    .B(_0562_));
 sg13g2_o21ai_1 _1346_ (.B1(net116),
    .Y(_0565_),
    .A1(net534),
    .A2(net121));
 sg13g2_a21oi_1 _1347_ (.A1(net121),
    .A2(_0564_),
    .Y(_0150_),
    .B1(_0565_));
 sg13g2_nand2_1 _1348_ (.Y(_0566_),
    .A(_0512_),
    .B(_0563_));
 sg13g2_xnor2_1 _1349_ (.Y(_0567_),
    .A(_0511_),
    .B(_0566_));
 sg13g2_o21ai_1 _1350_ (.B1(net116),
    .Y(_0568_),
    .A1(net537),
    .A2(net121));
 sg13g2_a21oi_1 _1351_ (.A1(net121),
    .A2(_0567_),
    .Y(_0151_),
    .B1(_0568_));
 sg13g2_nand2_1 _1352_ (.Y(_0569_),
    .A(_0524_),
    .B(_0529_));
 sg13g2_xnor2_1 _1353_ (.Y(_0570_),
    .A(_0524_),
    .B(_0529_));
 sg13g2_o21ai_1 _1354_ (.B1(net117),
    .Y(_0571_),
    .A1(net362),
    .A2(net123));
 sg13g2_a21oi_1 _1355_ (.A1(net123),
    .A2(_0570_),
    .Y(_0152_),
    .B1(_0571_));
 sg13g2_nand2_1 _1356_ (.Y(_0572_),
    .A(_0528_),
    .B(_0569_));
 sg13g2_xnor2_1 _1357_ (.Y(_0573_),
    .A(_0527_),
    .B(_0572_));
 sg13g2_o21ai_1 _1358_ (.B1(net117),
    .Y(_0574_),
    .A1(net548),
    .A2(net123));
 sg13g2_a21oi_1 _1359_ (.A1(net123),
    .A2(_0573_),
    .Y(_0153_),
    .B1(_0574_));
 sg13g2_o21ai_1 _1360_ (.B1(net116),
    .Y(_0575_),
    .A1(net539),
    .A2(_0533_));
 sg13g2_nor2_1 _1361_ (.A(_0534_),
    .B(_0575_),
    .Y(_0154_));
 sg13g2_o21ai_1 _1362_ (.B1(net116),
    .Y(_0576_),
    .A1(net510),
    .A2(_0534_));
 sg13g2_nor2_1 _1363_ (.A(_0535_),
    .B(net511),
    .Y(_0155_));
 sg13g2_and2_1 _1364_ (.A(net526),
    .B(_0535_),
    .X(_0577_));
 sg13g2_o21ai_1 _1365_ (.B1(net116),
    .Y(_0578_),
    .A1(net526),
    .A2(_0535_));
 sg13g2_nor2_1 _1366_ (.A(_0577_),
    .B(net527),
    .Y(_0156_));
 sg13g2_o21ai_1 _1367_ (.B1(net116),
    .Y(_0579_),
    .A1(net301),
    .A2(_0577_));
 sg13g2_a21oi_1 _1368_ (.A1(net301),
    .A2(_0577_),
    .Y(_0157_),
    .B1(_0579_));
 sg13g2_a21oi_1 _1369_ (.A1(net301),
    .A2(_0577_),
    .Y(_0580_),
    .B1(net332));
 sg13g2_nor3_1 _1370_ (.A(_0493_),
    .B(_0537_),
    .C(net333),
    .Y(_0158_));
 sg13g2_o21ai_1 _1371_ (.B1(net118),
    .Y(_0581_),
    .A1(net536),
    .A2(_0537_));
 sg13g2_nor2b_1 _1372_ (.A(_0581_),
    .B_N(_0538_),
    .Y(_0159_));
 sg13g2_xor2_1 _1373_ (.B(_0538_),
    .A(net476),
    .X(_0582_));
 sg13g2_nor2_1 _1374_ (.A(_0493_),
    .B(net477),
    .Y(_0160_));
 sg13g2_and2_1 _1375_ (.A(net530),
    .B(_0539_),
    .X(_0583_));
 sg13g2_o21ai_1 _1376_ (.B1(net118),
    .Y(_0584_),
    .A1(net530),
    .A2(_0539_));
 sg13g2_nor2_1 _1377_ (.A(_0583_),
    .B(_0584_),
    .Y(_0161_));
 sg13g2_o21ai_1 _1378_ (.B1(net118),
    .Y(_0585_),
    .A1(net524),
    .A2(_0583_));
 sg13g2_nor2_1 _1379_ (.A(net531),
    .B(_0585_),
    .Y(_0162_));
 sg13g2_o21ai_1 _1380_ (.B1(net118),
    .Y(_0586_),
    .A1(net505),
    .A2(_0540_));
 sg13g2_nor2_1 _1381_ (.A(net506),
    .B(_0586_),
    .Y(_0163_));
 sg13g2_xnor2_1 _1382_ (.Y(_0587_),
    .A(net374),
    .B(net506));
 sg13g2_nor2_1 _1383_ (.A(_0493_),
    .B(_0587_),
    .Y(_0164_));
 sg13g2_a21oi_1 _1384_ (.A1(\addr_in[20] ),
    .A2(_0541_),
    .Y(_0588_),
    .B1(net350));
 sg13g2_nor3_1 _1385_ (.A(_0493_),
    .B(_0542_),
    .C(net351),
    .Y(_0165_));
 sg13g2_o21ai_1 _1386_ (.B1(net118),
    .Y(_0589_),
    .A1(net323),
    .A2(_0542_));
 sg13g2_nor2b_1 _1387_ (.A(_0589_),
    .B_N(_0543_),
    .Y(_0166_));
 sg13g2_nor2b_1 _1388_ (.A(_0200_),
    .B_N(\i_display.h_count[9] ),
    .Y(_0590_));
 sg13g2_a21oi_1 _1389_ (.A1(\i_display.h_count[10] ),
    .A2(_0201_),
    .Y(_0591_),
    .B1(_0590_));
 sg13g2_nand3_1 _1390_ (.B(net129),
    .C(_0209_),
    .A(net386),
    .Y(_0592_));
 sg13g2_a21oi_1 _1391_ (.A1(_0591_),
    .A2(net387),
    .Y(_0167_),
    .B1(net167));
 sg13g2_nand3_1 _1392_ (.B(net168),
    .C(_0202_),
    .A(\i_display.h_count[10] ),
    .Y(_0593_));
 sg13g2_nand2_1 _1393_ (.Y(_0594_),
    .A(net358),
    .B(_0303_));
 sg13g2_nand2_1 _1394_ (.Y(_0168_),
    .A(_0593_),
    .B(_0594_));
 sg13g2_xnor2_1 _1395_ (.Y(_0595_),
    .A(net551),
    .B(_0294_));
 sg13g2_nand2_1 _1396_ (.Y(_0169_),
    .A(net169),
    .B(net552));
 sg13g2_a21oi_1 _1397_ (.A1(\i_display.v_state[0] ),
    .A2(_0294_),
    .Y(_0596_),
    .B1(net528));
 sg13g2_o21ai_1 _1398_ (.B1(net169),
    .Y(_0170_),
    .A1(_0295_),
    .A2(net529));
 sg13g2_xor2_1 _1399_ (.B(_0205_),
    .A(net554),
    .X(_0597_));
 sg13g2_nand2_1 _1400_ (.Y(_0171_),
    .A(_0193_),
    .B(net555));
 sg13g2_a21oi_1 _1401_ (.A1(net160),
    .A2(net130),
    .Y(_0598_),
    .B1(net159));
 sg13g2_a21oi_1 _1402_ (.A1(net169),
    .A2(_0598_),
    .Y(_0172_),
    .B1(_0303_));
 sg13g2_dfrbpq_2 _1403_ (.RESET_B(net33),
    .D(_0011_),
    .Q(\i_display.v_count[6] ),
    .CLK(clknet_5_22__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1404_ (.RESET_B(net212),
    .D(net373),
    .Q(\i_display.v_count[7] ),
    .CLK(clknet_5_21__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1405_ (.RESET_B(net210),
    .D(_0013_),
    .Q(\i_display.v_count[8] ),
    .CLK(clknet_5_20__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1406_ (.RESET_B(net208),
    .D(_0014_),
    .Q(\i_display.v_count[9] ),
    .CLK(clknet_5_21__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1407_ (.RESET_B(net206),
    .D(_0015_),
    .Q(\i_display.v_count[10] ),
    .CLK(clknet_5_20__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1408_ (.RESET_B(net204),
    .D(net403),
    .Q(\i_display.v_count[0] ),
    .CLK(clknet_5_19__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1409_ (.RESET_B(net203),
    .D(net533),
    .Q(\i_display.v_count[1] ),
    .CLK(clknet_5_19__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1410_ (.RESET_B(net202),
    .D(net514),
    .Q(\i_display.v_count[2] ),
    .CLK(clknet_5_22__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1411_ (.RESET_B(net201),
    .D(net544),
    .Q(\i_display.v_count[3] ),
    .CLK(clknet_5_19__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1412_ (.RESET_B(net200),
    .D(net419),
    .Q(\i_display.v_count[4] ),
    .CLK(clknet_5_22__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1413_ (.RESET_B(net199),
    .D(net523),
    .Q(\i_display.v_count[5] ),
    .CLK(clknet_5_22__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1414_ (.RESET_B(net198),
    .D(_0022_),
    .Q(uo_out[6]),
    .CLK(clknet_5_27__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1415_ (.RESET_B(net196),
    .D(_0023_),
    .Q(uo_out[2]),
    .CLK(clknet_5_25__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1416_ (.RESET_B(net194),
    .D(net415),
    .Q(uo_out[5]),
    .CLK(clknet_5_27__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1417_ (.RESET_B(net192),
    .D(_0025_),
    .Q(uo_out[1]),
    .CLK(clknet_5_25__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1418_ (.RESET_B(net190),
    .D(net407),
    .Q(uo_out[4]),
    .CLK(clknet_5_26__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1419_ (.RESET_B(net34),
    .D(_0027_),
    .Q(uo_out[0]),
    .CLK(clknet_5_26__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1420_ (.RESET_B(net70),
    .D(net282),
    .Q(hsync_r),
    .CLK(clknet_5_19__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1421_ (.RESET_B(net188),
    .D(net318),
    .Q(vsync_r),
    .CLK(clknet_5_7__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1422_ (.RESET_B(net186),
    .D(net365),
    .Q(\i_qpsi.addr[4] ),
    .CLK(clknet_5_14__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1423_ (.RESET_B(net185),
    .D(net292),
    .Q(\i_qpsi.addr[5] ),
    .CLK(clknet_5_12__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1424_ (.RESET_B(net184),
    .D(net290),
    .Q(\i_qpsi.addr[6] ),
    .CLK(clknet_5_9__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1425_ (.RESET_B(net183),
    .D(net308),
    .Q(\i_qpsi.addr[7] ),
    .CLK(clknet_5_8__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1426_ (.RESET_B(net182),
    .D(net363),
    .Q(\i_qpsi.addr[8] ),
    .CLK(clknet_5_12__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1427_ (.RESET_B(net181),
    .D(net300),
    .Q(\i_qpsi.addr[9] ),
    .CLK(clknet_5_9__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1428_ (.RESET_B(net180),
    .D(net296),
    .Q(\i_qpsi.addr[10] ),
    .CLK(clknet_5_8__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1429_ (.RESET_B(net179),
    .D(net312),
    .Q(\i_qpsi.addr[11] ),
    .CLK(clknet_5_8__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1430_ (.RESET_B(net178),
    .D(net316),
    .Q(\i_qpsi.addr[12] ),
    .CLK(clknet_5_14__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1431_ (.RESET_B(net177),
    .D(net286),
    .Q(\i_qpsi.addr[13] ),
    .CLK(clknet_5_14__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1432_ (.RESET_B(net176),
    .D(net322),
    .Q(\i_qpsi.addr[14] ),
    .CLK(clknet_5_8__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1433_ (.RESET_B(net175),
    .D(net306),
    .Q(\i_qpsi.addr[15] ),
    .CLK(clknet_5_10__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1434_ (.RESET_B(net174),
    .D(net298),
    .Q(\i_qpsi.addr[16] ),
    .CLK(clknet_5_14__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1435_ (.RESET_B(net173),
    .D(net280),
    .Q(\i_qpsi.addr[17] ),
    .CLK(clknet_5_14__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1436_ (.RESET_B(net115),
    .D(net288),
    .Q(\i_qpsi.addr[18] ),
    .CLK(clknet_5_11__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1437_ (.RESET_B(net114),
    .D(net310),
    .Q(\i_qpsi.addr[19] ),
    .CLK(clknet_5_10__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1438_ (.RESET_B(net113),
    .D(net375),
    .Q(\i_qpsi.addr[20] ),
    .CLK(clknet_5_15__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1439_ (.RESET_B(net112),
    .D(_0045_),
    .Q(\i_qpsi.addr[21] ),
    .CLK(clknet_5_15__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1440_ (.RESET_B(net111),
    .D(net324),
    .Q(\i_qpsi.addr[22] ),
    .CLK(clknet_5_11__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1441_ (.RESET_B(net110),
    .D(net320),
    .Q(\i_qpsi.addr[23] ),
    .CLK(clknet_5_10__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1442_ (.RESET_B(net109),
    .D(_0048_),
    .Q(\i_qpsi.spi_clk ),
    .CLK(clknet_5_15__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1443_ (.RESET_B(net107),
    .D(net546),
    .Q(\i_qpsi.bits_remaining[0] ),
    .CLK(clknet_5_13__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1444_ (.RESET_B(net105),
    .D(_0050_),
    .Q(\i_qpsi.bits_remaining[1] ),
    .CLK(clknet_5_24__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1445_ (.RESET_B(net103),
    .D(net445),
    .Q(\i_qpsi.bits_remaining[2] ),
    .CLK(clknet_5_24__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1446_ (.RESET_B(net101),
    .D(_0052_),
    .Q(\i_qpsi.fsm_state[0] ),
    .CLK(clknet_5_15__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1447_ (.RESET_B(net99),
    .D(_0053_),
    .Q(\i_qpsi.fsm_state[1] ),
    .CLK(clknet_5_15__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1448_ (.RESET_B(net97),
    .D(_0054_),
    .Q(\i_qpsi.fsm_state[2] ),
    .CLK(clknet_5_14__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1449_ (.RESET_B(net95),
    .D(net349),
    .Q(\i_qpsi.data[0] ),
    .CLK(clknet_5_31__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1450_ (.RESET_B(net94),
    .D(net377),
    .Q(\i_qpsi.data[1] ),
    .CLK(clknet_5_27__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1451_ (.RESET_B(net93),
    .D(_0057_),
    .Q(\i_qpsi.data[2] ),
    .CLK(clknet_5_27__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1452_ (.RESET_B(net92),
    .D(net355),
    .Q(\i_qpsi.data[3] ),
    .CLK(clknet_5_31__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1453_ (.RESET_B(net91),
    .D(net331),
    .Q(\i_qpsi.data[4] ),
    .CLK(clknet_5_30__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1454_ (.RESET_B(net90),
    .D(net304),
    .Q(\i_qpsi.data[5] ),
    .CLK(clknet_5_25__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1455_ (.RESET_B(net89),
    .D(net284),
    .Q(\i_qpsi.data[6] ),
    .CLK(clknet_5_30__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1456_ (.RESET_B(net71),
    .D(net314),
    .Q(\i_qpsi.data[7] ),
    .CLK(clknet_5_27__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1457_ (.RESET_B(net72),
    .D(\i_qpsi.spi_data_in[0] ),
    .Q(\i_qpsi.spi_miso_buf[0] ),
    .CLK(clknet_5_30__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1458_ (.RESET_B(net73),
    .D(\i_qpsi.spi_data_in[1] ),
    .Q(\i_qpsi.spi_miso_buf[1] ),
    .CLK(clknet_5_26__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1459_ (.RESET_B(net74),
    .D(net12),
    .Q(\i_qpsi.spi_miso_buf[2] ),
    .CLK(clknet_5_30__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1460_ (.RESET_B(net75),
    .D(net13),
    .Q(\i_qpsi.spi_miso_buf[3] ),
    .CLK(clknet_5_25__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1461_ (.RESET_B(net76),
    .D(net271),
    .Q(\i_qpsi.spi_miso_buf[4] ),
    .CLK(clknet_5_30__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1462_ (.RESET_B(net77),
    .D(net275),
    .Q(\i_qpsi.spi_miso_buf[5] ),
    .CLK(clknet_5_26__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1463_ (.RESET_B(net78),
    .D(net272),
    .Q(\i_qpsi.spi_miso_buf[6] ),
    .CLK(clknet_5_31__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1464_ (.RESET_B(net79),
    .D(net274),
    .Q(\i_qpsi.spi_miso_buf[7] ),
    .CLK(clknet_5_28__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1465_ (.RESET_B(net80),
    .D(net270),
    .Q(\i_qpsi.spi_miso_buf[8] ),
    .CLK(clknet_5_30__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1466_ (.RESET_B(net81),
    .D(net276),
    .Q(\i_qpsi.spi_miso_buf[9] ),
    .CLK(clknet_5_27__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1467_ (.RESET_B(net215),
    .D(net273),
    .Q(\i_qpsi.spi_miso_buf[10] ),
    .CLK(clknet_5_31__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1468_ (.RESET_B(net88),
    .D(net277),
    .Q(\i_qpsi.spi_miso_buf[11] ),
    .CLK(clknet_5_31__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1469_ (.RESET_B(net87),
    .D(_0063_),
    .Q(\i_display.cfg[0] ),
    .CLK(clknet_5_13__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1470_ (.RESET_B(net86),
    .D(net340),
    .Q(\i_display.cfg[1] ),
    .CLK(clknet_5_24__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1471_ (.RESET_B(net85),
    .D(_0065_),
    .Q(\i_display.cfg[2] ),
    .CLK(clknet_5_19__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1472_ (.RESET_B(net84),
    .D(_0066_),
    .Q(\i_display.cfg[3] ),
    .CLK(clknet_5_22__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1473_ (.RESET_B(net83),
    .D(net401),
    .Q(\i_display.cfg[4] ),
    .CLK(clknet_5_23__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1474_ (.RESET_B(net82),
    .D(net367),
    .Q(\i_display.cfg[5] ),
    .CLK(clknet_5_23__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1475_ (.RESET_B(net69),
    .D(_0069_),
    .Q(\i_display.cfg[6] ),
    .CLK(clknet_5_13__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1476_ (.RESET_B(net68),
    .D(_0070_),
    .Q(\i_display.cfg[7] ),
    .CLK(clknet_5_24__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1477_ (.RESET_B(net67),
    .D(_0071_),
    .Q(\i_display.cfg[8] ),
    .CLK(clknet_5_25__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1478_ (.RESET_B(net66),
    .D(net434),
    .Q(\i_display.cfg[9] ),
    .CLK(clknet_5_28__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1479_ (.RESET_B(net65),
    .D(_0073_),
    .Q(\i_display.cfg[10] ),
    .CLK(clknet_5_29__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1480_ (.RESET_B(net64),
    .D(_0074_),
    .Q(\i_display.cfg[11] ),
    .CLK(clknet_5_13__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1481_ (.RESET_B(net63),
    .D(_0075_),
    .Q(\i_display.cfg[12] ),
    .CLK(clknet_5_13__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1482_ (.RESET_B(net62),
    .D(net409),
    .Q(\i_display.cfg[13] ),
    .CLK(clknet_5_24__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1483_ (.RESET_B(net61),
    .D(_0077_),
    .Q(\i_display.cfg[14] ),
    .CLK(clknet_5_25__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1484_ (.RESET_B(net60),
    .D(net427),
    .Q(\i_display.cfg[15] ),
    .CLK(clknet_5_29__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1485_ (.RESET_B(net59),
    .D(net470),
    .Q(\i_display.cfg[16] ),
    .CLK(clknet_5_29__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1486_ (.RESET_B(net58),
    .D(net432),
    .Q(\i_display.cfg[17] ),
    .CLK(clknet_5_19__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1487_ (.RESET_B(net57),
    .D(_0081_),
    .Q(\i_display.cfg[18] ),
    .CLK(clknet_5_7__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1488_ (.RESET_B(net56),
    .D(net453),
    .Q(\i_display.cfg[19] ),
    .CLK(clknet_5_24__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1489_ (.RESET_B(net55),
    .D(_0083_),
    .Q(\i_display.cfg[20] ),
    .CLK(clknet_5_29__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1490_ (.RESET_B(net54),
    .D(net465),
    .Q(\i_display.cfg[21] ),
    .CLK(clknet_5_29__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1491_ (.RESET_B(net53),
    .D(net417),
    .Q(\i_display.cfg[22] ),
    .CLK(clknet_5_23__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1492_ (.RESET_B(net52),
    .D(_0086_),
    .Q(\i_display.cfg[23] ),
    .CLK(clknet_5_23__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1493_ (.RESET_B(net51),
    .D(_0087_),
    .Q(\i_display.cfg[24] ),
    .CLK(clknet_5_23__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1494_ (.RESET_B(net50),
    .D(net456),
    .Q(\i_display.cfg[25] ),
    .CLK(clknet_5_21__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1495_ (.RESET_B(net49),
    .D(_0089_),
    .Q(\i_display.cfg[26] ),
    .CLK(clknet_5_21__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1496_ (.RESET_B(net48),
    .D(net430),
    .Q(\i_display.cfg[27] ),
    .CLK(clknet_5_21__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1497_ (.RESET_B(net47),
    .D(_0091_),
    .Q(\i_display.cfg[28] ),
    .CLK(clknet_5_21__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1498_ (.RESET_B(net46),
    .D(net385),
    .Q(\i_display.cfg[29] ),
    .CLK(clknet_5_20__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1499_ (.RESET_B(net45),
    .D(net347),
    .Q(\i_display.cfg[30] ),
    .CLK(clknet_5_20__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1500_ (.RESET_B(net44),
    .D(_0094_),
    .Q(\i_display.cfg[31] ),
    .CLK(clknet_5_17__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1501_ (.RESET_B(net43),
    .D(net344),
    .Q(\i_display.cfg[32] ),
    .CLK(clknet_5_16__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1502_ (.RESET_B(net42),
    .D(_0096_),
    .Q(\i_display.cfg[33] ),
    .CLK(clknet_5_5__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1503_ (.RESET_B(net41),
    .D(_0097_),
    .Q(\i_display.cfg[34] ),
    .CLK(clknet_5_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1504_ (.RESET_B(net40),
    .D(_0098_),
    .Q(\i_display.cfg[35] ),
    .CLK(clknet_5_0__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1505_ (.RESET_B(net39),
    .D(_0099_),
    .Q(\i_display.cfg[36] ),
    .CLK(clknet_5_0__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1506_ (.RESET_B(net38),
    .D(net379),
    .Q(\i_display.cfg[37] ),
    .CLK(clknet_5_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1507_ (.RESET_B(net37),
    .D(net326),
    .Q(\i_display.cfg[38] ),
    .CLK(clknet_5_17__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1508_ (.RESET_B(net36),
    .D(_0102_),
    .Q(\i_display.cfg[39] ),
    .CLK(clknet_5_20__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1509_ (.RESET_B(net35),
    .D(_0103_),
    .Q(\i_display.cfg[40] ),
    .CLK(clknet_5_20__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1510_ (.RESET_B(net32),
    .D(net497),
    .Q(\i_display.cfg[41] ),
    .CLK(clknet_5_16__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1511_ (.RESET_B(net31),
    .D(net482),
    .Q(\i_display.cfg[42] ),
    .CLK(clknet_5_5__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1512_ (.RESET_B(net30),
    .D(_0106_),
    .Q(\i_display.cfg[43] ),
    .CLK(clknet_5_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1513_ (.RESET_B(net29),
    .D(net449),
    .Q(\i_display.cfg[44] ),
    .CLK(clknet_5_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1514_ (.RESET_B(net28),
    .D(_0108_),
    .Q(\i_display.cfg[45] ),
    .CLK(clknet_5_4__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1515_ (.RESET_B(net27),
    .D(_0109_),
    .Q(\i_display.cfg[46] ),
    .CLK(clknet_5_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1516_ (.RESET_B(net26),
    .D(_0110_),
    .Q(\i_display.cfg[47] ),
    .CLK(clknet_5_16__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1517_ (.RESET_B(net25),
    .D(net468),
    .Q(\i_display.cfg[48] ),
    .CLK(clknet_5_17__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1518_ (.RESET_B(net24),
    .D(_0112_),
    .Q(\i_display.cfg[49] ),
    .CLK(clknet_5_17__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1519_ (.RESET_B(net23),
    .D(net460),
    .Q(\i_display.cfg[50] ),
    .CLK(clknet_5_16__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1520_ (.RESET_B(net22),
    .D(_0114_),
    .Q(\i_display.cfg[51] ),
    .CLK(clknet_5_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1521_ (.RESET_B(net21),
    .D(net439),
    .Q(\i_display.cfg[52] ),
    .CLK(clknet_5_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1522_ (.RESET_B(net20),
    .D(net338),
    .Q(\i_display.cfg[53] ),
    .CLK(clknet_5_0__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1523_ (.RESET_B(net19),
    .D(_0117_),
    .Q(\i_display.cfg[54] ),
    .CLK(clknet_5_0__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1524_ (.RESET_B(net18),
    .D(_0118_),
    .Q(\i_display.cfg[55] ),
    .CLK(clknet_5_1__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1525_ (.RESET_B(net17),
    .D(_0119_),
    .Q(\i_display.cfg[56] ),
    .CLK(clknet_5_5__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1526_ (.RESET_B(net16),
    .D(_0120_),
    .Q(\i_display.cfg[57] ),
    .CLK(clknet_5_18__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1527_ (.RESET_B(net264),
    .D(_0121_),
    .Q(\i_display.cfg[58] ),
    .CLK(clknet_5_16__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1528_ (.RESET_B(net263),
    .D(_0122_),
    .Q(\i_display.cfg[59] ),
    .CLK(clknet_5_5__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1529_ (.RESET_B(net262),
    .D(net488),
    .Q(\i_display.cfg[60] ),
    .CLK(clknet_5_4__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1530_ (.RESET_B(net261),
    .D(net521),
    .Q(\i_display.cfg[61] ),
    .CLK(clknet_5_0__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1531_ (.RESET_B(net260),
    .D(net500),
    .Q(\i_display.cfg[62] ),
    .CLK(clknet_5_2__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1532_ (.RESET_B(net259),
    .D(net486),
    .Q(\i_display.cfg[63] ),
    .CLK(clknet_5_0__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1533_ (.RESET_B(net253),
    .D(_0127_),
    .Q(\i_display.cfg[64] ),
    .CLK(clknet_5_2__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1534_ (.RESET_B(net252),
    .D(_0128_),
    .Q(\i_display.cfg[65] ),
    .CLK(clknet_5_3__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1535_ (.RESET_B(net251),
    .D(_0129_),
    .Q(\i_display.cfg[66] ),
    .CLK(clknet_5_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1536_ (.RESET_B(net250),
    .D(_0130_),
    .Q(\i_display.cfg[67] ),
    .CLK(clknet_5_6__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1537_ (.RESET_B(net249),
    .D(_0131_),
    .Q(\i_display.cfg[68] ),
    .CLK(clknet_5_7__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1538_ (.RESET_B(net248),
    .D(_0132_),
    .Q(\i_display.cfg[69] ),
    .CLK(clknet_5_7__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1539_ (.RESET_B(net247),
    .D(_0133_),
    .Q(\i_display.cfg[70] ),
    .CLK(clknet_5_18__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1540_ (.RESET_B(net246),
    .D(net451),
    .Q(\i_display.cfg[71] ),
    .CLK(clknet_5_18__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1541_ (.RESET_B(net245),
    .D(_0135_),
    .Q(\i_display.cfg[72] ),
    .CLK(clknet_5_18__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1542_ (.RESET_B(net244),
    .D(net479),
    .Q(\i_display.cfg[73] ),
    .CLK(clknet_5_7__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1543_ (.RESET_B(net243),
    .D(net421),
    .Q(\i_display.cfg[74] ),
    .CLK(clknet_5_7__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1544_ (.RESET_B(net222),
    .D(\i_qpsi.spi_clk ),
    .Q(\i_qpsi.spi_clk_n ),
    .CLK(net267));
 sg13g2_dfrbpq_1 _1545_ (.RESET_B(net242),
    .D(_0009_),
    .Q(\i_qpsi.valid ),
    .CLK(clknet_5_26__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1546_ (.RESET_B(net241),
    .D(_0138_),
    .Q(\i_qpsi.spi_data_oe[0] ),
    .CLK(clknet_5_26__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1547_ (.RESET_B(net239),
    .D(_0139_),
    .Q(\i_qpsi.addr[0] ),
    .CLK(clknet_5_12__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1548_ (.RESET_B(net237),
    .D(_0140_),
    .Q(\i_qpsi.addr[1] ),
    .CLK(clknet_5_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1549_ (.RESET_B(net235),
    .D(_0141_),
    .Q(\i_qpsi.addr[2] ),
    .CLK(clknet_5_2__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1550_ (.RESET_B(net233),
    .D(_0142_),
    .Q(\i_qpsi.addr[3] ),
    .CLK(clknet_5_9__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1551_ (.RESET_B(net223),
    .D(_0143_),
    .Q(\addr_in[23] ),
    .CLK(clknet_5_10__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1552_ (.RESET_B(net224),
    .D(net462),
    .Q(\i_display.h_count[0] ),
    .CLK(clknet_5_17__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1553_ (.RESET_B(net225),
    .D(_0001_),
    .Q(\i_display.h_count[1] ),
    .CLK(clknet_5_18__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1554_ (.RESET_B(net226),
    .D(_0002_),
    .Q(\i_display.h_count[2] ),
    .CLK(clknet_5_16__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1555_ (.RESET_B(net227),
    .D(_0003_),
    .Q(\i_display.h_count[3] ),
    .CLK(clknet_5_5__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1556_ (.RESET_B(net228),
    .D(net357),
    .Q(\i_display.h_count[4] ),
    .CLK(clknet_5_5__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1557_ (.RESET_B(net229),
    .D(net390),
    .Q(\i_display.h_count[5] ),
    .CLK(clknet_5_4__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1558_ (.RESET_B(net230),
    .D(net516),
    .Q(\i_display.h_count[6] ),
    .CLK(clknet_5_1__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1559_ (.RESET_B(net254),
    .D(_0007_),
    .Q(\i_display.h_count[7] ),
    .CLK(clknet_5_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1560_ (.RESET_B(net231),
    .D(net411),
    .Q(\i_display.h_count[8] ),
    .CLK(clknet_5_6__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1561_ (.RESET_B(net221),
    .D(net294),
    .Q(\addr_in[0] ),
    .CLK(clknet_5_12__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1562_ (.RESET_B(net219),
    .D(_0145_),
    .Q(\addr_in[1] ),
    .CLK(clknet_5_13__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1563_ (.RESET_B(net217),
    .D(_0146_),
    .Q(\addr_in[2] ),
    .CLK(clknet_5_2__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1564_ (.RESET_B(net214),
    .D(_0147_),
    .Q(\addr_in[3] ),
    .CLK(clknet_5_2__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1565_ (.RESET_B(net211),
    .D(_0148_),
    .Q(\addr_in[4] ),
    .CLK(clknet_5_3__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1566_ (.RESET_B(net207),
    .D(_0149_),
    .Q(\addr_in[5] ),
    .CLK(clknet_5_3__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1567_ (.RESET_B(net197),
    .D(net535),
    .Q(\addr_in[6] ),
    .CLK(clknet_5_3__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1568_ (.RESET_B(net193),
    .D(_0151_),
    .Q(\addr_in[7] ),
    .CLK(clknet_5_2__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1569_ (.RESET_B(net189),
    .D(_0152_),
    .Q(\addr_in[8] ),
    .CLK(clknet_5_12__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1570_ (.RESET_B(net108),
    .D(_0153_),
    .Q(\addr_in[9] ),
    .CLK(clknet_5_6__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1571_ (.RESET_B(net104),
    .D(_0154_),
    .Q(\addr_in[10] ),
    .CLK(clknet_5_9__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1572_ (.RESET_B(net100),
    .D(net512),
    .Q(\addr_in[11] ),
    .CLK(clknet_5_9__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1573_ (.RESET_B(net96),
    .D(_0156_),
    .Q(\addr_in[12] ),
    .CLK(clknet_5_12__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1574_ (.RESET_B(net238),
    .D(net302),
    .Q(\addr_in[13] ),
    .CLK(clknet_5_9__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1575_ (.RESET_B(net234),
    .D(net334),
    .Q(\addr_in[14] ),
    .CLK(clknet_5_8__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1576_ (.RESET_B(net220),
    .D(_0159_),
    .Q(\addr_in[15] ),
    .CLK(clknet_5_8__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1577_ (.RESET_B(net216),
    .D(_0160_),
    .Q(\addr_in[16] ),
    .CLK(clknet_5_11__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1578_ (.RESET_B(net209),
    .D(_0161_),
    .Q(\addr_in[17] ),
    .CLK(clknet_5_11__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1579_ (.RESET_B(net195),
    .D(_0162_),
    .Q(\addr_in[18] ),
    .CLK(clknet_5_10__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1580_ (.RESET_B(net187),
    .D(_0163_),
    .Q(\addr_in[19] ),
    .CLK(clknet_5_10__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1581_ (.RESET_B(net102),
    .D(_0164_),
    .Q(\addr_in[20] ),
    .CLK(clknet_5_15__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1582_ (.RESET_B(net240),
    .D(net352),
    .Q(\addr_in[21] ),
    .CLK(clknet_5_11__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1583_ (.RESET_B(net255),
    .D(_0166_),
    .Q(\addr_in[22] ),
    .CLK(clknet_5_11__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1584_ (.RESET_B(net256),
    .D(net3),
    .Q(\i_display.cfg_data_sync[0] ),
    .CLK(clknet_5_29__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1585_ (.RESET_B(net257),
    .D(net268),
    .Q(\i_display.cfg_data_sync[1] ),
    .CLK(clknet_5_28__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1586_ (.RESET_B(net258),
    .D(net2),
    .Q(\i_display.cfg_clk_sync[0] ),
    .CLK(clknet_5_28__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1587_ (.RESET_B(net106),
    .D(net269),
    .Q(\i_display.cfg_clk_sync[1] ),
    .CLK(clknet_5_28__leaf_clk_regs));
 sg13g2_dfrbpq_1 _1588_ (.RESET_B(net232),
    .D(net278),
    .Q(\i_display.cfg_clk_sync[2] ),
    .CLK(clknet_5_28__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1589_ (.RESET_B(net213),
    .D(net388),
    .Q(\i_display.h_count[9] ),
    .CLK(clknet_5_6__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1590_ (.RESET_B(net205),
    .D(net359),
    .Q(\i_display.h_count[10] ),
    .CLK(clknet_5_6__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1591_ (.RESET_B(net191),
    .D(_0169_),
    .Q(\i_display.v_state[0] ),
    .CLK(clknet_5_22__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1592_ (.RESET_B(net98),
    .D(_0170_),
    .Q(\i_display.v_state[1] ),
    .CLK(clknet_5_23__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1593_ (.RESET_B(net218),
    .D(_0171_),
    .Q(\i_display.h_state[0] ),
    .CLK(clknet_5_17__leaf_clk_regs));
 sg13g2_dfrbpq_2 _1594_ (.RESET_B(net236),
    .D(_0172_),
    .Q(\i_display.h_state[1] ),
    .CLK(clknet_5_18__leaf_clk_regs));
 sg13g2_tiehi _1525__17 (.L_HI(net17));
 sg13g2_tiehi _1524__18 (.L_HI(net18));
 sg13g2_tiehi _1523__19 (.L_HI(net19));
 sg13g2_tiehi _1522__20 (.L_HI(net20));
 sg13g2_tiehi _1521__21 (.L_HI(net21));
 sg13g2_tiehi _1520__22 (.L_HI(net22));
 sg13g2_tiehi _1519__23 (.L_HI(net23));
 sg13g2_tiehi _1518__24 (.L_HI(net24));
 sg13g2_tiehi _1517__25 (.L_HI(net25));
 sg13g2_tiehi _1516__26 (.L_HI(net26));
 sg13g2_tiehi _1515__27 (.L_HI(net27));
 sg13g2_tiehi _1514__28 (.L_HI(net28));
 sg13g2_tiehi _1513__29 (.L_HI(net29));
 sg13g2_tiehi _1512__30 (.L_HI(net30));
 sg13g2_tiehi _1511__31 (.L_HI(net31));
 sg13g2_tiehi _1510__32 (.L_HI(net32));
 sg13g2_tiehi _1403__33 (.L_HI(net33));
 sg13g2_tiehi _1419__34 (.L_HI(net34));
 sg13g2_tiehi _1509__35 (.L_HI(net35));
 sg13g2_tiehi _1508__36 (.L_HI(net36));
 sg13g2_tiehi _1507__37 (.L_HI(net37));
 sg13g2_tiehi _1506__38 (.L_HI(net38));
 sg13g2_tiehi _1505__39 (.L_HI(net39));
 sg13g2_tiehi _1504__40 (.L_HI(net40));
 sg13g2_tiehi _1503__41 (.L_HI(net41));
 sg13g2_tiehi _1502__42 (.L_HI(net42));
 sg13g2_tiehi _1501__43 (.L_HI(net43));
 sg13g2_tiehi _1500__44 (.L_HI(net44));
 sg13g2_tiehi _1499__45 (.L_HI(net45));
 sg13g2_tiehi _1498__46 (.L_HI(net46));
 sg13g2_tiehi _1497__47 (.L_HI(net47));
 sg13g2_tiehi _1496__48 (.L_HI(net48));
 sg13g2_tiehi _1495__49 (.L_HI(net49));
 sg13g2_tiehi _1494__50 (.L_HI(net50));
 sg13g2_tiehi _1493__51 (.L_HI(net51));
 sg13g2_tiehi _1492__52 (.L_HI(net52));
 sg13g2_tiehi _1491__53 (.L_HI(net53));
 sg13g2_tiehi _1490__54 (.L_HI(net54));
 sg13g2_tiehi _1489__55 (.L_HI(net55));
 sg13g2_tiehi _1488__56 (.L_HI(net56));
 sg13g2_tiehi _1487__57 (.L_HI(net57));
 sg13g2_tiehi _1486__58 (.L_HI(net58));
 sg13g2_tiehi _1485__59 (.L_HI(net59));
 sg13g2_tiehi _1484__60 (.L_HI(net60));
 sg13g2_tiehi _1483__61 (.L_HI(net61));
 sg13g2_tiehi _1482__62 (.L_HI(net62));
 sg13g2_tiehi _1481__63 (.L_HI(net63));
 sg13g2_tiehi _1480__64 (.L_HI(net64));
 sg13g2_tiehi _1479__65 (.L_HI(net65));
 sg13g2_tiehi _1478__66 (.L_HI(net66));
 sg13g2_tiehi _1477__67 (.L_HI(net67));
 sg13g2_tiehi _1476__68 (.L_HI(net68));
 sg13g2_tiehi _1475__69 (.L_HI(net69));
 sg13g2_tiehi _1420__70 (.L_HI(net70));
 sg13g2_tiehi _1456__71 (.L_HI(net71));
 sg13g2_tiehi _1457__72 (.L_HI(net72));
 sg13g2_tiehi _1458__73 (.L_HI(net73));
 sg13g2_tiehi _1459__74 (.L_HI(net74));
 sg13g2_tiehi _1460__75 (.L_HI(net75));
 sg13g2_tiehi _1461__76 (.L_HI(net76));
 sg13g2_tiehi _1462__77 (.L_HI(net77));
 sg13g2_tiehi _1463__78 (.L_HI(net78));
 sg13g2_tiehi _1464__79 (.L_HI(net79));
 sg13g2_tiehi _1465__80 (.L_HI(net80));
 sg13g2_tiehi _1466__81 (.L_HI(net81));
 sg13g2_tiehi _1474__82 (.L_HI(net82));
 sg13g2_tiehi _1473__83 (.L_HI(net83));
 sg13g2_tiehi _1472__84 (.L_HI(net84));
 sg13g2_tiehi _1471__85 (.L_HI(net85));
 sg13g2_tiehi _1470__86 (.L_HI(net86));
 sg13g2_tiehi _1469__87 (.L_HI(net87));
 sg13g2_tiehi _1468__88 (.L_HI(net88));
 sg13g2_tiehi _1455__89 (.L_HI(net89));
 sg13g2_tiehi _1454__90 (.L_HI(net90));
 sg13g2_tiehi _1453__91 (.L_HI(net91));
 sg13g2_tiehi _1452__92 (.L_HI(net92));
 sg13g2_tiehi _1451__93 (.L_HI(net93));
 sg13g2_tiehi _1450__94 (.L_HI(net94));
 sg13g2_tiehi _1449__95 (.L_HI(net95));
 sg13g2_tiehi _1573__96 (.L_HI(net96));
 sg13g2_tiehi _1448__97 (.L_HI(net97));
 sg13g2_tiehi _1592__98 (.L_HI(net98));
 sg13g2_tiehi _1447__99 (.L_HI(net99));
 sg13g2_tiehi _1572__100 (.L_HI(net100));
 sg13g2_tiehi _1446__101 (.L_HI(net101));
 sg13g2_tiehi _1581__102 (.L_HI(net102));
 sg13g2_tiehi _1445__103 (.L_HI(net103));
 sg13g2_tiehi _1571__104 (.L_HI(net104));
 sg13g2_tiehi _1444__105 (.L_HI(net105));
 sg13g2_tiehi _1587__106 (.L_HI(net106));
 sg13g2_tiehi _1443__107 (.L_HI(net107));
 sg13g2_tiehi _1570__108 (.L_HI(net108));
 sg13g2_tiehi _1442__109 (.L_HI(net109));
 sg13g2_tiehi _1441__110 (.L_HI(net110));
 sg13g2_tiehi _1440__111 (.L_HI(net111));
 sg13g2_tiehi _1439__112 (.L_HI(net112));
 sg13g2_tiehi _1438__113 (.L_HI(net113));
 sg13g2_tiehi _1437__114 (.L_HI(net114));
 sg13g2_tiehi _1436__115 (.L_HI(net115));
 sg13g2_tiehi _1435__116 (.L_HI(net173));
 sg13g2_tiehi _1434__117 (.L_HI(net174));
 sg13g2_tiehi _1433__118 (.L_HI(net175));
 sg13g2_tiehi _1432__119 (.L_HI(net176));
 sg13g2_tiehi _1431__120 (.L_HI(net177));
 sg13g2_tiehi _1430__121 (.L_HI(net178));
 sg13g2_tiehi _1429__122 (.L_HI(net179));
 sg13g2_tiehi _1428__123 (.L_HI(net180));
 sg13g2_tiehi _1427__124 (.L_HI(net181));
 sg13g2_tiehi _1426__125 (.L_HI(net182));
 sg13g2_tiehi _1425__126 (.L_HI(net183));
 sg13g2_tiehi _1424__127 (.L_HI(net184));
 sg13g2_tiehi _1423__128 (.L_HI(net185));
 sg13g2_tiehi _1422__129 (.L_HI(net186));
 sg13g2_tiehi _1580__130 (.L_HI(net187));
 sg13g2_tiehi _1421__131 (.L_HI(net188));
 sg13g2_tiehi _1569__132 (.L_HI(net189));
 sg13g2_tiehi _1418__133 (.L_HI(net190));
 sg13g2_tiehi _1591__134 (.L_HI(net191));
 sg13g2_tiehi _1417__135 (.L_HI(net192));
 sg13g2_tiehi _1568__136 (.L_HI(net193));
 sg13g2_tiehi _1416__137 (.L_HI(net194));
 sg13g2_tiehi _1579__138 (.L_HI(net195));
 sg13g2_tiehi _1415__139 (.L_HI(net196));
 sg13g2_tiehi _1567__140 (.L_HI(net197));
 sg13g2_tiehi _1414__141 (.L_HI(net198));
 sg13g2_tiehi _1413__142 (.L_HI(net199));
 sg13g2_tiehi _1412__143 (.L_HI(net200));
 sg13g2_tiehi _1411__144 (.L_HI(net201));
 sg13g2_tiehi _1410__145 (.L_HI(net202));
 sg13g2_tiehi _1409__146 (.L_HI(net203));
 sg13g2_tiehi _1408__147 (.L_HI(net204));
 sg13g2_tiehi _1590__148 (.L_HI(net205));
 sg13g2_tiehi _1407__149 (.L_HI(net206));
 sg13g2_tiehi _1566__150 (.L_HI(net207));
 sg13g2_tiehi _1406__151 (.L_HI(net208));
 sg13g2_tiehi _1578__152 (.L_HI(net209));
 sg13g2_tiehi _1405__153 (.L_HI(net210));
 sg13g2_tiehi _1565__154 (.L_HI(net211));
 sg13g2_tiehi _1404__155 (.L_HI(net212));
 sg13g2_tiehi _1589__156 (.L_HI(net213));
 sg13g2_tiehi _1564__157 (.L_HI(net214));
 sg13g2_tiehi _1467__158 (.L_HI(net215));
 sg13g2_tiehi _1577__159 (.L_HI(net216));
 sg13g2_tiehi _1563__160 (.L_HI(net217));
 sg13g2_tiehi _1593__161 (.L_HI(net218));
 sg13g2_tiehi _1562__162 (.L_HI(net219));
 sg13g2_tiehi _1576__163 (.L_HI(net220));
 sg13g2_tiehi _1561__164 (.L_HI(net221));
 sg13g2_tiehi _1544__165 (.L_HI(net222));
 sg13g2_tiehi _1551__166 (.L_HI(net223));
 sg13g2_tiehi _1552__167 (.L_HI(net224));
 sg13g2_tiehi _1553__168 (.L_HI(net225));
 sg13g2_tiehi _1554__169 (.L_HI(net226));
 sg13g2_tiehi _1555__170 (.L_HI(net227));
 sg13g2_tiehi _1556__171 (.L_HI(net228));
 sg13g2_tiehi _1557__172 (.L_HI(net229));
 sg13g2_tiehi _1558__173 (.L_HI(net230));
 sg13g2_tiehi _1560__174 (.L_HI(net231));
 sg13g2_tiehi _1588__175 (.L_HI(net232));
 sg13g2_tiehi _1550__176 (.L_HI(net233));
 sg13g2_tiehi _1575__177 (.L_HI(net234));
 sg13g2_tiehi _1549__178 (.L_HI(net235));
 sg13g2_tiehi _1594__179 (.L_HI(net236));
 sg13g2_tiehi _1548__180 (.L_HI(net237));
 sg13g2_tiehi _1574__181 (.L_HI(net238));
 sg13g2_tiehi _1547__182 (.L_HI(net239));
 sg13g2_tiehi _1582__183 (.L_HI(net240));
 sg13g2_tiehi _1546__184 (.L_HI(net241));
 sg13g2_tiehi _1545__185 (.L_HI(net242));
 sg13g2_tiehi _1543__186 (.L_HI(net243));
 sg13g2_tiehi _1542__187 (.L_HI(net244));
 sg13g2_tiehi _1541__188 (.L_HI(net245));
 sg13g2_tiehi _1540__189 (.L_HI(net246));
 sg13g2_tiehi _1539__190 (.L_HI(net247));
 sg13g2_tiehi _1538__191 (.L_HI(net248));
 sg13g2_tiehi _1537__192 (.L_HI(net249));
 sg13g2_tiehi _1536__193 (.L_HI(net250));
 sg13g2_tiehi _1535__194 (.L_HI(net251));
 sg13g2_tiehi _1534__195 (.L_HI(net252));
 sg13g2_tiehi _1533__196 (.L_HI(net253));
 sg13g2_tiehi _1559__197 (.L_HI(net254));
 sg13g2_tiehi _1583__198 (.L_HI(net255));
 sg13g2_tiehi _1584__199 (.L_HI(net256));
 sg13g2_tiehi _1585__200 (.L_HI(net257));
 sg13g2_tiehi _1586__201 (.L_HI(net258));
 sg13g2_tiehi _1532__202 (.L_HI(net259));
 sg13g2_tiehi _1531__203 (.L_HI(net260));
 sg13g2_tiehi _1530__204 (.L_HI(net261));
 sg13g2_tiehi _1529__205 (.L_HI(net262));
 sg13g2_tiehi _1528__206 (.L_HI(net263));
 sg13g2_tiehi _1527__207 (.L_HI(net264));
 sg13g2_tiehi tt_um_MichaelBell_photo_frame_208 (.L_HI(net265));
 sg13g2_tiehi tt_um_MichaelBell_photo_frame_209 (.L_HI(net266));
 sg13g2_inv_1 _0805__1 (.Y(net267),
    .A(clknet_1_0__leaf_clk));
 sg13g2_tielo tt_um_MichaelBell_photo_frame_15 (.L_LO(net15));
 sg13g2_tiehi _1526__16 (.L_HI(net16));
 sg13g2_buf_1 _1791_ (.A(net172),
    .X(uio_oe[0]));
 sg13g2_buf_1 _1792_ (.A(net172),
    .X(uio_oe[6]));
 sg13g2_buf_1 _1793_ (.A(net172),
    .X(uio_oe[7]));
 sg13g2_buf_1 _1794_ (.A(\i_qpsi.spi_select ),
    .X(uio_out[0]));
 sg13g2_buf_1 _1795_ (.A(vsync_r),
    .X(uo_out[3]));
 sg13g2_buf_1 _1796_ (.A(hsync_r),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout116 (.A(net118),
    .X(net116));
 sg13g2_buf_1 fanout117 (.A(net118),
    .X(net117));
 sg13g2_buf_8 fanout118 (.A(_0494_),
    .X(net118));
 sg13g2_buf_8 fanout119 (.A(net120),
    .X(net119));
 sg13g2_buf_8 fanout120 (.A(_0370_),
    .X(net120));
 sg13g2_buf_8 fanout121 (.A(net122),
    .X(net121));
 sg13g2_buf_1 fanout122 (.A(net123),
    .X(net122));
 sg13g2_buf_8 fanout123 (.A(_0496_),
    .X(net123));
 sg13g2_buf_8 fanout124 (.A(net128),
    .X(net124));
 sg13g2_buf_8 fanout125 (.A(net128),
    .X(net125));
 sg13g2_buf_8 fanout126 (.A(net127),
    .X(net126));
 sg13g2_buf_8 fanout127 (.A(net128),
    .X(net127));
 sg13g2_buf_8 fanout128 (.A(_0366_),
    .X(net128));
 sg13g2_buf_8 fanout129 (.A(_0204_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_0204_),
    .X(net130));
 sg13g2_buf_8 fanout131 (.A(net132),
    .X(net131));
 sg13g2_buf_8 fanout132 (.A(_0283_),
    .X(net132));
 sg13g2_buf_8 fanout133 (.A(net134),
    .X(net133));
 sg13g2_buf_8 fanout134 (.A(net137),
    .X(net134));
 sg13g2_buf_8 fanout135 (.A(net136),
    .X(net135));
 sg13g2_buf_8 fanout136 (.A(net137),
    .X(net136));
 sg13g2_buf_8 fanout137 (.A(_0260_),
    .X(net137));
 sg13g2_buf_8 fanout138 (.A(net139),
    .X(net138));
 sg13g2_buf_8 fanout139 (.A(net140),
    .X(net139));
 sg13g2_buf_1 fanout140 (.A(_0189_),
    .X(net140));
 sg13g2_buf_8 fanout141 (.A(net143),
    .X(net141));
 sg13g2_buf_1 fanout142 (.A(net143),
    .X(net142));
 sg13g2_buf_8 fanout143 (.A(net144),
    .X(net143));
 sg13g2_buf_8 fanout144 (.A(net147),
    .X(net144));
 sg13g2_buf_8 fanout145 (.A(net146),
    .X(net145));
 sg13g2_buf_8 fanout146 (.A(net147),
    .X(net146));
 sg13g2_buf_8 fanout147 (.A(_0471_),
    .X(net147));
 sg13g2_buf_8 fanout148 (.A(net149),
    .X(net148));
 sg13g2_buf_8 fanout149 (.A(net150),
    .X(net149));
 sg13g2_buf_8 fanout150 (.A(_0471_),
    .X(net150));
 sg13g2_buf_8 fanout151 (.A(net152),
    .X(net151));
 sg13g2_buf_8 fanout152 (.A(net155),
    .X(net152));
 sg13g2_buf_8 fanout153 (.A(net154),
    .X(net153));
 sg13g2_buf_8 fanout154 (.A(net155),
    .X(net154));
 sg13g2_buf_8 fanout155 (.A(_0471_),
    .X(net155));
 sg13g2_buf_8 fanout156 (.A(net157),
    .X(net156));
 sg13g2_buf_8 fanout157 (.A(_0206_),
    .X(net157));
 sg13g2_buf_1 fanout158 (.A(_0206_),
    .X(net158));
 sg13g2_buf_8 fanout159 (.A(net558),
    .X(net159));
 sg13g2_buf_8 fanout160 (.A(net554),
    .X(net160));
 sg13g2_buf_8 fanout161 (.A(net559),
    .X(net161));
 sg13g2_buf_8 fanout162 (.A(\i_display.v_state[0] ),
    .X(net162));
 sg13g2_buf_8 fanout163 (.A(net164),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(\i_qpsi.valid ),
    .X(net164));
 sg13g2_buf_8 fanout165 (.A(net166),
    .X(net165));
 sg13g2_buf_8 fanout166 (.A(net167),
    .X(net166));
 sg13g2_buf_8 fanout167 (.A(_0194_),
    .X(net167));
 sg13g2_buf_8 fanout168 (.A(net169),
    .X(net168));
 sg13g2_buf_8 fanout169 (.A(_0193_),
    .X(net169));
 sg13g2_buf_8 fanout170 (.A(net171),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(ui_in[3]),
    .X(net171));
 sg13g2_buf_8 fanout172 (.A(net1),
    .X(net172));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[1]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[2]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[3]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[4]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[5]),
    .X(net13));
 sg13g2_tielo tt_um_MichaelBell_photo_frame_14 (.L_LO(net14));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(delaynet_0_clk));
 sg13g2_buf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_8 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_buf_8 clkbuf_5_0__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_0__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_1__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_1__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_2__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_2__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_3__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_3__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_4__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_4__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_5__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_5__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_6__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_6__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_7__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_7__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_8__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_8__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_9__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_9__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_10__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_10__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_11__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_12__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_12__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_13__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_13__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_14__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_14__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_15__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_15__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_16__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_16__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_17__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_17__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_18__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_18__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_19__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_20__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_20__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_21__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_21__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_22__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_22__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_23__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_23__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_24__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_24__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_25__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_26__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_26__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_27__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_27__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_28__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_28__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_29__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_29__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_30__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_30__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_31__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_31__leaf_clk_regs));
 sg13g2_buf_1 clkload0 (.A(clknet_5_1__leaf_clk_regs));
 sg13g2_buf_1 clkload1 (.A(clknet_5_4__leaf_clk_regs));
 sg13g2_buf_1 clkload2 (.A(clknet_5_7__leaf_clk_regs));
 sg13g2_buf_1 clkload3 (.A(clknet_5_8__leaf_clk_regs));
 sg13g2_buf_1 clkload4 (.A(clknet_5_10__leaf_clk_regs));
 sg13g2_buf_1 clkload5 (.A(clknet_5_13__leaf_clk_regs));
 sg13g2_buf_1 clkload6 (.A(clknet_5_14__leaf_clk_regs));
 sg13g2_buf_1 clkload7 (.A(clknet_5_17__leaf_clk_regs));
 sg13g2_buf_1 clkload8 (.A(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_1 clkload9 (.A(clknet_5_21__leaf_clk_regs));
 sg13g2_buf_1 clkload10 (.A(clknet_5_26__leaf_clk_regs));
 sg13g2_buf_1 clkload11 (.A(clknet_5_28__leaf_clk_regs));
 sg13g2_inv_1 clkload12 (.A(clknet_5_31__leaf_clk_regs));
 sg13g2_buf_8 delaybuf_0_clk (.A(delaynet_0_clk),
    .X(clknet_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\i_display.cfg_data_sync[0] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold2 (.A(\i_display.cfg_clk_sync[0] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold3 (.A(\i_qpsi.spi_miso_buf[4] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold4 (.A(\i_qpsi.spi_miso_buf[0] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold5 (.A(\i_qpsi.spi_miso_buf[2] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold6 (.A(\i_qpsi.spi_miso_buf[6] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold7 (.A(\i_qpsi.spi_miso_buf[3] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold8 (.A(\i_qpsi.spi_miso_buf[1] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold9 (.A(\i_qpsi.spi_miso_buf[5] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold10 (.A(\i_qpsi.spi_miso_buf[7] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold11 (.A(\i_display.cfg_clk_sync[1] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold12 (.A(\i_qpsi.addr[17] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0041_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold14 (.A(\i_display.cfg[68] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold15 (.A(hsync),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold16 (.A(\i_qpsi.data[6] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0061_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold18 (.A(\i_qpsi.addr[13] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0037_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold20 (.A(\i_qpsi.addr[18] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0042_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold22 (.A(\i_qpsi.addr[6] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0030_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold24 (.A(\i_qpsi.addr[5] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0029_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold26 (.A(\addr_in[0] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0144_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold28 (.A(\i_qpsi.addr[10] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0034_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold30 (.A(\i_qpsi.addr[16] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0040_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold32 (.A(\i_qpsi.addr[9] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0033_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold34 (.A(\addr_in[13] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0157_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold36 (.A(\i_qpsi.data[5] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0060_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold38 (.A(\i_qpsi.addr[15] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0039_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold40 (.A(\i_qpsi.addr[7] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0031_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold42 (.A(\i_qpsi.addr[19] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0043_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold44 (.A(\i_qpsi.addr[11] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0035_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold46 (.A(\i_qpsi.data[7] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0062_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold48 (.A(\i_qpsi.addr[12] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0036_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold50 (.A(\i_display.cfg[67] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold51 (.A(\i_display.vsync ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold52 (.A(\addr_in[23] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0047_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold54 (.A(\i_qpsi.addr[14] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0038_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold56 (.A(\addr_in[22] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0046_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold58 (.A(\i_display.cfg[38] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0101_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold60 (.A(\i_qpsi.addr[2] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0490_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold62 (.A(\i_qpsi.addr[0] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold63 (.A(\i_qpsi.data[4] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0059_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold65 (.A(\addr_in[14] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0580_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0158_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold68 (.A(\i_qpsi.addr[3] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0491_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold70 (.A(\i_display.cfg[53] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0116_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold72 (.A(\i_display.cfg[1] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0064_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold74 (.A(\i_qpsi.addr[1] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0489_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold76 (.A(\i_display.cfg[32] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0095_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold78 (.A(\i_display.cfg[54] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold79 (.A(\i_display.cfg[30] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0093_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold81 (.A(\i_qpsi.data[0] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0055_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold83 (.A(\addr_in[21] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0588_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0165_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold86 (.A(\i_qpsi.addr[21] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold87 (.A(\i_qpsi.data[3] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0058_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold89 (.A(\i_display.cfg[33] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0004_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold91 (.A(\i_display.cfg[66] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0168_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold93 (.A(\i_qpsi.data[2] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0352_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold95 (.A(\addr_in[8] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0032_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold97 (.A(\addr_in[4] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0028_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold99 (.A(\i_display.cfg[5] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0068_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold101 (.A(uo_out[6]),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0341_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0342_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold104 (.A(\i_display.v_count[7] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0288_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0012_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold107 (.A(\addr_in[20] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0044_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold109 (.A(\i_qpsi.data[1] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0056_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold111 (.A(\i_display.cfg[36] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0100_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold113 (.A(\i_display.cfg[35] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold114 (.A(\i_qpsi.spi_miso_buf[10] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold115 (.A(\i_qpsi.spi_data_oe[0] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0487_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold117 (.A(\i_display.cfg[28] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0092_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold119 (.A(\i_display.cfg[65] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0592_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0167_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold122 (.A(\i_display.cfg[34] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0005_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold124 (.A(uo_out[1]),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0347_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0348_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold127 (.A(\i_display.h_count[3] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0229_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0230_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold130 (.A(\i_display.cfg[31] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold131 (.A(\i_display.v_count[10] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0301_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold133 (.A(\i_display.cfg[3] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0067_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold135 (.A(\i_display.cfg[0] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0016_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold137 (.A(uo_out[4]),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0349_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0350_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0026_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold141 (.A(\i_display.cfg[12] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0076_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold143 (.A(\i_display.cfg[37] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0008_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold145 (.A(uo_out[5]),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0345_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0346_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0024_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold149 (.A(\i_display.cfg[22] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0085_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold151 (.A(\i_display.v_count[4] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0020_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold153 (.A(\i_display.cfg[74] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0137_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold155 (.A(uo_out[2]),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0343_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0344_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold158 (.A(\i_display.cfg[11] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold159 (.A(\i_display.cfg[14] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0078_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold161 (.A(\i_display.cfg[23] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold162 (.A(\i_display.cfg[26] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0090_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold164 (.A(\i_display.cfg[17] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0080_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold166 (.A(\i_display.cfg[8] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0072_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold168 (.A(\i_display.cfg[39] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold169 (.A(\i_display.cfg[13] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold170 (.A(\i_display.cfg[55] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold171 (.A(\i_display.cfg[51] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0115_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold173 (.A(\i_display.cfg[7] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold174 (.A(\i_display.cfg[6] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold175 (.A(\i_display.cfg_data_sync[1] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold176 (.A(\i_qpsi.bits_remaining[2] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0448_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0051_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold179 (.A(\i_display.h_count[7] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0253_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold181 (.A(\i_display.cfg[44] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0107_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold183 (.A(\i_display.cfg[70] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0134_),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold185 (.A(\i_display.cfg[19] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0082_),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold187 (.A(\i_display.cfg[27] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold188 (.A(\i_display.cfg[25] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0088_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold190 (.A(\i_display.cfg[69] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold191 (.A(\i_display.cfg[10] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold192 (.A(\i_display.cfg[50] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0113_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold194 (.A(\i_display.cfg[29] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0000_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold196 (.A(\i_display.cfg[45] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold197 (.A(\i_display.cfg[20] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0084_),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold199 (.A(\i_display.cfg[24] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold200 (.A(\i_display.cfg[48] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0111_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold202 (.A(\i_display.cfg[16] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0079_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold204 (.A(\i_display.cfg[46] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold205 (.A(\i_display.cfg[49] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold206 (.A(\i_display.v_count[6] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold207 (.A(\i_qpsi.fsm_state[2] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0457_),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold209 (.A(\addr_in[16] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0582_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold211 (.A(\i_display.cfg[72] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0136_),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold213 (.A(\i_display.cfg[47] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold214 (.A(\i_display.cfg[42] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0105_),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold216 (.A(\i_display.cfg[2] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold217 (.A(\i_display.cfg[64] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold218 (.A(\i_display.cfg[63] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0126_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold220 (.A(\i_display.cfg[59] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0123_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold222 (.A(\i_display.cfg[43] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold223 (.A(\i_display.cfg[18] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold224 (.A(\i_display.cfg[58] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0221_),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0223_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0225_),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold228 (.A(\i_display.cfg[57] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold229 (.A(\i_display.cfg[41] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0104_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold231 (.A(\i_display.cfg[40] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold232 (.A(\i_display.cfg[62] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0125_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold234 (.A(\i_display.cfg[9] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold235 (.A(\i_display.cfg[56] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold236 (.A(\i_display.h_count[1] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0216_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold238 (.A(\addr_in[19] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0541_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold240 (.A(\i_display.cfg[71] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold241 (.A(\i_qpsi.fsm_state[1] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0456_),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold243 (.A(\addr_in[11] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0576_),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0155_),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold246 (.A(\i_display.v_count[2] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0018_),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold248 (.A(\i_display.h_count[6] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0006_),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold250 (.A(\addr_in[1] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold251 (.A(\i_qpsi.spi_clk ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0430_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold253 (.A(\i_display.cfg[61] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0124_),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold255 (.A(\i_display.v_count[5] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0021_),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold257 (.A(\addr_in[18] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0541_),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold259 (.A(\addr_in[12] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0578_),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold261 (.A(\i_display.v_state[1] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0596_),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold263 (.A(\addr_in[17] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0540_),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold265 (.A(\i_display.v_count[1] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0017_),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold267 (.A(\addr_in[6] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0150_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold269 (.A(\addr_in[15] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold270 (.A(\addr_in[7] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0523_),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold272 (.A(\addr_in[10] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold273 (.A(\addr_in[3] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold274 (.A(_0509_),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold275 (.A(\addr_in[2] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold276 (.A(\i_display.v_count[3] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0019_),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold278 (.A(\i_qpsi.bits_remaining[0] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold279 (.A(_0049_),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold280 (.A(\addr_in[5] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold281 (.A(\addr_in[9] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold282 (.A(\i_display.v_count[8] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0292_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold284 (.A(\i_display.v_state[0] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0595_),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold286 (.A(\i_display.v_count[9] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold287 (.A(\i_display.h_state[0] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0597_),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold289 (.A(\i_qpsi.fsm_state[0] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold290 (.A(\i_qpsi.bits_remaining[1] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold291 (.A(\i_display.h_state[1] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold292 (.A(\i_display.v_state[1] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold293 (.A(\i_display.v_count[5] ),
    .X(net560));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_4 FILLER_0_56 ();
 sg13g2_decap_4 FILLER_0_97 ();
 sg13g2_decap_4 FILLER_0_111 ();
 sg13g2_fill_1 FILLER_0_115 ();
 sg13g2_decap_8 FILLER_0_120 ();
 sg13g2_fill_1 FILLER_0_127 ();
 sg13g2_decap_4 FILLER_0_138 ();
 sg13g2_decap_4 FILLER_0_146 ();
 sg13g2_fill_2 FILLER_0_150 ();
 sg13g2_decap_4 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_188 ();
 sg13g2_decap_4 FILLER_0_195 ();
 sg13g2_fill_1 FILLER_0_199 ();
 sg13g2_decap_4 FILLER_0_227 ();
 sg13g2_fill_1 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_276 ();
 sg13g2_decap_8 FILLER_0_283 ();
 sg13g2_decap_8 FILLER_0_290 ();
 sg13g2_decap_8 FILLER_0_297 ();
 sg13g2_decap_8 FILLER_0_304 ();
 sg13g2_decap_8 FILLER_0_311 ();
 sg13g2_decap_8 FILLER_0_318 ();
 sg13g2_decap_8 FILLER_0_325 ();
 sg13g2_decap_8 FILLER_0_332 ();
 sg13g2_decap_8 FILLER_0_339 ();
 sg13g2_decap_8 FILLER_0_346 ();
 sg13g2_decap_8 FILLER_0_353 ();
 sg13g2_decap_8 FILLER_0_360 ();
 sg13g2_decap_8 FILLER_0_367 ();
 sg13g2_decap_8 FILLER_0_374 ();
 sg13g2_decap_8 FILLER_0_381 ();
 sg13g2_decap_8 FILLER_0_388 ();
 sg13g2_decap_8 FILLER_0_395 ();
 sg13g2_decap_8 FILLER_0_402 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_4 FILLER_1_49 ();
 sg13g2_fill_2 FILLER_1_53 ();
 sg13g2_fill_1 FILLER_1_82 ();
 sg13g2_fill_2 FILLER_1_216 ();
 sg13g2_fill_2 FILLER_1_246 ();
 sg13g2_decap_4 FILLER_1_285 ();
 sg13g2_fill_1 FILLER_1_289 ();
 sg13g2_fill_1 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_304 ();
 sg13g2_decap_8 FILLER_1_311 ();
 sg13g2_decap_8 FILLER_1_318 ();
 sg13g2_decap_8 FILLER_1_325 ();
 sg13g2_decap_8 FILLER_1_332 ();
 sg13g2_decap_8 FILLER_1_339 ();
 sg13g2_decap_8 FILLER_1_346 ();
 sg13g2_decap_8 FILLER_1_353 ();
 sg13g2_decap_8 FILLER_1_360 ();
 sg13g2_decap_8 FILLER_1_367 ();
 sg13g2_decap_8 FILLER_1_374 ();
 sg13g2_decap_8 FILLER_1_381 ();
 sg13g2_decap_8 FILLER_1_388 ();
 sg13g2_decap_8 FILLER_1_395 ();
 sg13g2_decap_8 FILLER_1_402 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_fill_1 FILLER_2_49 ();
 sg13g2_fill_2 FILLER_2_58 ();
 sg13g2_fill_1 FILLER_2_60 ();
 sg13g2_fill_1 FILLER_2_83 ();
 sg13g2_fill_2 FILLER_2_97 ();
 sg13g2_fill_2 FILLER_2_118 ();
 sg13g2_fill_1 FILLER_2_120 ();
 sg13g2_decap_8 FILLER_2_130 ();
 sg13g2_decap_8 FILLER_2_137 ();
 sg13g2_fill_2 FILLER_2_157 ();
 sg13g2_fill_2 FILLER_2_253 ();
 sg13g2_fill_1 FILLER_2_255 ();
 sg13g2_fill_2 FILLER_2_283 ();
 sg13g2_decap_8 FILLER_2_312 ();
 sg13g2_decap_8 FILLER_2_319 ();
 sg13g2_decap_8 FILLER_2_326 ();
 sg13g2_decap_8 FILLER_2_333 ();
 sg13g2_decap_8 FILLER_2_340 ();
 sg13g2_decap_8 FILLER_2_347 ();
 sg13g2_decap_8 FILLER_2_354 ();
 sg13g2_decap_8 FILLER_2_361 ();
 sg13g2_decap_8 FILLER_2_368 ();
 sg13g2_decap_8 FILLER_2_375 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_4 FILLER_2_403 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_fill_2 FILLER_3_28 ();
 sg13g2_fill_1 FILLER_3_30 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_4 FILLER_3_42 ();
 sg13g2_fill_1 FILLER_3_46 ();
 sg13g2_fill_1 FILLER_3_139 ();
 sg13g2_fill_2 FILLER_3_168 ();
 sg13g2_fill_1 FILLER_3_170 ();
 sg13g2_decap_4 FILLER_3_194 ();
 sg13g2_fill_1 FILLER_3_198 ();
 sg13g2_fill_2 FILLER_3_240 ();
 sg13g2_fill_2 FILLER_3_254 ();
 sg13g2_fill_1 FILLER_3_256 ();
 sg13g2_fill_1 FILLER_3_266 ();
 sg13g2_fill_2 FILLER_3_285 ();
 sg13g2_fill_1 FILLER_3_296 ();
 sg13g2_fill_2 FILLER_3_302 ();
 sg13g2_fill_2 FILLER_3_339 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_4 FILLER_4_21 ();
 sg13g2_fill_1 FILLER_4_25 ();
 sg13g2_fill_1 FILLER_4_53 ();
 sg13g2_fill_1 FILLER_4_72 ();
 sg13g2_fill_2 FILLER_4_83 ();
 sg13g2_fill_1 FILLER_4_108 ();
 sg13g2_decap_8 FILLER_4_122 ();
 sg13g2_fill_2 FILLER_4_129 ();
 sg13g2_fill_2 FILLER_4_156 ();
 sg13g2_fill_1 FILLER_4_158 ();
 sg13g2_fill_1 FILLER_4_189 ();
 sg13g2_fill_2 FILLER_4_233 ();
 sg13g2_fill_1 FILLER_4_235 ();
 sg13g2_fill_2 FILLER_4_268 ();
 sg13g2_fill_1 FILLER_4_270 ();
 sg13g2_fill_1 FILLER_4_325 ();
 sg13g2_decap_8 FILLER_4_358 ();
 sg13g2_decap_8 FILLER_4_365 ();
 sg13g2_decap_8 FILLER_4_372 ();
 sg13g2_decap_8 FILLER_4_379 ();
 sg13g2_decap_8 FILLER_4_386 ();
 sg13g2_decap_8 FILLER_4_393 ();
 sg13g2_decap_8 FILLER_4_400 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_4 FILLER_5_28 ();
 sg13g2_fill_2 FILLER_5_153 ();
 sg13g2_decap_8 FILLER_5_183 ();
 sg13g2_fill_1 FILLER_5_190 ();
 sg13g2_fill_2 FILLER_5_219 ();
 sg13g2_fill_1 FILLER_5_221 ();
 sg13g2_fill_2 FILLER_5_296 ();
 sg13g2_fill_1 FILLER_5_311 ();
 sg13g2_fill_1 FILLER_5_344 ();
 sg13g2_fill_2 FILLER_5_359 ();
 sg13g2_decap_8 FILLER_5_369 ();
 sg13g2_decap_8 FILLER_5_376 ();
 sg13g2_decap_8 FILLER_5_383 ();
 sg13g2_decap_8 FILLER_5_390 ();
 sg13g2_decap_8 FILLER_5_397 ();
 sg13g2_decap_4 FILLER_5_404 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_4 FILLER_6_14 ();
 sg13g2_fill_2 FILLER_6_18 ();
 sg13g2_decap_4 FILLER_6_24 ();
 sg13g2_fill_1 FILLER_6_28 ();
 sg13g2_fill_1 FILLER_6_111 ();
 sg13g2_fill_1 FILLER_6_121 ();
 sg13g2_fill_1 FILLER_6_131 ();
 sg13g2_fill_1 FILLER_6_157 ();
 sg13g2_decap_8 FILLER_6_199 ();
 sg13g2_fill_2 FILLER_6_206 ();
 sg13g2_fill_1 FILLER_6_208 ();
 sg13g2_fill_1 FILLER_6_264 ();
 sg13g2_fill_2 FILLER_6_291 ();
 sg13g2_fill_1 FILLER_6_369 ();
 sg13g2_fill_2 FILLER_6_374 ();
 sg13g2_decap_4 FILLER_6_398 ();
 sg13g2_fill_1 FILLER_6_402 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_fill_1 FILLER_7_14 ();
 sg13g2_fill_1 FILLER_7_107 ();
 sg13g2_fill_1 FILLER_7_131 ();
 sg13g2_fill_2 FILLER_7_149 ();
 sg13g2_fill_2 FILLER_7_170 ();
 sg13g2_fill_1 FILLER_7_172 ();
 sg13g2_fill_2 FILLER_7_229 ();
 sg13g2_fill_2 FILLER_7_272 ();
 sg13g2_fill_2 FILLER_7_323 ();
 sg13g2_fill_1 FILLER_7_354 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_fill_1 FILLER_8_35 ();
 sg13g2_fill_1 FILLER_8_58 ();
 sg13g2_fill_1 FILLER_8_68 ();
 sg13g2_fill_2 FILLER_8_94 ();
 sg13g2_fill_2 FILLER_8_102 ();
 sg13g2_fill_2 FILLER_8_118 ();
 sg13g2_decap_8 FILLER_8_148 ();
 sg13g2_fill_1 FILLER_8_183 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_fill_1 FILLER_8_210 ();
 sg13g2_fill_1 FILLER_8_239 ();
 sg13g2_fill_1 FILLER_8_295 ();
 sg13g2_fill_2 FILLER_8_369 ();
 sg13g2_fill_1 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_fill_1 FILLER_9_14 ();
 sg13g2_fill_2 FILLER_9_53 ();
 sg13g2_fill_1 FILLER_9_104 ();
 sg13g2_fill_1 FILLER_9_117 ();
 sg13g2_fill_2 FILLER_9_123 ();
 sg13g2_decap_4 FILLER_9_135 ();
 sg13g2_fill_1 FILLER_9_139 ();
 sg13g2_decap_8 FILLER_9_144 ();
 sg13g2_fill_1 FILLER_9_209 ();
 sg13g2_fill_2 FILLER_9_214 ();
 sg13g2_fill_2 FILLER_9_235 ();
 sg13g2_fill_2 FILLER_9_243 ();
 sg13g2_fill_1 FILLER_9_245 ();
 sg13g2_fill_1 FILLER_9_273 ();
 sg13g2_fill_2 FILLER_9_306 ();
 sg13g2_fill_1 FILLER_9_325 ();
 sg13g2_fill_1 FILLER_9_355 ();
 sg13g2_fill_2 FILLER_9_388 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_4 FILLER_10_14 ();
 sg13g2_fill_2 FILLER_10_18 ();
 sg13g2_fill_2 FILLER_10_24 ();
 sg13g2_fill_2 FILLER_10_73 ();
 sg13g2_fill_1 FILLER_10_88 ();
 sg13g2_decap_4 FILLER_10_134 ();
 sg13g2_fill_1 FILLER_10_138 ();
 sg13g2_fill_2 FILLER_10_149 ();
 sg13g2_decap_4 FILLER_10_177 ();
 sg13g2_decap_4 FILLER_10_191 ();
 sg13g2_fill_2 FILLER_10_233 ();
 sg13g2_fill_1 FILLER_10_235 ();
 sg13g2_fill_2 FILLER_10_244 ();
 sg13g2_fill_2 FILLER_10_339 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_4 FILLER_11_21 ();
 sg13g2_fill_1 FILLER_11_25 ();
 sg13g2_fill_1 FILLER_11_39 ();
 sg13g2_fill_1 FILLER_11_50 ();
 sg13g2_decap_4 FILLER_11_102 ();
 sg13g2_fill_1 FILLER_11_106 ();
 sg13g2_fill_1 FILLER_11_116 ();
 sg13g2_fill_2 FILLER_11_132 ();
 sg13g2_fill_1 FILLER_11_134 ();
 sg13g2_fill_2 FILLER_11_167 ();
 sg13g2_fill_1 FILLER_11_169 ();
 sg13g2_fill_2 FILLER_11_190 ();
 sg13g2_fill_1 FILLER_11_225 ();
 sg13g2_fill_1 FILLER_11_259 ();
 sg13g2_decap_4 FILLER_11_299 ();
 sg13g2_fill_1 FILLER_11_303 ();
 sg13g2_fill_2 FILLER_11_320 ();
 sg13g2_fill_1 FILLER_11_322 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_fill_2 FILLER_12_21 ();
 sg13g2_fill_1 FILLER_12_23 ();
 sg13g2_fill_1 FILLER_12_88 ();
 sg13g2_fill_1 FILLER_12_114 ();
 sg13g2_fill_2 FILLER_12_135 ();
 sg13g2_fill_1 FILLER_12_137 ();
 sg13g2_fill_1 FILLER_12_148 ();
 sg13g2_decap_4 FILLER_12_185 ();
 sg13g2_fill_2 FILLER_12_206 ();
 sg13g2_fill_2 FILLER_12_233 ();
 sg13g2_fill_2 FILLER_12_322 ();
 sg13g2_fill_1 FILLER_12_324 ();
 sg13g2_fill_1 FILLER_12_336 ();
 sg13g2_fill_1 FILLER_12_351 ();
 sg13g2_fill_2 FILLER_12_379 ();
 sg13g2_fill_1 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_4 FILLER_13_28 ();
 sg13g2_fill_1 FILLER_13_32 ();
 sg13g2_decap_4 FILLER_13_42 ();
 sg13g2_fill_2 FILLER_13_91 ();
 sg13g2_decap_4 FILLER_13_117 ();
 sg13g2_fill_1 FILLER_13_121 ();
 sg13g2_fill_2 FILLER_13_137 ();
 sg13g2_fill_1 FILLER_13_139 ();
 sg13g2_fill_2 FILLER_13_152 ();
 sg13g2_fill_1 FILLER_13_181 ();
 sg13g2_fill_2 FILLER_13_191 ();
 sg13g2_fill_1 FILLER_13_193 ();
 sg13g2_fill_1 FILLER_13_217 ();
 sg13g2_fill_2 FILLER_13_228 ();
 sg13g2_decap_4 FILLER_13_238 ();
 sg13g2_fill_2 FILLER_13_264 ();
 sg13g2_fill_1 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_277 ();
 sg13g2_fill_2 FILLER_13_336 ();
 sg13g2_fill_1 FILLER_13_351 ();
 sg13g2_fill_1 FILLER_13_365 ();
 sg13g2_fill_2 FILLER_13_375 ();
 sg13g2_fill_1 FILLER_13_377 ();
 sg13g2_fill_1 FILLER_13_391 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_4 FILLER_14_42 ();
 sg13g2_fill_1 FILLER_14_46 ();
 sg13g2_decap_8 FILLER_14_52 ();
 sg13g2_fill_2 FILLER_14_59 ();
 sg13g2_fill_2 FILLER_14_89 ();
 sg13g2_fill_2 FILLER_14_128 ();
 sg13g2_fill_1 FILLER_14_130 ();
 sg13g2_fill_2 FILLER_14_166 ();
 sg13g2_fill_2 FILLER_14_205 ();
 sg13g2_fill_1 FILLER_14_234 ();
 sg13g2_decap_4 FILLER_14_272 ();
 sg13g2_fill_1 FILLER_14_276 ();
 sg13g2_fill_1 FILLER_14_296 ();
 sg13g2_fill_2 FILLER_14_341 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_fill_2 FILLER_15_28 ();
 sg13g2_decap_4 FILLER_15_66 ();
 sg13g2_fill_1 FILLER_15_70 ();
 sg13g2_fill_1 FILLER_15_88 ();
 sg13g2_decap_4 FILLER_15_177 ();
 sg13g2_decap_4 FILLER_15_185 ();
 sg13g2_fill_2 FILLER_15_202 ();
 sg13g2_fill_2 FILLER_15_221 ();
 sg13g2_fill_2 FILLER_15_236 ();
 sg13g2_fill_2 FILLER_15_286 ();
 sg13g2_fill_2 FILLER_15_337 ();
 sg13g2_fill_2 FILLER_15_348 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_fill_2 FILLER_16_14 ();
 sg13g2_decap_4 FILLER_16_20 ();
 sg13g2_fill_2 FILLER_16_24 ();
 sg13g2_fill_1 FILLER_16_52 ();
 sg13g2_fill_1 FILLER_16_75 ();
 sg13g2_fill_1 FILLER_16_81 ();
 sg13g2_decap_8 FILLER_16_122 ();
 sg13g2_fill_1 FILLER_16_134 ();
 sg13g2_fill_2 FILLER_16_141 ();
 sg13g2_fill_1 FILLER_16_143 ();
 sg13g2_decap_8 FILLER_16_158 ();
 sg13g2_fill_1 FILLER_16_165 ();
 sg13g2_decap_4 FILLER_16_231 ();
 sg13g2_fill_2 FILLER_16_282 ();
 sg13g2_fill_1 FILLER_16_298 ();
 sg13g2_fill_2 FILLER_16_316 ();
 sg13g2_fill_2 FILLER_16_332 ();
 sg13g2_fill_1 FILLER_16_334 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_70 ();
 sg13g2_fill_2 FILLER_17_87 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_fill_1 FILLER_17_132 ();
 sg13g2_fill_2 FILLER_17_138 ();
 sg13g2_fill_1 FILLER_17_140 ();
 sg13g2_decap_4 FILLER_17_145 ();
 sg13g2_decap_8 FILLER_17_176 ();
 sg13g2_decap_4 FILLER_17_183 ();
 sg13g2_fill_2 FILLER_17_187 ();
 sg13g2_decap_8 FILLER_17_193 ();
 sg13g2_decap_8 FILLER_17_214 ();
 sg13g2_fill_1 FILLER_17_221 ();
 sg13g2_decap_4 FILLER_17_255 ();
 sg13g2_fill_2 FILLER_17_259 ();
 sg13g2_fill_2 FILLER_17_288 ();
 sg13g2_fill_1 FILLER_17_290 ();
 sg13g2_fill_2 FILLER_17_360 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_50 ();
 sg13g2_fill_2 FILLER_18_74 ();
 sg13g2_fill_2 FILLER_18_102 ();
 sg13g2_fill_1 FILLER_18_104 ();
 sg13g2_fill_1 FILLER_18_113 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_fill_2 FILLER_18_140 ();
 sg13g2_fill_1 FILLER_18_142 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_158 ();
 sg13g2_fill_1 FILLER_18_165 ();
 sg13g2_fill_2 FILLER_18_170 ();
 sg13g2_fill_2 FILLER_18_227 ();
 sg13g2_fill_2 FILLER_18_273 ();
 sg13g2_fill_1 FILLER_18_275 ();
 sg13g2_fill_2 FILLER_18_293 ();
 sg13g2_fill_1 FILLER_18_308 ();
 sg13g2_fill_2 FILLER_18_319 ();
 sg13g2_fill_1 FILLER_18_321 ();
 sg13g2_fill_1 FILLER_18_344 ();
 sg13g2_fill_2 FILLER_18_358 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_fill_1 FILLER_19_30 ();
 sg13g2_fill_2 FILLER_19_40 ();
 sg13g2_fill_1 FILLER_19_85 ();
 sg13g2_fill_2 FILLER_19_99 ();
 sg13g2_decap_4 FILLER_19_124 ();
 sg13g2_fill_2 FILLER_19_128 ();
 sg13g2_fill_2 FILLER_19_166 ();
 sg13g2_decap_4 FILLER_19_189 ();
 sg13g2_fill_1 FILLER_19_193 ();
 sg13g2_decap_8 FILLER_19_219 ();
 sg13g2_fill_1 FILLER_19_226 ();
 sg13g2_decap_4 FILLER_19_235 ();
 sg13g2_fill_2 FILLER_19_244 ();
 sg13g2_fill_1 FILLER_19_246 ();
 sg13g2_fill_1 FILLER_19_276 ();
 sg13g2_fill_2 FILLER_19_308 ();
 sg13g2_fill_2 FILLER_19_328 ();
 sg13g2_fill_1 FILLER_19_330 ();
 sg13g2_fill_1 FILLER_19_371 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_65 ();
 sg13g2_fill_1 FILLER_20_67 ();
 sg13g2_fill_2 FILLER_20_77 ();
 sg13g2_fill_1 FILLER_20_88 ();
 sg13g2_fill_1 FILLER_20_124 ();
 sg13g2_decap_8 FILLER_20_146 ();
 sg13g2_fill_1 FILLER_20_153 ();
 sg13g2_decap_8 FILLER_20_184 ();
 sg13g2_fill_2 FILLER_20_191 ();
 sg13g2_fill_1 FILLER_20_205 ();
 sg13g2_fill_2 FILLER_20_219 ();
 sg13g2_fill_1 FILLER_20_221 ();
 sg13g2_fill_2 FILLER_20_227 ();
 sg13g2_fill_2 FILLER_20_239 ();
 sg13g2_fill_2 FILLER_20_246 ();
 sg13g2_fill_1 FILLER_20_248 ();
 sg13g2_fill_2 FILLER_20_277 ();
 sg13g2_fill_1 FILLER_20_322 ();
 sg13g2_fill_2 FILLER_20_367 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_2 ();
 sg13g2_fill_2 FILLER_21_28 ();
 sg13g2_fill_1 FILLER_21_30 ();
 sg13g2_fill_1 FILLER_21_41 ();
 sg13g2_fill_1 FILLER_21_57 ();
 sg13g2_fill_1 FILLER_21_103 ();
 sg13g2_decap_4 FILLER_21_116 ();
 sg13g2_fill_2 FILLER_21_120 ();
 sg13g2_fill_1 FILLER_21_143 ();
 sg13g2_fill_1 FILLER_21_154 ();
 sg13g2_fill_2 FILLER_21_168 ();
 sg13g2_fill_1 FILLER_21_174 ();
 sg13g2_decap_8 FILLER_21_179 ();
 sg13g2_fill_2 FILLER_21_186 ();
 sg13g2_fill_2 FILLER_21_201 ();
 sg13g2_decap_4 FILLER_21_230 ();
 sg13g2_fill_2 FILLER_21_234 ();
 sg13g2_fill_2 FILLER_21_253 ();
 sg13g2_fill_2 FILLER_21_259 ();
 sg13g2_fill_2 FILLER_21_356 ();
 sg13g2_fill_1 FILLER_21_358 ();
 sg13g2_fill_2 FILLER_21_369 ();
 sg13g2_fill_2 FILLER_22_31 ();
 sg13g2_fill_1 FILLER_22_42 ();
 sg13g2_fill_2 FILLER_22_52 ();
 sg13g2_fill_2 FILLER_22_67 ();
 sg13g2_fill_2 FILLER_22_74 ();
 sg13g2_fill_1 FILLER_22_76 ();
 sg13g2_fill_1 FILLER_22_81 ();
 sg13g2_fill_2 FILLER_22_90 ();
 sg13g2_fill_1 FILLER_22_102 ();
 sg13g2_decap_8 FILLER_22_108 ();
 sg13g2_fill_2 FILLER_22_142 ();
 sg13g2_fill_1 FILLER_22_144 ();
 sg13g2_decap_8 FILLER_22_149 ();
 sg13g2_fill_1 FILLER_22_156 ();
 sg13g2_fill_1 FILLER_22_189 ();
 sg13g2_fill_2 FILLER_22_261 ();
 sg13g2_fill_1 FILLER_22_263 ();
 sg13g2_fill_2 FILLER_22_277 ();
 sg13g2_fill_1 FILLER_22_279 ();
 sg13g2_fill_2 FILLER_22_294 ();
 sg13g2_fill_1 FILLER_22_338 ();
 sg13g2_fill_2 FILLER_22_356 ();
 sg13g2_fill_1 FILLER_22_358 ();
 sg13g2_fill_1 FILLER_23_31 ();
 sg13g2_fill_1 FILLER_23_83 ();
 sg13g2_fill_2 FILLER_23_124 ();
 sg13g2_fill_2 FILLER_23_200 ();
 sg13g2_fill_2 FILLER_23_242 ();
 sg13g2_fill_2 FILLER_23_276 ();
 sg13g2_fill_2 FILLER_23_321 ();
 sg13g2_fill_1 FILLER_23_323 ();
 sg13g2_fill_2 FILLER_23_375 ();
 sg13g2_fill_1 FILLER_23_381 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_50 ();
 sg13g2_fill_1 FILLER_24_57 ();
 sg13g2_fill_2 FILLER_24_120 ();
 sg13g2_fill_1 FILLER_24_140 ();
 sg13g2_fill_2 FILLER_24_150 ();
 sg13g2_fill_2 FILLER_24_189 ();
 sg13g2_fill_1 FILLER_24_191 ();
 sg13g2_fill_2 FILLER_24_205 ();
 sg13g2_fill_1 FILLER_24_207 ();
 sg13g2_fill_1 FILLER_24_314 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_fill_1 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_32 ();
 sg13g2_fill_1 FILLER_25_78 ();
 sg13g2_fill_2 FILLER_25_156 ();
 sg13g2_fill_1 FILLER_25_158 ();
 sg13g2_fill_2 FILLER_25_162 ();
 sg13g2_decap_8 FILLER_25_172 ();
 sg13g2_fill_2 FILLER_25_179 ();
 sg13g2_fill_1 FILLER_25_181 ();
 sg13g2_fill_1 FILLER_25_188 ();
 sg13g2_fill_1 FILLER_25_220 ();
 sg13g2_fill_2 FILLER_25_240 ();
 sg13g2_fill_1 FILLER_25_242 ();
 sg13g2_fill_2 FILLER_25_296 ();
 sg13g2_fill_2 FILLER_25_354 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_33 ();
 sg13g2_fill_1 FILLER_26_123 ();
 sg13g2_fill_2 FILLER_26_146 ();
 sg13g2_fill_1 FILLER_26_148 ();
 sg13g2_fill_2 FILLER_26_160 ();
 sg13g2_fill_1 FILLER_26_193 ();
 sg13g2_fill_2 FILLER_26_247 ();
 sg13g2_fill_1 FILLER_26_249 ();
 sg13g2_fill_2 FILLER_26_296 ();
 sg13g2_fill_2 FILLER_26_308 ();
 sg13g2_fill_1 FILLER_26_332 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_2 ();
 sg13g2_fill_2 FILLER_27_39 ();
 sg13g2_fill_2 FILLER_27_64 ();
 sg13g2_fill_2 FILLER_27_94 ();
 sg13g2_fill_2 FILLER_27_155 ();
 sg13g2_fill_1 FILLER_27_166 ();
 sg13g2_fill_1 FILLER_27_171 ();
 sg13g2_decap_4 FILLER_27_181 ();
 sg13g2_fill_1 FILLER_27_207 ();
 sg13g2_fill_2 FILLER_27_229 ();
 sg13g2_fill_2 FILLER_27_280 ();
 sg13g2_fill_1 FILLER_27_282 ();
 sg13g2_fill_2 FILLER_27_377 ();
 sg13g2_fill_1 FILLER_27_379 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_2 ();
 sg13g2_fill_2 FILLER_28_81 ();
 sg13g2_fill_1 FILLER_28_122 ();
 sg13g2_fill_2 FILLER_28_184 ();
 sg13g2_fill_1 FILLER_28_186 ();
 sg13g2_fill_1 FILLER_28_215 ();
 sg13g2_fill_1 FILLER_28_255 ();
 sg13g2_fill_2 FILLER_28_293 ();
 sg13g2_fill_1 FILLER_28_295 ();
 sg13g2_fill_2 FILLER_28_332 ();
 sg13g2_fill_1 FILLER_28_334 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_1 FILLER_29_57 ();
 sg13g2_fill_2 FILLER_29_76 ();
 sg13g2_fill_1 FILLER_29_78 ();
 sg13g2_fill_2 FILLER_29_114 ();
 sg13g2_fill_1 FILLER_29_116 ();
 sg13g2_fill_1 FILLER_29_175 ();
 sg13g2_fill_2 FILLER_29_201 ();
 sg13g2_fill_1 FILLER_29_216 ();
 sg13g2_fill_2 FILLER_29_258 ();
 sg13g2_fill_1 FILLER_29_272 ();
 sg13g2_fill_2 FILLER_29_314 ();
 sg13g2_fill_2 FILLER_29_374 ();
 sg13g2_fill_1 FILLER_29_381 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_2 ();
 sg13g2_fill_2 FILLER_30_44 ();
 sg13g2_fill_2 FILLER_30_55 ();
 sg13g2_fill_1 FILLER_30_71 ();
 sg13g2_fill_2 FILLER_30_104 ();
 sg13g2_fill_1 FILLER_30_106 ();
 sg13g2_fill_2 FILLER_30_120 ();
 sg13g2_fill_2 FILLER_30_186 ();
 sg13g2_fill_2 FILLER_30_224 ();
 sg13g2_fill_1 FILLER_30_226 ();
 sg13g2_fill_1 FILLER_30_237 ();
 sg13g2_fill_1 FILLER_30_266 ();
 sg13g2_fill_1 FILLER_30_363 ();
 sg13g2_fill_2 FILLER_31_34 ();
 sg13g2_fill_1 FILLER_31_36 ();
 sg13g2_fill_2 FILLER_31_77 ();
 sg13g2_fill_1 FILLER_31_79 ();
 sg13g2_fill_2 FILLER_31_110 ();
 sg13g2_fill_2 FILLER_31_160 ();
 sg13g2_fill_1 FILLER_31_162 ();
 sg13g2_fill_1 FILLER_31_171 ();
 sg13g2_fill_1 FILLER_31_204 ();
 sg13g2_fill_1 FILLER_31_215 ();
 sg13g2_fill_2 FILLER_31_234 ();
 sg13g2_fill_2 FILLER_31_257 ();
 sg13g2_fill_1 FILLER_31_313 ();
 sg13g2_fill_1 FILLER_31_337 ();
 sg13g2_fill_2 FILLER_31_365 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_2 ();
 sg13g2_fill_2 FILLER_32_45 ();
 sg13g2_fill_1 FILLER_32_57 ();
 sg13g2_fill_2 FILLER_32_68 ();
 sg13g2_fill_1 FILLER_32_235 ();
 sg13g2_fill_1 FILLER_32_268 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_fill_2 FILLER_33_73 ();
 sg13g2_fill_1 FILLER_33_75 ();
 sg13g2_fill_1 FILLER_33_115 ();
 sg13g2_fill_1 FILLER_33_133 ();
 sg13g2_fill_1 FILLER_33_178 ();
 sg13g2_fill_1 FILLER_33_192 ();
 sg13g2_fill_2 FILLER_33_263 ();
 sg13g2_fill_1 FILLER_33_269 ();
 sg13g2_fill_2 FILLER_33_275 ();
 sg13g2_fill_1 FILLER_33_277 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_fill_2 FILLER_34_41 ();
 sg13g2_fill_2 FILLER_34_97 ();
 sg13g2_fill_2 FILLER_34_113 ();
 sg13g2_fill_2 FILLER_34_155 ();
 sg13g2_fill_1 FILLER_34_157 ();
 sg13g2_fill_1 FILLER_34_203 ();
 sg13g2_fill_1 FILLER_34_236 ();
 sg13g2_fill_2 FILLER_34_245 ();
 sg13g2_fill_2 FILLER_34_257 ();
 sg13g2_fill_2 FILLER_34_374 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_2 ();
 sg13g2_fill_1 FILLER_35_51 ();
 sg13g2_fill_1 FILLER_35_84 ();
 sg13g2_fill_2 FILLER_35_126 ();
 sg13g2_fill_2 FILLER_35_147 ();
 sg13g2_fill_1 FILLER_35_149 ();
 sg13g2_fill_2 FILLER_35_228 ();
 sg13g2_fill_1 FILLER_35_230 ();
 sg13g2_fill_2 FILLER_35_253 ();
 sg13g2_fill_1 FILLER_35_255 ();
 sg13g2_fill_2 FILLER_35_398 ();
 sg13g2_fill_1 FILLER_36_79 ();
 sg13g2_fill_1 FILLER_36_107 ();
 sg13g2_fill_1 FILLER_36_118 ();
 sg13g2_fill_2 FILLER_36_155 ();
 sg13g2_fill_1 FILLER_36_157 ();
 sg13g2_fill_1 FILLER_36_171 ();
 sg13g2_fill_1 FILLER_36_231 ();
 sg13g2_fill_2 FILLER_36_246 ();
 sg13g2_fill_1 FILLER_36_248 ();
 sg13g2_fill_2 FILLER_36_271 ();
 sg13g2_fill_1 FILLER_36_317 ();
 sg13g2_fill_2 FILLER_36_374 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_39 ();
 sg13g2_fill_1 FILLER_37_62 ();
 sg13g2_fill_2 FILLER_37_122 ();
 sg13g2_fill_2 FILLER_37_128 ();
 sg13g2_fill_1 FILLER_37_130 ();
 sg13g2_fill_2 FILLER_37_135 ();
 sg13g2_fill_1 FILLER_37_137 ();
 sg13g2_fill_2 FILLER_37_198 ();
 sg13g2_fill_2 FILLER_37_239 ();
 sg13g2_fill_2 FILLER_37_299 ();
 sg13g2_fill_1 FILLER_37_301 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_114 ();
 sg13g2_fill_2 FILLER_38_169 ();
 sg13g2_fill_2 FILLER_38_217 ();
 sg13g2_fill_2 FILLER_38_263 ();
 sg13g2_fill_1 FILLER_38_313 ();
 sg13g2_fill_1 FILLER_38_323 ();
 sg13g2_fill_2 FILLER_38_333 ();
 sg13g2_fill_1 FILLER_38_335 ();
 sg13g2_fill_1 FILLER_38_345 ();
 assign uio_oe[4] = net14;
 assign uio_oe[5] = net15;
 assign uio_out[6] = net265;
 assign uio_out[7] = net266;
endmodule
