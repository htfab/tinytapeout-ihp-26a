module tt_um_dranoel06_SAP1 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire \cpu0.a_reg[0] ;
 wire \cpu0.a_reg[1] ;
 wire \cpu0.a_reg[2] ;
 wire \cpu0.a_reg[3] ;
 wire \cpu0.a_reg[4] ;
 wire \cpu0.a_reg[5] ;
 wire \cpu0.a_reg[6] ;
 wire \cpu0.a_reg[7] ;
 wire \cpu0.b_reg[0] ;
 wire \cpu0.b_reg[1] ;
 wire \cpu0.b_reg[2] ;
 wire \cpu0.b_reg[3] ;
 wire \cpu0.b_reg[4] ;
 wire \cpu0.b_reg[5] ;
 wire \cpu0.b_reg[6] ;
 wire \cpu0.b_reg[7] ;
 wire \cpu0.carry_flag ;
 wire \cpu0.ir[0] ;
 wire \cpu0.ir[1] ;
 wire \cpu0.ir[2] ;
 wire \cpu0.ir[3] ;
 wire \cpu0.ir[4] ;
 wire \cpu0.ir[5] ;
 wire \cpu0.ir[6] ;
 wire \cpu0.ir[7] ;
 wire \cpu0.mar[0] ;
 wire \cpu0.mar[1] ;
 wire \cpu0.mar[2] ;
 wire \cpu0.mar[3] ;
 wire \cpu0.pc[0] ;
 wire \cpu0.pc[1] ;
 wire \cpu0.pc[2] ;
 wire \cpu0.pc[3] ;
 wire \cpu0.ram[0][0] ;
 wire \cpu0.ram[0][1] ;
 wire \cpu0.ram[0][2] ;
 wire \cpu0.ram[0][3] ;
 wire \cpu0.ram[0][4] ;
 wire \cpu0.ram[0][5] ;
 wire \cpu0.ram[0][6] ;
 wire \cpu0.ram[0][7] ;
 wire \cpu0.ram[10][0] ;
 wire \cpu0.ram[10][1] ;
 wire \cpu0.ram[10][2] ;
 wire \cpu0.ram[10][3] ;
 wire \cpu0.ram[10][4] ;
 wire \cpu0.ram[10][5] ;
 wire \cpu0.ram[10][6] ;
 wire \cpu0.ram[10][7] ;
 wire \cpu0.ram[11][0] ;
 wire \cpu0.ram[11][1] ;
 wire \cpu0.ram[11][2] ;
 wire \cpu0.ram[11][3] ;
 wire \cpu0.ram[11][4] ;
 wire \cpu0.ram[11][5] ;
 wire \cpu0.ram[11][6] ;
 wire \cpu0.ram[11][7] ;
 wire \cpu0.ram[12][0] ;
 wire \cpu0.ram[12][1] ;
 wire \cpu0.ram[12][2] ;
 wire \cpu0.ram[12][3] ;
 wire \cpu0.ram[12][4] ;
 wire \cpu0.ram[12][5] ;
 wire \cpu0.ram[12][6] ;
 wire \cpu0.ram[12][7] ;
 wire \cpu0.ram[13][0] ;
 wire \cpu0.ram[13][1] ;
 wire \cpu0.ram[13][2] ;
 wire \cpu0.ram[13][3] ;
 wire \cpu0.ram[13][4] ;
 wire \cpu0.ram[13][5] ;
 wire \cpu0.ram[13][6] ;
 wire \cpu0.ram[13][7] ;
 wire \cpu0.ram[14][0] ;
 wire \cpu0.ram[14][1] ;
 wire \cpu0.ram[14][2] ;
 wire \cpu0.ram[14][3] ;
 wire \cpu0.ram[14][4] ;
 wire \cpu0.ram[14][5] ;
 wire \cpu0.ram[14][6] ;
 wire \cpu0.ram[14][7] ;
 wire \cpu0.ram[15][0] ;
 wire \cpu0.ram[15][1] ;
 wire \cpu0.ram[15][2] ;
 wire \cpu0.ram[15][3] ;
 wire \cpu0.ram[15][4] ;
 wire \cpu0.ram[15][5] ;
 wire \cpu0.ram[15][6] ;
 wire \cpu0.ram[15][7] ;
 wire \cpu0.ram[1][0] ;
 wire \cpu0.ram[1][1] ;
 wire \cpu0.ram[1][2] ;
 wire \cpu0.ram[1][3] ;
 wire \cpu0.ram[1][4] ;
 wire \cpu0.ram[1][5] ;
 wire \cpu0.ram[1][6] ;
 wire \cpu0.ram[1][7] ;
 wire \cpu0.ram[2][0] ;
 wire \cpu0.ram[2][1] ;
 wire \cpu0.ram[2][2] ;
 wire \cpu0.ram[2][3] ;
 wire \cpu0.ram[2][4] ;
 wire \cpu0.ram[2][5] ;
 wire \cpu0.ram[2][6] ;
 wire \cpu0.ram[2][7] ;
 wire \cpu0.ram[3][0] ;
 wire \cpu0.ram[3][1] ;
 wire \cpu0.ram[3][2] ;
 wire \cpu0.ram[3][3] ;
 wire \cpu0.ram[3][4] ;
 wire \cpu0.ram[3][5] ;
 wire \cpu0.ram[3][6] ;
 wire \cpu0.ram[3][7] ;
 wire \cpu0.ram[4][0] ;
 wire \cpu0.ram[4][1] ;
 wire \cpu0.ram[4][2] ;
 wire \cpu0.ram[4][3] ;
 wire \cpu0.ram[4][4] ;
 wire \cpu0.ram[4][5] ;
 wire \cpu0.ram[4][6] ;
 wire \cpu0.ram[4][7] ;
 wire \cpu0.ram[5][0] ;
 wire \cpu0.ram[5][1] ;
 wire \cpu0.ram[5][2] ;
 wire \cpu0.ram[5][3] ;
 wire \cpu0.ram[5][4] ;
 wire \cpu0.ram[5][5] ;
 wire \cpu0.ram[5][6] ;
 wire \cpu0.ram[5][7] ;
 wire \cpu0.ram[6][0] ;
 wire \cpu0.ram[6][1] ;
 wire \cpu0.ram[6][2] ;
 wire \cpu0.ram[6][3] ;
 wire \cpu0.ram[6][4] ;
 wire \cpu0.ram[6][5] ;
 wire \cpu0.ram[6][6] ;
 wire \cpu0.ram[6][7] ;
 wire \cpu0.ram[7][0] ;
 wire \cpu0.ram[7][1] ;
 wire \cpu0.ram[7][2] ;
 wire \cpu0.ram[7][3] ;
 wire \cpu0.ram[7][4] ;
 wire \cpu0.ram[7][5] ;
 wire \cpu0.ram[7][6] ;
 wire \cpu0.ram[7][7] ;
 wire \cpu0.ram[8][0] ;
 wire \cpu0.ram[8][1] ;
 wire \cpu0.ram[8][2] ;
 wire \cpu0.ram[8][3] ;
 wire \cpu0.ram[8][4] ;
 wire \cpu0.ram[8][5] ;
 wire \cpu0.ram[8][6] ;
 wire \cpu0.ram[8][7] ;
 wire \cpu0.ram[9][0] ;
 wire \cpu0.ram[9][1] ;
 wire \cpu0.ram[9][2] ;
 wire \cpu0.ram[9][3] ;
 wire \cpu0.ram[9][4] ;
 wire \cpu0.ram[9][5] ;
 wire \cpu0.ram[9][6] ;
 wire \cpu0.ram[9][7] ;
 wire \cpu0.step[0] ;
 wire \cpu0.step[1] ;
 wire \cpu0.step[2] ;
 wire \cpu0.zero_flag ;
 wire \uart0.bit_counter[0] ;
 wire \uart0.bit_counter[1] ;
 wire \uart0.bit_counter[2] ;
 wire \uart0.bit_counter[3] ;
 wire \uart0.tx ;
 wire \uart0.tx_en_prev ;
 wire \uart0.uart_state[0] ;
 wire \uart0.uart_state[1] ;
 wire \uart0.uart_state[2] ;
 wire \uart0.uart_state[3] ;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire clknet_0_clk;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;

 sg13g2_inv_1 _0804_ (.Y(_0191_),
    .A(net278));
 sg13g2_inv_1 _0805_ (.Y(_0192_),
    .A(net434));
 sg13g2_inv_1 _0806_ (.Y(_0193_),
    .A(net148));
 sg13g2_inv_1 _0807_ (.Y(_0194_),
    .A(\cpu0.ir[6] ));
 sg13g2_inv_1 _0808_ (.Y(_0195_),
    .A(\cpu0.ir[5] ));
 sg13g2_inv_1 _0809_ (.Y(_0196_),
    .A(\cpu0.ir[3] ));
 sg13g2_inv_1 _0810_ (.Y(_0197_),
    .A(\cpu0.ir[2] ));
 sg13g2_inv_1 _0811_ (.Y(_0198_),
    .A(\cpu0.a_reg[4] ));
 sg13g2_inv_1 _0812_ (.Y(_0199_),
    .A(net178));
 sg13g2_inv_1 _0813_ (.Y(_0200_),
    .A(\cpu0.step[2] ));
 sg13g2_inv_1 _0814_ (.Y(_0201_),
    .A(net487));
 sg13g2_inv_1 _0815_ (.Y(_0202_),
    .A(net455));
 sg13g2_inv_2 _0816_ (.Y(_0203_),
    .A(net157));
 sg13g2_inv_1 _0817_ (.Y(_0204_),
    .A(net153));
 sg13g2_inv_1 _0818_ (.Y(_0205_),
    .A(net289));
 sg13g2_inv_1 _0819_ (.Y(_0206_),
    .A(net288));
 sg13g2_inv_1 _0820_ (.Y(_0207_),
    .A(net291));
 sg13g2_inv_1 _0821_ (.Y(_0208_),
    .A(\cpu0.ram[14][2] ));
 sg13g2_inv_1 _0822_ (.Y(_0209_),
    .A(\cpu0.ram[4][3] ));
 sg13g2_inv_1 _0823_ (.Y(_0210_),
    .A(net290));
 sg13g2_inv_1 _0824_ (.Y(_0211_),
    .A(\cpu0.ram[13][6] ));
 sg13g2_inv_1 _0825_ (.Y(_0212_),
    .A(\cpu0.ram[15][7] ));
 sg13g2_nor2b_1 _0826_ (.A(net463),
    .B_N(\cpu0.step[0] ),
    .Y(_0213_));
 sg13g2_nand2_1 _0827_ (.Y(_0214_),
    .A(\cpu0.step[1] ),
    .B(\cpu0.step[0] ));
 sg13g2_nor2_2 _0828_ (.A(net463),
    .B(_0214_),
    .Y(_0215_));
 sg13g2_nor2_1 _0829_ (.A(net173),
    .B(\cpu0.step[2] ),
    .Y(_0216_));
 sg13g2_nand2_2 _0830_ (.Y(_0217_),
    .A(net177),
    .B(_0215_));
 sg13g2_nor2_1 _0831_ (.A(net148),
    .B(\cpu0.ir[6] ),
    .Y(_0218_));
 sg13g2_nand2_1 _0832_ (.Y(_0219_),
    .A(\cpu0.ir[5] ),
    .B(\cpu0.ir[4] ));
 sg13g2_or4_1 _0833_ (.A(net148),
    .B(\cpu0.ir[6] ),
    .C(_0217_),
    .D(_0219_),
    .X(_0220_));
 sg13g2_inv_2 _0834_ (.Y(_0185_),
    .A(net145));
 sg13g2_o21ai_1 _0835_ (.B1(\uart0.uart_state[0] ),
    .Y(_0221_),
    .A1(net276),
    .A2(net145));
 sg13g2_nand3b_1 _0836_ (.B(_0221_),
    .C(net178),
    .Y(_0006_),
    .A_N(net304));
 sg13g2_nand4_1 _0837_ (.B(net434),
    .C(\uart0.bit_counter[1] ),
    .A(_0191_),
    .Y(_0222_),
    .D(\uart0.bit_counter[0] ));
 sg13g2_a21oi_1 _0838_ (.A1(\uart0.uart_state[1] ),
    .A2(_0222_),
    .Y(_0223_),
    .B1(net292));
 sg13g2_nor2_1 _0839_ (.A(net174),
    .B(net293),
    .Y(_0007_));
 sg13g2_nor3_1 _0840_ (.A(_0202_),
    .B(net276),
    .C(net145),
    .Y(_0004_));
 sg13g2_nor3_1 _0841_ (.A(net174),
    .B(_0201_),
    .C(net435),
    .Y(_0005_));
 sg13g2_nor2b_2 _0842_ (.A(net148),
    .B_N(\cpu0.ir[6] ),
    .Y(_0224_));
 sg13g2_nor2b_2 _0843_ (.A(\cpu0.ir[5] ),
    .B_N(\cpu0.ir[4] ),
    .Y(_0225_));
 sg13g2_nor3_2 _0844_ (.A(\cpu0.step[1] ),
    .B(_0200_),
    .C(\cpu0.step[0] ),
    .Y(_0226_));
 sg13g2_nand4_1 _0845_ (.B(_0224_),
    .C(_0225_),
    .A(net177),
    .Y(_0227_),
    .D(_0226_));
 sg13g2_nand2b_2 _0846_ (.Y(_0228_),
    .B(_0227_),
    .A_N(net13));
 sg13g2_nor2_1 _0847_ (.A(net13),
    .B(_0227_),
    .Y(_0229_));
 sg13g2_mux2_1 _0848_ (.A0(net10),
    .A1(\cpu0.mar[1] ),
    .S(net143),
    .X(_0230_));
 sg13g2_nor2b_2 _0849_ (.A(_0230_),
    .B_N(_0228_),
    .Y(_0231_));
 sg13g2_nor2b_1 _0850_ (.A(net142),
    .B_N(net9),
    .Y(_0232_));
 sg13g2_a21oi_2 _0851_ (.B1(_0232_),
    .Y(_0233_),
    .A2(net143),
    .A1(\cpu0.mar[0] ));
 sg13g2_nand2b_2 _0852_ (.Y(_0234_),
    .B(_0231_),
    .A_N(_0233_));
 sg13g2_mux2_1 _0853_ (.A0(net11),
    .A1(\cpu0.mar[2] ),
    .S(net144),
    .X(_0235_));
 sg13g2_mux2_1 _0854_ (.A0(net12),
    .A1(\cpu0.mar[3] ),
    .S(net144),
    .X(_0236_));
 sg13g2_nand2b_1 _0855_ (.Y(_0237_),
    .B(_0235_),
    .A_N(_0236_));
 sg13g2_or2_1 _0856_ (.X(_0238_),
    .B(_0237_),
    .A(_0234_));
 sg13g2_nor2b_2 _0857_ (.A(net468),
    .B_N(\cpu0.step[0] ),
    .Y(_0239_));
 sg13g2_and2_1 _0858_ (.A(_0216_),
    .B(_0239_),
    .X(_0240_));
 sg13g2_nand2b_1 _0859_ (.Y(_0241_),
    .B(_0240_),
    .A_N(net477));
 sg13g2_nor2_1 _0860_ (.A(\cpu0.ir[5] ),
    .B(\cpu0.ir[4] ),
    .Y(_0242_));
 sg13g2_nor2b_1 _0861_ (.A(\cpu0.ir[6] ),
    .B_N(net148),
    .Y(_0243_));
 sg13g2_nand2_1 _0862_ (.Y(_0244_),
    .A(\cpu0.zero_flag ),
    .B(_0215_));
 sg13g2_nand2_1 _0863_ (.Y(_0245_),
    .A(_0242_),
    .B(_0244_));
 sg13g2_a22oi_1 _0864_ (.Y(_0246_),
    .B1(_0243_),
    .B2(_0245_),
    .A2(_0242_),
    .A1(_0224_));
 sg13g2_a21oi_1 _0865_ (.A1(\cpu0.carry_flag ),
    .A2(_0215_),
    .Y(_0247_),
    .B1(_0195_));
 sg13g2_nor3_1 _0866_ (.A(net448),
    .B(_0246_),
    .C(_0247_),
    .Y(_0248_));
 sg13g2_nand3b_1 _0867_ (.B(_0224_),
    .C(_0242_),
    .Y(_0249_),
    .A_N(_0215_));
 sg13g2_nor2_1 _0868_ (.A(\cpu0.ir[6] ),
    .B(_0219_),
    .Y(_0250_));
 sg13g2_or2_1 _0869_ (.X(_0251_),
    .B(_0242_),
    .A(\cpu0.ir[7] ));
 sg13g2_o21ai_1 _0870_ (.B1(_0249_),
    .Y(_0252_),
    .A1(_0250_),
    .A2(_0251_));
 sg13g2_inv_1 _0871_ (.Y(_0253_),
    .A(_0252_));
 sg13g2_nand2_1 _0872_ (.Y(_0254_),
    .A(_0225_),
    .B(_0243_));
 sg13g2_o21ai_1 _0873_ (.B1(_0254_),
    .Y(_0255_),
    .A1(_0250_),
    .A2(_0251_));
 sg13g2_nand2b_1 _0874_ (.Y(_0256_),
    .B(\cpu0.ir[5] ),
    .A_N(\cpu0.ir[4] ));
 sg13g2_nor3_1 _0875_ (.A(net148),
    .B(\cpu0.ir[6] ),
    .C(_0256_),
    .Y(_0257_));
 sg13g2_a22oi_1 _0876_ (.Y(_0258_),
    .B1(_0255_),
    .B2(_0215_),
    .A2(_0253_),
    .A1(_0248_));
 sg13g2_nor2_2 _0877_ (.A(net172),
    .B(_0258_),
    .Y(_0259_));
 sg13g2_nand2_1 _0878_ (.Y(_0260_),
    .A(net284),
    .B(_0259_));
 sg13g2_nor2b_2 _0879_ (.A(_0219_),
    .B_N(_0224_),
    .Y(_0261_));
 sg13g2_nor2_2 _0880_ (.A(_0257_),
    .B(_0261_),
    .Y(_0262_));
 sg13g2_a21oi_1 _0881_ (.A1(_0254_),
    .A2(_0262_),
    .Y(_0263_),
    .B1(net172));
 sg13g2_nand2_2 _0882_ (.Y(_0264_),
    .A(_0226_),
    .B(_0263_));
 sg13g2_inv_1 _0883_ (.Y(_0265_),
    .A(net141));
 sg13g2_nand4_1 _0884_ (.B(_0218_),
    .C(_0225_),
    .A(net177),
    .Y(_0266_),
    .D(_0226_));
 sg13g2_nor2b_2 _0885_ (.A(net485),
    .B_N(net468),
    .Y(_0267_));
 sg13g2_and2_1 _0886_ (.A(_0216_),
    .B(_0267_),
    .X(_0268_));
 sg13g2_nand2_2 _0887_ (.Y(_0269_),
    .A(_0216_),
    .B(_0267_));
 sg13g2_and3_2 _0888_ (.X(_0270_),
    .A(net141),
    .B(_0266_),
    .C(_0269_));
 sg13g2_nand3_1 _0889_ (.B(_0266_),
    .C(_0269_),
    .A(net141),
    .Y(_0271_));
 sg13g2_mux4_1 _0890_ (.S0(net163),
    .A0(\cpu0.ram[0][0] ),
    .A1(\cpu0.ram[1][0] ),
    .A2(\cpu0.ram[2][0] ),
    .A3(\cpu0.ram[3][0] ),
    .S1(net155),
    .X(_0272_));
 sg13g2_or2_1 _0891_ (.X(_0273_),
    .B(_0272_),
    .A(net152));
 sg13g2_mux4_1 _0892_ (.S0(net163),
    .A0(\cpu0.ram[4][0] ),
    .A1(\cpu0.ram[5][0] ),
    .A2(\cpu0.ram[6][0] ),
    .A3(\cpu0.ram[7][0] ),
    .S1(net155),
    .X(_0274_));
 sg13g2_o21ai_1 _0893_ (.B1(_0273_),
    .Y(_0275_),
    .A1(net146),
    .A2(_0274_));
 sg13g2_mux4_1 _0894_ (.S0(net162),
    .A0(\cpu0.ram[8][0] ),
    .A1(\cpu0.ram[9][0] ),
    .A2(\cpu0.ram[10][0] ),
    .A3(\cpu0.ram[11][0] ),
    .S1(net154),
    .X(_0276_));
 sg13g2_nor2_1 _0895_ (.A(net151),
    .B(_0276_),
    .Y(_0277_));
 sg13g2_mux4_1 _0896_ (.S0(net165),
    .A0(\cpu0.ram[12][0] ),
    .A1(\cpu0.ram[13][0] ),
    .A2(\cpu0.ram[14][0] ),
    .A3(\cpu0.ram[15][0] ),
    .S1(net157),
    .X(_0278_));
 sg13g2_o21ai_1 _0897_ (.B1(net150),
    .Y(_0279_),
    .A1(net146),
    .A2(_0278_));
 sg13g2_or2_1 _0898_ (.X(_0280_),
    .B(_0279_),
    .A(_0277_));
 sg13g2_o21ai_1 _0899_ (.B1(_0280_),
    .Y(_0281_),
    .A1(net149),
    .A2(_0275_));
 sg13g2_a21oi_1 _0900_ (.A1(_0271_),
    .A2(_0281_),
    .Y(_0282_),
    .B1(_0240_));
 sg13g2_nand2_2 _0901_ (.Y(_0283_),
    .A(net145),
    .B(_0227_));
 sg13g2_nor2b_1 _0902_ (.A(\cpu0.a_reg[0] ),
    .B_N(\cpu0.b_reg[0] ),
    .Y(_0284_));
 sg13g2_xor2_1 _0903_ (.B(\cpu0.a_reg[0] ),
    .A(\cpu0.b_reg[0] ),
    .X(_0285_));
 sg13g2_nand2_2 _0904_ (.Y(_0286_),
    .A(\cpu0.step[2] ),
    .B(_0267_));
 sg13g2_nor2_1 _0905_ (.A(_0262_),
    .B(_0286_),
    .Y(_0287_));
 sg13g2_nor3_2 _0906_ (.A(net172),
    .B(_0262_),
    .C(_0286_),
    .Y(_0288_));
 sg13g2_nand2_2 _0907_ (.Y(_0289_),
    .A(net175),
    .B(_0287_));
 sg13g2_a22oi_1 _0908_ (.Y(_0290_),
    .B1(_0285_),
    .B2(_0288_),
    .A2(_0283_),
    .A1(\cpu0.a_reg[0] ));
 sg13g2_nand3_1 _0909_ (.B(_0282_),
    .C(_0290_),
    .A(_0260_),
    .Y(_0291_));
 sg13g2_nand2_2 _0910_ (.Y(_0292_),
    .A(_0241_),
    .B(_0291_));
 sg13g2_inv_1 _0911_ (.Y(_0293_),
    .A(_0292_));
 sg13g2_nor2_1 _0912_ (.A(net1),
    .B(net142),
    .Y(_0294_));
 sg13g2_a21oi_2 _0913_ (.B1(_0294_),
    .Y(_0295_),
    .A2(_0292_),
    .A1(net144));
 sg13g2_mux2_1 _0914_ (.A0(net134),
    .A1(net345),
    .S(_0238_),
    .X(_0008_));
 sg13g2_and4_1 _0915_ (.A(\cpu0.step[2] ),
    .B(_0225_),
    .C(_0239_),
    .D(_0243_),
    .X(_0296_));
 sg13g2_nor2_2 _0916_ (.A(_0261_),
    .B(_0296_),
    .Y(_0297_));
 sg13g2_a21o_2 _0917_ (.A2(_0286_),
    .A1(_0261_),
    .B1(net172),
    .X(_0298_));
 sg13g2_or2_1 _0918_ (.X(_0299_),
    .B(_0298_),
    .A(_0297_));
 sg13g2_o21ai_1 _0919_ (.B1(\cpu0.b_reg[0] ),
    .Y(_0300_),
    .A1(_0297_),
    .A2(_0298_));
 sg13g2_xor2_1 _0920_ (.B(_0300_),
    .A(\cpu0.b_reg[1] ),
    .X(_0301_));
 sg13g2_nand2_1 _0921_ (.Y(_0302_),
    .A(\cpu0.a_reg[1] ),
    .B(_0301_));
 sg13g2_xnor2_1 _0922_ (.Y(_0303_),
    .A(\cpu0.a_reg[1] ),
    .B(_0301_));
 sg13g2_xor2_1 _0923_ (.B(_0303_),
    .A(_0284_),
    .X(_0304_));
 sg13g2_a21oi_1 _0924_ (.A1(\cpu0.ir[1] ),
    .A2(_0259_),
    .Y(_0305_),
    .B1(_0271_));
 sg13g2_a22oi_1 _0925_ (.Y(_0306_),
    .B1(_0288_),
    .B2(_0304_),
    .A2(_0283_),
    .A1(\cpu0.a_reg[1] ));
 sg13g2_nand2_1 _0926_ (.Y(_0307_),
    .A(_0305_),
    .B(_0306_));
 sg13g2_nand2b_1 _0927_ (.Y(_0308_),
    .B(net164),
    .A_N(\cpu0.ram[1][1] ));
 sg13g2_o21ai_1 _0928_ (.B1(_0308_),
    .Y(_0309_),
    .A1(net164),
    .A2(\cpu0.ram[0][1] ));
 sg13g2_mux2_1 _0929_ (.A0(\cpu0.ram[2][1] ),
    .A1(\cpu0.ram[3][1] ),
    .S(net163),
    .X(_0310_));
 sg13g2_a21oi_1 _0930_ (.A1(net156),
    .A2(_0310_),
    .Y(_0311_),
    .B1(net152));
 sg13g2_o21ai_1 _0931_ (.B1(_0311_),
    .Y(_0312_),
    .A1(net155),
    .A2(_0309_));
 sg13g2_nor2b_1 _0932_ (.A(net170),
    .B_N(\cpu0.ram[4][1] ),
    .Y(_0313_));
 sg13g2_a21oi_1 _0933_ (.A1(net170),
    .A2(\cpu0.ram[5][1] ),
    .Y(_0314_),
    .B1(_0313_));
 sg13g2_o21ai_1 _0934_ (.B1(net159),
    .Y(_0315_),
    .A1(net170),
    .A2(\cpu0.ram[6][1] ));
 sg13g2_a21oi_1 _0935_ (.A1(net170),
    .A2(_0205_),
    .Y(_0316_),
    .B1(_0315_));
 sg13g2_o21ai_1 _0936_ (.B1(net153),
    .Y(_0317_),
    .A1(net159),
    .A2(_0314_));
 sg13g2_o21ai_1 _0937_ (.B1(_0312_),
    .Y(_0318_),
    .A1(_0316_),
    .A2(_0317_));
 sg13g2_nor2b_1 _0938_ (.A(net160),
    .B_N(\cpu0.ram[8][1] ),
    .Y(_0319_));
 sg13g2_a21oi_1 _0939_ (.A1(net160),
    .A2(\cpu0.ram[9][1] ),
    .Y(_0320_),
    .B1(_0319_));
 sg13g2_mux2_1 _0940_ (.A0(\cpu0.ram[10][1] ),
    .A1(\cpu0.ram[11][1] ),
    .S(net160),
    .X(_0321_));
 sg13g2_a21oi_1 _0941_ (.A1(net154),
    .A2(_0321_),
    .Y(_0322_),
    .B1(net151));
 sg13g2_o21ai_1 _0942_ (.B1(_0322_),
    .Y(_0323_),
    .A1(net156),
    .A2(_0320_));
 sg13g2_a21oi_1 _0943_ (.A1(net167),
    .A2(_0206_),
    .Y(_0324_),
    .B1(net158));
 sg13g2_o21ai_1 _0944_ (.B1(_0324_),
    .Y(_0325_),
    .A1(net167),
    .A2(\cpu0.ram[12][1] ));
 sg13g2_mux2_1 _0945_ (.A0(\cpu0.ram[14][1] ),
    .A1(\cpu0.ram[15][1] ),
    .S(net167),
    .X(_0326_));
 sg13g2_a21oi_1 _0946_ (.A1(net157),
    .A2(_0326_),
    .Y(_0327_),
    .B1(net146));
 sg13g2_nand2_1 _0947_ (.Y(_0328_),
    .A(_0325_),
    .B(_0327_));
 sg13g2_nand3_1 _0948_ (.B(_0323_),
    .C(_0328_),
    .A(net150),
    .Y(_0329_));
 sg13g2_and2_1 _0949_ (.A(_0271_),
    .B(_0329_),
    .X(_0330_));
 sg13g2_o21ai_1 _0950_ (.B1(_0330_),
    .Y(_0331_),
    .A1(net149),
    .A2(_0318_));
 sg13g2_a22oi_1 _0951_ (.Y(_0332_),
    .B1(_0307_),
    .B2(_0331_),
    .A2(_0240_),
    .A1(\cpu0.pc[1] ));
 sg13g2_nor2_1 _0952_ (.A(net2),
    .B(net142),
    .Y(_0333_));
 sg13g2_a21oi_2 _0953_ (.B1(_0333_),
    .Y(_0334_),
    .A2(_0332_),
    .A1(net143));
 sg13g2_mux2_1 _0954_ (.A0(net132),
    .A1(net430),
    .S(_0238_),
    .X(_0009_));
 sg13g2_o21ai_1 _0955_ (.B1(_0302_),
    .Y(_0335_),
    .A1(_0284_),
    .A2(_0303_));
 sg13g2_or2_1 _0956_ (.X(_0336_),
    .B(\cpu0.b_reg[0] ),
    .A(\cpu0.b_reg[1] ));
 sg13g2_o21ai_1 _0957_ (.B1(_0336_),
    .Y(_0337_),
    .A1(_0297_),
    .A2(_0298_));
 sg13g2_xor2_1 _0958_ (.B(_0337_),
    .A(\cpu0.b_reg[2] ),
    .X(_0338_));
 sg13g2_and2_1 _0959_ (.A(\cpu0.a_reg[2] ),
    .B(_0338_),
    .X(_0339_));
 sg13g2_xnor2_1 _0960_ (.Y(_0340_),
    .A(\cpu0.a_reg[2] ),
    .B(_0338_));
 sg13g2_nand2b_1 _0961_ (.Y(_0341_),
    .B(_0340_),
    .A_N(_0335_));
 sg13g2_nand2b_1 _0962_ (.Y(_0342_),
    .B(_0335_),
    .A_N(_0340_));
 sg13g2_nand3_1 _0963_ (.B(_0341_),
    .C(_0342_),
    .A(_0288_),
    .Y(_0343_));
 sg13g2_a21oi_1 _0964_ (.A1(\cpu0.a_reg[2] ),
    .A2(_0283_),
    .Y(_0344_),
    .B1(_0259_));
 sg13g2_a221oi_1 _0965_ (.B2(_0344_),
    .C1(_0271_),
    .B1(_0343_),
    .A1(_0197_),
    .Y(_0345_),
    .A2(_0259_));
 sg13g2_a21oi_1 _0966_ (.A1(net167),
    .A2(\cpu0.ram[13][2] ),
    .Y(_0346_),
    .B1(net158));
 sg13g2_o21ai_1 _0967_ (.B1(_0346_),
    .Y(_0347_),
    .A1(net167),
    .A2(_0207_));
 sg13g2_a21oi_1 _0968_ (.A1(net168),
    .A2(\cpu0.ram[15][2] ),
    .Y(_0348_),
    .B1(net147));
 sg13g2_o21ai_1 _0969_ (.B1(_0348_),
    .Y(_0349_),
    .A1(net167),
    .A2(_0208_));
 sg13g2_nand3_1 _0970_ (.B(_0347_),
    .C(_0349_),
    .A(net153),
    .Y(_0350_));
 sg13g2_mux4_1 _0971_ (.S0(net162),
    .A0(\cpu0.ram[8][2] ),
    .A1(\cpu0.ram[9][2] ),
    .A2(\cpu0.ram[10][2] ),
    .A3(\cpu0.ram[11][2] ),
    .S1(net154),
    .X(_0351_));
 sg13g2_nand2_1 _0972_ (.Y(_0352_),
    .A(net146),
    .B(_0351_));
 sg13g2_nand3_1 _0973_ (.B(_0350_),
    .C(_0352_),
    .A(net150),
    .Y(_0353_));
 sg13g2_mux4_1 _0974_ (.S0(net163),
    .A0(\cpu0.ram[0][2] ),
    .A1(\cpu0.ram[1][2] ),
    .A2(\cpu0.ram[2][2] ),
    .A3(\cpu0.ram[3][2] ),
    .S1(net155),
    .X(_0354_));
 sg13g2_nand2_1 _0975_ (.Y(_0355_),
    .A(net146),
    .B(_0354_));
 sg13g2_nor2b_1 _0976_ (.A(net170),
    .B_N(\cpu0.ram[4][2] ),
    .Y(_0356_));
 sg13g2_a21oi_1 _0977_ (.A1(net170),
    .A2(\cpu0.ram[5][2] ),
    .Y(_0357_),
    .B1(_0356_));
 sg13g2_nand2b_1 _0978_ (.Y(_0358_),
    .B(\cpu0.ram[6][2] ),
    .A_N(net171));
 sg13g2_a21oi_1 _0979_ (.A1(net171),
    .A2(\cpu0.ram[7][2] ),
    .Y(_0359_),
    .B1(net147));
 sg13g2_a221oi_1 _0980_ (.B2(_0359_),
    .C1(net146),
    .B1(_0358_),
    .A1(net147),
    .Y(_0360_),
    .A2(_0357_));
 sg13g2_nor2_1 _0981_ (.A(net149),
    .B(_0360_),
    .Y(_0361_));
 sg13g2_a21oi_1 _0982_ (.A1(_0355_),
    .A2(_0361_),
    .Y(_0362_),
    .B1(_0270_));
 sg13g2_a221oi_1 _0983_ (.B2(_0362_),
    .C1(_0345_),
    .B1(_0353_),
    .A1(\cpu0.pc[2] ),
    .Y(_0363_),
    .A2(_0240_));
 sg13g2_nor2_1 _0984_ (.A(net3),
    .B(net142),
    .Y(_0364_));
 sg13g2_a21oi_2 _0985_ (.B1(_0364_),
    .Y(_0365_),
    .A2(_0363_),
    .A1(net143));
 sg13g2_mux2_1 _0986_ (.A0(net130),
    .A1(net376),
    .S(_0238_),
    .X(_0010_));
 sg13g2_a21oi_1 _0987_ (.A1(\cpu0.a_reg[3] ),
    .A2(_0283_),
    .Y(_0366_),
    .B1(_0259_));
 sg13g2_or2_1 _0988_ (.X(_0367_),
    .B(_0336_),
    .A(\cpu0.b_reg[2] ));
 sg13g2_o21ai_1 _0989_ (.B1(_0367_),
    .Y(_0368_),
    .A1(_0297_),
    .A2(_0298_));
 sg13g2_xnor2_1 _0990_ (.Y(_0369_),
    .A(\cpu0.b_reg[3] ),
    .B(_0368_));
 sg13g2_nand2b_1 _0991_ (.Y(_0370_),
    .B(_0369_),
    .A_N(\cpu0.a_reg[3] ));
 sg13g2_nor2b_1 _0992_ (.A(_0369_),
    .B_N(\cpu0.a_reg[3] ),
    .Y(_0371_));
 sg13g2_xnor2_1 _0993_ (.Y(_0372_),
    .A(\cpu0.a_reg[3] ),
    .B(_0369_));
 sg13g2_nand2b_1 _0994_ (.Y(_0373_),
    .B(_0342_),
    .A_N(_0339_));
 sg13g2_xnor2_1 _0995_ (.Y(_0374_),
    .A(_0372_),
    .B(_0373_));
 sg13g2_o21ai_1 _0996_ (.B1(_0366_),
    .Y(_0375_),
    .A1(_0289_),
    .A2(_0374_));
 sg13g2_a21oi_1 _0997_ (.A1(_0196_),
    .A2(_0259_),
    .Y(_0376_),
    .B1(_0271_));
 sg13g2_mux2_1 _0998_ (.A0(\cpu0.ram[12][3] ),
    .A1(\cpu0.ram[13][3] ),
    .S(net168),
    .X(_0377_));
 sg13g2_o21ai_1 _0999_ (.B1(net158),
    .Y(_0378_),
    .A1(net167),
    .A2(_0210_));
 sg13g2_a21oi_1 _1000_ (.A1(net167),
    .A2(\cpu0.ram[15][3] ),
    .Y(_0379_),
    .B1(_0378_));
 sg13g2_o21ai_1 _1001_ (.B1(net153),
    .Y(_0380_),
    .A1(net157),
    .A2(_0377_));
 sg13g2_nor2b_1 _1002_ (.A(net160),
    .B_N(\cpu0.ram[8][3] ),
    .Y(_0381_));
 sg13g2_a21oi_1 _1003_ (.A1(net161),
    .A2(\cpu0.ram[9][3] ),
    .Y(_0382_),
    .B1(_0381_));
 sg13g2_nand2b_1 _1004_ (.Y(_0383_),
    .B(\cpu0.ram[10][3] ),
    .A_N(net161));
 sg13g2_a21oi_1 _1005_ (.A1(net160),
    .A2(\cpu0.ram[11][3] ),
    .Y(_0384_),
    .B1(net147));
 sg13g2_a221oi_1 _1006_ (.B2(_0384_),
    .C1(net151),
    .B1(_0383_),
    .A1(net147),
    .Y(_0385_),
    .A2(_0382_));
 sg13g2_o21ai_1 _1007_ (.B1(net150),
    .Y(_0386_),
    .A1(_0379_),
    .A2(_0380_));
 sg13g2_nor2_1 _1008_ (.A(_0385_),
    .B(_0386_),
    .Y(_0387_));
 sg13g2_mux4_1 _1009_ (.S0(net164),
    .A0(\cpu0.ram[0][3] ),
    .A1(\cpu0.ram[1][3] ),
    .A2(\cpu0.ram[2][3] ),
    .A3(\cpu0.ram[3][3] ),
    .S1(net156),
    .X(_0388_));
 sg13g2_a21oi_1 _1010_ (.A1(net170),
    .A2(\cpu0.ram[5][3] ),
    .Y(_0389_),
    .B1(net159));
 sg13g2_o21ai_1 _1011_ (.B1(_0389_),
    .Y(_0390_),
    .A1(net170),
    .A2(_0209_));
 sg13g2_nor2b_1 _1012_ (.A(net168),
    .B_N(\cpu0.ram[6][3] ),
    .Y(_0391_));
 sg13g2_a21oi_1 _1013_ (.A1(net168),
    .A2(\cpu0.ram[7][3] ),
    .Y(_0392_),
    .B1(_0391_));
 sg13g2_a21oi_1 _1014_ (.A1(net159),
    .A2(_0392_),
    .Y(_0393_),
    .B1(net146));
 sg13g2_a221oi_1 _1015_ (.B2(_0393_),
    .C1(net150),
    .B1(_0390_),
    .A1(_0204_),
    .Y(_0394_),
    .A2(_0388_));
 sg13g2_nor3_1 _1016_ (.A(_0270_),
    .B(_0387_),
    .C(_0394_),
    .Y(_0395_));
 sg13g2_a221oi_1 _1017_ (.B2(_0376_),
    .C1(_0395_),
    .B1(_0375_),
    .A1(\cpu0.pc[3] ),
    .Y(_0396_),
    .A2(_0240_));
 sg13g2_nor2_1 _1018_ (.A(net4),
    .B(net142),
    .Y(_0397_));
 sg13g2_a21oi_2 _1019_ (.B1(_0397_),
    .Y(_0398_),
    .A2(_0396_),
    .A1(net143));
 sg13g2_mux2_1 _1020_ (.A0(net126),
    .A1(net360),
    .S(_0238_),
    .X(_0011_));
 sg13g2_mux4_1 _1021_ (.S0(net160),
    .A0(\cpu0.ram[12][4] ),
    .A1(\cpu0.ram[13][4] ),
    .A2(\cpu0.ram[14][4] ),
    .A3(\cpu0.ram[15][4] ),
    .S1(net154),
    .X(_0399_));
 sg13g2_mux4_1 _1022_ (.S0(net162),
    .A0(\cpu0.ram[8][4] ),
    .A1(\cpu0.ram[9][4] ),
    .A2(\cpu0.ram[10][4] ),
    .A3(\cpu0.ram[11][4] ),
    .S1(net154),
    .X(_0400_));
 sg13g2_mux4_1 _1023_ (.S0(net161),
    .A0(\cpu0.ram[4][4] ),
    .A1(\cpu0.ram[5][4] ),
    .A2(\cpu0.ram[6][4] ),
    .A3(\cpu0.ram[7][4] ),
    .S1(net154),
    .X(_0401_));
 sg13g2_mux4_1 _1024_ (.S0(net163),
    .A0(\cpu0.ram[0][4] ),
    .A1(\cpu0.ram[1][4] ),
    .A2(\cpu0.ram[2][4] ),
    .A3(\cpu0.ram[3][4] ),
    .S1(net155),
    .X(_0402_));
 sg13g2_mux4_1 _1025_ (.S0(net152),
    .A0(_0402_),
    .A1(_0401_),
    .A2(_0400_),
    .A3(_0399_),
    .S1(net149),
    .X(_0403_));
 sg13g2_nor2_1 _1026_ (.A(_0270_),
    .B(_0403_),
    .Y(_0404_));
 sg13g2_nor2b_1 _1027_ (.A(_0340_),
    .B_N(_0372_),
    .Y(_0405_));
 sg13g2_a221oi_1 _1028_ (.B2(_0335_),
    .C1(_0371_),
    .B1(_0405_),
    .A1(_0339_),
    .Y(_0406_),
    .A2(_0370_));
 sg13g2_or2_1 _1029_ (.X(_0407_),
    .B(_0367_),
    .A(\cpu0.b_reg[3] ));
 sg13g2_nand2_1 _1030_ (.Y(_0408_),
    .A(_0299_),
    .B(_0407_));
 sg13g2_xnor2_1 _1031_ (.Y(_0409_),
    .A(\cpu0.b_reg[4] ),
    .B(_0408_));
 sg13g2_or2_1 _1032_ (.X(_0410_),
    .B(_0409_),
    .A(_0198_));
 sg13g2_xnor2_1 _1033_ (.Y(_0411_),
    .A(_0198_),
    .B(_0409_));
 sg13g2_or2_1 _1034_ (.X(_0412_),
    .B(_0411_),
    .A(_0406_));
 sg13g2_a21oi_1 _1035_ (.A1(_0406_),
    .A2(_0411_),
    .Y(_0413_),
    .B1(_0289_));
 sg13g2_nand2_1 _1036_ (.Y(_0414_),
    .A(_0412_),
    .B(_0413_));
 sg13g2_a21oi_1 _1037_ (.A1(net337),
    .A2(_0283_),
    .Y(_0415_),
    .B1(_0271_));
 sg13g2_a21oi_2 _1038_ (.B1(_0404_),
    .Y(_0416_),
    .A2(_0415_),
    .A1(_0414_));
 sg13g2_mux2_1 _1039_ (.A0(net5),
    .A1(_0416_),
    .S(net144),
    .X(_0417_));
 sg13g2_mux2_1 _1040_ (.A0(net128),
    .A1(net397),
    .S(_0238_),
    .X(_0012_));
 sg13g2_nor2_1 _1041_ (.A(net6),
    .B(net142),
    .Y(_0418_));
 sg13g2_or2_1 _1042_ (.X(_0419_),
    .B(_0407_),
    .A(\cpu0.b_reg[4] ));
 sg13g2_nand2_1 _1043_ (.Y(_0420_),
    .A(_0299_),
    .B(_0419_));
 sg13g2_xnor2_1 _1044_ (.Y(_0421_),
    .A(\cpu0.b_reg[5] ),
    .B(_0420_));
 sg13g2_nand2b_1 _1045_ (.Y(_0422_),
    .B(\cpu0.a_reg[5] ),
    .A_N(_0421_));
 sg13g2_xor2_1 _1046_ (.B(_0421_),
    .A(\cpu0.a_reg[5] ),
    .X(_0423_));
 sg13g2_nand3_1 _1047_ (.B(_0412_),
    .C(_0423_),
    .A(_0410_),
    .Y(_0424_));
 sg13g2_nor2_1 _1048_ (.A(_0411_),
    .B(_0423_),
    .Y(_0425_));
 sg13g2_nor2b_1 _1049_ (.A(_0406_),
    .B_N(_0425_),
    .Y(_0426_));
 sg13g2_o21ai_1 _1050_ (.B1(_0288_),
    .Y(_0427_),
    .A1(_0410_),
    .A2(_0423_));
 sg13g2_nor2_1 _1051_ (.A(_0426_),
    .B(_0427_),
    .Y(_0428_));
 sg13g2_a221oi_1 _1052_ (.B2(_0428_),
    .C1(_0271_),
    .B1(_0424_),
    .A1(\cpu0.a_reg[5] ),
    .Y(_0429_),
    .A2(_0283_));
 sg13g2_mux4_1 _1053_ (.S0(net165),
    .A0(\cpu0.ram[12][5] ),
    .A1(\cpu0.ram[13][5] ),
    .A2(\cpu0.ram[14][5] ),
    .A3(\cpu0.ram[15][5] ),
    .S1(net158),
    .X(_0430_));
 sg13g2_mux4_1 _1054_ (.S0(net160),
    .A0(\cpu0.ram[8][5] ),
    .A1(\cpu0.ram[9][5] ),
    .A2(\cpu0.ram[10][5] ),
    .A3(\cpu0.ram[11][5] ),
    .S1(net156),
    .X(_0431_));
 sg13g2_mux2_1 _1055_ (.A0(_0430_),
    .A1(_0431_),
    .S(net146),
    .X(_0432_));
 sg13g2_mux4_1 _1056_ (.S0(net163),
    .A0(\cpu0.ram[0][5] ),
    .A1(\cpu0.ram[1][5] ),
    .A2(\cpu0.ram[2][5] ),
    .A3(\cpu0.ram[3][5] ),
    .S1(net155),
    .X(_0433_));
 sg13g2_mux2_1 _1057_ (.A0(\cpu0.ram[4][5] ),
    .A1(\cpu0.ram[5][5] ),
    .S(net168),
    .X(_0434_));
 sg13g2_nor2b_1 _1058_ (.A(\cpu0.ram[7][5] ),
    .B_N(net168),
    .Y(_0435_));
 sg13g2_o21ai_1 _1059_ (.B1(net158),
    .Y(_0436_),
    .A1(net168),
    .A2(\cpu0.ram[6][5] ));
 sg13g2_o21ai_1 _1060_ (.B1(net153),
    .Y(_0437_),
    .A1(_0435_),
    .A2(_0436_));
 sg13g2_a21oi_1 _1061_ (.A1(net147),
    .A2(_0434_),
    .Y(_0438_),
    .B1(_0437_));
 sg13g2_nor2_1 _1062_ (.A(net149),
    .B(_0438_),
    .Y(_0439_));
 sg13g2_o21ai_1 _1063_ (.B1(_0439_),
    .Y(_0440_),
    .A1(net152),
    .A2(_0433_));
 sg13g2_a21oi_1 _1064_ (.A1(net149),
    .A2(_0432_),
    .Y(_0441_),
    .B1(_0270_));
 sg13g2_a21o_2 _1065_ (.A2(_0441_),
    .A1(_0440_),
    .B1(_0429_),
    .X(_0442_));
 sg13g2_inv_1 _1066_ (.Y(_0443_),
    .A(_0442_));
 sg13g2_a21oi_2 _1067_ (.B1(_0418_),
    .Y(_0444_),
    .A2(_0442_),
    .A1(net142));
 sg13g2_mux2_1 _1068_ (.A0(net124),
    .A1(net336),
    .S(_0238_),
    .X(_0013_));
 sg13g2_o21ai_1 _1069_ (.B1(_0299_),
    .Y(_0445_),
    .A1(\cpu0.b_reg[5] ),
    .A2(_0419_));
 sg13g2_xor2_1 _1070_ (.B(_0445_),
    .A(\cpu0.b_reg[6] ),
    .X(_0446_));
 sg13g2_nand2_1 _1071_ (.Y(_0447_),
    .A(\cpu0.a_reg[6] ),
    .B(_0446_));
 sg13g2_xor2_1 _1072_ (.B(_0446_),
    .A(\cpu0.a_reg[6] ),
    .X(_0448_));
 sg13g2_o21ai_1 _1073_ (.B1(_0422_),
    .Y(_0449_),
    .A1(_0410_),
    .A2(_0423_));
 sg13g2_o21ai_1 _1074_ (.B1(_0448_),
    .Y(_0450_),
    .A1(_0426_),
    .A2(_0449_));
 sg13g2_nor3_1 _1075_ (.A(_0426_),
    .B(_0448_),
    .C(_0449_),
    .Y(_0451_));
 sg13g2_nor2_1 _1076_ (.A(_0289_),
    .B(_0451_),
    .Y(_0452_));
 sg13g2_a22oi_1 _1077_ (.Y(_0453_),
    .B1(_0450_),
    .B2(_0452_),
    .A2(_0283_),
    .A1(\cpu0.a_reg[6] ));
 sg13g2_mux4_1 _1078_ (.S0(net163),
    .A0(\cpu0.ram[0][6] ),
    .A1(\cpu0.ram[1][6] ),
    .A2(\cpu0.ram[2][6] ),
    .A3(\cpu0.ram[3][6] ),
    .S1(net155),
    .X(_0454_));
 sg13g2_mux2_1 _1079_ (.A0(\cpu0.ram[4][6] ),
    .A1(\cpu0.ram[5][6] ),
    .S(net165),
    .X(_0455_));
 sg13g2_nor2b_1 _1080_ (.A(\cpu0.ram[7][6] ),
    .B_N(net166),
    .Y(_0456_));
 sg13g2_o21ai_1 _1081_ (.B1(net157),
    .Y(_0457_),
    .A1(net166),
    .A2(\cpu0.ram[6][6] ));
 sg13g2_o21ai_1 _1082_ (.B1(net153),
    .Y(_0458_),
    .A1(_0456_),
    .A2(_0457_));
 sg13g2_a21oi_1 _1083_ (.A1(_0203_),
    .A2(_0455_),
    .Y(_0459_),
    .B1(_0458_));
 sg13g2_nor2_1 _1084_ (.A(net149),
    .B(_0459_),
    .Y(_0460_));
 sg13g2_o21ai_1 _1085_ (.B1(_0460_),
    .Y(_0461_),
    .A1(net151),
    .A2(_0454_));
 sg13g2_mux4_1 _1086_ (.S0(net162),
    .A0(\cpu0.ram[8][6] ),
    .A1(\cpu0.ram[9][6] ),
    .A2(\cpu0.ram[10][6] ),
    .A3(\cpu0.ram[11][6] ),
    .S1(net154),
    .X(_0462_));
 sg13g2_nor2_1 _1087_ (.A(net151),
    .B(_0462_),
    .Y(_0463_));
 sg13g2_o21ai_1 _1088_ (.B1(_0203_),
    .Y(_0464_),
    .A1(net165),
    .A2(\cpu0.ram[12][6] ));
 sg13g2_a21oi_1 _1089_ (.A1(net165),
    .A2(_0211_),
    .Y(_0465_),
    .B1(_0464_));
 sg13g2_nor2b_1 _1090_ (.A(\cpu0.ram[15][6] ),
    .B_N(net165),
    .Y(_0466_));
 sg13g2_o21ai_1 _1091_ (.B1(net157),
    .Y(_0467_),
    .A1(net165),
    .A2(\cpu0.ram[14][6] ));
 sg13g2_o21ai_1 _1092_ (.B1(_0002_),
    .Y(_0468_),
    .A1(_0466_),
    .A2(_0467_));
 sg13g2_o21ai_1 _1093_ (.B1(net150),
    .Y(_0469_),
    .A1(_0465_),
    .A2(_0468_));
 sg13g2_o21ai_1 _1094_ (.B1(_0461_),
    .Y(_0470_),
    .A1(_0463_),
    .A2(_0469_));
 sg13g2_nor2_1 _1095_ (.A(_0270_),
    .B(_0470_),
    .Y(_0471_));
 sg13g2_a21o_2 _1096_ (.A2(_0453_),
    .A1(_0270_),
    .B1(_0471_),
    .X(_0472_));
 sg13g2_nor2_1 _1097_ (.A(net7),
    .B(net142),
    .Y(_0473_));
 sg13g2_a21oi_2 _1098_ (.B1(_0473_),
    .Y(_0474_),
    .A2(_0472_),
    .A1(net144));
 sg13g2_mux2_1 _1099_ (.A0(net122),
    .A1(net413),
    .S(_0238_),
    .X(_0014_));
 sg13g2_nand2_1 _1100_ (.Y(_0475_),
    .A(\cpu0.b_reg[6] ),
    .B(_0299_));
 sg13g2_nand2_1 _1101_ (.Y(_0476_),
    .A(_0445_),
    .B(_0475_));
 sg13g2_xnor2_1 _1102_ (.Y(_0477_),
    .A(\cpu0.b_reg[7] ),
    .B(_0476_));
 sg13g2_nand2_1 _1103_ (.Y(_0478_),
    .A(\cpu0.a_reg[7] ),
    .B(_0477_));
 sg13g2_xnor2_1 _1104_ (.Y(_0479_),
    .A(\cpu0.a_reg[7] ),
    .B(_0477_));
 sg13g2_nand3_1 _1105_ (.B(_0450_),
    .C(_0479_),
    .A(_0447_),
    .Y(_0480_));
 sg13g2_a21o_1 _1106_ (.A2(_0450_),
    .A1(_0447_),
    .B1(_0479_),
    .X(_0481_));
 sg13g2_nand3_1 _1107_ (.B(_0480_),
    .C(_0481_),
    .A(_0288_),
    .Y(_0482_));
 sg13g2_a21oi_1 _1108_ (.A1(\cpu0.a_reg[7] ),
    .A2(_0283_),
    .Y(_0483_),
    .B1(_0271_));
 sg13g2_mux4_1 _1109_ (.S0(net163),
    .A0(\cpu0.ram[0][7] ),
    .A1(\cpu0.ram[1][7] ),
    .A2(\cpu0.ram[2][7] ),
    .A3(\cpu0.ram[3][7] ),
    .S1(net155),
    .X(_0484_));
 sg13g2_mux2_1 _1110_ (.A0(\cpu0.ram[4][7] ),
    .A1(\cpu0.ram[5][7] ),
    .S(net171),
    .X(_0485_));
 sg13g2_nor2b_1 _1111_ (.A(\cpu0.ram[7][7] ),
    .B_N(net171),
    .Y(_0486_));
 sg13g2_o21ai_1 _1112_ (.B1(net157),
    .Y(_0487_),
    .A1(net165),
    .A2(\cpu0.ram[6][7] ));
 sg13g2_o21ai_1 _1113_ (.B1(net152),
    .Y(_0488_),
    .A1(_0486_),
    .A2(_0487_));
 sg13g2_a21oi_1 _1114_ (.A1(net147),
    .A2(_0485_),
    .Y(_0489_),
    .B1(_0488_));
 sg13g2_nor2_1 _1115_ (.A(net149),
    .B(_0489_),
    .Y(_0490_));
 sg13g2_o21ai_1 _1116_ (.B1(_0490_),
    .Y(_0491_),
    .A1(net151),
    .A2(_0484_));
 sg13g2_mux4_1 _1117_ (.S0(net162),
    .A0(\cpu0.ram[8][7] ),
    .A1(\cpu0.ram[9][7] ),
    .A2(\cpu0.ram[10][7] ),
    .A3(\cpu0.ram[11][7] ),
    .S1(net154),
    .X(_0492_));
 sg13g2_nor2_1 _1118_ (.A(net151),
    .B(_0492_),
    .Y(_0493_));
 sg13g2_nor2b_1 _1119_ (.A(\cpu0.ram[13][7] ),
    .B_N(net160),
    .Y(_0494_));
 sg13g2_o21ai_1 _1120_ (.B1(net147),
    .Y(_0495_),
    .A1(net161),
    .A2(\cpu0.ram[12][7] ));
 sg13g2_o21ai_1 _1121_ (.B1(net157),
    .Y(_0496_),
    .A1(net166),
    .A2(\cpu0.ram[14][7] ));
 sg13g2_a21oi_1 _1122_ (.A1(net166),
    .A2(_0212_),
    .Y(_0497_),
    .B1(_0496_));
 sg13g2_o21ai_1 _1123_ (.B1(net151),
    .Y(_0498_),
    .A1(_0494_),
    .A2(_0495_));
 sg13g2_o21ai_1 _1124_ (.B1(net150),
    .Y(_0499_),
    .A1(_0497_),
    .A2(_0498_));
 sg13g2_nor2_1 _1125_ (.A(_0493_),
    .B(_0499_),
    .Y(_0500_));
 sg13g2_nor2_1 _1126_ (.A(_0270_),
    .B(_0500_),
    .Y(_0501_));
 sg13g2_a22oi_1 _1127_ (.Y(_0502_),
    .B1(_0491_),
    .B2(_0501_),
    .A2(_0483_),
    .A1(_0482_));
 sg13g2_mux2_1 _1128_ (.A0(net8),
    .A1(_0502_),
    .S(net144),
    .X(_0503_));
 sg13g2_mux2_1 _1129_ (.A0(net120),
    .A1(net394),
    .S(_0238_),
    .X(_0015_));
 sg13g2_o21ai_1 _1130_ (.B1(_0225_),
    .Y(_0504_),
    .A1(_0193_),
    .A2(_0194_));
 sg13g2_a21oi_1 _1131_ (.A1(_0262_),
    .A2(_0504_),
    .Y(_0505_),
    .B1(_0217_));
 sg13g2_or2_1 _1132_ (.X(_0506_),
    .B(_0505_),
    .A(_0240_));
 sg13g2_o21ai_1 _1133_ (.B1(net175),
    .Y(_0507_),
    .A1(net482),
    .A2(net139));
 sg13g2_a21oi_1 _1134_ (.A1(_0292_),
    .A2(net139),
    .Y(_0016_),
    .B1(_0507_));
 sg13g2_o21ai_1 _1135_ (.B1(net175),
    .Y(_0508_),
    .A1(net479),
    .A2(net139));
 sg13g2_a21oi_1 _1136_ (.A1(_0332_),
    .A2(net140),
    .Y(_0017_),
    .B1(_0508_));
 sg13g2_o21ai_1 _1137_ (.B1(net175),
    .Y(_0509_),
    .A1(net475),
    .A2(net139));
 sg13g2_a21oi_1 _1138_ (.A1(_0363_),
    .A2(net139),
    .Y(_0018_),
    .B1(_0509_));
 sg13g2_o21ai_1 _1139_ (.B1(net177),
    .Y(_0510_),
    .A1(net467),
    .A2(net140));
 sg13g2_a21oi_1 _1140_ (.A1(_0396_),
    .A2(net140),
    .Y(_0019_),
    .B1(_0510_));
 sg13g2_nor2_2 _1141_ (.A(_0235_),
    .B(_0236_),
    .Y(_0511_));
 sg13g2_nand2_1 _1142_ (.Y(_0512_),
    .A(_0228_),
    .B(_0230_));
 sg13g2_nand3_1 _1143_ (.B(_0230_),
    .C(_0233_),
    .A(_0228_),
    .Y(_0513_));
 sg13g2_nand4_1 _1144_ (.B(_0230_),
    .C(_0233_),
    .A(_0228_),
    .Y(_0514_),
    .D(_0511_));
 sg13g2_mux2_1 _1145_ (.A0(net133),
    .A1(net416),
    .S(_0514_),
    .X(_0020_));
 sg13g2_mux2_1 _1146_ (.A0(net131),
    .A1(net329),
    .S(_0514_),
    .X(_0021_));
 sg13g2_mux2_1 _1147_ (.A0(net129),
    .A1(net392),
    .S(_0514_),
    .X(_0022_));
 sg13g2_mux2_1 _1148_ (.A0(net125),
    .A1(net440),
    .S(_0514_),
    .X(_0023_));
 sg13g2_mux2_1 _1149_ (.A0(net127),
    .A1(net390),
    .S(_0514_),
    .X(_0024_));
 sg13g2_mux2_1 _1150_ (.A0(net123),
    .A1(net363),
    .S(_0514_),
    .X(_0025_));
 sg13g2_mux2_1 _1151_ (.A0(net121),
    .A1(net388),
    .S(_0514_),
    .X(_0026_));
 sg13g2_mux2_1 _1152_ (.A0(net119),
    .A1(net402),
    .S(_0514_),
    .X(_0027_));
 sg13g2_o21ai_1 _1153_ (.B1(net177),
    .Y(_0515_),
    .A1(net469),
    .A2(_0267_));
 sg13g2_inv_1 _1154_ (.Y(_0028_),
    .A(_0515_));
 sg13g2_nand3_1 _1155_ (.B(net463),
    .C(_0214_),
    .A(net177),
    .Y(_0516_));
 sg13g2_nand2_1 _1156_ (.Y(_0029_),
    .A(_0217_),
    .B(net464));
 sg13g2_nand2_1 _1157_ (.Y(_0517_),
    .A(_0231_),
    .B(_0233_));
 sg13g2_or2_1 _1158_ (.X(_0518_),
    .B(_0517_),
    .A(_0237_));
 sg13g2_mux2_1 _1159_ (.A0(net134),
    .A1(net343),
    .S(_0518_),
    .X(_0030_));
 sg13g2_mux2_1 _1160_ (.A0(net132),
    .A1(net372),
    .S(_0518_),
    .X(_0031_));
 sg13g2_mux2_1 _1161_ (.A0(net130),
    .A1(net317),
    .S(_0518_),
    .X(_0032_));
 sg13g2_mux2_1 _1162_ (.A0(net126),
    .A1(net365),
    .S(_0518_),
    .X(_0033_));
 sg13g2_mux2_1 _1163_ (.A0(net128),
    .A1(net355),
    .S(_0518_),
    .X(_0034_));
 sg13g2_mux2_1 _1164_ (.A0(net124),
    .A1(net404),
    .S(_0518_),
    .X(_0035_));
 sg13g2_mux2_1 _1165_ (.A0(net122),
    .A1(net421),
    .S(_0518_),
    .X(_0036_));
 sg13g2_mux2_1 _1166_ (.A0(net120),
    .A1(net322),
    .S(_0518_),
    .X(_0037_));
 sg13g2_nor2_2 _1167_ (.A(_0233_),
    .B(_0512_),
    .Y(_0519_));
 sg13g2_nand2_2 _1168_ (.Y(_0520_),
    .A(_0511_),
    .B(_0519_));
 sg13g2_mux2_1 _1169_ (.A0(net133),
    .A1(net359),
    .S(_0520_),
    .X(_0038_));
 sg13g2_mux2_1 _1170_ (.A0(net131),
    .A1(net442),
    .S(_0520_),
    .X(_0039_));
 sg13g2_mux2_1 _1171_ (.A0(net129),
    .A1(net391),
    .S(_0520_),
    .X(_0040_));
 sg13g2_mux2_1 _1172_ (.A0(net125),
    .A1(net371),
    .S(_0520_),
    .X(_0041_));
 sg13g2_mux2_1 _1173_ (.A0(net127),
    .A1(net342),
    .S(_0520_),
    .X(_0042_));
 sg13g2_mux2_1 _1174_ (.A0(net123),
    .A1(net326),
    .S(_0520_),
    .X(_0043_));
 sg13g2_mux2_1 _1175_ (.A0(net121),
    .A1(net403),
    .S(_0520_),
    .X(_0044_));
 sg13g2_mux2_1 _1176_ (.A0(net119),
    .A1(net374),
    .S(_0520_),
    .X(_0045_));
 sg13g2_nand2_1 _1177_ (.Y(_0521_),
    .A(_0235_),
    .B(_0236_));
 sg13g2_inv_2 _1178_ (.Y(_0522_),
    .A(_0521_));
 sg13g2_nand2_2 _1179_ (.Y(_0523_),
    .A(_0519_),
    .B(_0522_));
 sg13g2_mux2_1 _1180_ (.A0(net134),
    .A1(net315),
    .S(_0523_),
    .X(_0046_));
 sg13g2_mux2_1 _1181_ (.A0(net132),
    .A1(net407),
    .S(_0523_),
    .X(_0047_));
 sg13g2_mux2_1 _1182_ (.A0(net130),
    .A1(net415),
    .S(_0523_),
    .X(_0048_));
 sg13g2_mux2_1 _1183_ (.A0(net126),
    .A1(net439),
    .S(_0523_),
    .X(_0049_));
 sg13g2_mux2_1 _1184_ (.A0(net128),
    .A1(net330),
    .S(_0523_),
    .X(_0050_));
 sg13g2_mux2_1 _1185_ (.A0(net124),
    .A1(net400),
    .S(_0523_),
    .X(_0051_));
 sg13g2_mux2_1 _1186_ (.A0(net122),
    .A1(net321),
    .S(_0523_),
    .X(_0052_));
 sg13g2_mux2_1 _1187_ (.A0(net120),
    .A1(net429),
    .S(_0523_),
    .X(_0053_));
 sg13g2_nand2b_2 _1188_ (.Y(_0524_),
    .B(_0511_),
    .A_N(_0234_));
 sg13g2_mux2_1 _1189_ (.A0(net133),
    .A1(net353),
    .S(_0524_),
    .X(_0054_));
 sg13g2_mux2_1 _1190_ (.A0(net131),
    .A1(net314),
    .S(_0524_),
    .X(_0055_));
 sg13g2_mux2_1 _1191_ (.A0(net129),
    .A1(net362),
    .S(_0524_),
    .X(_0056_));
 sg13g2_mux2_1 _1192_ (.A0(net125),
    .A1(net444),
    .S(_0524_),
    .X(_0057_));
 sg13g2_mux2_1 _1193_ (.A0(net127),
    .A1(net395),
    .S(_0524_),
    .X(_0058_));
 sg13g2_mux2_1 _1194_ (.A0(net123),
    .A1(net347),
    .S(_0524_),
    .X(_0059_));
 sg13g2_mux2_1 _1195_ (.A0(net121),
    .A1(net358),
    .S(_0524_),
    .X(_0060_));
 sg13g2_mux2_1 _1196_ (.A0(net119),
    .A1(net428),
    .S(_0524_),
    .X(_0061_));
 sg13g2_nand2b_2 _1197_ (.Y(_0525_),
    .B(_0522_),
    .A_N(_0513_));
 sg13g2_mux2_1 _1198_ (.A0(net134),
    .A1(net328),
    .S(net138),
    .X(_0062_));
 sg13g2_mux2_1 _1199_ (.A0(net132),
    .A1(net316),
    .S(net138),
    .X(_0063_));
 sg13g2_mux2_1 _1200_ (.A0(net130),
    .A1(net327),
    .S(net138),
    .X(_0064_));
 sg13g2_nor2_1 _1201_ (.A(net126),
    .B(net138),
    .Y(_0526_));
 sg13g2_a21oi_1 _1202_ (.A1(_0210_),
    .A2(_0525_),
    .Y(_0065_),
    .B1(_0526_));
 sg13g2_mux2_1 _1203_ (.A0(net128),
    .A1(net356),
    .S(net138),
    .X(_0066_));
 sg13g2_mux2_1 _1204_ (.A0(net124),
    .A1(net370),
    .S(net138),
    .X(_0067_));
 sg13g2_mux2_1 _1205_ (.A0(net122),
    .A1(net351),
    .S(net138),
    .X(_0068_));
 sg13g2_mux2_1 _1206_ (.A0(net120),
    .A1(net433),
    .S(net138),
    .X(_0069_));
 sg13g2_nand2_2 _1207_ (.Y(_0527_),
    .A(_0266_),
    .B(_0289_));
 sg13g2_nor4_1 _1208_ (.A(net148),
    .B(_0194_),
    .C(_0217_),
    .D(_0256_),
    .Y(_0528_));
 sg13g2_nor2_2 _1209_ (.A(_0527_),
    .B(_0528_),
    .Y(_0529_));
 sg13g2_or2_1 _1210_ (.X(_0530_),
    .B(_0528_),
    .A(_0527_));
 sg13g2_o21ai_1 _1211_ (.B1(net176),
    .Y(_0531_),
    .A1(net473),
    .A2(_0530_));
 sg13g2_a21oi_1 _1212_ (.A1(_0292_),
    .A2(_0530_),
    .Y(_0070_),
    .B1(_0531_));
 sg13g2_o21ai_1 _1213_ (.B1(net176),
    .Y(_0532_),
    .A1(net471),
    .A2(_0530_));
 sg13g2_a21oi_1 _1214_ (.A1(_0332_),
    .A2(_0530_),
    .Y(_0071_),
    .B1(_0532_));
 sg13g2_o21ai_1 _1215_ (.B1(net176),
    .Y(_0533_),
    .A1(net466),
    .A2(_0530_));
 sg13g2_a21oi_1 _1216_ (.A1(_0363_),
    .A2(_0530_),
    .Y(_0072_),
    .B1(_0533_));
 sg13g2_o21ai_1 _1217_ (.B1(net176),
    .Y(_0534_),
    .A1(net476),
    .A2(_0530_));
 sg13g2_a21oi_1 _1218_ (.A1(_0396_),
    .A2(_0530_),
    .Y(_0073_),
    .B1(_0534_));
 sg13g2_a22oi_1 _1219_ (.Y(_0535_),
    .B1(_0529_),
    .B2(net337),
    .A2(_0527_),
    .A1(_0416_));
 sg13g2_nor2_1 _1220_ (.A(net173),
    .B(_0535_),
    .Y(_0074_));
 sg13g2_a22oi_1 _1221_ (.Y(_0536_),
    .B1(_0529_),
    .B2(net457),
    .A2(_0527_),
    .A1(_0443_));
 sg13g2_nor2_1 _1222_ (.A(net173),
    .B(_0536_),
    .Y(_0075_));
 sg13g2_nand2b_1 _1223_ (.Y(_0537_),
    .B(_0527_),
    .A_N(_0472_));
 sg13g2_nand2_1 _1224_ (.Y(_0538_),
    .A(net437),
    .B(_0529_));
 sg13g2_a21oi_1 _1225_ (.A1(_0537_),
    .A2(_0538_),
    .Y(_0076_),
    .B1(net173));
 sg13g2_a22oi_1 _1226_ (.Y(_0539_),
    .B1(_0529_),
    .B2(net462),
    .A2(_0527_),
    .A1(_0502_));
 sg13g2_nor2_1 _1227_ (.A(net173),
    .B(_0539_),
    .Y(_0077_));
 sg13g2_nor2_2 _1228_ (.A(net172),
    .B(_0268_),
    .Y(_0540_));
 sg13g2_nand2_1 _1229_ (.Y(_0541_),
    .A(net284),
    .B(_0540_));
 sg13g2_o21ai_1 _1230_ (.B1(_0541_),
    .Y(_0078_),
    .A1(_0269_),
    .A2(_0292_));
 sg13g2_nand2_1 _1231_ (.Y(_0542_),
    .A(net286),
    .B(_0540_));
 sg13g2_o21ai_1 _1232_ (.B1(_0542_),
    .Y(_0079_),
    .A1(_0269_),
    .A2(_0332_));
 sg13g2_nand2_1 _1233_ (.Y(_0543_),
    .A(net280),
    .B(_0540_));
 sg13g2_o21ai_1 _1234_ (.B1(_0543_),
    .Y(_0080_),
    .A1(_0269_),
    .A2(_0363_));
 sg13g2_nand2_1 _1235_ (.Y(_0544_),
    .A(net282),
    .B(_0540_));
 sg13g2_o21ai_1 _1236_ (.B1(_0544_),
    .Y(_0081_),
    .A1(_0269_),
    .A2(_0396_));
 sg13g2_a22oi_1 _1237_ (.Y(_0545_),
    .B1(_0540_),
    .B2(net448),
    .A2(_0403_),
    .A1(_0268_));
 sg13g2_inv_1 _1238_ (.Y(_0082_),
    .A(_0545_));
 sg13g2_nand2_1 _1239_ (.Y(_0546_),
    .A(net453),
    .B(_0540_));
 sg13g2_o21ai_1 _1240_ (.B1(_0546_),
    .Y(_0083_),
    .A1(_0269_),
    .A2(_0442_));
 sg13g2_nand2_1 _1241_ (.Y(_0547_),
    .A(net450),
    .B(_0540_));
 sg13g2_o21ai_1 _1242_ (.B1(_0547_),
    .Y(_0084_),
    .A1(_0269_),
    .A2(_0472_));
 sg13g2_a22oi_1 _1243_ (.Y(_0548_),
    .B1(_0540_),
    .B2(net148),
    .A2(_0502_),
    .A1(_0268_));
 sg13g2_inv_1 _1244_ (.Y(_0085_),
    .A(_0548_));
 sg13g2_and3_2 _1245_ (.X(_0549_),
    .A(net175),
    .B(_0248_),
    .C(_0249_));
 sg13g2_nor2_1 _1246_ (.A(_0268_),
    .B(_0549_),
    .Y(_0550_));
 sg13g2_nand2b_1 _1247_ (.Y(_0551_),
    .B(_0268_),
    .A_N(net477));
 sg13g2_a22oi_1 _1248_ (.Y(_0552_),
    .B1(_0550_),
    .B2(net477),
    .A2(_0549_),
    .A1(_0293_));
 sg13g2_a21oi_1 _1249_ (.A1(_0551_),
    .A2(_0552_),
    .Y(_0090_),
    .B1(net172));
 sg13g2_nand2b_1 _1250_ (.Y(_0553_),
    .B(_0549_),
    .A_N(_0332_));
 sg13g2_xor2_1 _1251_ (.B(net477),
    .A(net480),
    .X(_0554_));
 sg13g2_a22oi_1 _1252_ (.Y(_0555_),
    .B1(_0554_),
    .B2(_0268_),
    .A2(_0550_),
    .A1(net480));
 sg13g2_a21oi_1 _1253_ (.A1(_0553_),
    .A2(_0555_),
    .Y(_0091_),
    .B1(net172));
 sg13g2_and3_1 _1254_ (.X(_0556_),
    .A(net480),
    .B(net477),
    .C(_0268_));
 sg13g2_or3_1 _1255_ (.A(net478),
    .B(_0549_),
    .C(_0556_),
    .X(_0557_));
 sg13g2_nand2_1 _1256_ (.Y(_0558_),
    .A(net478),
    .B(_0556_));
 sg13g2_nand3_1 _1257_ (.B(_0557_),
    .C(_0558_),
    .A(net175),
    .Y(_0559_));
 sg13g2_a21oi_1 _1258_ (.A1(_0363_),
    .A2(_0549_),
    .Y(_0092_),
    .B1(_0559_));
 sg13g2_xnor2_1 _1259_ (.Y(_0560_),
    .A(net472),
    .B(_0558_));
 sg13g2_nand2_1 _1260_ (.Y(_0561_),
    .A(_0396_),
    .B(_0549_));
 sg13g2_o21ai_1 _1261_ (.B1(_0561_),
    .Y(_0562_),
    .A1(_0549_),
    .A2(_0560_));
 sg13g2_nor2_1 _1262_ (.A(net172),
    .B(_0562_),
    .Y(_0093_));
 sg13g2_nor2_2 _1263_ (.A(net174),
    .B(_0185_),
    .Y(_0563_));
 sg13g2_nand2_1 _1264_ (.Y(_0564_),
    .A(net334),
    .B(_0563_));
 sg13g2_o21ai_1 _1265_ (.B1(_0564_),
    .Y(_0094_),
    .A1(net145),
    .A2(_0292_));
 sg13g2_nand2_1 _1266_ (.Y(_0565_),
    .A(net323),
    .B(_0563_));
 sg13g2_o21ai_1 _1267_ (.B1(_0565_),
    .Y(_0095_),
    .A1(net145),
    .A2(_0332_));
 sg13g2_nand2_1 _1268_ (.Y(_0566_),
    .A(net300),
    .B(_0563_));
 sg13g2_o21ai_1 _1269_ (.B1(_0566_),
    .Y(_0096_),
    .A1(_0220_),
    .A2(_0363_));
 sg13g2_nand2_1 _1270_ (.Y(_0567_),
    .A(net296),
    .B(_0563_));
 sg13g2_o21ai_1 _1271_ (.B1(_0567_),
    .Y(_0097_),
    .A1(_0220_),
    .A2(_0396_));
 sg13g2_a22oi_1 _1272_ (.Y(_0568_),
    .B1(_0563_),
    .B2(net449),
    .A2(_0416_),
    .A1(_0185_));
 sg13g2_inv_1 _1273_ (.Y(_0098_),
    .A(_0568_));
 sg13g2_nand2_1 _1274_ (.Y(_0569_),
    .A(net306),
    .B(_0563_));
 sg13g2_o21ai_1 _1275_ (.B1(_0569_),
    .Y(_0099_),
    .A1(net145),
    .A2(_0442_));
 sg13g2_nand2_1 _1276_ (.Y(_0570_),
    .A(net339),
    .B(_0563_));
 sg13g2_o21ai_1 _1277_ (.B1(_0570_),
    .Y(_0100_),
    .A1(net145),
    .A2(_0472_));
 sg13g2_a22oi_1 _1278_ (.Y(_0571_),
    .B1(_0563_),
    .B2(net446),
    .A2(_0502_),
    .A1(_0185_));
 sg13g2_inv_1 _1279_ (.Y(_0101_),
    .A(_0571_));
 sg13g2_nand3_1 _1280_ (.B(_0233_),
    .C(_0511_),
    .A(_0231_),
    .Y(_0572_));
 sg13g2_mux2_1 _1281_ (.A0(net133),
    .A1(net350),
    .S(_0572_),
    .X(_0102_));
 sg13g2_mux2_1 _1282_ (.A0(net131),
    .A1(net405),
    .S(_0572_),
    .X(_0103_));
 sg13g2_mux2_1 _1283_ (.A0(net129),
    .A1(net352),
    .S(_0572_),
    .X(_0104_));
 sg13g2_mux2_1 _1284_ (.A0(net125),
    .A1(net409),
    .S(_0572_),
    .X(_0105_));
 sg13g2_mux2_1 _1285_ (.A0(net127),
    .A1(net318),
    .S(_0572_),
    .X(_0106_));
 sg13g2_mux2_1 _1286_ (.A0(net123),
    .A1(net361),
    .S(_0572_),
    .X(_0107_));
 sg13g2_mux2_1 _1287_ (.A0(net121),
    .A1(net367),
    .S(_0572_),
    .X(_0108_));
 sg13g2_mux2_1 _1288_ (.A0(net119),
    .A1(net385),
    .S(_0572_),
    .X(_0109_));
 sg13g2_nor2b_2 _1289_ (.A(_0235_),
    .B_N(_0236_),
    .Y(_0573_));
 sg13g2_nand3_1 _1290_ (.B(_0233_),
    .C(_0573_),
    .A(_0231_),
    .Y(_0574_));
 sg13g2_mux2_1 _1291_ (.A0(net133),
    .A1(net422),
    .S(_0574_),
    .X(_0110_));
 sg13g2_mux2_1 _1292_ (.A0(net131),
    .A1(net313),
    .S(_0574_),
    .X(_0111_));
 sg13g2_mux2_1 _1293_ (.A0(net129),
    .A1(net441),
    .S(_0574_),
    .X(_0112_));
 sg13g2_mux2_1 _1294_ (.A0(net125),
    .A1(net331),
    .S(_0574_),
    .X(_0113_));
 sg13g2_mux2_1 _1295_ (.A0(net127),
    .A1(net412),
    .S(_0574_),
    .X(_0114_));
 sg13g2_mux2_1 _1296_ (.A0(net123),
    .A1(net379),
    .S(_0574_),
    .X(_0115_));
 sg13g2_mux2_1 _1297_ (.A0(net121),
    .A1(net420),
    .S(_0574_),
    .X(_0116_));
 sg13g2_mux2_1 _1298_ (.A0(net119),
    .A1(net349),
    .S(_0574_),
    .X(_0117_));
 sg13g2_nand2b_2 _1299_ (.Y(_0575_),
    .B(_0519_),
    .A_N(_0237_));
 sg13g2_mux2_1 _1300_ (.A0(net134),
    .A1(net414),
    .S(net137),
    .X(_0118_));
 sg13g2_nor2_1 _1301_ (.A(net132),
    .B(net137),
    .Y(_0576_));
 sg13g2_a21oi_1 _1302_ (.A1(_0205_),
    .A2(net137),
    .Y(_0119_),
    .B1(_0576_));
 sg13g2_mux2_1 _1303_ (.A0(net130),
    .A1(net445),
    .S(net137),
    .X(_0120_));
 sg13g2_mux2_1 _1304_ (.A0(net126),
    .A1(net432),
    .S(net137),
    .X(_0121_));
 sg13g2_mux2_1 _1305_ (.A0(net128),
    .A1(net424),
    .S(net137),
    .X(_0122_));
 sg13g2_mux2_1 _1306_ (.A0(net124),
    .A1(net338),
    .S(net137),
    .X(_0123_));
 sg13g2_mux2_1 _1307_ (.A0(net122),
    .A1(net377),
    .S(_0575_),
    .X(_0124_));
 sg13g2_mux2_1 _1308_ (.A0(net120),
    .A1(net354),
    .S(net137),
    .X(_0125_));
 sg13g2_nand2b_2 _1309_ (.Y(_0577_),
    .B(_0573_),
    .A_N(_0513_));
 sg13g2_mux2_1 _1310_ (.A0(net133),
    .A1(net411),
    .S(_0577_),
    .X(_0126_));
 sg13g2_mux2_1 _1311_ (.A0(net131),
    .A1(net320),
    .S(_0577_),
    .X(_0127_));
 sg13g2_mux2_1 _1312_ (.A0(net129),
    .A1(net348),
    .S(_0577_),
    .X(_0128_));
 sg13g2_mux2_1 _1313_ (.A0(net125),
    .A1(net426),
    .S(_0577_),
    .X(_0129_));
 sg13g2_mux2_1 _1314_ (.A0(net127),
    .A1(net387),
    .S(_0577_),
    .X(_0130_));
 sg13g2_mux2_1 _1315_ (.A0(net123),
    .A1(net324),
    .S(_0577_),
    .X(_0131_));
 sg13g2_mux2_1 _1316_ (.A0(net121),
    .A1(net378),
    .S(_0577_),
    .X(_0132_));
 sg13g2_mux2_1 _1317_ (.A0(net119),
    .A1(net364),
    .S(_0577_),
    .X(_0133_));
 sg13g2_nand2_2 _1318_ (.Y(_0578_),
    .A(_0519_),
    .B(_0573_));
 sg13g2_mux2_1 _1319_ (.A0(net133),
    .A1(net333),
    .S(_0578_),
    .X(_0134_));
 sg13g2_mux2_1 _1320_ (.A0(net131),
    .A1(net368),
    .S(_0578_),
    .X(_0135_));
 sg13g2_mux2_1 _1321_ (.A0(net129),
    .A1(net399),
    .S(_0578_),
    .X(_0136_));
 sg13g2_mux2_1 _1322_ (.A0(net125),
    .A1(net383),
    .S(_0578_),
    .X(_0137_));
 sg13g2_mux2_1 _1323_ (.A0(net127),
    .A1(net366),
    .S(_0578_),
    .X(_0138_));
 sg13g2_mux2_1 _1324_ (.A0(net123),
    .A1(net389),
    .S(_0578_),
    .X(_0139_));
 sg13g2_mux2_1 _1325_ (.A0(net121),
    .A1(net427),
    .S(_0578_),
    .X(_0140_));
 sg13g2_mux2_1 _1326_ (.A0(net119),
    .A1(net375),
    .S(_0578_),
    .X(_0141_));
 sg13g2_nand2b_2 _1327_ (.Y(_0579_),
    .B(_0522_),
    .A_N(_0517_));
 sg13g2_mux2_1 _1328_ (.A0(net134),
    .A1(net425),
    .S(net136),
    .X(_0142_));
 sg13g2_mux2_1 _1329_ (.A0(net132),
    .A1(net384),
    .S(net136),
    .X(_0143_));
 sg13g2_nor2_1 _1330_ (.A(net130),
    .B(net136),
    .Y(_0580_));
 sg13g2_a21oi_1 _1331_ (.A1(_0207_),
    .A2(net136),
    .Y(_0144_),
    .B1(_0580_));
 sg13g2_mux2_1 _1332_ (.A0(net126),
    .A1(net380),
    .S(_0579_),
    .X(_0145_));
 sg13g2_mux2_1 _1333_ (.A0(net128),
    .A1(net408),
    .S(net136),
    .X(_0146_));
 sg13g2_mux2_1 _1334_ (.A0(net124),
    .A1(net319),
    .S(net136),
    .X(_0147_));
 sg13g2_mux2_1 _1335_ (.A0(net122),
    .A1(net401),
    .S(net136),
    .X(_0148_));
 sg13g2_mux2_1 _1336_ (.A0(net120),
    .A1(net369),
    .S(net136),
    .X(_0149_));
 sg13g2_nand2b_2 _1337_ (.Y(_0581_),
    .B(_0573_),
    .A_N(_0234_));
 sg13g2_mux2_1 _1338_ (.A0(net133),
    .A1(net373),
    .S(_0581_),
    .X(_0150_));
 sg13g2_mux2_1 _1339_ (.A0(net131),
    .A1(net398),
    .S(_0581_),
    .X(_0151_));
 sg13g2_mux2_1 _1340_ (.A0(net129),
    .A1(net431),
    .S(_0581_),
    .X(_0152_));
 sg13g2_mux2_1 _1341_ (.A0(net125),
    .A1(net382),
    .S(_0581_),
    .X(_0153_));
 sg13g2_mux2_1 _1342_ (.A0(net127),
    .A1(net438),
    .S(_0581_),
    .X(_0154_));
 sg13g2_mux2_1 _1343_ (.A0(net123),
    .A1(net419),
    .S(_0581_),
    .X(_0155_));
 sg13g2_mux2_1 _1344_ (.A0(net121),
    .A1(net443),
    .S(_0581_),
    .X(_0156_));
 sg13g2_mux2_1 _1345_ (.A0(net119),
    .A1(net325),
    .S(_0581_),
    .X(_0157_));
 sg13g2_nor2_2 _1346_ (.A(net174),
    .B(_0265_),
    .Y(_0582_));
 sg13g2_nand2_1 _1347_ (.Y(_0583_),
    .A(net311),
    .B(_0582_));
 sg13g2_o21ai_1 _1348_ (.B1(_0583_),
    .Y(_0158_),
    .A1(net141),
    .A2(_0292_));
 sg13g2_nand2_1 _1349_ (.Y(_0584_),
    .A(net298),
    .B(_0582_));
 sg13g2_o21ai_1 _1350_ (.B1(_0584_),
    .Y(_0159_),
    .A1(net141),
    .A2(_0332_));
 sg13g2_nand2_1 _1351_ (.Y(_0585_),
    .A(net309),
    .B(_0582_));
 sg13g2_o21ai_1 _1352_ (.B1(_0585_),
    .Y(_0160_),
    .A1(net141),
    .A2(_0363_));
 sg13g2_nand2_1 _1353_ (.Y(_0586_),
    .A(net302),
    .B(_0582_));
 sg13g2_o21ai_1 _1354_ (.B1(_0586_),
    .Y(_0161_),
    .A1(_0264_),
    .A2(_0396_));
 sg13g2_a22oi_1 _1355_ (.Y(_0587_),
    .B1(_0582_),
    .B2(net447),
    .A2(_0403_),
    .A1(_0265_));
 sg13g2_inv_1 _1356_ (.Y(_0162_),
    .A(_0587_));
 sg13g2_nand2_1 _1357_ (.Y(_0588_),
    .A(net307),
    .B(_0582_));
 sg13g2_o21ai_1 _1358_ (.B1(_0588_),
    .Y(_0163_),
    .A1(net141),
    .A2(_0442_));
 sg13g2_nand2_1 _1359_ (.Y(_0589_),
    .A(net294),
    .B(_0582_));
 sg13g2_o21ai_1 _1360_ (.B1(_0589_),
    .Y(_0164_),
    .A1(net141),
    .A2(_0472_));
 sg13g2_a22oi_1 _1361_ (.Y(_0590_),
    .B1(_0582_),
    .B2(net452),
    .A2(_0502_),
    .A1(_0265_));
 sg13g2_inv_1 _1362_ (.Y(_0165_),
    .A(_0590_));
 sg13g2_or2_1 _1363_ (.X(_0591_),
    .B(_0296_),
    .A(_0287_));
 sg13g2_inv_1 _1364_ (.Y(_0592_),
    .A(_0591_));
 sg13g2_nor2_1 _1365_ (.A(_0285_),
    .B(_0592_),
    .Y(_0593_));
 sg13g2_nand4_1 _1366_ (.B(_0425_),
    .C(_0448_),
    .A(_0405_),
    .Y(_0594_),
    .D(_0593_));
 sg13g2_nor3_1 _1367_ (.A(_0304_),
    .B(_0479_),
    .C(_0594_),
    .Y(_0595_));
 sg13g2_a21o_1 _1368_ (.A2(_0592_),
    .A1(net481),
    .B1(_0595_),
    .X(_0596_));
 sg13g2_and2_1 _1369_ (.A(net175),
    .B(_0596_),
    .X(_0166_));
 sg13g2_o21ai_1 _1370_ (.B1(_0299_),
    .Y(_0597_),
    .A1(net452),
    .A2(_0476_));
 sg13g2_nand3_1 _1371_ (.B(_0450_),
    .C(_0478_),
    .A(_0447_),
    .Y(_0598_));
 sg13g2_o21ai_1 _1372_ (.B1(_0598_),
    .Y(_0599_),
    .A1(\cpu0.a_reg[7] ),
    .A2(_0477_));
 sg13g2_xor2_1 _1373_ (.B(_0599_),
    .A(_0597_),
    .X(_0600_));
 sg13g2_o21ai_1 _1374_ (.B1(net175),
    .Y(_0601_),
    .A1(net458),
    .A2(_0591_));
 sg13g2_a21oi_1 _1375_ (.A1(_0591_),
    .A2(_0600_),
    .Y(_0167_),
    .B1(_0601_));
 sg13g2_nand2b_2 _1376_ (.Y(_0602_),
    .B(_0522_),
    .A_N(_0234_));
 sg13g2_mux2_1 _1377_ (.A0(net134),
    .A1(net417),
    .S(net135),
    .X(_0168_));
 sg13g2_nor2_1 _1378_ (.A(net132),
    .B(net135),
    .Y(_0603_));
 sg13g2_a21oi_1 _1379_ (.A1(_0206_),
    .A2(net135),
    .Y(_0169_),
    .B1(_0603_));
 sg13g2_mux2_1 _1380_ (.A0(net130),
    .A1(net340),
    .S(net135),
    .X(_0170_));
 sg13g2_mux2_1 _1381_ (.A0(net126),
    .A1(net386),
    .S(_0602_),
    .X(_0171_));
 sg13g2_mux2_1 _1382_ (.A0(net128),
    .A1(net357),
    .S(net135),
    .X(_0172_));
 sg13g2_mux2_1 _1383_ (.A0(net124),
    .A1(net418),
    .S(net135),
    .X(_0173_));
 sg13g2_mux2_1 _1384_ (.A0(net122),
    .A1(net332),
    .S(net135),
    .X(_0174_));
 sg13g2_mux2_1 _1385_ (.A0(net120),
    .A1(net346),
    .S(net135),
    .X(_0175_));
 sg13g2_mux4_1 _1386_ (.S0(\uart0.bit_counter[0] ),
    .A0(uo_out[4]),
    .A1(uo_out[5]),
    .A2(uo_out[6]),
    .A3(uo_out[7]),
    .S1(\uart0.bit_counter[1] ),
    .X(_0604_));
 sg13g2_mux4_1 _1387_ (.S0(\uart0.bit_counter[0] ),
    .A0(uo_out[0]),
    .A1(uo_out[1]),
    .A2(uo_out[2]),
    .A3(uo_out[3]),
    .S1(\uart0.bit_counter[1] ),
    .X(_0605_));
 sg13g2_a21o_1 _1388_ (.A2(_0605_),
    .A1(_0192_),
    .B1(_0201_),
    .X(_0606_));
 sg13g2_a21oi_1 _1389_ (.A1(net434),
    .A2(_0604_),
    .Y(_0607_),
    .B1(_0606_));
 sg13g2_nor3_1 _1390_ (.A(\uart0.tx ),
    .B(\uart0.uart_state[1] ),
    .C(net304),
    .Y(_0608_));
 sg13g2_or3_1 _1391_ (.A(net292),
    .B(_0607_),
    .C(_0608_),
    .X(_0609_));
 sg13g2_nand3_1 _1392_ (.B(_0202_),
    .C(_0609_),
    .A(net178),
    .Y(_0176_));
 sg13g2_or2_1 _1393_ (.X(_0610_),
    .B(_0513_),
    .A(_0237_));
 sg13g2_mux2_1 _1394_ (.A0(net134),
    .A1(net381),
    .S(_0610_),
    .X(_0177_));
 sg13g2_mux2_1 _1395_ (.A0(net132),
    .A1(net423),
    .S(_0610_),
    .X(_0178_));
 sg13g2_mux2_1 _1396_ (.A0(net130),
    .A1(net396),
    .S(_0610_),
    .X(_0179_));
 sg13g2_mux2_1 _1397_ (.A0(net126),
    .A1(net341),
    .S(_0610_),
    .X(_0180_));
 sg13g2_mux2_1 _1398_ (.A0(net128),
    .A1(net344),
    .S(_0610_),
    .X(_0181_));
 sg13g2_mux2_1 _1399_ (.A0(net124),
    .A1(net406),
    .S(_0610_),
    .X(_0182_));
 sg13g2_mux2_1 _1400_ (.A0(net122),
    .A1(net393),
    .S(_0610_),
    .X(_0183_));
 sg13g2_mux2_1 _1401_ (.A0(net120),
    .A1(net410),
    .S(_0610_),
    .X(_0184_));
 sg13g2_nor3_1 _1402_ (.A(net292),
    .B(_0201_),
    .C(net455),
    .Y(_0611_));
 sg13g2_or2_1 _1403_ (.X(_0612_),
    .B(_0611_),
    .A(net483));
 sg13g2_nand2_1 _1404_ (.Y(_0613_),
    .A(net483),
    .B(_0611_));
 sg13g2_and3_1 _1405_ (.X(_0186_),
    .A(net178),
    .B(_0612_),
    .C(_0613_));
 sg13g2_nand2b_1 _1406_ (.Y(_0614_),
    .B(net484),
    .A_N(net460));
 sg13g2_nand3_1 _1407_ (.B(\uart0.bit_counter[0] ),
    .C(_0611_),
    .A(net460),
    .Y(_0615_));
 sg13g2_and3_1 _1408_ (.X(_0187_),
    .A(net178),
    .B(_0614_),
    .C(net461));
 sg13g2_o21ai_1 _1409_ (.B1(net178),
    .Y(_0616_),
    .A1(_0192_),
    .A2(net461));
 sg13g2_a21oi_1 _1410_ (.A1(_0192_),
    .A2(net461),
    .Y(_0188_),
    .B1(_0616_));
 sg13g2_nor2_1 _1411_ (.A(_0191_),
    .B(_0616_),
    .Y(_0189_));
 sg13g2_nor3_1 _1412_ (.A(net173),
    .B(_0213_),
    .C(net469),
    .Y(_0190_));
 sg13g2_a21oi_1 _1413_ (.A1(_0292_),
    .A2(net139),
    .Y(_0086_),
    .B1(_0507_));
 sg13g2_a21oi_1 _1414_ (.A1(_0332_),
    .A2(net139),
    .Y(_0087_),
    .B1(_0508_));
 sg13g2_a21oi_1 _1415_ (.A1(_0363_),
    .A2(net139),
    .Y(_0088_),
    .B1(_0509_));
 sg13g2_a21oi_1 _1416_ (.A1(_0396_),
    .A2(net140),
    .Y(_0089_),
    .B1(_0510_));
 sg13g2_dfrbpq_1 _1417_ (.RESET_B(net50),
    .D(_0008_),
    .Q(\cpu0.ram[5][0] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1418_ (.RESET_B(net232),
    .D(_0009_),
    .Q(\cpu0.ram[5][1] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1419_ (.RESET_B(net231),
    .D(_0010_),
    .Q(\cpu0.ram[5][2] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1420_ (.RESET_B(net230),
    .D(_0011_),
    .Q(\cpu0.ram[5][3] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1421_ (.RESET_B(net229),
    .D(_0012_),
    .Q(\cpu0.ram[5][4] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1422_ (.RESET_B(net228),
    .D(_0013_),
    .Q(\cpu0.ram[5][5] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1423_ (.RESET_B(net227),
    .D(_0014_),
    .Q(\cpu0.ram[5][6] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1424_ (.RESET_B(net226),
    .D(_0015_),
    .Q(\cpu0.ram[5][7] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 _1425_ (.RESET_B(net225),
    .D(_0016_),
    .Q(_0000_),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 _1426_ (.RESET_B(net224),
    .D(_0017_),
    .Q(_0001_),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 _1427_ (.RESET_B(net223),
    .D(_0018_),
    .Q(_0002_),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1428_ (.RESET_B(net222),
    .D(_0019_),
    .Q(_0003_),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1429_ (.RESET_B(net221),
    .D(_0020_),
    .Q(\cpu0.ram[2][0] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1430_ (.RESET_B(net220),
    .D(_0021_),
    .Q(\cpu0.ram[2][1] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1431_ (.RESET_B(net219),
    .D(_0022_),
    .Q(\cpu0.ram[2][2] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1432_ (.RESET_B(net218),
    .D(_0023_),
    .Q(\cpu0.ram[2][3] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1433_ (.RESET_B(net217),
    .D(_0024_),
    .Q(\cpu0.ram[2][4] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1434_ (.RESET_B(net216),
    .D(_0025_),
    .Q(\cpu0.ram[2][5] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1435_ (.RESET_B(net215),
    .D(_0026_),
    .Q(\cpu0.ram[2][6] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1436_ (.RESET_B(net214),
    .D(_0027_),
    .Q(\cpu0.ram[2][7] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _1437_ (.RESET_B(net213),
    .D(_0028_),
    .Q(\cpu0.step[1] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _1438_ (.RESET_B(net51),
    .D(net465),
    .Q(\cpu0.step[2] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1439_ (.RESET_B(net52),
    .D(net305),
    .Q(\uart0.uart_state[0] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1440_ (.RESET_B(net53),
    .D(_0007_),
    .Q(\uart0.uart_state[1] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1441_ (.RESET_B(net80),
    .D(net277),
    .Q(\uart0.uart_state[2] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1442_ (.RESET_B(net212),
    .D(net436),
    .Q(\uart0.uart_state[3] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1443_ (.RESET_B(net211),
    .D(_0030_),
    .Q(\cpu0.ram[4][0] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1444_ (.RESET_B(net210),
    .D(_0031_),
    .Q(\cpu0.ram[4][1] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1445_ (.RESET_B(net209),
    .D(_0032_),
    .Q(\cpu0.ram[4][2] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1446_ (.RESET_B(net208),
    .D(_0033_),
    .Q(\cpu0.ram[4][3] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1447_ (.RESET_B(net207),
    .D(_0034_),
    .Q(\cpu0.ram[4][4] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1448_ (.RESET_B(net206),
    .D(_0035_),
    .Q(\cpu0.ram[4][5] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1449_ (.RESET_B(net205),
    .D(_0036_),
    .Q(\cpu0.ram[4][6] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1450_ (.RESET_B(net204),
    .D(_0037_),
    .Q(\cpu0.ram[4][7] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1451_ (.RESET_B(net203),
    .D(_0038_),
    .Q(\cpu0.ram[3][0] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1452_ (.RESET_B(net202),
    .D(_0039_),
    .Q(\cpu0.ram[3][1] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1453_ (.RESET_B(net201),
    .D(_0040_),
    .Q(\cpu0.ram[3][2] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1454_ (.RESET_B(net200),
    .D(_0041_),
    .Q(\cpu0.ram[3][3] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1455_ (.RESET_B(net199),
    .D(_0042_),
    .Q(\cpu0.ram[3][4] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1456_ (.RESET_B(net198),
    .D(_0043_),
    .Q(\cpu0.ram[3][5] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1457_ (.RESET_B(net197),
    .D(_0044_),
    .Q(\cpu0.ram[3][6] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1458_ (.RESET_B(net196),
    .D(_0045_),
    .Q(\cpu0.ram[3][7] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1459_ (.RESET_B(net195),
    .D(_0046_),
    .Q(\cpu0.ram[15][0] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1460_ (.RESET_B(net194),
    .D(_0047_),
    .Q(\cpu0.ram[15][1] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1461_ (.RESET_B(net193),
    .D(_0048_),
    .Q(\cpu0.ram[15][2] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1462_ (.RESET_B(net192),
    .D(_0049_),
    .Q(\cpu0.ram[15][3] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1463_ (.RESET_B(net191),
    .D(_0050_),
    .Q(\cpu0.ram[15][4] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1464_ (.RESET_B(net190),
    .D(_0051_),
    .Q(\cpu0.ram[15][5] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1465_ (.RESET_B(net189),
    .D(_0052_),
    .Q(\cpu0.ram[15][6] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1466_ (.RESET_B(net188),
    .D(_0053_),
    .Q(\cpu0.ram[15][7] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1467_ (.RESET_B(net187),
    .D(_0054_),
    .Q(\cpu0.ram[1][0] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1468_ (.RESET_B(net186),
    .D(_0055_),
    .Q(\cpu0.ram[1][1] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1469_ (.RESET_B(net185),
    .D(_0056_),
    .Q(\cpu0.ram[1][2] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1470_ (.RESET_B(net184),
    .D(_0057_),
    .Q(\cpu0.ram[1][3] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1471_ (.RESET_B(net183),
    .D(_0058_),
    .Q(\cpu0.ram[1][4] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1472_ (.RESET_B(net182),
    .D(_0059_),
    .Q(\cpu0.ram[1][5] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1473_ (.RESET_B(net181),
    .D(_0060_),
    .Q(\cpu0.ram[1][6] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1474_ (.RESET_B(net180),
    .D(_0061_),
    .Q(\cpu0.ram[1][7] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1475_ (.RESET_B(net179),
    .D(_0062_),
    .Q(\cpu0.ram[14][0] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1476_ (.RESET_B(net118),
    .D(_0063_),
    .Q(\cpu0.ram[14][1] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1477_ (.RESET_B(net117),
    .D(_0064_),
    .Q(\cpu0.ram[14][2] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1478_ (.RESET_B(net116),
    .D(_0065_),
    .Q(\cpu0.ram[14][3] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1479_ (.RESET_B(net115),
    .D(_0066_),
    .Q(\cpu0.ram[14][4] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1480_ (.RESET_B(net114),
    .D(_0067_),
    .Q(\cpu0.ram[14][5] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1481_ (.RESET_B(net113),
    .D(_0068_),
    .Q(\cpu0.ram[14][6] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1482_ (.RESET_B(net112),
    .D(_0069_),
    .Q(\cpu0.ram[14][7] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _1483_ (.RESET_B(net111),
    .D(net474),
    .Q(\cpu0.a_reg[0] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _1484_ (.RESET_B(net109),
    .D(_0071_),
    .Q(\cpu0.a_reg[1] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_2 _1485_ (.RESET_B(net107),
    .D(_0072_),
    .Q(\cpu0.a_reg[2] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _1486_ (.RESET_B(net105),
    .D(_0073_),
    .Q(\cpu0.a_reg[3] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1487_ (.RESET_B(net103),
    .D(_0074_),
    .Q(\cpu0.a_reg[4] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 _1488_ (.RESET_B(net101),
    .D(_0075_),
    .Q(\cpu0.a_reg[5] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 _1489_ (.RESET_B(net99),
    .D(_0076_),
    .Q(\cpu0.a_reg[6] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 _1490_ (.RESET_B(net97),
    .D(_0077_),
    .Q(\cpu0.a_reg[7] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1491_ (.RESET_B(net95),
    .D(net285),
    .Q(\cpu0.ir[0] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1492_ (.RESET_B(net93),
    .D(net287),
    .Q(\cpu0.ir[1] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1493_ (.RESET_B(net91),
    .D(net281),
    .Q(\cpu0.ir[2] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1494_ (.RESET_B(net89),
    .D(net283),
    .Q(\cpu0.ir[3] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 _1495_ (.RESET_B(net87),
    .D(_0082_),
    .Q(\cpu0.ir[4] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _1496_ (.RESET_B(net85),
    .D(net454),
    .Q(\cpu0.ir[5] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _1497_ (.RESET_B(net83),
    .D(net451),
    .Q(\cpu0.ir[6] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1498_ (.RESET_B(net81),
    .D(_0085_),
    .Q(\cpu0.ir[7] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _1499_ (.RESET_B(net79),
    .D(_0086_),
    .Q(\cpu0.mar[0] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1500_ (.RESET_B(net77),
    .D(_0087_),
    .Q(\cpu0.mar[1] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1501_ (.RESET_B(net75),
    .D(_0088_),
    .Q(\cpu0.mar[2] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1502_ (.RESET_B(net73),
    .D(_0089_),
    .Q(\cpu0.mar[3] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 _1503_ (.RESET_B(net71),
    .D(_0090_),
    .Q(\cpu0.pc[0] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _1504_ (.RESET_B(net69),
    .D(_0091_),
    .Q(\cpu0.pc[1] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1505_ (.RESET_B(net67),
    .D(_0092_),
    .Q(\cpu0.pc[2] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1506_ (.RESET_B(net65),
    .D(_0093_),
    .Q(\cpu0.pc[3] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _1507_ (.RESET_B(net63),
    .D(net335),
    .Q(uo_out[0]),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _1508_ (.RESET_B(net61),
    .D(_0095_),
    .Q(uo_out[1]),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _1509_ (.RESET_B(net59),
    .D(net301),
    .Q(uo_out[2]),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _1510_ (.RESET_B(net57),
    .D(net297),
    .Q(uo_out[3]),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _1511_ (.RESET_B(net55),
    .D(_0098_),
    .Q(uo_out[4]),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 _1512_ (.RESET_B(net49),
    .D(_0099_),
    .Q(uo_out[5]),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 _1513_ (.RESET_B(net47),
    .D(_0100_),
    .Q(uo_out[6]),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _1514_ (.RESET_B(net45),
    .D(_0101_),
    .Q(uo_out[7]),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1515_ (.RESET_B(net43),
    .D(_0102_),
    .Q(\cpu0.ram[0][0] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1516_ (.RESET_B(net42),
    .D(_0103_),
    .Q(\cpu0.ram[0][1] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1517_ (.RESET_B(net41),
    .D(_0104_),
    .Q(\cpu0.ram[0][2] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1518_ (.RESET_B(net40),
    .D(_0105_),
    .Q(\cpu0.ram[0][3] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1519_ (.RESET_B(net39),
    .D(_0106_),
    .Q(\cpu0.ram[0][4] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1520_ (.RESET_B(net38),
    .D(_0107_),
    .Q(\cpu0.ram[0][5] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1521_ (.RESET_B(net37),
    .D(_0108_),
    .Q(\cpu0.ram[0][6] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1522_ (.RESET_B(net36),
    .D(_0109_),
    .Q(\cpu0.ram[0][7] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1523_ (.RESET_B(net35),
    .D(_0110_),
    .Q(\cpu0.ram[8][0] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1524_ (.RESET_B(net34),
    .D(_0111_),
    .Q(\cpu0.ram[8][1] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1525_ (.RESET_B(net33),
    .D(_0112_),
    .Q(\cpu0.ram[8][2] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1526_ (.RESET_B(net32),
    .D(_0113_),
    .Q(\cpu0.ram[8][3] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1527_ (.RESET_B(net31),
    .D(_0114_),
    .Q(\cpu0.ram[8][4] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1528_ (.RESET_B(net30),
    .D(_0115_),
    .Q(\cpu0.ram[8][5] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1529_ (.RESET_B(net29),
    .D(_0116_),
    .Q(\cpu0.ram[8][6] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1530_ (.RESET_B(net28),
    .D(_0117_),
    .Q(\cpu0.ram[8][7] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1531_ (.RESET_B(net274),
    .D(_0118_),
    .Q(\cpu0.ram[7][0] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1532_ (.RESET_B(net273),
    .D(_0119_),
    .Q(\cpu0.ram[7][1] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1533_ (.RESET_B(net272),
    .D(_0120_),
    .Q(\cpu0.ram[7][2] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1534_ (.RESET_B(net271),
    .D(_0121_),
    .Q(\cpu0.ram[7][3] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1535_ (.RESET_B(net270),
    .D(_0122_),
    .Q(\cpu0.ram[7][4] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1536_ (.RESET_B(net269),
    .D(_0123_),
    .Q(\cpu0.ram[7][5] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1537_ (.RESET_B(net268),
    .D(_0124_),
    .Q(\cpu0.ram[7][6] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1538_ (.RESET_B(net267),
    .D(_0125_),
    .Q(\cpu0.ram[7][7] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1539_ (.RESET_B(net266),
    .D(_0126_),
    .Q(\cpu0.ram[10][0] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1540_ (.RESET_B(net265),
    .D(_0127_),
    .Q(\cpu0.ram[10][1] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1541_ (.RESET_B(net264),
    .D(_0128_),
    .Q(\cpu0.ram[10][2] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1542_ (.RESET_B(net263),
    .D(_0129_),
    .Q(\cpu0.ram[10][3] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1543_ (.RESET_B(net262),
    .D(_0130_),
    .Q(\cpu0.ram[10][4] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1544_ (.RESET_B(net261),
    .D(_0131_),
    .Q(\cpu0.ram[10][5] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1545_ (.RESET_B(net260),
    .D(_0132_),
    .Q(\cpu0.ram[10][6] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1546_ (.RESET_B(net259),
    .D(_0133_),
    .Q(\cpu0.ram[10][7] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1547_ (.RESET_B(net258),
    .D(_0134_),
    .Q(\cpu0.ram[11][0] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1548_ (.RESET_B(net257),
    .D(_0135_),
    .Q(\cpu0.ram[11][1] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1549_ (.RESET_B(net256),
    .D(_0136_),
    .Q(\cpu0.ram[11][2] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1550_ (.RESET_B(net255),
    .D(_0137_),
    .Q(\cpu0.ram[11][3] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1551_ (.RESET_B(net254),
    .D(_0138_),
    .Q(\cpu0.ram[11][4] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1552_ (.RESET_B(net253),
    .D(_0139_),
    .Q(\cpu0.ram[11][5] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1553_ (.RESET_B(net252),
    .D(_0140_),
    .Q(\cpu0.ram[11][6] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1554_ (.RESET_B(net251),
    .D(_0141_),
    .Q(\cpu0.ram[11][7] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1555_ (.RESET_B(net250),
    .D(_0142_),
    .Q(\cpu0.ram[12][0] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1556_ (.RESET_B(net249),
    .D(_0143_),
    .Q(\cpu0.ram[12][1] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1557_ (.RESET_B(net248),
    .D(_0144_),
    .Q(\cpu0.ram[12][2] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1558_ (.RESET_B(net247),
    .D(_0145_),
    .Q(\cpu0.ram[12][3] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1559_ (.RESET_B(net246),
    .D(_0146_),
    .Q(\cpu0.ram[12][4] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1560_ (.RESET_B(net245),
    .D(_0147_),
    .Q(\cpu0.ram[12][5] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1561_ (.RESET_B(net244),
    .D(_0148_),
    .Q(\cpu0.ram[12][6] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1562_ (.RESET_B(net243),
    .D(_0149_),
    .Q(\cpu0.ram[12][7] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1563_ (.RESET_B(net242),
    .D(_0150_),
    .Q(\cpu0.ram[9][0] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1564_ (.RESET_B(net241),
    .D(_0151_),
    .Q(\cpu0.ram[9][1] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1565_ (.RESET_B(net240),
    .D(_0152_),
    .Q(\cpu0.ram[9][2] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1566_ (.RESET_B(net239),
    .D(_0153_),
    .Q(\cpu0.ram[9][3] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1567_ (.RESET_B(net238),
    .D(_0154_),
    .Q(\cpu0.ram[9][4] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1568_ (.RESET_B(net237),
    .D(_0155_),
    .Q(\cpu0.ram[9][5] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1569_ (.RESET_B(net236),
    .D(_0156_),
    .Q(\cpu0.ram[9][6] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1570_ (.RESET_B(net235),
    .D(_0157_),
    .Q(\cpu0.ram[9][7] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_2 _1571_ (.RESET_B(net234),
    .D(net312),
    .Q(\cpu0.b_reg[0] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _1572_ (.RESET_B(net110),
    .D(net299),
    .Q(\cpu0.b_reg[1] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1573_ (.RESET_B(net106),
    .D(net310),
    .Q(\cpu0.b_reg[2] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1574_ (.RESET_B(net102),
    .D(net303),
    .Q(\cpu0.b_reg[3] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1575_ (.RESET_B(net98),
    .D(_0162_),
    .Q(\cpu0.b_reg[4] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1576_ (.RESET_B(net94),
    .D(net308),
    .Q(\cpu0.b_reg[5] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1577_ (.RESET_B(net90),
    .D(net295),
    .Q(\cpu0.b_reg[6] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1578_ (.RESET_B(net86),
    .D(_0165_),
    .Q(\cpu0.b_reg[7] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1579_ (.RESET_B(net82),
    .D(_0166_),
    .Q(\cpu0.zero_flag ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1580_ (.RESET_B(net78),
    .D(net459),
    .Q(\cpu0.carry_flag ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1581_ (.RESET_B(net74),
    .D(_0168_),
    .Q(\cpu0.ram[13][0] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1582_ (.RESET_B(net72),
    .D(_0169_),
    .Q(\cpu0.ram[13][1] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1583_ (.RESET_B(net70),
    .D(_0170_),
    .Q(\cpu0.ram[13][2] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1584_ (.RESET_B(net68),
    .D(_0171_),
    .Q(\cpu0.ram[13][3] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1585_ (.RESET_B(net66),
    .D(_0172_),
    .Q(\cpu0.ram[13][4] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1586_ (.RESET_B(net64),
    .D(_0173_),
    .Q(\cpu0.ram[13][5] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1587_ (.RESET_B(net62),
    .D(_0174_),
    .Q(\cpu0.ram[13][6] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1588_ (.RESET_B(net60),
    .D(_0175_),
    .Q(\cpu0.ram[13][7] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1589_ (.RESET_B(net58),
    .D(net456),
    .Q(\uart0.tx ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1590_ (.RESET_B(net54),
    .D(_0177_),
    .Q(\cpu0.ram[6][0] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1591_ (.RESET_B(net48),
    .D(_0178_),
    .Q(\cpu0.ram[6][1] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1592_ (.RESET_B(net46),
    .D(_0179_),
    .Q(\cpu0.ram[6][2] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1593_ (.RESET_B(net44),
    .D(_0180_),
    .Q(\cpu0.ram[6][3] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1594_ (.RESET_B(net233),
    .D(_0181_),
    .Q(\cpu0.ram[6][4] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1595_ (.RESET_B(net108),
    .D(_0182_),
    .Q(\cpu0.ram[6][5] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1596_ (.RESET_B(net104),
    .D(_0183_),
    .Q(\cpu0.ram[6][6] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1597_ (.RESET_B(net100),
    .D(_0184_),
    .Q(\cpu0.ram[6][7] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1598_ (.RESET_B(net96),
    .D(_0185_),
    .Q(\uart0.tx_en_prev ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_2 _1599_ (.RESET_B(net92),
    .D(_0186_),
    .Q(\uart0.bit_counter[0] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_2 _1600_ (.RESET_B(net84),
    .D(_0187_),
    .Q(\uart0.bit_counter[1] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1601_ (.RESET_B(net76),
    .D(_0188_),
    .Q(\uart0.bit_counter[2] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1602_ (.RESET_B(net88),
    .D(net279),
    .Q(\uart0.bit_counter[3] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _1603_ (.RESET_B(net56),
    .D(net470),
    .Q(\cpu0.step[0] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_tiehi _1529__29 (.L_HI(net29));
 sg13g2_tiehi _1528__30 (.L_HI(net30));
 sg13g2_tiehi _1527__31 (.L_HI(net31));
 sg13g2_tiehi _1526__32 (.L_HI(net32));
 sg13g2_tiehi _1525__33 (.L_HI(net33));
 sg13g2_tiehi _1524__34 (.L_HI(net34));
 sg13g2_tiehi _1523__35 (.L_HI(net35));
 sg13g2_tiehi _1522__36 (.L_HI(net36));
 sg13g2_tiehi _1521__37 (.L_HI(net37));
 sg13g2_tiehi _1520__38 (.L_HI(net38));
 sg13g2_tiehi _1519__39 (.L_HI(net39));
 sg13g2_tiehi _1518__40 (.L_HI(net40));
 sg13g2_tiehi _1517__41 (.L_HI(net41));
 sg13g2_tiehi _1516__42 (.L_HI(net42));
 sg13g2_tiehi _1515__43 (.L_HI(net43));
 sg13g2_tiehi _1593__44 (.L_HI(net44));
 sg13g2_tiehi _1514__45 (.L_HI(net45));
 sg13g2_tiehi _1592__46 (.L_HI(net46));
 sg13g2_tiehi _1513__47 (.L_HI(net47));
 sg13g2_tiehi _1591__48 (.L_HI(net48));
 sg13g2_tiehi _1512__49 (.L_HI(net49));
 sg13g2_tiehi _1417__50 (.L_HI(net50));
 sg13g2_tiehi _1438__51 (.L_HI(net51));
 sg13g2_tiehi _1439__52 (.L_HI(net52));
 sg13g2_tiehi _1440__53 (.L_HI(net53));
 sg13g2_tiehi _1590__54 (.L_HI(net54));
 sg13g2_tiehi _1511__55 (.L_HI(net55));
 sg13g2_tiehi _1603__56 (.L_HI(net56));
 sg13g2_tiehi _1510__57 (.L_HI(net57));
 sg13g2_tiehi _1589__58 (.L_HI(net58));
 sg13g2_tiehi _1509__59 (.L_HI(net59));
 sg13g2_tiehi _1588__60 (.L_HI(net60));
 sg13g2_tiehi _1508__61 (.L_HI(net61));
 sg13g2_tiehi _1587__62 (.L_HI(net62));
 sg13g2_tiehi _1507__63 (.L_HI(net63));
 sg13g2_tiehi _1586__64 (.L_HI(net64));
 sg13g2_tiehi _1506__65 (.L_HI(net65));
 sg13g2_tiehi _1585__66 (.L_HI(net66));
 sg13g2_tiehi _1505__67 (.L_HI(net67));
 sg13g2_tiehi _1584__68 (.L_HI(net68));
 sg13g2_tiehi _1504__69 (.L_HI(net69));
 sg13g2_tiehi _1583__70 (.L_HI(net70));
 sg13g2_tiehi _1503__71 (.L_HI(net71));
 sg13g2_tiehi _1582__72 (.L_HI(net72));
 sg13g2_tiehi _1502__73 (.L_HI(net73));
 sg13g2_tiehi _1581__74 (.L_HI(net74));
 sg13g2_tiehi _1501__75 (.L_HI(net75));
 sg13g2_tiehi _1601__76 (.L_HI(net76));
 sg13g2_tiehi _1500__77 (.L_HI(net77));
 sg13g2_tiehi _1580__78 (.L_HI(net78));
 sg13g2_tiehi _1499__79 (.L_HI(net79));
 sg13g2_tiehi _1441__80 (.L_HI(net80));
 sg13g2_tiehi _1498__81 (.L_HI(net81));
 sg13g2_tiehi _1579__82 (.L_HI(net82));
 sg13g2_tiehi _1497__83 (.L_HI(net83));
 sg13g2_tiehi _1600__84 (.L_HI(net84));
 sg13g2_tiehi _1496__85 (.L_HI(net85));
 sg13g2_tiehi _1578__86 (.L_HI(net86));
 sg13g2_tiehi _1495__87 (.L_HI(net87));
 sg13g2_tiehi _1602__88 (.L_HI(net88));
 sg13g2_tiehi _1494__89 (.L_HI(net89));
 sg13g2_tiehi _1577__90 (.L_HI(net90));
 sg13g2_tiehi _1493__91 (.L_HI(net91));
 sg13g2_tiehi _1599__92 (.L_HI(net92));
 sg13g2_tiehi _1492__93 (.L_HI(net93));
 sg13g2_tiehi _1576__94 (.L_HI(net94));
 sg13g2_tiehi _1491__95 (.L_HI(net95));
 sg13g2_tiehi _1598__96 (.L_HI(net96));
 sg13g2_tiehi _1490__97 (.L_HI(net97));
 sg13g2_tiehi _1575__98 (.L_HI(net98));
 sg13g2_tiehi _1489__99 (.L_HI(net99));
 sg13g2_tiehi _1597__100 (.L_HI(net100));
 sg13g2_tiehi _1488__101 (.L_HI(net101));
 sg13g2_tiehi _1574__102 (.L_HI(net102));
 sg13g2_tiehi _1487__103 (.L_HI(net103));
 sg13g2_tiehi _1596__104 (.L_HI(net104));
 sg13g2_tiehi _1486__105 (.L_HI(net105));
 sg13g2_tiehi _1573__106 (.L_HI(net106));
 sg13g2_tiehi _1485__107 (.L_HI(net107));
 sg13g2_tiehi _1595__108 (.L_HI(net108));
 sg13g2_tiehi _1484__109 (.L_HI(net109));
 sg13g2_tiehi _1572__110 (.L_HI(net110));
 sg13g2_tiehi _1483__111 (.L_HI(net111));
 sg13g2_tiehi _1482__112 (.L_HI(net112));
 sg13g2_tiehi _1481__113 (.L_HI(net113));
 sg13g2_tiehi _1480__114 (.L_HI(net114));
 sg13g2_tiehi _1479__115 (.L_HI(net115));
 sg13g2_tiehi _1478__116 (.L_HI(net116));
 sg13g2_tiehi _1477__117 (.L_HI(net117));
 sg13g2_tiehi _1476__118 (.L_HI(net118));
 sg13g2_tiehi _1475__119 (.L_HI(net179));
 sg13g2_tiehi _1474__120 (.L_HI(net180));
 sg13g2_tiehi _1473__121 (.L_HI(net181));
 sg13g2_tiehi _1472__122 (.L_HI(net182));
 sg13g2_tiehi _1471__123 (.L_HI(net183));
 sg13g2_tiehi _1470__124 (.L_HI(net184));
 sg13g2_tiehi _1469__125 (.L_HI(net185));
 sg13g2_tiehi _1468__126 (.L_HI(net186));
 sg13g2_tiehi _1467__127 (.L_HI(net187));
 sg13g2_tiehi _1466__128 (.L_HI(net188));
 sg13g2_tiehi _1465__129 (.L_HI(net189));
 sg13g2_tiehi _1464__130 (.L_HI(net190));
 sg13g2_tiehi _1463__131 (.L_HI(net191));
 sg13g2_tiehi _1462__132 (.L_HI(net192));
 sg13g2_tiehi _1461__133 (.L_HI(net193));
 sg13g2_tiehi _1460__134 (.L_HI(net194));
 sg13g2_tiehi _1459__135 (.L_HI(net195));
 sg13g2_tiehi _1458__136 (.L_HI(net196));
 sg13g2_tiehi _1457__137 (.L_HI(net197));
 sg13g2_tiehi _1456__138 (.L_HI(net198));
 sg13g2_tiehi _1455__139 (.L_HI(net199));
 sg13g2_tiehi _1454__140 (.L_HI(net200));
 sg13g2_tiehi _1453__141 (.L_HI(net201));
 sg13g2_tiehi _1452__142 (.L_HI(net202));
 sg13g2_tiehi _1451__143 (.L_HI(net203));
 sg13g2_tiehi _1450__144 (.L_HI(net204));
 sg13g2_tiehi _1449__145 (.L_HI(net205));
 sg13g2_tiehi _1448__146 (.L_HI(net206));
 sg13g2_tiehi _1447__147 (.L_HI(net207));
 sg13g2_tiehi _1446__148 (.L_HI(net208));
 sg13g2_tiehi _1445__149 (.L_HI(net209));
 sg13g2_tiehi _1444__150 (.L_HI(net210));
 sg13g2_tiehi _1443__151 (.L_HI(net211));
 sg13g2_tiehi _1442__152 (.L_HI(net212));
 sg13g2_tiehi _1437__153 (.L_HI(net213));
 sg13g2_tiehi _1436__154 (.L_HI(net214));
 sg13g2_tiehi _1435__155 (.L_HI(net215));
 sg13g2_tiehi _1434__156 (.L_HI(net216));
 sg13g2_tiehi _1433__157 (.L_HI(net217));
 sg13g2_tiehi _1432__158 (.L_HI(net218));
 sg13g2_tiehi _1431__159 (.L_HI(net219));
 sg13g2_tiehi _1430__160 (.L_HI(net220));
 sg13g2_tiehi _1429__161 (.L_HI(net221));
 sg13g2_tiehi _1428__162 (.L_HI(net222));
 sg13g2_tiehi _1427__163 (.L_HI(net223));
 sg13g2_tiehi _1426__164 (.L_HI(net224));
 sg13g2_tiehi _1425__165 (.L_HI(net225));
 sg13g2_tiehi _1424__166 (.L_HI(net226));
 sg13g2_tiehi _1423__167 (.L_HI(net227));
 sg13g2_tiehi _1422__168 (.L_HI(net228));
 sg13g2_tiehi _1421__169 (.L_HI(net229));
 sg13g2_tiehi _1420__170 (.L_HI(net230));
 sg13g2_tiehi _1419__171 (.L_HI(net231));
 sg13g2_tiehi _1418__172 (.L_HI(net232));
 sg13g2_tiehi _1594__173 (.L_HI(net233));
 sg13g2_tiehi _1571__174 (.L_HI(net234));
 sg13g2_tiehi _1570__175 (.L_HI(net235));
 sg13g2_tiehi _1569__176 (.L_HI(net236));
 sg13g2_tiehi _1568__177 (.L_HI(net237));
 sg13g2_tiehi _1567__178 (.L_HI(net238));
 sg13g2_tiehi _1566__179 (.L_HI(net239));
 sg13g2_tiehi _1565__180 (.L_HI(net240));
 sg13g2_tiehi _1564__181 (.L_HI(net241));
 sg13g2_tiehi _1563__182 (.L_HI(net242));
 sg13g2_tiehi _1562__183 (.L_HI(net243));
 sg13g2_tiehi _1561__184 (.L_HI(net244));
 sg13g2_tiehi _1560__185 (.L_HI(net245));
 sg13g2_tiehi _1559__186 (.L_HI(net246));
 sg13g2_tiehi _1558__187 (.L_HI(net247));
 sg13g2_tiehi _1557__188 (.L_HI(net248));
 sg13g2_tiehi _1556__189 (.L_HI(net249));
 sg13g2_tiehi _1555__190 (.L_HI(net250));
 sg13g2_tiehi _1554__191 (.L_HI(net251));
 sg13g2_tiehi _1553__192 (.L_HI(net252));
 sg13g2_tiehi _1552__193 (.L_HI(net253));
 sg13g2_tiehi _1551__194 (.L_HI(net254));
 sg13g2_tiehi _1550__195 (.L_HI(net255));
 sg13g2_tiehi _1549__196 (.L_HI(net256));
 sg13g2_tiehi _1548__197 (.L_HI(net257));
 sg13g2_tiehi _1547__198 (.L_HI(net258));
 sg13g2_tiehi _1546__199 (.L_HI(net259));
 sg13g2_tiehi _1545__200 (.L_HI(net260));
 sg13g2_tiehi _1544__201 (.L_HI(net261));
 sg13g2_tiehi _1543__202 (.L_HI(net262));
 sg13g2_tiehi _1542__203 (.L_HI(net263));
 sg13g2_tiehi _1541__204 (.L_HI(net264));
 sg13g2_tiehi _1540__205 (.L_HI(net265));
 sg13g2_tiehi _1539__206 (.L_HI(net266));
 sg13g2_tiehi _1538__207 (.L_HI(net267));
 sg13g2_tiehi _1537__208 (.L_HI(net268));
 sg13g2_tiehi _1536__209 (.L_HI(net269));
 sg13g2_tiehi _1535__210 (.L_HI(net270));
 sg13g2_tiehi _1534__211 (.L_HI(net271));
 sg13g2_tiehi _1533__212 (.L_HI(net272));
 sg13g2_tiehi _1532__213 (.L_HI(net273));
 sg13g2_tiehi _1531__214 (.L_HI(net274));
 sg13g2_tiehi tt_um_dranoel06_SAP1_215 (.L_HI(net275));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_dranoel06_SAP1_15 (.L_LO(net15));
 sg13g2_tielo tt_um_dranoel06_SAP1_16 (.L_LO(net16));
 sg13g2_tielo tt_um_dranoel06_SAP1_17 (.L_LO(net17));
 sg13g2_tielo tt_um_dranoel06_SAP1_18 (.L_LO(net18));
 sg13g2_tielo tt_um_dranoel06_SAP1_19 (.L_LO(net19));
 sg13g2_tielo tt_um_dranoel06_SAP1_20 (.L_LO(net20));
 sg13g2_tielo tt_um_dranoel06_SAP1_21 (.L_LO(net21));
 sg13g2_tielo tt_um_dranoel06_SAP1_22 (.L_LO(net22));
 sg13g2_tielo tt_um_dranoel06_SAP1_23 (.L_LO(net23));
 sg13g2_tielo tt_um_dranoel06_SAP1_24 (.L_LO(net24));
 sg13g2_tielo tt_um_dranoel06_SAP1_25 (.L_LO(net25));
 sg13g2_tielo tt_um_dranoel06_SAP1_26 (.L_LO(net26));
 sg13g2_tielo tt_um_dranoel06_SAP1_27 (.L_LO(net27));
 sg13g2_tiehi _1530__28 (.L_HI(net28));
 sg13g2_buf_1 _1806_ (.A(\uart0.tx ),
    .X(uio_out[6]));
 sg13g2_buf_8 fanout119 (.A(_0503_),
    .X(net119));
 sg13g2_buf_8 fanout120 (.A(_0503_),
    .X(net120));
 sg13g2_buf_8 fanout121 (.A(_0474_),
    .X(net121));
 sg13g2_buf_8 fanout122 (.A(_0474_),
    .X(net122));
 sg13g2_buf_8 fanout123 (.A(_0444_),
    .X(net123));
 sg13g2_buf_8 fanout124 (.A(_0444_),
    .X(net124));
 sg13g2_buf_8 fanout125 (.A(_0398_),
    .X(net125));
 sg13g2_buf_8 fanout126 (.A(_0398_),
    .X(net126));
 sg13g2_buf_8 fanout127 (.A(_0417_),
    .X(net127));
 sg13g2_buf_8 fanout128 (.A(_0417_),
    .X(net128));
 sg13g2_buf_8 fanout129 (.A(_0365_),
    .X(net129));
 sg13g2_buf_8 fanout130 (.A(_0365_),
    .X(net130));
 sg13g2_buf_8 fanout131 (.A(_0334_),
    .X(net131));
 sg13g2_buf_8 fanout132 (.A(_0334_),
    .X(net132));
 sg13g2_buf_8 fanout133 (.A(_0295_),
    .X(net133));
 sg13g2_buf_8 fanout134 (.A(_0295_),
    .X(net134));
 sg13g2_buf_8 fanout135 (.A(_0602_),
    .X(net135));
 sg13g2_buf_8 fanout136 (.A(_0579_),
    .X(net136));
 sg13g2_buf_8 fanout137 (.A(_0575_),
    .X(net137));
 sg13g2_buf_8 fanout138 (.A(_0525_),
    .X(net138));
 sg13g2_buf_8 fanout139 (.A(net140),
    .X(net139));
 sg13g2_buf_8 fanout140 (.A(_0506_),
    .X(net140));
 sg13g2_buf_8 fanout141 (.A(_0264_),
    .X(net141));
 sg13g2_buf_8 fanout142 (.A(net143),
    .X(net142));
 sg13g2_buf_8 fanout143 (.A(net144),
    .X(net143));
 sg13g2_buf_8 fanout144 (.A(_0229_),
    .X(net144));
 sg13g2_buf_8 fanout145 (.A(_0220_),
    .X(net145));
 sg13g2_buf_8 fanout146 (.A(_0204_),
    .X(net146));
 sg13g2_buf_8 fanout147 (.A(_0203_),
    .X(net147));
 sg13g2_buf_8 fanout148 (.A(net486),
    .X(net148));
 sg13g2_buf_8 fanout149 (.A(net150),
    .X(net149));
 sg13g2_buf_8 fanout150 (.A(_0003_),
    .X(net150));
 sg13g2_buf_8 fanout151 (.A(net153),
    .X(net151));
 sg13g2_buf_8 fanout152 (.A(net153),
    .X(net152));
 sg13g2_buf_8 fanout153 (.A(_0002_),
    .X(net153));
 sg13g2_buf_8 fanout154 (.A(net156),
    .X(net154));
 sg13g2_buf_8 fanout155 (.A(net156),
    .X(net155));
 sg13g2_buf_8 fanout156 (.A(_0001_),
    .X(net156));
 sg13g2_buf_8 fanout157 (.A(net159),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(net159),
    .X(net158));
 sg13g2_buf_8 fanout159 (.A(_0001_),
    .X(net159));
 sg13g2_buf_8 fanout160 (.A(net162),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(net162),
    .X(net161));
 sg13g2_buf_8 fanout162 (.A(net164),
    .X(net162));
 sg13g2_buf_8 fanout163 (.A(net164),
    .X(net163));
 sg13g2_buf_8 fanout164 (.A(_0000_),
    .X(net164));
 sg13g2_buf_8 fanout165 (.A(net169),
    .X(net165));
 sg13g2_buf_1 fanout166 (.A(net169),
    .X(net166));
 sg13g2_buf_8 fanout167 (.A(net169),
    .X(net167));
 sg13g2_buf_8 fanout168 (.A(net169),
    .X(net168));
 sg13g2_buf_8 fanout169 (.A(_0000_),
    .X(net169));
 sg13g2_buf_8 fanout170 (.A(net171),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_0000_),
    .X(net171));
 sg13g2_buf_8 fanout172 (.A(net173),
    .X(net172));
 sg13g2_buf_8 fanout173 (.A(net174),
    .X(net173));
 sg13g2_buf_8 fanout174 (.A(_0199_),
    .X(net174));
 sg13g2_buf_8 fanout175 (.A(net177),
    .X(net175));
 sg13g2_buf_1 fanout176 (.A(net177),
    .X(net176));
 sg13g2_buf_8 fanout177 (.A(net178),
    .X(net177));
 sg13g2_buf_8 fanout178 (.A(rst_n),
    .X(net178));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[7]),
    .X(net13));
 sg13g2_tielo tt_um_dranoel06_SAP1_14 (.L_LO(net14));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_8 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_8 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_8 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_8 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_8 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_8 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_8 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_8 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_8 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_8 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_8 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_8 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_8 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_8 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_8 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_8 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_8 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_8 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_8 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_8 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_8 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_8 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_8 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_8 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_8 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_8 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_8 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_8 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_8 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_8 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_8 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_5_12__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_5_18__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_23__leaf_clk));
 sg13g2_buf_1 clkload6 (.A(clknet_5_24__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkload8 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\uart0.tx_en_prev ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0004_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold3 (.A(\uart0.bit_counter[3] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0189_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold5 (.A(\cpu0.ir[2] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0080_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold7 (.A(\cpu0.ir[3] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0081_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold9 (.A(\cpu0.ir[0] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0078_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold11 (.A(\cpu0.ir[1] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0079_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold13 (.A(\cpu0.ram[13][1] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold14 (.A(\cpu0.ram[7][1] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold15 (.A(\cpu0.ram[14][3] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold16 (.A(\cpu0.ram[12][2] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold17 (.A(\uart0.uart_state[2] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0223_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold19 (.A(\cpu0.b_reg[6] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0164_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold21 (.A(uo_out[3]),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0097_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold23 (.A(\cpu0.b_reg[1] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0159_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold25 (.A(uo_out[2]),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0096_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold27 (.A(\cpu0.b_reg[3] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0161_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold29 (.A(\uart0.uart_state[3] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0006_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold31 (.A(uo_out[5]),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold32 (.A(\cpu0.b_reg[5] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0163_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold34 (.A(\cpu0.b_reg[2] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0160_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold36 (.A(\cpu0.b_reg[0] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0158_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold38 (.A(\cpu0.ram[8][1] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold39 (.A(\cpu0.ram[1][1] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold40 (.A(\cpu0.ram[15][0] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold41 (.A(\cpu0.ram[14][1] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold42 (.A(\cpu0.ram[4][2] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold43 (.A(\cpu0.ram[0][4] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold44 (.A(\cpu0.ram[12][5] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold45 (.A(\cpu0.ram[10][1] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold46 (.A(\cpu0.ram[15][6] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold47 (.A(\cpu0.ram[4][7] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold48 (.A(uo_out[1]),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold49 (.A(\cpu0.ram[10][5] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold50 (.A(\cpu0.ram[9][7] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold51 (.A(\cpu0.ram[3][5] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold52 (.A(\cpu0.ram[14][2] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold53 (.A(\cpu0.ram[14][0] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold54 (.A(\cpu0.ram[2][1] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold55 (.A(\cpu0.ram[15][4] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold56 (.A(\cpu0.ram[8][3] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold57 (.A(\cpu0.ram[13][6] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold58 (.A(\cpu0.ram[11][0] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold59 (.A(uo_out[0]),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0094_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold61 (.A(\cpu0.ram[5][5] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold62 (.A(\cpu0.a_reg[4] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold63 (.A(\cpu0.ram[7][5] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold64 (.A(uo_out[6]),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold65 (.A(\cpu0.ram[13][2] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold66 (.A(\cpu0.ram[6][3] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold67 (.A(\cpu0.ram[3][4] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold68 (.A(\cpu0.ram[4][0] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold69 (.A(\cpu0.ram[6][4] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold70 (.A(\cpu0.ram[5][0] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold71 (.A(\cpu0.ram[13][7] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold72 (.A(\cpu0.ram[1][5] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold73 (.A(\cpu0.ram[10][2] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold74 (.A(\cpu0.ram[8][7] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold75 (.A(\cpu0.ram[0][0] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold76 (.A(\cpu0.ram[14][6] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold77 (.A(\cpu0.ram[0][2] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold78 (.A(\cpu0.ram[1][0] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold79 (.A(\cpu0.ram[7][7] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold80 (.A(\cpu0.ram[4][4] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold81 (.A(\cpu0.ram[14][4] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold82 (.A(\cpu0.ram[13][4] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold83 (.A(\cpu0.ram[1][6] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold84 (.A(\cpu0.ram[3][0] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold85 (.A(\cpu0.ram[5][3] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold86 (.A(\cpu0.ram[0][5] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold87 (.A(\cpu0.ram[1][2] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold88 (.A(\cpu0.ram[2][5] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold89 (.A(\cpu0.ram[10][7] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold90 (.A(\cpu0.ram[4][3] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold91 (.A(\cpu0.ram[11][4] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold92 (.A(\cpu0.ram[0][6] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold93 (.A(\cpu0.ram[11][1] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold94 (.A(\cpu0.ram[12][7] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold95 (.A(\cpu0.ram[14][5] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold96 (.A(\cpu0.ram[3][3] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold97 (.A(\cpu0.ram[4][1] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold98 (.A(\cpu0.ram[9][0] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold99 (.A(\cpu0.ram[3][7] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold100 (.A(\cpu0.ram[11][7] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold101 (.A(\cpu0.ram[5][2] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold102 (.A(\cpu0.ram[7][6] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold103 (.A(\cpu0.ram[10][6] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold104 (.A(\cpu0.ram[8][5] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold105 (.A(\cpu0.ram[12][3] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold106 (.A(\cpu0.ram[6][0] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold107 (.A(\cpu0.ram[9][3] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold108 (.A(\cpu0.ram[11][3] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold109 (.A(\cpu0.ram[12][1] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold110 (.A(\cpu0.ram[0][7] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold111 (.A(\cpu0.ram[13][3] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold112 (.A(\cpu0.ram[10][4] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold113 (.A(\cpu0.ram[2][6] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold114 (.A(\cpu0.ram[11][5] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold115 (.A(\cpu0.ram[2][4] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold116 (.A(\cpu0.ram[3][2] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold117 (.A(\cpu0.ram[2][2] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold118 (.A(\cpu0.ram[6][6] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold119 (.A(\cpu0.ram[5][7] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold120 (.A(\cpu0.ram[1][4] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold121 (.A(\cpu0.ram[6][2] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold122 (.A(\cpu0.ram[5][4] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold123 (.A(\cpu0.ram[9][1] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold124 (.A(\cpu0.ram[11][2] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold125 (.A(\cpu0.ram[15][5] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold126 (.A(\cpu0.ram[12][6] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold127 (.A(\cpu0.ram[2][7] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold128 (.A(\cpu0.ram[3][6] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold129 (.A(\cpu0.ram[4][5] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold130 (.A(\cpu0.ram[0][1] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold131 (.A(\cpu0.ram[6][5] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold132 (.A(\cpu0.ram[15][1] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold133 (.A(\cpu0.ram[12][4] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold134 (.A(\cpu0.ram[0][3] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold135 (.A(\cpu0.ram[6][7] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold136 (.A(\cpu0.ram[10][0] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold137 (.A(\cpu0.ram[8][4] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold138 (.A(\cpu0.ram[5][6] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold139 (.A(\cpu0.ram[7][0] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold140 (.A(\cpu0.ram[15][2] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold141 (.A(\cpu0.ram[2][0] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold142 (.A(\cpu0.ram[13][0] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold143 (.A(\cpu0.ram[13][5] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold144 (.A(\cpu0.ram[9][5] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold145 (.A(\cpu0.ram[8][6] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold146 (.A(\cpu0.ram[4][6] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold147 (.A(\cpu0.ram[8][0] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold148 (.A(\cpu0.ram[6][1] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold149 (.A(\cpu0.ram[7][4] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold150 (.A(\cpu0.ram[12][0] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold151 (.A(\cpu0.ram[10][3] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold152 (.A(\cpu0.ram[11][6] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold153 (.A(\cpu0.ram[1][7] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold154 (.A(\cpu0.ram[15][7] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold155 (.A(\cpu0.ram[5][1] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold156 (.A(\cpu0.ram[9][2] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold157 (.A(\cpu0.ram[7][3] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold158 (.A(\cpu0.ram[14][7] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold159 (.A(\uart0.bit_counter[2] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0222_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0005_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold162 (.A(\cpu0.a_reg[6] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold163 (.A(\cpu0.ram[9][4] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold164 (.A(\cpu0.ram[15][3] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold165 (.A(\cpu0.ram[2][3] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold166 (.A(\cpu0.ram[8][2] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold167 (.A(\cpu0.ram[3][1] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold168 (.A(\cpu0.ram[9][6] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold169 (.A(\cpu0.ram[1][3] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold170 (.A(\cpu0.ram[7][2] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold171 (.A(uo_out[7]),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold172 (.A(\cpu0.b_reg[4] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold173 (.A(\cpu0.ir[4] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold174 (.A(uo_out[4]),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold175 (.A(\cpu0.ir[6] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0084_),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold177 (.A(\cpu0.b_reg[7] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold178 (.A(\cpu0.ir[5] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0083_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold180 (.A(\uart0.uart_state[0] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0176_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold182 (.A(\cpu0.a_reg[5] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold183 (.A(\cpu0.carry_flag ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0167_),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold185 (.A(\uart0.bit_counter[1] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0615_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold187 (.A(\cpu0.a_reg[7] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold188 (.A(\cpu0.step[2] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0516_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0029_),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold191 (.A(\cpu0.a_reg[2] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold192 (.A(\cpu0.mar[3] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold193 (.A(\cpu0.step[1] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0239_),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0190_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold196 (.A(\cpu0.a_reg[1] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold197 (.A(\cpu0.pc[3] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold198 (.A(\cpu0.a_reg[0] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0070_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold200 (.A(\cpu0.mar[2] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold201 (.A(\cpu0.a_reg[3] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold202 (.A(\cpu0.pc[0] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold203 (.A(\cpu0.pc[2] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold204 (.A(\cpu0.mar[1] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold205 (.A(\cpu0.pc[1] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold206 (.A(\cpu0.zero_flag ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold207 (.A(\cpu0.mar[0] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold208 (.A(\uart0.bit_counter[0] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0613_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold210 (.A(\cpu0.step[0] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold211 (.A(\cpu0.ir[7] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold212 (.A(\uart0.uart_state[1] ),
    .X(net487));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_fill_2 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_194 ();
 sg13g2_decap_8 FILLER_0_201 ();
 sg13g2_fill_2 FILLER_0_208 ();
 sg13g2_fill_1 FILLER_0_210 ();
 sg13g2_fill_1 FILLER_0_215 ();
 sg13g2_decap_4 FILLER_0_234 ();
 sg13g2_fill_2 FILLER_0_238 ();
 sg13g2_fill_1 FILLER_0_244 ();
 sg13g2_fill_2 FILLER_0_255 ();
 sg13g2_decap_4 FILLER_0_267 ();
 sg13g2_fill_2 FILLER_0_275 ();
 sg13g2_decap_8 FILLER_0_286 ();
 sg13g2_decap_8 FILLER_0_293 ();
 sg13g2_decap_4 FILLER_0_300 ();
 sg13g2_decap_4 FILLER_0_314 ();
 sg13g2_fill_2 FILLER_0_318 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_4 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_141 ();
 sg13g2_decap_8 FILLER_1_148 ();
 sg13g2_decap_8 FILLER_1_155 ();
 sg13g2_decap_4 FILLER_1_162 ();
 sg13g2_fill_2 FILLER_1_166 ();
 sg13g2_fill_1 FILLER_1_195 ();
 sg13g2_fill_2 FILLER_1_233 ();
 sg13g2_decap_4 FILLER_1_262 ();
 sg13g2_decap_8 FILLER_1_293 ();
 sg13g2_decap_4 FILLER_1_300 ();
 sg13g2_fill_1 FILLER_1_304 ();
 sg13g2_decap_8 FILLER_1_332 ();
 sg13g2_fill_2 FILLER_1_339 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_fill_2 FILLER_2_49 ();
 sg13g2_fill_1 FILLER_2_51 ();
 sg13g2_decap_4 FILLER_2_62 ();
 sg13g2_decap_8 FILLER_2_75 ();
 sg13g2_decap_8 FILLER_2_82 ();
 sg13g2_decap_8 FILLER_2_89 ();
 sg13g2_decap_8 FILLER_2_96 ();
 sg13g2_decap_8 FILLER_2_103 ();
 sg13g2_fill_1 FILLER_2_110 ();
 sg13g2_decap_8 FILLER_2_115 ();
 sg13g2_decap_8 FILLER_2_122 ();
 sg13g2_fill_2 FILLER_2_129 ();
 sg13g2_fill_1 FILLER_2_131 ();
 sg13g2_decap_4 FILLER_2_168 ();
 sg13g2_fill_1 FILLER_2_172 ();
 sg13g2_decap_8 FILLER_2_177 ();
 sg13g2_decap_8 FILLER_2_184 ();
 sg13g2_fill_1 FILLER_2_191 ();
 sg13g2_decap_8 FILLER_2_242 ();
 sg13g2_decap_8 FILLER_2_295 ();
 sg13g2_decap_8 FILLER_2_302 ();
 sg13g2_fill_1 FILLER_2_309 ();
 sg13g2_decap_8 FILLER_2_314 ();
 sg13g2_decap_8 FILLER_2_358 ();
 sg13g2_decap_8 FILLER_2_365 ();
 sg13g2_decap_8 FILLER_2_372 ();
 sg13g2_decap_8 FILLER_2_379 ();
 sg13g2_decap_8 FILLER_2_386 ();
 sg13g2_decap_8 FILLER_2_393 ();
 sg13g2_decap_8 FILLER_2_400 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_fill_2 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_40 ();
 sg13g2_fill_2 FILLER_3_47 ();
 sg13g2_decap_8 FILLER_3_76 ();
 sg13g2_fill_1 FILLER_3_143 ();
 sg13g2_fill_1 FILLER_3_167 ();
 sg13g2_fill_2 FILLER_3_216 ();
 sg13g2_fill_1 FILLER_3_218 ();
 sg13g2_fill_2 FILLER_3_228 ();
 sg13g2_fill_2 FILLER_3_253 ();
 sg13g2_fill_2 FILLER_3_276 ();
 sg13g2_decap_8 FILLER_3_324 ();
 sg13g2_fill_1 FILLER_3_331 ();
 sg13g2_decap_4 FILLER_3_346 ();
 sg13g2_fill_2 FILLER_3_354 ();
 sg13g2_decap_8 FILLER_3_365 ();
 sg13g2_decap_8 FILLER_3_372 ();
 sg13g2_decap_8 FILLER_3_379 ();
 sg13g2_decap_8 FILLER_3_386 ();
 sg13g2_decap_8 FILLER_3_393 ();
 sg13g2_decap_8 FILLER_3_400 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_fill_1 FILLER_4_21 ();
 sg13g2_fill_2 FILLER_4_66 ();
 sg13g2_fill_1 FILLER_4_105 ();
 sg13g2_fill_1 FILLER_4_110 ();
 sg13g2_fill_2 FILLER_4_176 ();
 sg13g2_decap_8 FILLER_4_191 ();
 sg13g2_fill_1 FILLER_4_198 ();
 sg13g2_fill_2 FILLER_4_236 ();
 sg13g2_fill_1 FILLER_4_280 ();
 sg13g2_fill_1 FILLER_4_306 ();
 sg13g2_decap_8 FILLER_4_337 ();
 sg13g2_fill_1 FILLER_4_344 ();
 sg13g2_decap_4 FILLER_4_372 ();
 sg13g2_decap_8 FILLER_4_380 ();
 sg13g2_decap_8 FILLER_4_387 ();
 sg13g2_decap_8 FILLER_4_394 ();
 sg13g2_decap_8 FILLER_4_401 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_fill_2 FILLER_5_7 ();
 sg13g2_fill_1 FILLER_5_9 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_4 FILLER_5_21 ();
 sg13g2_fill_1 FILLER_5_44 ();
 sg13g2_decap_8 FILLER_5_93 ();
 sg13g2_fill_2 FILLER_5_144 ();
 sg13g2_fill_1 FILLER_5_146 ();
 sg13g2_decap_4 FILLER_5_205 ();
 sg13g2_fill_2 FILLER_5_209 ();
 sg13g2_fill_2 FILLER_5_234 ();
 sg13g2_fill_1 FILLER_5_236 ();
 sg13g2_fill_1 FILLER_5_246 ();
 sg13g2_fill_2 FILLER_5_270 ();
 sg13g2_fill_2 FILLER_5_309 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_4 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_401 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_4 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_4 ();
 sg13g2_fill_2 FILLER_6_32 ();
 sg13g2_fill_1 FILLER_6_34 ();
 sg13g2_fill_2 FILLER_6_49 ();
 sg13g2_decap_4 FILLER_6_81 ();
 sg13g2_fill_2 FILLER_6_89 ();
 sg13g2_fill_2 FILLER_6_138 ();
 sg13g2_fill_1 FILLER_6_145 ();
 sg13g2_decap_4 FILLER_6_191 ();
 sg13g2_fill_1 FILLER_6_222 ();
 sg13g2_fill_1 FILLER_6_250 ();
 sg13g2_fill_2 FILLER_6_278 ();
 sg13g2_fill_2 FILLER_6_290 ();
 sg13g2_fill_2 FILLER_6_301 ();
 sg13g2_fill_2 FILLER_6_340 ();
 sg13g2_fill_2 FILLER_6_395 ();
 sg13g2_fill_1 FILLER_6_397 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_4 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_31 ();
 sg13g2_fill_1 FILLER_7_33 ();
 sg13g2_fill_2 FILLER_7_78 ();
 sg13g2_decap_4 FILLER_7_107 ();
 sg13g2_fill_1 FILLER_7_138 ();
 sg13g2_fill_2 FILLER_7_149 ();
 sg13g2_fill_1 FILLER_7_151 ();
 sg13g2_decap_4 FILLER_7_183 ();
 sg13g2_fill_2 FILLER_7_187 ();
 sg13g2_fill_2 FILLER_7_203 ();
 sg13g2_fill_1 FILLER_7_205 ();
 sg13g2_decap_8 FILLER_7_215 ();
 sg13g2_fill_2 FILLER_7_227 ();
 sg13g2_fill_1 FILLER_7_229 ();
 sg13g2_decap_4 FILLER_7_235 ();
 sg13g2_fill_2 FILLER_7_263 ();
 sg13g2_fill_1 FILLER_7_274 ();
 sg13g2_fill_2 FILLER_7_312 ();
 sg13g2_fill_1 FILLER_7_314 ();
 sg13g2_fill_2 FILLER_7_332 ();
 sg13g2_fill_2 FILLER_7_344 ();
 sg13g2_fill_1 FILLER_7_346 ();
 sg13g2_fill_2 FILLER_7_369 ();
 sg13g2_fill_1 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_13 ();
 sg13g2_fill_1 FILLER_8_20 ();
 sg13g2_fill_1 FILLER_8_114 ();
 sg13g2_fill_2 FILLER_8_125 ();
 sg13g2_fill_1 FILLER_8_127 ();
 sg13g2_fill_1 FILLER_8_147 ();
 sg13g2_decap_4 FILLER_8_179 ();
 sg13g2_decap_8 FILLER_8_215 ();
 sg13g2_fill_2 FILLER_8_253 ();
 sg13g2_fill_2 FILLER_8_273 ();
 sg13g2_fill_2 FILLER_8_288 ();
 sg13g2_fill_2 FILLER_8_312 ();
 sg13g2_fill_2 FILLER_8_332 ();
 sg13g2_fill_1 FILLER_8_348 ();
 sg13g2_decap_4 FILLER_8_404 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_47 ();
 sg13g2_decap_4 FILLER_9_78 ();
 sg13g2_fill_1 FILLER_9_82 ();
 sg13g2_fill_1 FILLER_9_146 ();
 sg13g2_fill_2 FILLER_9_157 ();
 sg13g2_fill_1 FILLER_9_159 ();
 sg13g2_decap_8 FILLER_9_179 ();
 sg13g2_fill_1 FILLER_9_186 ();
 sg13g2_fill_2 FILLER_9_197 ();
 sg13g2_fill_1 FILLER_9_199 ();
 sg13g2_decap_4 FILLER_9_213 ();
 sg13g2_fill_1 FILLER_9_217 ();
 sg13g2_fill_1 FILLER_9_231 ();
 sg13g2_fill_2 FILLER_9_260 ();
 sg13g2_fill_2 FILLER_9_289 ();
 sg13g2_fill_1 FILLER_9_291 ();
 sg13g2_fill_1 FILLER_9_319 ();
 sg13g2_fill_1 FILLER_9_366 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_85 ();
 sg13g2_decap_4 FILLER_10_102 ();
 sg13g2_fill_2 FILLER_10_106 ();
 sg13g2_decap_8 FILLER_10_117 ();
 sg13g2_decap_4 FILLER_10_128 ();
 sg13g2_decap_4 FILLER_10_217 ();
 sg13g2_fill_2 FILLER_10_231 ();
 sg13g2_fill_1 FILLER_10_233 ();
 sg13g2_fill_2 FILLER_10_273 ();
 sg13g2_fill_2 FILLER_10_370 ();
 sg13g2_decap_4 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_4 ();
 sg13g2_fill_2 FILLER_11_107 ();
 sg13g2_fill_1 FILLER_11_109 ();
 sg13g2_fill_1 FILLER_11_120 ();
 sg13g2_fill_2 FILLER_11_125 ();
 sg13g2_fill_2 FILLER_11_174 ();
 sg13g2_decap_4 FILLER_11_180 ();
 sg13g2_fill_1 FILLER_11_184 ();
 sg13g2_fill_2 FILLER_11_220 ();
 sg13g2_fill_2 FILLER_11_248 ();
 sg13g2_fill_2 FILLER_11_300 ();
 sg13g2_fill_1 FILLER_11_302 ();
 sg13g2_fill_2 FILLER_11_336 ();
 sg13g2_fill_2 FILLER_11_378 ();
 sg13g2_fill_1 FILLER_11_380 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_4 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_4 ();
 sg13g2_fill_2 FILLER_12_69 ();
 sg13g2_fill_1 FILLER_12_71 ();
 sg13g2_fill_1 FILLER_12_143 ();
 sg13g2_fill_1 FILLER_12_152 ();
 sg13g2_fill_2 FILLER_12_168 ();
 sg13g2_fill_1 FILLER_12_170 ();
 sg13g2_fill_1 FILLER_12_222 ();
 sg13g2_fill_1 FILLER_12_232 ();
 sg13g2_decap_8 FILLER_12_243 ();
 sg13g2_fill_1 FILLER_12_250 ();
 sg13g2_fill_1 FILLER_12_270 ();
 sg13g2_decap_8 FILLER_12_302 ();
 sg13g2_decap_4 FILLER_12_309 ();
 sg13g2_fill_1 FILLER_12_313 ();
 sg13g2_fill_1 FILLER_12_327 ();
 sg13g2_fill_2 FILLER_12_338 ();
 sg13g2_fill_1 FILLER_12_340 ();
 sg13g2_fill_2 FILLER_12_355 ();
 sg13g2_fill_2 FILLER_12_367 ();
 sg13g2_fill_1 FILLER_12_369 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_7 ();
 sg13g2_fill_1 FILLER_13_9 ();
 sg13g2_decap_4 FILLER_13_18 ();
 sg13g2_fill_1 FILLER_13_22 ();
 sg13g2_fill_2 FILLER_13_33 ();
 sg13g2_fill_1 FILLER_13_35 ();
 sg13g2_decap_4 FILLER_13_74 ();
 sg13g2_fill_1 FILLER_13_78 ();
 sg13g2_decap_4 FILLER_13_106 ();
 sg13g2_fill_2 FILLER_13_110 ();
 sg13g2_fill_1 FILLER_13_116 ();
 sg13g2_fill_2 FILLER_13_126 ();
 sg13g2_decap_4 FILLER_13_177 ();
 sg13g2_decap_4 FILLER_13_206 ();
 sg13g2_fill_1 FILLER_13_210 ();
 sg13g2_fill_1 FILLER_13_265 ();
 sg13g2_decap_4 FILLER_13_329 ();
 sg13g2_fill_2 FILLER_13_360 ();
 sg13g2_fill_1 FILLER_13_381 ();
 sg13g2_decap_4 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_31 ();
 sg13g2_fill_2 FILLER_14_82 ();
 sg13g2_fill_1 FILLER_14_134 ();
 sg13g2_fill_2 FILLER_14_148 ();
 sg13g2_fill_1 FILLER_14_150 ();
 sg13g2_decap_4 FILLER_14_162 ();
 sg13g2_fill_1 FILLER_14_166 ();
 sg13g2_fill_1 FILLER_14_171 ();
 sg13g2_decap_4 FILLER_14_191 ();
 sg13g2_fill_2 FILLER_14_209 ();
 sg13g2_fill_1 FILLER_14_241 ();
 sg13g2_fill_2 FILLER_14_246 ();
 sg13g2_fill_1 FILLER_14_248 ();
 sg13g2_fill_1 FILLER_14_288 ();
 sg13g2_fill_2 FILLER_14_311 ();
 sg13g2_fill_1 FILLER_14_313 ();
 sg13g2_fill_2 FILLER_14_332 ();
 sg13g2_fill_1 FILLER_14_334 ();
 sg13g2_decap_4 FILLER_14_348 ();
 sg13g2_fill_2 FILLER_14_352 ();
 sg13g2_fill_2 FILLER_14_369 ();
 sg13g2_fill_1 FILLER_14_381 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_13 ();
 sg13g2_fill_1 FILLER_15_20 ();
 sg13g2_fill_2 FILLER_15_108 ();
 sg13g2_fill_2 FILLER_15_142 ();
 sg13g2_fill_1 FILLER_15_157 ();
 sg13g2_fill_2 FILLER_15_225 ();
 sg13g2_decap_4 FILLER_15_268 ();
 sg13g2_fill_1 FILLER_15_272 ();
 sg13g2_fill_2 FILLER_15_286 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_fill_2 FILLER_15_322 ();
 sg13g2_fill_1 FILLER_15_324 ();
 sg13g2_fill_2 FILLER_15_343 ();
 sg13g2_fill_2 FILLER_15_363 ();
 sg13g2_fill_2 FILLER_15_375 ();
 sg13g2_fill_1 FILLER_15_377 ();
 sg13g2_decap_4 FILLER_16_31 ();
 sg13g2_fill_2 FILLER_16_80 ();
 sg13g2_fill_2 FILLER_16_92 ();
 sg13g2_fill_1 FILLER_16_94 ();
 sg13g2_fill_2 FILLER_16_108 ();
 sg13g2_fill_2 FILLER_16_160 ();
 sg13g2_fill_1 FILLER_16_162 ();
 sg13g2_decap_8 FILLER_16_167 ();
 sg13g2_fill_1 FILLER_16_174 ();
 sg13g2_decap_4 FILLER_16_188 ();
 sg13g2_fill_1 FILLER_16_219 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_fill_2 FILLER_16_299 ();
 sg13g2_fill_2 FILLER_16_338 ();
 sg13g2_fill_1 FILLER_16_340 ();
 sg13g2_fill_2 FILLER_16_368 ();
 sg13g2_fill_1 FILLER_16_370 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_2 ();
 sg13g2_fill_1 FILLER_17_35 ();
 sg13g2_fill_2 FILLER_17_50 ();
 sg13g2_fill_1 FILLER_17_52 ();
 sg13g2_decap_4 FILLER_17_62 ();
 sg13g2_fill_2 FILLER_17_87 ();
 sg13g2_fill_1 FILLER_17_89 ();
 sg13g2_decap_8 FILLER_17_117 ();
 sg13g2_fill_2 FILLER_17_152 ();
 sg13g2_fill_1 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_177 ();
 sg13g2_decap_8 FILLER_17_184 ();
 sg13g2_fill_1 FILLER_17_191 ();
 sg13g2_decap_8 FILLER_17_213 ();
 sg13g2_decap_4 FILLER_17_220 ();
 sg13g2_fill_2 FILLER_17_256 ();
 sg13g2_fill_1 FILLER_17_286 ();
 sg13g2_fill_2 FILLER_17_369 ();
 sg13g2_fill_2 FILLER_17_389 ();
 sg13g2_fill_1 FILLER_17_391 ();
 sg13g2_decap_4 FILLER_17_405 ();
 sg13g2_decap_4 FILLER_18_48 ();
 sg13g2_fill_2 FILLER_18_52 ();
 sg13g2_fill_1 FILLER_18_68 ();
 sg13g2_decap_8 FILLER_18_114 ();
 sg13g2_fill_1 FILLER_18_121 ();
 sg13g2_fill_2 FILLER_18_165 ();
 sg13g2_decap_4 FILLER_18_194 ();
 sg13g2_fill_1 FILLER_18_198 ();
 sg13g2_decap_4 FILLER_18_209 ();
 sg13g2_fill_2 FILLER_18_213 ();
 sg13g2_fill_2 FILLER_18_266 ();
 sg13g2_fill_1 FILLER_18_268 ();
 sg13g2_fill_2 FILLER_18_273 ();
 sg13g2_fill_1 FILLER_18_288 ();
 sg13g2_decap_4 FILLER_18_336 ();
 sg13g2_fill_2 FILLER_18_380 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_4 ();
 sg13g2_fill_1 FILLER_19_9 ();
 sg13g2_fill_1 FILLER_19_29 ();
 sg13g2_decap_4 FILLER_19_84 ();
 sg13g2_fill_2 FILLER_19_88 ();
 sg13g2_decap_4 FILLER_19_131 ();
 sg13g2_fill_2 FILLER_19_144 ();
 sg13g2_fill_1 FILLER_19_146 ();
 sg13g2_fill_1 FILLER_19_160 ();
 sg13g2_decap_8 FILLER_19_165 ();
 sg13g2_fill_1 FILLER_19_172 ();
 sg13g2_fill_2 FILLER_19_183 ();
 sg13g2_fill_2 FILLER_19_195 ();
 sg13g2_fill_2 FILLER_19_237 ();
 sg13g2_fill_1 FILLER_19_248 ();
 sg13g2_fill_1 FILLER_19_263 ();
 sg13g2_fill_2 FILLER_19_291 ();
 sg13g2_fill_2 FILLER_19_307 ();
 sg13g2_decap_4 FILLER_19_339 ();
 sg13g2_fill_2 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_fill_1 FILLER_19_385 ();
 sg13g2_fill_1 FILLER_19_390 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_4 FILLER_20_27 ();
 sg13g2_fill_2 FILLER_20_31 ();
 sg13g2_decap_4 FILLER_20_56 ();
 sg13g2_fill_1 FILLER_20_60 ();
 sg13g2_decap_8 FILLER_20_65 ();
 sg13g2_fill_1 FILLER_20_72 ();
 sg13g2_fill_2 FILLER_20_93 ();
 sg13g2_fill_1 FILLER_20_99 ();
 sg13g2_decap_8 FILLER_20_144 ();
 sg13g2_fill_1 FILLER_20_204 ();
 sg13g2_fill_1 FILLER_20_218 ();
 sg13g2_decap_4 FILLER_20_256 ();
 sg13g2_fill_2 FILLER_20_260 ();
 sg13g2_fill_2 FILLER_20_275 ();
 sg13g2_fill_1 FILLER_20_277 ();
 sg13g2_decap_8 FILLER_20_338 ();
 sg13g2_fill_2 FILLER_20_345 ();
 sg13g2_fill_1 FILLER_20_347 ();
 sg13g2_fill_2 FILLER_20_368 ();
 sg13g2_fill_1 FILLER_20_380 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_fill_1 FILLER_21_14 ();
 sg13g2_decap_4 FILLER_21_52 ();
 sg13g2_decap_4 FILLER_21_83 ();
 sg13g2_fill_1 FILLER_21_150 ();
 sg13g2_fill_2 FILLER_21_177 ();
 sg13g2_fill_2 FILLER_21_212 ();
 sg13g2_fill_2 FILLER_21_224 ();
 sg13g2_fill_1 FILLER_21_226 ();
 sg13g2_decap_4 FILLER_21_253 ();
 sg13g2_decap_4 FILLER_21_270 ();
 sg13g2_fill_2 FILLER_21_274 ();
 sg13g2_fill_2 FILLER_21_302 ();
 sg13g2_fill_1 FILLER_21_304 ();
 sg13g2_fill_1 FILLER_21_309 ();
 sg13g2_fill_2 FILLER_21_314 ();
 sg13g2_fill_2 FILLER_21_326 ();
 sg13g2_fill_1 FILLER_21_328 ();
 sg13g2_fill_1 FILLER_21_371 ();
 sg13g2_fill_2 FILLER_22_27 ();
 sg13g2_decap_8 FILLER_22_52 ();
 sg13g2_fill_2 FILLER_22_59 ();
 sg13g2_decap_4 FILLER_22_70 ();
 sg13g2_fill_1 FILLER_22_74 ();
 sg13g2_decap_8 FILLER_22_107 ();
 sg13g2_decap_8 FILLER_22_114 ();
 sg13g2_fill_2 FILLER_22_121 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_fill_1 FILLER_22_140 ();
 sg13g2_fill_1 FILLER_22_154 ();
 sg13g2_fill_1 FILLER_22_160 ();
 sg13g2_fill_2 FILLER_22_209 ();
 sg13g2_fill_1 FILLER_22_211 ();
 sg13g2_fill_1 FILLER_22_225 ();
 sg13g2_fill_2 FILLER_22_239 ();
 sg13g2_fill_2 FILLER_22_286 ();
 sg13g2_fill_1 FILLER_22_288 ();
 sg13g2_decap_4 FILLER_22_334 ();
 sg13g2_fill_2 FILLER_22_338 ();
 sg13g2_fill_1 FILLER_22_381 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_4 ();
 sg13g2_decap_8 FILLER_23_9 ();
 sg13g2_fill_2 FILLER_23_16 ();
 sg13g2_fill_2 FILLER_23_76 ();
 sg13g2_fill_1 FILLER_23_78 ();
 sg13g2_fill_1 FILLER_23_92 ();
 sg13g2_fill_2 FILLER_23_97 ();
 sg13g2_fill_2 FILLER_23_149 ();
 sg13g2_fill_1 FILLER_23_151 ();
 sg13g2_decap_4 FILLER_23_177 ();
 sg13g2_fill_2 FILLER_23_244 ();
 sg13g2_fill_2 FILLER_23_256 ();
 sg13g2_fill_1 FILLER_23_272 ();
 sg13g2_fill_2 FILLER_23_343 ();
 sg13g2_fill_1 FILLER_23_353 ();
 sg13g2_fill_1 FILLER_23_381 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_40 ();
 sg13g2_fill_2 FILLER_24_47 ();
 sg13g2_decap_8 FILLER_24_62 ();
 sg13g2_decap_8 FILLER_24_69 ();
 sg13g2_fill_2 FILLER_24_76 ();
 sg13g2_fill_1 FILLER_24_78 ();
 sg13g2_decap_8 FILLER_24_106 ();
 sg13g2_fill_1 FILLER_24_113 ();
 sg13g2_fill_1 FILLER_24_118 ();
 sg13g2_decap_8 FILLER_24_128 ();
 sg13g2_fill_2 FILLER_24_135 ();
 sg13g2_fill_1 FILLER_24_153 ();
 sg13g2_fill_2 FILLER_24_171 ();
 sg13g2_fill_1 FILLER_24_173 ();
 sg13g2_decap_8 FILLER_24_197 ();
 sg13g2_decap_8 FILLER_24_204 ();
 sg13g2_decap_8 FILLER_24_211 ();
 sg13g2_decap_4 FILLER_24_218 ();
 sg13g2_fill_1 FILLER_24_226 ();
 sg13g2_decap_4 FILLER_24_231 ();
 sg13g2_fill_2 FILLER_24_244 ();
 sg13g2_fill_1 FILLER_24_246 ();
 sg13g2_fill_2 FILLER_24_274 ();
 sg13g2_fill_1 FILLER_24_276 ();
 sg13g2_fill_2 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_309 ();
 sg13g2_fill_2 FILLER_24_316 ();
 sg13g2_fill_1 FILLER_24_332 ();
 sg13g2_fill_2 FILLER_24_354 ();
 sg13g2_fill_2 FILLER_24_365 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_fill_2 FILLER_25_36 ();
 sg13g2_fill_1 FILLER_25_38 ();
 sg13g2_decap_4 FILLER_25_66 ();
 sg13g2_fill_1 FILLER_25_80 ();
 sg13g2_fill_2 FILLER_25_107 ();
 sg13g2_fill_1 FILLER_25_109 ();
 sg13g2_fill_2 FILLER_25_120 ();
 sg13g2_decap_4 FILLER_25_135 ();
 sg13g2_fill_1 FILLER_25_139 ();
 sg13g2_fill_2 FILLER_25_162 ();
 sg13g2_decap_8 FILLER_25_176 ();
 sg13g2_decap_8 FILLER_25_183 ();
 sg13g2_fill_2 FILLER_25_190 ();
 sg13g2_fill_1 FILLER_25_229 ();
 sg13g2_decap_4 FILLER_25_234 ();
 sg13g2_fill_2 FILLER_25_247 ();
 sg13g2_fill_1 FILLER_25_249 ();
 sg13g2_fill_1 FILLER_25_273 ();
 sg13g2_fill_1 FILLER_25_289 ();
 sg13g2_fill_2 FILLER_25_367 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_39 ();
 sg13g2_fill_1 FILLER_26_41 ();
 sg13g2_fill_1 FILLER_26_56 ();
 sg13g2_fill_2 FILLER_26_105 ();
 sg13g2_fill_2 FILLER_26_155 ();
 sg13g2_fill_1 FILLER_26_180 ();
 sg13g2_decap_4 FILLER_26_185 ();
 sg13g2_fill_2 FILLER_26_189 ();
 sg13g2_fill_2 FILLER_26_206 ();
 sg13g2_decap_4 FILLER_26_212 ();
 sg13g2_fill_1 FILLER_26_216 ();
 sg13g2_fill_2 FILLER_26_234 ();
 sg13g2_fill_2 FILLER_26_268 ();
 sg13g2_fill_1 FILLER_26_290 ();
 sg13g2_decap_8 FILLER_26_312 ();
 sg13g2_decap_8 FILLER_26_319 ();
 sg13g2_decap_8 FILLER_26_326 ();
 sg13g2_fill_1 FILLER_26_342 ();
 sg13g2_fill_2 FILLER_26_348 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_11 ();
 sg13g2_fill_1 FILLER_27_15 ();
 sg13g2_decap_4 FILLER_27_46 ();
 sg13g2_fill_1 FILLER_27_50 ();
 sg13g2_fill_2 FILLER_27_87 ();
 sg13g2_fill_1 FILLER_27_98 ();
 sg13g2_fill_2 FILLER_27_143 ();
 sg13g2_fill_1 FILLER_27_149 ();
 sg13g2_fill_2 FILLER_27_159 ();
 sg13g2_fill_1 FILLER_27_167 ();
 sg13g2_decap_8 FILLER_27_212 ();
 sg13g2_decap_4 FILLER_27_219 ();
 sg13g2_fill_1 FILLER_27_223 ();
 sg13g2_decap_8 FILLER_27_230 ();
 sg13g2_fill_1 FILLER_27_237 ();
 sg13g2_fill_1 FILLER_27_266 ();
 sg13g2_fill_2 FILLER_27_287 ();
 sg13g2_fill_1 FILLER_27_289 ();
 sg13g2_fill_2 FILLER_27_295 ();
 sg13g2_fill_1 FILLER_27_297 ();
 sg13g2_fill_1 FILLER_27_310 ();
 sg13g2_fill_2 FILLER_27_315 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_28 ();
 sg13g2_decap_4 FILLER_28_39 ();
 sg13g2_decap_4 FILLER_28_47 ();
 sg13g2_fill_2 FILLER_28_51 ();
 sg13g2_fill_2 FILLER_28_80 ();
 sg13g2_fill_1 FILLER_28_82 ();
 sg13g2_fill_2 FILLER_28_114 ();
 sg13g2_fill_1 FILLER_28_116 ();
 sg13g2_fill_2 FILLER_28_127 ();
 sg13g2_fill_1 FILLER_28_129 ();
 sg13g2_fill_1 FILLER_28_167 ();
 sg13g2_decap_4 FILLER_28_195 ();
 sg13g2_fill_2 FILLER_28_199 ();
 sg13g2_decap_8 FILLER_28_218 ();
 sg13g2_fill_1 FILLER_28_225 ();
 sg13g2_decap_4 FILLER_28_239 ();
 sg13g2_decap_8 FILLER_28_247 ();
 sg13g2_fill_2 FILLER_28_254 ();
 sg13g2_fill_1 FILLER_28_256 ();
 sg13g2_fill_2 FILLER_28_297 ();
 sg13g2_fill_1 FILLER_28_299 ();
 sg13g2_fill_2 FILLER_28_341 ();
 sg13g2_fill_2 FILLER_28_379 ();
 sg13g2_decap_4 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_4 ();
 sg13g2_fill_2 FILLER_29_29 ();
 sg13g2_fill_1 FILLER_29_31 ();
 sg13g2_fill_1 FILLER_29_69 ();
 sg13g2_decap_4 FILLER_29_101 ();
 sg13g2_fill_1 FILLER_29_141 ();
 sg13g2_fill_1 FILLER_29_159 ();
 sg13g2_fill_1 FILLER_29_169 ();
 sg13g2_fill_2 FILLER_29_183 ();
 sg13g2_fill_1 FILLER_29_185 ();
 sg13g2_fill_1 FILLER_29_195 ();
 sg13g2_fill_2 FILLER_29_212 ();
 sg13g2_fill_1 FILLER_29_232 ();
 sg13g2_decap_4 FILLER_29_248 ();
 sg13g2_fill_2 FILLER_29_252 ();
 sg13g2_fill_1 FILLER_29_312 ();
 sg13g2_fill_1 FILLER_29_330 ();
 sg13g2_fill_1 FILLER_29_339 ();
 sg13g2_fill_1 FILLER_29_345 ();
 sg13g2_fill_1 FILLER_29_356 ();
 sg13g2_fill_1 FILLER_29_379 ();
 sg13g2_fill_2 FILLER_29_389 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_2 ();
 sg13g2_fill_2 FILLER_30_39 ();
 sg13g2_fill_1 FILLER_30_46 ();
 sg13g2_fill_1 FILLER_30_51 ();
 sg13g2_decap_4 FILLER_30_122 ();
 sg13g2_fill_1 FILLER_30_126 ();
 sg13g2_fill_1 FILLER_30_180 ();
 sg13g2_decap_4 FILLER_30_195 ();
 sg13g2_fill_2 FILLER_30_199 ();
 sg13g2_fill_2 FILLER_30_228 ();
 sg13g2_fill_1 FILLER_30_230 ();
 sg13g2_decap_4 FILLER_30_287 ();
 sg13g2_fill_2 FILLER_30_291 ();
 sg13g2_fill_2 FILLER_30_304 ();
 sg13g2_fill_2 FILLER_30_326 ();
 sg13g2_fill_1 FILLER_30_341 ();
 sg13g2_fill_2 FILLER_30_360 ();
 sg13g2_fill_1 FILLER_30_362 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_127 ();
 sg13g2_fill_2 FILLER_31_156 ();
 sg13g2_fill_2 FILLER_31_173 ();
 sg13g2_decap_8 FILLER_31_209 ();
 sg13g2_fill_2 FILLER_31_245 ();
 sg13g2_fill_1 FILLER_31_247 ();
 sg13g2_decap_4 FILLER_31_252 ();
 sg13g2_fill_1 FILLER_31_265 ();
 sg13g2_decap_4 FILLER_31_282 ();
 sg13g2_fill_1 FILLER_31_286 ();
 sg13g2_fill_2 FILLER_31_303 ();
 sg13g2_fill_1 FILLER_31_305 ();
 sg13g2_fill_2 FILLER_31_323 ();
 sg13g2_fill_1 FILLER_31_325 ();
 sg13g2_fill_2 FILLER_31_332 ();
 sg13g2_fill_2 FILLER_31_360 ();
 sg13g2_fill_1 FILLER_31_398 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_74 ();
 sg13g2_fill_2 FILLER_32_91 ();
 sg13g2_fill_1 FILLER_32_119 ();
 sg13g2_fill_1 FILLER_32_132 ();
 sg13g2_fill_2 FILLER_32_138 ();
 sg13g2_fill_1 FILLER_32_199 ();
 sg13g2_decap_8 FILLER_32_212 ();
 sg13g2_fill_2 FILLER_32_219 ();
 sg13g2_fill_1 FILLER_32_221 ();
 sg13g2_fill_2 FILLER_32_252 ();
 sg13g2_fill_1 FILLER_32_254 ();
 sg13g2_fill_1 FILLER_32_260 ();
 sg13g2_fill_1 FILLER_32_282 ();
 sg13g2_fill_2 FILLER_32_310 ();
 sg13g2_fill_1 FILLER_32_320 ();
 sg13g2_fill_1 FILLER_32_326 ();
 sg13g2_fill_2 FILLER_32_351 ();
 sg13g2_fill_2 FILLER_32_369 ();
 sg13g2_fill_1 FILLER_32_371 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_2 ();
 sg13g2_fill_1 FILLER_33_30 ();
 sg13g2_fill_1 FILLER_33_58 ();
 sg13g2_fill_1 FILLER_33_151 ();
 sg13g2_fill_1 FILLER_33_169 ();
 sg13g2_fill_1 FILLER_33_220 ();
 sg13g2_fill_2 FILLER_33_229 ();
 sg13g2_fill_2 FILLER_33_236 ();
 sg13g2_fill_1 FILLER_33_238 ();
 sg13g2_fill_1 FILLER_33_295 ();
 sg13g2_fill_2 FILLER_33_301 ();
 sg13g2_fill_2 FILLER_33_314 ();
 sg13g2_fill_2 FILLER_33_344 ();
 sg13g2_fill_1 FILLER_33_346 ();
 sg13g2_fill_1 FILLER_33_378 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_44 ();
 sg13g2_fill_2 FILLER_34_119 ();
 sg13g2_fill_2 FILLER_34_161 ();
 sg13g2_fill_2 FILLER_34_204 ();
 sg13g2_fill_2 FILLER_34_222 ();
 sg13g2_fill_1 FILLER_34_224 ();
 sg13g2_fill_2 FILLER_34_230 ();
 sg13g2_fill_2 FILLER_34_240 ();
 sg13g2_fill_1 FILLER_34_307 ();
 sg13g2_fill_2 FILLER_34_327 ();
 sg13g2_fill_1 FILLER_34_357 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_fill_1 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_83 ();
 sg13g2_fill_1 FILLER_35_149 ();
 sg13g2_fill_1 FILLER_35_167 ();
 sg13g2_fill_1 FILLER_35_237 ();
 sg13g2_fill_1 FILLER_35_242 ();
 sg13g2_fill_2 FILLER_35_252 ();
 sg13g2_fill_1 FILLER_35_311 ();
 sg13g2_fill_2 FILLER_35_325 ();
 sg13g2_fill_1 FILLER_35_327 ();
 sg13g2_fill_1 FILLER_35_342 ();
 sg13g2_fill_2 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_4 FILLER_36_7 ();
 sg13g2_fill_2 FILLER_36_58 ();
 sg13g2_fill_2 FILLER_36_67 ();
 sg13g2_fill_1 FILLER_36_123 ();
 sg13g2_fill_1 FILLER_36_169 ();
 sg13g2_fill_2 FILLER_36_206 ();
 sg13g2_fill_1 FILLER_36_302 ();
 sg13g2_fill_1 FILLER_36_321 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_4 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_4 ();
 sg13g2_fill_2 FILLER_37_79 ();
 sg13g2_fill_2 FILLER_37_90 ();
 sg13g2_fill_1 FILLER_37_92 ();
 sg13g2_fill_2 FILLER_37_130 ();
 sg13g2_fill_1 FILLER_37_132 ();
 sg13g2_fill_1 FILLER_37_187 ();
 sg13g2_fill_1 FILLER_37_219 ();
 sg13g2_fill_2 FILLER_37_238 ();
 sg13g2_fill_2 FILLER_37_270 ();
 sg13g2_fill_2 FILLER_37_293 ();
 sg13g2_fill_1 FILLER_37_388 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_7 ();
 sg13g2_fill_1 FILLER_38_9 ();
 sg13g2_fill_2 FILLER_38_88 ();
 sg13g2_fill_1 FILLER_38_143 ();
 sg13g2_fill_2 FILLER_38_190 ();
 sg13g2_fill_2 FILLER_38_201 ();
 sg13g2_fill_1 FILLER_38_203 ();
 sg13g2_fill_2 FILLER_38_208 ();
 sg13g2_fill_1 FILLER_38_210 ();
 sg13g2_fill_2 FILLER_38_305 ();
 assign uio_oe[0] = net14;
 assign uio_oe[1] = net15;
 assign uio_oe[2] = net16;
 assign uio_oe[3] = net17;
 assign uio_oe[4] = net18;
 assign uio_oe[5] = net19;
 assign uio_oe[6] = net275;
 assign uio_oe[7] = net20;
 assign uio_out[0] = net21;
 assign uio_out[1] = net22;
 assign uio_out[2] = net23;
 assign uio_out[3] = net24;
 assign uio_out[4] = net25;
 assign uio_out[5] = net26;
 assign uio_out[7] = net27;
endmodule
