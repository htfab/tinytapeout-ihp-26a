module tt_um_snake_game (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire eat;
 wire failure;
 wire \game_inst.apple_inst.apple_x[0] ;
 wire \game_inst.apple_inst.apple_x[1] ;
 wire \game_inst.apple_inst.apple_x[2] ;
 wire \game_inst.apple_inst.apple_x[3] ;
 wire \game_inst.apple_inst.apple_x[4] ;
 wire \game_inst.apple_inst.apple_y[0] ;
 wire \game_inst.apple_inst.apple_y[1] ;
 wire \game_inst.apple_inst.apple_y[2] ;
 wire \game_inst.apple_inst.apple_y[3] ;
 wire \game_inst.apple_inst.i_snake_valid ;
 wire \game_inst.apple_inst.i_snake_x[0] ;
 wire \game_inst.apple_inst.i_snake_x[1] ;
 wire \game_inst.apple_inst.i_snake_x[2] ;
 wire \game_inst.apple_inst.i_snake_x[3] ;
 wire \game_inst.apple_inst.i_snake_x[4] ;
 wire \game_inst.apple_inst.i_snake_y[0] ;
 wire \game_inst.apple_inst.i_snake_y[1] ;
 wire \game_inst.apple_inst.i_snake_y[2] ;
 wire \game_inst.apple_inst.i_snake_y[3] ;
 wire \game_inst.apple_inst.o_ready ;
 wire \game_inst.apple_inst.random_inst.lfsr4[0] ;
 wire \game_inst.apple_inst.random_inst.lfsr4[1] ;
 wire \game_inst.apple_inst.random_inst.lfsr4[2] ;
 wire \game_inst.apple_inst.random_inst.lfsr4[3] ;
 wire \game_inst.apple_inst.random_inst.lfsr5[0] ;
 wire \game_inst.apple_inst.random_inst.lfsr5[1] ;
 wire \game_inst.apple_inst.random_inst.lfsr5[2] ;
 wire \game_inst.apple_inst.random_inst.lfsr5[3] ;
 wire \game_inst.apple_inst.random_inst.lfsr5[4] ;
 wire \game_inst.apple_inst.test ;
 wire \game_inst.colorblind ;
 wire \game_inst.control_inst.backwards[1] ;
 wire \game_inst.control_inst.dir[0] ;
 wire \game_inst.control_inst.dir[1] ;
 wire \game_inst.control_inst.i_head_dir[0] ;
 wire \game_inst.control_inst.o_start ;
 wire \game_inst.head_x[0] ;
 wire \game_inst.head_x[1] ;
 wire \game_inst.head_x[2] ;
 wire \game_inst.head_x[3] ;
 wire \game_inst.head_x[4] ;
 wire \game_inst.head_y[0] ;
 wire \game_inst.head_y[1] ;
 wire \game_inst.head_y[2] ;
 wire \game_inst.head_y[3] ;
 wire \game_inst.o_success ;
 wire \game_inst.o_vga_hsync ;
 wire \game_inst.o_vga_vsync ;
 wire \game_inst.snake_inst.dir_first[0] ;
 wire \game_inst.snake_inst.dir_first[1] ;
 wire \game_inst.snake_inst.dir_out[0] ;
 wire \game_inst.snake_inst.dir_out[1] ;
 wire \game_inst.snake_inst.length[0] ;
 wire \game_inst.snake_inst.length[1] ;
 wire \game_inst.snake_inst.length[2] ;
 wire \game_inst.snake_inst.length[3] ;
 wire \game_inst.snake_inst.length[4] ;
 wire \game_inst.snake_inst.length[5] ;
 wire \game_inst.snake_inst.length[6] ;
 wire \game_inst.snake_inst.length[7] ;
 wire \game_inst.snake_inst.pos[0] ;
 wire \game_inst.snake_inst.pos[1] ;
 wire \game_inst.snake_inst.pos[2] ;
 wire \game_inst.snake_inst.pos[3] ;
 wire \game_inst.snake_inst.pos[4] ;
 wire \game_inst.snake_inst.pos[5] ;
 wire \game_inst.snake_inst.pos[6] ;
 wire \game_inst.snake_inst.pos[7] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[100][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[100][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[101][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[101][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[102][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[102][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[103][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[103][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[104][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[104][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[105][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[105][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[106][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[106][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[107][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[107][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[108][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[108][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[109][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[109][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[10][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[10][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[110][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[110][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[111][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[111][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[112][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[112][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[113][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[113][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[114][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[114][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[115][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[115][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[116][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[116][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[117][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[117][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[118][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[118][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[119][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[119][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[11][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[11][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[120][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[120][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[121][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[121][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[122][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[122][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[123][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[123][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[124][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[124][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[125][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[125][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[126][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[126][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[127][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[127][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[128][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[128][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[129][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[129][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[12][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[12][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[130][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[130][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[131][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[131][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[132][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[132][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[133][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[133][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[134][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[134][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[135][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[135][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[136][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[136][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[137][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[137][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[138][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[138][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[139][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[139][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[13][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[13][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[140][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[140][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[141][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[141][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[142][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[142][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[143][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[143][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[144][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[144][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[145][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[145][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[146][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[146][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[147][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[147][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[148][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[148][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[149][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[149][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[14][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[14][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[150][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[150][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[151][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[151][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[152][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[152][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[153][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[153][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[154][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[154][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[155][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[155][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[156][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[156][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[157][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[157][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[158][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[158][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[159][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[159][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[15][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[15][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[160][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[160][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[161][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[161][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[162][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[162][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[163][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[163][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[164][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[164][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[165][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[165][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[166][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[166][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[167][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[167][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[168][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[168][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[169][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[169][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[16][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[16][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[170][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[170][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[171][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[171][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[172][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[172][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[173][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[173][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[174][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[174][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[175][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[175][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[176][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[176][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[177][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[177][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[178][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[178][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[179][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[179][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[17][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[17][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[180][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[180][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[181][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[181][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[182][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[182][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[183][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[183][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[184][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[184][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[185][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[185][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[186][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[186][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[187][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[187][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[188][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[188][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[189][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[189][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[18][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[18][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[190][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[190][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[191][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[191][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[192][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[192][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[193][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[193][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[194][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[194][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[195][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[195][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[196][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[196][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[197][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[197][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[198][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[198][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[199][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[199][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[19][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[19][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[1][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[1][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[200][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[200][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[201][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[201][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[202][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[202][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[203][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[203][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[204][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[204][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[205][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[205][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[206][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[206][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[207][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[207][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[208][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[208][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[209][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[209][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[20][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[20][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[210][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[210][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[211][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[211][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[212][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[212][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[213][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[213][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[214][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[214][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[215][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[215][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[216][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[216][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[217][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[217][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[218][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[218][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[219][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[219][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[21][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[21][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[220][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[220][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[221][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[221][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[222][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[222][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[223][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[223][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[224][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[224][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[225][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[225][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[226][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[226][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[227][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[227][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[228][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[228][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[229][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[229][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[22][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[22][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[230][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[230][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[231][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[231][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[232][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[232][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[23][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[23][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[24][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[24][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[25][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[25][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[26][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[26][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[27][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[27][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[28][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[28][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[29][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[29][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[2][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[2][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[30][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[30][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[31][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[31][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[32][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[32][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[33][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[33][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[34][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[34][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[35][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[35][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[36][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[36][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[37][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[37][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[38][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[38][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[39][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[39][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[3][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[3][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[40][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[40][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[41][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[41][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[42][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[42][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[43][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[43][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[44][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[44][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[45][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[45][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[46][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[46][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[47][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[47][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[48][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[48][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[49][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[49][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[4][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[4][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[50][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[50][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[51][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[51][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[52][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[52][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[53][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[53][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[54][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[54][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[55][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[55][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[56][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[56][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[57][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[57][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[58][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[58][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[59][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[59][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[5][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[5][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[60][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[60][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[61][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[61][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[62][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[62][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[63][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[63][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[64][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[64][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[65][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[65][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[66][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[66][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[67][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[67][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[68][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[68][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[69][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[69][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[6][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[6][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[70][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[70][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[71][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[71][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[72][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[72][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[73][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[73][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[74][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[74][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[75][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[75][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[76][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[76][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[77][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[77][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[78][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[78][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[79][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[79][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[7][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[7][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[80][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[80][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[81][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[81][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[82][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[82][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[83][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[83][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[84][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[84][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[85][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[85][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[86][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[86][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[87][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[87][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[88][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[88][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[89][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[89][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[8][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[8][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[90][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[90][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[91][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[91][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[92][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[92][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[93][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[93][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[94][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[94][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[95][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[95][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[96][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[96][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[97][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[97][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[98][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[98][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[99][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[99][1] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[9][0] ;
 wire \game_inst.snake_inst.shiftreg_inst.memory[9][1] ;
 wire \game_inst.tick ;
 wire \game_inst.tickgen_inst.counter[0] ;
 wire \game_inst.tickgen_inst.counter[1] ;
 wire \game_inst.tickgen_inst.counter[2] ;
 wire \game_inst.tickgen_inst.counter[3] ;
 wire \game_inst.tickgen_inst.counter[4] ;
 wire \game_inst.tickgen_inst.counter_max[0] ;
 wire \game_inst.tickgen_inst.counter_max[1] ;
 wire \game_inst.tickgen_inst.counter_max[2] ;
 wire \game_inst.tickgen_inst.counter_max[3] ;
 wire \game_inst.tickgen_inst.counter_max[4] ;
 wire \game_inst.tickgen_inst.i_vsync ;
 wire \game_inst.tickgen_inst.prev_user_input ;
 wire \game_inst.tickgen_inst.prev_vsync ;
 wire \game_inst.vga_inst.pos_counter[0] ;
 wire \game_inst.vga_inst.pos_counter[1] ;
 wire \game_inst.vga_inst.px[0] ;
 wire \game_inst.vga_inst.px[1] ;
 wire \game_inst.vga_inst.px[2] ;
 wire \game_inst.vga_inst.px[3] ;
 wire \game_inst.vga_inst.px[4] ;
 wire \game_inst.vga_inst.px[5] ;
 wire \game_inst.vga_inst.px[6] ;
 wire \game_inst.vga_inst.px[7] ;
 wire \game_inst.vga_inst.px[8] ;
 wire \game_inst.vga_inst.px[9] ;
 wire \game_inst.vga_inst.py[0] ;
 wire \game_inst.vga_inst.py[1] ;
 wire \game_inst.vga_inst.py[2] ;
 wire \game_inst.vga_inst.py[3] ;
 wire \game_inst.vga_inst.py[4] ;
 wire \game_inst.vga_inst.py[5] ;
 wire \game_inst.vga_inst.py[6] ;
 wire \game_inst.vga_inst.py[7] ;
 wire \game_inst.vga_inst.py[8] ;
 wire \game_inst.vga_inst.py[9] ;
 wire \game_inst.vga_inst.row_buffer[0][0] ;
 wire \game_inst.vga_inst.row_buffer[0][1] ;
 wire \game_inst.vga_inst.row_buffer[10][0] ;
 wire \game_inst.vga_inst.row_buffer[10][1] ;
 wire \game_inst.vga_inst.row_buffer[11][0] ;
 wire \game_inst.vga_inst.row_buffer[11][1] ;
 wire \game_inst.vga_inst.row_buffer[12][0] ;
 wire \game_inst.vga_inst.row_buffer[12][1] ;
 wire \game_inst.vga_inst.row_buffer[13][0] ;
 wire \game_inst.vga_inst.row_buffer[13][1] ;
 wire \game_inst.vga_inst.row_buffer[14][0] ;
 wire \game_inst.vga_inst.row_buffer[14][1] ;
 wire \game_inst.vga_inst.row_buffer[15][0] ;
 wire \game_inst.vga_inst.row_buffer[15][1] ;
 wire \game_inst.vga_inst.row_buffer[16][0] ;
 wire \game_inst.vga_inst.row_buffer[16][1] ;
 wire \game_inst.vga_inst.row_buffer[17][0] ;
 wire \game_inst.vga_inst.row_buffer[17][1] ;
 wire \game_inst.vga_inst.row_buffer[1][0] ;
 wire \game_inst.vga_inst.row_buffer[1][1] ;
 wire \game_inst.vga_inst.row_buffer[2][0] ;
 wire \game_inst.vga_inst.row_buffer[2][1] ;
 wire \game_inst.vga_inst.row_buffer[3][0] ;
 wire \game_inst.vga_inst.row_buffer[3][1] ;
 wire \game_inst.vga_inst.row_buffer[4][0] ;
 wire \game_inst.vga_inst.row_buffer[4][1] ;
 wire \game_inst.vga_inst.row_buffer[5][0] ;
 wire \game_inst.vga_inst.row_buffer[5][1] ;
 wire \game_inst.vga_inst.row_buffer[6][0] ;
 wire \game_inst.vga_inst.row_buffer[6][1] ;
 wire \game_inst.vga_inst.row_buffer[7][0] ;
 wire \game_inst.vga_inst.row_buffer[7][1] ;
 wire \game_inst.vga_inst.row_buffer[8][0] ;
 wire \game_inst.vga_inst.row_buffer[8][1] ;
 wire \game_inst.vga_inst.row_buffer[9][0] ;
 wire \game_inst.vga_inst.row_buffer[9][1] ;
 wire net669;
 wire net670;
 wire clknet_leaf_0_clk;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;

 sg13g2_inv_1 _1333_ (.Y(_0161_),
    .A(net1310));
 sg13g2_inv_1 _1334_ (.Y(_0162_),
    .A(\game_inst.tickgen_inst.counter[1] ));
 sg13g2_inv_1 _1335_ (.Y(_0163_),
    .A(\game_inst.tickgen_inst.counter[0] ));
 sg13g2_inv_1 _1336_ (.Y(_0164_),
    .A(net1144));
 sg13g2_inv_1 _1337_ (.Y(_0165_),
    .A(\game_inst.tickgen_inst.counter_max[1] ));
 sg13g2_inv_1 _1338_ (.Y(_0166_),
    .A(net1285));
 sg13g2_inv_1 _1339_ (.Y(_0167_),
    .A(net1148));
 sg13g2_inv_1 _1340_ (.Y(_0168_),
    .A(\game_inst.colorblind ));
 sg13g2_inv_1 _1341_ (.Y(_0169_),
    .A(\game_inst.apple_inst.i_snake_valid ));
 sg13g2_inv_2 _1342_ (.Y(_0170_),
    .A(net1283));
 sg13g2_inv_1 _1343_ (.Y(_0171_),
    .A(net119));
 sg13g2_inv_1 _1344_ (.Y(_0172_),
    .A(net120));
 sg13g2_inv_1 _1345_ (.Y(_0173_),
    .A(\game_inst.head_y[0] ));
 sg13g2_inv_2 _1346_ (.Y(_0174_),
    .A(net1284));
 sg13g2_inv_1 _1347_ (.Y(_0175_),
    .A(net121));
 sg13g2_inv_2 _1348_ (.Y(_0176_),
    .A(\game_inst.head_x[1] ));
 sg13g2_inv_2 _1349_ (.Y(_0177_),
    .A(\game_inst.head_x[0] ));
 sg13g2_inv_2 _1350_ (.Y(_0178_),
    .A(net1325));
 sg13g2_inv_1 _1351_ (.Y(_0179_),
    .A(net1213));
 sg13g2_inv_1 _1352_ (.Y(_0180_),
    .A(net1154));
 sg13g2_inv_1 _1353_ (.Y(_0181_),
    .A(net1223));
 sg13g2_inv_1 _1354_ (.Y(_0182_),
    .A(net1164));
 sg13g2_inv_1 _1355_ (.Y(_0183_),
    .A(net1162));
 sg13g2_inv_1 _1356_ (.Y(_0184_),
    .A(net1192));
 sg13g2_inv_1 _1357_ (.Y(_0185_),
    .A(net1150));
 sg13g2_inv_2 _1358_ (.Y(_0186_),
    .A(\game_inst.vga_inst.py[7] ));
 sg13g2_inv_2 _1359_ (.Y(_0187_),
    .A(net122));
 sg13g2_inv_1 _1360_ (.Y(_0188_),
    .A(\game_inst.snake_inst.pos[1] ));
 sg13g2_inv_1 _1361_ (.Y(_0189_),
    .A(net1168));
 sg13g2_inv_1 _1362_ (.Y(_0190_),
    .A(\game_inst.snake_inst.pos[6] ));
 sg13g2_inv_1 _1363_ (.Y(_0191_),
    .A(net1257));
 sg13g2_inv_1 _1364_ (.Y(_0192_),
    .A(net1171));
 sg13g2_inv_1 _1365_ (.Y(_0193_),
    .A(net1));
 sg13g2_inv_1 _1366_ (.Y(_0194_),
    .A(\game_inst.snake_inst.length[0] ));
 sg13g2_inv_1 _1367_ (.Y(_0195_),
    .A(\game_inst.snake_inst.length[1] ));
 sg13g2_inv_1 _1368_ (.Y(_0196_),
    .A(\game_inst.snake_inst.length[3] ));
 sg13g2_inv_1 _1369_ (.Y(_0197_),
    .A(net1322));
 sg13g2_inv_1 _1370_ (.Y(_0198_),
    .A(\game_inst.snake_inst.length[6] ));
 sg13g2_inv_1 _1371_ (.Y(_0199_),
    .A(\game_inst.apple_inst.apple_x[0] ));
 sg13g2_inv_2 _1372_ (.Y(_0200_),
    .A(net117));
 sg13g2_inv_1 _1373_ (.Y(_0201_),
    .A(net1323));
 sg13g2_inv_1 _1374_ (.Y(_0202_),
    .A(\game_inst.apple_inst.apple_x[2] ));
 sg13g2_inv_2 _1375_ (.Y(_0203_),
    .A(net1309));
 sg13g2_inv_1 _1376_ (.Y(_0204_),
    .A(\game_inst.apple_inst.apple_x[3] ));
 sg13g2_inv_2 _1377_ (.Y(_0205_),
    .A(net1318));
 sg13g2_inv_1 _1378_ (.Y(_0206_),
    .A(\game_inst.apple_inst.apple_x[4] ));
 sg13g2_inv_2 _1379_ (.Y(_0207_),
    .A(net1313));
 sg13g2_inv_1 _1380_ (.Y(_0208_),
    .A(\game_inst.apple_inst.i_snake_y[0] ));
 sg13g2_inv_1 _1381_ (.Y(_0209_),
    .A(\game_inst.apple_inst.apple_y[0] ));
 sg13g2_inv_2 _1382_ (.Y(_0210_),
    .A(net1307));
 sg13g2_inv_1 _1383_ (.Y(_0211_),
    .A(net1273));
 sg13g2_inv_1 _1384_ (.Y(_0212_),
    .A(\game_inst.apple_inst.apple_y[2] ));
 sg13g2_inv_1 _1385_ (.Y(_0213_),
    .A(net1294));
 sg13g2_inv_2 _1386_ (.Y(_0214_),
    .A(net128));
 sg13g2_inv_2 _1387_ (.Y(_0215_),
    .A(\game_inst.vga_inst.px[6] ));
 sg13g2_inv_4 _1388_ (.A(net1327),
    .Y(_0216_));
 sg13g2_inv_1 _1389_ (.Y(_0217_),
    .A(net123));
 sg13g2_inv_1 _1390_ (.Y(_0218_),
    .A(\game_inst.vga_inst.row_buffer[11][0] ));
 sg13g2_inv_1 _1391_ (.Y(_0219_),
    .A(\game_inst.vga_inst.row_buffer[9][1] ));
 sg13g2_nor2b_1 _1392_ (.A(net6),
    .B_N(net1140),
    .Y(\game_inst.tickgen_inst.i_vsync ));
 sg13g2_xor2_1 _1393_ (.B(\game_inst.apple_inst.apple_y[3] ),
    .A(\game_inst.apple_inst.i_snake_y[3] ),
    .X(_0220_));
 sg13g2_xnor2_1 _1394_ (.Y(_0221_),
    .A(\game_inst.apple_inst.i_snake_y[1] ),
    .B(\game_inst.apple_inst.apple_y[1] ));
 sg13g2_xnor2_1 _1395_ (.Y(_0222_),
    .A(\game_inst.apple_inst.i_snake_y[2] ),
    .B(\game_inst.apple_inst.apple_y[2] ));
 sg13g2_a22oi_1 _1396_ (.Y(_0223_),
    .B1(\game_inst.apple_inst.apple_x[3] ),
    .B2(_0205_),
    .A2(\game_inst.apple_inst.i_snake_x[2] ),
    .A1(_0202_));
 sg13g2_xor2_1 _1397_ (.B(\game_inst.apple_inst.i_snake_x[1] ),
    .A(\game_inst.apple_inst.apple_x[1] ),
    .X(_0224_));
 sg13g2_a22oi_1 _1398_ (.Y(_0225_),
    .B1(\game_inst.apple_inst.i_snake_y[0] ),
    .B2(_0209_),
    .A2(_0203_),
    .A1(\game_inst.apple_inst.apple_x[2] ));
 sg13g2_a221oi_1 _1399_ (.B2(\game_inst.apple_inst.i_snake_x[4] ),
    .C1(_0224_),
    .B1(_0206_),
    .A1(\game_inst.apple_inst.apple_x[0] ),
    .Y(_0226_),
    .A2(_0200_));
 sg13g2_a221oi_1 _1400_ (.B2(_0207_),
    .C1(_0220_),
    .B1(\game_inst.apple_inst.apple_x[4] ),
    .A1(_0199_),
    .Y(_0227_),
    .A2(net117));
 sg13g2_nand4_1 _1401_ (.B(_0225_),
    .C(_0226_),
    .A(_0223_),
    .Y(_0228_),
    .D(_0227_));
 sg13g2_a22oi_1 _1402_ (.Y(_0229_),
    .B1(_0208_),
    .B2(\game_inst.apple_inst.apple_y[0] ),
    .A2(\game_inst.apple_inst.i_snake_x[3] ),
    .A1(_0204_));
 sg13g2_nand3_1 _1403_ (.B(_0222_),
    .C(_0229_),
    .A(_0221_),
    .Y(_0230_));
 sg13g2_nor4_1 _1404_ (.A(net1168),
    .B(\game_inst.snake_inst.pos[5] ),
    .C(\game_inst.snake_inst.pos[6] ),
    .D(\game_inst.snake_inst.pos[7] ),
    .Y(_0231_));
 sg13g2_nor2_1 _1405_ (.A(net1305),
    .B(net1206),
    .Y(_0232_));
 sg13g2_nor4_1 _1406_ (.A(\game_inst.snake_inst.pos[1] ),
    .B(\game_inst.snake_inst.pos[0] ),
    .C(\game_inst.snake_inst.pos[2] ),
    .D(\game_inst.snake_inst.pos[3] ),
    .Y(_0233_));
 sg13g2_and2_1 _1407_ (.A(_0231_),
    .B(_0233_),
    .X(_0234_));
 sg13g2_nand2_2 _1408_ (.Y(_0235_),
    .A(_0231_),
    .B(_0233_));
 sg13g2_nand2_1 _1409_ (.Y(_0236_),
    .A(net1180),
    .B(_0234_));
 sg13g2_nor3_2 _1410_ (.A(_0228_),
    .B(_0230_),
    .C(_0236_),
    .Y(eat));
 sg13g2_and2_1 _1411_ (.A(\game_inst.vga_inst.py[7] ),
    .B(\game_inst.vga_inst.py[6] ),
    .X(_0237_));
 sg13g2_nand2_1 _1412_ (.Y(_0238_),
    .A(\game_inst.vga_inst.py[8] ),
    .B(_0237_));
 sg13g2_nand3_1 _1413_ (.B(net122),
    .C(_0237_),
    .A(net1271),
    .Y(_0239_));
 sg13g2_and2_1 _1414_ (.A(net1166),
    .B(net1182),
    .X(_0240_));
 sg13g2_nand2b_1 _1415_ (.Y(_0241_),
    .B(net1166),
    .A_N(net1225));
 sg13g2_nand2b_1 _1416_ (.Y(_0242_),
    .B(net1185),
    .A_N(net1217));
 sg13g2_nor4_2 _1417_ (.A(net1272),
    .B(_0240_),
    .C(_0241_),
    .Y(_0002_),
    .D(_0242_));
 sg13g2_nor2_1 _1418_ (.A(net129),
    .B(net127),
    .Y(_0243_));
 sg13g2_or2_1 _1419_ (.X(_0244_),
    .B(net127),
    .A(net129));
 sg13g2_nor2_1 _1420_ (.A(net1289),
    .B(net114),
    .Y(_0245_));
 sg13g2_nor2_2 _1421_ (.A(net116),
    .B(net115),
    .Y(_0246_));
 sg13g2_nand2_1 _1422_ (.Y(_0247_),
    .A(net129),
    .B(net127));
 sg13g2_a21oi_1 _1423_ (.A1(net1289),
    .A2(net111),
    .Y(_0248_),
    .B1(_0245_));
 sg13g2_and4_1 _1424_ (.A(net126),
    .B(net1327),
    .C(_0217_),
    .D(_0248_),
    .X(_0001_));
 sg13g2_or2_1 _1425_ (.X(_0249_),
    .B(net123),
    .A(net125));
 sg13g2_a21oi_1 _1426_ (.A1(\game_inst.vga_inst.px[9] ),
    .A2(_0249_),
    .Y(_0250_),
    .B1(\game_inst.vga_inst.py[9] ));
 sg13g2_nand2_2 _1427_ (.Y(_0251_),
    .A(_0239_),
    .B(_0250_));
 sg13g2_inv_1 _1428_ (.Y(_0252_),
    .A(_0251_));
 sg13g2_xnor2_1 _1429_ (.Y(_0253_),
    .A(\game_inst.head_x[2] ),
    .B(net125));
 sg13g2_nor2_1 _1430_ (.A(net7),
    .B(net135),
    .Y(_0254_));
 sg13g2_nand2b_1 _1431_ (.Y(_0255_),
    .B(net139),
    .A_N(net7));
 sg13g2_xor2_1 _1432_ (.B(\game_inst.vga_inst.py[6] ),
    .A(net120),
    .X(_0256_));
 sg13g2_xnor2_1 _1433_ (.Y(_0257_),
    .A(\game_inst.head_y[3] ),
    .B(\game_inst.vga_inst.py[8] ));
 sg13g2_a22oi_1 _1434_ (.Y(_0258_),
    .B1(_0217_),
    .B2(net121),
    .A2(_0216_),
    .A1(\game_inst.head_x[4] ));
 sg13g2_a22oi_1 _1435_ (.Y(_0259_),
    .B1(_0187_),
    .B2(\game_inst.head_y[0] ),
    .A2(_0186_),
    .A1(net119));
 sg13g2_nand4_1 _1436_ (.B(_0257_),
    .C(_0258_),
    .A(_0253_),
    .Y(_0260_),
    .D(_0259_));
 sg13g2_a221oi_1 _1437_ (.B2(\game_inst.head_x[1] ),
    .C1(net130),
    .B1(_0215_),
    .A1(_0173_),
    .Y(_0261_),
    .A2(net122));
 sg13g2_a221oi_1 _1438_ (.B2(_0175_),
    .C1(_0256_),
    .B1(net123),
    .A1(_0177_),
    .Y(_0262_),
    .A2(net128));
 sg13g2_a22oi_1 _1439_ (.Y(_0263_),
    .B1(\game_inst.vga_inst.px[9] ),
    .B2(_0174_),
    .A2(\game_inst.vga_inst.py[7] ),
    .A1(_0171_));
 sg13g2_a22oi_1 _1440_ (.Y(_0264_),
    .B1(net127),
    .B2(_0176_),
    .A2(_0214_),
    .A1(\game_inst.head_x[0] ));
 sg13g2_nand4_1 _1441_ (.B(_0262_),
    .C(_0263_),
    .A(_0261_),
    .Y(_0265_),
    .D(_0264_));
 sg13g2_or2_1 _1442_ (.X(_0266_),
    .B(_0265_),
    .A(_0260_));
 sg13g2_and2_1 _1443_ (.A(_0252_),
    .B(_0266_),
    .X(_0267_));
 sg13g2_nor2_2 _1444_ (.A(net125),
    .B(net114),
    .Y(_0268_));
 sg13g2_nor2_1 _1445_ (.A(net114),
    .B(_0249_),
    .Y(_0269_));
 sg13g2_o21ai_1 _1446_ (.B1(_0216_),
    .Y(_0270_),
    .A1(net114),
    .A2(_0249_));
 sg13g2_o21ai_1 _1447_ (.B1(\game_inst.vga_inst.px[9] ),
    .Y(_0271_),
    .A1(_0247_),
    .A2(_0249_));
 sg13g2_nor3_1 _1448_ (.A(\game_inst.vga_inst.py[8] ),
    .B(\game_inst.vga_inst.py[7] ),
    .C(\game_inst.vga_inst.py[6] ),
    .Y(_0272_));
 sg13g2_a21o_1 _1449_ (.A2(_0237_),
    .A1(\game_inst.vga_inst.py[8] ),
    .B1(_0272_),
    .X(_0273_));
 sg13g2_a22oi_1 _1450_ (.Y(_0274_),
    .B1(_0273_),
    .B2(_0187_),
    .A2(_0271_),
    .A1(_0270_));
 sg13g2_nor2b_2 _1451_ (.A(failure),
    .B_N(\game_inst.o_success ),
    .Y(_0275_));
 sg13g2_nor2_2 _1452_ (.A(_0191_),
    .B(\game_inst.o_success ),
    .Y(_0276_));
 sg13g2_nor2_1 _1453_ (.A(_0275_),
    .B(_0276_),
    .Y(_0277_));
 sg13g2_o21ai_1 _1454_ (.B1(_0267_),
    .Y(_0278_),
    .A1(_0274_),
    .A2(_0277_));
 sg13g2_nor2_1 _1455_ (.A(\game_inst.vga_inst.row_buffer[3][0] ),
    .B(net114),
    .Y(_0279_));
 sg13g2_a221oi_1 _1456_ (.B2(net115),
    .C1(net125),
    .B1(\game_inst.vga_inst.row_buffer[0][0] ),
    .A1(net116),
    .Y(_0280_),
    .A2(\game_inst.vga_inst.row_buffer[1][0] ));
 sg13g2_a21oi_1 _1457_ (.A1(\game_inst.vga_inst.row_buffer[2][0] ),
    .A2(net111),
    .Y(_0281_),
    .B1(net124));
 sg13g2_o21ai_1 _1458_ (.B1(_0281_),
    .Y(_0282_),
    .A1(_0279_),
    .A2(_0280_));
 sg13g2_xnor2_1 _1459_ (.Y(_0283_),
    .A(net124),
    .B(_0268_));
 sg13g2_xor2_1 _1460_ (.B(_0268_),
    .A(net124),
    .X(_0284_));
 sg13g2_nand2b_1 _1461_ (.Y(_0285_),
    .B(net124),
    .A_N(\game_inst.vga_inst.row_buffer[7][0] ));
 sg13g2_nand2_2 _1462_ (.Y(_0286_),
    .A(net126),
    .B(net114));
 sg13g2_a22oi_1 _1463_ (.Y(_0287_),
    .B1(\game_inst.vga_inst.row_buffer[4][0] ),
    .B2(net115),
    .A2(\game_inst.vga_inst.row_buffer[5][0] ),
    .A1(net116));
 sg13g2_nand2b_1 _1464_ (.Y(_0288_),
    .B(_0287_),
    .A_N(_0286_));
 sg13g2_a22oi_1 _1465_ (.Y(_0289_),
    .B1(_0285_),
    .B2(_0288_),
    .A2(net111),
    .A1(\game_inst.vga_inst.row_buffer[6][0] ));
 sg13g2_nor2_1 _1466_ (.A(_0284_),
    .B(_0289_),
    .Y(_0290_));
 sg13g2_a22oi_1 _1467_ (.Y(_0291_),
    .B1(\game_inst.vga_inst.row_buffer[12][0] ),
    .B2(net129),
    .A2(\game_inst.vga_inst.row_buffer[13][0] ),
    .A1(net127));
 sg13g2_nor2_1 _1468_ (.A(net111),
    .B(_0291_),
    .Y(_0292_));
 sg13g2_nand2b_2 _1469_ (.Y(_0293_),
    .B(_0286_),
    .A_N(_0268_));
 sg13g2_a221oi_1 _1470_ (.B2(\game_inst.vga_inst.row_buffer[14][0] ),
    .C1(_0292_),
    .B1(net111),
    .A1(\game_inst.vga_inst.row_buffer[15][0] ),
    .Y(_0294_),
    .A2(_0243_));
 sg13g2_a21oi_1 _1471_ (.A1(net115),
    .A2(\game_inst.vga_inst.row_buffer[8][0] ),
    .Y(_0295_),
    .B1(net116));
 sg13g2_a21oi_1 _1472_ (.A1(_0218_),
    .A2(_0243_),
    .Y(_0296_),
    .B1(_0295_));
 sg13g2_o21ai_1 _1473_ (.B1(_0296_),
    .Y(_0297_),
    .A1(net115),
    .A2(\game_inst.vga_inst.row_buffer[9][0] ));
 sg13g2_a21oi_1 _1474_ (.A1(\game_inst.vga_inst.row_buffer[10][0] ),
    .A2(_0246_),
    .Y(_0298_),
    .B1(_0293_));
 sg13g2_a22oi_1 _1475_ (.Y(_0299_),
    .B1(_0297_),
    .B2(_0298_),
    .A2(_0294_),
    .A1(_0293_));
 sg13g2_xnor2_1 _1476_ (.Y(_0300_),
    .A(_0216_),
    .B(_0269_));
 sg13g2_a221oi_1 _1477_ (.B2(_0284_),
    .C1(_0300_),
    .B1(_0299_),
    .A1(_0282_),
    .Y(_0301_),
    .A2(_0290_));
 sg13g2_and2_1 _1478_ (.A(net128),
    .B(\game_inst.vga_inst.row_buffer[16][0] ),
    .X(_0302_));
 sg13g2_a21oi_1 _1479_ (.A1(net116),
    .A2(\game_inst.vga_inst.row_buffer[17][0] ),
    .Y(_0303_),
    .B1(_0302_));
 sg13g2_nand2_1 _1480_ (.Y(_0304_),
    .A(_0300_),
    .B(_0303_));
 sg13g2_xor2_1 _1481_ (.B(\game_inst.apple_inst.apple_y[3] ),
    .A(\game_inst.vga_inst.py[8] ),
    .X(_0305_));
 sg13g2_nor2b_1 _1482_ (.A(\game_inst.apple_inst.apple_x[2] ),
    .B_N(net125),
    .Y(_0306_));
 sg13g2_nand2b_1 _1483_ (.Y(_0307_),
    .B(\game_inst.apple_inst.apple_x[2] ),
    .A_N(net126));
 sg13g2_o21ai_1 _1484_ (.B1(_0307_),
    .Y(_0308_),
    .A1(_0204_),
    .A2(net123));
 sg13g2_a221oi_1 _1485_ (.B2(_0204_),
    .C1(_0308_),
    .B1(net123),
    .A1(_0187_),
    .Y(_0309_),
    .A2(\game_inst.apple_inst.apple_y[0] ));
 sg13g2_xor2_1 _1486_ (.B(\game_inst.apple_inst.apple_y[1] ),
    .A(\game_inst.vga_inst.py[6] ),
    .X(_0310_));
 sg13g2_a221oi_1 _1487_ (.B2(\game_inst.vga_inst.py[7] ),
    .C1(_0310_),
    .B1(_0212_),
    .A1(net122),
    .Y(_0311_),
    .A2(_0209_));
 sg13g2_a221oi_1 _1488_ (.B2(_0199_),
    .C1(_0306_),
    .B1(net128),
    .A1(_0186_),
    .Y(_0312_),
    .A2(\game_inst.apple_inst.apple_y[2] ));
 sg13g2_xor2_1 _1489_ (.B(net127),
    .A(\game_inst.apple_inst.apple_x[1] ),
    .X(_0313_));
 sg13g2_o21ai_1 _1490_ (.B1(\game_inst.apple_inst.o_ready ),
    .Y(_0314_),
    .A1(_0199_),
    .A2(\game_inst.vga_inst.px[5] ));
 sg13g2_xor2_1 _1491_ (.B(\game_inst.vga_inst.px[9] ),
    .A(\game_inst.apple_inst.apple_x[4] ),
    .X(_0315_));
 sg13g2_nor4_1 _1492_ (.A(_0305_),
    .B(_0313_),
    .C(_0314_),
    .D(_0315_),
    .Y(_0316_));
 sg13g2_nand4_1 _1493_ (.B(_0311_),
    .C(_0312_),
    .A(_0309_),
    .Y(_0317_),
    .D(_0316_));
 sg13g2_nand2_1 _1494_ (.Y(_0318_),
    .A(_0304_),
    .B(_0317_));
 sg13g2_o21ai_1 _1495_ (.B1(_0274_),
    .Y(_0319_),
    .A1(_0301_),
    .A2(_0318_));
 sg13g2_nor2b_1 _1496_ (.A(_0278_),
    .B_N(_0319_),
    .Y(_0320_));
 sg13g2_inv_1 _1497_ (.Y(_0321_),
    .A(_0320_));
 sg13g2_nand2b_1 _1498_ (.Y(_0322_),
    .B(_0267_),
    .A_N(_0274_));
 sg13g2_nor3_1 _1499_ (.A(_0275_),
    .B(_0276_),
    .C(_0322_),
    .Y(_0323_));
 sg13g2_nand2_1 _1500_ (.Y(_0324_),
    .A(_0168_),
    .B(_0323_));
 sg13g2_o21ai_1 _1501_ (.B1(_0324_),
    .Y(uo_out[6]),
    .A1(_0168_),
    .A2(_0321_));
 sg13g2_nand2_1 _1502_ (.Y(_0325_),
    .A(\game_inst.vga_inst.row_buffer[6][1] ),
    .B(_0246_));
 sg13g2_nor2b_1 _1503_ (.A(\game_inst.vga_inst.row_buffer[7][1] ),
    .B_N(net124),
    .Y(_0326_));
 sg13g2_a221oi_1 _1504_ (.B2(net115),
    .C1(_0286_),
    .B1(\game_inst.vga_inst.row_buffer[4][1] ),
    .A1(net116),
    .Y(_0327_),
    .A2(\game_inst.vga_inst.row_buffer[5][1] ));
 sg13g2_o21ai_1 _1505_ (.B1(_0325_),
    .Y(_0328_),
    .A1(_0326_),
    .A2(_0327_));
 sg13g2_nor2_1 _1506_ (.A(\game_inst.vga_inst.row_buffer[3][1] ),
    .B(net114),
    .Y(_0329_));
 sg13g2_a221oi_1 _1507_ (.B2(net115),
    .C1(net125),
    .B1(\game_inst.vga_inst.row_buffer[0][1] ),
    .A1(net116),
    .Y(_0330_),
    .A2(\game_inst.vga_inst.row_buffer[1][1] ));
 sg13g2_a21oi_1 _1508_ (.A1(\game_inst.vga_inst.row_buffer[2][1] ),
    .A2(net111),
    .Y(_0331_),
    .B1(net124));
 sg13g2_o21ai_1 _1509_ (.B1(_0331_),
    .Y(_0332_),
    .A1(_0329_),
    .A2(_0330_));
 sg13g2_nand3_1 _1510_ (.B(_0328_),
    .C(_0332_),
    .A(_0283_),
    .Y(_0333_));
 sg13g2_o21ai_1 _1511_ (.B1(net115),
    .Y(_0334_),
    .A1(net116),
    .A2(\game_inst.vga_inst.row_buffer[8][1] ));
 sg13g2_o21ai_1 _1512_ (.B1(_0334_),
    .Y(_0335_),
    .A1(net128),
    .A2(_0219_));
 sg13g2_o21ai_1 _1513_ (.B1(_0335_),
    .Y(_0336_),
    .A1(\game_inst.vga_inst.row_buffer[11][1] ),
    .A2(net114));
 sg13g2_a21oi_1 _1514_ (.A1(\game_inst.vga_inst.row_buffer[10][1] ),
    .A2(_0246_),
    .Y(_0337_),
    .B1(_0293_));
 sg13g2_a22oi_1 _1515_ (.Y(_0338_),
    .B1(\game_inst.vga_inst.row_buffer[12][1] ),
    .B2(net129),
    .A2(\game_inst.vga_inst.row_buffer[13][1] ),
    .A1(net127));
 sg13g2_nor2_1 _1516_ (.A(net111),
    .B(_0338_),
    .Y(_0339_));
 sg13g2_a221oi_1 _1517_ (.B2(\game_inst.vga_inst.row_buffer[14][1] ),
    .C1(_0339_),
    .B1(net111),
    .A1(\game_inst.vga_inst.row_buffer[15][1] ),
    .Y(_0340_),
    .A2(_0243_));
 sg13g2_a22oi_1 _1518_ (.Y(_0341_),
    .B1(_0340_),
    .B2(_0293_),
    .A2(_0337_),
    .A1(_0336_));
 sg13g2_a21oi_1 _1519_ (.A1(_0284_),
    .A2(_0341_),
    .Y(_0342_),
    .B1(_0300_));
 sg13g2_nand2_1 _1520_ (.Y(_0343_),
    .A(_0274_),
    .B(_0317_));
 sg13g2_nor2b_1 _1521_ (.A(net128),
    .B_N(\game_inst.vga_inst.row_buffer[17][1] ),
    .Y(_0344_));
 sg13g2_a21oi_1 _1522_ (.A1(net128),
    .A2(\game_inst.vga_inst.row_buffer[16][1] ),
    .Y(_0345_),
    .B1(_0344_));
 sg13g2_a221oi_1 _1523_ (.B2(_0300_),
    .C1(_0343_),
    .B1(_0345_),
    .A1(_0333_),
    .Y(_0346_),
    .A2(_0342_));
 sg13g2_o21ai_1 _1524_ (.B1(_0266_),
    .Y(_0347_),
    .A1(_0274_),
    .A2(_0276_));
 sg13g2_o21ai_1 _1525_ (.B1(_0252_),
    .Y(_0348_),
    .A1(_0346_),
    .A2(_0347_));
 sg13g2_o21ai_1 _1526_ (.B1(_0324_),
    .Y(uo_out[2]),
    .A1(_0168_),
    .A2(_0348_));
 sg13g2_nor2b_2 _1527_ (.A(_0278_),
    .B_N(_0343_),
    .Y(uo_out[4]));
 sg13g2_nand2b_1 _1528_ (.Y(_0349_),
    .B(_0275_),
    .A_N(_0274_));
 sg13g2_nand2_1 _1529_ (.Y(_0350_),
    .A(_0343_),
    .B(_0349_));
 sg13g2_a21oi_2 _1530_ (.B1(_0251_),
    .Y(uo_out[0]),
    .A2(_0350_),
    .A1(_0266_));
 sg13g2_nand2_1 _1531_ (.Y(_0351_),
    .A(\game_inst.colorblind ),
    .B(_0323_));
 sg13g2_o21ai_1 _1532_ (.B1(_0351_),
    .Y(uo_out[5]),
    .A1(\game_inst.colorblind ),
    .A2(_0321_));
 sg13g2_o21ai_1 _1533_ (.B1(_0351_),
    .Y(uo_out[1]),
    .A1(\game_inst.colorblind ),
    .A2(_0348_));
 sg13g2_nor2_1 _1534_ (.A(net3),
    .B(net136),
    .Y(_0352_));
 sg13g2_nand2b_1 _1535_ (.Y(_0000_),
    .B(_0352_),
    .A_N(net5));
 sg13g2_and4_1 _1536_ (.A(net1166),
    .B(net1182),
    .C(net1185),
    .D(\game_inst.vga_inst.py[0] ),
    .X(_0353_));
 sg13g2_nand3_1 _1537_ (.B(\game_inst.vga_inst.py[0] ),
    .C(_0240_),
    .A(\game_inst.vga_inst.py[1] ),
    .Y(_0354_));
 sg13g2_nand2_2 _1538_ (.Y(_0355_),
    .A(net1225),
    .B(_0353_));
 sg13g2_and2_1 _1539_ (.A(net122),
    .B(\game_inst.vga_inst.py[4] ),
    .X(_0356_));
 sg13g2_and2_1 _1540_ (.A(_0353_),
    .B(_0356_),
    .X(_0357_));
 sg13g2_xnor2_1 _1541_ (.Y(_0358_),
    .A(\game_inst.vga_inst.py[5] ),
    .B(_0355_));
 sg13g2_xnor2_1 _1542_ (.Y(_0359_),
    .A(\game_inst.apple_inst.i_snake_y[0] ),
    .B(_0358_));
 sg13g2_nor2b_1 _1543_ (.A(\game_inst.vga_inst.px[6] ),
    .B_N(\game_inst.apple_inst.i_snake_x[1] ),
    .Y(_0360_));
 sg13g2_nor3_1 _1544_ (.A(net117),
    .B(_0214_),
    .C(_0360_),
    .Y(_0361_));
 sg13g2_nand2b_1 _1545_ (.Y(_0362_),
    .B(\game_inst.vga_inst.px[6] ),
    .A_N(\game_inst.apple_inst.i_snake_x[1] ));
 sg13g2_nand2b_1 _1546_ (.Y(_0363_),
    .B(\game_inst.vga_inst.px[8] ),
    .A_N(\game_inst.apple_inst.i_snake_x[3] ));
 sg13g2_nand2b_1 _1547_ (.Y(_0364_),
    .B(net126),
    .A_N(\game_inst.apple_inst.i_snake_x[2] ));
 sg13g2_nand3_1 _1548_ (.B(_0363_),
    .C(_0364_),
    .A(_0362_),
    .Y(_0365_));
 sg13g2_nor2b_1 _1549_ (.A(net126),
    .B_N(\game_inst.apple_inst.i_snake_x[2] ),
    .Y(_0366_));
 sg13g2_nor2b_1 _1550_ (.A(net124),
    .B_N(\game_inst.apple_inst.i_snake_x[3] ),
    .Y(_0367_));
 sg13g2_a221oi_1 _1551_ (.B2(_0366_),
    .C1(_0367_),
    .B1(_0363_),
    .A1(\game_inst.apple_inst.i_snake_x[4] ),
    .Y(_0368_),
    .A2(_0216_));
 sg13g2_o21ai_1 _1552_ (.B1(_0368_),
    .Y(_0369_),
    .A1(_0361_),
    .A2(_0365_));
 sg13g2_a21oi_1 _1553_ (.A1(_0207_),
    .A2(\game_inst.vga_inst.px[9] ),
    .Y(_0370_),
    .B1(_0355_));
 sg13g2_a21oi_1 _1554_ (.A1(_0369_),
    .A2(_0370_),
    .Y(_0371_),
    .B1(_0169_));
 sg13g2_nand3_1 _1555_ (.B(_0353_),
    .C(_0356_),
    .A(\game_inst.vga_inst.py[6] ),
    .Y(_0372_));
 sg13g2_a21o_1 _1556_ (.A2(_0356_),
    .A1(_0353_),
    .B1(\game_inst.vga_inst.py[6] ),
    .X(_0373_));
 sg13g2_and3_1 _1557_ (.X(_0374_),
    .A(_0210_),
    .B(_0372_),
    .C(_0373_));
 sg13g2_a21oi_1 _1558_ (.A1(_0372_),
    .A2(_0373_),
    .Y(_0375_),
    .B1(_0210_));
 sg13g2_and2_1 _1559_ (.A(_0186_),
    .B(_0372_),
    .X(_0376_));
 sg13g2_and2_1 _1560_ (.A(_0237_),
    .B(_0357_),
    .X(_0377_));
 sg13g2_a221oi_1 _1561_ (.B2(_0186_),
    .C1(\game_inst.apple_inst.i_snake_y[2] ),
    .B1(_0372_),
    .A1(_0237_),
    .Y(_0378_),
    .A2(_0357_));
 sg13g2_o21ai_1 _1562_ (.B1(\game_inst.apple_inst.i_snake_y[2] ),
    .Y(_0379_),
    .A1(_0376_),
    .A2(_0377_));
 sg13g2_nand2b_2 _1563_ (.Y(_0380_),
    .B(_0357_),
    .A_N(_0238_));
 sg13g2_o21ai_1 _1564_ (.B1(_0380_),
    .Y(_0381_),
    .A1(\game_inst.vga_inst.py[8] ),
    .A2(_0377_));
 sg13g2_xnor2_1 _1565_ (.Y(_0382_),
    .A(\game_inst.apple_inst.i_snake_y[3] ),
    .B(_0381_));
 sg13g2_nor3_1 _1566_ (.A(_0374_),
    .B(_0375_),
    .C(_0378_),
    .Y(_0383_));
 sg13g2_nand4_1 _1567_ (.B(_0371_),
    .C(_0379_),
    .A(_0359_),
    .Y(_0384_),
    .D(_0383_));
 sg13g2_nor2_1 _1568_ (.A(_0382_),
    .B(_0384_),
    .Y(_0385_));
 sg13g2_and3_1 _1569_ (.X(_0386_),
    .A(net1136),
    .B(\game_inst.vga_inst.px[1] ),
    .C(net1141));
 sg13g2_and2_1 _1570_ (.A(net1229),
    .B(_0386_),
    .X(_0387_));
 sg13g2_and2_1 _1571_ (.A(net1289),
    .B(_0387_),
    .X(_0388_));
 sg13g2_nand2_1 _1572_ (.Y(_0389_),
    .A(net1289),
    .B(_0387_));
 sg13g2_nor3_2 _1573_ (.A(_0251_),
    .B(_0355_),
    .C(_0389_),
    .Y(_0390_));
 sg13g2_nor3_2 _1574_ (.A(_0382_),
    .B(_0384_),
    .C(_0390_),
    .Y(_0391_));
 sg13g2_nor3_2 _1575_ (.A(net117),
    .B(\game_inst.apple_inst.i_snake_x[1] ),
    .C(\game_inst.apple_inst.i_snake_x[2] ),
    .Y(_0392_));
 sg13g2_and2_1 _1576_ (.A(_0205_),
    .B(_0392_),
    .X(_0393_));
 sg13g2_xnor2_1 _1577_ (.Y(_0394_),
    .A(_0207_),
    .B(_0393_));
 sg13g2_mux2_1 _1578_ (.A0(_0300_),
    .A1(_0394_),
    .S(net102),
    .X(_0395_));
 sg13g2_xnor2_1 _1579_ (.Y(_0396_),
    .A(\game_inst.apple_inst.i_snake_x[3] ),
    .B(_0392_));
 sg13g2_inv_1 _1580_ (.Y(_0397_),
    .A(_0396_));
 sg13g2_mux2_1 _1581_ (.A0(_0283_),
    .A1(_0396_),
    .S(net102),
    .X(_0398_));
 sg13g2_mux2_1 _1582_ (.A0(_0284_),
    .A1(_0397_),
    .S(net102),
    .X(_0399_));
 sg13g2_o21ai_1 _1583_ (.B1(\game_inst.apple_inst.i_snake_x[2] ),
    .Y(_0400_),
    .A1(net117),
    .A2(\game_inst.apple_inst.i_snake_x[1] ));
 sg13g2_nor2b_2 _1584_ (.A(_0392_),
    .B_N(_0400_),
    .Y(_0401_));
 sg13g2_inv_1 _1585_ (.Y(_0402_),
    .A(_0401_));
 sg13g2_or4_1 _1586_ (.A(_0382_),
    .B(_0384_),
    .C(_0390_),
    .D(_0402_),
    .X(_0403_));
 sg13g2_o21ai_1 _1587_ (.B1(_0403_),
    .Y(_0404_),
    .A1(_0293_),
    .A2(net102));
 sg13g2_mux2_1 _1588_ (.A0(_0293_),
    .A1(_0402_),
    .S(net102),
    .X(_0405_));
 sg13g2_nand3b_1 _1589_ (.B(_0398_),
    .C(_0404_),
    .Y(_0406_),
    .A_N(_0395_));
 sg13g2_nor2_2 _1590_ (.A(_0385_),
    .B(_0390_),
    .Y(_0407_));
 sg13g2_mux2_1 _1591_ (.A0(net128),
    .A1(net117),
    .S(net102),
    .X(_0408_));
 sg13g2_nand2_1 _1592_ (.Y(_0409_),
    .A(_0244_),
    .B(_0247_));
 sg13g2_xor2_1 _1593_ (.B(\game_inst.apple_inst.i_snake_x[1] ),
    .A(net117),
    .X(_0410_));
 sg13g2_inv_1 _1594_ (.Y(_0411_),
    .A(_0410_));
 sg13g2_or4_1 _1595_ (.A(_0382_),
    .B(_0384_),
    .C(_0390_),
    .D(_0411_),
    .X(_0412_));
 sg13g2_o21ai_1 _1596_ (.B1(_0412_),
    .Y(_0413_),
    .A1(net102),
    .A2(_0409_));
 sg13g2_mux2_1 _1597_ (.A0(_0409_),
    .A1(_0411_),
    .S(net102),
    .X(_0414_));
 sg13g2_nand3b_1 _1598_ (.B(_0408_),
    .C(_0413_),
    .Y(_0415_),
    .A_N(_0407_));
 sg13g2_nor2_1 _1599_ (.A(_0406_),
    .B(_0415_),
    .Y(_0416_));
 sg13g2_and2_1 _1600_ (.A(net1137),
    .B(_0391_),
    .X(_0417_));
 sg13g2_mux2_1 _1601_ (.A0(net1236),
    .A1(net99),
    .S(_0416_),
    .X(_0003_));
 sg13g2_nand2b_1 _1602_ (.Y(_0418_),
    .B(net1137),
    .A_N(net1158));
 sg13g2_and2_1 _1603_ (.A(_0391_),
    .B(_0418_),
    .X(_0419_));
 sg13g2_mux2_1 _1604_ (.A0(net1215),
    .A1(net96),
    .S(_0416_),
    .X(_0004_));
 sg13g2_nor3_1 _1605_ (.A(_0395_),
    .B(_0398_),
    .C(_0405_),
    .Y(_0420_));
 sg13g2_nand3b_1 _1606_ (.B(_0399_),
    .C(_0404_),
    .Y(_0421_),
    .A_N(_0395_));
 sg13g2_nand3b_1 _1607_ (.B(_0408_),
    .C(_0414_),
    .Y(_0422_),
    .A_N(_0407_));
 sg13g2_nor2_1 _1608_ (.A(_0421_),
    .B(_0422_),
    .Y(_0423_));
 sg13g2_mux2_1 _1609_ (.A0(net1222),
    .A1(net100),
    .S(_0423_),
    .X(_0005_));
 sg13g2_mux2_1 _1610_ (.A0(net1195),
    .A1(net97),
    .S(_0423_),
    .X(_0006_));
 sg13g2_nor3_2 _1611_ (.A(_0395_),
    .B(_0399_),
    .C(_0404_),
    .Y(_0424_));
 sg13g2_nor3_2 _1612_ (.A(_0407_),
    .B(_0408_),
    .C(_0413_),
    .Y(_0425_));
 sg13g2_nand2_1 _1613_ (.Y(_0426_),
    .A(_0424_),
    .B(_0425_));
 sg13g2_mux2_1 _1614_ (.A0(net100),
    .A1(net1177),
    .S(_0426_),
    .X(_0007_));
 sg13g2_mux2_1 _1615_ (.A0(net97),
    .A1(net1202),
    .S(_0426_),
    .X(_0008_));
 sg13g2_nor2b_1 _1616_ (.A(_0422_),
    .B_N(_0424_),
    .Y(_0427_));
 sg13g2_mux2_1 _1617_ (.A0(net1211),
    .A1(net100),
    .S(_0427_),
    .X(_0009_));
 sg13g2_mux2_1 _1618_ (.A0(net1190),
    .A1(net97),
    .S(_0427_),
    .X(_0010_));
 sg13g2_nor2b_1 _1619_ (.A(net1259),
    .B_N(\game_inst.snake_inst.pos[3] ),
    .Y(_0428_));
 sg13g2_nand4_1 _1620_ (.B(net1180),
    .C(_0232_),
    .A(net1148),
    .Y(_0429_),
    .D(_0428_));
 sg13g2_or3_1 _1621_ (.A(net1257),
    .B(net1246),
    .C(_0192_),
    .X(_0430_));
 sg13g2_nand4_1 _1622_ (.B(net1304),
    .C(net1298),
    .A(_0189_),
    .Y(_0431_),
    .D(net1312));
 sg13g2_nor3_2 _1623_ (.A(_0429_),
    .B(_0430_),
    .C(_0431_),
    .Y(_0432_));
 sg13g2_or3_1 _1624_ (.A(_0429_),
    .B(_0430_),
    .C(_0431_),
    .X(_0433_));
 sg13g2_o21ai_1 _1625_ (.B1(net113),
    .Y(_0011_),
    .A1(net1206),
    .A2(_0432_));
 sg13g2_nand3_1 _1626_ (.B(\game_inst.snake_inst.pos[0] ),
    .C(_0428_),
    .A(_0188_),
    .Y(_0434_));
 sg13g2_or2_1 _1627_ (.X(_0435_),
    .B(_0434_),
    .A(_0431_));
 sg13g2_and2_1 _1628_ (.A(net110),
    .B(_0435_),
    .X(_0436_));
 sg13g2_nand2_2 _1629_ (.Y(_0437_),
    .A(net110),
    .B(_0435_));
 sg13g2_and2_1 _1630_ (.A(net1305),
    .B(net1206),
    .X(_0438_));
 sg13g2_and2_1 _1631_ (.A(net1259),
    .B(_0438_),
    .X(_0439_));
 sg13g2_xnor2_1 _1632_ (.Y(_0440_),
    .A(net1317),
    .B(_0439_));
 sg13g2_o21ai_1 _1633_ (.B1(net112),
    .Y(_0012_),
    .A1(_0437_),
    .A2(_0440_));
 sg13g2_and3_1 _1634_ (.X(_0441_),
    .A(net1317),
    .B(net1168),
    .C(_0439_));
 sg13g2_and2_1 _1635_ (.A(net1304),
    .B(_0441_),
    .X(_0442_));
 sg13g2_o21ai_1 _1636_ (.B1(_0436_),
    .Y(_0443_),
    .A1(net1304),
    .A2(_0441_));
 sg13g2_o21ai_1 _1637_ (.B1(net112),
    .Y(_0013_),
    .A1(_0442_),
    .A2(_0443_));
 sg13g2_nand2_1 _1638_ (.Y(_0444_),
    .A(net1298),
    .B(_0442_));
 sg13g2_nor2_1 _1639_ (.A(net1298),
    .B(_0442_),
    .Y(_0445_));
 sg13g2_nand2_1 _1640_ (.Y(_0446_),
    .A(_0436_),
    .B(_0444_));
 sg13g2_o21ai_1 _1641_ (.B1(net113),
    .Y(_0014_),
    .A1(_0445_),
    .A2(_0446_));
 sg13g2_xor2_1 _1642_ (.B(_0444_),
    .A(net1312),
    .X(_0447_));
 sg13g2_o21ai_1 _1643_ (.B1(net112),
    .Y(_0015_),
    .A1(_0437_),
    .A2(_0447_));
 sg13g2_nor2_1 _1644_ (.A(_0415_),
    .B(_0421_),
    .Y(_0448_));
 sg13g2_mux2_1 _1645_ (.A0(net1203),
    .A1(net100),
    .S(_0448_),
    .X(_0016_));
 sg13g2_mux2_1 _1646_ (.A0(net1194),
    .A1(net97),
    .S(_0448_),
    .X(_0017_));
 sg13g2_nand4_1 _1647_ (.B(net123),
    .C(_0268_),
    .A(\game_inst.vga_inst.px[9] ),
    .Y(_0449_),
    .D(_0388_));
 sg13g2_inv_2 _1648_ (.Y(_0450_),
    .A(_0449_));
 sg13g2_nor2_2 _1649_ (.A(net134),
    .B(_0450_),
    .Y(_0451_));
 sg13g2_nand2_2 _1650_ (.Y(_0452_),
    .A(net137),
    .B(_0449_));
 sg13g2_nor2_1 _1651_ (.A(net1136),
    .B(_0452_),
    .Y(_0018_));
 sg13g2_xnor2_1 _1652_ (.Y(_0453_),
    .A(net1136),
    .B(net1238));
 sg13g2_nor2_1 _1653_ (.A(_0452_),
    .B(_0453_),
    .Y(_0019_));
 sg13g2_a21oi_1 _1654_ (.A1(net1136),
    .A2(\game_inst.vga_inst.px[1] ),
    .Y(_0454_),
    .B1(net1141));
 sg13g2_nor3_1 _1655_ (.A(net134),
    .B(_0386_),
    .C(net1142),
    .Y(_0020_));
 sg13g2_o21ai_1 _1656_ (.B1(net137),
    .Y(_0455_),
    .A1(net1229),
    .A2(_0386_));
 sg13g2_nor2_1 _1657_ (.A(_0387_),
    .B(net1230),
    .Y(_0021_));
 sg13g2_o21ai_1 _1658_ (.B1(net137),
    .Y(_0456_),
    .A1(net1289),
    .A2(_0387_));
 sg13g2_nor2_1 _1659_ (.A(_0388_),
    .B(_0456_),
    .Y(_0022_));
 sg13g2_o21ai_1 _1660_ (.B1(_0451_),
    .Y(_0457_),
    .A1(net129),
    .A2(_0388_));
 sg13g2_a21oi_1 _1661_ (.A1(net129),
    .A2(_0388_),
    .Y(_0023_),
    .B1(_0457_));
 sg13g2_a21oi_1 _1662_ (.A1(net129),
    .A2(_0388_),
    .Y(_0458_),
    .B1(net127));
 sg13g2_nor2_1 _1663_ (.A(_0247_),
    .B(_0389_),
    .Y(_0459_));
 sg13g2_nor3_1 _1664_ (.A(_0452_),
    .B(_0458_),
    .C(_0459_),
    .Y(_0024_));
 sg13g2_nor2_1 _1665_ (.A(net125),
    .B(_0459_),
    .Y(_0460_));
 sg13g2_and2_1 _1666_ (.A(net125),
    .B(_0459_),
    .X(_0461_));
 sg13g2_nor3_1 _1667_ (.A(_0452_),
    .B(_0460_),
    .C(_0461_),
    .Y(_0025_));
 sg13g2_nand2_1 _1668_ (.Y(_0462_),
    .A(net123),
    .B(_0461_));
 sg13g2_o21ai_1 _1669_ (.B1(_0451_),
    .Y(_0463_),
    .A1(net123),
    .A2(_0461_));
 sg13g2_nor2b_1 _1670_ (.A(_0463_),
    .B_N(_0462_),
    .Y(_0026_));
 sg13g2_xnor2_1 _1671_ (.Y(_0464_),
    .A(_0216_),
    .B(_0462_));
 sg13g2_nor2_1 _1672_ (.A(_0452_),
    .B(_0464_),
    .Y(_0027_));
 sg13g2_nor2b_2 _1673_ (.A(_0415_),
    .B_N(_0424_),
    .Y(_0465_));
 sg13g2_mux2_1 _1674_ (.A0(net1243),
    .A1(net101),
    .S(_0465_),
    .X(_0028_));
 sg13g2_mux2_1 _1675_ (.A0(net1235),
    .A1(net98),
    .S(_0465_),
    .X(_0029_));
 sg13g2_nand3_1 _1676_ (.B(_0398_),
    .C(_0404_),
    .A(_0395_),
    .Y(_0466_));
 sg13g2_nor3_2 _1677_ (.A(_0407_),
    .B(_0408_),
    .C(_0414_),
    .Y(_0467_));
 sg13g2_nand2b_1 _1678_ (.Y(_0468_),
    .B(_0467_),
    .A_N(_0466_));
 sg13g2_mux2_1 _1679_ (.A0(net100),
    .A1(net1189),
    .S(_0468_),
    .X(_0030_));
 sg13g2_mux2_1 _1680_ (.A0(net97),
    .A1(net1173),
    .S(_0468_),
    .X(_0031_));
 sg13g2_nand2_1 _1681_ (.Y(_0469_),
    .A(_0424_),
    .B(_0467_));
 sg13g2_mux2_1 _1682_ (.A0(net100),
    .A1(net1219),
    .S(_0469_),
    .X(_0032_));
 sg13g2_mux2_1 _1683_ (.A0(net97),
    .A1(net1208),
    .S(_0469_),
    .X(_0033_));
 sg13g2_nor3_1 _1684_ (.A(_0395_),
    .B(_0398_),
    .C(_0404_),
    .Y(_0470_));
 sg13g2_nand3b_1 _1685_ (.B(_0399_),
    .C(_0405_),
    .Y(_0471_),
    .A_N(_0395_));
 sg13g2_nand2_1 _1686_ (.Y(_0472_),
    .A(_0467_),
    .B(_0470_));
 sg13g2_mux2_1 _1687_ (.A0(net99),
    .A1(net1210),
    .S(_0472_),
    .X(_0034_));
 sg13g2_mux2_1 _1688_ (.A0(net96),
    .A1(net1212),
    .S(_0472_),
    .X(_0035_));
 sg13g2_nand2_1 _1689_ (.Y(_0473_),
    .A(_0420_),
    .B(_0467_));
 sg13g2_mux2_1 _1690_ (.A0(net100),
    .A1(net1209),
    .S(_0473_),
    .X(_0036_));
 sg13g2_mux2_1 _1691_ (.A0(net97),
    .A1(net1184),
    .S(_0473_),
    .X(_0037_));
 sg13g2_nand2_1 _1692_ (.Y(_0474_),
    .A(net1152),
    .B(net110));
 sg13g2_nand2_1 _1693_ (.Y(_0475_),
    .A(\game_inst.control_inst.dir[0] ),
    .B(_0432_));
 sg13g2_a21oi_1 _1694_ (.A1(_0474_),
    .A2(_0475_),
    .Y(_0038_),
    .B1(net132));
 sg13g2_nor2_2 _1695_ (.A(_0178_),
    .B(net109),
    .Y(_0476_));
 sg13g2_a21oi_1 _1696_ (.A1(net1160),
    .A2(net109),
    .Y(_0477_),
    .B1(_0476_));
 sg13g2_nor2_1 _1697_ (.A(net133),
    .B(net1161),
    .Y(_0039_));
 sg13g2_nand2_1 _1698_ (.Y(_0478_),
    .A(_0425_),
    .B(_0470_));
 sg13g2_mux2_1 _1699_ (.A0(net99),
    .A1(net1224),
    .S(_0478_),
    .X(_0040_));
 sg13g2_mux2_1 _1700_ (.A0(net96),
    .A1(net1204),
    .S(_0478_),
    .X(_0041_));
 sg13g2_nand2_1 _1701_ (.Y(_0042_),
    .A(net1137),
    .B(_0235_));
 sg13g2_nand2b_1 _1702_ (.Y(_0479_),
    .B(net1158),
    .A_N(net1137));
 sg13g2_a21oi_1 _1703_ (.A1(_0418_),
    .A2(_0479_),
    .Y(_0043_),
    .B1(_0234_));
 sg13g2_nor3_1 _1704_ (.A(\game_inst.vga_inst.py[4] ),
    .B(\game_inst.vga_inst.py[1] ),
    .C(\game_inst.vga_inst.py[0] ),
    .Y(_0480_));
 sg13g2_and4_1 _1705_ (.A(\game_inst.vga_inst.py[9] ),
    .B(_0187_),
    .C(_0240_),
    .D(_0480_),
    .X(_0481_));
 sg13g2_a21oi_1 _1706_ (.A1(_0272_),
    .A2(_0481_),
    .Y(_0482_),
    .B1(_0449_));
 sg13g2_and2_1 _1707_ (.A(net1306),
    .B(_0450_),
    .X(_0483_));
 sg13g2_o21ai_1 _1708_ (.B1(net137),
    .Y(_0484_),
    .A1(net1306),
    .A2(_0482_));
 sg13g2_nor2_1 _1709_ (.A(_0483_),
    .B(_0484_),
    .Y(_0044_));
 sg13g2_o21ai_1 _1710_ (.B1(net137),
    .Y(_0485_),
    .A1(net1185),
    .A2(_0483_));
 sg13g2_a21oi_1 _1711_ (.A1(net1185),
    .A2(_0483_),
    .Y(_0045_),
    .B1(_0485_));
 sg13g2_nand2_1 _1712_ (.Y(_0486_),
    .A(net1182),
    .B(_0451_));
 sg13g2_a21oi_1 _1713_ (.A1(\game_inst.vga_inst.py[1] ),
    .A2(\game_inst.vga_inst.py[0] ),
    .Y(_0487_),
    .B1(net1182));
 sg13g2_and3_1 _1714_ (.X(_0488_),
    .A(net1182),
    .B(\game_inst.vga_inst.py[1] ),
    .C(\game_inst.vga_inst.py[0] ));
 sg13g2_or2_1 _1715_ (.X(_0489_),
    .B(_0488_),
    .A(_0487_));
 sg13g2_nand2_1 _1716_ (.Y(_0490_),
    .A(net137),
    .B(_0482_));
 sg13g2_o21ai_1 _1717_ (.B1(_0486_),
    .Y(_0046_),
    .A1(_0489_),
    .A2(_0490_));
 sg13g2_nand2_1 _1718_ (.Y(_0491_),
    .A(net1166),
    .B(_0451_));
 sg13g2_o21ai_1 _1719_ (.B1(_0354_),
    .Y(_0492_),
    .A1(net1166),
    .A2(_0488_));
 sg13g2_o21ai_1 _1720_ (.B1(_0491_),
    .Y(_0047_),
    .A1(_0490_),
    .A2(_0492_));
 sg13g2_a21oi_1 _1721_ (.A1(_0353_),
    .A2(_0450_),
    .Y(_0493_),
    .B1(net1225));
 sg13g2_nor2_2 _1722_ (.A(_0355_),
    .B(_0449_),
    .Y(_0494_));
 sg13g2_nor3_1 _1723_ (.A(net134),
    .B(net1226),
    .C(_0494_),
    .Y(_0048_));
 sg13g2_o21ai_1 _1724_ (.B1(net137),
    .Y(_0495_),
    .A1(net122),
    .A2(_0494_));
 sg13g2_a21oi_1 _1725_ (.A1(net122),
    .A2(_0494_),
    .Y(_0049_),
    .B1(_0495_));
 sg13g2_a21oi_1 _1726_ (.A1(net122),
    .A2(_0494_),
    .Y(_0496_),
    .B1(net1287));
 sg13g2_nor2_2 _1727_ (.A(_0372_),
    .B(_0449_),
    .Y(_0497_));
 sg13g2_nor3_1 _1728_ (.A(net134),
    .B(net1288),
    .C(_0497_),
    .Y(_0050_));
 sg13g2_o21ai_1 _1729_ (.B1(net137),
    .Y(_0498_),
    .A1(net1241),
    .A2(_0497_));
 sg13g2_a21oi_1 _1730_ (.A1(net1241),
    .A2(_0497_),
    .Y(_0051_),
    .B1(_0498_));
 sg13g2_a21oi_1 _1731_ (.A1(net1241),
    .A2(_0497_),
    .Y(_0499_),
    .B1(net1271));
 sg13g2_o21ai_1 _1732_ (.B1(net138),
    .Y(_0500_),
    .A1(_0380_),
    .A2(_0449_));
 sg13g2_nor2_1 _1733_ (.A(_0499_),
    .B(_0500_),
    .Y(_0052_));
 sg13g2_nand2_1 _1734_ (.Y(_0501_),
    .A(net1217),
    .B(_0451_));
 sg13g2_xor2_1 _1735_ (.B(_0380_),
    .A(net1217),
    .X(_0502_));
 sg13g2_o21ai_1 _1736_ (.B1(_0501_),
    .Y(_0053_),
    .A1(_0490_),
    .A2(_0502_));
 sg13g2_nand4_1 _1737_ (.B(\game_inst.snake_inst.length[5] ),
    .C(\game_inst.snake_inst.length[6] ),
    .A(_0197_),
    .Y(_0503_),
    .D(net1146));
 sg13g2_nand2_1 _1738_ (.Y(_0504_),
    .A(\game_inst.snake_inst.length[0] ),
    .B(net1174));
 sg13g2_nor4_1 _1739_ (.A(net1198),
    .B(\game_inst.snake_inst.length[2] ),
    .C(_0503_),
    .D(_0504_),
    .Y(_0505_));
 sg13g2_nor2_1 _1740_ (.A(net1246),
    .B(_0505_),
    .Y(_0506_));
 sg13g2_nor2_1 _1741_ (.A(net131),
    .B(net1247),
    .Y(_0054_));
 sg13g2_a21oi_1 _1742_ (.A1(\game_inst.apple_inst.o_ready ),
    .A2(_0234_),
    .Y(_0507_),
    .B1(\game_inst.apple_inst.i_snake_valid ));
 sg13g2_nor3_1 _1743_ (.A(_0228_),
    .B(_0230_),
    .C(_0507_),
    .Y(_0508_));
 sg13g2_and3_1 _1744_ (.X(_0509_),
    .A(\game_inst.apple_inst.apple_y[1] ),
    .B(\game_inst.apple_inst.apple_y[2] ),
    .C(\game_inst.apple_inst.apple_y[3] ));
 sg13g2_nand2_1 _1745_ (.Y(_0510_),
    .A(\game_inst.apple_inst.apple_x[0] ),
    .B(\game_inst.apple_inst.apple_x[1] ));
 sg13g2_nor2_1 _1746_ (.A(\game_inst.apple_inst.apple_x[2] ),
    .B(\game_inst.apple_inst.apple_x[3] ),
    .Y(_0511_));
 sg13g2_a21oi_1 _1747_ (.A1(_0510_),
    .A2(_0511_),
    .Y(_0512_),
    .B1(_0206_));
 sg13g2_or4_1 _1748_ (.A(net130),
    .B(_0508_),
    .C(_0509_),
    .D(_0512_),
    .X(_0513_));
 sg13g2_nor2_1 _1749_ (.A(\game_inst.apple_inst.apple_x[0] ),
    .B(net103),
    .Y(_0514_));
 sg13g2_a21oi_1 _1750_ (.A1(_0184_),
    .A2(net103),
    .Y(_0055_),
    .B1(_0514_));
 sg13g2_nor2_1 _1751_ (.A(\game_inst.apple_inst.apple_x[1] ),
    .B(net103),
    .Y(_0515_));
 sg13g2_a21oi_1 _1752_ (.A1(_0183_),
    .A2(net103),
    .Y(_0056_),
    .B1(_0515_));
 sg13g2_nand2_1 _1753_ (.Y(_0516_),
    .A(net1178),
    .B(net105));
 sg13g2_o21ai_1 _1754_ (.B1(_0516_),
    .Y(_0057_),
    .A1(_0202_),
    .A2(net104));
 sg13g2_nor2_1 _1755_ (.A(\game_inst.apple_inst.apple_x[3] ),
    .B(net103),
    .Y(_0517_));
 sg13g2_a21oi_1 _1756_ (.A1(_0182_),
    .A2(net103),
    .Y(_0058_),
    .B1(_0517_));
 sg13g2_nor2_1 _1757_ (.A(net1234),
    .B(net103),
    .Y(_0518_));
 sg13g2_a21oi_1 _1758_ (.A1(_0181_),
    .A2(net103),
    .Y(_0059_),
    .B1(_0518_));
 sg13g2_nor2_1 _1759_ (.A(net1263),
    .B(_0185_),
    .Y(_0519_));
 sg13g2_a21oi_1 _1760_ (.A1(_0235_),
    .A2(_0519_),
    .Y(_0520_),
    .B1(net1180));
 sg13g2_nor2_1 _1761_ (.A(net105),
    .B(net1264),
    .Y(_0060_));
 sg13g2_a21oi_1 _1762_ (.A1(_0185_),
    .A2(_0235_),
    .Y(_0061_),
    .B1(net104));
 sg13g2_nor2_1 _1763_ (.A(net1156),
    .B(net1171),
    .Y(_0521_));
 sg13g2_o21ai_1 _1764_ (.B1(net136),
    .Y(_0522_),
    .A1(net1248),
    .A2(_0521_));
 sg13g2_nand2b_1 _1765_ (.Y(_0523_),
    .B(net4),
    .A_N(net1248));
 sg13g2_nand3_1 _1766_ (.B(_0522_),
    .C(_0523_),
    .A(net118),
    .Y(_0524_));
 sg13g2_nand2b_1 _1767_ (.Y(_0525_),
    .B(net5),
    .A_N(net1248));
 sg13g2_nand2_1 _1768_ (.Y(_0526_),
    .A(net1248),
    .B(net3));
 sg13g2_nand3b_1 _1769_ (.B(_0525_),
    .C(_0526_),
    .Y(_0527_),
    .A_N(net118));
 sg13g2_nand3_1 _1770_ (.B(_0523_),
    .C(_0527_),
    .A(_0522_),
    .Y(_0528_));
 sg13g2_nand2b_1 _1771_ (.Y(_0529_),
    .B(_0528_),
    .A_N(net118));
 sg13g2_nand3_1 _1772_ (.B(_0523_),
    .C(_0525_),
    .A(_0178_),
    .Y(_0530_));
 sg13g2_nand3_1 _1773_ (.B(_0526_),
    .C(_0530_),
    .A(_0522_),
    .Y(_0531_));
 sg13g2_xnor2_1 _1774_ (.Y(_0532_),
    .A(\game_inst.control_inst.dir[1] ),
    .B(_0531_));
 sg13g2_a21oi_1 _1775_ (.A1(_0524_),
    .A2(_0529_),
    .Y(_0533_),
    .B1(_0532_));
 sg13g2_nor2_1 _1776_ (.A(net1180),
    .B(_0533_),
    .Y(_0534_));
 sg13g2_a21oi_1 _1777_ (.A1(\game_inst.apple_inst.o_ready ),
    .A2(_0533_),
    .Y(_0535_),
    .B1(net105));
 sg13g2_nor2b_2 _1778_ (.A(_0534_),
    .B_N(_0535_),
    .Y(_0536_));
 sg13g2_xnor2_1 _1779_ (.Y(_0537_),
    .A(net1223),
    .B(net1178));
 sg13g2_a21oi_1 _1780_ (.A1(net1192),
    .A2(net95),
    .Y(_0538_),
    .B1(net134));
 sg13g2_o21ai_1 _1781_ (.B1(_0538_),
    .Y(_0062_),
    .A1(net94),
    .A2(_0537_));
 sg13g2_a21oi_1 _1782_ (.A1(net1162),
    .A2(net94),
    .Y(_0539_),
    .B1(net134));
 sg13g2_o21ai_1 _1783_ (.B1(_0539_),
    .Y(_0063_),
    .A1(_0184_),
    .A2(net94));
 sg13g2_a21oi_1 _1784_ (.A1(net1178),
    .A2(net94),
    .Y(_0540_),
    .B1(net134));
 sg13g2_o21ai_1 _1785_ (.B1(_0540_),
    .Y(_0064_),
    .A1(_0183_),
    .A2(net94));
 sg13g2_o21ai_1 _1786_ (.B1(net138),
    .Y(_0541_),
    .A1(net1178),
    .A2(net95));
 sg13g2_a21oi_1 _1787_ (.A1(_0182_),
    .A2(net94),
    .Y(_0065_),
    .B1(_0541_));
 sg13g2_o21ai_1 _1788_ (.B1(net138),
    .Y(_0542_),
    .A1(net1164),
    .A2(net94));
 sg13g2_a21oi_1 _1789_ (.A1(_0181_),
    .A2(net94),
    .Y(_0066_),
    .B1(_0542_));
 sg13g2_nand2b_1 _1790_ (.Y(_0543_),
    .B(\game_inst.apple_inst.random_inst.lfsr4[3] ),
    .A_N(net95));
 sg13g2_a21oi_1 _1791_ (.A1(net1154),
    .A2(_0543_),
    .Y(_0544_),
    .B1(net135));
 sg13g2_o21ai_1 _1792_ (.B1(_0544_),
    .Y(_0067_),
    .A1(net1154),
    .A2(_0543_));
 sg13g2_a21oi_1 _1793_ (.A1(net1227),
    .A2(net95),
    .Y(_0545_),
    .B1(net134));
 sg13g2_o21ai_1 _1794_ (.B1(_0545_),
    .Y(_0068_),
    .A1(_0180_),
    .A2(net1181));
 sg13g2_o21ai_1 _1795_ (.B1(net139),
    .Y(_0546_),
    .A1(net1227),
    .A2(net95));
 sg13g2_a21oi_1 _1796_ (.A1(_0179_),
    .A2(net95),
    .Y(_0069_),
    .B1(_0546_));
 sg13g2_a21oi_1 _1797_ (.A1(net1233),
    .A2(net95),
    .Y(_0547_),
    .B1(net135));
 sg13g2_o21ai_1 _1798_ (.B1(_0547_),
    .Y(_0070_),
    .A1(_0179_),
    .A2(net1181));
 sg13g2_nor2_1 _1799_ (.A(_0406_),
    .B(_0422_),
    .Y(_0548_));
 sg13g2_mux2_1 _1800_ (.A0(net1221),
    .A1(net99),
    .S(_0548_),
    .X(_0071_));
 sg13g2_mux2_1 _1801_ (.A0(net1239),
    .A1(net96),
    .S(_0548_),
    .X(_0072_));
 sg13g2_nand2b_2 _1802_ (.Y(_0549_),
    .B(_0425_),
    .A_N(_0406_));
 sg13g2_mux2_1 _1803_ (.A0(net99),
    .A1(net1244),
    .S(_0549_),
    .X(_0073_));
 sg13g2_mux2_1 _1804_ (.A0(net96),
    .A1(net1237),
    .S(_0549_),
    .X(_0074_));
 sg13g2_nor2_1 _1805_ (.A(_0422_),
    .B(_0471_),
    .Y(_0550_));
 sg13g2_mux2_1 _1806_ (.A0(net1232),
    .A1(net99),
    .S(_0550_),
    .X(_0075_));
 sg13g2_mux2_1 _1807_ (.A0(net1228),
    .A1(net96),
    .S(_0550_),
    .X(_0076_));
 sg13g2_nor2_1 _1808_ (.A(_0415_),
    .B(_0471_),
    .Y(_0551_));
 sg13g2_mux2_1 _1809_ (.A0(net1201),
    .A1(net99),
    .S(_0551_),
    .X(_0077_));
 sg13g2_mux2_1 _1810_ (.A0(net1191),
    .A1(net96),
    .S(_0551_),
    .X(_0078_));
 sg13g2_nand2_1 _1811_ (.Y(_0552_),
    .A(net1156),
    .B(net110));
 sg13g2_a21oi_1 _1812_ (.A1(_0475_),
    .A2(_0552_),
    .Y(_0079_),
    .B1(net132));
 sg13g2_nor2_1 _1813_ (.A(net1248),
    .B(_0432_),
    .Y(_0553_));
 sg13g2_nor2_2 _1814_ (.A(net1336),
    .B(net110),
    .Y(_0554_));
 sg13g2_nor3_1 _1815_ (.A(net131),
    .B(net1249),
    .C(_0554_),
    .Y(_0080_));
 sg13g2_nand2_1 _1816_ (.Y(_0555_),
    .A(net1320),
    .B(net108));
 sg13g2_xnor2_1 _1817_ (.Y(_0556_),
    .A(net1320),
    .B(net1325));
 sg13g2_nor2_1 _1818_ (.A(net108),
    .B(_0556_),
    .Y(_0557_));
 sg13g2_nand3b_1 _1819_ (.B(net113),
    .C(_0555_),
    .Y(_0081_),
    .A_N(_0557_));
 sg13g2_nand2_1 _1820_ (.Y(_0558_),
    .A(net1291),
    .B(net108));
 sg13g2_and2_1 _1821_ (.A(\game_inst.control_inst.dir[1] ),
    .B(net118),
    .X(_0559_));
 sg13g2_nand2_1 _1822_ (.Y(_0560_),
    .A(\game_inst.head_x[1] ),
    .B(_0559_));
 sg13g2_xnor2_1 _1823_ (.Y(_0561_),
    .A(_0176_),
    .B(_0559_));
 sg13g2_nand2_1 _1824_ (.Y(_0562_),
    .A(\game_inst.head_x[0] ),
    .B(_0561_));
 sg13g2_xnor2_1 _1825_ (.Y(_0563_),
    .A(_0177_),
    .B(_0561_));
 sg13g2_a22oi_1 _1826_ (.Y(_0564_),
    .B1(_0563_),
    .B2(_0476_),
    .A2(_0554_),
    .A1(net1291));
 sg13g2_a21oi_1 _1827_ (.A1(_0558_),
    .A2(_0564_),
    .Y(_0082_),
    .B1(net130));
 sg13g2_nand2_1 _1828_ (.Y(_0565_),
    .A(net1297),
    .B(net108));
 sg13g2_xnor2_1 _1829_ (.Y(_0566_),
    .A(\game_inst.head_x[2] ),
    .B(_0559_));
 sg13g2_nand3_1 _1830_ (.B(_0562_),
    .C(_0566_),
    .A(_0560_),
    .Y(_0567_));
 sg13g2_a21oi_1 _1831_ (.A1(_0560_),
    .A2(_0562_),
    .Y(_0568_),
    .B1(_0566_));
 sg13g2_nor2b_1 _1832_ (.A(_0568_),
    .B_N(_0476_),
    .Y(_0569_));
 sg13g2_a22oi_1 _1833_ (.Y(_0570_),
    .B1(_0567_),
    .B2(_0569_),
    .A2(_0554_),
    .A1(net1297));
 sg13g2_a21oi_1 _1834_ (.A1(_0565_),
    .A2(_0570_),
    .Y(_0083_),
    .B1(net130));
 sg13g2_a21oi_1 _1835_ (.A1(net121),
    .A2(net108),
    .Y(_0571_),
    .B1(net130));
 sg13g2_a21oi_1 _1836_ (.A1(\game_inst.head_x[2] ),
    .A2(_0559_),
    .Y(_0572_),
    .B1(_0568_));
 sg13g2_nor2b_1 _1837_ (.A(_0572_),
    .B_N(net121),
    .Y(_0573_));
 sg13g2_nor2b_1 _1838_ (.A(net121),
    .B_N(_0572_),
    .Y(_0574_));
 sg13g2_nor2_1 _1839_ (.A(_0573_),
    .B(_0574_),
    .Y(_0575_));
 sg13g2_xor2_1 _1840_ (.B(_0575_),
    .A(net118),
    .X(_0576_));
 sg13g2_a22oi_1 _1841_ (.Y(_0577_),
    .B1(_0576_),
    .B2(_0476_),
    .A2(_0554_),
    .A1(net121));
 sg13g2_nand2_1 _1842_ (.Y(_0084_),
    .A(_0571_),
    .B(_0577_));
 sg13g2_nand2_1 _1843_ (.Y(_0578_),
    .A(net1284),
    .B(net108));
 sg13g2_nor2_1 _1844_ (.A(_0178_),
    .B(net118),
    .Y(_0579_));
 sg13g2_a22oi_1 _1845_ (.Y(_0580_),
    .B1(_0579_),
    .B2(_0573_),
    .A2(_0574_),
    .A1(_0559_));
 sg13g2_a21oi_1 _1846_ (.A1(_0174_),
    .A2(_0580_),
    .Y(_0581_),
    .B1(net108));
 sg13g2_o21ai_1 _1847_ (.B1(_0581_),
    .Y(_0582_),
    .A1(_0174_),
    .A2(_0580_));
 sg13g2_a21oi_1 _1848_ (.A1(_0578_),
    .A2(_0582_),
    .Y(_0085_),
    .B1(net130));
 sg13g2_nand2_1 _1849_ (.Y(_0583_),
    .A(net1314),
    .B(net109));
 sg13g2_xnor2_1 _1850_ (.Y(_0584_),
    .A(net1314),
    .B(net1325));
 sg13g2_nand2_1 _1851_ (.Y(_0585_),
    .A(_0432_),
    .B(_0584_));
 sg13g2_a21oi_1 _1852_ (.A1(_0583_),
    .A2(_0585_),
    .Y(_0086_),
    .B1(net130));
 sg13g2_nand2_1 _1853_ (.Y(_0586_),
    .A(net1292),
    .B(net109));
 sg13g2_nor2b_2 _1854_ (.A(\game_inst.control_inst.dir[1] ),
    .B_N(\game_inst.control_inst.dir[0] ),
    .Y(_0587_));
 sg13g2_or2_1 _1855_ (.X(_0588_),
    .B(_0587_),
    .A(net120));
 sg13g2_and2_1 _1856_ (.A(net120),
    .B(_0587_),
    .X(_0589_));
 sg13g2_xnor2_1 _1857_ (.Y(_0590_),
    .A(net120),
    .B(_0587_));
 sg13g2_xnor2_1 _1858_ (.Y(_0591_),
    .A(\game_inst.head_y[0] ),
    .B(_0590_));
 sg13g2_a22oi_1 _1859_ (.Y(_0592_),
    .B1(_0554_),
    .B2(_0591_),
    .A2(_0476_),
    .A1(net1292));
 sg13g2_nand3_1 _1860_ (.B(_0586_),
    .C(_0592_),
    .A(net113),
    .Y(_0087_));
 sg13g2_nand2_1 _1861_ (.Y(_0593_),
    .A(net119),
    .B(net109));
 sg13g2_nand2_1 _1862_ (.Y(_0594_),
    .A(net113),
    .B(_0593_));
 sg13g2_a21oi_1 _1863_ (.A1(\game_inst.head_y[0] ),
    .A2(_0588_),
    .Y(_0595_),
    .B1(_0589_));
 sg13g2_nor2b_1 _1864_ (.A(net119),
    .B_N(net118),
    .Y(_0596_));
 sg13g2_xnor2_1 _1865_ (.Y(_0597_),
    .A(net119),
    .B(_0587_));
 sg13g2_nand2_1 _1866_ (.Y(_0598_),
    .A(_0595_),
    .B(_0597_));
 sg13g2_nor2_1 _1867_ (.A(_0595_),
    .B(_0597_),
    .Y(_0599_));
 sg13g2_nand2_1 _1868_ (.Y(_0600_),
    .A(_0554_),
    .B(_0598_));
 sg13g2_nand2_1 _1869_ (.Y(_0601_),
    .A(net119),
    .B(_0476_));
 sg13g2_o21ai_1 _1870_ (.B1(_0601_),
    .Y(_0602_),
    .A1(_0599_),
    .A2(_0600_));
 sg13g2_or2_1 _1871_ (.X(_0088_),
    .B(_0602_),
    .A(_0594_));
 sg13g2_or2_1 _1872_ (.X(_0603_),
    .B(_0599_),
    .A(_0596_));
 sg13g2_nand2_1 _1873_ (.Y(_0604_),
    .A(net118),
    .B(_0599_));
 sg13g2_nand3_1 _1874_ (.B(_0603_),
    .C(_0604_),
    .A(_0178_),
    .Y(_0605_));
 sg13g2_o21ai_1 _1875_ (.B1(_0432_),
    .Y(_0606_),
    .A1(_0170_),
    .A2(_0605_));
 sg13g2_a21oi_1 _1876_ (.A1(_0170_),
    .A2(_0605_),
    .Y(_0607_),
    .B1(_0606_));
 sg13g2_a21oi_1 _1877_ (.A1(net1283),
    .A2(net109),
    .Y(_0608_),
    .B1(_0607_));
 sg13g2_nor2_1 _1878_ (.A(net130),
    .B(_0608_),
    .Y(_0089_));
 sg13g2_nand2_1 _1879_ (.Y(_0090_),
    .A(net113),
    .B(_0528_));
 sg13g2_nor2_1 _1880_ (.A(net131),
    .B(_0531_),
    .Y(_0091_));
 sg13g2_nor2_2 _1881_ (.A(net1139),
    .B(net106),
    .Y(_0609_));
 sg13g2_a22oi_1 _1882_ (.Y(_0610_),
    .B1(net106),
    .B2(_0555_),
    .A2(net107),
    .A1(net1326));
 sg13g2_nor2_1 _1883_ (.A(_0557_),
    .B(_0610_),
    .Y(_0611_));
 sg13g2_xnor2_1 _1884_ (.Y(_0092_),
    .A(_0609_),
    .B(_0611_));
 sg13g2_nor2_1 _1885_ (.A(net107),
    .B(_0558_),
    .Y(_0612_));
 sg13g2_nand2_2 _1886_ (.Y(_0613_),
    .A(\game_inst.snake_inst.dir_first[1] ),
    .B(\game_inst.snake_inst.dir_first[0] ));
 sg13g2_nor2_1 _1887_ (.A(_0410_),
    .B(_0613_),
    .Y(_0614_));
 sg13g2_xnor2_1 _1888_ (.Y(_0615_),
    .A(_0410_),
    .B(_0613_));
 sg13g2_a21oi_1 _1889_ (.A1(net1139),
    .A2(_0615_),
    .Y(_0616_),
    .B1(net106));
 sg13g2_nor2_1 _1890_ (.A(_0612_),
    .B(_0616_),
    .Y(_0617_));
 sg13g2_a22oi_1 _1891_ (.Y(_0093_),
    .B1(_0617_),
    .B2(_0564_),
    .A2(_0609_),
    .A1(_0201_));
 sg13g2_xor2_1 _1892_ (.B(_0614_),
    .A(_0401_),
    .X(_0618_));
 sg13g2_a22oi_1 _1893_ (.Y(_0619_),
    .B1(_0618_),
    .B2(net107),
    .A2(_0565_),
    .A1(net106));
 sg13g2_nor2_1 _1894_ (.A(_0609_),
    .B(_0619_),
    .Y(_0620_));
 sg13g2_a22oi_1 _1895_ (.Y(_0094_),
    .B1(_0620_),
    .B2(_0570_),
    .A2(_0609_),
    .A1(_0203_));
 sg13g2_a21o_1 _1896_ (.A2(net108),
    .A1(net121),
    .B1(_0436_),
    .X(_0621_));
 sg13g2_nand2_1 _1897_ (.Y(_0622_),
    .A(_0397_),
    .B(_0613_));
 sg13g2_nor3_1 _1898_ (.A(_0200_),
    .B(_0201_),
    .C(_0203_),
    .Y(_0623_));
 sg13g2_a21oi_1 _1899_ (.A1(\game_inst.apple_inst.i_snake_x[3] ),
    .A2(_0623_),
    .Y(_0624_),
    .B1(_0613_));
 sg13g2_o21ai_1 _1900_ (.B1(_0624_),
    .Y(_0625_),
    .A1(\game_inst.apple_inst.i_snake_x[3] ),
    .A2(_0623_));
 sg13g2_nand3_1 _1901_ (.B(_0622_),
    .C(_0625_),
    .A(net107),
    .Y(_0626_));
 sg13g2_o21ai_1 _1902_ (.B1(_0621_),
    .Y(_0627_),
    .A1(_0609_),
    .A2(_0626_));
 sg13g2_a22oi_1 _1903_ (.Y(_0095_),
    .B1(_0627_),
    .B2(_0577_),
    .A2(_0609_),
    .A1(_0205_));
 sg13g2_nor2b_1 _1904_ (.A(_0393_),
    .B_N(_0613_),
    .Y(_0628_));
 sg13g2_nor2_1 _1905_ (.A(_0624_),
    .B(_0628_),
    .Y(_0629_));
 sg13g2_xnor2_1 _1906_ (.Y(_0630_),
    .A(net1313),
    .B(_0629_));
 sg13g2_a22oi_1 _1907_ (.Y(_0631_),
    .B1(_0630_),
    .B2(net107),
    .A2(_0578_),
    .A1(net106));
 sg13g2_nor2_1 _1908_ (.A(_0609_),
    .B(_0631_),
    .Y(_0632_));
 sg13g2_a22oi_1 _1909_ (.Y(_0096_),
    .B1(_0632_),
    .B2(_0582_),
    .A2(_0609_),
    .A1(_0207_));
 sg13g2_a22oi_1 _1910_ (.Y(_0633_),
    .B1(net1265),
    .B2(_0190_),
    .A2(_0196_),
    .A1(\game_inst.snake_inst.pos[3] ));
 sg13g2_xnor2_1 _1911_ (.Y(_0634_),
    .A(net1259),
    .B(net1274));
 sg13g2_a22oi_1 _1912_ (.Y(_0635_),
    .B1(net1198),
    .B2(_0188_),
    .A2(_0194_),
    .A1(\game_inst.snake_inst.pos[0] ));
 sg13g2_xnor2_1 _1913_ (.Y(_0636_),
    .A(\game_inst.snake_inst.pos[5] ),
    .B(net1277));
 sg13g2_nand4_1 _1914_ (.B(_0634_),
    .C(_0635_),
    .A(_0633_),
    .Y(_0637_),
    .D(_0636_));
 sg13g2_xnor2_1 _1915_ (.Y(_0638_),
    .A(\game_inst.snake_inst.pos[7] ),
    .B(net1146));
 sg13g2_a22oi_1 _1916_ (.Y(_0639_),
    .B1(_0198_),
    .B2(net1298),
    .A2(\game_inst.snake_inst.length[4] ),
    .A1(_0189_));
 sg13g2_nand2b_1 _1917_ (.Y(_0640_),
    .B(\game_inst.snake_inst.length[0] ),
    .A_N(\game_inst.snake_inst.pos[0] ));
 sg13g2_o21ai_1 _1918_ (.B1(_0640_),
    .Y(_0641_),
    .A1(\game_inst.snake_inst.pos[3] ),
    .A2(_0196_));
 sg13g2_a221oi_1 _1919_ (.B2(net1168),
    .C1(_0641_),
    .B1(_0197_),
    .A1(\game_inst.snake_inst.pos[1] ),
    .Y(_0642_),
    .A2(_0195_));
 sg13g2_nand3_1 _1920_ (.B(net1299),
    .C(_0642_),
    .A(_0638_),
    .Y(_0643_));
 sg13g2_o21ai_1 _1921_ (.B1(net1263),
    .Y(_0644_),
    .A1(_0637_),
    .A2(net1300));
 sg13g2_a21oi_1 _1922_ (.A1(_0436_),
    .A2(net1301),
    .Y(_0097_),
    .B1(net132));
 sg13g2_and2_1 _1923_ (.A(net1139),
    .B(_0436_),
    .X(_0645_));
 sg13g2_nand2_1 _1924_ (.Y(_0646_),
    .A(net1139),
    .B(_0436_));
 sg13g2_a22oi_1 _1925_ (.Y(_0647_),
    .B1(net106),
    .B2(_0583_),
    .A2(_0435_),
    .A1(net1334));
 sg13g2_a21oi_1 _1926_ (.A1(_0432_),
    .A2(_0584_),
    .Y(_0648_),
    .B1(_0647_));
 sg13g2_xnor2_1 _1927_ (.Y(_0098_),
    .A(_0645_),
    .B(_0648_));
 sg13g2_nand2b_2 _1928_ (.Y(_0649_),
    .B(\game_inst.snake_inst.dir_first[0] ),
    .A_N(\game_inst.snake_inst.dir_first[1] ));
 sg13g2_and2_1 _1929_ (.A(\game_inst.apple_inst.i_snake_y[1] ),
    .B(_0649_),
    .X(_0650_));
 sg13g2_xnor2_1 _1930_ (.Y(_0651_),
    .A(_0210_),
    .B(_0649_));
 sg13g2_xor2_1 _1931_ (.B(_0651_),
    .A(\game_inst.apple_inst.i_snake_y[0] ),
    .X(_0652_));
 sg13g2_o21ai_1 _1932_ (.B1(_0436_),
    .Y(_0653_),
    .A1(net1139),
    .A2(_0652_));
 sg13g2_o21ai_1 _1933_ (.B1(_0653_),
    .Y(_0654_),
    .A1(net107),
    .A2(_0586_));
 sg13g2_inv_1 _1934_ (.Y(_0655_),
    .A(_0654_));
 sg13g2_a22oi_1 _1935_ (.Y(_0099_),
    .B1(_0655_),
    .B2(_0592_),
    .A2(_0645_),
    .A1(_0210_));
 sg13g2_nor2_1 _1936_ (.A(\game_inst.apple_inst.i_snake_y[2] ),
    .B(_0649_),
    .Y(_0656_));
 sg13g2_nand2_1 _1937_ (.Y(_0657_),
    .A(\game_inst.apple_inst.i_snake_y[2] ),
    .B(_0649_));
 sg13g2_nor2b_1 _1938_ (.A(_0656_),
    .B_N(_0657_),
    .Y(_0658_));
 sg13g2_a21oi_1 _1939_ (.A1(\game_inst.apple_inst.i_snake_y[0] ),
    .A2(_0651_),
    .Y(_0659_),
    .B1(_0650_));
 sg13g2_xor2_1 _1940_ (.B(_0659_),
    .A(_0658_),
    .X(_0660_));
 sg13g2_a22oi_1 _1941_ (.Y(_0661_),
    .B1(_0660_),
    .B2(net107),
    .A2(_0593_),
    .A1(net106));
 sg13g2_nor3_1 _1942_ (.A(_0602_),
    .B(_0645_),
    .C(_0661_),
    .Y(_0662_));
 sg13g2_a21oi_1 _1943_ (.A1(_0211_),
    .A2(_0645_),
    .Y(_0100_),
    .B1(_0662_));
 sg13g2_o21ai_1 _1944_ (.B1(_0657_),
    .Y(_0663_),
    .A1(_0656_),
    .A2(_0659_));
 sg13g2_xnor2_1 _1945_ (.Y(_0664_),
    .A(_0213_),
    .B(_0649_));
 sg13g2_xnor2_1 _1946_ (.Y(_0665_),
    .A(_0663_),
    .B(_0664_));
 sg13g2_nand3_1 _1947_ (.B(_0646_),
    .C(_0665_),
    .A(net107),
    .Y(_0666_));
 sg13g2_o21ai_1 _1948_ (.B1(net106),
    .Y(_0667_),
    .A1(_0170_),
    .A2(_0432_));
 sg13g2_a21oi_1 _1949_ (.A1(_0666_),
    .A2(_0667_),
    .Y(_0668_),
    .B1(_0607_));
 sg13g2_a21oi_1 _1950_ (.A1(_0213_),
    .A2(_0645_),
    .Y(_0101_),
    .B1(_0668_));
 sg13g2_xnor2_1 _1951_ (.Y(_0669_),
    .A(net1296),
    .B(eat));
 sg13g2_nand2_1 _1952_ (.Y(_0102_),
    .A(net112),
    .B(_0669_));
 sg13g2_a21oi_1 _1953_ (.A1(\game_inst.snake_inst.length[0] ),
    .A2(eat),
    .Y(_0670_),
    .B1(net1198));
 sg13g2_and3_2 _1954_ (.X(_0671_),
    .A(\game_inst.snake_inst.length[0] ),
    .B(net1198),
    .C(eat));
 sg13g2_nor3_1 _1955_ (.A(net131),
    .B(net1199),
    .C(_0671_),
    .Y(_0103_));
 sg13g2_xnor2_1 _1956_ (.Y(_0672_),
    .A(net1274),
    .B(_0671_));
 sg13g2_nor2_1 _1957_ (.A(net131),
    .B(net1275),
    .Y(_0104_));
 sg13g2_a21oi_1 _1958_ (.A1(\game_inst.snake_inst.length[2] ),
    .A2(_0671_),
    .Y(_0673_),
    .B1(net1174));
 sg13g2_nand3_1 _1959_ (.B(net1174),
    .C(_0671_),
    .A(net1274),
    .Y(_0674_));
 sg13g2_nand2_1 _1960_ (.Y(_0675_),
    .A(net112),
    .B(_0674_));
 sg13g2_nor2_1 _1961_ (.A(net1175),
    .B(_0675_),
    .Y(_0105_));
 sg13g2_and2_1 _1962_ (.A(_0197_),
    .B(_0674_),
    .X(_0676_));
 sg13g2_and4_1 _1963_ (.A(net1274),
    .B(net1174),
    .C(net1322),
    .D(_0671_),
    .X(_0677_));
 sg13g2_nor3_1 _1964_ (.A(net131),
    .B(_0676_),
    .C(_0677_),
    .Y(_0106_));
 sg13g2_and2_1 _1965_ (.A(net1277),
    .B(_0677_),
    .X(_0678_));
 sg13g2_o21ai_1 _1966_ (.B1(net112),
    .Y(_0679_),
    .A1(net1277),
    .A2(_0677_));
 sg13g2_nor2_1 _1967_ (.A(_0678_),
    .B(net1278),
    .Y(_0107_));
 sg13g2_nor2_1 _1968_ (.A(net1265),
    .B(_0678_),
    .Y(_0680_));
 sg13g2_and2_1 _1969_ (.A(net1265),
    .B(_0678_),
    .X(_0681_));
 sg13g2_nor3_1 _1970_ (.A(net131),
    .B(net1266),
    .C(_0681_),
    .Y(_0108_));
 sg13g2_o21ai_1 _1971_ (.B1(net112),
    .Y(_0682_),
    .A1(net1146),
    .A2(_0681_));
 sg13g2_a21oi_1 _1972_ (.A1(net1146),
    .A2(_0681_),
    .Y(_0109_),
    .B1(_0682_));
 sg13g2_nand2_1 _1973_ (.Y(_0683_),
    .A(net112),
    .B(_0436_));
 sg13g2_nor3_1 _1974_ (.A(_0232_),
    .B(_0438_),
    .C(_0683_),
    .Y(_0110_));
 sg13g2_nor2_1 _1975_ (.A(net1259),
    .B(_0438_),
    .Y(_0684_));
 sg13g2_nor3_1 _1976_ (.A(_0439_),
    .B(_0683_),
    .C(net1260),
    .Y(_0111_));
 sg13g2_a21oi_1 _1977_ (.A1(\game_inst.snake_inst.pos[3] ),
    .A2(_0439_),
    .Y(_0685_),
    .B1(net1168));
 sg13g2_nor3_1 _1978_ (.A(_0441_),
    .B(_0683_),
    .C(net1169),
    .Y(_0112_));
 sg13g2_nand2b_1 _1979_ (.Y(_0686_),
    .B(_0467_),
    .A_N(_0406_));
 sg13g2_mux2_1 _1980_ (.A0(net99),
    .A1(net1216),
    .S(_0686_),
    .X(_0113_));
 sg13g2_mux2_1 _1981_ (.A0(net96),
    .A1(net1187),
    .S(_0686_),
    .X(_0114_));
 sg13g2_nand2_1 _1982_ (.Y(_0687_),
    .A(_0420_),
    .B(_0425_));
 sg13g2_mux2_1 _1983_ (.A0(net101),
    .A1(net1197),
    .S(_0687_),
    .X(_0115_));
 sg13g2_mux2_1 _1984_ (.A0(net98),
    .A1(net1205),
    .S(_0687_),
    .X(_0116_));
 sg13g2_nor2_1 _1985_ (.A(net1220),
    .B(net104),
    .Y(_0688_));
 sg13g2_a21oi_1 _1986_ (.A1(_0180_),
    .A2(net104),
    .Y(_0117_),
    .B1(_0688_));
 sg13g2_mux2_1 _1987_ (.A0(net1245),
    .A1(net1227),
    .S(net104),
    .X(_0118_));
 sg13g2_nor2_1 _1988_ (.A(\game_inst.apple_inst.apple_y[2] ),
    .B(net104),
    .Y(_0689_));
 sg13g2_a21oi_1 _1989_ (.A1(_0179_),
    .A2(net104),
    .Y(_0119_),
    .B1(_0689_));
 sg13g2_mux2_1 _1990_ (.A0(net1240),
    .A1(net1233),
    .S(net104),
    .X(_0120_));
 sg13g2_a21oi_1 _1991_ (.A1(_0192_),
    .A2(_0587_),
    .Y(_0121_),
    .B1(net132));
 sg13g2_nor2_1 _1992_ (.A(_0415_),
    .B(_0466_),
    .Y(_0690_));
 sg13g2_mux2_1 _1993_ (.A0(net1188),
    .A1(net100),
    .S(_0690_),
    .X(_0122_));
 sg13g2_mux2_1 _1994_ (.A0(net1196),
    .A1(net97),
    .S(_0690_),
    .X(_0123_));
 sg13g2_nor2b_2 _1995_ (.A(\game_inst.tickgen_inst.prev_user_input ),
    .B_N(net7),
    .Y(_0691_));
 sg13g2_a21oi_1 _1996_ (.A1(net5),
    .A2(_0691_),
    .Y(_0692_),
    .B1(net1268));
 sg13g2_and3_1 _1997_ (.X(_0693_),
    .A(net1268),
    .B(net5),
    .C(_0691_));
 sg13g2_nor3_1 _1998_ (.A(net135),
    .B(net1269),
    .C(_0693_),
    .Y(_0124_));
 sg13g2_nor2b_2 _1999_ (.A(\game_inst.tickgen_inst.prev_vsync ),
    .B_N(\game_inst.tickgen_inst.i_vsync ),
    .Y(_0694_));
 sg13g2_xor2_1 _2000_ (.B(\game_inst.tickgen_inst.counter_max[3] ),
    .A(\game_inst.tickgen_inst.counter[3] ),
    .X(_0695_));
 sg13g2_a221oi_1 _2001_ (.B2(_0163_),
    .C1(_0695_),
    .B1(\game_inst.tickgen_inst.counter_max[0] ),
    .A1(\game_inst.tickgen_inst.counter[4] ),
    .Y(_0696_),
    .A2(_0164_));
 sg13g2_xor2_1 _2002_ (.B(\game_inst.tickgen_inst.counter_max[2] ),
    .A(\game_inst.tickgen_inst.counter[2] ),
    .X(_0697_));
 sg13g2_a221oi_1 _2003_ (.B2(_0162_),
    .C1(_0697_),
    .B1(\game_inst.tickgen_inst.counter_max[1] ),
    .A1(_0161_),
    .Y(_0698_),
    .A2(net1144));
 sg13g2_a22oi_1 _2004_ (.Y(_0699_),
    .B1(_0166_),
    .B2(\game_inst.tickgen_inst.counter[0] ),
    .A2(_0165_),
    .A1(\game_inst.tickgen_inst.counter[1] ));
 sg13g2_nand4_1 _2005_ (.B(_0696_),
    .C(_0698_),
    .A(_0694_),
    .Y(_0700_),
    .D(_0699_));
 sg13g2_o21ai_1 _2006_ (.B1(net139),
    .Y(_0701_),
    .A1(_0235_),
    .A2(_0694_));
 sg13g2_a21oi_1 _2007_ (.A1(_0167_),
    .A2(_0700_),
    .Y(_0125_),
    .B1(_0701_));
 sg13g2_nand2b_2 _2008_ (.Y(_0702_),
    .B(_0691_),
    .A_N(_0352_));
 sg13g2_o21ai_1 _2009_ (.B1(net139),
    .Y(_0703_),
    .A1(_0166_),
    .A2(_0702_));
 sg13g2_a21oi_1 _2010_ (.A1(_0166_),
    .A2(_0702_),
    .Y(_0126_),
    .B1(_0703_));
 sg13g2_nor2_1 _2011_ (.A(_0165_),
    .B(net136),
    .Y(_0704_));
 sg13g2_xnor2_1 _2012_ (.Y(_0705_),
    .A(net1280),
    .B(net136));
 sg13g2_a21oi_1 _2013_ (.A1(\game_inst.tickgen_inst.counter_max[0] ),
    .A2(_0705_),
    .Y(_0706_),
    .B1(_0702_));
 sg13g2_o21ai_1 _2014_ (.B1(_0706_),
    .Y(_0707_),
    .A1(\game_inst.tickgen_inst.counter_max[0] ),
    .A2(_0705_));
 sg13g2_a21oi_1 _2015_ (.A1(net1280),
    .A2(_0702_),
    .Y(_0708_),
    .B1(net135));
 sg13g2_nand2_1 _2016_ (.Y(_0127_),
    .A(_0707_),
    .B(net1281));
 sg13g2_nand2b_1 _2017_ (.Y(_0709_),
    .B(\game_inst.tickgen_inst.counter_max[2] ),
    .A_N(net136));
 sg13g2_xor2_1 _2018_ (.B(net136),
    .A(net1302),
    .X(_0710_));
 sg13g2_a21oi_1 _2019_ (.A1(net1285),
    .A2(_0705_),
    .Y(_0711_),
    .B1(_0704_));
 sg13g2_or2_1 _2020_ (.X(_0712_),
    .B(_0711_),
    .A(_0710_));
 sg13g2_a21oi_1 _2021_ (.A1(_0710_),
    .A2(_0711_),
    .Y(_0713_),
    .B1(_0702_));
 sg13g2_a22oi_1 _2022_ (.Y(_0714_),
    .B1(_0712_),
    .B2(_0713_),
    .A2(_0702_),
    .A1(net1302));
 sg13g2_nand2_1 _2023_ (.Y(_0128_),
    .A(net139),
    .B(net1303));
 sg13g2_and2_1 _2024_ (.A(_0709_),
    .B(_0712_),
    .X(_0715_));
 sg13g2_nor2_1 _2025_ (.A(net136),
    .B(_0715_),
    .Y(_0716_));
 sg13g2_or2_1 _2026_ (.X(_0717_),
    .B(_0716_),
    .A(_0702_));
 sg13g2_a21oi_1 _2027_ (.A1(net136),
    .A2(_0712_),
    .Y(_0718_),
    .B1(_0717_));
 sg13g2_xnor2_1 _2028_ (.Y(_0719_),
    .A(net1276),
    .B(_0718_));
 sg13g2_nand2_1 _2029_ (.Y(_0129_),
    .A(net139),
    .B(_0719_));
 sg13g2_mux2_1 _2030_ (.A0(net2),
    .A1(_0715_),
    .S(\game_inst.tickgen_inst.counter_max[3] ),
    .X(_0720_));
 sg13g2_nor2_1 _2031_ (.A(_0717_),
    .B(_0720_),
    .Y(_0721_));
 sg13g2_o21ai_1 _2032_ (.B1(net139),
    .Y(_0722_),
    .A1(net1144),
    .A2(_0721_));
 sg13g2_a21oi_1 _2033_ (.A1(net1144),
    .A2(_0721_),
    .Y(_0130_),
    .B1(_0722_));
 sg13g2_nand2_2 _2034_ (.Y(_0723_),
    .A(net1),
    .B(_0700_));
 sg13g2_inv_1 _2035_ (.Y(_0724_),
    .A(_0723_));
 sg13g2_and2_1 _2036_ (.A(net1254),
    .B(_0694_),
    .X(_0725_));
 sg13g2_nor2_1 _2037_ (.A(net1254),
    .B(_0694_),
    .Y(_0726_));
 sg13g2_nor3_1 _2038_ (.A(_0723_),
    .B(_0725_),
    .C(net1255),
    .Y(_0131_));
 sg13g2_and2_1 _2039_ (.A(net1251),
    .B(_0725_),
    .X(_0727_));
 sg13g2_nor2_1 _2040_ (.A(net1251),
    .B(_0725_),
    .Y(_0728_));
 sg13g2_nor3_1 _2041_ (.A(_0723_),
    .B(_0727_),
    .C(net1252),
    .Y(_0132_));
 sg13g2_and2_1 _2042_ (.A(net1262),
    .B(_0727_),
    .X(_0137_));
 sg13g2_nor2_1 _2043_ (.A(net1262),
    .B(_0727_),
    .Y(_0138_));
 sg13g2_nor3_1 _2044_ (.A(_0723_),
    .B(_0137_),
    .C(_0138_),
    .Y(_0133_));
 sg13g2_nand2_1 _2045_ (.Y(_0139_),
    .A(net1290),
    .B(_0137_));
 sg13g2_o21ai_1 _2046_ (.B1(_0724_),
    .Y(_0140_),
    .A1(net1290),
    .A2(_0137_));
 sg13g2_nor2b_1 _2047_ (.A(_0140_),
    .B_N(_0139_),
    .Y(_0134_));
 sg13g2_xnor2_1 _2048_ (.Y(_0141_),
    .A(_0161_),
    .B(_0139_));
 sg13g2_nor2_1 _2049_ (.A(_0723_),
    .B(_0141_),
    .Y(_0135_));
 sg13g2_xnor2_1 _2050_ (.Y(_0142_),
    .A(\game_inst.head_x[2] ),
    .B(\game_inst.apple_inst.i_snake_x[2] ));
 sg13g2_xor2_1 _2051_ (.B(\game_inst.apple_inst.i_snake_y[2] ),
    .A(net119),
    .X(_0143_));
 sg13g2_xor2_1 _2052_ (.B(\game_inst.apple_inst.i_snake_y[3] ),
    .A(\game_inst.head_y[3] ),
    .X(_0144_));
 sg13g2_xor2_1 _2053_ (.B(\game_inst.apple_inst.i_snake_y[0] ),
    .A(\game_inst.head_y[0] ),
    .X(_0145_));
 sg13g2_a221oi_1 _2054_ (.B2(_0176_),
    .C1(_0144_),
    .B1(\game_inst.apple_inst.i_snake_x[1] ),
    .A1(_0177_),
    .Y(_0146_),
    .A2(net117));
 sg13g2_xor2_1 _2055_ (.B(\game_inst.apple_inst.i_snake_x[3] ),
    .A(net121),
    .X(_0147_));
 sg13g2_a22oi_1 _2056_ (.Y(_0148_),
    .B1(\game_inst.apple_inst.i_snake_y[1] ),
    .B2(_0172_),
    .A2(_0201_),
    .A1(\game_inst.head_x[1] ));
 sg13g2_xnor2_1 _2057_ (.Y(_0149_),
    .A(\game_inst.head_x[4] ),
    .B(\game_inst.apple_inst.i_snake_x[4] ));
 sg13g2_a22oi_1 _2058_ (.Y(_0150_),
    .B1(_0210_),
    .B2(net120),
    .A2(_0200_),
    .A1(\game_inst.head_x[0] ));
 sg13g2_nand4_1 _2059_ (.B(_0148_),
    .C(_0149_),
    .A(_0142_),
    .Y(_0151_),
    .D(_0150_));
 sg13g2_nor4_1 _2060_ (.A(_0143_),
    .B(_0145_),
    .C(_0147_),
    .D(_0151_),
    .Y(_0152_));
 sg13g2_a21oi_1 _2061_ (.A1(\game_inst.head_x[1] ),
    .A2(\game_inst.head_x[0] ),
    .Y(_0153_),
    .B1(_0174_));
 sg13g2_a21oi_1 _2062_ (.A1(_0176_),
    .A2(_0177_),
    .Y(_0154_),
    .B1(\game_inst.head_x[4] ));
 sg13g2_nor4_1 _2063_ (.A(\game_inst.head_x[3] ),
    .B(\game_inst.head_x[2] ),
    .C(_0153_),
    .D(_0154_),
    .Y(_0155_));
 sg13g2_o21ai_1 _2064_ (.B1(_0170_),
    .Y(_0156_),
    .A1(net119),
    .A2(net120));
 sg13g2_nand2_1 _2065_ (.Y(_0157_),
    .A(\game_inst.head_y[2] ),
    .B(net120));
 sg13g2_a21oi_1 _2066_ (.A1(\game_inst.head_y[3] ),
    .A2(_0157_),
    .Y(_0158_),
    .B1(\game_inst.head_y[0] ));
 sg13g2_a221oi_1 _2067_ (.B2(_0158_),
    .C1(_0155_),
    .B1(_0156_),
    .A1(_0146_),
    .Y(_0159_),
    .A2(_0152_));
 sg13g2_nand3b_1 _2068_ (.B(\game_inst.apple_inst.i_snake_valid ),
    .C(_0235_),
    .Y(_0160_),
    .A_N(_0159_));
 sg13g2_a21oi_1 _2069_ (.A1(_0191_),
    .A2(_0160_),
    .Y(_0136_),
    .B1(net131));
 sg13g2_dfrbpq_1 _2070_ (.RESET_B(net59),
    .D(_0003_),
    .Q(\game_inst.vga_inst.row_buffer[0][0] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _2071_ (.RESET_B(net91),
    .D(_0004_),
    .Q(\game_inst.vga_inst.row_buffer[0][1] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _2072_ (.RESET_B(net90),
    .D(_0005_),
    .Q(\game_inst.vga_inst.row_buffer[10][0] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2073_ (.RESET_B(net89),
    .D(_0006_),
    .Q(\game_inst.vga_inst.row_buffer[10][1] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2074_ (.RESET_B(net88),
    .D(_0007_),
    .Q(\game_inst.vga_inst.row_buffer[7][0] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2075_ (.RESET_B(net87),
    .D(_0008_),
    .Q(\game_inst.vga_inst.row_buffer[7][1] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2076_ (.RESET_B(net86),
    .D(_0009_),
    .Q(\game_inst.vga_inst.row_buffer[6][0] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2077_ (.RESET_B(net85),
    .D(_0010_),
    .Q(\game_inst.vga_inst.row_buffer[6][1] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _2078_ (.RESET_B(net84),
    .D(net1207),
    .Q(\game_inst.snake_inst.pos[0] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _2079_ (.RESET_B(net83),
    .D(_0012_),
    .Q(\game_inst.snake_inst.pos[3] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _2080_ (.RESET_B(net82),
    .D(_0013_),
    .Q(\game_inst.snake_inst.pos[5] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _2081_ (.RESET_B(net81),
    .D(_0014_),
    .Q(\game_inst.snake_inst.pos[6] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _2082_ (.RESET_B(net80),
    .D(_0015_),
    .Q(\game_inst.snake_inst.pos[7] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2083_ (.RESET_B(net79),
    .D(_0016_),
    .Q(\game_inst.vga_inst.row_buffer[8][0] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2084_ (.RESET_B(net78),
    .D(_0017_),
    .Q(\game_inst.vga_inst.row_buffer[8][1] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _2085_ (.RESET_B(net77),
    .D(_0018_),
    .Q(\game_inst.vga_inst.px[0] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _2086_ (.RESET_B(net76),
    .D(_0019_),
    .Q(\game_inst.vga_inst.px[1] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _2087_ (.RESET_B(net75),
    .D(net1143),
    .Q(\game_inst.vga_inst.px[2] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _2088_ (.RESET_B(net74),
    .D(net1231),
    .Q(\game_inst.vga_inst.px[3] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _2089_ (.RESET_B(net73),
    .D(_0022_),
    .Q(\game_inst.vga_inst.px[4] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _2090_ (.RESET_B(net72),
    .D(_0023_),
    .Q(\game_inst.vga_inst.px[5] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _2091_ (.RESET_B(net71),
    .D(_0024_),
    .Q(\game_inst.vga_inst.px[6] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _2092_ (.RESET_B(net69),
    .D(_0025_),
    .Q(\game_inst.vga_inst.px[7] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _2093_ (.RESET_B(net68),
    .D(_0026_),
    .Q(\game_inst.vga_inst.px[8] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _2094_ (.RESET_B(net67),
    .D(_0027_),
    .Q(\game_inst.vga_inst.px[9] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _2095_ (.RESET_B(net66),
    .D(_0028_),
    .Q(\game_inst.vga_inst.row_buffer[4][0] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2096_ (.RESET_B(net65),
    .D(_0029_),
    .Q(\game_inst.vga_inst.row_buffer[4][1] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2097_ (.RESET_B(net64),
    .D(_0030_),
    .Q(\game_inst.vga_inst.row_buffer[17][0] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2098_ (.RESET_B(net63),
    .D(_0031_),
    .Q(\game_inst.vga_inst.row_buffer[17][1] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2099_ (.RESET_B(net62),
    .D(_0032_),
    .Q(\game_inst.vga_inst.row_buffer[5][0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2100_ (.RESET_B(net61),
    .D(_0033_),
    .Q(\game_inst.vga_inst.row_buffer[5][1] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2101_ (.RESET_B(net60),
    .D(_0034_),
    .Q(\game_inst.vga_inst.row_buffer[13][0] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _2102_ (.RESET_B(net58),
    .D(_0035_),
    .Q(\game_inst.vga_inst.row_buffer[13][1] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _2103_ (.RESET_B(net57),
    .D(_0036_),
    .Q(\game_inst.vga_inst.row_buffer[9][0] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2104_ (.RESET_B(net56),
    .D(_0037_),
    .Q(\game_inst.vga_inst.row_buffer[9][1] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _2105_ (.RESET_B(net55),
    .D(net1153),
    .Q(\game_inst.snake_inst.dir_first[0] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _2106_ (.RESET_B(net54),
    .D(_0039_),
    .Q(\game_inst.snake_inst.dir_first[1] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _2107_ (.RESET_B(net53),
    .D(_0040_),
    .Q(\game_inst.vga_inst.row_buffer[15][0] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _2108_ (.RESET_B(net52),
    .D(_0041_),
    .Q(\game_inst.vga_inst.row_buffer[15][1] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2109_ (.RESET_B(net51),
    .D(net1138),
    .Q(\game_inst.vga_inst.pos_counter[0] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2110_ (.RESET_B(net70),
    .D(net1159),
    .Q(\game_inst.vga_inst.pos_counter[1] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2111_ (.RESET_B(net50),
    .D(net1328),
    .Q(\game_inst.o_vga_hsync ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _2112_ (.RESET_B(net49),
    .D(_0044_),
    .Q(\game_inst.vga_inst.py[0] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _2113_ (.RESET_B(net47),
    .D(net1186),
    .Q(\game_inst.vga_inst.py[1] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _2114_ (.RESET_B(net45),
    .D(net1183),
    .Q(\game_inst.vga_inst.py[2] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _2115_ (.RESET_B(net43),
    .D(net1167),
    .Q(\game_inst.vga_inst.py[3] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _2116_ (.RESET_B(net41),
    .D(_0048_),
    .Q(\game_inst.vga_inst.py[4] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _2117_ (.RESET_B(net39),
    .D(_0049_),
    .Q(\game_inst.vga_inst.py[5] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _2118_ (.RESET_B(net37),
    .D(_0050_),
    .Q(\game_inst.vga_inst.py[6] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _2119_ (.RESET_B(net35),
    .D(net1242),
    .Q(\game_inst.vga_inst.py[7] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _2120_ (.RESET_B(net33),
    .D(_0052_),
    .Q(\game_inst.vga_inst.py[8] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _2121_ (.RESET_B(net173),
    .D(net1218),
    .Q(\game_inst.vga_inst.py[9] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _2122_ (.RESET_B(net31),
    .D(_0002_),
    .Q(\game_inst.o_vga_vsync ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _2123_ (.RESET_B(net29),
    .D(_0054_),
    .Q(\game_inst.o_success ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _2124_ (.RESET_B(net28),
    .D(net1193),
    .Q(\game_inst.apple_inst.apple_x[0] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _2125_ (.RESET_B(net27),
    .D(net1163),
    .Q(\game_inst.apple_inst.apple_x[1] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _2126_ (.RESET_B(net26),
    .D(net1179),
    .Q(\game_inst.apple_inst.apple_x[2] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _2127_ (.RESET_B(net25),
    .D(net1165),
    .Q(\game_inst.apple_inst.apple_x[3] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _2128_ (.RESET_B(net24),
    .D(_0059_),
    .Q(\game_inst.apple_inst.apple_x[4] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _2129_ (.RESET_B(net23),
    .D(_0060_),
    .Q(\game_inst.apple_inst.o_ready ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _2130_ (.RESET_B(net21),
    .D(net1151),
    .Q(\game_inst.apple_inst.test ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _2131_ (.RESET_B(net19),
    .D(_0062_),
    .Q(\game_inst.apple_inst.random_inst.lfsr5[0] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _2132_ (.RESET_B(net667),
    .D(_0063_),
    .Q(\game_inst.apple_inst.random_inst.lfsr5[1] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _2133_ (.RESET_B(net665),
    .D(_0064_),
    .Q(\game_inst.apple_inst.random_inst.lfsr5[2] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _2134_ (.RESET_B(net663),
    .D(_0065_),
    .Q(\game_inst.apple_inst.random_inst.lfsr5[3] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _2135_ (.RESET_B(net661),
    .D(_0066_),
    .Q(\game_inst.apple_inst.random_inst.lfsr5[4] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _2136_ (.RESET_B(net659),
    .D(net1155),
    .Q(\game_inst.apple_inst.random_inst.lfsr4[0] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _2137_ (.RESET_B(net657),
    .D(_0068_),
    .Q(\game_inst.apple_inst.random_inst.lfsr4[1] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _2138_ (.RESET_B(net653),
    .D(_0069_),
    .Q(\game_inst.apple_inst.random_inst.lfsr4[2] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _2139_ (.RESET_B(net651),
    .D(_0070_),
    .Q(\game_inst.apple_inst.random_inst.lfsr4[3] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _2140_ (.RESET_B(net649),
    .D(_0071_),
    .Q(\game_inst.vga_inst.row_buffer[2][0] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _2141_ (.RESET_B(net648),
    .D(_0072_),
    .Q(\game_inst.vga_inst.row_buffer[2][1] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _2142_ (.RESET_B(net647),
    .D(_0073_),
    .Q(\game_inst.vga_inst.row_buffer[3][0] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _2143_ (.RESET_B(net646),
    .D(_0074_),
    .Q(\game_inst.vga_inst.row_buffer[3][1] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _2144_ (.RESET_B(net645),
    .D(_0075_),
    .Q(\game_inst.vga_inst.row_buffer[14][0] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2145_ (.RESET_B(net644),
    .D(_0076_),
    .Q(\game_inst.vga_inst.row_buffer[14][1] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2146_ (.RESET_B(net643),
    .D(_0077_),
    .Q(\game_inst.vga_inst.row_buffer[12][0] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _2147_ (.RESET_B(net642),
    .D(_0078_),
    .Q(\game_inst.vga_inst.row_buffer[12][1] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _2148_ (.RESET_B(net641),
    .D(net1157),
    .Q(\game_inst.control_inst.i_head_dir[0] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _2149_ (.RESET_B(net639),
    .D(net1250),
    .Q(\game_inst.control_inst.backwards[1] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _2150_ (.RESET_B(net171),
    .D(net1321),
    .Q(\game_inst.head_x[0] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _2151_ (.RESET_B(net169),
    .D(_0082_),
    .Q(\game_inst.head_x[1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _2152_ (.RESET_B(net167),
    .D(_0083_),
    .Q(\game_inst.head_x[2] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2153_ (.RESET_B(net165),
    .D(net1332),
    .Q(\game_inst.head_x[3] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _2154_ (.RESET_B(net163),
    .D(_0085_),
    .Q(\game_inst.head_x[4] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _2155_ (.RESET_B(net161),
    .D(net1315),
    .Q(\game_inst.head_y[0] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _2156_ (.RESET_B(net159),
    .D(net1293),
    .Q(\game_inst.head_y[1] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _2157_ (.RESET_B(net157),
    .D(_0088_),
    .Q(\game_inst.head_y[2] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _2158_ (.RESET_B(net155),
    .D(_0089_),
    .Q(\game_inst.head_y[3] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _2159_ (.RESET_B(net153),
    .D(_0090_),
    .Q(\game_inst.control_inst.dir[0] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _2160_ (.RESET_B(net152),
    .D(_0091_),
    .Q(\game_inst.control_inst.dir[1] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _2161_ (.RESET_B(net151),
    .D(_0092_),
    .Q(\game_inst.apple_inst.i_snake_x[0] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _2162_ (.RESET_B(net150),
    .D(net1324),
    .Q(\game_inst.apple_inst.i_snake_x[1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _2163_ (.RESET_B(net149),
    .D(_0094_),
    .Q(\game_inst.apple_inst.i_snake_x[2] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _2164_ (.RESET_B(net148),
    .D(net1319),
    .Q(\game_inst.apple_inst.i_snake_x[3] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _2165_ (.RESET_B(net147),
    .D(_0096_),
    .Q(\game_inst.apple_inst.i_snake_x[4] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _2166_ (.RESET_B(net146),
    .D(_0097_),
    .Q(\game_inst.apple_inst.i_snake_valid ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _2167_ (.RESET_B(net144),
    .D(_0098_),
    .Q(\game_inst.apple_inst.i_snake_y[0] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _2168_ (.RESET_B(net143),
    .D(net1308),
    .Q(\game_inst.apple_inst.i_snake_y[1] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _2169_ (.RESET_B(net142),
    .D(_0100_),
    .Q(\game_inst.apple_inst.i_snake_y[2] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _2170_ (.RESET_B(net141),
    .D(_0101_),
    .Q(\game_inst.apple_inst.i_snake_y[3] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _2171_ (.RESET_B(net140),
    .D(_0102_),
    .Q(\game_inst.snake_inst.length[0] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _2172_ (.RESET_B(net93),
    .D(net1200),
    .Q(\game_inst.snake_inst.length[1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _2173_ (.RESET_B(net92),
    .D(_0104_),
    .Q(\game_inst.snake_inst.length[2] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _2174_ (.RESET_B(net48),
    .D(net1176),
    .Q(\game_inst.snake_inst.length[3] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _2175_ (.RESET_B(net46),
    .D(_0106_),
    .Q(\game_inst.snake_inst.length[4] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _2176_ (.RESET_B(net44),
    .D(net1279),
    .Q(\game_inst.snake_inst.length[5] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _2177_ (.RESET_B(net42),
    .D(net1267),
    .Q(\game_inst.snake_inst.length[6] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _2178_ (.RESET_B(net174),
    .D(net1147),
    .Q(\game_inst.snake_inst.length[7] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _2179_ (.RESET_B(net175),
    .D(net1026),
    .Q(\game_inst.snake_inst.dir_out[0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2180_ (.RESET_B(net176),
    .D(net1059),
    .Q(\game_inst.snake_inst.dir_out[1] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _2181_ (.RESET_B(net177),
    .D(net762),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[232][0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2182_ (.RESET_B(net178),
    .D(net820),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[232][1] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _2183_ (.RESET_B(net179),
    .D(net1060),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[231][0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2184_ (.RESET_B(net180),
    .D(net955),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[231][1] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _2185_ (.RESET_B(net181),
    .D(net1028),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[230][0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2186_ (.RESET_B(net182),
    .D(net847),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[230][1] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _2187_ (.RESET_B(net183),
    .D(net1040),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[229][0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2188_ (.RESET_B(net184),
    .D(net676),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[229][1] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _2189_ (.RESET_B(net185),
    .D(net714),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[228][0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2190_ (.RESET_B(net186),
    .D(net876),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[228][1] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _2191_ (.RESET_B(net187),
    .D(net1080),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[227][0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2192_ (.RESET_B(net188),
    .D(net807),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[227][1] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _2193_ (.RESET_B(net189),
    .D(net819),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[226][0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _2194_ (.RESET_B(net190),
    .D(net718),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[226][1] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _2195_ (.RESET_B(net191),
    .D(net708),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[225][0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _2196_ (.RESET_B(net192),
    .D(net1102),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[225][1] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _2197_ (.RESET_B(net193),
    .D(net986),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[224][0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _2198_ (.RESET_B(net194),
    .D(net679),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[224][1] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _2199_ (.RESET_B(net195),
    .D(net1000),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[223][0] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _2200_ (.RESET_B(net196),
    .D(net1054),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[223][1] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _2201_ (.RESET_B(net197),
    .D(net865),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[222][0] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _2202_ (.RESET_B(net198),
    .D(net674),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[222][1] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _2203_ (.RESET_B(net199),
    .D(net1083),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[221][0] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _2204_ (.RESET_B(net200),
    .D(net1070),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[221][1] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _2205_ (.RESET_B(net201),
    .D(net1076),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[220][0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _2206_ (.RESET_B(net202),
    .D(net868),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[220][1] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _2207_ (.RESET_B(net203),
    .D(net879),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[219][0] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _2208_ (.RESET_B(net204),
    .D(net1114),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[219][1] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _2209_ (.RESET_B(net205),
    .D(net944),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[218][0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _2210_ (.RESET_B(net206),
    .D(net751),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[218][1] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _2211_ (.RESET_B(net207),
    .D(net1090),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[217][0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _2212_ (.RESET_B(net208),
    .D(net801),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[217][1] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _2213_ (.RESET_B(net209),
    .D(net937),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[216][0] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _2214_ (.RESET_B(net210),
    .D(net886),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[216][1] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _2215_ (.RESET_B(net211),
    .D(net683),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[215][0] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _2216_ (.RESET_B(net212),
    .D(net949),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[215][1] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _2217_ (.RESET_B(net213),
    .D(net1111),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[214][0] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _2218_ (.RESET_B(net214),
    .D(net1093),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[214][1] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _2219_ (.RESET_B(net215),
    .D(net760),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[213][0] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _2220_ (.RESET_B(net216),
    .D(net772),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[213][1] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _2221_ (.RESET_B(net217),
    .D(net763),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[212][0] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _2222_ (.RESET_B(net218),
    .D(net979),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[212][1] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _2223_ (.RESET_B(net219),
    .D(net952),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[211][0] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _2224_ (.RESET_B(net220),
    .D(net837),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[211][1] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _2225_ (.RESET_B(net221),
    .D(net903),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[210][0] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _2226_ (.RESET_B(net222),
    .D(net1017),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[210][1] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _2227_ (.RESET_B(net223),
    .D(net705),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[209][0] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _2228_ (.RESET_B(net224),
    .D(net730),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[209][1] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _2229_ (.RESET_B(net225),
    .D(net1031),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[208][0] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _2230_ (.RESET_B(net226),
    .D(net905),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[208][1] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _2231_ (.RESET_B(net227),
    .D(net971),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[207][0] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _2232_ (.RESET_B(net228),
    .D(net1096),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[207][1] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _2233_ (.RESET_B(net229),
    .D(net1039),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[206][0] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _2234_ (.RESET_B(net230),
    .D(net817),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[206][1] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _2235_ (.RESET_B(net231),
    .D(net699),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[205][0] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _2236_ (.RESET_B(net232),
    .D(net934),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[205][1] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _2237_ (.RESET_B(net233),
    .D(net1038),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[204][0] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _2238_ (.RESET_B(net234),
    .D(net832),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[204][1] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _2239_ (.RESET_B(net235),
    .D(net884),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[203][0] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _2240_ (.RESET_B(net236),
    .D(net977),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[203][1] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _2241_ (.RESET_B(net237),
    .D(net672),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[202][0] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _2242_ (.RESET_B(net238),
    .D(net1072),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[202][1] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _2243_ (.RESET_B(net239),
    .D(net912),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[201][0] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _2244_ (.RESET_B(net240),
    .D(net1032),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[201][1] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _2245_ (.RESET_B(net241),
    .D(net1033),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[200][0] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _2246_ (.RESET_B(net242),
    .D(net1056),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[200][1] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _2247_ (.RESET_B(net243),
    .D(net798),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[199][0] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _2248_ (.RESET_B(net244),
    .D(net716),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[199][1] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _2249_ (.RESET_B(net245),
    .D(net966),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[198][0] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _2250_ (.RESET_B(net246),
    .D(net1109),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[198][1] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _2251_ (.RESET_B(net247),
    .D(net956),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[197][0] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _2252_ (.RESET_B(net248),
    .D(net928),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[197][1] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _2253_ (.RESET_B(net249),
    .D(net929),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[196][0] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _2254_ (.RESET_B(net250),
    .D(net1029),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[196][1] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _2255_ (.RESET_B(net251),
    .D(net1020),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[195][0] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _2256_ (.RESET_B(net252),
    .D(net824),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[195][1] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _2257_ (.RESET_B(net253),
    .D(net945),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[194][0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _2258_ (.RESET_B(net254),
    .D(net997),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[194][1] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _2259_ (.RESET_B(net255),
    .D(net904),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[193][0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _2260_ (.RESET_B(net256),
    .D(net1089),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[193][1] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _2261_ (.RESET_B(net257),
    .D(net900),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[192][0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _2262_ (.RESET_B(net258),
    .D(net1021),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[192][1] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _2263_ (.RESET_B(net259),
    .D(net1097),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[191][0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _2264_ (.RESET_B(net260),
    .D(net1008),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[191][1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _2265_ (.RESET_B(net261),
    .D(net787),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[190][0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _2266_ (.RESET_B(net262),
    .D(net698),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[190][1] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _2267_ (.RESET_B(net263),
    .D(net834),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[189][0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _2268_ (.RESET_B(net264),
    .D(net777),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[189][1] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _2269_ (.RESET_B(net265),
    .D(net1081),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[188][0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _2270_ (.RESET_B(net266),
    .D(net684),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[188][1] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _2271_ (.RESET_B(net267),
    .D(net704),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[187][0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _2272_ (.RESET_B(net268),
    .D(net1098),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[187][1] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _2273_ (.RESET_B(net269),
    .D(net933),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[186][0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _2274_ (.RESET_B(net270),
    .D(net747),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[186][1] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _2275_ (.RESET_B(net271),
    .D(net715),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[185][0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _2276_ (.RESET_B(net272),
    .D(net753),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[185][1] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _2277_ (.RESET_B(net273),
    .D(net1117),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[184][0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _2278_ (.RESET_B(net274),
    .D(net703),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[184][1] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _2279_ (.RESET_B(net275),
    .D(net802),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[183][0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _2280_ (.RESET_B(net276),
    .D(net1132),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[183][1] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _2281_ (.RESET_B(net277),
    .D(net736),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[182][0] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _2282_ (.RESET_B(net278),
    .D(net738),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[182][1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _2283_ (.RESET_B(net279),
    .D(net982),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[181][0] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _2284_ (.RESET_B(net280),
    .D(net836),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[181][1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _2285_ (.RESET_B(net281),
    .D(net675),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[180][0] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _2286_ (.RESET_B(net282),
    .D(net992),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[180][1] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _2287_ (.RESET_B(net283),
    .D(net804),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[179][0] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _2288_ (.RESET_B(net284),
    .D(net913),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[179][1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _2289_ (.RESET_B(net285),
    .D(net853),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[178][0] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _2290_ (.RESET_B(net286),
    .D(net752),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[178][1] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _2291_ (.RESET_B(net287),
    .D(net961),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[177][0] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _2292_ (.RESET_B(net288),
    .D(net788),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[177][1] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _2293_ (.RESET_B(net289),
    .D(net980),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[176][0] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _2294_ (.RESET_B(net290),
    .D(net692),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[176][1] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _2295_ (.RESET_B(net291),
    .D(net862),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[175][0] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _2296_ (.RESET_B(net292),
    .D(net1122),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[175][1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _2297_ (.RESET_B(net293),
    .D(net843),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[174][0] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _2298_ (.RESET_B(net294),
    .D(net938),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[174][1] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _2299_ (.RESET_B(net295),
    .D(net1053),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[173][0] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _2300_ (.RESET_B(net296),
    .D(net895),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[173][1] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _2301_ (.RESET_B(net297),
    .D(net1037),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[172][0] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _2302_ (.RESET_B(net298),
    .D(net790),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[172][1] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _2303_ (.RESET_B(net299),
    .D(net924),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[171][0] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _2304_ (.RESET_B(net300),
    .D(net840),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[171][1] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _2305_ (.RESET_B(net301),
    .D(net726),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[170][0] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _2306_ (.RESET_B(net302),
    .D(net693),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[170][1] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _2307_ (.RESET_B(net303),
    .D(net789),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[169][0] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _2308_ (.RESET_B(net304),
    .D(net936),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[169][1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _2309_ (.RESET_B(net305),
    .D(net1001),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[168][0] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _2310_ (.RESET_B(net306),
    .D(net1124),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[168][1] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _2311_ (.RESET_B(net307),
    .D(net782),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[167][0] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _2312_ (.RESET_B(net308),
    .D(net1061),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[167][1] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _2313_ (.RESET_B(net309),
    .D(net885),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[166][0] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _2314_ (.RESET_B(net310),
    .D(net880),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[166][1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _2315_ (.RESET_B(net311),
    .D(net869),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[165][0] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _2316_ (.RESET_B(net312),
    .D(net901),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[165][1] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _2317_ (.RESET_B(net313),
    .D(net794),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[164][0] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _2318_ (.RESET_B(net314),
    .D(net1023),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[164][1] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _2319_ (.RESET_B(net315),
    .D(net816),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[163][0] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _2320_ (.RESET_B(net316),
    .D(net799),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[163][1] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _2321_ (.RESET_B(net317),
    .D(net963),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[162][0] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _2322_ (.RESET_B(net318),
    .D(net848),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[162][1] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _2323_ (.RESET_B(net319),
    .D(net1058),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[161][0] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _2324_ (.RESET_B(net320),
    .D(net774),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[161][1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _2325_ (.RESET_B(net321),
    .D(net915),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[160][0] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _2326_ (.RESET_B(net322),
    .D(net779),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[160][1] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _2327_ (.RESET_B(net323),
    .D(net998),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[159][0] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _2328_ (.RESET_B(net324),
    .D(net1041),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[159][1] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _2329_ (.RESET_B(net325),
    .D(net682),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[158][0] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _2330_ (.RESET_B(net326),
    .D(net764),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[158][1] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _2331_ (.RESET_B(net327),
    .D(net996),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[157][0] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _2332_ (.RESET_B(net328),
    .D(net737),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[157][1] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _2333_ (.RESET_B(net329),
    .D(net671),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[156][0] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _2334_ (.RESET_B(net330),
    .D(net854),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[156][1] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _2335_ (.RESET_B(net331),
    .D(net825),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[155][0] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _2336_ (.RESET_B(net332),
    .D(net920),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[155][1] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _2337_ (.RESET_B(net333),
    .D(net1074),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[154][0] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _2338_ (.RESET_B(net334),
    .D(net780),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[154][1] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _2339_ (.RESET_B(net335),
    .D(net909),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[153][0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2340_ (.RESET_B(net336),
    .D(net770),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[153][1] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _2341_ (.RESET_B(net337),
    .D(net828),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[152][0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2342_ (.RESET_B(net338),
    .D(net803),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[152][1] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _2343_ (.RESET_B(net339),
    .D(net707),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[151][0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2344_ (.RESET_B(net340),
    .D(net756),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[151][1] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _2345_ (.RESET_B(net341),
    .D(net891),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[150][0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2346_ (.RESET_B(net342),
    .D(net983),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[150][1] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _2347_ (.RESET_B(net343),
    .D(net947),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[149][0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2348_ (.RESET_B(net344),
    .D(net1130),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[149][1] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _2349_ (.RESET_B(net345),
    .D(net870),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[148][0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2350_ (.RESET_B(net346),
    .D(net942),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[148][1] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _2351_ (.RESET_B(net347),
    .D(net742),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[147][0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2352_ (.RESET_B(net348),
    .D(net1126),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[147][1] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _2353_ (.RESET_B(net349),
    .D(net1003),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[146][0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2354_ (.RESET_B(net350),
    .D(net1016),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[146][1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _2355_ (.RESET_B(net351),
    .D(net739),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[145][0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2356_ (.RESET_B(net352),
    .D(net972),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[145][1] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _2357_ (.RESET_B(net353),
    .D(net1123),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[144][0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2358_ (.RESET_B(net354),
    .D(net1128),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[144][1] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _2359_ (.RESET_B(net355),
    .D(net1065),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[143][0] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _2360_ (.RESET_B(net356),
    .D(net898),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[143][1] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _2361_ (.RESET_B(net357),
    .D(net728),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[142][0] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _2362_ (.RESET_B(net358),
    .D(net866),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[142][1] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _2363_ (.RESET_B(net359),
    .D(net914),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[141][0] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _2364_ (.RESET_B(net360),
    .D(net927),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[141][1] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _2365_ (.RESET_B(net361),
    .D(net1066),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[140][0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2366_ (.RESET_B(net362),
    .D(net769),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[140][1] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _2367_ (.RESET_B(net363),
    .D(net1034),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[139][0] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _2368_ (.RESET_B(net364),
    .D(net946),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[139][1] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _2369_ (.RESET_B(net365),
    .D(net1004),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[138][0] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _2370_ (.RESET_B(net366),
    .D(net932),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[138][1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _2371_ (.RESET_B(net367),
    .D(net758),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[137][0] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _2372_ (.RESET_B(net368),
    .D(net781),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[137][1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _2373_ (.RESET_B(net369),
    .D(net1134),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[136][0] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _2374_ (.RESET_B(net370),
    .D(net999),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[136][1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _2375_ (.RESET_B(net371),
    .D(net987),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[135][0] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _2376_ (.RESET_B(net372),
    .D(net878),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[135][1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _2377_ (.RESET_B(net373),
    .D(net896),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[134][0] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _2378_ (.RESET_B(net374),
    .D(net873),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[134][1] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _2379_ (.RESET_B(net375),
    .D(net1046),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[133][0] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _2380_ (.RESET_B(net376),
    .D(net925),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[133][1] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _2381_ (.RESET_B(net377),
    .D(net785),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[132][0] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _2382_ (.RESET_B(net378),
    .D(net1024),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[132][1] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _2383_ (.RESET_B(net379),
    .D(net821),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[131][0] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _2384_ (.RESET_B(net380),
    .D(net822),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[131][1] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _2385_ (.RESET_B(net381),
    .D(net797),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[130][0] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _2386_ (.RESET_B(net382),
    .D(net805),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[130][1] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _2387_ (.RESET_B(net383),
    .D(net839),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[129][0] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _2388_ (.RESET_B(net384),
    .D(net871),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[129][1] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _2389_ (.RESET_B(net385),
    .D(net985),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[128][0] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _2390_ (.RESET_B(net386),
    .D(net976),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[128][1] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _2391_ (.RESET_B(net387),
    .D(net917),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[127][0] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _2392_ (.RESET_B(net388),
    .D(net867),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[127][1] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _2393_ (.RESET_B(net389),
    .D(net1010),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[126][0] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _2394_ (.RESET_B(net390),
    .D(net890),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[126][1] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _2395_ (.RESET_B(net391),
    .D(net791),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[125][0] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _2396_ (.RESET_B(net392),
    .D(net858),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[125][1] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _2397_ (.RESET_B(net393),
    .D(net735),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[124][0] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _2398_ (.RESET_B(net394),
    .D(net889),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[124][1] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _2399_ (.RESET_B(net395),
    .D(net893),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[123][0] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _2400_ (.RESET_B(net396),
    .D(net697),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[123][1] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _2401_ (.RESET_B(net397),
    .D(net741),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[122][0] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _2402_ (.RESET_B(net398),
    .D(net995),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[122][1] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _2403_ (.RESET_B(net399),
    .D(net970),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[121][0] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _2404_ (.RESET_B(net400),
    .D(net882),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[121][1] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _2405_ (.RESET_B(net401),
    .D(net851),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[120][0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2406_ (.RESET_B(net402),
    .D(net731),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[120][1] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _2407_ (.RESET_B(net403),
    .D(net856),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[119][0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2408_ (.RESET_B(net404),
    .D(net965),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[119][1] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _2409_ (.RESET_B(net405),
    .D(net740),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[118][0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2410_ (.RESET_B(net406),
    .D(net935),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[118][1] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _2411_ (.RESET_B(net407),
    .D(net1044),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[117][0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2412_ (.RESET_B(net408),
    .D(net713),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[117][1] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _2413_ (.RESET_B(net409),
    .D(net823),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[116][0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2414_ (.RESET_B(net410),
    .D(net930),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[116][1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _2415_ (.RESET_B(net411),
    .D(net844),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[115][0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2416_ (.RESET_B(net412),
    .D(net991),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[115][1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _2417_ (.RESET_B(net413),
    .D(net864),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[114][0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2418_ (.RESET_B(net414),
    .D(net887),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[114][1] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _2419_ (.RESET_B(net415),
    .D(net1133),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[113][0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2420_ (.RESET_B(net416),
    .D(net734),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[113][1] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _2421_ (.RESET_B(net417),
    .D(net1105),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[112][0] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _2422_ (.RESET_B(net418),
    .D(net916),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[112][1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _2423_ (.RESET_B(net419),
    .D(net700),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[111][0] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _2424_ (.RESET_B(net420),
    .D(net1022),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[111][1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _2425_ (.RESET_B(net421),
    .D(net950),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[110][0] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _2426_ (.RESET_B(net422),
    .D(net811),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[110][1] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2427_ (.RESET_B(net423),
    .D(net830),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[109][0] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _2428_ (.RESET_B(net424),
    .D(net892),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[109][1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _2429_ (.RESET_B(net425),
    .D(net857),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[108][0] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _2430_ (.RESET_B(net426),
    .D(net1116),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[108][1] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2431_ (.RESET_B(net427),
    .D(net1087),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[107][0] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _2432_ (.RESET_B(net428),
    .D(net1131),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[107][1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _2433_ (.RESET_B(net429),
    .D(net744),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[106][0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2434_ (.RESET_B(net430),
    .D(net773),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[106][1] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _2435_ (.RESET_B(net431),
    .D(net685),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[105][0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2436_ (.RESET_B(net432),
    .D(net846),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[105][1] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _2437_ (.RESET_B(net433),
    .D(net1049),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[104][0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2438_ (.RESET_B(net434),
    .D(net775),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[104][1] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _2439_ (.RESET_B(net435),
    .D(net694),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[103][0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2440_ (.RESET_B(net436),
    .D(net771),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[103][1] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _2441_ (.RESET_B(net437),
    .D(net712),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[102][0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2442_ (.RESET_B(net438),
    .D(net778),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[102][1] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _2443_ (.RESET_B(net439),
    .D(net695),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[101][0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2444_ (.RESET_B(net440),
    .D(net1125),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[101][1] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _2445_ (.RESET_B(net441),
    .D(net1009),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[100][0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2446_ (.RESET_B(net442),
    .D(net765),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[100][1] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _2447_ (.RESET_B(net443),
    .D(net702),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[99][0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2448_ (.RESET_B(net444),
    .D(net1005),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[99][1] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2449_ (.RESET_B(net445),
    .D(net1036),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[98][0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2450_ (.RESET_B(net446),
    .D(net1012),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[98][1] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2451_ (.RESET_B(net447),
    .D(net919),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[97][0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2452_ (.RESET_B(net448),
    .D(net958),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[97][1] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2453_ (.RESET_B(net449),
    .D(net1079),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[96][0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2454_ (.RESET_B(net450),
    .D(net1018),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[96][1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2455_ (.RESET_B(net451),
    .D(net1062),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[95][0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2456_ (.RESET_B(net452),
    .D(net1110),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[95][1] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2457_ (.RESET_B(net453),
    .D(net690),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[94][0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2458_ (.RESET_B(net454),
    .D(net727),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[94][1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2459_ (.RESET_B(net455),
    .D(net967),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[93][0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2460_ (.RESET_B(net456),
    .D(net1127),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[93][1] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2461_ (.RESET_B(net457),
    .D(net729),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[92][0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2462_ (.RESET_B(net458),
    .D(net748),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[92][1] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2463_ (.RESET_B(net459),
    .D(net1092),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[91][0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2464_ (.RESET_B(net460),
    .D(net964),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[91][1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2465_ (.RESET_B(net461),
    .D(net940),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[90][0] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2466_ (.RESET_B(net462),
    .D(net1064),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[90][1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2467_ (.RESET_B(net463),
    .D(net796),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[89][0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2468_ (.RESET_B(net464),
    .D(net1120),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[89][1] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2469_ (.RESET_B(net465),
    .D(net1118),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[88][0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2470_ (.RESET_B(net466),
    .D(net1035),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[88][1] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2471_ (.RESET_B(net467),
    .D(net923),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[87][0] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2472_ (.RESET_B(net468),
    .D(net688),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[87][1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2473_ (.RESET_B(net469),
    .D(net786),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[86][0] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2474_ (.RESET_B(net470),
    .D(net750),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[86][1] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2475_ (.RESET_B(net471),
    .D(net859),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[85][0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2476_ (.RESET_B(net472),
    .D(net1025),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[85][1] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2477_ (.RESET_B(net473),
    .D(net1050),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[84][0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2478_ (.RESET_B(net474),
    .D(net767),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[84][1] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2479_ (.RESET_B(net475),
    .D(net907),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[83][0] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2480_ (.RESET_B(net476),
    .D(net1042),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[83][1] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2481_ (.RESET_B(net477),
    .D(net841),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[82][0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2482_ (.RESET_B(net478),
    .D(net1071),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[82][1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2483_ (.RESET_B(net479),
    .D(net800),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[81][0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2484_ (.RESET_B(net480),
    .D(net1030),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[81][1] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2485_ (.RESET_B(net481),
    .D(net911),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[80][0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2486_ (.RESET_B(net482),
    .D(net1075),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[80][1] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2487_ (.RESET_B(net483),
    .D(net1057),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[79][0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2488_ (.RESET_B(net484),
    .D(net721),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[79][1] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2489_ (.RESET_B(net485),
    .D(net724),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[78][0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2490_ (.RESET_B(net486),
    .D(net921),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[78][1] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2491_ (.RESET_B(net487),
    .D(net989),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[77][0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2492_ (.RESET_B(net488),
    .D(net957),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[77][1] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2493_ (.RESET_B(net489),
    .D(net689),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[76][0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2494_ (.RESET_B(net490),
    .D(net931),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[76][1] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2495_ (.RESET_B(net491),
    .D(net1104),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[75][0] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2496_ (.RESET_B(net492),
    .D(net723),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[75][1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2497_ (.RESET_B(net493),
    .D(net761),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[74][0] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2498_ (.RESET_B(net494),
    .D(net827),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[74][1] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2499_ (.RESET_B(net495),
    .D(net813),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[73][0] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2500_ (.RESET_B(net496),
    .D(net1094),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[73][1] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2501_ (.RESET_B(net497),
    .D(net709),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[72][0] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2502_ (.RESET_B(net498),
    .D(net910),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[72][1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2503_ (.RESET_B(net499),
    .D(net746),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[71][0] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2504_ (.RESET_B(net500),
    .D(net863),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[71][1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2505_ (.RESET_B(net501),
    .D(net719),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[70][0] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2506_ (.RESET_B(net502),
    .D(net974),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[70][1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2507_ (.RESET_B(net503),
    .D(net1112),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[69][0] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2508_ (.RESET_B(net504),
    .D(net792),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[69][1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2509_ (.RESET_B(net505),
    .D(net1086),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[68][0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2510_ (.RESET_B(net506),
    .D(net1067),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[68][1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2511_ (.RESET_B(net507),
    .D(net831),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[67][0] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2512_ (.RESET_B(net508),
    .D(net883),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[67][1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2513_ (.RESET_B(net509),
    .D(net1011),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[66][0] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2514_ (.RESET_B(net510),
    .D(net706),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[66][1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2515_ (.RESET_B(net511),
    .D(net1095),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[65][0] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2516_ (.RESET_B(net512),
    .D(net793),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[65][1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2517_ (.RESET_B(net513),
    .D(net954),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[64][0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2518_ (.RESET_B(net514),
    .D(net1045),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[64][1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2519_ (.RESET_B(net515),
    .D(net815),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[63][0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2520_ (.RESET_B(net516),
    .D(net829),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[63][1] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2521_ (.RESET_B(net517),
    .D(net990),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[62][0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2522_ (.RESET_B(net518),
    .D(net1108),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[62][1] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2523_ (.RESET_B(net519),
    .D(net918),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[61][0] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2524_ (.RESET_B(net520),
    .D(net784),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[61][1] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2525_ (.RESET_B(net521),
    .D(net1015),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[60][0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2526_ (.RESET_B(net522),
    .D(net722),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[60][1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2527_ (.RESET_B(net523),
    .D(net835),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[59][0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _2528_ (.RESET_B(net524),
    .D(net711),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[59][1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2529_ (.RESET_B(net525),
    .D(net1073),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[58][0] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2530_ (.RESET_B(net526),
    .D(net766),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[58][1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2531_ (.RESET_B(net527),
    .D(net850),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[57][0] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2532_ (.RESET_B(net528),
    .D(net1078),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[57][1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2533_ (.RESET_B(net529),
    .D(net973),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[56][0] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2534_ (.RESET_B(net530),
    .D(net717),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[56][1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2535_ (.RESET_B(net531),
    .D(net1099),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[55][0] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2536_ (.RESET_B(net532),
    .D(net720),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[55][1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2537_ (.RESET_B(net533),
    .D(net733),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[54][0] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _2538_ (.RESET_B(net534),
    .D(net1027),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[54][1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2539_ (.RESET_B(net535),
    .D(net795),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[53][0] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2540_ (.RESET_B(net536),
    .D(net978),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[53][1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2541_ (.RESET_B(net537),
    .D(net1082),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[52][0] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2542_ (.RESET_B(net538),
    .D(net696),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[52][1] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _2543_ (.RESET_B(net539),
    .D(net1129),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[51][0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2544_ (.RESET_B(net540),
    .D(net845),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[51][1] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _2545_ (.RESET_B(net541),
    .D(net1077),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[50][0] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2546_ (.RESET_B(net542),
    .D(net1084),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[50][1] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _2547_ (.RESET_B(net543),
    .D(net1007),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[49][0] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2548_ (.RESET_B(net544),
    .D(net838),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[49][1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2549_ (.RESET_B(net545),
    .D(net874),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[48][0] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2550_ (.RESET_B(net546),
    .D(net808),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[48][1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2551_ (.RESET_B(net547),
    .D(net960),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[47][0] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _2552_ (.RESET_B(net548),
    .D(net814),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[47][1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2553_ (.RESET_B(net549),
    .D(net673),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[46][0] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _2554_ (.RESET_B(net550),
    .D(net1103),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[46][1] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _2555_ (.RESET_B(net551),
    .D(net993),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[45][0] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _2556_ (.RESET_B(net552),
    .D(net941),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[45][1] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _2557_ (.RESET_B(net553),
    .D(net710),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[44][0] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _2558_ (.RESET_B(net554),
    .D(net768),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[44][1] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2559_ (.RESET_B(net555),
    .D(net1006),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[43][0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _2560_ (.RESET_B(net556),
    .D(net1013),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[43][1] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2561_ (.RESET_B(net557),
    .D(net1069),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[42][0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _2562_ (.RESET_B(net558),
    .D(net969),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[42][1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2563_ (.RESET_B(net559),
    .D(net725),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[41][0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _2564_ (.RESET_B(net560),
    .D(net975),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[41][1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2565_ (.RESET_B(net561),
    .D(net939),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[40][0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _2566_ (.RESET_B(net562),
    .D(net743),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[40][1] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _2567_ (.RESET_B(net563),
    .D(net1048),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[39][0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _2568_ (.RESET_B(net564),
    .D(net849),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[39][1] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _2569_ (.RESET_B(net565),
    .D(net877),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[38][0] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2570_ (.RESET_B(net566),
    .D(net691),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[38][1] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _2571_ (.RESET_B(net567),
    .D(net899),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[37][0] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2572_ (.RESET_B(net568),
    .D(net1107),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[37][1] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _2573_ (.RESET_B(net569),
    .D(net745),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[36][0] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2574_ (.RESET_B(net570),
    .D(net1047),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[36][1] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _2575_ (.RESET_B(net571),
    .D(net888),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[35][0] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2576_ (.RESET_B(net572),
    .D(net1055),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[35][1] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2577_ (.RESET_B(net573),
    .D(net812),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[34][0] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2578_ (.RESET_B(net574),
    .D(net981),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[34][1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2579_ (.RESET_B(net575),
    .D(net902),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[33][0] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2580_ (.RESET_B(net576),
    .D(net681),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[33][1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2581_ (.RESET_B(net577),
    .D(net757),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[32][0] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2582_ (.RESET_B(net578),
    .D(net1101),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[32][1] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2583_ (.RESET_B(net579),
    .D(net1106),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[31][0] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2584_ (.RESET_B(net580),
    .D(net776),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[31][1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2585_ (.RESET_B(net581),
    .D(net833),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[30][0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2586_ (.RESET_B(net582),
    .D(net953),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[30][1] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2587_ (.RESET_B(net583),
    .D(net783),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[29][0] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2588_ (.RESET_B(net584),
    .D(net906),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[29][1] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _2589_ (.RESET_B(net585),
    .D(net988),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[28][0] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2590_ (.RESET_B(net586),
    .D(net1085),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[28][1] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _2591_ (.RESET_B(net587),
    .D(net1052),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[27][0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2592_ (.RESET_B(net588),
    .D(net1014),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[27][1] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _2593_ (.RESET_B(net589),
    .D(net818),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[26][0] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2594_ (.RESET_B(net590),
    .D(net809),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[26][1] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _2595_ (.RESET_B(net591),
    .D(net984),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[25][0] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2596_ (.RESET_B(net592),
    .D(net948),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[25][1] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _2597_ (.RESET_B(net593),
    .D(net1113),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[24][0] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2598_ (.RESET_B(net594),
    .D(net678),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[24][1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _2599_ (.RESET_B(net595),
    .D(net994),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[23][0] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2600_ (.RESET_B(net596),
    .D(net943),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[23][1] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _2601_ (.RESET_B(net597),
    .D(net749),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[22][0] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2602_ (.RESET_B(net598),
    .D(net755),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[22][1] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _2603_ (.RESET_B(net599),
    .D(net826),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[21][0] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2604_ (.RESET_B(net600),
    .D(net1100),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[21][1] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _2605_ (.RESET_B(net601),
    .D(net1002),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[20][0] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2606_ (.RESET_B(net602),
    .D(net1119),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[20][1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2607_ (.RESET_B(net603),
    .D(net1115),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[19][0] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2608_ (.RESET_B(net604),
    .D(net732),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[19][1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _2609_ (.RESET_B(net605),
    .D(net968),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[18][0] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2610_ (.RESET_B(net606),
    .D(net680),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[18][1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _2611_ (.RESET_B(net607),
    .D(net686),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[17][0] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2612_ (.RESET_B(net608),
    .D(net1063),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[17][1] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _2613_ (.RESET_B(net609),
    .D(net806),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[16][0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2614_ (.RESET_B(net610),
    .D(net701),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[16][1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _2615_ (.RESET_B(net611),
    .D(net951),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[15][0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2616_ (.RESET_B(net612),
    .D(net1043),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[15][1] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _2617_ (.RESET_B(net613),
    .D(net842),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[14][0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2618_ (.RESET_B(net614),
    .D(net677),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[14][1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _2619_ (.RESET_B(net615),
    .D(net894),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[13][0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2620_ (.RESET_B(net616),
    .D(net1068),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[13][1] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _2621_ (.RESET_B(net617),
    .D(net759),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[12][0] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2622_ (.RESET_B(net618),
    .D(net1121),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[12][1] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _2623_ (.RESET_B(net619),
    .D(net959),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[11][0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2624_ (.RESET_B(net620),
    .D(net922),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[11][1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2625_ (.RESET_B(net621),
    .D(net926),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[10][0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2626_ (.RESET_B(net622),
    .D(net810),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[10][1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2627_ (.RESET_B(net623),
    .D(net754),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[9][0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2628_ (.RESET_B(net624),
    .D(net852),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[9][1] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _2629_ (.RESET_B(net625),
    .D(net861),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[8][0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2630_ (.RESET_B(net626),
    .D(net897),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[8][1] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _2631_ (.RESET_B(net627),
    .D(net860),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[7][0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2632_ (.RESET_B(net628),
    .D(net872),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[7][1] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _2633_ (.RESET_B(net629),
    .D(net1091),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[6][0] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2634_ (.RESET_B(net630),
    .D(net875),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[6][1] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _2635_ (.RESET_B(net631),
    .D(net1051),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[5][0] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2636_ (.RESET_B(net632),
    .D(net1019),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[5][1] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _2637_ (.RESET_B(net633),
    .D(net962),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[4][0] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2638_ (.RESET_B(net634),
    .D(net687),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[4][1] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _2639_ (.RESET_B(net635),
    .D(net881),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[3][0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2640_ (.RESET_B(net636),
    .D(net1088),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[3][1] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _2641_ (.RESET_B(net637),
    .D(net908),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[2][0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2642_ (.RESET_B(net638),
    .D(net855),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[2][1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2643_ (.RESET_B(net655),
    .D(net1135),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[1][0] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2644_ (.RESET_B(net40),
    .D(net1139),
    .Q(\game_inst.snake_inst.shiftreg_inst.memory[1][1] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _2645_ (.RESET_B(net38),
    .D(_0110_),
    .Q(\game_inst.snake_inst.pos[1] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _2646_ (.RESET_B(net36),
    .D(net1261),
    .Q(\game_inst.snake_inst.pos[2] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _2647_ (.RESET_B(net34),
    .D(net1170),
    .Q(\game_inst.snake_inst.pos[4] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _2648_ (.RESET_B(net32),
    .D(_0113_),
    .Q(\game_inst.vga_inst.row_buffer[1][0] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _2649_ (.RESET_B(net30),
    .D(_0114_),
    .Q(\game_inst.vga_inst.row_buffer[1][1] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _2650_ (.RESET_B(net22),
    .D(_0115_),
    .Q(\game_inst.vga_inst.row_buffer[11][0] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2651_ (.RESET_B(net20),
    .D(_0116_),
    .Q(\game_inst.vga_inst.row_buffer[11][1] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _2652_ (.RESET_B(net18),
    .D(_0117_),
    .Q(\game_inst.apple_inst.apple_y[0] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _2653_ (.RESET_B(net666),
    .D(_0118_),
    .Q(\game_inst.apple_inst.apple_y[1] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _2654_ (.RESET_B(net664),
    .D(net1214),
    .Q(\game_inst.apple_inst.apple_y[2] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _2655_ (.RESET_B(net662),
    .D(_0120_),
    .Q(\game_inst.apple_inst.apple_y[3] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _2656_ (.RESET_B(net660),
    .D(net1172),
    .Q(\game_inst.control_inst.o_start ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _2657_ (.RESET_B(net658),
    .D(_0122_),
    .Q(\game_inst.vga_inst.row_buffer[16][0] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2658_ (.RESET_B(net654),
    .D(_0123_),
    .Q(\game_inst.vga_inst.row_buffer[16][1] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _2659_ (.RESET_B(net652),
    .D(net1270),
    .Q(\game_inst.colorblind ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _2660_ (.RESET_B(net656),
    .D(net1149),
    .Q(\game_inst.tick ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _2661_ (.RESET_B(net156),
    .D(\game_inst.tickgen_inst.i_vsync ),
    .Q(\game_inst.tickgen_inst.prev_vsync ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _2662_ (.RESET_B(net640),
    .D(_0000_),
    .Q(\game_inst.tickgen_inst.prev_user_input ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _2663_ (.RESET_B(net170),
    .D(net1286),
    .Q(\game_inst.tickgen_inst.counter_max[0] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _2664_ (.RESET_B(net166),
    .D(net1282),
    .Q(\game_inst.tickgen_inst.counter_max[1] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _2665_ (.RESET_B(net162),
    .D(_0128_),
    .Q(\game_inst.tickgen_inst.counter_max[2] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _2666_ (.RESET_B(net158),
    .D(_0129_),
    .Q(\game_inst.tickgen_inst.counter_max[3] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _2667_ (.RESET_B(net154),
    .D(net1145),
    .Q(\game_inst.tickgen_inst.counter_max[4] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _2668_ (.RESET_B(net650),
    .D(net1256),
    .Q(\game_inst.tickgen_inst.counter[0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2669_ (.RESET_B(net168),
    .D(net1253),
    .Q(\game_inst.tickgen_inst.counter[1] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _2670_ (.RESET_B(net160),
    .D(_0133_),
    .Q(\game_inst.tickgen_inst.counter[2] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _2671_ (.RESET_B(net145),
    .D(_0134_),
    .Q(\game_inst.tickgen_inst.counter[3] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _2672_ (.RESET_B(net164),
    .D(net1311),
    .Q(\game_inst.tickgen_inst.counter[4] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _2673_ (.RESET_B(net172),
    .D(net1258),
    .Q(failure),
    .CLK(clknet_leaf_33_clk));
 sg13g2_tiehi _2131__19 (.L_HI(net19));
 sg13g2_tiehi _2651__20 (.L_HI(net20));
 sg13g2_tiehi _2130__21 (.L_HI(net21));
 sg13g2_tiehi _2650__22 (.L_HI(net22));
 sg13g2_tiehi _2129__23 (.L_HI(net23));
 sg13g2_tiehi _2128__24 (.L_HI(net24));
 sg13g2_tiehi _2127__25 (.L_HI(net25));
 sg13g2_tiehi _2126__26 (.L_HI(net26));
 sg13g2_tiehi _2125__27 (.L_HI(net27));
 sg13g2_tiehi _2124__28 (.L_HI(net28));
 sg13g2_tiehi _2123__29 (.L_HI(net29));
 sg13g2_tiehi _2649__30 (.L_HI(net30));
 sg13g2_tiehi _2122__31 (.L_HI(net31));
 sg13g2_tiehi _2648__32 (.L_HI(net32));
 sg13g2_tiehi _2120__33 (.L_HI(net33));
 sg13g2_tiehi _2647__34 (.L_HI(net34));
 sg13g2_tiehi _2119__35 (.L_HI(net35));
 sg13g2_tiehi _2646__36 (.L_HI(net36));
 sg13g2_tiehi _2118__37 (.L_HI(net37));
 sg13g2_tiehi _2645__38 (.L_HI(net38));
 sg13g2_tiehi _2117__39 (.L_HI(net39));
 sg13g2_tiehi _2644__40 (.L_HI(net40));
 sg13g2_tiehi _2116__41 (.L_HI(net41));
 sg13g2_tiehi _2177__42 (.L_HI(net42));
 sg13g2_tiehi _2115__43 (.L_HI(net43));
 sg13g2_tiehi _2176__44 (.L_HI(net44));
 sg13g2_tiehi _2114__45 (.L_HI(net45));
 sg13g2_tiehi _2175__46 (.L_HI(net46));
 sg13g2_tiehi _2113__47 (.L_HI(net47));
 sg13g2_tiehi _2174__48 (.L_HI(net48));
 sg13g2_tiehi _2112__49 (.L_HI(net49));
 sg13g2_tiehi _2111__50 (.L_HI(net50));
 sg13g2_tiehi _2109__51 (.L_HI(net51));
 sg13g2_tiehi _2108__52 (.L_HI(net52));
 sg13g2_tiehi _2107__53 (.L_HI(net53));
 sg13g2_tiehi _2106__54 (.L_HI(net54));
 sg13g2_tiehi _2105__55 (.L_HI(net55));
 sg13g2_tiehi _2104__56 (.L_HI(net56));
 sg13g2_tiehi _2103__57 (.L_HI(net57));
 sg13g2_tiehi _2102__58 (.L_HI(net58));
 sg13g2_tiehi _2070__59 (.L_HI(net59));
 sg13g2_tiehi _2101__60 (.L_HI(net60));
 sg13g2_tiehi _2100__61 (.L_HI(net61));
 sg13g2_tiehi _2099__62 (.L_HI(net62));
 sg13g2_tiehi _2098__63 (.L_HI(net63));
 sg13g2_tiehi _2097__64 (.L_HI(net64));
 sg13g2_tiehi _2096__65 (.L_HI(net65));
 sg13g2_tiehi _2095__66 (.L_HI(net66));
 sg13g2_tiehi _2094__67 (.L_HI(net67));
 sg13g2_tiehi _2093__68 (.L_HI(net68));
 sg13g2_tiehi _2092__69 (.L_HI(net69));
 sg13g2_tiehi _2110__70 (.L_HI(net70));
 sg13g2_tiehi _2091__71 (.L_HI(net71));
 sg13g2_tiehi _2090__72 (.L_HI(net72));
 sg13g2_tiehi _2089__73 (.L_HI(net73));
 sg13g2_tiehi _2088__74 (.L_HI(net74));
 sg13g2_tiehi _2087__75 (.L_HI(net75));
 sg13g2_tiehi _2086__76 (.L_HI(net76));
 sg13g2_tiehi _2085__77 (.L_HI(net77));
 sg13g2_tiehi _2084__78 (.L_HI(net78));
 sg13g2_tiehi _2083__79 (.L_HI(net79));
 sg13g2_tiehi _2082__80 (.L_HI(net80));
 sg13g2_tiehi _2081__81 (.L_HI(net81));
 sg13g2_tiehi _2080__82 (.L_HI(net82));
 sg13g2_tiehi _2079__83 (.L_HI(net83));
 sg13g2_tiehi _2078__84 (.L_HI(net84));
 sg13g2_tiehi _2077__85 (.L_HI(net85));
 sg13g2_tiehi _2076__86 (.L_HI(net86));
 sg13g2_tiehi _2075__87 (.L_HI(net87));
 sg13g2_tiehi _2074__88 (.L_HI(net88));
 sg13g2_tiehi _2073__89 (.L_HI(net89));
 sg13g2_tiehi _2072__90 (.L_HI(net90));
 sg13g2_tiehi _2071__91 (.L_HI(net91));
 sg13g2_tiehi _2173__92 (.L_HI(net92));
 sg13g2_tiehi _2172__93 (.L_HI(net93));
 sg13g2_tiehi _2171__94 (.L_HI(net140));
 sg13g2_tiehi _2170__95 (.L_HI(net141));
 sg13g2_tiehi _2169__96 (.L_HI(net142));
 sg13g2_tiehi _2168__97 (.L_HI(net143));
 sg13g2_tiehi _2167__98 (.L_HI(net144));
 sg13g2_tiehi _2671__99 (.L_HI(net145));
 sg13g2_tiehi _2166__100 (.L_HI(net146));
 sg13g2_tiehi _2165__101 (.L_HI(net147));
 sg13g2_tiehi _2164__102 (.L_HI(net148));
 sg13g2_tiehi _2163__103 (.L_HI(net149));
 sg13g2_tiehi _2162__104 (.L_HI(net150));
 sg13g2_tiehi _2161__105 (.L_HI(net151));
 sg13g2_tiehi _2160__106 (.L_HI(net152));
 sg13g2_tiehi _2159__107 (.L_HI(net153));
 sg13g2_tiehi _2667__108 (.L_HI(net154));
 sg13g2_tiehi _2158__109 (.L_HI(net155));
 sg13g2_tiehi _2661__110 (.L_HI(net156));
 sg13g2_tiehi _2157__111 (.L_HI(net157));
 sg13g2_tiehi _2666__112 (.L_HI(net158));
 sg13g2_tiehi _2156__113 (.L_HI(net159));
 sg13g2_tiehi _2670__114 (.L_HI(net160));
 sg13g2_tiehi _2155__115 (.L_HI(net161));
 sg13g2_tiehi _2665__116 (.L_HI(net162));
 sg13g2_tiehi _2154__117 (.L_HI(net163));
 sg13g2_tiehi _2672__118 (.L_HI(net164));
 sg13g2_tiehi _2153__119 (.L_HI(net165));
 sg13g2_tiehi _2664__120 (.L_HI(net166));
 sg13g2_tiehi _2152__121 (.L_HI(net167));
 sg13g2_tiehi _2669__122 (.L_HI(net168));
 sg13g2_tiehi _2151__123 (.L_HI(net169));
 sg13g2_tiehi _2663__124 (.L_HI(net170));
 sg13g2_tiehi _2150__125 (.L_HI(net171));
 sg13g2_tiehi _2673__126 (.L_HI(net172));
 sg13g2_tiehi _2121__127 (.L_HI(net173));
 sg13g2_tiehi _2178__128 (.L_HI(net174));
 sg13g2_tiehi _2179__129 (.L_HI(net175));
 sg13g2_tiehi _2180__130 (.L_HI(net176));
 sg13g2_tiehi _2181__131 (.L_HI(net177));
 sg13g2_tiehi _2182__132 (.L_HI(net178));
 sg13g2_tiehi _2183__133 (.L_HI(net179));
 sg13g2_tiehi _2184__134 (.L_HI(net180));
 sg13g2_tiehi _2185__135 (.L_HI(net181));
 sg13g2_tiehi _2186__136 (.L_HI(net182));
 sg13g2_tiehi _2187__137 (.L_HI(net183));
 sg13g2_tiehi _2188__138 (.L_HI(net184));
 sg13g2_tiehi _2189__139 (.L_HI(net185));
 sg13g2_tiehi _2190__140 (.L_HI(net186));
 sg13g2_tiehi _2191__141 (.L_HI(net187));
 sg13g2_tiehi _2192__142 (.L_HI(net188));
 sg13g2_tiehi _2193__143 (.L_HI(net189));
 sg13g2_tiehi _2194__144 (.L_HI(net190));
 sg13g2_tiehi _2195__145 (.L_HI(net191));
 sg13g2_tiehi _2196__146 (.L_HI(net192));
 sg13g2_tiehi _2197__147 (.L_HI(net193));
 sg13g2_tiehi _2198__148 (.L_HI(net194));
 sg13g2_tiehi _2199__149 (.L_HI(net195));
 sg13g2_tiehi _2200__150 (.L_HI(net196));
 sg13g2_tiehi _2201__151 (.L_HI(net197));
 sg13g2_tiehi _2202__152 (.L_HI(net198));
 sg13g2_tiehi _2203__153 (.L_HI(net199));
 sg13g2_tiehi _2204__154 (.L_HI(net200));
 sg13g2_tiehi _2205__155 (.L_HI(net201));
 sg13g2_tiehi _2206__156 (.L_HI(net202));
 sg13g2_tiehi _2207__157 (.L_HI(net203));
 sg13g2_tiehi _2208__158 (.L_HI(net204));
 sg13g2_tiehi _2209__159 (.L_HI(net205));
 sg13g2_tiehi _2210__160 (.L_HI(net206));
 sg13g2_tiehi _2211__161 (.L_HI(net207));
 sg13g2_tiehi _2212__162 (.L_HI(net208));
 sg13g2_tiehi _2213__163 (.L_HI(net209));
 sg13g2_tiehi _2214__164 (.L_HI(net210));
 sg13g2_tiehi _2215__165 (.L_HI(net211));
 sg13g2_tiehi _2216__166 (.L_HI(net212));
 sg13g2_tiehi _2217__167 (.L_HI(net213));
 sg13g2_tiehi _2218__168 (.L_HI(net214));
 sg13g2_tiehi _2219__169 (.L_HI(net215));
 sg13g2_tiehi _2220__170 (.L_HI(net216));
 sg13g2_tiehi _2221__171 (.L_HI(net217));
 sg13g2_tiehi _2222__172 (.L_HI(net218));
 sg13g2_tiehi _2223__173 (.L_HI(net219));
 sg13g2_tiehi _2224__174 (.L_HI(net220));
 sg13g2_tiehi _2225__175 (.L_HI(net221));
 sg13g2_tiehi _2226__176 (.L_HI(net222));
 sg13g2_tiehi _2227__177 (.L_HI(net223));
 sg13g2_tiehi _2228__178 (.L_HI(net224));
 sg13g2_tiehi _2229__179 (.L_HI(net225));
 sg13g2_tiehi _2230__180 (.L_HI(net226));
 sg13g2_tiehi _2231__181 (.L_HI(net227));
 sg13g2_tiehi _2232__182 (.L_HI(net228));
 sg13g2_tiehi _2233__183 (.L_HI(net229));
 sg13g2_tiehi _2234__184 (.L_HI(net230));
 sg13g2_tiehi _2235__185 (.L_HI(net231));
 sg13g2_tiehi _2236__186 (.L_HI(net232));
 sg13g2_tiehi _2237__187 (.L_HI(net233));
 sg13g2_tiehi _2238__188 (.L_HI(net234));
 sg13g2_tiehi _2239__189 (.L_HI(net235));
 sg13g2_tiehi _2240__190 (.L_HI(net236));
 sg13g2_tiehi _2241__191 (.L_HI(net237));
 sg13g2_tiehi _2242__192 (.L_HI(net238));
 sg13g2_tiehi _2243__193 (.L_HI(net239));
 sg13g2_tiehi _2244__194 (.L_HI(net240));
 sg13g2_tiehi _2245__195 (.L_HI(net241));
 sg13g2_tiehi _2246__196 (.L_HI(net242));
 sg13g2_tiehi _2247__197 (.L_HI(net243));
 sg13g2_tiehi _2248__198 (.L_HI(net244));
 sg13g2_tiehi _2249__199 (.L_HI(net245));
 sg13g2_tiehi _2250__200 (.L_HI(net246));
 sg13g2_tiehi _2251__201 (.L_HI(net247));
 sg13g2_tiehi _2252__202 (.L_HI(net248));
 sg13g2_tiehi _2253__203 (.L_HI(net249));
 sg13g2_tiehi _2254__204 (.L_HI(net250));
 sg13g2_tiehi _2255__205 (.L_HI(net251));
 sg13g2_tiehi _2256__206 (.L_HI(net252));
 sg13g2_tiehi _2257__207 (.L_HI(net253));
 sg13g2_tiehi _2258__208 (.L_HI(net254));
 sg13g2_tiehi _2259__209 (.L_HI(net255));
 sg13g2_tiehi _2260__210 (.L_HI(net256));
 sg13g2_tiehi _2261__211 (.L_HI(net257));
 sg13g2_tiehi _2262__212 (.L_HI(net258));
 sg13g2_tiehi _2263__213 (.L_HI(net259));
 sg13g2_tiehi _2264__214 (.L_HI(net260));
 sg13g2_tiehi _2265__215 (.L_HI(net261));
 sg13g2_tiehi _2266__216 (.L_HI(net262));
 sg13g2_tiehi _2267__217 (.L_HI(net263));
 sg13g2_tiehi _2268__218 (.L_HI(net264));
 sg13g2_tiehi _2269__219 (.L_HI(net265));
 sg13g2_tiehi _2270__220 (.L_HI(net266));
 sg13g2_tiehi _2271__221 (.L_HI(net267));
 sg13g2_tiehi _2272__222 (.L_HI(net268));
 sg13g2_tiehi _2273__223 (.L_HI(net269));
 sg13g2_tiehi _2274__224 (.L_HI(net270));
 sg13g2_tiehi _2275__225 (.L_HI(net271));
 sg13g2_tiehi _2276__226 (.L_HI(net272));
 sg13g2_tiehi _2277__227 (.L_HI(net273));
 sg13g2_tiehi _2278__228 (.L_HI(net274));
 sg13g2_tiehi _2279__229 (.L_HI(net275));
 sg13g2_tiehi _2280__230 (.L_HI(net276));
 sg13g2_tiehi _2281__231 (.L_HI(net277));
 sg13g2_tiehi _2282__232 (.L_HI(net278));
 sg13g2_tiehi _2283__233 (.L_HI(net279));
 sg13g2_tiehi _2284__234 (.L_HI(net280));
 sg13g2_tiehi _2285__235 (.L_HI(net281));
 sg13g2_tiehi _2286__236 (.L_HI(net282));
 sg13g2_tiehi _2287__237 (.L_HI(net283));
 sg13g2_tiehi _2288__238 (.L_HI(net284));
 sg13g2_tiehi _2289__239 (.L_HI(net285));
 sg13g2_tiehi _2290__240 (.L_HI(net286));
 sg13g2_tiehi _2291__241 (.L_HI(net287));
 sg13g2_tiehi _2292__242 (.L_HI(net288));
 sg13g2_tiehi _2293__243 (.L_HI(net289));
 sg13g2_tiehi _2294__244 (.L_HI(net290));
 sg13g2_tiehi _2295__245 (.L_HI(net291));
 sg13g2_tiehi _2296__246 (.L_HI(net292));
 sg13g2_tiehi _2297__247 (.L_HI(net293));
 sg13g2_tiehi _2298__248 (.L_HI(net294));
 sg13g2_tiehi _2299__249 (.L_HI(net295));
 sg13g2_tiehi _2300__250 (.L_HI(net296));
 sg13g2_tiehi _2301__251 (.L_HI(net297));
 sg13g2_tiehi _2302__252 (.L_HI(net298));
 sg13g2_tiehi _2303__253 (.L_HI(net299));
 sg13g2_tiehi _2304__254 (.L_HI(net300));
 sg13g2_tiehi _2305__255 (.L_HI(net301));
 sg13g2_tiehi _2306__256 (.L_HI(net302));
 sg13g2_tiehi _2307__257 (.L_HI(net303));
 sg13g2_tiehi _2308__258 (.L_HI(net304));
 sg13g2_tiehi _2309__259 (.L_HI(net305));
 sg13g2_tiehi _2310__260 (.L_HI(net306));
 sg13g2_tiehi _2311__261 (.L_HI(net307));
 sg13g2_tiehi _2312__262 (.L_HI(net308));
 sg13g2_tiehi _2313__263 (.L_HI(net309));
 sg13g2_tiehi _2314__264 (.L_HI(net310));
 sg13g2_tiehi _2315__265 (.L_HI(net311));
 sg13g2_tiehi _2316__266 (.L_HI(net312));
 sg13g2_tiehi _2317__267 (.L_HI(net313));
 sg13g2_tiehi _2318__268 (.L_HI(net314));
 sg13g2_tiehi _2319__269 (.L_HI(net315));
 sg13g2_tiehi _2320__270 (.L_HI(net316));
 sg13g2_tiehi _2321__271 (.L_HI(net317));
 sg13g2_tiehi _2322__272 (.L_HI(net318));
 sg13g2_tiehi _2323__273 (.L_HI(net319));
 sg13g2_tiehi _2324__274 (.L_HI(net320));
 sg13g2_tiehi _2325__275 (.L_HI(net321));
 sg13g2_tiehi _2326__276 (.L_HI(net322));
 sg13g2_tiehi _2327__277 (.L_HI(net323));
 sg13g2_tiehi _2328__278 (.L_HI(net324));
 sg13g2_tiehi _2329__279 (.L_HI(net325));
 sg13g2_tiehi _2330__280 (.L_HI(net326));
 sg13g2_tiehi _2331__281 (.L_HI(net327));
 sg13g2_tiehi _2332__282 (.L_HI(net328));
 sg13g2_tiehi _2333__283 (.L_HI(net329));
 sg13g2_tiehi _2334__284 (.L_HI(net330));
 sg13g2_tiehi _2335__285 (.L_HI(net331));
 sg13g2_tiehi _2336__286 (.L_HI(net332));
 sg13g2_tiehi _2337__287 (.L_HI(net333));
 sg13g2_tiehi _2338__288 (.L_HI(net334));
 sg13g2_tiehi _2339__289 (.L_HI(net335));
 sg13g2_tiehi _2340__290 (.L_HI(net336));
 sg13g2_tiehi _2341__291 (.L_HI(net337));
 sg13g2_tiehi _2342__292 (.L_HI(net338));
 sg13g2_tiehi _2343__293 (.L_HI(net339));
 sg13g2_tiehi _2344__294 (.L_HI(net340));
 sg13g2_tiehi _2345__295 (.L_HI(net341));
 sg13g2_tiehi _2346__296 (.L_HI(net342));
 sg13g2_tiehi _2347__297 (.L_HI(net343));
 sg13g2_tiehi _2348__298 (.L_HI(net344));
 sg13g2_tiehi _2349__299 (.L_HI(net345));
 sg13g2_tiehi _2350__300 (.L_HI(net346));
 sg13g2_tiehi _2351__301 (.L_HI(net347));
 sg13g2_tiehi _2352__302 (.L_HI(net348));
 sg13g2_tiehi _2353__303 (.L_HI(net349));
 sg13g2_tiehi _2354__304 (.L_HI(net350));
 sg13g2_tiehi _2355__305 (.L_HI(net351));
 sg13g2_tiehi _2356__306 (.L_HI(net352));
 sg13g2_tiehi _2357__307 (.L_HI(net353));
 sg13g2_tiehi _2358__308 (.L_HI(net354));
 sg13g2_tiehi _2359__309 (.L_HI(net355));
 sg13g2_tiehi _2360__310 (.L_HI(net356));
 sg13g2_tiehi _2361__311 (.L_HI(net357));
 sg13g2_tiehi _2362__312 (.L_HI(net358));
 sg13g2_tiehi _2363__313 (.L_HI(net359));
 sg13g2_tiehi _2364__314 (.L_HI(net360));
 sg13g2_tiehi _2365__315 (.L_HI(net361));
 sg13g2_tiehi _2366__316 (.L_HI(net362));
 sg13g2_tiehi _2367__317 (.L_HI(net363));
 sg13g2_tiehi _2368__318 (.L_HI(net364));
 sg13g2_tiehi _2369__319 (.L_HI(net365));
 sg13g2_tiehi _2370__320 (.L_HI(net366));
 sg13g2_tiehi _2371__321 (.L_HI(net367));
 sg13g2_tiehi _2372__322 (.L_HI(net368));
 sg13g2_tiehi _2373__323 (.L_HI(net369));
 sg13g2_tiehi _2374__324 (.L_HI(net370));
 sg13g2_tiehi _2375__325 (.L_HI(net371));
 sg13g2_tiehi _2376__326 (.L_HI(net372));
 sg13g2_tiehi _2377__327 (.L_HI(net373));
 sg13g2_tiehi _2378__328 (.L_HI(net374));
 sg13g2_tiehi _2379__329 (.L_HI(net375));
 sg13g2_tiehi _2380__330 (.L_HI(net376));
 sg13g2_tiehi _2381__331 (.L_HI(net377));
 sg13g2_tiehi _2382__332 (.L_HI(net378));
 sg13g2_tiehi _2383__333 (.L_HI(net379));
 sg13g2_tiehi _2384__334 (.L_HI(net380));
 sg13g2_tiehi _2385__335 (.L_HI(net381));
 sg13g2_tiehi _2386__336 (.L_HI(net382));
 sg13g2_tiehi _2387__337 (.L_HI(net383));
 sg13g2_tiehi _2388__338 (.L_HI(net384));
 sg13g2_tiehi _2389__339 (.L_HI(net385));
 sg13g2_tiehi _2390__340 (.L_HI(net386));
 sg13g2_tiehi _2391__341 (.L_HI(net387));
 sg13g2_tiehi _2392__342 (.L_HI(net388));
 sg13g2_tiehi _2393__343 (.L_HI(net389));
 sg13g2_tiehi _2394__344 (.L_HI(net390));
 sg13g2_tiehi _2395__345 (.L_HI(net391));
 sg13g2_tiehi _2396__346 (.L_HI(net392));
 sg13g2_tiehi _2397__347 (.L_HI(net393));
 sg13g2_tiehi _2398__348 (.L_HI(net394));
 sg13g2_tiehi _2399__349 (.L_HI(net395));
 sg13g2_tiehi _2400__350 (.L_HI(net396));
 sg13g2_tiehi _2401__351 (.L_HI(net397));
 sg13g2_tiehi _2402__352 (.L_HI(net398));
 sg13g2_tiehi _2403__353 (.L_HI(net399));
 sg13g2_tiehi _2404__354 (.L_HI(net400));
 sg13g2_tiehi _2405__355 (.L_HI(net401));
 sg13g2_tiehi _2406__356 (.L_HI(net402));
 sg13g2_tiehi _2407__357 (.L_HI(net403));
 sg13g2_tiehi _2408__358 (.L_HI(net404));
 sg13g2_tiehi _2409__359 (.L_HI(net405));
 sg13g2_tiehi _2410__360 (.L_HI(net406));
 sg13g2_tiehi _2411__361 (.L_HI(net407));
 sg13g2_tiehi _2412__362 (.L_HI(net408));
 sg13g2_tiehi _2413__363 (.L_HI(net409));
 sg13g2_tiehi _2414__364 (.L_HI(net410));
 sg13g2_tiehi _2415__365 (.L_HI(net411));
 sg13g2_tiehi _2416__366 (.L_HI(net412));
 sg13g2_tiehi _2417__367 (.L_HI(net413));
 sg13g2_tiehi _2418__368 (.L_HI(net414));
 sg13g2_tiehi _2419__369 (.L_HI(net415));
 sg13g2_tiehi _2420__370 (.L_HI(net416));
 sg13g2_tiehi _2421__371 (.L_HI(net417));
 sg13g2_tiehi _2422__372 (.L_HI(net418));
 sg13g2_tiehi _2423__373 (.L_HI(net419));
 sg13g2_tiehi _2424__374 (.L_HI(net420));
 sg13g2_tiehi _2425__375 (.L_HI(net421));
 sg13g2_tiehi _2426__376 (.L_HI(net422));
 sg13g2_tiehi _2427__377 (.L_HI(net423));
 sg13g2_tiehi _2428__378 (.L_HI(net424));
 sg13g2_tiehi _2429__379 (.L_HI(net425));
 sg13g2_tiehi _2430__380 (.L_HI(net426));
 sg13g2_tiehi _2431__381 (.L_HI(net427));
 sg13g2_tiehi _2432__382 (.L_HI(net428));
 sg13g2_tiehi _2433__383 (.L_HI(net429));
 sg13g2_tiehi _2434__384 (.L_HI(net430));
 sg13g2_tiehi _2435__385 (.L_HI(net431));
 sg13g2_tiehi _2436__386 (.L_HI(net432));
 sg13g2_tiehi _2437__387 (.L_HI(net433));
 sg13g2_tiehi _2438__388 (.L_HI(net434));
 sg13g2_tiehi _2439__389 (.L_HI(net435));
 sg13g2_tiehi _2440__390 (.L_HI(net436));
 sg13g2_tiehi _2441__391 (.L_HI(net437));
 sg13g2_tiehi _2442__392 (.L_HI(net438));
 sg13g2_tiehi _2443__393 (.L_HI(net439));
 sg13g2_tiehi _2444__394 (.L_HI(net440));
 sg13g2_tiehi _2445__395 (.L_HI(net441));
 sg13g2_tiehi _2446__396 (.L_HI(net442));
 sg13g2_tiehi _2447__397 (.L_HI(net443));
 sg13g2_tiehi _2448__398 (.L_HI(net444));
 sg13g2_tiehi _2449__399 (.L_HI(net445));
 sg13g2_tiehi _2450__400 (.L_HI(net446));
 sg13g2_tiehi _2451__401 (.L_HI(net447));
 sg13g2_tiehi _2452__402 (.L_HI(net448));
 sg13g2_tiehi _2453__403 (.L_HI(net449));
 sg13g2_tiehi _2454__404 (.L_HI(net450));
 sg13g2_tiehi _2455__405 (.L_HI(net451));
 sg13g2_tiehi _2456__406 (.L_HI(net452));
 sg13g2_tiehi _2457__407 (.L_HI(net453));
 sg13g2_tiehi _2458__408 (.L_HI(net454));
 sg13g2_tiehi _2459__409 (.L_HI(net455));
 sg13g2_tiehi _2460__410 (.L_HI(net456));
 sg13g2_tiehi _2461__411 (.L_HI(net457));
 sg13g2_tiehi _2462__412 (.L_HI(net458));
 sg13g2_tiehi _2463__413 (.L_HI(net459));
 sg13g2_tiehi _2464__414 (.L_HI(net460));
 sg13g2_tiehi _2465__415 (.L_HI(net461));
 sg13g2_tiehi _2466__416 (.L_HI(net462));
 sg13g2_tiehi _2467__417 (.L_HI(net463));
 sg13g2_tiehi _2468__418 (.L_HI(net464));
 sg13g2_tiehi _2469__419 (.L_HI(net465));
 sg13g2_tiehi _2470__420 (.L_HI(net466));
 sg13g2_tiehi _2471__421 (.L_HI(net467));
 sg13g2_tiehi _2472__422 (.L_HI(net468));
 sg13g2_tiehi _2473__423 (.L_HI(net469));
 sg13g2_tiehi _2474__424 (.L_HI(net470));
 sg13g2_tiehi _2475__425 (.L_HI(net471));
 sg13g2_tiehi _2476__426 (.L_HI(net472));
 sg13g2_tiehi _2477__427 (.L_HI(net473));
 sg13g2_tiehi _2478__428 (.L_HI(net474));
 sg13g2_tiehi _2479__429 (.L_HI(net475));
 sg13g2_tiehi _2480__430 (.L_HI(net476));
 sg13g2_tiehi _2481__431 (.L_HI(net477));
 sg13g2_tiehi _2482__432 (.L_HI(net478));
 sg13g2_tiehi _2483__433 (.L_HI(net479));
 sg13g2_tiehi _2484__434 (.L_HI(net480));
 sg13g2_tiehi _2485__435 (.L_HI(net481));
 sg13g2_tiehi _2486__436 (.L_HI(net482));
 sg13g2_tiehi _2487__437 (.L_HI(net483));
 sg13g2_tiehi _2488__438 (.L_HI(net484));
 sg13g2_tiehi _2489__439 (.L_HI(net485));
 sg13g2_tiehi _2490__440 (.L_HI(net486));
 sg13g2_tiehi _2491__441 (.L_HI(net487));
 sg13g2_tiehi _2492__442 (.L_HI(net488));
 sg13g2_tiehi _2493__443 (.L_HI(net489));
 sg13g2_tiehi _2494__444 (.L_HI(net490));
 sg13g2_tiehi _2495__445 (.L_HI(net491));
 sg13g2_tiehi _2496__446 (.L_HI(net492));
 sg13g2_tiehi _2497__447 (.L_HI(net493));
 sg13g2_tiehi _2498__448 (.L_HI(net494));
 sg13g2_tiehi _2499__449 (.L_HI(net495));
 sg13g2_tiehi _2500__450 (.L_HI(net496));
 sg13g2_tiehi _2501__451 (.L_HI(net497));
 sg13g2_tiehi _2502__452 (.L_HI(net498));
 sg13g2_tiehi _2503__453 (.L_HI(net499));
 sg13g2_tiehi _2504__454 (.L_HI(net500));
 sg13g2_tiehi _2505__455 (.L_HI(net501));
 sg13g2_tiehi _2506__456 (.L_HI(net502));
 sg13g2_tiehi _2507__457 (.L_HI(net503));
 sg13g2_tiehi _2508__458 (.L_HI(net504));
 sg13g2_tiehi _2509__459 (.L_HI(net505));
 sg13g2_tiehi _2510__460 (.L_HI(net506));
 sg13g2_tiehi _2511__461 (.L_HI(net507));
 sg13g2_tiehi _2512__462 (.L_HI(net508));
 sg13g2_tiehi _2513__463 (.L_HI(net509));
 sg13g2_tiehi _2514__464 (.L_HI(net510));
 sg13g2_tiehi _2515__465 (.L_HI(net511));
 sg13g2_tiehi _2516__466 (.L_HI(net512));
 sg13g2_tiehi _2517__467 (.L_HI(net513));
 sg13g2_tiehi _2518__468 (.L_HI(net514));
 sg13g2_tiehi _2519__469 (.L_HI(net515));
 sg13g2_tiehi _2520__470 (.L_HI(net516));
 sg13g2_tiehi _2521__471 (.L_HI(net517));
 sg13g2_tiehi _2522__472 (.L_HI(net518));
 sg13g2_tiehi _2523__473 (.L_HI(net519));
 sg13g2_tiehi _2524__474 (.L_HI(net520));
 sg13g2_tiehi _2525__475 (.L_HI(net521));
 sg13g2_tiehi _2526__476 (.L_HI(net522));
 sg13g2_tiehi _2527__477 (.L_HI(net523));
 sg13g2_tiehi _2528__478 (.L_HI(net524));
 sg13g2_tiehi _2529__479 (.L_HI(net525));
 sg13g2_tiehi _2530__480 (.L_HI(net526));
 sg13g2_tiehi _2531__481 (.L_HI(net527));
 sg13g2_tiehi _2532__482 (.L_HI(net528));
 sg13g2_tiehi _2533__483 (.L_HI(net529));
 sg13g2_tiehi _2534__484 (.L_HI(net530));
 sg13g2_tiehi _2535__485 (.L_HI(net531));
 sg13g2_tiehi _2536__486 (.L_HI(net532));
 sg13g2_tiehi _2537__487 (.L_HI(net533));
 sg13g2_tiehi _2538__488 (.L_HI(net534));
 sg13g2_tiehi _2539__489 (.L_HI(net535));
 sg13g2_tiehi _2540__490 (.L_HI(net536));
 sg13g2_tiehi _2541__491 (.L_HI(net537));
 sg13g2_tiehi _2542__492 (.L_HI(net538));
 sg13g2_tiehi _2543__493 (.L_HI(net539));
 sg13g2_tiehi _2544__494 (.L_HI(net540));
 sg13g2_tiehi _2545__495 (.L_HI(net541));
 sg13g2_tiehi _2546__496 (.L_HI(net542));
 sg13g2_tiehi _2547__497 (.L_HI(net543));
 sg13g2_tiehi _2548__498 (.L_HI(net544));
 sg13g2_tiehi _2549__499 (.L_HI(net545));
 sg13g2_tiehi _2550__500 (.L_HI(net546));
 sg13g2_tiehi _2551__501 (.L_HI(net547));
 sg13g2_tiehi _2552__502 (.L_HI(net548));
 sg13g2_tiehi _2553__503 (.L_HI(net549));
 sg13g2_tiehi _2554__504 (.L_HI(net550));
 sg13g2_tiehi _2555__505 (.L_HI(net551));
 sg13g2_tiehi _2556__506 (.L_HI(net552));
 sg13g2_tiehi _2557__507 (.L_HI(net553));
 sg13g2_tiehi _2558__508 (.L_HI(net554));
 sg13g2_tiehi _2559__509 (.L_HI(net555));
 sg13g2_tiehi _2560__510 (.L_HI(net556));
 sg13g2_tiehi _2561__511 (.L_HI(net557));
 sg13g2_tiehi _2562__512 (.L_HI(net558));
 sg13g2_tiehi _2563__513 (.L_HI(net559));
 sg13g2_tiehi _2564__514 (.L_HI(net560));
 sg13g2_tiehi _2565__515 (.L_HI(net561));
 sg13g2_tiehi _2566__516 (.L_HI(net562));
 sg13g2_tiehi _2567__517 (.L_HI(net563));
 sg13g2_tiehi _2568__518 (.L_HI(net564));
 sg13g2_tiehi _2569__519 (.L_HI(net565));
 sg13g2_tiehi _2570__520 (.L_HI(net566));
 sg13g2_tiehi _2571__521 (.L_HI(net567));
 sg13g2_tiehi _2572__522 (.L_HI(net568));
 sg13g2_tiehi _2573__523 (.L_HI(net569));
 sg13g2_tiehi _2574__524 (.L_HI(net570));
 sg13g2_tiehi _2575__525 (.L_HI(net571));
 sg13g2_tiehi _2576__526 (.L_HI(net572));
 sg13g2_tiehi _2577__527 (.L_HI(net573));
 sg13g2_tiehi _2578__528 (.L_HI(net574));
 sg13g2_tiehi _2579__529 (.L_HI(net575));
 sg13g2_tiehi _2580__530 (.L_HI(net576));
 sg13g2_tiehi _2581__531 (.L_HI(net577));
 sg13g2_tiehi _2582__532 (.L_HI(net578));
 sg13g2_tiehi _2583__533 (.L_HI(net579));
 sg13g2_tiehi _2584__534 (.L_HI(net580));
 sg13g2_tiehi _2585__535 (.L_HI(net581));
 sg13g2_tiehi _2586__536 (.L_HI(net582));
 sg13g2_tiehi _2587__537 (.L_HI(net583));
 sg13g2_tiehi _2588__538 (.L_HI(net584));
 sg13g2_tiehi _2589__539 (.L_HI(net585));
 sg13g2_tiehi _2590__540 (.L_HI(net586));
 sg13g2_tiehi _2591__541 (.L_HI(net587));
 sg13g2_tiehi _2592__542 (.L_HI(net588));
 sg13g2_tiehi _2593__543 (.L_HI(net589));
 sg13g2_tiehi _2594__544 (.L_HI(net590));
 sg13g2_tiehi _2595__545 (.L_HI(net591));
 sg13g2_tiehi _2596__546 (.L_HI(net592));
 sg13g2_tiehi _2597__547 (.L_HI(net593));
 sg13g2_tiehi _2598__548 (.L_HI(net594));
 sg13g2_tiehi _2599__549 (.L_HI(net595));
 sg13g2_tiehi _2600__550 (.L_HI(net596));
 sg13g2_tiehi _2601__551 (.L_HI(net597));
 sg13g2_tiehi _2602__552 (.L_HI(net598));
 sg13g2_tiehi _2603__553 (.L_HI(net599));
 sg13g2_tiehi _2604__554 (.L_HI(net600));
 sg13g2_tiehi _2605__555 (.L_HI(net601));
 sg13g2_tiehi _2606__556 (.L_HI(net602));
 sg13g2_tiehi _2607__557 (.L_HI(net603));
 sg13g2_tiehi _2608__558 (.L_HI(net604));
 sg13g2_tiehi _2609__559 (.L_HI(net605));
 sg13g2_tiehi _2610__560 (.L_HI(net606));
 sg13g2_tiehi _2611__561 (.L_HI(net607));
 sg13g2_tiehi _2612__562 (.L_HI(net608));
 sg13g2_tiehi _2613__563 (.L_HI(net609));
 sg13g2_tiehi _2614__564 (.L_HI(net610));
 sg13g2_tiehi _2615__565 (.L_HI(net611));
 sg13g2_tiehi _2616__566 (.L_HI(net612));
 sg13g2_tiehi _2617__567 (.L_HI(net613));
 sg13g2_tiehi _2618__568 (.L_HI(net614));
 sg13g2_tiehi _2619__569 (.L_HI(net615));
 sg13g2_tiehi _2620__570 (.L_HI(net616));
 sg13g2_tiehi _2621__571 (.L_HI(net617));
 sg13g2_tiehi _2622__572 (.L_HI(net618));
 sg13g2_tiehi _2623__573 (.L_HI(net619));
 sg13g2_tiehi _2624__574 (.L_HI(net620));
 sg13g2_tiehi _2625__575 (.L_HI(net621));
 sg13g2_tiehi _2626__576 (.L_HI(net622));
 sg13g2_tiehi _2627__577 (.L_HI(net623));
 sg13g2_tiehi _2628__578 (.L_HI(net624));
 sg13g2_tiehi _2629__579 (.L_HI(net625));
 sg13g2_tiehi _2630__580 (.L_HI(net626));
 sg13g2_tiehi _2631__581 (.L_HI(net627));
 sg13g2_tiehi _2632__582 (.L_HI(net628));
 sg13g2_tiehi _2633__583 (.L_HI(net629));
 sg13g2_tiehi _2634__584 (.L_HI(net630));
 sg13g2_tiehi _2635__585 (.L_HI(net631));
 sg13g2_tiehi _2636__586 (.L_HI(net632));
 sg13g2_tiehi _2637__587 (.L_HI(net633));
 sg13g2_tiehi _2638__588 (.L_HI(net634));
 sg13g2_tiehi _2639__589 (.L_HI(net635));
 sg13g2_tiehi _2640__590 (.L_HI(net636));
 sg13g2_tiehi _2641__591 (.L_HI(net637));
 sg13g2_tiehi _2642__592 (.L_HI(net638));
 sg13g2_tiehi _2149__593 (.L_HI(net639));
 sg13g2_tiehi _2662__594 (.L_HI(net640));
 sg13g2_tiehi _2148__595 (.L_HI(net641));
 sg13g2_tiehi _2147__596 (.L_HI(net642));
 sg13g2_tiehi _2146__597 (.L_HI(net643));
 sg13g2_tiehi _2145__598 (.L_HI(net644));
 sg13g2_tiehi _2144__599 (.L_HI(net645));
 sg13g2_tiehi _2143__600 (.L_HI(net646));
 sg13g2_tiehi _2142__601 (.L_HI(net647));
 sg13g2_tiehi _2141__602 (.L_HI(net648));
 sg13g2_tiehi _2140__603 (.L_HI(net649));
 sg13g2_tiehi _2668__604 (.L_HI(net650));
 sg13g2_tiehi _2139__605 (.L_HI(net651));
 sg13g2_tiehi _2659__606 (.L_HI(net652));
 sg13g2_tiehi _2138__607 (.L_HI(net653));
 sg13g2_tiehi _2658__608 (.L_HI(net654));
 sg13g2_tiehi _2643__609 (.L_HI(net655));
 sg13g2_tiehi _2660__610 (.L_HI(net656));
 sg13g2_tiehi _2137__611 (.L_HI(net657));
 sg13g2_tiehi _2657__612 (.L_HI(net658));
 sg13g2_tiehi _2136__613 (.L_HI(net659));
 sg13g2_tiehi _2656__614 (.L_HI(net660));
 sg13g2_tiehi _2135__615 (.L_HI(net661));
 sg13g2_tiehi _2655__616 (.L_HI(net662));
 sg13g2_tiehi _2134__617 (.L_HI(net663));
 sg13g2_tiehi _2654__618 (.L_HI(net664));
 sg13g2_tiehi _2133__619 (.L_HI(net665));
 sg13g2_tiehi _2653__620 (.L_HI(net666));
 sg13g2_tiehi _2132__621 (.L_HI(net667));
 sg13g2_tiehi tt_um_snake_game_622 (.L_HI(net668));
 sg13g2_tiehi tt_um_snake_game_623 (.L_HI(net669));
 sg13g2_tiehi tt_um_snake_game_624 (.L_HI(net670));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_snake_game_9 (.L_LO(net9));
 sg13g2_tielo tt_um_snake_game_10 (.L_LO(net10));
 sg13g2_tielo tt_um_snake_game_11 (.L_LO(net11));
 sg13g2_tielo tt_um_snake_game_12 (.L_LO(net12));
 sg13g2_tielo tt_um_snake_game_13 (.L_LO(net13));
 sg13g2_tielo tt_um_snake_game_14 (.L_LO(net14));
 sg13g2_tielo tt_um_snake_game_15 (.L_LO(net15));
 sg13g2_tielo tt_um_snake_game_16 (.L_LO(net16));
 sg13g2_tielo tt_um_snake_game_17 (.L_LO(net17));
 sg13g2_tiehi _2652__18 (.L_HI(net18));
 sg13g2_buf_1 _3291_ (.A(failure),
    .X(uio_out[0]));
 sg13g2_buf_1 _3292_ (.A(\game_inst.o_success ),
    .X(uio_out[1]));
 sg13g2_buf_1 _3293_ (.A(eat),
    .X(uio_out[2]));
 sg13g2_buf_1 _3294_ (.A(\game_inst.o_vga_vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _3295_ (.A(\game_inst.o_vga_hsync ),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout94 (.A(net95),
    .X(net94));
 sg13g2_buf_8 fanout95 (.A(_0536_),
    .X(net95));
 sg13g2_buf_8 fanout96 (.A(net98),
    .X(net96));
 sg13g2_buf_8 fanout97 (.A(net98),
    .X(net97));
 sg13g2_buf_8 fanout98 (.A(_0419_),
    .X(net98));
 sg13g2_buf_8 fanout99 (.A(net101),
    .X(net99));
 sg13g2_buf_8 fanout100 (.A(net101),
    .X(net100));
 sg13g2_buf_8 fanout101 (.A(_0417_),
    .X(net101));
 sg13g2_buf_8 fanout102 (.A(_0391_),
    .X(net102));
 sg13g2_buf_8 fanout103 (.A(net105),
    .X(net103));
 sg13g2_buf_8 fanout104 (.A(net105),
    .X(net104));
 sg13g2_buf_8 fanout105 (.A(_0513_),
    .X(net105));
 sg13g2_buf_8 fanout106 (.A(_0437_),
    .X(net106));
 sg13g2_buf_8 fanout107 (.A(_0435_),
    .X(net107));
 sg13g2_buf_8 fanout108 (.A(net109),
    .X(net108));
 sg13g2_buf_8 fanout109 (.A(net110),
    .X(net109));
 sg13g2_buf_8 fanout110 (.A(_0433_),
    .X(net110));
 sg13g2_buf_8 fanout111 (.A(_0246_),
    .X(net111));
 sg13g2_buf_8 fanout112 (.A(net113),
    .X(net112));
 sg13g2_buf_8 fanout113 (.A(_0254_),
    .X(net113));
 sg13g2_buf_8 fanout114 (.A(_0244_),
    .X(net114));
 sg13g2_buf_8 fanout115 (.A(_0215_),
    .X(net115));
 sg13g2_buf_8 fanout116 (.A(_0214_),
    .X(net116));
 sg13g2_buf_8 fanout117 (.A(\game_inst.apple_inst.i_snake_x[0] ),
    .X(net117));
 sg13g2_buf_8 fanout118 (.A(\game_inst.control_inst.dir[0] ),
    .X(net118));
 sg13g2_buf_8 fanout119 (.A(net1335),
    .X(net119));
 sg13g2_buf_8 fanout120 (.A(\game_inst.head_y[1] ),
    .X(net120));
 sg13g2_buf_8 fanout121 (.A(net1331),
    .X(net121));
 sg13g2_buf_8 fanout122 (.A(net1295),
    .X(net122));
 sg13g2_buf_8 fanout123 (.A(net124),
    .X(net123));
 sg13g2_buf_8 fanout124 (.A(net1333),
    .X(net124));
 sg13g2_buf_8 fanout125 (.A(net1329),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(\game_inst.vga_inst.px[7] ),
    .X(net126));
 sg13g2_buf_8 fanout127 (.A(net1330),
    .X(net127));
 sg13g2_buf_8 fanout128 (.A(\game_inst.vga_inst.px[5] ),
    .X(net128));
 sg13g2_buf_8 fanout129 (.A(net1316),
    .X(net129));
 sg13g2_buf_8 fanout130 (.A(net133),
    .X(net130));
 sg13g2_buf_8 fanout131 (.A(net133),
    .X(net131));
 sg13g2_buf_1 fanout132 (.A(net133),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_0255_),
    .X(net133));
 sg13g2_buf_8 fanout134 (.A(net135),
    .X(net134));
 sg13g2_buf_8 fanout135 (.A(_0193_),
    .X(net135));
 sg13g2_buf_8 fanout136 (.A(net2),
    .X(net136));
 sg13g2_buf_8 fanout137 (.A(net138),
    .X(net137));
 sg13g2_buf_1 fanout138 (.A(net139),
    .X(net138));
 sg13g2_buf_8 fanout139 (.A(net1),
    .X(net139));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_tielo tt_um_snake_game_8 (.L_LO(net8));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_4_7_0_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_4_11_0_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_4_15_0_clk));
 sg13g2_inv_2 clkload4 (.A(clknet_leaf_75_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_leaf_10_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_37_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\game_inst.snake_inst.shiftreg_inst.memory[155][0] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold2 (.A(\game_inst.snake_inst.shiftreg_inst.memory[201][0] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold3 (.A(\game_inst.snake_inst.shiftreg_inst.memory[45][0] ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold4 (.A(\game_inst.snake_inst.shiftreg_inst.memory[221][1] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold5 (.A(\game_inst.snake_inst.shiftreg_inst.memory[179][0] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold6 (.A(\game_inst.snake_inst.shiftreg_inst.memory[228][1] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold7 (.A(\game_inst.snake_inst.shiftreg_inst.memory[13][1] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold8 (.A(\game_inst.snake_inst.shiftreg_inst.memory[23][1] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold9 (.A(\game_inst.snake_inst.shiftreg_inst.memory[223][1] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold10 (.A(\game_inst.snake_inst.shiftreg_inst.memory[17][1] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold11 (.A(\game_inst.snake_inst.shiftreg_inst.memory[32][1] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold12 (.A(\game_inst.snake_inst.shiftreg_inst.memory[157][0] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold13 (.A(\game_inst.snake_inst.shiftreg_inst.memory[214][0] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold14 (.A(\game_inst.snake_inst.shiftreg_inst.memory[187][1] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold15 (.A(\game_inst.snake_inst.shiftreg_inst.memory[104][0] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold16 (.A(\game_inst.snake_inst.shiftreg_inst.memory[16][0] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold17 (.A(\game_inst.snake_inst.shiftreg_inst.memory[3][1] ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold18 (.A(\game_inst.snake_inst.shiftreg_inst.memory[86][1] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold19 (.A(\game_inst.snake_inst.shiftreg_inst.memory[75][0] ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold20 (.A(\game_inst.snake_inst.shiftreg_inst.memory[93][0] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold21 (.A(\game_inst.snake_inst.shiftreg_inst.memory[37][1] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold22 (.A(\game_inst.snake_inst.shiftreg_inst.memory[175][1] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold23 (.A(\game_inst.snake_inst.shiftreg_inst.memory[169][1] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold24 (.A(\game_inst.snake_inst.shiftreg_inst.memory[102][0] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold25 (.A(\game_inst.snake_inst.shiftreg_inst.memory[100][0] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold26 (.A(\game_inst.snake_inst.shiftreg_inst.memory[51][1] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold27 (.A(\game_inst.snake_inst.shiftreg_inst.memory[122][1] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold28 (.A(\game_inst.snake_inst.shiftreg_inst.memory[189][1] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold29 (.A(\game_inst.snake_inst.shiftreg_inst.memory[204][0] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold30 (.A(\game_inst.snake_inst.shiftreg_inst.memory[110][0] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold31 (.A(\game_inst.snake_inst.shiftreg_inst.memory[15][1] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold32 (.A(\game_inst.snake_inst.shiftreg_inst.memory[98][0] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold33 (.A(\game_inst.snake_inst.shiftreg_inst.memory[183][1] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold34 (.A(\game_inst.snake_inst.shiftreg_inst.memory[186][0] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold35 (.A(\game_inst.snake_inst.shiftreg_inst.memory[208][0] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold36 (.A(\game_inst.snake_inst.shiftreg_inst.memory[65][1] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold37 (.A(\game_inst.snake_inst.shiftreg_inst.memory[150][0] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold38 (.A(\game_inst.snake_inst.shiftreg_inst.memory[224][0] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold39 (.A(\game_inst.snake_inst.shiftreg_inst.memory[71][0] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold40 (.A(\game_inst.snake_inst.shiftreg_inst.memory[43][0] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold41 (.A(\game_inst.snake_inst.shiftreg_inst.memory[58][1] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold42 (.A(\game_inst.snake_inst.shiftreg_inst.memory[101][0] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold43 (.A(\game_inst.snake_inst.shiftreg_inst.memory[116][1] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold44 (.A(\game_inst.snake_inst.shiftreg_inst.memory[227][0] ),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold45 (.A(\game_inst.snake_inst.shiftreg_inst.memory[184][0] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold46 (.A(\game_inst.snake_inst.shiftreg_inst.memory[198][1] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold47 (.A(\game_inst.snake_inst.shiftreg_inst.memory[55][1] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold48 (.A(\game_inst.snake_inst.shiftreg_inst.memory[225][1] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold49 (.A(\game_inst.snake_inst.shiftreg_inst.memory[69][0] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold50 (.A(\game_inst.snake_inst.shiftreg_inst.memory[54][1] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold51 (.A(\game_inst.snake_inst.shiftreg_inst.memory[78][1] ),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold52 (.A(\game_inst.snake_inst.shiftreg_inst.memory[59][1] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold53 (.A(\game_inst.snake_inst.shiftreg_inst.memory[74][1] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold54 (.A(\game_inst.snake_inst.shiftreg_inst.memory[77][0] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold55 (.A(\game_inst.snake_inst.shiftreg_inst.memory[40][0] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold56 (.A(\game_inst.snake_inst.shiftreg_inst.memory[169][0] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold57 (.A(\game_inst.snake_inst.shiftreg_inst.memory[93][1] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold58 (.A(\game_inst.snake_inst.shiftreg_inst.memory[141][0] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold59 (.A(\game_inst.snake_inst.shiftreg_inst.memory[91][0] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold60 (.A(\game_inst.snake_inst.shiftreg_inst.memory[208][1] ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold61 (.A(\game_inst.snake_inst.shiftreg_inst.memory[119][1] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold62 (.A(\game_inst.snake_inst.shiftreg_inst.memory[18][1] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold63 (.A(\game_inst.snake_inst.shiftreg_inst.memory[53][0] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold64 (.A(\game_inst.snake_inst.shiftreg_inst.memory[112][1] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold65 (.A(\game_inst.snake_inst.shiftreg_inst.memory[123][0] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold66 (.A(\game_inst.snake_inst.shiftreg_inst.memory[181][0] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold67 (.A(\game_inst.snake_inst.shiftreg_inst.memory[156][1] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold68 (.A(\game_inst.snake_inst.shiftreg_inst.memory[181][1] ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold69 (.A(\game_inst.snake_inst.shiftreg_inst.memory[144][0] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold70 (.A(\game_inst.snake_inst.shiftreg_inst.memory[117][0] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold71 (.A(\game_inst.snake_inst.shiftreg_inst.memory[121][0] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold72 (.A(\game_inst.snake_inst.shiftreg_inst.memory[146][0] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold73 (.A(\game_inst.snake_inst.shiftreg_inst.memory[39][1] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold74 (.A(\game_inst.snake_inst.shiftreg_inst.memory[105][0] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold75 (.A(\game_inst.snake_inst.shiftreg_inst.memory[35][0] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold76 (.A(\game_inst.snake_inst.shiftreg_inst.memory[70][0] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold77 (.A(\game_inst.snake_inst.shiftreg_inst.memory[185][1] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold78 (.A(\game_inst.snake_inst.shiftreg_inst.memory[91][1] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold79 (.A(\game_inst.snake_inst.shiftreg_inst.memory[21][0] ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold80 (.A(\game_inst.snake_inst.shiftreg_inst.memory[85][1] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold81 (.A(\game_inst.snake_inst.shiftreg_inst.memory[217][1] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold82 (.A(\game_inst.snake_inst.shiftreg_inst.memory[177][1] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold83 (.A(\game_inst.snake_inst.shiftreg_inst.memory[184][1] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold84 (.A(\game_inst.snake_inst.shiftreg_inst.memory[8][0] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold85 (.A(\game_inst.snake_inst.shiftreg_inst.memory[21][1] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold86 (.A(\game_inst.snake_inst.shiftreg_inst.memory[150][1] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold87 (.A(\game_inst.snake_inst.shiftreg_inst.memory[31][0] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold88 (.A(\game_inst.snake_inst.shiftreg_inst.memory[136][0] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold89 (.A(\game_inst.snake_inst.shiftreg_inst.memory[11][0] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold90 (.A(\game_inst.snake_inst.shiftreg_inst.memory[212][0] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold91 (.A(\game_inst.snake_inst.shiftreg_inst.memory[73][0] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold92 (.A(\game_inst.snake_inst.shiftreg_inst.memory[231][0] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold93 (.A(\game_inst.snake_inst.shiftreg_inst.memory[211][0] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold94 (.A(\game_inst.snake_inst.shiftreg_inst.memory[157][1] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold95 (.A(\game_inst.snake_inst.shiftreg_inst.memory[99][1] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold96 (.A(\game_inst.snake_inst.shiftreg_inst.memory[57][1] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold97 (.A(\game_inst.snake_inst.shiftreg_inst.memory[83][1] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold98 (.A(\game_inst.snake_inst.shiftreg_inst.memory[43][1] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold99 (.A(\game_inst.snake_inst.shiftreg_inst.memory[139][1] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold100 (.A(\game_inst.snake_inst.shiftreg_inst.memory[152][1] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold101 (.A(\game_inst.snake_inst.shiftreg_inst.memory[102][1] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold102 (.A(\game_inst.snake_inst.shiftreg_inst.memory[212][1] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold103 (.A(\game_inst.snake_inst.shiftreg_inst.memory[105][1] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold104 (.A(\game_inst.snake_inst.shiftreg_inst.memory[160][1] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold105 (.A(\game_inst.snake_inst.shiftreg_inst.memory[103][1] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold106 (.A(\game_inst.snake_inst.shiftreg_inst.memory[30][1] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold107 (.A(\game_inst.snake_inst.shiftreg_inst.memory[188][1] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold108 (.A(\game_inst.snake_inst.shiftreg_inst.memory[101][1] ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold109 (.A(\game_inst.snake_inst.shiftreg_inst.memory[159][1] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold110 (.A(\game_inst.snake_inst.shiftreg_inst.memory[153][1] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold111 (.A(\game_inst.snake_inst.shiftreg_inst.memory[136][1] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold112 (.A(\game_inst.snake_inst.shiftreg_inst.memory[166][0] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold113 (.A(\game_inst.snake_inst.shiftreg_inst.memory[28][0] ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold114 (.A(\game_inst.snake_inst.shiftreg_inst.memory[60][1] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold115 (.A(\game_inst.snake_inst.shiftreg_inst.memory[131][0] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold116 (.A(\game_inst.snake_inst.shiftreg_inst.memory[85][0] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold117 (.A(\game_inst.snake_inst.shiftreg_inst.memory[189][0] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold118 (.A(\game_inst.snake_inst.shiftreg_inst.memory[176][1] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold119 (.A(\game_inst.snake_inst.shiftreg_inst.memory[168][0] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold120 (.A(\game_inst.snake_inst.shiftreg_inst.memory[171][1] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold121 (.A(\game_inst.snake_inst.shiftreg_inst.memory[124][0] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold122 (.A(\game_inst.snake_inst.shiftreg_inst.memory[68][1] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold123 (.A(\game_inst.snake_inst.shiftreg_inst.memory[64][1] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold124 (.A(\game_inst.snake_inst.shiftreg_inst.memory[163][0] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold125 (.A(\game_inst.snake_inst.shiftreg_inst.memory[52][0] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold126 (.A(\game_inst.snake_inst.shiftreg_inst.memory[88][0] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold127 (.A(\game_inst.snake_inst.shiftreg_inst.memory[129][0] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold128 (.A(\game_inst.snake_inst.shiftreg_inst.memory[198][0] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold129 (.A(\game_inst.snake_inst.shiftreg_inst.memory[162][1] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold130 (.A(\game_inst.snake_inst.shiftreg_inst.memory[80][0] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold131 (.A(\game_inst.snake_inst.shiftreg_inst.memory[216][1] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold132 (.A(\game_inst.snake_inst.shiftreg_inst.memory[182][0] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold133 (.A(\game_inst.snake_inst.shiftreg_inst.memory[151][1] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold134 (.A(\game_inst.snake_inst.shiftreg_inst.memory[178][0] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold135 (.A(\game_inst.snake_inst.shiftreg_inst.memory[129][1] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold136 (.A(\game_inst.snake_inst.shiftreg_inst.memory[15][0] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold137 (.A(\game_inst.snake_inst.shiftreg_inst.memory[226][1] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold138 (.A(\game_inst.snake_inst.shiftreg_inst.memory[47][1] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold139 (.A(\game_inst.snake_inst.shiftreg_inst.memory[25][1] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold140 (.A(\game_inst.snake_inst.shiftreg_inst.memory[9][1] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold141 (.A(\game_inst.snake_inst.shiftreg_inst.memory[109][1] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold142 (.A(\game_inst.snake_inst.shiftreg_inst.memory[33][0] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold143 (.A(\game_inst.snake_inst.shiftreg_inst.memory[72][0] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold144 (.A(\game_inst.snake_inst.shiftreg_inst.memory[46][1] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold145 (.A(\game_inst.snake_inst.shiftreg_inst.memory[62][0] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold146 (.A(\game_inst.snake_inst.shiftreg_inst.memory[162][0] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold147 (.A(\game_inst.snake_inst.shiftreg_inst.memory[205][1] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold148 (.A(\game_inst.snake_inst.shiftreg_inst.memory[25][0] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold149 (.A(\game_inst.snake_inst.shiftreg_inst.memory[225][0] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold150 (.A(\game_inst.snake_inst.shiftreg_inst.memory[231][1] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold151 (.A(\game_inst.snake_inst.shiftreg_inst.memory[130][0] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold152 (.A(\game_inst.snake_inst.shiftreg_inst.memory[130][1] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold153 (.A(\game_inst.snake_inst.shiftreg_inst.memory[115][0] ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold154 (.A(\game_inst.snake_inst.shiftreg_inst.memory[194][1] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold155 (.A(\game_inst.snake_inst.shiftreg_inst.memory[154][0] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold156 (.A(\game_inst.snake_inst.shiftreg_inst.memory[20][0] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold157 (.A(\game_inst.snake_inst.shiftreg_inst.memory[73][1] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold158 (.A(\game_inst.snake_inst.shiftreg_inst.memory[151][0] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold159 (.A(\game_inst.snake_inst.shiftreg_inst.memory[62][1] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold160 (.A(\game_inst.snake_inst.shiftreg_inst.memory[108][0] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold161 (.A(\game_inst.snake_inst.shiftreg_inst.memory[66][0] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold162 (.A(\game_inst.snake_inst.shiftreg_inst.memory[203][1] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold163 (.A(\game_inst.snake_inst.shiftreg_inst.memory[29][0] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold164 (.A(\game_inst.snake_inst.shiftreg_inst.memory[188][0] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold165 (.A(\game_inst.snake_inst.shiftreg_inst.memory[58][0] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold166 (.A(\game_inst.snake_inst.shiftreg_inst.memory[180][1] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold167 (.A(\game_inst.snake_inst.shiftreg_inst.memory[210][1] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold168 (.A(\game_inst.snake_inst.shiftreg_inst.memory[48][1] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold169 (.A(\game_inst.snake_inst.shiftreg_inst.memory[128][0] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold170 (.A(\game_inst.snake_inst.shiftreg_inst.memory[170][1] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold171 (.A(\game_inst.snake_inst.shiftreg_inst.memory[81][0] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold172 (.A(\game_inst.snake_inst.shiftreg_inst.memory[13][0] ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold173 (.A(\game_inst.snake_inst.shiftreg_inst.memory[173][0] ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold174 (.A(\game_inst.snake_inst.shiftreg_inst.memory[114][0] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold175 (.A(\game_inst.snake_inst.shiftreg_inst.memory[50][1] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold176 (.A(\game_inst.snake_inst.shiftreg_inst.memory[104][1] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold177 (.A(\game_inst.snake_inst.shiftreg_inst.memory[229][1] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold178 (.A(\game_inst.snake_inst.shiftreg_inst.memory[161][1] ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold179 (.A(\game_inst.snake_inst.shiftreg_inst.memory[38][1] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold180 (.A(\game_inst.snake_inst.shiftreg_inst.memory[56][0] ),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold181 (.A(\game_inst.snake_inst.shiftreg_inst.memory[119][0] ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold182 (.A(\game_inst.snake_inst.shiftreg_inst.memory[8][1] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold183 (.A(\game_inst.snake_inst.shiftreg_inst.memory[177][0] ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold184 (.A(\game_inst.snake_inst.shiftreg_inst.memory[155][1] ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold185 (.A(\game_inst.snake_inst.shiftreg_inst.memory[1][1] ),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold186 (.A(\game_inst.snake_inst.shiftreg_inst.memory[118][0] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold187 (.A(\game_inst.snake_inst.shiftreg_inst.memory[107][0] ),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold188 (.A(\game_inst.snake_inst.shiftreg_inst.memory[124][1] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold189 (.A(\game_inst.snake_inst.shiftreg_inst.memory[84][0] ),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold190 (.A(\game_inst.snake_inst.shiftreg_inst.memory[6][0] ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold191 (.A(\game_inst.snake_inst.shiftreg_inst.memory[7][0] ),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold192 (.A(\game_inst.snake_inst.shiftreg_inst.memory[174][0] ),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold193 (.A(\game_inst.snake_inst.shiftreg_inst.memory[70][1] ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold194 (.A(\game_inst.snake_inst.shiftreg_inst.memory[113][0] ),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold195 (.A(\game_inst.snake_inst.shiftreg_inst.memory[221][0] ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold196 (.A(\game_inst.snake_inst.shiftreg_inst.memory[141][1] ),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold197 (.A(\game_inst.snake_inst.shiftreg_inst.memory[126][1] ),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold198 (.A(\game_inst.snake_inst.shiftreg_inst.memory[219][1] ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold199 (.A(\game_inst.snake_inst.shiftreg_inst.memory[164][0] ),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold200 (.A(\game_inst.snake_inst.shiftreg_inst.memory[147][0] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold201 (.A(\game_inst.snake_inst.shiftreg_inst.memory[128][1] ),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold202 (.A(\game_inst.snake_inst.shiftreg_inst.memory[6][1] ),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold203 (.A(\game_inst.snake_inst.shiftreg_inst.memory[133][1] ),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold204 (.A(\game_inst.snake_inst.shiftreg_inst.memory[47][0] ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold205 (.A(\game_inst.snake_inst.shiftreg_inst.memory[5][1] ),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold206 (.A(\game_inst.snake_inst.shiftreg_inst.memory[227][1] ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold207 (.A(\game_inst.snake_inst.shiftreg_inst.memory[37][0] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold208 (.A(\game_inst.snake_inst.shiftreg_inst.memory[134][1] ),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold209 (.A(\game_inst.snake_inst.shiftreg_inst.memory[218][0] ),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold210 (.A(\game_inst.snake_inst.shiftreg_inst.memory[165][1] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold211 (.A(\game_inst.snake_inst.shiftreg_inst.memory[2][0] ),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold212 (.A(\game_inst.snake_inst.shiftreg_inst.memory[120][1] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold213 (.A(\game_inst.snake_inst.shiftreg_inst.memory[66][1] ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold214 (.A(\game_inst.snake_inst.shiftreg_inst.memory[202][0] ),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold215 (.A(\game_inst.snake_inst.shiftreg_inst.memory[165][0] ),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold216 (.A(\game_inst.snake_inst.shiftreg_inst.memory[215][1] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold217 (.A(\game_inst.snake_inst.shiftreg_inst.memory[113][1] ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold218 (.A(\game_inst.snake_inst.shiftreg_inst.memory[34][0] ),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold219 (.A(\game_inst.snake_inst.shiftreg_inst.memory[123][1] ),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold220 (.A(\game_inst.snake_inst.shiftreg_inst.memory[125][1] ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold221 (.A(\game_inst.snake_inst.shiftreg_inst.memory[149][0] ),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold222 (.A(\game_inst.snake_inst.shiftreg_inst.memory[108][1] ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold223 (.A(\game_inst.snake_inst.shiftreg_inst.memory[122][0] ),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold224 (.A(\game_inst.snake_inst.shiftreg_inst.memory[12][0] ),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold225 (.A(\game_inst.snake_inst.shiftreg_inst.memory[172][1] ),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold226 (.A(\game_inst.snake_inst.shiftreg_inst.memory[133][0] ),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold227 (.A(\game_inst.snake_inst.shiftreg_inst.memory[7][1] ),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold228 (.A(\game_inst.snake_inst.shiftreg_inst.memory[142][1] ),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold229 (.A(\game_inst.snake_inst.shiftreg_inst.memory[36][0] ),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold230 (.A(\game_inst.snake_inst.shiftreg_inst.memory[191][0] ),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold231 (.A(\game_inst.snake_inst.shiftreg_inst.memory[164][1] ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold232 (.A(\game_inst.snake_inst.shiftreg_inst.memory[32][0] ),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold233 (.A(\game_inst.snake_inst.shiftreg_inst.memory[209][0] ),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold234 (.A(\game_inst.snake_inst.shiftreg_inst.memory[192][0] ),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold235 (.A(\game_inst.snake_inst.shiftreg_inst.memory[207][1] ),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold236 (.A(\game_inst.snake_inst.shiftreg_inst.memory[28][1] ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold237 (.A(\game_inst.snake_inst.shiftreg_inst.memory[82][0] ),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold238 (.A(\game_inst.snake_inst.shiftreg_inst.memory[1][0] ),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold239 (.A(\game_inst.snake_inst.shiftreg_inst.memory[152][0] ),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold240 (.A(\game_inst.snake_inst.shiftreg_inst.memory[71][1] ),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold241 (.A(\game_inst.snake_inst.shiftreg_inst.memory[79][0] ),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold242 (.A(\game_inst.snake_inst.shiftreg_inst.memory[200][0] ),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold243 (.A(\game_inst.snake_inst.shiftreg_inst.memory[178][1] ),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold244 (.A(\game_inst.snake_inst.shiftreg_inst.memory[140][0] ),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold245 (.A(\game_inst.snake_inst.shiftreg_inst.memory[159][0] ),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold246 (.A(\game_inst.snake_inst.shiftreg_inst.memory[111][1] ),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold247 (.A(\game_inst.snake_inst.shiftreg_inst.memory[126][0] ),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold248 (.A(\game_inst.snake_inst.shiftreg_inst.memory[60][0] ),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold249 (.A(\game_inst.snake_inst.shiftreg_inst.memory[96][0] ),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold250 (.A(\game_inst.snake_inst.shiftreg_inst.memory[154][1] ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold251 (.A(\game_inst.snake_inst.shiftreg_inst.memory[77][1] ),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold252 (.A(\game_inst.snake_inst.shiftreg_inst.memory[10][1] ),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold253 (.A(\game_inst.snake_inst.shiftreg_inst.memory[86][0] ),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold254 (.A(\game_inst.snake_inst.shiftreg_inst.memory[170][0] ),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold255 (.A(\game_inst.snake_inst.shiftreg_inst.memory[132][1] ),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold256 (.A(\game_inst.snake_inst.shiftreg_inst.memory[9][0] ),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold257 (.A(\game_inst.snake_inst.shiftreg_inst.memory[140][1] ),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold258 (.A(\game_inst.snake_inst.shiftreg_inst.memory[196][1] ),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold259 (.A(\game_inst.snake_inst.shiftreg_inst.memory[195][0] ),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold260 (.A(\game_inst.snake_inst.shiftreg_inst.memory[115][1] ),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold261 (.A(\game_inst.snake_inst.shiftreg_inst.memory[75][1] ),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold262 (.A(\game_inst.snake_inst.shiftreg_inst.memory[137][1] ),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold263 (.A(\game_inst.snake_inst.shiftreg_inst.memory[185][0] ),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold264 (.A(\game_inst.snake_inst.shiftreg_inst.memory[204][1] ),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold265 (.A(\game_inst.snake_inst.shiftreg_inst.memory[117][1] ),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold266 (.A(\game_inst.snake_inst.shiftreg_inst.memory[168][1] ),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold267 (.A(\game_inst.snake_inst.shiftreg_inst.memory[215][0] ),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold268 (.A(\game_inst.snake_inst.shiftreg_inst.memory[173][1] ),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold269 (.A(\game_inst.snake_inst.shiftreg_inst.memory[39][0] ),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold270 (.A(\game_inst.snake_inst.shiftreg_inst.memory[89][0] ),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold271 (.A(\game_inst.snake_inst.shiftreg_inst.memory[44][1] ),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold272 (.A(\game_inst.snake_inst.shiftreg_inst.memory[147][1] ),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold273 (.A(\game_inst.snake_inst.shiftreg_inst.memory[22][1] ),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold274 (.A(\game_inst.snake_inst.shiftreg_inst.memory[217][0] ),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold275 (.A(\game_inst.snake_inst.shiftreg_inst.memory[193][0] ),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold276 (.A(\game_inst.snake_inst.shiftreg_inst.memory[138][1] ),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold277 (.A(\game_inst.snake_inst.shiftreg_inst.memory[148][0] ),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold278 (.A(\game_inst.snake_inst.shiftreg_inst.memory[24][1] ),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold279 (.A(\game_inst.snake_inst.shiftreg_inst.memory[214][1] ),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold280 (.A(\game_inst.snake_inst.shiftreg_inst.memory[109][0] ),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold281 (.A(\game_inst.snake_inst.shiftreg_inst.memory[14][0] ),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold282 (.A(\game_inst.snake_inst.shiftreg_inst.memory[210][0] ),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold283 (.A(\game_inst.snake_inst.shiftreg_inst.memory[29][1] ),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold284 (.A(\game_inst.snake_inst.shiftreg_inst.memory[63][0] ),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold285 (.A(\game_inst.snake_inst.shiftreg_inst.memory[230][1] ),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold286 (.A(\game_inst.snake_inst.shiftreg_inst.memory[196][0] ),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold287 (.A(\game_inst.snake_inst.shiftreg_inst.memory[76][1] ),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold288 (.A(\game_inst.snake_inst.shiftreg_inst.memory[96][1] ),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold289 (.A(\game_inst.snake_inst.shiftreg_inst.memory[10][0] ),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold290 (.A(\game_inst.snake_inst.shiftreg_inst.memory[46][0] ),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold291 (.A(\game_inst.snake_inst.shiftreg_inst.memory[176][0] ),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold292 (.A(\game_inst.snake_inst.shiftreg_inst.memory[3][0] ),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold293 (.A(\game_inst.snake_inst.shiftreg_inst.memory[161][0] ),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold294 (.A(\game_inst.snake_inst.shiftreg_inst.memory[90][1] ),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold295 (.A(\game_inst.snake_inst.shiftreg_inst.memory[118][1] ),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold296 (.A(\game_inst.snake_inst.shiftreg_inst.memory[197][0] ),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold297 (.A(\game_inst.snake_inst.shiftreg_inst.memory[92][0] ),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold298 (.A(\game_inst.snake_inst.shiftreg_inst.memory[17][0] ),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold299 (.A(\game_inst.snake_inst.shiftreg_inst.memory[41][1] ),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold300 (.A(\game_inst.snake_inst.shiftreg_inst.memory[120][0] ),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold301 (.A(\game_inst.snake_inst.shiftreg_inst.memory[206][0] ),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold302 (.A(\game_inst.snake_inst.shiftreg_inst.memory[144][1] ),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold303 (.A(\game_inst.snake_inst.shiftreg_inst.memory[55][0] ),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold304 (.A(\game_inst.snake_inst.shiftreg_inst.memory[69][1] ),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold305 (.A(\game_inst.snake_inst.shiftreg_inst.memory[40][1] ),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold306 (.A(\game_inst.snake_inst.shiftreg_inst.memory[127][1] ),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold307 (.A(\game_inst.snake_inst.shiftreg_inst.memory[202][1] ),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold308 (.A(\game_inst.snake_inst.shiftreg_inst.memory[52][1] ),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold309 (.A(\game_inst.snake_inst.shiftreg_inst.memory[211][1] ),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold310 (.A(\game_inst.snake_inst.shiftreg_inst.memory[175][0] ),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold311 (.A(\game_inst.snake_inst.shiftreg_inst.memory[33][1] ),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold312 (.A(\game_inst.snake_inst.shiftreg_inst.memory[180][0] ),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold313 (.A(\game_inst.snake_inst.shiftreg_inst.memory[149][1] ),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold314 (.A(\game_inst.snake_inst.shiftreg_inst.memory[24][0] ),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold315 (.A(\game_inst.snake_inst.shiftreg_inst.memory[127][0] ),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold316 (.A(\game_inst.snake_inst.shiftreg_inst.memory[223][0] ),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold317 (.A(\game_inst.snake_inst.shiftreg_inst.memory[134][0] ),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold318 (.A(\game_inst.snake_inst.shiftreg_inst.memory[27][0] ),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold319 (.A(\game_inst.snake_inst.shiftreg_inst.memory[76][0] ),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold320 (.A(\game_inst.snake_inst.shiftreg_inst.memory[61][0] ),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold321 (.A(\game_inst.snake_inst.shiftreg_inst.memory[114][1] ),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold322 (.A(\game_inst.snake_inst.shiftreg_inst.memory[179][1] ),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold323 (.A(\game_inst.snake_inst.shiftreg_inst.memory[44][0] ),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold324 (.A(\game_inst.snake_inst.shiftreg_inst.memory[22][0] ),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold325 (.A(\game_inst.snake_inst.shiftreg_inst.memory[121][1] ),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold326 (.A(\game_inst.snake_inst.shiftreg_inst.memory[156][0] ),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold327 (.A(\game_inst.snake_inst.shiftreg_inst.memory[193][1] ),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold328 (.A(\game_inst.snake_inst.shiftreg_inst.memory[158][0] ),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold329 (.A(\game_inst.snake_inst.shiftreg_inst.memory[135][1] ),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold330 (.A(\game_inst.snake_inst.shiftreg_inst.memory[222][0] ),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold331 (.A(\game_inst.snake_inst.shiftreg_inst.memory[167][0] ),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold332 (.A(\game_inst.snake_inst.shiftreg_inst.memory[19][0] ),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold333 (.A(\game_inst.snake_inst.shiftreg_inst.memory[145][0] ),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold334 (.A(\game_inst.snake_inst.shiftreg_inst.memory[137][0] ),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold335 (.A(\game_inst.snake_inst.shiftreg_inst.memory[98][1] ),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold336 (.A(\game_inst.snake_inst.shiftreg_inst.memory[42][0] ),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold337 (.A(\game_inst.snake_inst.shiftreg_inst.memory[48][0] ),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold338 (.A(\game_inst.snake_inst.shiftreg_inst.memory[190][1] ),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold339 (.A(\game_inst.snake_inst.shiftreg_inst.memory[99][0] ),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold340 (.A(\game_inst.snake_inst.shiftreg_inst.memory[125][0] ),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold341 (.A(\game_inst.snake_inst.shiftreg_inst.memory[65][0] ),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold342 (.A(\game_inst.snake_inst.shiftreg_inst.memory[97][1] ),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold343 (.A(\game_inst.snake_inst.shiftreg_inst.memory[42][1] ),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold344 (.A(\game_inst.snake_inst.shiftreg_inst.memory[26][1] ),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold345 (.A(\game_inst.snake_inst.shiftreg_inst.memory[59][0] ),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold346 (.A(\game_inst.snake_inst.shiftreg_inst.memory[145][1] ),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold347 (.A(\game_inst.snake_inst.shiftreg_inst.memory[209][1] ),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold348 (.A(\game_inst.snake_inst.shiftreg_inst.memory[95][1] ),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold349 (.A(\game_inst.snake_inst.shiftreg_inst.memory[4][1] ),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold350 (.A(\game_inst.snake_inst.shiftreg_inst.memory[194][0] ),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold351 (.A(\game_inst.snake_inst.shiftreg_inst.memory[191][1] ),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold352 (.A(\game_inst.snake_inst.shiftreg_inst.memory[110][1] ),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold353 (.A(\game_inst.snake_inst.shiftreg_inst.memory[163][1] ),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold354 (.A(\game_inst.snake_inst.shiftreg_inst.memory[131][1] ),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold355 (.A(\game_inst.snake_inst.shiftreg_inst.memory[84][1] ),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold356 (.A(\game_inst.snake_inst.shiftreg_inst.memory[232][0] ),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold357 (.A(\game_inst.snake_inst.shiftreg_inst.memory[53][1] ),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold358 (.A(\game_inst.snake_inst.shiftreg_inst.memory[229][0] ),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold359 (.A(\game_inst.snake_inst.shiftreg_inst.memory[195][1] ),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold360 (.A(\game_inst.snake_inst.shiftreg_inst.memory[80][1] ),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold361 (.A(\game_inst.snake_inst.shiftreg_inst.memory[207][0] ),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold362 (.A(\game_inst.snake_inst.shiftreg_inst.memory[200][1] ),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold363 (.A(\game_inst.snake_inst.shiftreg_inst.memory[199][0] ),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold364 (.A(\game_inst.snake_inst.shiftreg_inst.memory[138][0] ),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold365 (.A(\game_inst.snake_inst.shiftreg_inst.memory[87][1] ),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold366 (.A(\game_inst.snake_inst.shiftreg_inst.memory[97][0] ),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold367 (.A(\game_inst.snake_inst.shiftreg_inst.memory[171][0] ),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold368 (.A(\game_inst.snake_inst.shiftreg_inst.memory[203][0] ),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold369 (.A(\game_inst.snake_inst.shiftreg_inst.memory[205][0] ),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold370 (.A(\game_inst.snake_inst.shiftreg_inst.memory[228][0] ),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold371 (.A(\game_inst.snake_inst.shiftreg_inst.memory[158][1] ),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold372 (.A(\game_inst.snake_inst.shiftreg_inst.memory[82][1] ),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold373 (.A(\game_inst.snake_inst.shiftreg_inst.memory[14][1] ),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold374 (.A(\game_inst.snake_inst.shiftreg_inst.memory[116][0] ),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold375 (.A(\game_inst.snake_inst.shiftreg_inst.memory[63][1] ),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold376 (.A(\game_inst.snake_inst.shiftreg_inst.memory[132][0] ),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold377 (.A(\game_inst.snake_inst.shiftreg_inst.memory[35][1] ),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold378 (.A(\game_inst.snake_inst.shiftreg_inst.memory[38][0] ),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold379 (.A(\game_inst.snake_inst.shiftreg_inst.memory[103][0] ),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold380 (.A(\game_inst.snake_inst.shiftreg_inst.memory[83][0] ),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold381 (.A(\game_inst.snake_inst.shiftreg_inst.memory[4][0] ),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold382 (.A(\game_inst.snake_inst.shiftreg_inst.memory[26][0] ),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold383 (.A(\game_inst.snake_inst.shiftreg_inst.memory[172][0] ),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold384 (.A(\game_inst.snake_inst.shiftreg_inst.memory[222][1] ),
    .X(net1054));
 sg13g2_dlygate4sd3_1 hold385 (.A(\game_inst.snake_inst.shiftreg_inst.memory[34][1] ),
    .X(net1055));
 sg13g2_dlygate4sd3_1 hold386 (.A(\game_inst.snake_inst.shiftreg_inst.memory[199][1] ),
    .X(net1056));
 sg13g2_dlygate4sd3_1 hold387 (.A(\game_inst.snake_inst.shiftreg_inst.memory[78][0] ),
    .X(net1057));
 sg13g2_dlygate4sd3_1 hold388 (.A(\game_inst.snake_inst.shiftreg_inst.memory[160][0] ),
    .X(net1058));
 sg13g2_dlygate4sd3_1 hold389 (.A(\game_inst.snake_inst.shiftreg_inst.memory[232][1] ),
    .X(net1059));
 sg13g2_dlygate4sd3_1 hold390 (.A(\game_inst.snake_inst.shiftreg_inst.memory[230][0] ),
    .X(net1060));
 sg13g2_dlygate4sd3_1 hold391 (.A(\game_inst.snake_inst.shiftreg_inst.memory[166][1] ),
    .X(net1061));
 sg13g2_dlygate4sd3_1 hold392 (.A(\game_inst.snake_inst.shiftreg_inst.memory[94][0] ),
    .X(net1062));
 sg13g2_dlygate4sd3_1 hold393 (.A(\game_inst.snake_inst.shiftreg_inst.memory[16][1] ),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold394 (.A(\game_inst.snake_inst.shiftreg_inst.memory[89][1] ),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold395 (.A(\game_inst.snake_inst.shiftreg_inst.memory[142][0] ),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold396 (.A(\game_inst.snake_inst.shiftreg_inst.memory[139][0] ),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold397 (.A(\game_inst.snake_inst.shiftreg_inst.memory[67][1] ),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold398 (.A(\game_inst.snake_inst.shiftreg_inst.memory[12][1] ),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold399 (.A(\game_inst.snake_inst.shiftreg_inst.memory[41][0] ),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold400 (.A(\game_inst.snake_inst.shiftreg_inst.memory[220][1] ),
    .X(net1070));
 sg13g2_dlygate4sd3_1 hold401 (.A(\game_inst.snake_inst.shiftreg_inst.memory[81][1] ),
    .X(net1071));
 sg13g2_dlygate4sd3_1 hold402 (.A(\game_inst.snake_inst.shiftreg_inst.memory[201][1] ),
    .X(net1072));
 sg13g2_dlygate4sd3_1 hold403 (.A(\game_inst.snake_inst.shiftreg_inst.memory[57][0] ),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold404 (.A(\game_inst.snake_inst.shiftreg_inst.memory[153][0] ),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold405 (.A(\game_inst.snake_inst.shiftreg_inst.memory[79][1] ),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold406 (.A(\game_inst.snake_inst.shiftreg_inst.memory[219][0] ),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold407 (.A(\game_inst.snake_inst.shiftreg_inst.memory[49][0] ),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold408 (.A(\game_inst.snake_inst.shiftreg_inst.memory[56][1] ),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold409 (.A(\game_inst.snake_inst.shiftreg_inst.memory[95][0] ),
    .X(net1079));
 sg13g2_dlygate4sd3_1 hold410 (.A(\game_inst.snake_inst.shiftreg_inst.memory[226][0] ),
    .X(net1080));
 sg13g2_dlygate4sd3_1 hold411 (.A(\game_inst.snake_inst.shiftreg_inst.memory[187][0] ),
    .X(net1081));
 sg13g2_dlygate4sd3_1 hold412 (.A(\game_inst.snake_inst.shiftreg_inst.memory[51][0] ),
    .X(net1082));
 sg13g2_dlygate4sd3_1 hold413 (.A(\game_inst.snake_inst.shiftreg_inst.memory[220][0] ),
    .X(net1083));
 sg13g2_dlygate4sd3_1 hold414 (.A(\game_inst.snake_inst.shiftreg_inst.memory[49][1] ),
    .X(net1084));
 sg13g2_dlygate4sd3_1 hold415 (.A(\game_inst.snake_inst.shiftreg_inst.memory[27][1] ),
    .X(net1085));
 sg13g2_dlygate4sd3_1 hold416 (.A(\game_inst.snake_inst.shiftreg_inst.memory[67][0] ),
    .X(net1086));
 sg13g2_dlygate4sd3_1 hold417 (.A(\game_inst.snake_inst.shiftreg_inst.memory[106][0] ),
    .X(net1087));
 sg13g2_dlygate4sd3_1 hold418 (.A(\game_inst.snake_inst.shiftreg_inst.memory[2][1] ),
    .X(net1088));
 sg13g2_dlygate4sd3_1 hold419 (.A(\game_inst.snake_inst.shiftreg_inst.memory[192][1] ),
    .X(net1089));
 sg13g2_dlygate4sd3_1 hold420 (.A(\game_inst.snake_inst.shiftreg_inst.memory[216][0] ),
    .X(net1090));
 sg13g2_dlygate4sd3_1 hold421 (.A(\game_inst.snake_inst.shiftreg_inst.memory[5][0] ),
    .X(net1091));
 sg13g2_dlygate4sd3_1 hold422 (.A(\game_inst.snake_inst.shiftreg_inst.memory[90][0] ),
    .X(net1092));
 sg13g2_dlygate4sd3_1 hold423 (.A(\game_inst.snake_inst.shiftreg_inst.memory[213][1] ),
    .X(net1093));
 sg13g2_dlygate4sd3_1 hold424 (.A(\game_inst.snake_inst.shiftreg_inst.memory[72][1] ),
    .X(net1094));
 sg13g2_dlygate4sd3_1 hold425 (.A(\game_inst.snake_inst.shiftreg_inst.memory[64][0] ),
    .X(net1095));
 sg13g2_dlygate4sd3_1 hold426 (.A(\game_inst.snake_inst.shiftreg_inst.memory[206][1] ),
    .X(net1096));
 sg13g2_dlygate4sd3_1 hold427 (.A(\game_inst.snake_inst.shiftreg_inst.memory[190][0] ),
    .X(net1097));
 sg13g2_dlygate4sd3_1 hold428 (.A(\game_inst.snake_inst.shiftreg_inst.memory[186][1] ),
    .X(net1098));
 sg13g2_dlygate4sd3_1 hold429 (.A(\game_inst.snake_inst.shiftreg_inst.memory[54][0] ),
    .X(net1099));
 sg13g2_dlygate4sd3_1 hold430 (.A(\game_inst.snake_inst.shiftreg_inst.memory[20][1] ),
    .X(net1100));
 sg13g2_dlygate4sd3_1 hold431 (.A(\game_inst.snake_inst.shiftreg_inst.memory[31][1] ),
    .X(net1101));
 sg13g2_dlygate4sd3_1 hold432 (.A(\game_inst.snake_inst.shiftreg_inst.memory[224][1] ),
    .X(net1102));
 sg13g2_dlygate4sd3_1 hold433 (.A(\game_inst.snake_inst.shiftreg_inst.memory[45][1] ),
    .X(net1103));
 sg13g2_dlygate4sd3_1 hold434 (.A(\game_inst.snake_inst.shiftreg_inst.memory[74][0] ),
    .X(net1104));
 sg13g2_dlygate4sd3_1 hold435 (.A(\game_inst.snake_inst.shiftreg_inst.memory[111][0] ),
    .X(net1105));
 sg13g2_dlygate4sd3_1 hold436 (.A(\game_inst.snake_inst.shiftreg_inst.memory[30][0] ),
    .X(net1106));
 sg13g2_dlygate4sd3_1 hold437 (.A(\game_inst.snake_inst.shiftreg_inst.memory[36][1] ),
    .X(net1107));
 sg13g2_dlygate4sd3_1 hold438 (.A(\game_inst.snake_inst.shiftreg_inst.memory[61][1] ),
    .X(net1108));
 sg13g2_dlygate4sd3_1 hold439 (.A(\game_inst.snake_inst.shiftreg_inst.memory[197][1] ),
    .X(net1109));
 sg13g2_dlygate4sd3_1 hold440 (.A(\game_inst.snake_inst.shiftreg_inst.memory[94][1] ),
    .X(net1110));
 sg13g2_dlygate4sd3_1 hold441 (.A(\game_inst.snake_inst.shiftreg_inst.memory[213][0] ),
    .X(net1111));
 sg13g2_dlygate4sd3_1 hold442 (.A(\game_inst.snake_inst.shiftreg_inst.memory[68][0] ),
    .X(net1112));
 sg13g2_dlygate4sd3_1 hold443 (.A(\game_inst.snake_inst.shiftreg_inst.memory[23][0] ),
    .X(net1113));
 sg13g2_dlygate4sd3_1 hold444 (.A(\game_inst.snake_inst.shiftreg_inst.memory[218][1] ),
    .X(net1114));
 sg13g2_dlygate4sd3_1 hold445 (.A(\game_inst.snake_inst.shiftreg_inst.memory[18][0] ),
    .X(net1115));
 sg13g2_dlygate4sd3_1 hold446 (.A(\game_inst.snake_inst.shiftreg_inst.memory[107][1] ),
    .X(net1116));
 sg13g2_dlygate4sd3_1 hold447 (.A(\game_inst.snake_inst.shiftreg_inst.memory[183][0] ),
    .X(net1117));
 sg13g2_dlygate4sd3_1 hold448 (.A(\game_inst.snake_inst.shiftreg_inst.memory[87][0] ),
    .X(net1118));
 sg13g2_dlygate4sd3_1 hold449 (.A(\game_inst.snake_inst.shiftreg_inst.memory[19][1] ),
    .X(net1119));
 sg13g2_dlygate4sd3_1 hold450 (.A(\game_inst.snake_inst.shiftreg_inst.memory[88][1] ),
    .X(net1120));
 sg13g2_dlygate4sd3_1 hold451 (.A(\game_inst.snake_inst.shiftreg_inst.memory[11][1] ),
    .X(net1121));
 sg13g2_dlygate4sd3_1 hold452 (.A(\game_inst.snake_inst.shiftreg_inst.memory[174][1] ),
    .X(net1122));
 sg13g2_dlygate4sd3_1 hold453 (.A(\game_inst.snake_inst.shiftreg_inst.memory[143][0] ),
    .X(net1123));
 sg13g2_dlygate4sd3_1 hold454 (.A(\game_inst.snake_inst.shiftreg_inst.memory[167][1] ),
    .X(net1124));
 sg13g2_dlygate4sd3_1 hold455 (.A(\game_inst.snake_inst.shiftreg_inst.memory[100][1] ),
    .X(net1125));
 sg13g2_dlygate4sd3_1 hold456 (.A(\game_inst.snake_inst.shiftreg_inst.memory[146][1] ),
    .X(net1126));
 sg13g2_dlygate4sd3_1 hold457 (.A(\game_inst.snake_inst.shiftreg_inst.memory[92][1] ),
    .X(net1127));
 sg13g2_dlygate4sd3_1 hold458 (.A(\game_inst.snake_inst.shiftreg_inst.memory[143][1] ),
    .X(net1128));
 sg13g2_dlygate4sd3_1 hold459 (.A(\game_inst.snake_inst.shiftreg_inst.memory[50][0] ),
    .X(net1129));
 sg13g2_dlygate4sd3_1 hold460 (.A(\game_inst.snake_inst.shiftreg_inst.memory[148][1] ),
    .X(net1130));
 sg13g2_dlygate4sd3_1 hold461 (.A(\game_inst.snake_inst.shiftreg_inst.memory[106][1] ),
    .X(net1131));
 sg13g2_dlygate4sd3_1 hold462 (.A(\game_inst.snake_inst.shiftreg_inst.memory[182][1] ),
    .X(net1132));
 sg13g2_dlygate4sd3_1 hold463 (.A(\game_inst.snake_inst.shiftreg_inst.memory[112][0] ),
    .X(net1133));
 sg13g2_dlygate4sd3_1 hold464 (.A(\game_inst.snake_inst.shiftreg_inst.memory[135][0] ),
    .X(net1134));
 sg13g2_dlygate4sd3_1 hold465 (.A(\game_inst.snake_inst.dir_first[0] ),
    .X(net1135));
 sg13g2_dlygate4sd3_1 hold466 (.A(\game_inst.vga_inst.px[0] ),
    .X(net1136));
 sg13g2_dlygate4sd3_1 hold467 (.A(\game_inst.vga_inst.pos_counter[0] ),
    .X(net1137));
 sg13g2_dlygate4sd3_1 hold468 (.A(_0042_),
    .X(net1138));
 sg13g2_dlygate4sd3_1 hold469 (.A(\game_inst.snake_inst.dir_first[1] ),
    .X(net1139));
 sg13g2_dlygate4sd3_1 hold470 (.A(\game_inst.o_vga_vsync ),
    .X(net1140));
 sg13g2_dlygate4sd3_1 hold471 (.A(\game_inst.vga_inst.px[2] ),
    .X(net1141));
 sg13g2_dlygate4sd3_1 hold472 (.A(_0454_),
    .X(net1142));
 sg13g2_dlygate4sd3_1 hold473 (.A(_0020_),
    .X(net1143));
 sg13g2_dlygate4sd3_1 hold474 (.A(\game_inst.tickgen_inst.counter_max[4] ),
    .X(net1144));
 sg13g2_dlygate4sd3_1 hold475 (.A(_0130_),
    .X(net1145));
 sg13g2_dlygate4sd3_1 hold476 (.A(\game_inst.snake_inst.length[7] ),
    .X(net1146));
 sg13g2_dlygate4sd3_1 hold477 (.A(_0109_),
    .X(net1147));
 sg13g2_dlygate4sd3_1 hold478 (.A(\game_inst.tick ),
    .X(net1148));
 sg13g2_dlygate4sd3_1 hold479 (.A(_0125_),
    .X(net1149));
 sg13g2_dlygate4sd3_1 hold480 (.A(\game_inst.apple_inst.test ),
    .X(net1150));
 sg13g2_dlygate4sd3_1 hold481 (.A(_0061_),
    .X(net1151));
 sg13g2_dlygate4sd3_1 hold482 (.A(\game_inst.snake_inst.dir_out[0] ),
    .X(net1152));
 sg13g2_dlygate4sd3_1 hold483 (.A(_0038_),
    .X(net1153));
 sg13g2_dlygate4sd3_1 hold484 (.A(\game_inst.apple_inst.random_inst.lfsr4[0] ),
    .X(net1154));
 sg13g2_dlygate4sd3_1 hold485 (.A(_0067_),
    .X(net1155));
 sg13g2_dlygate4sd3_1 hold486 (.A(\game_inst.control_inst.i_head_dir[0] ),
    .X(net1156));
 sg13g2_dlygate4sd3_1 hold487 (.A(_0079_),
    .X(net1157));
 sg13g2_dlygate4sd3_1 hold488 (.A(\game_inst.vga_inst.pos_counter[1] ),
    .X(net1158));
 sg13g2_dlygate4sd3_1 hold489 (.A(_0043_),
    .X(net1159));
 sg13g2_dlygate4sd3_1 hold490 (.A(\game_inst.snake_inst.dir_out[1] ),
    .X(net1160));
 sg13g2_dlygate4sd3_1 hold491 (.A(_0477_),
    .X(net1161));
 sg13g2_dlygate4sd3_1 hold492 (.A(\game_inst.apple_inst.random_inst.lfsr5[1] ),
    .X(net1162));
 sg13g2_dlygate4sd3_1 hold493 (.A(_0056_),
    .X(net1163));
 sg13g2_dlygate4sd3_1 hold494 (.A(\game_inst.apple_inst.random_inst.lfsr5[3] ),
    .X(net1164));
 sg13g2_dlygate4sd3_1 hold495 (.A(_0058_),
    .X(net1165));
 sg13g2_dlygate4sd3_1 hold496 (.A(\game_inst.vga_inst.py[3] ),
    .X(net1166));
 sg13g2_dlygate4sd3_1 hold497 (.A(_0047_),
    .X(net1167));
 sg13g2_dlygate4sd3_1 hold498 (.A(\game_inst.snake_inst.pos[4] ),
    .X(net1168));
 sg13g2_dlygate4sd3_1 hold499 (.A(_0685_),
    .X(net1169));
 sg13g2_dlygate4sd3_1 hold500 (.A(_0112_),
    .X(net1170));
 sg13g2_dlygate4sd3_1 hold501 (.A(\game_inst.control_inst.o_start ),
    .X(net1171));
 sg13g2_dlygate4sd3_1 hold502 (.A(_0121_),
    .X(net1172));
 sg13g2_dlygate4sd3_1 hold503 (.A(\game_inst.vga_inst.row_buffer[17][1] ),
    .X(net1173));
 sg13g2_dlygate4sd3_1 hold504 (.A(\game_inst.snake_inst.length[3] ),
    .X(net1174));
 sg13g2_dlygate4sd3_1 hold505 (.A(_0673_),
    .X(net1175));
 sg13g2_dlygate4sd3_1 hold506 (.A(_0105_),
    .X(net1176));
 sg13g2_dlygate4sd3_1 hold507 (.A(\game_inst.vga_inst.row_buffer[7][0] ),
    .X(net1177));
 sg13g2_dlygate4sd3_1 hold508 (.A(\game_inst.apple_inst.random_inst.lfsr5[2] ),
    .X(net1178));
 sg13g2_dlygate4sd3_1 hold509 (.A(_0057_),
    .X(net1179));
 sg13g2_dlygate4sd3_1 hold510 (.A(\game_inst.apple_inst.o_ready ),
    .X(net1180));
 sg13g2_dlygate4sd3_1 hold511 (.A(_0536_),
    .X(net1181));
 sg13g2_dlygate4sd3_1 hold512 (.A(\game_inst.vga_inst.py[2] ),
    .X(net1182));
 sg13g2_dlygate4sd3_1 hold513 (.A(_0046_),
    .X(net1183));
 sg13g2_dlygate4sd3_1 hold514 (.A(\game_inst.vga_inst.row_buffer[9][1] ),
    .X(net1184));
 sg13g2_dlygate4sd3_1 hold515 (.A(\game_inst.vga_inst.py[1] ),
    .X(net1185));
 sg13g2_dlygate4sd3_1 hold516 (.A(_0045_),
    .X(net1186));
 sg13g2_dlygate4sd3_1 hold517 (.A(\game_inst.vga_inst.row_buffer[1][1] ),
    .X(net1187));
 sg13g2_dlygate4sd3_1 hold518 (.A(\game_inst.vga_inst.row_buffer[16][0] ),
    .X(net1188));
 sg13g2_dlygate4sd3_1 hold519 (.A(\game_inst.vga_inst.row_buffer[17][0] ),
    .X(net1189));
 sg13g2_dlygate4sd3_1 hold520 (.A(\game_inst.vga_inst.row_buffer[6][1] ),
    .X(net1190));
 sg13g2_dlygate4sd3_1 hold521 (.A(\game_inst.vga_inst.row_buffer[12][1] ),
    .X(net1191));
 sg13g2_dlygate4sd3_1 hold522 (.A(\game_inst.apple_inst.random_inst.lfsr5[0] ),
    .X(net1192));
 sg13g2_dlygate4sd3_1 hold523 (.A(_0055_),
    .X(net1193));
 sg13g2_dlygate4sd3_1 hold524 (.A(\game_inst.vga_inst.row_buffer[8][1] ),
    .X(net1194));
 sg13g2_dlygate4sd3_1 hold525 (.A(\game_inst.vga_inst.row_buffer[10][1] ),
    .X(net1195));
 sg13g2_dlygate4sd3_1 hold526 (.A(\game_inst.vga_inst.row_buffer[16][1] ),
    .X(net1196));
 sg13g2_dlygate4sd3_1 hold527 (.A(\game_inst.vga_inst.row_buffer[11][0] ),
    .X(net1197));
 sg13g2_dlygate4sd3_1 hold528 (.A(\game_inst.snake_inst.length[1] ),
    .X(net1198));
 sg13g2_dlygate4sd3_1 hold529 (.A(_0670_),
    .X(net1199));
 sg13g2_dlygate4sd3_1 hold530 (.A(_0103_),
    .X(net1200));
 sg13g2_dlygate4sd3_1 hold531 (.A(\game_inst.vga_inst.row_buffer[12][0] ),
    .X(net1201));
 sg13g2_dlygate4sd3_1 hold532 (.A(\game_inst.vga_inst.row_buffer[7][1] ),
    .X(net1202));
 sg13g2_dlygate4sd3_1 hold533 (.A(\game_inst.vga_inst.row_buffer[8][0] ),
    .X(net1203));
 sg13g2_dlygate4sd3_1 hold534 (.A(\game_inst.vga_inst.row_buffer[15][1] ),
    .X(net1204));
 sg13g2_dlygate4sd3_1 hold535 (.A(\game_inst.vga_inst.row_buffer[11][1] ),
    .X(net1205));
 sg13g2_dlygate4sd3_1 hold536 (.A(\game_inst.snake_inst.pos[0] ),
    .X(net1206));
 sg13g2_dlygate4sd3_1 hold537 (.A(_0011_),
    .X(net1207));
 sg13g2_dlygate4sd3_1 hold538 (.A(\game_inst.vga_inst.row_buffer[5][1] ),
    .X(net1208));
 sg13g2_dlygate4sd3_1 hold539 (.A(\game_inst.vga_inst.row_buffer[9][0] ),
    .X(net1209));
 sg13g2_dlygate4sd3_1 hold540 (.A(\game_inst.vga_inst.row_buffer[13][0] ),
    .X(net1210));
 sg13g2_dlygate4sd3_1 hold541 (.A(\game_inst.vga_inst.row_buffer[6][0] ),
    .X(net1211));
 sg13g2_dlygate4sd3_1 hold542 (.A(\game_inst.vga_inst.row_buffer[13][1] ),
    .X(net1212));
 sg13g2_dlygate4sd3_1 hold543 (.A(\game_inst.apple_inst.random_inst.lfsr4[2] ),
    .X(net1213));
 sg13g2_dlygate4sd3_1 hold544 (.A(_0119_),
    .X(net1214));
 sg13g2_dlygate4sd3_1 hold545 (.A(\game_inst.vga_inst.row_buffer[0][1] ),
    .X(net1215));
 sg13g2_dlygate4sd3_1 hold546 (.A(\game_inst.vga_inst.row_buffer[1][0] ),
    .X(net1216));
 sg13g2_dlygate4sd3_1 hold547 (.A(\game_inst.vga_inst.py[9] ),
    .X(net1217));
 sg13g2_dlygate4sd3_1 hold548 (.A(_0053_),
    .X(net1218));
 sg13g2_dlygate4sd3_1 hold549 (.A(\game_inst.vga_inst.row_buffer[5][0] ),
    .X(net1219));
 sg13g2_dlygate4sd3_1 hold550 (.A(\game_inst.apple_inst.apple_y[0] ),
    .X(net1220));
 sg13g2_dlygate4sd3_1 hold551 (.A(\game_inst.vga_inst.row_buffer[2][0] ),
    .X(net1221));
 sg13g2_dlygate4sd3_1 hold552 (.A(\game_inst.vga_inst.row_buffer[10][0] ),
    .X(net1222));
 sg13g2_dlygate4sd3_1 hold553 (.A(\game_inst.apple_inst.random_inst.lfsr5[4] ),
    .X(net1223));
 sg13g2_dlygate4sd3_1 hold554 (.A(\game_inst.vga_inst.row_buffer[15][0] ),
    .X(net1224));
 sg13g2_dlygate4sd3_1 hold555 (.A(\game_inst.vga_inst.py[4] ),
    .X(net1225));
 sg13g2_dlygate4sd3_1 hold556 (.A(_0493_),
    .X(net1226));
 sg13g2_dlygate4sd3_1 hold557 (.A(\game_inst.apple_inst.random_inst.lfsr4[1] ),
    .X(net1227));
 sg13g2_dlygate4sd3_1 hold558 (.A(\game_inst.vga_inst.row_buffer[14][1] ),
    .X(net1228));
 sg13g2_dlygate4sd3_1 hold559 (.A(\game_inst.vga_inst.px[3] ),
    .X(net1229));
 sg13g2_dlygate4sd3_1 hold560 (.A(_0455_),
    .X(net1230));
 sg13g2_dlygate4sd3_1 hold561 (.A(_0021_),
    .X(net1231));
 sg13g2_dlygate4sd3_1 hold562 (.A(\game_inst.vga_inst.row_buffer[14][0] ),
    .X(net1232));
 sg13g2_dlygate4sd3_1 hold563 (.A(\game_inst.apple_inst.random_inst.lfsr4[3] ),
    .X(net1233));
 sg13g2_dlygate4sd3_1 hold564 (.A(\game_inst.apple_inst.apple_x[4] ),
    .X(net1234));
 sg13g2_dlygate4sd3_1 hold565 (.A(\game_inst.vga_inst.row_buffer[4][1] ),
    .X(net1235));
 sg13g2_dlygate4sd3_1 hold566 (.A(\game_inst.vga_inst.row_buffer[0][0] ),
    .X(net1236));
 sg13g2_dlygate4sd3_1 hold567 (.A(\game_inst.vga_inst.row_buffer[3][1] ),
    .X(net1237));
 sg13g2_dlygate4sd3_1 hold568 (.A(\game_inst.vga_inst.px[1] ),
    .X(net1238));
 sg13g2_dlygate4sd3_1 hold569 (.A(\game_inst.vga_inst.row_buffer[2][1] ),
    .X(net1239));
 sg13g2_dlygate4sd3_1 hold570 (.A(\game_inst.apple_inst.apple_y[3] ),
    .X(net1240));
 sg13g2_dlygate4sd3_1 hold571 (.A(\game_inst.vga_inst.py[7] ),
    .X(net1241));
 sg13g2_dlygate4sd3_1 hold572 (.A(_0051_),
    .X(net1242));
 sg13g2_dlygate4sd3_1 hold573 (.A(\game_inst.vga_inst.row_buffer[4][0] ),
    .X(net1243));
 sg13g2_dlygate4sd3_1 hold574 (.A(\game_inst.vga_inst.row_buffer[3][0] ),
    .X(net1244));
 sg13g2_dlygate4sd3_1 hold575 (.A(\game_inst.apple_inst.apple_y[1] ),
    .X(net1245));
 sg13g2_dlygate4sd3_1 hold576 (.A(\game_inst.o_success ),
    .X(net1246));
 sg13g2_dlygate4sd3_1 hold577 (.A(_0506_),
    .X(net1247));
 sg13g2_dlygate4sd3_1 hold578 (.A(\game_inst.control_inst.backwards[1] ),
    .X(net1248));
 sg13g2_dlygate4sd3_1 hold579 (.A(_0553_),
    .X(net1249));
 sg13g2_dlygate4sd3_1 hold580 (.A(_0080_),
    .X(net1250));
 sg13g2_dlygate4sd3_1 hold581 (.A(\game_inst.tickgen_inst.counter[1] ),
    .X(net1251));
 sg13g2_dlygate4sd3_1 hold582 (.A(_0728_),
    .X(net1252));
 sg13g2_dlygate4sd3_1 hold583 (.A(_0132_),
    .X(net1253));
 sg13g2_dlygate4sd3_1 hold584 (.A(\game_inst.tickgen_inst.counter[0] ),
    .X(net1254));
 sg13g2_dlygate4sd3_1 hold585 (.A(_0726_),
    .X(net1255));
 sg13g2_dlygate4sd3_1 hold586 (.A(_0131_),
    .X(net1256));
 sg13g2_dlygate4sd3_1 hold587 (.A(failure),
    .X(net1257));
 sg13g2_dlygate4sd3_1 hold588 (.A(_0136_),
    .X(net1258));
 sg13g2_dlygate4sd3_1 hold589 (.A(\game_inst.snake_inst.pos[2] ),
    .X(net1259));
 sg13g2_dlygate4sd3_1 hold590 (.A(_0684_),
    .X(net1260));
 sg13g2_dlygate4sd3_1 hold591 (.A(_0111_),
    .X(net1261));
 sg13g2_dlygate4sd3_1 hold592 (.A(\game_inst.tickgen_inst.counter[2] ),
    .X(net1262));
 sg13g2_dlygate4sd3_1 hold593 (.A(\game_inst.apple_inst.i_snake_valid ),
    .X(net1263));
 sg13g2_dlygate4sd3_1 hold594 (.A(_0520_),
    .X(net1264));
 sg13g2_dlygate4sd3_1 hold595 (.A(\game_inst.snake_inst.length[6] ),
    .X(net1265));
 sg13g2_dlygate4sd3_1 hold596 (.A(_0680_),
    .X(net1266));
 sg13g2_dlygate4sd3_1 hold597 (.A(_0108_),
    .X(net1267));
 sg13g2_dlygate4sd3_1 hold598 (.A(\game_inst.colorblind ),
    .X(net1268));
 sg13g2_dlygate4sd3_1 hold599 (.A(_0692_),
    .X(net1269));
 sg13g2_dlygate4sd3_1 hold600 (.A(_0124_),
    .X(net1270));
 sg13g2_dlygate4sd3_1 hold601 (.A(\game_inst.vga_inst.py[8] ),
    .X(net1271));
 sg13g2_dlygate4sd3_1 hold602 (.A(_0239_),
    .X(net1272));
 sg13g2_dlygate4sd3_1 hold603 (.A(\game_inst.apple_inst.i_snake_y[2] ),
    .X(net1273));
 sg13g2_dlygate4sd3_1 hold604 (.A(\game_inst.snake_inst.length[2] ),
    .X(net1274));
 sg13g2_dlygate4sd3_1 hold605 (.A(_0672_),
    .X(net1275));
 sg13g2_dlygate4sd3_1 hold606 (.A(\game_inst.tickgen_inst.counter_max[3] ),
    .X(net1276));
 sg13g2_dlygate4sd3_1 hold607 (.A(\game_inst.snake_inst.length[5] ),
    .X(net1277));
 sg13g2_dlygate4sd3_1 hold608 (.A(_0679_),
    .X(net1278));
 sg13g2_dlygate4sd3_1 hold609 (.A(_0107_),
    .X(net1279));
 sg13g2_dlygate4sd3_1 hold610 (.A(\game_inst.tickgen_inst.counter_max[1] ),
    .X(net1280));
 sg13g2_dlygate4sd3_1 hold611 (.A(_0708_),
    .X(net1281));
 sg13g2_dlygate4sd3_1 hold612 (.A(_0127_),
    .X(net1282));
 sg13g2_dlygate4sd3_1 hold613 (.A(\game_inst.head_y[3] ),
    .X(net1283));
 sg13g2_dlygate4sd3_1 hold614 (.A(\game_inst.head_x[4] ),
    .X(net1284));
 sg13g2_dlygate4sd3_1 hold615 (.A(\game_inst.tickgen_inst.counter_max[0] ),
    .X(net1285));
 sg13g2_dlygate4sd3_1 hold616 (.A(_0126_),
    .X(net1286));
 sg13g2_dlygate4sd3_1 hold617 (.A(\game_inst.vga_inst.py[6] ),
    .X(net1287));
 sg13g2_dlygate4sd3_1 hold618 (.A(_0496_),
    .X(net1288));
 sg13g2_dlygate4sd3_1 hold619 (.A(\game_inst.vga_inst.px[4] ),
    .X(net1289));
 sg13g2_dlygate4sd3_1 hold620 (.A(\game_inst.tickgen_inst.counter[3] ),
    .X(net1290));
 sg13g2_dlygate4sd3_1 hold621 (.A(\game_inst.head_x[1] ),
    .X(net1291));
 sg13g2_dlygate4sd3_1 hold622 (.A(\game_inst.head_y[1] ),
    .X(net1292));
 sg13g2_dlygate4sd3_1 hold623 (.A(_0087_),
    .X(net1293));
 sg13g2_dlygate4sd3_1 hold624 (.A(\game_inst.apple_inst.i_snake_y[3] ),
    .X(net1294));
 sg13g2_dlygate4sd3_1 hold625 (.A(\game_inst.vga_inst.py[5] ),
    .X(net1295));
 sg13g2_dlygate4sd3_1 hold626 (.A(\game_inst.snake_inst.length[0] ),
    .X(net1296));
 sg13g2_dlygate4sd3_1 hold627 (.A(\game_inst.head_x[2] ),
    .X(net1297));
 sg13g2_dlygate4sd3_1 hold628 (.A(\game_inst.snake_inst.pos[6] ),
    .X(net1298));
 sg13g2_dlygate4sd3_1 hold629 (.A(_0639_),
    .X(net1299));
 sg13g2_dlygate4sd3_1 hold630 (.A(_0643_),
    .X(net1300));
 sg13g2_dlygate4sd3_1 hold631 (.A(_0644_),
    .X(net1301));
 sg13g2_dlygate4sd3_1 hold632 (.A(\game_inst.tickgen_inst.counter_max[2] ),
    .X(net1302));
 sg13g2_dlygate4sd3_1 hold633 (.A(_0714_),
    .X(net1303));
 sg13g2_dlygate4sd3_1 hold634 (.A(\game_inst.snake_inst.pos[5] ),
    .X(net1304));
 sg13g2_dlygate4sd3_1 hold635 (.A(\game_inst.snake_inst.pos[1] ),
    .X(net1305));
 sg13g2_dlygate4sd3_1 hold636 (.A(\game_inst.vga_inst.py[0] ),
    .X(net1306));
 sg13g2_dlygate4sd3_1 hold637 (.A(\game_inst.apple_inst.i_snake_y[1] ),
    .X(net1307));
 sg13g2_dlygate4sd3_1 hold638 (.A(_0099_),
    .X(net1308));
 sg13g2_dlygate4sd3_1 hold639 (.A(\game_inst.apple_inst.i_snake_x[2] ),
    .X(net1309));
 sg13g2_dlygate4sd3_1 hold640 (.A(\game_inst.tickgen_inst.counter[4] ),
    .X(net1310));
 sg13g2_dlygate4sd3_1 hold641 (.A(_0135_),
    .X(net1311));
 sg13g2_dlygate4sd3_1 hold642 (.A(\game_inst.snake_inst.pos[7] ),
    .X(net1312));
 sg13g2_dlygate4sd3_1 hold643 (.A(\game_inst.apple_inst.i_snake_x[4] ),
    .X(net1313));
 sg13g2_dlygate4sd3_1 hold644 (.A(\game_inst.head_y[0] ),
    .X(net1314));
 sg13g2_dlygate4sd3_1 hold645 (.A(_0086_),
    .X(net1315));
 sg13g2_dlygate4sd3_1 hold646 (.A(\game_inst.vga_inst.px[5] ),
    .X(net1316));
 sg13g2_dlygate4sd3_1 hold647 (.A(\game_inst.snake_inst.pos[3] ),
    .X(net1317));
 sg13g2_dlygate4sd3_1 hold648 (.A(\game_inst.apple_inst.i_snake_x[3] ),
    .X(net1318));
 sg13g2_dlygate4sd3_1 hold649 (.A(_0095_),
    .X(net1319));
 sg13g2_dlygate4sd3_1 hold650 (.A(\game_inst.head_x[0] ),
    .X(net1320));
 sg13g2_dlygate4sd3_1 hold651 (.A(_0081_),
    .X(net1321));
 sg13g2_dlygate4sd3_1 hold652 (.A(\game_inst.snake_inst.length[4] ),
    .X(net1322));
 sg13g2_dlygate4sd3_1 hold653 (.A(\game_inst.apple_inst.i_snake_x[1] ),
    .X(net1323));
 sg13g2_dlygate4sd3_1 hold654 (.A(_0093_),
    .X(net1324));
 sg13g2_dlygate4sd3_1 hold655 (.A(\game_inst.control_inst.dir[1] ),
    .X(net1325));
 sg13g2_dlygate4sd3_1 hold656 (.A(\game_inst.apple_inst.i_snake_x[0] ),
    .X(net1326));
 sg13g2_dlygate4sd3_1 hold657 (.A(\game_inst.vga_inst.px[9] ),
    .X(net1327));
 sg13g2_dlygate4sd3_1 hold658 (.A(_0001_),
    .X(net1328));
 sg13g2_dlygate4sd3_1 hold659 (.A(\game_inst.vga_inst.px[7] ),
    .X(net1329));
 sg13g2_dlygate4sd3_1 hold660 (.A(\game_inst.vga_inst.px[6] ),
    .X(net1330));
 sg13g2_dlygate4sd3_1 hold661 (.A(\game_inst.head_x[3] ),
    .X(net1331));
 sg13g2_dlygate4sd3_1 hold662 (.A(_0084_),
    .X(net1332));
 sg13g2_dlygate4sd3_1 hold663 (.A(\game_inst.vga_inst.px[8] ),
    .X(net1333));
 sg13g2_dlygate4sd3_1 hold664 (.A(\game_inst.apple_inst.i_snake_y[0] ),
    .X(net1334));
 sg13g2_dlygate4sd3_1 hold665 (.A(\game_inst.head_y[2] ),
    .X(net1335));
 sg13g2_dlygate4sd3_1 hold666 (.A(\game_inst.control_inst.dir[1] ),
    .X(net1336));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_fill_2 FILLER_0_112 ();
 sg13g2_fill_1 FILLER_0_114 ();
 sg13g2_fill_2 FILLER_0_136 ();
 sg13g2_fill_1 FILLER_0_138 ();
 sg13g2_fill_2 FILLER_0_215 ();
 sg13g2_fill_2 FILLER_0_238 ();
 sg13g2_fill_2 FILLER_0_257 ();
 sg13g2_fill_1 FILLER_0_259 ();
 sg13g2_fill_2 FILLER_0_336 ();
 sg13g2_fill_2 FILLER_0_387 ();
 sg13g2_fill_1 FILLER_0_389 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_fill_2 FILLER_1_105 ();
 sg13g2_fill_1 FILLER_1_107 ();
 sg13g2_fill_2 FILLER_1_306 ();
 sg13g2_fill_1 FILLER_1_308 ();
 sg13g2_fill_1 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_4 FILLER_2_91 ();
 sg13g2_fill_2 FILLER_2_95 ();
 sg13g2_fill_2 FILLER_2_105 ();
 sg13g2_fill_2 FILLER_2_272 ();
 sg13g2_fill_1 FILLER_2_355 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_fill_1 FILLER_3_91 ();
 sg13g2_fill_1 FILLER_3_222 ();
 sg13g2_fill_2 FILLER_3_312 ();
 sg13g2_fill_1 FILLER_3_341 ();
 sg13g2_fill_2 FILLER_3_369 ();
 sg13g2_fill_1 FILLER_3_371 ();
 sg13g2_fill_1 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_4 FILLER_4_70 ();
 sg13g2_fill_2 FILLER_4_78 ();
 sg13g2_fill_1 FILLER_4_133 ();
 sg13g2_fill_1 FILLER_4_161 ();
 sg13g2_fill_1 FILLER_4_201 ();
 sg13g2_fill_1 FILLER_4_237 ();
 sg13g2_fill_2 FILLER_4_287 ();
 sg13g2_fill_2 FILLER_4_347 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_fill_1 FILLER_5_35 ();
 sg13g2_decap_4 FILLER_5_40 ();
 sg13g2_fill_2 FILLER_5_44 ();
 sg13g2_fill_1 FILLER_5_59 ();
 sg13g2_fill_1 FILLER_5_68 ();
 sg13g2_fill_2 FILLER_5_86 ();
 sg13g2_fill_1 FILLER_5_88 ();
 sg13g2_fill_1 FILLER_5_152 ();
 sg13g2_fill_2 FILLER_5_184 ();
 sg13g2_fill_1 FILLER_5_186 ();
 sg13g2_fill_1 FILLER_5_214 ();
 sg13g2_fill_2 FILLER_5_228 ();
 sg13g2_fill_2 FILLER_5_243 ();
 sg13g2_fill_2 FILLER_5_315 ();
 sg13g2_fill_1 FILLER_5_317 ();
 sg13g2_fill_2 FILLER_5_380 ();
 sg13g2_decap_4 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_4 ();
 sg13g2_decap_8 FILLER_6_17 ();
 sg13g2_decap_8 FILLER_6_24 ();
 sg13g2_fill_1 FILLER_6_58 ();
 sg13g2_fill_1 FILLER_6_108 ();
 sg13g2_fill_1 FILLER_6_201 ();
 sg13g2_fill_2 FILLER_6_363 ();
 sg13g2_fill_1 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_32 ();
 sg13g2_fill_2 FILLER_7_96 ();
 sg13g2_fill_1 FILLER_7_161 ();
 sg13g2_fill_1 FILLER_7_202 ();
 sg13g2_fill_2 FILLER_7_270 ();
 sg13g2_fill_1 FILLER_7_317 ();
 sg13g2_fill_2 FILLER_7_376 ();
 sg13g2_fill_1 FILLER_7_378 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_fill_1 FILLER_8_44 ();
 sg13g2_fill_2 FILLER_8_85 ();
 sg13g2_fill_1 FILLER_8_87 ();
 sg13g2_fill_2 FILLER_8_115 ();
 sg13g2_fill_2 FILLER_8_148 ();
 sg13g2_fill_1 FILLER_8_150 ();
 sg13g2_fill_1 FILLER_8_182 ();
 sg13g2_fill_1 FILLER_8_210 ();
 sg13g2_fill_2 FILLER_8_259 ();
 sg13g2_fill_1 FILLER_8_261 ();
 sg13g2_fill_2 FILLER_8_355 ();
 sg13g2_fill_1 FILLER_8_357 ();
 sg13g2_fill_2 FILLER_8_398 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_42 ();
 sg13g2_fill_1 FILLER_9_127 ();
 sg13g2_fill_2 FILLER_9_132 ();
 sg13g2_fill_1 FILLER_9_152 ();
 sg13g2_fill_1 FILLER_9_166 ();
 sg13g2_fill_2 FILLER_9_216 ();
 sg13g2_fill_2 FILLER_9_272 ();
 sg13g2_fill_1 FILLER_9_274 ();
 sg13g2_fill_1 FILLER_9_310 ();
 sg13g2_fill_2 FILLER_9_377 ();
 sg13g2_fill_1 FILLER_9_379 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_2 ();
 sg13g2_fill_1 FILLER_10_42 ();
 sg13g2_fill_2 FILLER_10_110 ();
 sg13g2_fill_2 FILLER_10_143 ();
 sg13g2_fill_1 FILLER_10_145 ();
 sg13g2_fill_1 FILLER_10_159 ();
 sg13g2_fill_2 FILLER_10_191 ();
 sg13g2_fill_1 FILLER_10_193 ();
 sg13g2_fill_2 FILLER_10_230 ();
 sg13g2_fill_2 FILLER_10_259 ();
 sg13g2_fill_1 FILLER_10_265 ();
 sg13g2_fill_2 FILLER_10_310 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_fill_1 FILLER_11_147 ();
 sg13g2_fill_2 FILLER_11_250 ();
 sg13g2_fill_1 FILLER_11_252 ();
 sg13g2_fill_2 FILLER_11_280 ();
 sg13g2_fill_1 FILLER_11_282 ();
 sg13g2_fill_2 FILLER_11_310 ();
 sg13g2_fill_1 FILLER_11_312 ();
 sg13g2_fill_1 FILLER_11_370 ();
 sg13g2_fill_2 FILLER_11_380 ();
 sg13g2_fill_1 FILLER_12_72 ();
 sg13g2_fill_1 FILLER_12_209 ();
 sg13g2_fill_1 FILLER_12_245 ();
 sg13g2_fill_2 FILLER_12_303 ();
 sg13g2_fill_1 FILLER_12_305 ();
 sg13g2_fill_2 FILLER_12_355 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_86 ();
 sg13g2_fill_2 FILLER_13_128 ();
 sg13g2_fill_1 FILLER_13_130 ();
 sg13g2_fill_1 FILLER_13_167 ();
 sg13g2_fill_1 FILLER_13_203 ();
 sg13g2_fill_2 FILLER_13_231 ();
 sg13g2_fill_1 FILLER_13_277 ();
 sg13g2_fill_1 FILLER_13_291 ();
 sg13g2_fill_2 FILLER_13_319 ();
 sg13g2_fill_1 FILLER_13_321 ();
 sg13g2_fill_1 FILLER_13_349 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_fill_1 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_126 ();
 sg13g2_fill_1 FILLER_14_159 ();
 sg13g2_fill_1 FILLER_14_381 ();
 sg13g2_fill_2 FILLER_15_31 ();
 sg13g2_fill_1 FILLER_15_33 ();
 sg13g2_fill_1 FILLER_15_91 ();
 sg13g2_fill_1 FILLER_15_185 ();
 sg13g2_fill_1 FILLER_15_217 ();
 sg13g2_fill_2 FILLER_15_245 ();
 sg13g2_fill_1 FILLER_15_306 ();
 sg13g2_fill_1 FILLER_15_338 ();
 sg13g2_fill_1 FILLER_15_388 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_fill_2 FILLER_16_161 ();
 sg13g2_fill_2 FILLER_16_172 ();
 sg13g2_fill_2 FILLER_16_219 ();
 sg13g2_fill_2 FILLER_16_234 ();
 sg13g2_fill_1 FILLER_16_236 ();
 sg13g2_fill_1 FILLER_16_257 ();
 sg13g2_fill_1 FILLER_16_347 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_fill_2 FILLER_17_31 ();
 sg13g2_fill_2 FILLER_17_46 ();
 sg13g2_fill_2 FILLER_17_111 ();
 sg13g2_fill_1 FILLER_17_113 ();
 sg13g2_fill_2 FILLER_17_136 ();
 sg13g2_fill_2 FILLER_17_210 ();
 sg13g2_fill_1 FILLER_17_212 ();
 sg13g2_fill_2 FILLER_17_273 ();
 sg13g2_fill_1 FILLER_17_288 ();
 sg13g2_fill_1 FILLER_18_40 ();
 sg13g2_fill_2 FILLER_18_50 ();
 sg13g2_fill_1 FILLER_18_52 ();
 sg13g2_fill_1 FILLER_18_75 ();
 sg13g2_fill_2 FILLER_18_130 ();
 sg13g2_fill_2 FILLER_18_208 ();
 sg13g2_fill_1 FILLER_18_210 ();
 sg13g2_fill_1 FILLER_18_215 ();
 sg13g2_fill_2 FILLER_18_243 ();
 sg13g2_fill_2 FILLER_18_254 ();
 sg13g2_fill_2 FILLER_18_284 ();
 sg13g2_fill_1 FILLER_18_286 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_fill_1 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_14 ();
 sg13g2_fill_1 FILLER_19_69 ();
 sg13g2_fill_2 FILLER_19_101 ();
 sg13g2_fill_2 FILLER_19_160 ();
 sg13g2_fill_1 FILLER_19_162 ();
 sg13g2_fill_1 FILLER_19_176 ();
 sg13g2_fill_2 FILLER_19_193 ();
 sg13g2_fill_1 FILLER_19_195 ();
 sg13g2_fill_2 FILLER_19_312 ();
 sg13g2_fill_2 FILLER_19_332 ();
 sg13g2_fill_1 FILLER_19_365 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_2 ();
 sg13g2_fill_1 FILLER_20_12 ();
 sg13g2_fill_2 FILLER_20_76 ();
 sg13g2_fill_1 FILLER_20_78 ();
 sg13g2_decap_8 FILLER_20_101 ();
 sg13g2_decap_4 FILLER_20_108 ();
 sg13g2_fill_1 FILLER_20_116 ();
 sg13g2_fill_2 FILLER_20_176 ();
 sg13g2_fill_1 FILLER_20_205 ();
 sg13g2_fill_1 FILLER_20_224 ();
 sg13g2_fill_1 FILLER_20_261 ();
 sg13g2_fill_2 FILLER_20_305 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_2 ();
 sg13g2_fill_2 FILLER_21_30 ();
 sg13g2_fill_1 FILLER_21_32 ();
 sg13g2_fill_2 FILLER_21_73 ();
 sg13g2_fill_1 FILLER_21_75 ();
 sg13g2_decap_4 FILLER_21_121 ();
 sg13g2_fill_1 FILLER_21_125 ();
 sg13g2_fill_1 FILLER_21_135 ();
 sg13g2_fill_2 FILLER_21_176 ();
 sg13g2_fill_1 FILLER_21_209 ();
 sg13g2_fill_2 FILLER_21_220 ();
 sg13g2_fill_1 FILLER_21_222 ();
 sg13g2_fill_2 FILLER_21_232 ();
 sg13g2_fill_1 FILLER_21_234 ();
 sg13g2_fill_1 FILLER_21_242 ();
 sg13g2_fill_1 FILLER_21_263 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_65 ();
 sg13g2_fill_1 FILLER_22_67 ();
 sg13g2_fill_1 FILLER_22_131 ();
 sg13g2_fill_2 FILLER_22_173 ();
 sg13g2_fill_2 FILLER_22_185 ();
 sg13g2_fill_1 FILLER_22_228 ();
 sg13g2_fill_2 FILLER_22_262 ();
 sg13g2_fill_1 FILLER_22_306 ();
 sg13g2_fill_1 FILLER_22_351 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_42 ();
 sg13g2_fill_1 FILLER_23_44 ();
 sg13g2_fill_1 FILLER_23_112 ();
 sg13g2_fill_1 FILLER_23_161 ();
 sg13g2_fill_1 FILLER_23_168 ();
 sg13g2_fill_2 FILLER_23_201 ();
 sg13g2_fill_1 FILLER_23_203 ();
 sg13g2_fill_1 FILLER_23_255 ();
 sg13g2_fill_2 FILLER_23_383 ();
 sg13g2_fill_1 FILLER_23_385 ();
 sg13g2_fill_1 FILLER_23_399 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_decap_4 FILLER_24_122 ();
 sg13g2_fill_1 FILLER_24_177 ();
 sg13g2_fill_2 FILLER_24_228 ();
 sg13g2_fill_1 FILLER_24_230 ();
 sg13g2_fill_1 FILLER_24_253 ();
 sg13g2_fill_1 FILLER_24_282 ();
 sg13g2_fill_2 FILLER_24_319 ();
 sg13g2_fill_2 FILLER_24_348 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_2 ();
 sg13g2_fill_1 FILLER_25_11 ();
 sg13g2_fill_1 FILLER_25_24 ();
 sg13g2_fill_1 FILLER_25_52 ();
 sg13g2_fill_1 FILLER_25_66 ();
 sg13g2_fill_2 FILLER_25_80 ();
 sg13g2_fill_1 FILLER_25_147 ();
 sg13g2_fill_2 FILLER_25_162 ();
 sg13g2_fill_1 FILLER_25_164 ();
 sg13g2_fill_2 FILLER_25_224 ();
 sg13g2_fill_1 FILLER_25_226 ();
 sg13g2_fill_2 FILLER_25_345 ();
 sg13g2_fill_1 FILLER_25_347 ();
 sg13g2_fill_2 FILLER_25_379 ();
 sg13g2_fill_1 FILLER_25_381 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_4 ();
 sg13g2_fill_1 FILLER_26_9 ();
 sg13g2_fill_1 FILLER_26_54 ();
 sg13g2_fill_2 FILLER_26_236 ();
 sg13g2_fill_1 FILLER_26_238 ();
 sg13g2_fill_1 FILLER_26_270 ();
 sg13g2_fill_2 FILLER_26_357 ();
 sg13g2_fill_1 FILLER_26_359 ();
 sg13g2_fill_2 FILLER_26_378 ();
 sg13g2_fill_1 FILLER_26_380 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_4 ();
 sg13g2_fill_1 FILLER_27_14 ();
 sg13g2_fill_1 FILLER_27_132 ();
 sg13g2_fill_1 FILLER_27_170 ();
 sg13g2_fill_1 FILLER_27_212 ();
 sg13g2_fill_1 FILLER_27_217 ();
 sg13g2_fill_2 FILLER_27_228 ();
 sg13g2_fill_2 FILLER_27_304 ();
 sg13g2_fill_1 FILLER_27_306 ();
 sg13g2_fill_1 FILLER_27_399 ();
 sg13g2_fill_1 FILLER_28_31 ();
 sg13g2_fill_2 FILLER_28_72 ();
 sg13g2_fill_1 FILLER_28_74 ();
 sg13g2_fill_2 FILLER_28_133 ();
 sg13g2_fill_1 FILLER_28_172 ();
 sg13g2_fill_1 FILLER_28_187 ();
 sg13g2_fill_2 FILLER_28_192 ();
 sg13g2_fill_2 FILLER_28_247 ();
 sg13g2_fill_2 FILLER_28_295 ();
 sg13g2_fill_2 FILLER_28_342 ();
 sg13g2_fill_1 FILLER_28_380 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_76 ();
 sg13g2_fill_2 FILLER_29_127 ();
 sg13g2_fill_1 FILLER_29_129 ();
 sg13g2_fill_2 FILLER_29_189 ();
 sg13g2_fill_2 FILLER_29_200 ();
 sg13g2_fill_1 FILLER_29_202 ();
 sg13g2_fill_1 FILLER_29_295 ();
 sg13g2_fill_2 FILLER_29_363 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_43 ();
 sg13g2_fill_1 FILLER_30_67 ();
 sg13g2_fill_1 FILLER_30_77 ();
 sg13g2_fill_1 FILLER_30_114 ();
 sg13g2_fill_1 FILLER_30_195 ();
 sg13g2_fill_2 FILLER_30_294 ();
 sg13g2_fill_2 FILLER_30_346 ();
 sg13g2_fill_2 FILLER_30_379 ();
 sg13g2_fill_1 FILLER_30_381 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_81 ();
 sg13g2_fill_2 FILLER_31_173 ();
 sg13g2_fill_1 FILLER_31_207 ();
 sg13g2_fill_2 FILLER_31_226 ();
 sg13g2_fill_1 FILLER_31_246 ();
 sg13g2_fill_1 FILLER_31_258 ();
 sg13g2_fill_2 FILLER_31_362 ();
 sg13g2_fill_1 FILLER_31_364 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_4 FILLER_32_20 ();
 sg13g2_fill_2 FILLER_32_24 ();
 sg13g2_fill_2 FILLER_32_129 ();
 sg13g2_fill_1 FILLER_32_159 ();
 sg13g2_fill_2 FILLER_32_173 ();
 sg13g2_fill_1 FILLER_32_216 ();
 sg13g2_fill_2 FILLER_32_254 ();
 sg13g2_fill_1 FILLER_32_256 ();
 sg13g2_fill_2 FILLER_32_285 ();
 sg13g2_fill_1 FILLER_32_287 ();
 sg13g2_fill_1 FILLER_32_315 ();
 sg13g2_fill_1 FILLER_32_356 ();
 sg13g2_fill_2 FILLER_32_396 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_fill_2 FILLER_33_21 ();
 sg13g2_fill_1 FILLER_33_23 ();
 sg13g2_fill_2 FILLER_33_189 ();
 sg13g2_fill_1 FILLER_33_213 ();
 sg13g2_fill_2 FILLER_33_230 ();
 sg13g2_fill_2 FILLER_33_243 ();
 sg13g2_fill_1 FILLER_33_245 ();
 sg13g2_fill_2 FILLER_33_253 ();
 sg13g2_fill_2 FILLER_33_301 ();
 sg13g2_fill_1 FILLER_33_303 ();
 sg13g2_fill_1 FILLER_33_326 ();
 sg13g2_fill_2 FILLER_33_367 ();
 sg13g2_fill_1 FILLER_33_369 ();
 sg13g2_fill_1 FILLER_33_374 ();
 sg13g2_decap_8 FILLER_33_387 ();
 sg13g2_decap_8 FILLER_33_394 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_14 ();
 sg13g2_fill_1 FILLER_34_131 ();
 sg13g2_fill_2 FILLER_34_172 ();
 sg13g2_fill_1 FILLER_34_184 ();
 sg13g2_fill_2 FILLER_34_199 ();
 sg13g2_decap_4 FILLER_34_232 ();
 sg13g2_fill_1 FILLER_34_236 ();
 sg13g2_fill_1 FILLER_34_275 ();
 sg13g2_fill_1 FILLER_34_313 ();
 sg13g2_fill_2 FILLER_34_345 ();
 sg13g2_decap_8 FILLER_34_383 ();
 sg13g2_decap_4 FILLER_34_390 ();
 sg13g2_fill_2 FILLER_34_394 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_83 ();
 sg13g2_fill_1 FILLER_35_94 ();
 sg13g2_fill_1 FILLER_35_99 ();
 sg13g2_fill_2 FILLER_35_187 ();
 sg13g2_decap_8 FILLER_35_201 ();
 sg13g2_fill_2 FILLER_35_208 ();
 sg13g2_fill_2 FILLER_35_223 ();
 sg13g2_decap_8 FILLER_35_243 ();
 sg13g2_fill_1 FILLER_35_274 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_4 ();
 sg13g2_fill_2 FILLER_36_32 ();
 sg13g2_fill_1 FILLER_36_34 ();
 sg13g2_fill_2 FILLER_36_84 ();
 sg13g2_fill_1 FILLER_36_86 ();
 sg13g2_fill_2 FILLER_36_109 ();
 sg13g2_decap_8 FILLER_36_197 ();
 sg13g2_decap_8 FILLER_36_204 ();
 sg13g2_fill_2 FILLER_36_211 ();
 sg13g2_decap_8 FILLER_36_235 ();
 sg13g2_decap_4 FILLER_36_247 ();
 sg13g2_fill_1 FILLER_36_251 ();
 sg13g2_fill_1 FILLER_36_257 ();
 sg13g2_decap_8 FILLER_36_267 ();
 sg13g2_decap_4 FILLER_36_274 ();
 sg13g2_fill_2 FILLER_36_278 ();
 sg13g2_fill_1 FILLER_36_339 ();
 sg13g2_decap_8 FILLER_36_402 ();
 sg13g2_fill_2 FILLER_37_88 ();
 sg13g2_fill_1 FILLER_37_90 ();
 sg13g2_fill_1 FILLER_37_190 ();
 sg13g2_fill_2 FILLER_37_196 ();
 sg13g2_fill_2 FILLER_37_202 ();
 sg13g2_fill_2 FILLER_37_216 ();
 sg13g2_fill_2 FILLER_37_221 ();
 sg13g2_fill_1 FILLER_37_228 ();
 sg13g2_fill_1 FILLER_37_233 ();
 sg13g2_decap_8 FILLER_37_276 ();
 sg13g2_fill_2 FILLER_37_283 ();
 sg13g2_fill_2 FILLER_37_332 ();
 sg13g2_fill_1 FILLER_37_334 ();
 sg13g2_decap_8 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_15 ();
 sg13g2_fill_1 FILLER_38_17 ();
 sg13g2_fill_2 FILLER_38_116 ();
 sg13g2_fill_1 FILLER_38_164 ();
 sg13g2_fill_2 FILLER_38_191 ();
 sg13g2_fill_1 FILLER_38_201 ();
 sg13g2_fill_2 FILLER_38_207 ();
 sg13g2_fill_1 FILLER_38_238 ();
 sg13g2_fill_2 FILLER_38_250 ();
 sg13g2_fill_1 FILLER_38_283 ();
 sg13g2_fill_1 FILLER_38_311 ();
 sg13g2_fill_2 FILLER_38_321 ();
 sg13g2_decap_4 FILLER_38_391 ();
 sg13g2_fill_2 FILLER_38_395 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_fill_2 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_37 ();
 sg13g2_fill_2 FILLER_39_74 ();
 sg13g2_fill_1 FILLER_39_76 ();
 sg13g2_fill_2 FILLER_39_113 ();
 sg13g2_fill_1 FILLER_39_115 ();
 sg13g2_fill_1 FILLER_39_125 ();
 sg13g2_decap_4 FILLER_39_193 ();
 sg13g2_fill_2 FILLER_39_276 ();
 sg13g2_fill_1 FILLER_39_342 ();
 sg13g2_fill_2 FILLER_39_351 ();
 sg13g2_decap_8 FILLER_39_366 ();
 sg13g2_decap_4 FILLER_39_373 ();
 sg13g2_fill_1 FILLER_39_377 ();
 sg13g2_decap_4 FILLER_39_405 ();
 sg13g2_decap_4 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_4 ();
 sg13g2_fill_2 FILLER_40_64 ();
 sg13g2_fill_1 FILLER_40_66 ();
 sg13g2_decap_8 FILLER_40_103 ();
 sg13g2_decap_4 FILLER_40_110 ();
 sg13g2_decap_4 FILLER_40_169 ();
 sg13g2_fill_2 FILLER_40_205 ();
 sg13g2_fill_1 FILLER_40_220 ();
 sg13g2_fill_1 FILLER_40_239 ();
 sg13g2_fill_1 FILLER_40_288 ();
 sg13g2_decap_8 FILLER_40_399 ();
 sg13g2_fill_2 FILLER_40_406 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_7 ();
 sg13g2_fill_1 FILLER_41_9 ();
 sg13g2_decap_8 FILLER_41_94 ();
 sg13g2_fill_2 FILLER_41_101 ();
 sg13g2_fill_1 FILLER_41_103 ();
 sg13g2_decap_8 FILLER_41_108 ();
 sg13g2_decap_4 FILLER_41_115 ();
 sg13g2_fill_2 FILLER_41_127 ();
 sg13g2_fill_2 FILLER_41_179 ();
 sg13g2_fill_1 FILLER_41_181 ();
 sg13g2_fill_2 FILLER_41_190 ();
 sg13g2_fill_1 FILLER_41_192 ();
 sg13g2_fill_1 FILLER_41_213 ();
 sg13g2_fill_2 FILLER_41_227 ();
 sg13g2_fill_1 FILLER_41_235 ();
 sg13g2_fill_1 FILLER_41_361 ();
 sg13g2_decap_8 FILLER_41_389 ();
 sg13g2_decap_8 FILLER_41_396 ();
 sg13g2_decap_4 FILLER_41_403 ();
 sg13g2_fill_2 FILLER_41_407 ();
 sg13g2_fill_2 FILLER_42_31 ();
 sg13g2_fill_1 FILLER_42_33 ();
 sg13g2_fill_2 FILLER_42_65 ();
 sg13g2_fill_1 FILLER_42_67 ();
 sg13g2_fill_1 FILLER_42_81 ();
 sg13g2_fill_2 FILLER_42_104 ();
 sg13g2_decap_8 FILLER_42_115 ();
 sg13g2_decap_8 FILLER_42_122 ();
 sg13g2_decap_4 FILLER_42_129 ();
 sg13g2_fill_2 FILLER_42_182 ();
 sg13g2_fill_1 FILLER_42_184 ();
 sg13g2_fill_1 FILLER_42_210 ();
 sg13g2_fill_1 FILLER_42_226 ();
 sg13g2_fill_2 FILLER_42_263 ();
 sg13g2_fill_1 FILLER_42_281 ();
 sg13g2_fill_2 FILLER_42_323 ();
 sg13g2_fill_2 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_2 ();
 sg13g2_fill_2 FILLER_43_91 ();
 sg13g2_fill_1 FILLER_43_93 ();
 sg13g2_decap_8 FILLER_43_121 ();
 sg13g2_decap_8 FILLER_43_128 ();
 sg13g2_fill_1 FILLER_43_150 ();
 sg13g2_decap_4 FILLER_43_175 ();
 sg13g2_fill_2 FILLER_43_179 ();
 sg13g2_fill_1 FILLER_43_257 ();
 sg13g2_fill_1 FILLER_43_264 ();
 sg13g2_decap_4 FILLER_43_278 ();
 sg13g2_fill_2 FILLER_43_303 ();
 sg13g2_fill_2 FILLER_43_363 ();
 sg13g2_fill_1 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_32 ();
 sg13g2_fill_1 FILLER_44_34 ();
 sg13g2_fill_1 FILLER_44_166 ();
 sg13g2_fill_2 FILLER_44_202 ();
 sg13g2_decap_4 FILLER_44_225 ();
 sg13g2_fill_2 FILLER_44_229 ();
 sg13g2_decap_4 FILLER_44_251 ();
 sg13g2_fill_1 FILLER_44_255 ();
 sg13g2_decap_8 FILLER_44_278 ();
 sg13g2_decap_4 FILLER_44_285 ();
 sg13g2_fill_1 FILLER_44_289 ();
 sg13g2_fill_2 FILLER_44_376 ();
 sg13g2_fill_1 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_14 ();
 sg13g2_fill_2 FILLER_45_42 ();
 sg13g2_fill_1 FILLER_45_44 ();
 sg13g2_fill_1 FILLER_45_171 ();
 sg13g2_decap_4 FILLER_45_196 ();
 sg13g2_fill_1 FILLER_45_200 ();
 sg13g2_decap_8 FILLER_45_204 ();
 sg13g2_decap_8 FILLER_45_215 ();
 sg13g2_decap_8 FILLER_45_222 ();
 sg13g2_decap_4 FILLER_45_229 ();
 sg13g2_fill_2 FILLER_45_233 ();
 sg13g2_decap_8 FILLER_45_242 ();
 sg13g2_decap_8 FILLER_45_249 ();
 sg13g2_decap_4 FILLER_45_256 ();
 sg13g2_fill_2 FILLER_45_260 ();
 sg13g2_fill_2 FILLER_45_266 ();
 sg13g2_decap_8 FILLER_45_281 ();
 sg13g2_fill_1 FILLER_45_288 ();
 sg13g2_fill_1 FILLER_45_323 ();
 sg13g2_fill_2 FILLER_45_357 ();
 sg13g2_fill_1 FILLER_45_359 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_2 ();
 sg13g2_fill_1 FILLER_46_66 ();
 sg13g2_fill_1 FILLER_46_121 ();
 sg13g2_fill_1 FILLER_46_153 ();
 sg13g2_fill_2 FILLER_46_181 ();
 sg13g2_decap_8 FILLER_46_189 ();
 sg13g2_decap_8 FILLER_46_196 ();
 sg13g2_decap_4 FILLER_46_203 ();
 sg13g2_decap_8 FILLER_46_212 ();
 sg13g2_decap_8 FILLER_46_219 ();
 sg13g2_fill_2 FILLER_46_226 ();
 sg13g2_fill_1 FILLER_46_232 ();
 sg13g2_fill_1 FILLER_46_250 ();
 sg13g2_decap_8 FILLER_46_261 ();
 sg13g2_decap_4 FILLER_46_268 ();
 sg13g2_fill_1 FILLER_46_272 ();
 sg13g2_fill_2 FILLER_46_315 ();
 sg13g2_fill_1 FILLER_46_317 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_fill_2 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_2 ();
 sg13g2_fill_2 FILLER_47_61 ();
 sg13g2_fill_1 FILLER_47_76 ();
 sg13g2_fill_1 FILLER_47_121 ();
 sg13g2_fill_1 FILLER_47_131 ();
 sg13g2_decap_4 FILLER_47_192 ();
 sg13g2_fill_2 FILLER_47_209 ();
 sg13g2_fill_1 FILLER_47_251 ();
 sg13g2_fill_2 FILLER_47_261 ();
 sg13g2_fill_1 FILLER_47_263 ();
 sg13g2_fill_1 FILLER_47_309 ();
 sg13g2_fill_1 FILLER_47_358 ();
 sg13g2_fill_1 FILLER_47_381 ();
 sg13g2_fill_1 FILLER_48_98 ();
 sg13g2_decap_4 FILLER_48_136 ();
 sg13g2_fill_2 FILLER_48_140 ();
 sg13g2_fill_1 FILLER_48_179 ();
 sg13g2_fill_2 FILLER_48_229 ();
 sg13g2_decap_4 FILLER_48_266 ();
 sg13g2_fill_1 FILLER_48_287 ();
 sg13g2_fill_1 FILLER_48_347 ();
 sg13g2_fill_1 FILLER_48_375 ();
 sg13g2_fill_2 FILLER_48_407 ();
 sg13g2_fill_2 FILLER_49_58 ();
 sg13g2_fill_1 FILLER_49_60 ();
 sg13g2_fill_1 FILLER_49_219 ();
 sg13g2_fill_1 FILLER_49_279 ();
 sg13g2_fill_1 FILLER_49_325 ();
 sg13g2_fill_2 FILLER_49_353 ();
 sg13g2_fill_1 FILLER_49_355 ();
 sg13g2_fill_2 FILLER_50_31 ();
 sg13g2_fill_1 FILLER_50_131 ();
 sg13g2_fill_2 FILLER_50_159 ();
 sg13g2_fill_2 FILLER_50_220 ();
 sg13g2_fill_1 FILLER_50_222 ();
 sg13g2_fill_1 FILLER_50_256 ();
 sg13g2_fill_2 FILLER_50_406 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_fill_1 FILLER_51_31 ();
 sg13g2_fill_2 FILLER_51_81 ();
 sg13g2_fill_2 FILLER_51_96 ();
 sg13g2_fill_1 FILLER_51_98 ();
 sg13g2_fill_1 FILLER_51_246 ();
 sg13g2_fill_1 FILLER_51_320 ();
 sg13g2_fill_2 FILLER_51_338 ();
 sg13g2_fill_2 FILLER_51_376 ();
 sg13g2_fill_1 FILLER_52_4 ();
 sg13g2_fill_1 FILLER_52_14 ();
 sg13g2_fill_1 FILLER_52_77 ();
 sg13g2_fill_1 FILLER_52_87 ();
 sg13g2_fill_1 FILLER_52_115 ();
 sg13g2_fill_2 FILLER_52_129 ();
 sg13g2_fill_2 FILLER_52_154 ();
 sg13g2_fill_2 FILLER_52_194 ();
 sg13g2_fill_1 FILLER_52_196 ();
 sg13g2_fill_1 FILLER_52_203 ();
 sg13g2_fill_2 FILLER_52_221 ();
 sg13g2_fill_1 FILLER_52_223 ();
 sg13g2_fill_2 FILLER_52_260 ();
 sg13g2_fill_2 FILLER_52_278 ();
 sg13g2_fill_1 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_54 ();
 sg13g2_fill_1 FILLER_53_56 ();
 sg13g2_fill_1 FILLER_53_93 ();
 sg13g2_fill_1 FILLER_53_103 ();
 sg13g2_fill_1 FILLER_53_148 ();
 sg13g2_fill_2 FILLER_53_208 ();
 sg13g2_fill_1 FILLER_53_210 ();
 sg13g2_fill_2 FILLER_53_259 ();
 sg13g2_fill_1 FILLER_53_261 ();
 sg13g2_fill_1 FILLER_53_378 ();
 sg13g2_fill_2 FILLER_54_40 ();
 sg13g2_fill_1 FILLER_54_42 ();
 sg13g2_fill_1 FILLER_54_110 ();
 sg13g2_fill_2 FILLER_54_138 ();
 sg13g2_fill_2 FILLER_54_149 ();
 sg13g2_fill_1 FILLER_54_151 ();
 sg13g2_fill_2 FILLER_54_193 ();
 sg13g2_fill_1 FILLER_54_195 ();
 sg13g2_fill_1 FILLER_54_350 ();
 sg13g2_fill_2 FILLER_54_378 ();
 sg13g2_fill_2 FILLER_54_398 ();
 sg13g2_fill_1 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_57 ();
 sg13g2_fill_1 FILLER_55_59 ();
 sg13g2_fill_1 FILLER_55_123 ();
 sg13g2_fill_2 FILLER_55_164 ();
 sg13g2_fill_1 FILLER_55_192 ();
 sg13g2_fill_2 FILLER_55_205 ();
 sg13g2_fill_2 FILLER_55_225 ();
 sg13g2_fill_1 FILLER_55_227 ();
 sg13g2_fill_1 FILLER_55_288 ();
 sg13g2_fill_2 FILLER_55_357 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_29 ();
 sg13g2_fill_1 FILLER_56_31 ();
 sg13g2_fill_1 FILLER_56_103 ();
 sg13g2_fill_2 FILLER_56_170 ();
 sg13g2_fill_2 FILLER_56_274 ();
 sg13g2_fill_2 FILLER_56_295 ();
 sg13g2_fill_1 FILLER_56_306 ();
 sg13g2_fill_1 FILLER_56_347 ();
 sg13g2_fill_2 FILLER_56_375 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_121 ();
 sg13g2_fill_2 FILLER_57_150 ();
 sg13g2_fill_1 FILLER_57_175 ();
 sg13g2_fill_1 FILLER_57_195 ();
 sg13g2_fill_1 FILLER_57_201 ();
 sg13g2_fill_1 FILLER_57_255 ();
 sg13g2_fill_2 FILLER_57_274 ();
 sg13g2_fill_1 FILLER_57_294 ();
 sg13g2_fill_2 FILLER_57_304 ();
 sg13g2_fill_1 FILLER_57_306 ();
 sg13g2_fill_2 FILLER_57_316 ();
 sg13g2_fill_1 FILLER_57_318 ();
 sg13g2_fill_2 FILLER_57_328 ();
 sg13g2_fill_2 FILLER_57_357 ();
 sg13g2_fill_1 FILLER_57_359 ();
 sg13g2_fill_2 FILLER_58_18 ();
 sg13g2_fill_1 FILLER_58_20 ();
 sg13g2_fill_2 FILLER_58_57 ();
 sg13g2_fill_2 FILLER_58_108 ();
 sg13g2_fill_1 FILLER_58_146 ();
 sg13g2_fill_2 FILLER_58_161 ();
 sg13g2_fill_1 FILLER_58_163 ();
 sg13g2_fill_1 FILLER_58_196 ();
 sg13g2_fill_2 FILLER_58_251 ();
 sg13g2_fill_2 FILLER_58_258 ();
 sg13g2_fill_1 FILLER_58_260 ();
 sg13g2_fill_2 FILLER_58_266 ();
 sg13g2_fill_1 FILLER_58_273 ();
 sg13g2_fill_2 FILLER_58_288 ();
 sg13g2_fill_1 FILLER_58_290 ();
 sg13g2_fill_2 FILLER_58_319 ();
 sg13g2_fill_1 FILLER_58_321 ();
 sg13g2_fill_2 FILLER_58_362 ();
 sg13g2_fill_1 FILLER_58_364 ();
 sg13g2_fill_1 FILLER_59_31 ();
 sg13g2_fill_1 FILLER_59_68 ();
 sg13g2_fill_1 FILLER_59_100 ();
 sg13g2_fill_1 FILLER_59_114 ();
 sg13g2_fill_2 FILLER_59_128 ();
 sg13g2_fill_1 FILLER_59_130 ();
 sg13g2_fill_2 FILLER_59_149 ();
 sg13g2_fill_1 FILLER_59_151 ();
 sg13g2_fill_1 FILLER_59_239 ();
 sg13g2_fill_2 FILLER_59_267 ();
 sg13g2_fill_1 FILLER_59_287 ();
 sg13g2_fill_2 FILLER_59_302 ();
 sg13g2_fill_1 FILLER_59_374 ();
 sg13g2_fill_2 FILLER_59_406 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_fill_1 FILLER_60_31 ();
 sg13g2_fill_2 FILLER_60_81 ();
 sg13g2_fill_2 FILLER_60_119 ();
 sg13g2_fill_1 FILLER_60_121 ();
 sg13g2_fill_2 FILLER_60_158 ();
 sg13g2_fill_2 FILLER_60_169 ();
 sg13g2_fill_1 FILLER_60_171 ();
 sg13g2_fill_1 FILLER_60_189 ();
 sg13g2_fill_2 FILLER_60_217 ();
 sg13g2_fill_2 FILLER_60_228 ();
 sg13g2_fill_1 FILLER_60_238 ();
 sg13g2_fill_2 FILLER_60_297 ();
 sg13g2_fill_2 FILLER_60_339 ();
 sg13g2_fill_1 FILLER_60_399 ();
 sg13g2_fill_1 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_32 ();
 sg13g2_fill_2 FILLER_61_64 ();
 sg13g2_fill_1 FILLER_61_66 ();
 sg13g2_fill_2 FILLER_61_186 ();
 sg13g2_fill_1 FILLER_61_188 ();
 sg13g2_fill_2 FILLER_61_198 ();
 sg13g2_fill_2 FILLER_61_286 ();
 sg13g2_fill_1 FILLER_61_288 ();
 sg13g2_fill_1 FILLER_61_310 ();
 sg13g2_fill_2 FILLER_61_348 ();
 sg13g2_fill_1 FILLER_61_350 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_2 ();
 sg13g2_fill_1 FILLER_62_57 ();
 sg13g2_fill_2 FILLER_62_134 ();
 sg13g2_fill_1 FILLER_62_190 ();
 sg13g2_fill_2 FILLER_62_199 ();
 sg13g2_fill_1 FILLER_62_209 ();
 sg13g2_fill_2 FILLER_62_285 ();
 sg13g2_fill_1 FILLER_62_300 ();
 sg13g2_fill_1 FILLER_62_315 ();
 sg13g2_fill_2 FILLER_62_334 ();
 sg13g2_fill_2 FILLER_62_345 ();
 sg13g2_fill_2 FILLER_63_0 ();
 sg13g2_fill_2 FILLER_63_33 ();
 sg13g2_fill_2 FILLER_63_146 ();
 sg13g2_fill_1 FILLER_63_148 ();
 sg13g2_fill_2 FILLER_63_212 ();
 sg13g2_fill_2 FILLER_63_223 ();
 sg13g2_fill_2 FILLER_63_262 ();
 sg13g2_fill_2 FILLER_63_313 ();
 sg13g2_fill_2 FILLER_63_333 ();
 sg13g2_fill_2 FILLER_63_344 ();
 sg13g2_fill_1 FILLER_63_346 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_2 ();
 sg13g2_fill_2 FILLER_64_140 ();
 sg13g2_fill_2 FILLER_64_164 ();
 sg13g2_fill_2 FILLER_64_188 ();
 sg13g2_fill_1 FILLER_64_218 ();
 sg13g2_fill_1 FILLER_64_322 ();
 sg13g2_fill_2 FILLER_64_359 ();
 sg13g2_fill_2 FILLER_65_36 ();
 sg13g2_fill_1 FILLER_65_38 ();
 sg13g2_fill_2 FILLER_65_66 ();
 sg13g2_fill_2 FILLER_65_104 ();
 sg13g2_fill_1 FILLER_65_106 ();
 sg13g2_fill_1 FILLER_65_169 ();
 sg13g2_fill_2 FILLER_65_188 ();
 sg13g2_fill_1 FILLER_65_190 ();
 sg13g2_fill_2 FILLER_65_196 ();
 sg13g2_fill_2 FILLER_65_239 ();
 sg13g2_fill_2 FILLER_65_275 ();
 sg13g2_fill_1 FILLER_65_290 ();
 sg13g2_fill_1 FILLER_65_309 ();
 sg13g2_fill_2 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_149 ();
 sg13g2_fill_1 FILLER_66_151 ();
 sg13g2_fill_1 FILLER_66_187 ();
 sg13g2_fill_2 FILLER_66_209 ();
 sg13g2_fill_2 FILLER_66_231 ();
 sg13g2_fill_2 FILLER_66_383 ();
 sg13g2_fill_2 FILLER_66_398 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_2 ();
 sg13g2_fill_2 FILLER_67_34 ();
 sg13g2_fill_1 FILLER_67_36 ();
 sg13g2_fill_1 FILLER_67_64 ();
 sg13g2_fill_1 FILLER_67_194 ();
 sg13g2_fill_2 FILLER_67_223 ();
 sg13g2_fill_2 FILLER_67_258 ();
 sg13g2_fill_1 FILLER_67_283 ();
 sg13g2_fill_1 FILLER_67_356 ();
 sg13g2_fill_2 FILLER_67_406 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_fill_2 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_2 ();
 sg13g2_fill_2 FILLER_68_34 ();
 sg13g2_fill_1 FILLER_68_72 ();
 sg13g2_fill_2 FILLER_68_122 ();
 sg13g2_fill_1 FILLER_68_269 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_fill_1 FILLER_69_53 ();
 sg13g2_fill_2 FILLER_69_90 ();
 sg13g2_fill_1 FILLER_69_92 ();
 sg13g2_fill_1 FILLER_69_155 ();
 sg13g2_fill_2 FILLER_69_307 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_fill_2 FILLER_70_106 ();
 sg13g2_fill_1 FILLER_70_108 ();
 sg13g2_fill_2 FILLER_70_127 ();
 sg13g2_fill_2 FILLER_70_199 ();
 sg13g2_fill_2 FILLER_70_288 ();
 sg13g2_fill_2 FILLER_71_31 ();
 sg13g2_fill_1 FILLER_71_33 ();
 sg13g2_fill_1 FILLER_71_74 ();
 sg13g2_fill_2 FILLER_71_132 ();
 sg13g2_fill_1 FILLER_71_134 ();
 sg13g2_fill_1 FILLER_71_175 ();
 sg13g2_fill_2 FILLER_71_241 ();
 sg13g2_fill_1 FILLER_71_252 ();
 sg13g2_fill_2 FILLER_71_276 ();
 sg13g2_fill_2 FILLER_71_322 ();
 sg13g2_fill_1 FILLER_72_0 ();
 sg13g2_fill_1 FILLER_72_295 ();
 sg13g2_fill_1 FILLER_72_324 ();
 sg13g2_fill_2 FILLER_72_364 ();
 sg13g2_fill_2 FILLER_73_49 ();
 sg13g2_fill_1 FILLER_73_123 ();
 sg13g2_fill_1 FILLER_73_151 ();
 sg13g2_fill_1 FILLER_73_221 ();
 sg13g2_fill_1 FILLER_73_239 ();
 sg13g2_fill_2 FILLER_73_302 ();
 sg13g2_fill_2 FILLER_73_407 ();
 sg13g2_fill_2 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_29 ();
 sg13g2_fill_2 FILLER_74_136 ();
 sg13g2_fill_2 FILLER_74_169 ();
 sg13g2_fill_1 FILLER_74_171 ();
 sg13g2_fill_2 FILLER_74_190 ();
 sg13g2_fill_1 FILLER_74_311 ();
 sg13g2_fill_2 FILLER_74_325 ();
 sg13g2_fill_2 FILLER_74_380 ();
 sg13g2_fill_2 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_2 ();
 sg13g2_fill_2 FILLER_75_106 ();
 sg13g2_fill_1 FILLER_75_108 ();
 sg13g2_fill_1 FILLER_75_127 ();
 sg13g2_fill_2 FILLER_75_155 ();
 sg13g2_fill_1 FILLER_75_184 ();
 sg13g2_fill_2 FILLER_75_194 ();
 sg13g2_fill_1 FILLER_75_331 ();
 sg13g2_fill_2 FILLER_75_380 ();
 sg13g2_fill_2 FILLER_76_13 ();
 sg13g2_fill_2 FILLER_76_46 ();
 sg13g2_fill_1 FILLER_76_48 ();
 sg13g2_fill_2 FILLER_76_154 ();
 sg13g2_fill_1 FILLER_76_156 ();
 sg13g2_fill_1 FILLER_76_197 ();
 sg13g2_fill_1 FILLER_76_239 ();
 sg13g2_fill_1 FILLER_76_340 ();
 sg13g2_fill_1 FILLER_76_377 ();
 sg13g2_fill_1 FILLER_77_0 ();
 sg13g2_fill_2 FILLER_77_131 ();
 sg13g2_fill_2 FILLER_77_182 ();
 sg13g2_fill_1 FILLER_77_184 ();
 sg13g2_fill_1 FILLER_77_285 ();
 sg13g2_fill_2 FILLER_77_372 ();
 sg13g2_fill_1 FILLER_77_399 ();
 sg13g2_fill_1 FILLER_78_0 ();
 sg13g2_fill_2 FILLER_78_32 ();
 sg13g2_fill_2 FILLER_78_97 ();
 sg13g2_fill_1 FILLER_78_99 ();
 sg13g2_fill_2 FILLER_78_185 ();
 sg13g2_fill_1 FILLER_78_187 ();
 sg13g2_fill_2 FILLER_78_288 ();
 sg13g2_fill_1 FILLER_78_301 ();
 sg13g2_fill_2 FILLER_78_389 ();
 sg13g2_fill_2 FILLER_79_0 ();
 sg13g2_fill_2 FILLER_79_15 ();
 sg13g2_fill_1 FILLER_79_17 ();
 sg13g2_fill_2 FILLER_79_113 ();
 sg13g2_fill_1 FILLER_79_115 ();
 sg13g2_fill_2 FILLER_79_243 ();
 sg13g2_fill_1 FILLER_79_272 ();
 sg13g2_fill_2 FILLER_79_281 ();
 sg13g2_fill_2 FILLER_79_287 ();
 sg13g2_fill_1 FILLER_79_289 ();
 sg13g2_fill_2 FILLER_79_337 ();
 sg13g2_fill_1 FILLER_79_343 ();
 sg13g2_fill_2 FILLER_79_364 ();
 sg13g2_fill_1 FILLER_79_394 ();
 sg13g2_fill_2 FILLER_79_407 ();
 sg13g2_fill_2 FILLER_80_0 ();
 sg13g2_fill_1 FILLER_80_2 ();
 sg13g2_fill_2 FILLER_80_7 ();
 sg13g2_fill_2 FILLER_80_145 ();
 sg13g2_fill_1 FILLER_80_156 ();
 sg13g2_fill_2 FILLER_80_206 ();
 sg13g2_fill_2 FILLER_80_231 ();
 sg13g2_fill_1 FILLER_80_233 ();
 sg13g2_fill_2 FILLER_80_243 ();
 sg13g2_fill_1 FILLER_80_284 ();
 sg13g2_fill_1 FILLER_80_289 ();
 sg13g2_fill_2 FILLER_80_302 ();
 sg13g2_fill_1 FILLER_80_304 ();
 sg13g2_decap_8 FILLER_80_392 ();
 sg13g2_decap_8 FILLER_80_399 ();
 sg13g2_fill_2 FILLER_80_406 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net668;
 assign uio_oe[1] = net669;
 assign uio_oe[2] = net670;
 assign uio_oe[3] = net8;
 assign uio_oe[4] = net9;
 assign uio_oe[5] = net10;
 assign uio_oe[6] = net11;
 assign uio_oe[7] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
endmodule
