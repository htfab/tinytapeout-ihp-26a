module tt_um_sujanreddy_synapse (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire \controller_inst.bit_cnt[0] ;
 wire \controller_inst.bit_cnt[1] ;
 wire \controller_inst.bit_cnt[2] ;
 wire \controller_inst.byte_ready ;
 wire \controller_inst.cmd_reg[0] ;
 wire \controller_inst.cmd_reg[1] ;
 wire \controller_inst.cmd_reg[2] ;
 wire \controller_inst.cmd_reg[3] ;
 wire \controller_inst.cmd_reg[4] ;
 wire \controller_inst.cmd_reg[5] ;
 wire \controller_inst.cmd_reg[6] ;
 wire \controller_inst.cmd_reg[7] ;
 wire \controller_inst.data_reg1[0] ;
 wire \controller_inst.data_reg1[1] ;
 wire \controller_inst.data_reg1[2] ;
 wire \controller_inst.data_reg1[3] ;
 wire \controller_inst.data_reg1[4] ;
 wire \controller_inst.data_reg1[5] ;
 wire \controller_inst.data_reg1[6] ;
 wire \controller_inst.data_reg1[7] ;
 wire \controller_inst.data_reg2[0] ;
 wire \controller_inst.data_reg2[1] ;
 wire \controller_inst.data_reg2[2] ;
 wire \controller_inst.data_reg2[3] ;
 wire \controller_inst.data_reg2[4] ;
 wire \controller_inst.data_reg2[5] ;
 wire \controller_inst.data_reg2[6] ;
 wire \controller_inst.data_reg2[7] ;
 wire \controller_inst.error ;
 wire \controller_inst.prog_done ;
 wire \controller_inst.pulse_counter[0] ;
 wire \controller_inst.pulse_counter[10] ;
 wire \controller_inst.pulse_counter[11] ;
 wire \controller_inst.pulse_counter[12] ;
 wire \controller_inst.pulse_counter[13] ;
 wire \controller_inst.pulse_counter[14] ;
 wire \controller_inst.pulse_counter[15] ;
 wire \controller_inst.pulse_counter[1] ;
 wire \controller_inst.pulse_counter[2] ;
 wire \controller_inst.pulse_counter[3] ;
 wire \controller_inst.pulse_counter[4] ;
 wire \controller_inst.pulse_counter[5] ;
 wire \controller_inst.pulse_counter[6] ;
 wire \controller_inst.pulse_counter[7] ;
 wire \controller_inst.pulse_counter[8] ;
 wire \controller_inst.pulse_counter[9] ;
 wire \controller_inst.pulse_width[0] ;
 wire \controller_inst.pulse_width[10] ;
 wire \controller_inst.pulse_width[11] ;
 wire \controller_inst.pulse_width[12] ;
 wire \controller_inst.pulse_width[13] ;
 wire \controller_inst.pulse_width[14] ;
 wire \controller_inst.pulse_width[15] ;
 wire \controller_inst.pulse_width[1] ;
 wire \controller_inst.pulse_width[2] ;
 wire \controller_inst.pulse_width[4] ;
 wire \controller_inst.ready ;
 wire \controller_inst.sck_d1 ;
 wire \controller_inst.sck_d2 ;
 wire \controller_inst.sck_d3 ;
 wire \controller_inst.shift_reg_in[0] ;
 wire \controller_inst.shift_reg_in[1] ;
 wire \controller_inst.shift_reg_in[2] ;
 wire \controller_inst.shift_reg_in[3] ;
 wire \controller_inst.shift_reg_in[4] ;
 wire \controller_inst.shift_reg_in[5] ;
 wire \controller_inst.shift_reg_in[6] ;
 wire \controller_inst.shift_reg_in[7] ;
 wire \controller_inst.shift_reg_out[0] ;
 wire \controller_inst.shift_reg_out[1] ;
 wire \controller_inst.shift_reg_out[2] ;
 wire \controller_inst.shift_reg_out[3] ;
 wire \controller_inst.shift_reg_out[5] ;
 wire \controller_inst.shift_reg_out[6] ;
 wire \controller_inst.shift_reg_out[7] ;
 wire \controller_inst.spi_miso ;
 wire \controller_inst.state[0] ;
 wire \controller_inst.state[1] ;
 wire \controller_inst.state[2] ;
 wire \controller_inst.state[3] ;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire clknet_0_clk;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;

 sg13g2_inv_1 _0795_ (.Y(_0010_),
    .A(net1));
 sg13g2_inv_1 _0796_ (.Y(\controller_inst.ready ),
    .A(net55));
 sg13g2_inv_2 _0797_ (.Y(_0102_),
    .A(net156));
 sg13g2_inv_1 _0798_ (.Y(_0103_),
    .A(net4));
 sg13g2_inv_1 _0799_ (.Y(_0104_),
    .A(net217));
 sg13g2_inv_1 _0800_ (.Y(_0105_),
    .A(net90));
 sg13g2_inv_1 _0801_ (.Y(_0106_),
    .A(net61));
 sg13g2_inv_1 _0802_ (.Y(_0107_),
    .A(net46));
 sg13g2_inv_1 _0803_ (.Y(_0108_),
    .A(net77));
 sg13g2_inv_1 _0804_ (.Y(_0109_),
    .A(net134));
 sg13g2_inv_1 _0805_ (.Y(_0110_),
    .A(net102));
 sg13g2_inv_1 _0806_ (.Y(_0111_),
    .A(net118));
 sg13g2_inv_1 _0807_ (.Y(_0112_),
    .A(net92));
 sg13g2_inv_1 _0808_ (.Y(_0113_),
    .A(net98));
 sg13g2_inv_1 _0809_ (.Y(_0114_),
    .A(net100));
 sg13g2_inv_1 _0810_ (.Y(_0115_),
    .A(net124));
 sg13g2_inv_1 _0811_ (.Y(_0116_),
    .A(net94));
 sg13g2_inv_1 _0812_ (.Y(_0117_),
    .A(net79));
 sg13g2_inv_1 _0813_ (.Y(_0118_),
    .A(net73));
 sg13g2_inv_2 _0814_ (.Y(_0119_),
    .A(net51));
 sg13g2_inv_1 _0815_ (.Y(_0120_),
    .A(\controller_inst.bit_cnt[2] ));
 sg13g2_inv_1 _0816_ (.Y(_0121_),
    .A(net31));
 sg13g2_inv_1 _0817_ (.Y(_0122_),
    .A(net32));
 sg13g2_inv_1 _0818_ (.Y(_0123_),
    .A(net34));
 sg13g2_inv_1 _0819_ (.Y(_0124_),
    .A(net33));
 sg13g2_inv_1 _0820_ (.Y(_0125_),
    .A(net155));
 sg13g2_nand2_1 _0821_ (.Y(_0126_),
    .A(net48),
    .B(net53));
 sg13g2_nand3_1 _0822_ (.B(net48),
    .C(net53),
    .A(net213),
    .Y(_0127_));
 sg13g2_nor2b_2 _0823_ (.A(net130),
    .B_N(net22),
    .Y(_0128_));
 sg13g2_nand2_2 _0824_ (.Y(_0129_),
    .A(net155),
    .B(_0128_));
 sg13g2_nor2_1 _0825_ (.A(_0127_),
    .B(net154),
    .Y(_0000_));
 sg13g2_nor2b_2 _0826_ (.A(\controller_inst.state[3] ),
    .B_N(\controller_inst.state[2] ),
    .Y(_0130_));
 sg13g2_inv_1 _0827_ (.Y(_0131_),
    .A(_0130_));
 sg13g2_and2_1 _0828_ (.A(\controller_inst.state[1] ),
    .B(_0130_),
    .X(_0132_));
 sg13g2_nand2_2 _0829_ (.Y(_0133_),
    .A(\controller_inst.state[1] ),
    .B(_0130_));
 sg13g2_nand2_2 _0830_ (.Y(_0134_),
    .A(net156),
    .B(_0132_));
 sg13g2_nor2_2 _0831_ (.A(\controller_inst.state[1] ),
    .B(net87),
    .Y(_0135_));
 sg13g2_nand2b_2 _0832_ (.Y(_0136_),
    .B(_0135_),
    .A_N(\controller_inst.state[3] ));
 sg13g2_nor2_2 _0833_ (.A(_0102_),
    .B(_0136_),
    .Y(_0137_));
 sg13g2_or4_1 _0834_ (.A(\controller_inst.cmd_reg[5] ),
    .B(\controller_inst.cmd_reg[4] ),
    .C(\controller_inst.cmd_reg[7] ),
    .D(\controller_inst.cmd_reg[6] ),
    .X(_0138_));
 sg13g2_nor2_1 _0835_ (.A(\controller_inst.cmd_reg[1] ),
    .B(_0138_),
    .Y(_0139_));
 sg13g2_inv_1 _0836_ (.Y(_0140_),
    .A(_0139_));
 sg13g2_nand2b_2 _0837_ (.Y(_0141_),
    .B(\controller_inst.cmd_reg[2] ),
    .A_N(\controller_inst.cmd_reg[3] ));
 sg13g2_nor3_2 _0838_ (.A(net129),
    .B(_0140_),
    .C(_0141_),
    .Y(_0142_));
 sg13g2_nor2b_1 _0839_ (.A(\controller_inst.cmd_reg[0] ),
    .B_N(\controller_inst.cmd_reg[1] ),
    .Y(_0143_));
 sg13g2_nor3_1 _0840_ (.A(\controller_inst.cmd_reg[3] ),
    .B(\controller_inst.cmd_reg[2] ),
    .C(_0138_),
    .Y(_0144_));
 sg13g2_a21o_1 _0841_ (.A2(_0144_),
    .A1(_0143_),
    .B1(_0142_),
    .X(_0145_));
 sg13g2_nand2_1 _0842_ (.Y(_0146_),
    .A(_0137_),
    .B(_0145_));
 sg13g2_nand2_1 _0843_ (.Y(_0147_),
    .A(_0134_),
    .B(_0146_));
 sg13g2_nor4_1 _0844_ (.A(\controller_inst.pulse_counter[13] ),
    .B(\controller_inst.pulse_counter[12] ),
    .C(\controller_inst.pulse_counter[15] ),
    .D(\controller_inst.pulse_counter[14] ),
    .Y(_0148_));
 sg13g2_nor4_1 _0845_ (.A(\controller_inst.pulse_counter[7] ),
    .B(\controller_inst.pulse_counter[6] ),
    .C(\controller_inst.pulse_counter[11] ),
    .D(\controller_inst.pulse_counter[10] ),
    .Y(_0149_));
 sg13g2_nor4_1 _0846_ (.A(\controller_inst.pulse_counter[3] ),
    .B(\controller_inst.pulse_counter[2] ),
    .C(\controller_inst.pulse_counter[5] ),
    .D(net46),
    .Y(_0150_));
 sg13g2_nor4_1 _0847_ (.A(_0104_),
    .B(\controller_inst.pulse_counter[1] ),
    .C(\controller_inst.pulse_counter[9] ),
    .D(\controller_inst.pulse_counter[8] ),
    .Y(_0151_));
 sg13g2_nand4_1 _0848_ (.B(_0149_),
    .C(_0150_),
    .A(_0148_),
    .Y(_0152_),
    .D(_0151_));
 sg13g2_nand2b_2 _0849_ (.Y(_0153_),
    .B(_0152_),
    .A_N(_0134_));
 sg13g2_and2_1 _0850_ (.A(_0147_),
    .B(_0153_),
    .X(_0154_));
 sg13g2_nand2_2 _0851_ (.Y(_0155_),
    .A(_0134_),
    .B(_0142_));
 sg13g2_nand3_1 _0852_ (.B(net138),
    .C(_0155_),
    .A(net5),
    .Y(_0156_));
 sg13g2_o21ai_1 _0853_ (.B1(_0156_),
    .Y(_0012_),
    .A1(_0124_),
    .A2(net138));
 sg13g2_nand3_1 _0854_ (.B(net138),
    .C(_0155_),
    .A(net6),
    .Y(_0157_));
 sg13g2_o21ai_1 _0855_ (.B1(_0157_),
    .Y(_0013_),
    .A1(_0123_),
    .A2(net138));
 sg13g2_nand3_1 _0856_ (.B(net138),
    .C(_0155_),
    .A(net7),
    .Y(_0158_));
 sg13g2_o21ai_1 _0857_ (.B1(_0158_),
    .Y(_0014_),
    .A1(_0122_),
    .A2(_0154_));
 sg13g2_nand3_1 _0858_ (.B(_0154_),
    .C(_0155_),
    .A(net8),
    .Y(_0159_));
 sg13g2_o21ai_1 _0859_ (.B1(_0159_),
    .Y(_0015_),
    .A1(_0121_),
    .A2(_0154_));
 sg13g2_nor2_1 _0860_ (.A(_0118_),
    .B(_0155_),
    .Y(_0160_));
 sg13g2_mux2_1 _0861_ (.A0(net41),
    .A1(_0160_),
    .S(net138),
    .X(_0016_));
 sg13g2_and3_1 _0862_ (.X(_0161_),
    .A(\controller_inst.error ),
    .B(_0134_),
    .C(_0142_));
 sg13g2_mux2_1 _0863_ (.A0(net63),
    .A1(_0161_),
    .S(net138),
    .X(_0017_));
 sg13g2_nor2_1 _0864_ (.A(net55),
    .B(_0155_),
    .Y(_0162_));
 sg13g2_mux2_1 _0865_ (.A0(net43),
    .A1(_0162_),
    .S(net138),
    .X(_0018_));
 sg13g2_nand2_1 _0866_ (.Y(_0163_),
    .A(\controller_inst.cmd_reg[0] ),
    .B(_0139_));
 sg13g2_nor3_1 _0867_ (.A(\controller_inst.cmd_reg[3] ),
    .B(\controller_inst.cmd_reg[2] ),
    .C(_0163_),
    .Y(_0164_));
 sg13g2_nor2_1 _0868_ (.A(_0138_),
    .B(_0141_),
    .Y(_0165_));
 sg13g2_nand3_1 _0869_ (.B(\controller_inst.cmd_reg[0] ),
    .C(_0165_),
    .A(\controller_inst.cmd_reg[1] ),
    .Y(_0166_));
 sg13g2_inv_1 _0870_ (.Y(_0167_),
    .A(_0166_));
 sg13g2_nand2b_1 _0871_ (.Y(_0168_),
    .B(_0166_),
    .A_N(_0164_));
 sg13g2_nand2_2 _0872_ (.Y(_0169_),
    .A(_0143_),
    .B(_0165_));
 sg13g2_nand3_1 _0873_ (.B(\controller_inst.cmd_reg[0] ),
    .C(_0144_),
    .A(\controller_inst.cmd_reg[1] ),
    .Y(_0170_));
 sg13g2_o21ai_1 _0874_ (.B1(_0170_),
    .Y(_0171_),
    .A1(_0141_),
    .A2(_0163_));
 sg13g2_nor2_1 _0875_ (.A(_0168_),
    .B(_0171_),
    .Y(_0172_));
 sg13g2_nand2_1 _0876_ (.Y(_0173_),
    .A(net120),
    .B(_0137_));
 sg13g2_a221oi_1 _0877_ (.B2(_0169_),
    .C1(_0173_),
    .B1(_0172_),
    .A1(_0103_),
    .Y(_0174_),
    .A2(_0171_));
 sg13g2_mux2_1 _0878_ (.A0(net25),
    .A1(net108),
    .S(net145),
    .X(_0019_));
 sg13g2_mux2_1 _0879_ (.A0(net27),
    .A1(net131),
    .S(net145),
    .X(_0020_));
 sg13g2_mux2_1 _0880_ (.A0(net116),
    .A1(net121),
    .S(_0174_),
    .X(_0021_));
 sg13g2_mux2_1 _0881_ (.A0(net112),
    .A1(net37),
    .S(net145),
    .X(_0022_));
 sg13g2_mux2_1 _0882_ (.A0(net109),
    .A1(\controller_inst.shift_reg_in[4] ),
    .S(net145),
    .X(_0023_));
 sg13g2_mux2_1 _0883_ (.A0(net185),
    .A1(net39),
    .S(net145),
    .X(_0024_));
 sg13g2_mux2_1 _0884_ (.A0(net184),
    .A1(net57),
    .S(net145),
    .X(_0025_));
 sg13g2_nand2_1 _0885_ (.Y(_0175_),
    .A(net29),
    .B(net145));
 sg13g2_o21ai_1 _0886_ (.B1(_0175_),
    .Y(_0026_),
    .A1(_0119_),
    .A2(net145));
 sg13g2_nand2b_2 _0887_ (.Y(_0176_),
    .B(net155),
    .A_N(_0128_));
 sg13g2_a21oi_1 _0888_ (.A1(net155),
    .A2(_0128_),
    .Y(_0177_),
    .B1(net53));
 sg13g2_a21oi_1 _0889_ (.A1(net53),
    .A2(_0176_),
    .Y(_0027_),
    .B1(_0177_));
 sg13g2_a21oi_1 _0890_ (.A1(\controller_inst.bit_cnt[0] ),
    .A2(_0176_),
    .Y(_0178_),
    .B1(net48));
 sg13g2_nand2_1 _0891_ (.Y(_0179_),
    .A(_0009_),
    .B(_0126_));
 sg13g2_a21oi_1 _0892_ (.A1(_0176_),
    .A2(_0179_),
    .Y(_0028_),
    .B1(net49));
 sg13g2_nand2b_1 _0893_ (.Y(_0180_),
    .B(_0176_),
    .A_N(_0126_));
 sg13g2_nand2_1 _0894_ (.Y(_0181_),
    .A(net67),
    .B(_0127_));
 sg13g2_a22oi_1 _0895_ (.Y(_0029_),
    .B1(net68),
    .B2(_0176_),
    .A2(_0180_),
    .A1(_0120_));
 sg13g2_nor2_1 _0896_ (.A(\controller_inst.pulse_counter[0] ),
    .B(\controller_inst.pulse_counter[1] ),
    .Y(_0182_));
 sg13g2_nor3_1 _0897_ (.A(\controller_inst.pulse_counter[0] ),
    .B(net90),
    .C(\controller_inst.pulse_counter[2] ),
    .Y(_0183_));
 sg13g2_nand2b_1 _0898_ (.Y(_0184_),
    .B(_0183_),
    .A_N(\controller_inst.pulse_counter[3] ));
 sg13g2_nand2_1 _0899_ (.Y(_0185_),
    .A(_0150_),
    .B(_0182_));
 sg13g2_nand4_1 _0900_ (.B(_0109_),
    .C(_0150_),
    .A(_0108_),
    .Y(_0186_),
    .D(_0182_));
 sg13g2_nand3b_1 _0901_ (.B(_0111_),
    .C(_0110_),
    .Y(_0187_),
    .A_N(_0186_));
 sg13g2_nor3_2 _0902_ (.A(net92),
    .B(net98),
    .C(_0187_),
    .Y(_0188_));
 sg13g2_inv_1 _0903_ (.Y(_0189_),
    .A(_0188_));
 sg13g2_nand2_2 _0904_ (.Y(_0190_),
    .A(_0115_),
    .B(_0188_));
 sg13g2_nor3_1 _0905_ (.A(\controller_inst.pulse_counter[13] ),
    .B(net79),
    .C(_0190_),
    .Y(_0191_));
 sg13g2_and2_1 _0906_ (.A(_0148_),
    .B(_0188_),
    .X(_0192_));
 sg13g2_nor2_2 _0907_ (.A(net156),
    .B(\controller_inst.state[3] ),
    .Y(_0193_));
 sg13g2_nand2_1 _0908_ (.Y(_0194_),
    .A(net221),
    .B(_0193_));
 sg13g2_nor2_1 _0909_ (.A(net156),
    .B(_0133_),
    .Y(_0195_));
 sg13g2_nand2_1 _0910_ (.Y(_0196_),
    .A(_0192_),
    .B(_0195_));
 sg13g2_nor3_2 _0911_ (.A(_0102_),
    .B(\controller_inst.state[1] ),
    .C(_0131_),
    .Y(_0197_));
 sg13g2_o21ai_1 _0912_ (.B1(_0196_),
    .Y(_0030_),
    .A1(_0118_),
    .A2(_0197_));
 sg13g2_mux2_1 _0913_ (.A0(net3),
    .A1(net108),
    .S(_0129_),
    .X(_0031_));
 sg13g2_mux2_1 _0914_ (.A0(net108),
    .A1(net131),
    .S(net154),
    .X(_0032_));
 sg13g2_mux2_1 _0915_ (.A0(net131),
    .A1(net121),
    .S(net154),
    .X(_0033_));
 sg13g2_mux2_1 _0916_ (.A0(net121),
    .A1(net37),
    .S(net154),
    .X(_0034_));
 sg13g2_mux2_1 _0917_ (.A0(net37),
    .A1(net205),
    .S(net154),
    .X(_0035_));
 sg13g2_mux2_1 _0918_ (.A0(net205),
    .A1(net39),
    .S(net154),
    .X(_0036_));
 sg13g2_mux2_1 _0919_ (.A0(net39),
    .A1(net57),
    .S(net154),
    .X(_0037_));
 sg13g2_mux2_1 _0920_ (.A0(net57),
    .A1(net29),
    .S(net154),
    .X(_0038_));
 sg13g2_or2_1 _0921_ (.X(_0198_),
    .B(_0170_),
    .A(_0103_));
 sg13g2_nand3_1 _0922_ (.B(_0169_),
    .C(_0198_),
    .A(_0166_),
    .Y(_0199_));
 sg13g2_nor3_1 _0923_ (.A(_0103_),
    .B(_0141_),
    .C(_0163_),
    .Y(_0200_));
 sg13g2_or2_1 _0924_ (.X(_0201_),
    .B(_0200_),
    .A(_0168_));
 sg13g2_nor4_1 _0925_ (.A(\controller_inst.cmd_reg[0] ),
    .B(\controller_inst.cmd_reg[3] ),
    .C(\controller_inst.cmd_reg[2] ),
    .D(_0140_),
    .Y(_0202_));
 sg13g2_nand2b_1 _0926_ (.Y(_0203_),
    .B(_0137_),
    .A_N(_0202_));
 sg13g2_nor4_1 _0927_ (.A(_0145_),
    .B(_0199_),
    .C(_0201_),
    .D(_0203_),
    .Y(_0204_));
 sg13g2_nor2_1 _0928_ (.A(\controller_inst.error ),
    .B(_0204_),
    .Y(_0205_));
 sg13g2_a21oi_1 _0929_ (.A1(net23),
    .A2(_0125_),
    .Y(_0039_),
    .B1(_0205_));
 sg13g2_nor2b_1 _0930_ (.A(_0192_),
    .B_N(_0195_),
    .Y(_0206_));
 sg13g2_nand4_1 _0931_ (.B(net202),
    .C(net155),
    .A(_0102_),
    .Y(_0207_),
    .D(_0135_));
 sg13g2_nor2_1 _0932_ (.A(net87),
    .B(_0194_),
    .Y(_0208_));
 sg13g2_nand2b_1 _0933_ (.Y(_0209_),
    .B(_0208_),
    .A_N(\controller_inst.byte_ready ));
 sg13g2_nand3b_1 _0934_ (.B(_0207_),
    .C(_0209_),
    .Y(_0210_),
    .A_N(_0206_));
 sg13g2_nor4_1 _0935_ (.A(net156),
    .B(\controller_inst.state[1] ),
    .C(_0131_),
    .D(_0164_),
    .Y(_0211_));
 sg13g2_nand2_1 _0936_ (.Y(_0212_),
    .A(_0169_),
    .B(_0208_));
 sg13g2_a21oi_1 _0937_ (.A1(_0102_),
    .A2(_0135_),
    .Y(_0213_),
    .B1(_0193_));
 sg13g2_nand2_1 _0938_ (.Y(_0214_),
    .A(_0136_),
    .B(_0213_));
 sg13g2_nand2_1 _0939_ (.Y(_0215_),
    .A(_0212_),
    .B(_0214_));
 sg13g2_nor3_1 _0940_ (.A(_0210_),
    .B(_0211_),
    .C(_0215_),
    .Y(_0216_));
 sg13g2_o21ai_1 _0941_ (.B1(_0203_),
    .Y(_0040_),
    .A1(\controller_inst.ready ),
    .A2(_0216_));
 sg13g2_and3_2 _0942_ (.X(_0217_),
    .A(net156),
    .B(\controller_inst.state[3] ),
    .C(_0135_));
 sg13g2_nand3_1 _0943_ (.B(\controller_inst.state[3] ),
    .C(_0135_),
    .A(net156),
    .Y(_0218_));
 sg13g2_nor2_2 _0944_ (.A(_0197_),
    .B(_0217_),
    .Y(_0219_));
 sg13g2_nor2_2 _0945_ (.A(_0132_),
    .B(_0217_),
    .Y(_0220_));
 sg13g2_nand2_2 _0946_ (.Y(_0221_),
    .A(_0133_),
    .B(_0218_));
 sg13g2_nor2_1 _0947_ (.A(_0197_),
    .B(_0221_),
    .Y(_0222_));
 sg13g2_nand2_2 _0948_ (.Y(_0223_),
    .A(_0133_),
    .B(_0219_));
 sg13g2_nand2_2 _0949_ (.Y(_0224_),
    .A(_0196_),
    .B(_0223_));
 sg13g2_a21o_2 _0950_ (.A2(_0192_),
    .A1(\controller_inst.state[0] ),
    .B1(_0133_),
    .X(_0225_));
 sg13g2_a21oi_2 _0951_ (.B1(_0133_),
    .Y(_0226_),
    .A2(_0192_),
    .A1(\controller_inst.state[0] ));
 sg13g2_nand2_1 _0952_ (.Y(_0227_),
    .A(_0104_),
    .B(_0226_));
 sg13g2_nand3_1 _0953_ (.B(net215),
    .C(net153),
    .A(net172),
    .Y(_0228_));
 sg13g2_nor2b_1 _0954_ (.A(net143),
    .B_N(_0228_),
    .Y(_0229_));
 sg13g2_a22oi_1 _0955_ (.Y(_0041_),
    .B1(_0227_),
    .B2(_0229_),
    .A2(net144),
    .A1(_0104_));
 sg13g2_xnor2_1 _0956_ (.Y(_0230_),
    .A(\controller_inst.pulse_counter[0] ),
    .B(net90));
 sg13g2_and4_1 _0957_ (.A(net172),
    .B(\controller_inst.pulse_width[0] ),
    .C(net181),
    .D(net169),
    .X(_0231_));
 sg13g2_a22oi_1 _0958_ (.Y(_0232_),
    .B1(net168),
    .B2(\controller_inst.pulse_width[0] ),
    .A2(net181),
    .A1(net173));
 sg13g2_nor2_1 _0959_ (.A(_0231_),
    .B(_0232_),
    .Y(_0233_));
 sg13g2_a221oi_1 _0960_ (.B2(net153),
    .C1(net143),
    .B1(_0233_),
    .A1(_0132_),
    .Y(_0234_),
    .A2(_0230_));
 sg13g2_a21oi_1 _0961_ (.A1(_0105_),
    .A2(net143),
    .Y(_0042_),
    .B1(_0234_));
 sg13g2_xnor2_1 _0962_ (.Y(_0235_),
    .A(net122),
    .B(_0182_));
 sg13g2_nand2_1 _0963_ (.Y(_0236_),
    .A(net183),
    .B(net166));
 sg13g2_and2_1 _0964_ (.A(net173),
    .B(net180),
    .X(_0237_));
 sg13g2_nand2_1 _0965_ (.Y(_0238_),
    .A(net182),
    .B(net169));
 sg13g2_nand3_1 _0966_ (.B(net169),
    .C(_0237_),
    .A(net182),
    .Y(_0239_));
 sg13g2_xor2_1 _0967_ (.B(_0238_),
    .A(_0237_),
    .X(_0240_));
 sg13g2_xor2_1 _0968_ (.B(_0240_),
    .A(_0236_),
    .X(_0241_));
 sg13g2_and2_1 _0969_ (.A(_0231_),
    .B(_0241_),
    .X(_0242_));
 sg13g2_o21ai_1 _0970_ (.B1(_0220_),
    .Y(_0243_),
    .A1(_0231_),
    .A2(_0241_));
 sg13g2_or2_1 _0971_ (.X(_0244_),
    .B(_0243_),
    .A(_0242_));
 sg13g2_o21ai_1 _0972_ (.B1(_0244_),
    .Y(_0245_),
    .A1(_0225_),
    .A2(_0235_));
 sg13g2_mux2_1 _0973_ (.A0(_0245_),
    .A1(net122),
    .S(net143),
    .X(_0043_));
 sg13g2_xnor2_1 _0974_ (.Y(_0246_),
    .A(net96),
    .B(_0183_));
 sg13g2_nand2_1 _0975_ (.Y(_0247_),
    .A(net183),
    .B(net163));
 sg13g2_o21ai_1 _0976_ (.B1(_0239_),
    .Y(_0248_),
    .A1(_0236_),
    .A2(_0240_));
 sg13g2_nand2_1 _0977_ (.Y(_0249_),
    .A(net182),
    .B(net166));
 sg13g2_nor2b_2 _0978_ (.A(net179),
    .B_N(net168),
    .Y(_0250_));
 sg13g2_nor2b_1 _0979_ (.A(net179),
    .B_N(net172),
    .Y(_0251_));
 sg13g2_nand2_1 _0980_ (.Y(_0252_),
    .A(_0237_),
    .B(_0250_));
 sg13g2_a21oi_1 _0981_ (.A1(net169),
    .A2(net180),
    .Y(_0253_),
    .B1(_0251_));
 sg13g2_a21oi_1 _0982_ (.A1(_0237_),
    .A2(_0250_),
    .Y(_0254_),
    .B1(_0253_));
 sg13g2_xnor2_1 _0983_ (.Y(_0255_),
    .A(_0249_),
    .B(_0254_));
 sg13g2_nand2_1 _0984_ (.Y(_0256_),
    .A(_0248_),
    .B(_0255_));
 sg13g2_xnor2_1 _0985_ (.Y(_0257_),
    .A(_0248_),
    .B(_0255_));
 sg13g2_xor2_1 _0986_ (.B(_0257_),
    .A(_0247_),
    .X(_0258_));
 sg13g2_nand2_1 _0987_ (.Y(_0259_),
    .A(_0242_),
    .B(_0258_));
 sg13g2_xnor2_1 _0988_ (.Y(_0260_),
    .A(_0242_),
    .B(_0258_));
 sg13g2_a221oi_1 _0989_ (.B2(net153),
    .C1(net143),
    .B1(_0260_),
    .A1(_0132_),
    .Y(_0261_),
    .A2(_0246_));
 sg13g2_a21o_1 _0990_ (.A2(net143),
    .A1(net96),
    .B1(_0261_),
    .X(_0044_));
 sg13g2_xnor2_1 _0991_ (.Y(_0262_),
    .A(net46),
    .B(_0184_));
 sg13g2_a22oi_1 _0992_ (.Y(_0263_),
    .B1(net161),
    .B2(net183),
    .A2(net163),
    .A1(net182));
 sg13g2_nand4_1 _0993_ (.B(net181),
    .C(net163),
    .A(net183),
    .Y(_0264_),
    .D(net161));
 sg13g2_nand2b_1 _0994_ (.Y(_0265_),
    .B(_0264_),
    .A_N(_0263_));
 sg13g2_o21ai_1 _0995_ (.B1(_0252_),
    .Y(_0266_),
    .A1(_0249_),
    .A2(_0253_));
 sg13g2_nand2_1 _0996_ (.Y(_0267_),
    .A(net180),
    .B(net166));
 sg13g2_nand2_1 _0997_ (.Y(_0268_),
    .A(net168),
    .B(\controller_inst.pulse_width[4] ));
 sg13g2_nand2_1 _0998_ (.Y(_0269_),
    .A(net172),
    .B(\controller_inst.pulse_width[4] ));
 sg13g2_nand3_1 _0999_ (.B(net178),
    .C(_0251_),
    .A(net168),
    .Y(_0270_));
 sg13g2_nor2b_1 _1000_ (.A(_0250_),
    .B_N(_0269_),
    .Y(_0271_));
 sg13g2_xnor2_1 _1001_ (.Y(_0272_),
    .A(_0250_),
    .B(_0269_));
 sg13g2_xnor2_1 _1002_ (.Y(_0273_),
    .A(_0267_),
    .B(_0272_));
 sg13g2_nand2_1 _1003_ (.Y(_0274_),
    .A(_0266_),
    .B(_0273_));
 sg13g2_xnor2_1 _1004_ (.Y(_0275_),
    .A(_0266_),
    .B(_0273_));
 sg13g2_xor2_1 _1005_ (.B(_0275_),
    .A(_0265_),
    .X(_0276_));
 sg13g2_o21ai_1 _1006_ (.B1(_0256_),
    .Y(_0277_),
    .A1(_0247_),
    .A2(_0257_));
 sg13g2_nand2_1 _1007_ (.Y(_0278_),
    .A(_0276_),
    .B(_0277_));
 sg13g2_xnor2_1 _1008_ (.Y(_0279_),
    .A(_0276_),
    .B(_0277_));
 sg13g2_or2_1 _1009_ (.X(_0280_),
    .B(_0279_),
    .A(_0259_));
 sg13g2_a21oi_1 _1010_ (.A1(_0259_),
    .A2(_0279_),
    .Y(_0281_),
    .B1(_0221_));
 sg13g2_a221oi_1 _1011_ (.B2(_0281_),
    .C1(net143),
    .B1(_0280_),
    .A1(_0226_),
    .Y(_0282_),
    .A2(_0262_));
 sg13g2_a21oi_1 _1012_ (.A1(_0107_),
    .A2(net144),
    .Y(_0045_),
    .B1(_0282_));
 sg13g2_o21ai_1 _1013_ (.B1(_0274_),
    .Y(_0283_),
    .A1(_0265_),
    .A2(_0275_));
 sg13g2_nand2_1 _1014_ (.Y(_0284_),
    .A(net183),
    .B(net159));
 sg13g2_nand2_1 _1015_ (.Y(_0285_),
    .A(net180),
    .B(net161));
 sg13g2_and4_1 _1016_ (.A(net181),
    .B(\controller_inst.pulse_width[2] ),
    .C(net163),
    .D(net161),
    .X(_0286_));
 sg13g2_a22oi_1 _1017_ (.Y(_0287_),
    .B1(net161),
    .B2(net181),
    .A2(net163),
    .A1(\controller_inst.pulse_width[2] ));
 sg13g2_nor3_1 _1018_ (.A(_0284_),
    .B(_0286_),
    .C(_0287_),
    .Y(_0288_));
 sg13g2_o21ai_1 _1019_ (.B1(_0284_),
    .Y(_0289_),
    .A1(_0286_),
    .A2(_0287_));
 sg13g2_nor2b_1 _1020_ (.A(_0288_),
    .B_N(_0289_),
    .Y(_0290_));
 sg13g2_o21ai_1 _1021_ (.B1(_0270_),
    .Y(_0291_),
    .A1(_0267_),
    .A2(_0271_));
 sg13g2_nor2b_1 _1022_ (.A(net179),
    .B_N(net166),
    .Y(_0292_));
 sg13g2_nor2b_1 _1023_ (.A(net177),
    .B_N(net168),
    .Y(_0293_));
 sg13g2_nand2b_1 _1024_ (.Y(_0294_),
    .B(net168),
    .A_N(net177));
 sg13g2_nor2b_1 _1025_ (.A(_0003_),
    .B_N(net173),
    .Y(_0295_));
 sg13g2_nor2_1 _1026_ (.A(_0269_),
    .B(_0294_),
    .Y(_0296_));
 sg13g2_xnor2_1 _1027_ (.Y(_0297_),
    .A(_0268_),
    .B(_0295_));
 sg13g2_xor2_1 _1028_ (.B(_0297_),
    .A(_0292_),
    .X(_0298_));
 sg13g2_and2_1 _1029_ (.A(_0291_),
    .B(_0298_),
    .X(_0299_));
 sg13g2_xor2_1 _1030_ (.B(_0298_),
    .A(_0291_),
    .X(_0300_));
 sg13g2_xnor2_1 _1031_ (.Y(_0301_),
    .A(_0290_),
    .B(_0300_));
 sg13g2_nand2b_1 _1032_ (.Y(_0302_),
    .B(_0283_),
    .A_N(_0301_));
 sg13g2_xor2_1 _1033_ (.B(_0301_),
    .A(_0283_),
    .X(_0303_));
 sg13g2_xor2_1 _1034_ (.B(_0303_),
    .A(_0264_),
    .X(_0304_));
 sg13g2_nand2b_1 _1035_ (.Y(_0305_),
    .B(_0304_),
    .A_N(_0278_));
 sg13g2_xor2_1 _1036_ (.B(_0304_),
    .A(_0278_),
    .X(_0306_));
 sg13g2_or2_1 _1037_ (.X(_0307_),
    .B(_0306_),
    .A(_0280_));
 sg13g2_a21oi_1 _1038_ (.A1(_0280_),
    .A2(_0306_),
    .Y(_0308_),
    .B1(_0221_));
 sg13g2_o21ai_1 _1039_ (.B1(net61),
    .Y(_0309_),
    .A1(net46),
    .A2(_0184_));
 sg13g2_a21o_1 _1040_ (.A2(_0309_),
    .A1(_0185_),
    .B1(_0225_),
    .X(_0310_));
 sg13g2_a21oi_1 _1041_ (.A1(_0307_),
    .A2(_0308_),
    .Y(_0311_),
    .B1(net143));
 sg13g2_a22oi_1 _1042_ (.Y(_0046_),
    .B1(_0310_),
    .B2(_0311_),
    .A2(net144),
    .A1(_0106_));
 sg13g2_o21ai_1 _1043_ (.B1(_0302_),
    .Y(_0312_),
    .A1(_0264_),
    .A2(_0303_));
 sg13g2_or2_1 _1044_ (.X(_0313_),
    .B(_0288_),
    .A(_0286_));
 sg13g2_nand2_1 _1045_ (.Y(_0314_),
    .A(net183),
    .B(net158));
 sg13g2_nand2b_1 _1046_ (.Y(_0315_),
    .B(_0313_),
    .A_N(_0314_));
 sg13g2_inv_1 _1047_ (.Y(_0316_),
    .A(_0315_));
 sg13g2_xnor2_1 _1048_ (.Y(_0317_),
    .A(_0313_),
    .B(_0314_));
 sg13g2_a21oi_1 _1049_ (.A1(_0290_),
    .A2(_0300_),
    .Y(_0318_),
    .B1(_0299_));
 sg13g2_nand2_1 _1050_ (.Y(_0319_),
    .A(net181),
    .B(net159));
 sg13g2_nand2b_1 _1051_ (.Y(_0320_),
    .B(net162),
    .A_N(net179));
 sg13g2_nand2b_1 _1052_ (.Y(_0321_),
    .B(\controller_inst.data_reg2[3] ),
    .A_N(_0002_));
 sg13g2_xor2_1 _1053_ (.B(_0321_),
    .A(_0285_),
    .X(_0322_));
 sg13g2_nand2b_1 _1054_ (.Y(_0323_),
    .B(_0322_),
    .A_N(_0319_));
 sg13g2_xnor2_1 _1055_ (.Y(_0324_),
    .A(_0319_),
    .B(_0322_));
 sg13g2_a21oi_1 _1056_ (.A1(_0292_),
    .A2(_0297_),
    .Y(_0325_),
    .B1(_0296_));
 sg13g2_nand2_1 _1057_ (.Y(_0326_),
    .A(net166),
    .B(net178));
 sg13g2_nand2b_1 _1058_ (.Y(_0327_),
    .B(net168),
    .A_N(net176));
 sg13g2_nor2b_2 _1059_ (.A(net176),
    .B_N(net171),
    .Y(_0328_));
 sg13g2_nand2_1 _1060_ (.Y(_0329_),
    .A(_0293_),
    .B(_0328_));
 sg13g2_nor2_1 _1061_ (.A(_0293_),
    .B(_0328_),
    .Y(_0330_));
 sg13g2_xnor2_1 _1062_ (.Y(_0331_),
    .A(_0294_),
    .B(_0328_));
 sg13g2_xnor2_1 _1063_ (.Y(_0332_),
    .A(_0326_),
    .B(_0331_));
 sg13g2_nor2b_1 _1064_ (.A(_0325_),
    .B_N(_0332_),
    .Y(_0333_));
 sg13g2_xnor2_1 _1065_ (.Y(_0334_),
    .A(_0325_),
    .B(_0332_));
 sg13g2_xnor2_1 _1066_ (.Y(_0335_),
    .A(_0324_),
    .B(_0334_));
 sg13g2_nor2_1 _1067_ (.A(_0318_),
    .B(_0335_),
    .Y(_0336_));
 sg13g2_xor2_1 _1068_ (.B(_0335_),
    .A(_0318_),
    .X(_0337_));
 sg13g2_xnor2_1 _1069_ (.Y(_0338_),
    .A(_0317_),
    .B(_0337_));
 sg13g2_nand2b_1 _1070_ (.Y(_0339_),
    .B(_0312_),
    .A_N(_0338_));
 sg13g2_xor2_1 _1071_ (.B(_0338_),
    .A(_0312_),
    .X(_0340_));
 sg13g2_or2_1 _1072_ (.X(_0341_),
    .B(_0340_),
    .A(_0305_));
 sg13g2_xnor2_1 _1073_ (.Y(_0342_),
    .A(_0305_),
    .B(_0340_));
 sg13g2_a21oi_1 _1074_ (.A1(_0307_),
    .A2(_0342_),
    .Y(_0343_),
    .B1(_0221_));
 sg13g2_o21ai_1 _1075_ (.B1(_0343_),
    .Y(_0344_),
    .A1(_0307_),
    .A2(_0342_));
 sg13g2_xnor2_1 _1076_ (.Y(_0345_),
    .A(net134),
    .B(_0185_));
 sg13g2_a21oi_1 _1077_ (.A1(_0226_),
    .A2(_0345_),
    .Y(_0346_),
    .B1(net144));
 sg13g2_a22oi_1 _1078_ (.Y(_0047_),
    .B1(_0344_),
    .B2(_0346_),
    .A2(net144),
    .A1(_0109_));
 sg13g2_o21ai_1 _1079_ (.B1(_0341_),
    .Y(_0347_),
    .A1(_0307_),
    .A2(_0342_));
 sg13g2_a21oi_1 _1080_ (.A1(_0317_),
    .A2(_0337_),
    .Y(_0348_),
    .B1(_0336_));
 sg13g2_nand2_1 _1081_ (.Y(_0349_),
    .A(net183),
    .B(net157));
 sg13g2_o21ai_1 _1082_ (.B1(_0323_),
    .Y(_0350_),
    .A1(_0285_),
    .A2(_0321_));
 sg13g2_nand2_1 _1083_ (.Y(_0351_),
    .A(net181),
    .B(net158));
 sg13g2_nand2b_1 _1084_ (.Y(_0352_),
    .B(_0350_),
    .A_N(_0351_));
 sg13g2_xor2_1 _1085_ (.B(_0351_),
    .A(_0350_),
    .X(_0353_));
 sg13g2_xor2_1 _1086_ (.B(_0353_),
    .A(_0349_),
    .X(_0354_));
 sg13g2_a21oi_1 _1087_ (.A1(_0324_),
    .A2(_0334_),
    .Y(_0355_),
    .B1(_0333_));
 sg13g2_nand2_1 _1088_ (.Y(_0356_),
    .A(net180),
    .B(net160));
 sg13g2_nand2_1 _1089_ (.Y(_0357_),
    .A(net178),
    .B(net161));
 sg13g2_nand2_1 _1090_ (.Y(_0358_),
    .A(net163),
    .B(net178));
 sg13g2_xor2_1 _1091_ (.B(_0358_),
    .A(_0320_),
    .X(_0359_));
 sg13g2_nand2b_1 _1092_ (.Y(_0360_),
    .B(_0359_),
    .A_N(_0356_));
 sg13g2_xnor2_1 _1093_ (.Y(_0361_),
    .A(_0356_),
    .B(_0359_));
 sg13g2_inv_1 _1094_ (.Y(_0362_),
    .A(_0361_));
 sg13g2_o21ai_1 _1095_ (.B1(_0329_),
    .Y(_0363_),
    .A1(_0326_),
    .A2(_0330_));
 sg13g2_nor2b_1 _1096_ (.A(_0003_),
    .B_N(net165),
    .Y(_0364_));
 sg13g2_nor2b_1 _1097_ (.A(net175),
    .B_N(net167),
    .Y(_0365_));
 sg13g2_nor2b_1 _1098_ (.A(net175),
    .B_N(net171),
    .Y(_0366_));
 sg13g2_xnor2_1 _1099_ (.Y(_0367_),
    .A(_0327_),
    .B(_0366_));
 sg13g2_xor2_1 _1100_ (.B(_0367_),
    .A(_0364_),
    .X(_0368_));
 sg13g2_nand2_1 _1101_ (.Y(_0369_),
    .A(_0363_),
    .B(_0368_));
 sg13g2_xnor2_1 _1102_ (.Y(_0370_),
    .A(_0363_),
    .B(_0368_));
 sg13g2_xnor2_1 _1103_ (.Y(_0371_),
    .A(_0362_),
    .B(_0370_));
 sg13g2_nor2_1 _1104_ (.A(_0355_),
    .B(_0371_),
    .Y(_0372_));
 sg13g2_xor2_1 _1105_ (.B(_0371_),
    .A(_0355_),
    .X(_0373_));
 sg13g2_xnor2_1 _1106_ (.Y(_0374_),
    .A(_0354_),
    .B(_0373_));
 sg13g2_nor2_1 _1107_ (.A(_0348_),
    .B(_0374_),
    .Y(_0375_));
 sg13g2_or2_1 _1108_ (.X(_0376_),
    .B(_0374_),
    .A(_0348_));
 sg13g2_xor2_1 _1109_ (.B(_0374_),
    .A(_0348_),
    .X(_0377_));
 sg13g2_nand2_1 _1110_ (.Y(_0378_),
    .A(_0316_),
    .B(_0377_));
 sg13g2_xnor2_1 _1111_ (.Y(_0379_),
    .A(_0315_),
    .B(_0377_));
 sg13g2_nor2b_1 _1112_ (.A(_0339_),
    .B_N(_0379_),
    .Y(_0380_));
 sg13g2_xnor2_1 _1113_ (.Y(_0381_),
    .A(_0339_),
    .B(_0379_));
 sg13g2_o21ai_1 _1114_ (.B1(_0220_),
    .Y(_0382_),
    .A1(_0347_),
    .A2(_0381_));
 sg13g2_a21oi_1 _1115_ (.A1(_0347_),
    .A2(_0381_),
    .Y(_0383_),
    .B1(_0382_));
 sg13g2_o21ai_1 _1116_ (.B1(net77),
    .Y(_0384_),
    .A1(\controller_inst.pulse_counter[6] ),
    .A2(_0185_));
 sg13g2_a21oi_1 _1117_ (.A1(_0186_),
    .A2(_0384_),
    .Y(_0385_),
    .B1(_0225_));
 sg13g2_nand3_1 _1118_ (.B(_0218_),
    .C(_0223_),
    .A(_0196_),
    .Y(_0386_));
 sg13g2_nor3_1 _1119_ (.A(_0383_),
    .B(_0385_),
    .C(_0386_),
    .Y(_0387_));
 sg13g2_a21oi_1 _1120_ (.A1(_0108_),
    .A2(net144),
    .Y(_0048_),
    .B1(_0387_));
 sg13g2_a21oi_2 _1121_ (.B1(_0380_),
    .Y(_0388_),
    .A2(_0381_),
    .A1(_0347_));
 sg13g2_o21ai_1 _1122_ (.B1(_0352_),
    .Y(_0389_),
    .A1(_0349_),
    .A2(_0353_));
 sg13g2_a21oi_1 _1123_ (.A1(_0354_),
    .A2(_0373_),
    .Y(_0390_),
    .B1(_0372_));
 sg13g2_nand2_1 _1124_ (.Y(_0391_),
    .A(net181),
    .B(net157));
 sg13g2_o21ai_1 _1125_ (.B1(_0360_),
    .Y(_0392_),
    .A1(_0320_),
    .A2(_0358_));
 sg13g2_nand2_1 _1126_ (.Y(_0393_),
    .A(net180),
    .B(net158));
 sg13g2_nand2b_1 _1127_ (.Y(_0394_),
    .B(_0392_),
    .A_N(_0393_));
 sg13g2_xor2_1 _1128_ (.B(_0393_),
    .A(_0392_),
    .X(_0395_));
 sg13g2_xor2_1 _1129_ (.B(_0395_),
    .A(_0391_),
    .X(_0396_));
 sg13g2_o21ai_1 _1130_ (.B1(_0369_),
    .Y(_0397_),
    .A1(_0362_),
    .A2(_0370_));
 sg13g2_nor2b_1 _1131_ (.A(net179),
    .B_N(net160),
    .Y(_0398_));
 sg13g2_nand2b_1 _1132_ (.Y(_0399_),
    .B(net161),
    .A_N(net177));
 sg13g2_nand2b_1 _1133_ (.Y(_0400_),
    .B(net163),
    .A_N(net177));
 sg13g2_nor2_1 _1134_ (.A(_0358_),
    .B(_0399_),
    .Y(_0401_));
 sg13g2_xor2_1 _1135_ (.B(_0400_),
    .A(_0357_),
    .X(_0402_));
 sg13g2_xor2_1 _1136_ (.B(_0402_),
    .A(_0398_),
    .X(_0403_));
 sg13g2_a22oi_1 _1137_ (.Y(_0404_),
    .B1(_0367_),
    .B2(_0364_),
    .A2(_0365_),
    .A1(_0328_));
 sg13g2_nor2b_1 _1138_ (.A(net176),
    .B_N(net166),
    .Y(_0405_));
 sg13g2_nor2b_1 _1139_ (.A(net174),
    .B_N(net167),
    .Y(_0406_));
 sg13g2_nor2b_1 _1140_ (.A(net174),
    .B_N(net172),
    .Y(_0407_));
 sg13g2_xor2_1 _1141_ (.B(_0407_),
    .A(_0365_),
    .X(_0408_));
 sg13g2_xor2_1 _1142_ (.B(_0408_),
    .A(_0405_),
    .X(_0409_));
 sg13g2_nor2b_1 _1143_ (.A(_0404_),
    .B_N(_0409_),
    .Y(_0410_));
 sg13g2_xnor2_1 _1144_ (.Y(_0411_),
    .A(_0404_),
    .B(_0409_));
 sg13g2_xor2_1 _1145_ (.B(_0411_),
    .A(_0403_),
    .X(_0412_));
 sg13g2_and2_1 _1146_ (.A(_0397_),
    .B(_0412_),
    .X(_0413_));
 sg13g2_xor2_1 _1147_ (.B(_0412_),
    .A(_0397_),
    .X(_0414_));
 sg13g2_xnor2_1 _1148_ (.Y(_0415_),
    .A(_0396_),
    .B(_0414_));
 sg13g2_nor2_1 _1149_ (.A(_0390_),
    .B(_0415_),
    .Y(_0416_));
 sg13g2_xor2_1 _1150_ (.B(_0415_),
    .A(_0390_),
    .X(_0417_));
 sg13g2_xnor2_1 _1151_ (.Y(_0418_),
    .A(_0389_),
    .B(_0417_));
 sg13g2_a21oi_1 _1152_ (.A1(_0316_),
    .A2(_0377_),
    .Y(_0419_),
    .B1(_0375_));
 sg13g2_or2_1 _1153_ (.X(_0420_),
    .B(_0419_),
    .A(_0418_));
 sg13g2_xnor2_1 _1154_ (.Y(_0421_),
    .A(_0418_),
    .B(_0419_));
 sg13g2_or2_1 _1155_ (.X(_0422_),
    .B(_0421_),
    .A(_0388_));
 sg13g2_a21oi_1 _1156_ (.A1(_0388_),
    .A2(_0421_),
    .Y(_0423_),
    .B1(_0221_));
 sg13g2_xnor2_1 _1157_ (.Y(_0424_),
    .A(net118),
    .B(_0186_));
 sg13g2_a221oi_1 _1158_ (.B2(_0226_),
    .C1(_0386_),
    .B1(_0424_),
    .A1(_0422_),
    .Y(_0425_),
    .A2(_0423_));
 sg13g2_a21oi_1 _1159_ (.A1(_0111_),
    .A2(net142),
    .Y(_0049_),
    .B1(_0425_));
 sg13g2_a21oi_1 _1160_ (.A1(_0389_),
    .A2(_0417_),
    .Y(_0426_),
    .B1(_0416_));
 sg13g2_o21ai_1 _1161_ (.B1(_0394_),
    .Y(_0427_),
    .A1(_0391_),
    .A2(_0395_));
 sg13g2_a21oi_1 _1162_ (.A1(_0396_),
    .A2(_0414_),
    .Y(_0428_),
    .B1(_0413_));
 sg13g2_nand2_1 _1163_ (.Y(_0429_),
    .A(net180),
    .B(net157));
 sg13g2_a21oi_1 _1164_ (.A1(_0398_),
    .A2(_0402_),
    .Y(_0430_),
    .B1(_0401_));
 sg13g2_nand2b_1 _1165_ (.Y(_0431_),
    .B(\controller_inst.data_reg2[6] ),
    .A_N(net179));
 sg13g2_xor2_1 _1166_ (.B(_0431_),
    .A(_0430_),
    .X(_0432_));
 sg13g2_nand2b_1 _1167_ (.Y(_0433_),
    .B(_0432_),
    .A_N(_0429_));
 sg13g2_xnor2_1 _1168_ (.Y(_0434_),
    .A(_0429_),
    .B(_0432_));
 sg13g2_a21oi_1 _1169_ (.A1(_0403_),
    .A2(_0411_),
    .Y(_0435_),
    .B1(_0410_));
 sg13g2_nand2_1 _1170_ (.Y(_0436_),
    .A(net178),
    .B(net160));
 sg13g2_nand2b_2 _1171_ (.Y(_0437_),
    .B(net161),
    .A_N(net176));
 sg13g2_nor2b_1 _1172_ (.A(_0004_),
    .B_N(net163),
    .Y(_0438_));
 sg13g2_xnor2_1 _1173_ (.Y(_0439_),
    .A(_0399_),
    .B(_0438_));
 sg13g2_nand2b_1 _1174_ (.Y(_0440_),
    .B(_0439_),
    .A_N(_0436_));
 sg13g2_xnor2_1 _1175_ (.Y(_0441_),
    .A(_0436_),
    .B(_0439_));
 sg13g2_a22oi_1 _1176_ (.Y(_0442_),
    .B1(_0408_),
    .B2(_0405_),
    .A2(_0406_),
    .A1(_0366_));
 sg13g2_nor2b_1 _1177_ (.A(net175),
    .B_N(net166),
    .Y(_0443_));
 sg13g2_nor2b_1 _1178_ (.A(_0007_),
    .B_N(net170),
    .Y(_0444_));
 sg13g2_nor2b_1 _1179_ (.A(_0007_),
    .B_N(net172),
    .Y(_0445_));
 sg13g2_xor2_1 _1180_ (.B(_0445_),
    .A(_0406_),
    .X(_0446_));
 sg13g2_xor2_1 _1181_ (.B(_0446_),
    .A(_0443_),
    .X(_0447_));
 sg13g2_nor2b_1 _1182_ (.A(_0442_),
    .B_N(_0447_),
    .Y(_0448_));
 sg13g2_xnor2_1 _1183_ (.Y(_0449_),
    .A(_0442_),
    .B(_0447_));
 sg13g2_xnor2_1 _1184_ (.Y(_0450_),
    .A(_0441_),
    .B(_0449_));
 sg13g2_nor2_1 _1185_ (.A(_0435_),
    .B(_0450_),
    .Y(_0451_));
 sg13g2_xor2_1 _1186_ (.B(_0450_),
    .A(_0435_),
    .X(_0452_));
 sg13g2_xnor2_1 _1187_ (.Y(_0453_),
    .A(_0434_),
    .B(_0452_));
 sg13g2_or2_1 _1188_ (.X(_0454_),
    .B(_0453_),
    .A(_0428_));
 sg13g2_xor2_1 _1189_ (.B(_0453_),
    .A(_0428_),
    .X(_0455_));
 sg13g2_nand2_1 _1190_ (.Y(_0456_),
    .A(_0427_),
    .B(_0455_));
 sg13g2_xnor2_1 _1191_ (.Y(_0457_),
    .A(_0427_),
    .B(_0455_));
 sg13g2_nor2_1 _1192_ (.A(_0426_),
    .B(_0457_),
    .Y(_0458_));
 sg13g2_xnor2_1 _1193_ (.Y(_0459_),
    .A(_0426_),
    .B(_0457_));
 sg13g2_nand3_1 _1194_ (.B(_0422_),
    .C(_0459_),
    .A(_0420_),
    .Y(_0460_));
 sg13g2_a21o_1 _1195_ (.A2(_0422_),
    .A1(_0420_),
    .B1(_0459_),
    .X(_0461_));
 sg13g2_nand3_1 _1196_ (.B(_0460_),
    .C(_0461_),
    .A(net153),
    .Y(_0462_));
 sg13g2_o21ai_1 _1197_ (.B1(net102),
    .Y(_0463_),
    .A1(\controller_inst.pulse_counter[8] ),
    .A2(_0186_));
 sg13g2_a21oi_1 _1198_ (.A1(_0187_),
    .A2(_0463_),
    .Y(_0464_),
    .B1(_0225_));
 sg13g2_nor2_1 _1199_ (.A(_0386_),
    .B(_0464_),
    .Y(_0465_));
 sg13g2_a22oi_1 _1200_ (.Y(_0050_),
    .B1(_0462_),
    .B2(_0465_),
    .A2(net142),
    .A1(_0110_));
 sg13g2_o21ai_1 _1201_ (.B1(_0433_),
    .Y(_0466_),
    .A1(_0430_),
    .A2(_0431_));
 sg13g2_a21oi_1 _1202_ (.A1(_0434_),
    .A2(_0452_),
    .Y(_0467_),
    .B1(_0451_));
 sg13g2_nand2b_1 _1203_ (.Y(_0468_),
    .B(\controller_inst.data_reg2[7] ),
    .A_N(net179));
 sg13g2_o21ai_1 _1204_ (.B1(_0440_),
    .Y(_0469_),
    .A1(_0400_),
    .A2(_0437_));
 sg13g2_nand2_1 _1205_ (.Y(_0470_),
    .A(net178),
    .B(\controller_inst.data_reg2[6] ));
 sg13g2_nand2b_1 _1206_ (.Y(_0471_),
    .B(_0469_),
    .A_N(_0470_));
 sg13g2_xor2_1 _1207_ (.B(_0470_),
    .A(_0469_),
    .X(_0472_));
 sg13g2_xor2_1 _1208_ (.B(_0472_),
    .A(_0468_),
    .X(_0473_));
 sg13g2_a21oi_1 _1209_ (.A1(_0441_),
    .A2(_0449_),
    .Y(_0474_),
    .B1(_0448_));
 sg13g2_nand2b_1 _1210_ (.Y(_0475_),
    .B(net160),
    .A_N(net177));
 sg13g2_nand2b_1 _1211_ (.Y(_0476_),
    .B(net162),
    .A_N(net175));
 sg13g2_nand2b_2 _1212_ (.Y(_0477_),
    .B(net164),
    .A_N(_0005_));
 sg13g2_xor2_1 _1213_ (.B(_0477_),
    .A(_0437_),
    .X(_0478_));
 sg13g2_nand2b_1 _1214_ (.Y(_0479_),
    .B(_0478_),
    .A_N(_0475_));
 sg13g2_xnor2_1 _1215_ (.Y(_0480_),
    .A(_0475_),
    .B(_0478_));
 sg13g2_a22oi_1 _1216_ (.Y(_0481_),
    .B1(_0446_),
    .B2(_0443_),
    .A2(_0444_),
    .A1(_0407_));
 sg13g2_nor2b_1 _1217_ (.A(net174),
    .B_N(net165),
    .Y(_0482_));
 sg13g2_and2_1 _1218_ (.A(net170),
    .B(\controller_inst.pulse_width[10] ),
    .X(_0483_));
 sg13g2_nand2_1 _1219_ (.Y(_0484_),
    .A(net167),
    .B(\controller_inst.pulse_width[10] ));
 sg13g2_nand2_1 _1220_ (.Y(_0485_),
    .A(net172),
    .B(\controller_inst.pulse_width[10] ));
 sg13g2_xnor2_1 _1221_ (.Y(_0486_),
    .A(_0444_),
    .B(_0485_));
 sg13g2_xor2_1 _1222_ (.B(_0486_),
    .A(_0482_),
    .X(_0487_));
 sg13g2_nor2b_1 _1223_ (.A(_0481_),
    .B_N(_0487_),
    .Y(_0488_));
 sg13g2_xnor2_1 _1224_ (.Y(_0489_),
    .A(_0481_),
    .B(_0487_));
 sg13g2_xor2_1 _1225_ (.B(_0489_),
    .A(_0480_),
    .X(_0490_));
 sg13g2_nor2b_1 _1226_ (.A(_0474_),
    .B_N(_0490_),
    .Y(_0491_));
 sg13g2_xnor2_1 _1227_ (.Y(_0492_),
    .A(_0474_),
    .B(_0490_));
 sg13g2_xnor2_1 _1228_ (.Y(_0493_),
    .A(_0473_),
    .B(_0492_));
 sg13g2_nor2_1 _1229_ (.A(_0467_),
    .B(_0493_),
    .Y(_0494_));
 sg13g2_xor2_1 _1230_ (.B(_0493_),
    .A(_0467_),
    .X(_0495_));
 sg13g2_xnor2_1 _1231_ (.Y(_0496_),
    .A(_0466_),
    .B(_0495_));
 sg13g2_a21oi_1 _1232_ (.A1(_0454_),
    .A2(_0456_),
    .Y(_0497_),
    .B1(_0496_));
 sg13g2_nand3_1 _1233_ (.B(_0456_),
    .C(_0496_),
    .A(_0454_),
    .Y(_0498_));
 sg13g2_nand2b_1 _1234_ (.Y(_0499_),
    .B(_0498_),
    .A_N(_0497_));
 sg13g2_or2_1 _1235_ (.X(_0500_),
    .B(_0459_),
    .A(_0421_));
 sg13g2_or2_1 _1236_ (.X(_0501_),
    .B(_0500_),
    .A(_0388_));
 sg13g2_a221oi_1 _1237_ (.B2(_0457_),
    .C1(_0418_),
    .B1(_0426_),
    .A1(_0376_),
    .Y(_0502_),
    .A2(_0378_));
 sg13g2_nor2_1 _1238_ (.A(_0458_),
    .B(_0502_),
    .Y(_0503_));
 sg13g2_a21oi_1 _1239_ (.A1(_0501_),
    .A2(_0503_),
    .Y(_0504_),
    .B1(_0499_));
 sg13g2_nand3_1 _1240_ (.B(_0501_),
    .C(_0503_),
    .A(_0499_),
    .Y(_0505_));
 sg13g2_nor2_1 _1241_ (.A(_0221_),
    .B(_0504_),
    .Y(_0506_));
 sg13g2_xnor2_1 _1242_ (.Y(_0507_),
    .A(net98),
    .B(_0187_));
 sg13g2_a221oi_1 _1243_ (.B2(_0226_),
    .C1(net142),
    .B1(_0507_),
    .A1(_0505_),
    .Y(_0508_),
    .A2(_0506_));
 sg13g2_a21oi_1 _1244_ (.A1(_0113_),
    .A2(net142),
    .Y(_0051_),
    .B1(_0508_));
 sg13g2_a21oi_1 _1245_ (.A1(_0466_),
    .A2(_0495_),
    .Y(_0509_),
    .B1(_0494_));
 sg13g2_o21ai_1 _1246_ (.B1(_0471_),
    .Y(_0510_),
    .A1(_0468_),
    .A2(_0472_));
 sg13g2_a21oi_1 _1247_ (.A1(_0473_),
    .A2(_0492_),
    .Y(_0511_),
    .B1(_0491_));
 sg13g2_nand2_1 _1248_ (.Y(_0512_),
    .A(net178),
    .B(\controller_inst.data_reg2[7] ));
 sg13g2_o21ai_1 _1249_ (.B1(_0479_),
    .Y(_0513_),
    .A1(_0437_),
    .A2(_0477_));
 sg13g2_nor2b_1 _1250_ (.A(net177),
    .B_N(\controller_inst.data_reg2[6] ),
    .Y(_0514_));
 sg13g2_nand2_1 _1251_ (.Y(_0515_),
    .A(_0513_),
    .B(_0514_));
 sg13g2_nor2_1 _1252_ (.A(_0513_),
    .B(_0514_),
    .Y(_0516_));
 sg13g2_xor2_1 _1253_ (.B(_0514_),
    .A(_0513_),
    .X(_0517_));
 sg13g2_xnor2_1 _1254_ (.Y(_0518_),
    .A(_0512_),
    .B(_0517_));
 sg13g2_a21oi_1 _1255_ (.A1(_0480_),
    .A2(_0489_),
    .Y(_0519_),
    .B1(_0488_));
 sg13g2_nand2b_1 _1256_ (.Y(_0520_),
    .B(net159),
    .A_N(net176));
 sg13g2_nand2b_2 _1257_ (.Y(_0521_),
    .B(net162),
    .A_N(net174));
 sg13g2_nor2b_1 _1258_ (.A(net174),
    .B_N(net164),
    .Y(_0522_));
 sg13g2_xnor2_1 _1259_ (.Y(_0523_),
    .A(_0476_),
    .B(_0522_));
 sg13g2_nand2b_1 _1260_ (.Y(_0524_),
    .B(_0523_),
    .A_N(_0520_));
 sg13g2_xnor2_1 _1261_ (.Y(_0525_),
    .A(_0520_),
    .B(_0523_));
 sg13g2_a22oi_1 _1262_ (.Y(_0526_),
    .B1(_0486_),
    .B2(_0482_),
    .A2(_0483_),
    .A1(_0445_));
 sg13g2_nand2b_1 _1263_ (.Y(_0527_),
    .B(net165),
    .A_N(_0007_));
 sg13g2_nand2_1 _1264_ (.Y(_0528_),
    .A(net171),
    .B(\controller_inst.pulse_width[11] ));
 sg13g2_or2_1 _1265_ (.X(_0529_),
    .B(_0528_),
    .A(_0484_));
 sg13g2_and2_1 _1266_ (.A(_0484_),
    .B(_0528_),
    .X(_0530_));
 sg13g2_xnor2_1 _1267_ (.Y(_0531_),
    .A(_0483_),
    .B(_0528_));
 sg13g2_xnor2_1 _1268_ (.Y(_0532_),
    .A(_0527_),
    .B(_0531_));
 sg13g2_nor2b_1 _1269_ (.A(_0526_),
    .B_N(_0532_),
    .Y(_0533_));
 sg13g2_xnor2_1 _1270_ (.Y(_0534_),
    .A(_0526_),
    .B(_0532_));
 sg13g2_xor2_1 _1271_ (.B(_0534_),
    .A(_0525_),
    .X(_0535_));
 sg13g2_nor2b_1 _1272_ (.A(_0519_),
    .B_N(_0535_),
    .Y(_0536_));
 sg13g2_xnor2_1 _1273_ (.Y(_0537_),
    .A(_0519_),
    .B(_0535_));
 sg13g2_xnor2_1 _1274_ (.Y(_0538_),
    .A(_0518_),
    .B(_0537_));
 sg13g2_nor2_1 _1275_ (.A(_0511_),
    .B(_0538_),
    .Y(_0539_));
 sg13g2_xor2_1 _1276_ (.B(_0538_),
    .A(_0511_),
    .X(_0540_));
 sg13g2_xnor2_1 _1277_ (.Y(_0541_),
    .A(_0510_),
    .B(_0540_));
 sg13g2_nor2_1 _1278_ (.A(_0509_),
    .B(_0541_),
    .Y(_0542_));
 sg13g2_nand2_1 _1279_ (.Y(_0543_),
    .A(_0509_),
    .B(_0541_));
 sg13g2_nor2b_1 _1280_ (.A(_0542_),
    .B_N(_0543_),
    .Y(_0544_));
 sg13g2_o21ai_1 _1281_ (.B1(_0544_),
    .Y(_0545_),
    .A1(_0497_),
    .A2(_0504_));
 sg13g2_nor3_1 _1282_ (.A(_0497_),
    .B(_0504_),
    .C(_0544_),
    .Y(_0546_));
 sg13g2_nand3b_1 _1283_ (.B(net153),
    .C(_0545_),
    .Y(_0547_),
    .A_N(_0546_));
 sg13g2_o21ai_1 _1284_ (.B1(net92),
    .Y(_0548_),
    .A1(\controller_inst.pulse_counter[10] ),
    .A2(_0187_));
 sg13g2_a21oi_1 _1285_ (.A1(_0189_),
    .A2(_0548_),
    .Y(_0549_),
    .B1(_0225_));
 sg13g2_nor2_1 _1286_ (.A(net142),
    .B(_0549_),
    .Y(_0550_));
 sg13g2_a22oi_1 _1287_ (.Y(_0052_),
    .B1(_0547_),
    .B2(_0550_),
    .A2(net141),
    .A1(_0112_));
 sg13g2_a221oi_1 _1288_ (.B2(_0541_),
    .C1(_0496_),
    .B1(_0509_),
    .A1(_0454_),
    .Y(_0551_),
    .A2(_0456_));
 sg13g2_nor4_1 _1289_ (.A(_0458_),
    .B(_0502_),
    .C(_0542_),
    .D(_0551_),
    .Y(_0552_));
 sg13g2_o21ai_1 _1290_ (.B1(_0552_),
    .Y(_0553_),
    .A1(_0388_),
    .A2(_0500_));
 sg13g2_a21o_1 _1291_ (.A2(_0543_),
    .A1(_0498_),
    .B1(_0542_),
    .X(_0554_));
 sg13g2_o21ai_1 _1292_ (.B1(_0515_),
    .Y(_0555_),
    .A1(_0512_),
    .A2(_0516_));
 sg13g2_a21oi_1 _1293_ (.A1(_0518_),
    .A2(_0537_),
    .Y(_0556_),
    .B1(_0536_));
 sg13g2_a21oi_1 _1294_ (.A1(_0525_),
    .A2(_0534_),
    .Y(_0557_),
    .B1(_0533_));
 sg13g2_o21ai_1 _1295_ (.B1(_0529_),
    .Y(_0558_),
    .A1(_0527_),
    .A2(_0530_));
 sg13g2_nand2_1 _1296_ (.Y(_0559_),
    .A(net165),
    .B(\controller_inst.pulse_width[10] ));
 sg13g2_nand2_1 _1297_ (.Y(_0560_),
    .A(net167),
    .B(\controller_inst.pulse_width[12] ));
 sg13g2_and4_1 _1298_ (.A(net171),
    .B(net167),
    .C(\controller_inst.pulse_width[11] ),
    .D(\controller_inst.pulse_width[12] ),
    .X(_0561_));
 sg13g2_a22oi_1 _1299_ (.Y(_0562_),
    .B1(\controller_inst.pulse_width[12] ),
    .B2(net171),
    .A2(\controller_inst.pulse_width[11] ),
    .A1(net167));
 sg13g2_nor3_1 _1300_ (.A(_0559_),
    .B(_0561_),
    .C(_0562_),
    .Y(_0563_));
 sg13g2_o21ai_1 _1301_ (.B1(_0559_),
    .Y(_0564_),
    .A1(_0561_),
    .A2(_0562_));
 sg13g2_nor2b_1 _1302_ (.A(_0563_),
    .B_N(_0564_),
    .Y(_0565_));
 sg13g2_nand2_1 _1303_ (.Y(_0566_),
    .A(_0558_),
    .B(_0565_));
 sg13g2_xnor2_1 _1304_ (.Y(_0567_),
    .A(_0558_),
    .B(_0565_));
 sg13g2_nor2b_1 _1305_ (.A(net175),
    .B_N(net159),
    .Y(_0568_));
 sg13g2_nor2b_1 _1306_ (.A(_0007_),
    .B_N(net162),
    .Y(_0569_));
 sg13g2_nand2b_2 _1307_ (.Y(_0570_),
    .B(net164),
    .A_N(_0007_));
 sg13g2_xor2_1 _1308_ (.B(_0570_),
    .A(_0521_),
    .X(_0571_));
 sg13g2_nand2_1 _1309_ (.Y(_0572_),
    .A(_0568_),
    .B(_0571_));
 sg13g2_xnor2_1 _1310_ (.Y(_0573_),
    .A(_0568_),
    .B(_0571_));
 sg13g2_xor2_1 _1311_ (.B(_0573_),
    .A(_0567_),
    .X(_0574_));
 sg13g2_nor2b_1 _1312_ (.A(_0557_),
    .B_N(_0574_),
    .Y(_0575_));
 sg13g2_xnor2_1 _1313_ (.Y(_0576_),
    .A(_0557_),
    .B(_0574_));
 sg13g2_nand2b_1 _1314_ (.Y(_0577_),
    .B(net157),
    .A_N(net177));
 sg13g2_o21ai_1 _1315_ (.B1(_0524_),
    .Y(_0578_),
    .A1(_0477_),
    .A2(_0521_));
 sg13g2_nor2b_1 _1316_ (.A(net176),
    .B_N(net158),
    .Y(_0579_));
 sg13g2_nand2_1 _1317_ (.Y(_0580_),
    .A(_0578_),
    .B(_0579_));
 sg13g2_nor2_1 _1318_ (.A(_0578_),
    .B(_0579_),
    .Y(_0581_));
 sg13g2_xor2_1 _1319_ (.B(_0579_),
    .A(_0578_),
    .X(_0582_));
 sg13g2_xnor2_1 _1320_ (.Y(_0583_),
    .A(_0577_),
    .B(_0582_));
 sg13g2_xnor2_1 _1321_ (.Y(_0584_),
    .A(_0576_),
    .B(_0583_));
 sg13g2_or2_1 _1322_ (.X(_0585_),
    .B(_0584_),
    .A(_0556_));
 sg13g2_xor2_1 _1323_ (.B(_0584_),
    .A(_0556_),
    .X(_0586_));
 sg13g2_nand2_1 _1324_ (.Y(_0587_),
    .A(_0555_),
    .B(_0586_));
 sg13g2_xnor2_1 _1325_ (.Y(_0588_),
    .A(_0555_),
    .B(_0586_));
 sg13g2_a21oi_1 _1326_ (.A1(_0510_),
    .A2(_0540_),
    .Y(_0589_),
    .B1(_0539_));
 sg13g2_nor2_1 _1327_ (.A(_0588_),
    .B(_0589_),
    .Y(_0590_));
 sg13g2_xnor2_1 _1328_ (.Y(_0591_),
    .A(_0588_),
    .B(_0589_));
 sg13g2_inv_1 _1329_ (.Y(_0592_),
    .A(_0591_));
 sg13g2_nand3_1 _1330_ (.B(_0554_),
    .C(_0592_),
    .A(_0553_),
    .Y(_0593_));
 sg13g2_a21oi_1 _1331_ (.A1(_0553_),
    .A2(_0554_),
    .Y(_0594_),
    .B1(_0592_));
 sg13g2_nor2_1 _1332_ (.A(_0221_),
    .B(_0594_),
    .Y(_0595_));
 sg13g2_nand2_1 _1333_ (.Y(_0596_),
    .A(net124),
    .B(_0189_));
 sg13g2_a21o_1 _1334_ (.A2(_0596_),
    .A1(_0190_),
    .B1(_0225_),
    .X(_0597_));
 sg13g2_a21oi_1 _1335_ (.A1(_0593_),
    .A2(_0595_),
    .Y(_0598_),
    .B1(_0386_));
 sg13g2_a22oi_1 _1336_ (.Y(_0053_),
    .B1(_0597_),
    .B2(_0598_),
    .A2(net141),
    .A1(_0115_));
 sg13g2_o21ai_1 _1337_ (.B1(_0580_),
    .Y(_0599_),
    .A1(_0577_),
    .A2(_0581_));
 sg13g2_a21oi_1 _1338_ (.A1(_0576_),
    .A2(_0583_),
    .Y(_0600_),
    .B1(_0575_));
 sg13g2_o21ai_1 _1339_ (.B1(_0566_),
    .Y(_0601_),
    .A1(_0567_),
    .A2(_0573_));
 sg13g2_or2_1 _1340_ (.X(_0602_),
    .B(_0563_),
    .A(_0561_));
 sg13g2_nand2_1 _1341_ (.Y(_0603_),
    .A(net165),
    .B(\controller_inst.pulse_width[11] ));
 sg13g2_nand2_1 _1342_ (.Y(_0604_),
    .A(net167),
    .B(\controller_inst.pulse_width[13] ));
 sg13g2_nand2_1 _1343_ (.Y(_0605_),
    .A(net171),
    .B(\controller_inst.pulse_width[13] ));
 sg13g2_xor2_1 _1344_ (.B(_0605_),
    .A(_0560_),
    .X(_0606_));
 sg13g2_nand2b_1 _1345_ (.Y(_0607_),
    .B(_0606_),
    .A_N(_0603_));
 sg13g2_xnor2_1 _1346_ (.Y(_0608_),
    .A(_0603_),
    .B(_0606_));
 sg13g2_xnor2_1 _1347_ (.Y(_0609_),
    .A(_0602_),
    .B(_0608_));
 sg13g2_nor2b_1 _1348_ (.A(net174),
    .B_N(net159),
    .Y(_0610_));
 sg13g2_nand2_1 _1349_ (.Y(_0611_),
    .A(net162),
    .B(\controller_inst.pulse_width[10] ));
 sg13g2_nand2_1 _1350_ (.Y(_0612_),
    .A(net164),
    .B(\controller_inst.pulse_width[10] ));
 sg13g2_nor2_1 _1351_ (.A(_0570_),
    .B(_0611_),
    .Y(_0613_));
 sg13g2_xnor2_1 _1352_ (.Y(_0614_),
    .A(_0569_),
    .B(_0612_));
 sg13g2_xor2_1 _1353_ (.B(_0614_),
    .A(_0610_),
    .X(_0615_));
 sg13g2_nor2b_1 _1354_ (.A(_0609_),
    .B_N(_0615_),
    .Y(_0616_));
 sg13g2_xnor2_1 _1355_ (.Y(_0617_),
    .A(_0609_),
    .B(_0615_));
 sg13g2_nand2_1 _1356_ (.Y(_0618_),
    .A(_0601_),
    .B(_0617_));
 sg13g2_xnor2_1 _1357_ (.Y(_0619_),
    .A(_0601_),
    .B(_0617_));
 sg13g2_nor2b_1 _1358_ (.A(net176),
    .B_N(net157),
    .Y(_0620_));
 sg13g2_o21ai_1 _1359_ (.B1(_0572_),
    .Y(_0621_),
    .A1(_0521_),
    .A2(_0570_));
 sg13g2_nor2b_1 _1360_ (.A(net175),
    .B_N(net158),
    .Y(_0622_));
 sg13g2_and2_1 _1361_ (.A(_0621_),
    .B(_0622_),
    .X(_0623_));
 sg13g2_xor2_1 _1362_ (.B(_0622_),
    .A(_0621_),
    .X(_0624_));
 sg13g2_xnor2_1 _1363_ (.Y(_0625_),
    .A(_0620_),
    .B(_0624_));
 sg13g2_xor2_1 _1364_ (.B(_0625_),
    .A(_0619_),
    .X(_0626_));
 sg13g2_nor2b_1 _1365_ (.A(_0600_),
    .B_N(_0626_),
    .Y(_0627_));
 sg13g2_xnor2_1 _1366_ (.Y(_0628_),
    .A(_0600_),
    .B(_0626_));
 sg13g2_xnor2_1 _1367_ (.Y(_0629_),
    .A(_0599_),
    .B(_0628_));
 sg13g2_a21oi_1 _1368_ (.A1(_0585_),
    .A2(_0587_),
    .Y(_0630_),
    .B1(_0629_));
 sg13g2_nand3_1 _1369_ (.B(_0587_),
    .C(_0629_),
    .A(_0585_),
    .Y(_0631_));
 sg13g2_nand2b_1 _1370_ (.Y(_0632_),
    .B(_0631_),
    .A_N(_0630_));
 sg13g2_nor2b_1 _1371_ (.A(_0590_),
    .B_N(_0593_),
    .Y(_0633_));
 sg13g2_o21ai_1 _1372_ (.B1(net153),
    .Y(_0634_),
    .A1(_0632_),
    .A2(_0633_));
 sg13g2_a21o_1 _1373_ (.A2(_0633_),
    .A1(_0632_),
    .B1(_0634_),
    .X(_0635_));
 sg13g2_xnor2_1 _1374_ (.Y(_0636_),
    .A(net100),
    .B(_0190_));
 sg13g2_a21oi_1 _1375_ (.A1(_0226_),
    .A2(_0636_),
    .Y(_0637_),
    .B1(net141));
 sg13g2_a22oi_1 _1376_ (.Y(_0054_),
    .B1(_0635_),
    .B2(_0637_),
    .A2(net141),
    .A1(_0114_));
 sg13g2_nor2_1 _1377_ (.A(_0591_),
    .B(_0632_),
    .Y(_0638_));
 sg13g2_nand3_1 _1378_ (.B(_0554_),
    .C(_0638_),
    .A(_0553_),
    .Y(_0639_));
 sg13g2_a21oi_1 _1379_ (.A1(_0590_),
    .A2(_0631_),
    .Y(_0640_),
    .B1(_0630_));
 sg13g2_a21oi_1 _1380_ (.A1(_0620_),
    .A2(_0624_),
    .Y(_0641_),
    .B1(_0623_));
 sg13g2_o21ai_1 _1381_ (.B1(_0618_),
    .Y(_0642_),
    .A1(_0619_),
    .A2(_0625_));
 sg13g2_a21o_1 _1382_ (.A2(_0608_),
    .A1(_0602_),
    .B1(_0616_),
    .X(_0643_));
 sg13g2_o21ai_1 _1383_ (.B1(_0607_),
    .Y(_0644_),
    .A1(_0560_),
    .A2(_0605_));
 sg13g2_nand2_1 _1384_ (.Y(_0645_),
    .A(net165),
    .B(\controller_inst.pulse_width[12] ));
 sg13g2_nand2_1 _1385_ (.Y(_0646_),
    .A(net167),
    .B(\controller_inst.pulse_width[14] ));
 sg13g2_nand2_1 _1386_ (.Y(_0647_),
    .A(net171),
    .B(\controller_inst.pulse_width[14] ));
 sg13g2_xor2_1 _1387_ (.B(_0647_),
    .A(_0604_),
    .X(_0648_));
 sg13g2_nand2b_1 _1388_ (.Y(_0649_),
    .B(_0648_),
    .A_N(_0645_));
 sg13g2_xnor2_1 _1389_ (.Y(_0650_),
    .A(_0645_),
    .B(_0648_));
 sg13g2_xnor2_1 _1390_ (.Y(_0651_),
    .A(_0644_),
    .B(_0650_));
 sg13g2_nand2b_1 _1391_ (.Y(_0652_),
    .B(net159),
    .A_N(_0007_));
 sg13g2_nand2_1 _1392_ (.Y(_0653_),
    .A(net162),
    .B(\controller_inst.pulse_width[11] ));
 sg13g2_nand2_1 _1393_ (.Y(_0654_),
    .A(net164),
    .B(\controller_inst.pulse_width[11] ));
 sg13g2_xor2_1 _1394_ (.B(_0654_),
    .A(_0611_),
    .X(_0655_));
 sg13g2_nand2b_1 _1395_ (.Y(_0656_),
    .B(_0655_),
    .A_N(_0652_));
 sg13g2_xnor2_1 _1396_ (.Y(_0657_),
    .A(_0652_),
    .B(_0655_));
 sg13g2_nor2b_1 _1397_ (.A(_0651_),
    .B_N(_0657_),
    .Y(_0658_));
 sg13g2_xnor2_1 _1398_ (.Y(_0659_),
    .A(_0651_),
    .B(_0657_));
 sg13g2_xnor2_1 _1399_ (.Y(_0660_),
    .A(_0643_),
    .B(_0659_));
 sg13g2_nand2b_1 _1400_ (.Y(_0661_),
    .B(net157),
    .A_N(net175));
 sg13g2_a21oi_1 _1401_ (.A1(_0610_),
    .A2(_0614_),
    .Y(_0662_),
    .B1(_0613_));
 sg13g2_nand2b_1 _1402_ (.Y(_0663_),
    .B(net158),
    .A_N(net174));
 sg13g2_xor2_1 _1403_ (.B(_0663_),
    .A(_0662_),
    .X(_0664_));
 sg13g2_nand2b_1 _1404_ (.Y(_0665_),
    .B(_0664_),
    .A_N(_0661_));
 sg13g2_xnor2_1 _1405_ (.Y(_0666_),
    .A(_0661_),
    .B(_0664_));
 sg13g2_nor2b_1 _1406_ (.A(_0660_),
    .B_N(_0666_),
    .Y(_0667_));
 sg13g2_xnor2_1 _1407_ (.Y(_0668_),
    .A(_0660_),
    .B(_0666_));
 sg13g2_nand2_1 _1408_ (.Y(_0669_),
    .A(_0642_),
    .B(_0668_));
 sg13g2_xnor2_1 _1409_ (.Y(_0670_),
    .A(_0642_),
    .B(_0668_));
 sg13g2_xnor2_1 _1410_ (.Y(_0671_),
    .A(_0641_),
    .B(_0670_));
 sg13g2_a21o_2 _1411_ (.A2(_0628_),
    .A1(_0599_),
    .B1(_0627_),
    .X(_0672_));
 sg13g2_nor2b_1 _1412_ (.A(_0671_),
    .B_N(_0672_),
    .Y(_0673_));
 sg13g2_xor2_1 _1413_ (.B(_0672_),
    .A(_0671_),
    .X(_0674_));
 sg13g2_a21oi_1 _1414_ (.A1(_0639_),
    .A2(_0640_),
    .Y(_0675_),
    .B1(_0674_));
 sg13g2_nand3_1 _1415_ (.B(_0640_),
    .C(_0674_),
    .A(_0639_),
    .Y(_0676_));
 sg13g2_nand3b_1 _1416_ (.B(_0676_),
    .C(net153),
    .Y(_0677_),
    .A_N(_0675_));
 sg13g2_o21ai_1 _1417_ (.B1(net79),
    .Y(_0678_),
    .A1(\controller_inst.pulse_counter[13] ),
    .A2(_0190_));
 sg13g2_nand2b_1 _1418_ (.Y(_0679_),
    .B(_0678_),
    .A_N(_0191_));
 sg13g2_a21oi_1 _1419_ (.A1(_0226_),
    .A2(_0679_),
    .Y(_0680_),
    .B1(net141));
 sg13g2_a22oi_1 _1420_ (.Y(_0055_),
    .B1(_0677_),
    .B2(_0680_),
    .A2(net141),
    .A1(_0117_));
 sg13g2_o21ai_1 _1421_ (.B1(_0669_),
    .Y(_0681_),
    .A1(_0641_),
    .A2(_0670_));
 sg13g2_o21ai_1 _1422_ (.B1(_0665_),
    .Y(_0682_),
    .A1(_0662_),
    .A2(_0663_));
 sg13g2_a21oi_1 _1423_ (.A1(_0643_),
    .A2(_0659_),
    .Y(_0683_),
    .B1(_0667_));
 sg13g2_nand2_1 _1424_ (.Y(_0684_),
    .A(net159),
    .B(\controller_inst.pulse_width[10] ));
 sg13g2_o21ai_1 _1425_ (.B1(_0649_),
    .Y(_0685_),
    .A1(_0604_),
    .A2(_0647_));
 sg13g2_xnor2_1 _1426_ (.Y(_0686_),
    .A(_0684_),
    .B(_0685_));
 sg13g2_o21ai_1 _1427_ (.B1(_0656_),
    .Y(_0687_),
    .A1(_0612_),
    .A2(_0653_));
 sg13g2_nor2b_1 _1428_ (.A(_0007_),
    .B_N(net158),
    .Y(_0688_));
 sg13g2_xnor2_1 _1429_ (.Y(_0689_),
    .A(_0687_),
    .B(_0688_));
 sg13g2_nand2_1 _1430_ (.Y(_0690_),
    .A(net165),
    .B(\controller_inst.pulse_width[13] ));
 sg13g2_nand2_1 _1431_ (.Y(_0691_),
    .A(net171),
    .B(\controller_inst.pulse_width[15] ));
 sg13g2_xor2_1 _1432_ (.B(_0691_),
    .A(_0646_),
    .X(_0692_));
 sg13g2_nand2_1 _1433_ (.Y(_0693_),
    .A(net164),
    .B(\controller_inst.pulse_width[12] ));
 sg13g2_xor2_1 _1434_ (.B(_0693_),
    .A(_0653_),
    .X(_0694_));
 sg13g2_xnor2_1 _1435_ (.Y(_0695_),
    .A(_0692_),
    .B(_0694_));
 sg13g2_xnor2_1 _1436_ (.Y(_0696_),
    .A(_0690_),
    .B(_0695_));
 sg13g2_xnor2_1 _1437_ (.Y(_0697_),
    .A(_0689_),
    .B(_0696_));
 sg13g2_xnor2_1 _1438_ (.Y(_0698_),
    .A(_0686_),
    .B(_0697_));
 sg13g2_a21oi_1 _1439_ (.A1(_0644_),
    .A2(_0650_),
    .Y(_0699_),
    .B1(_0658_));
 sg13g2_nand2b_1 _1440_ (.Y(_0700_),
    .B(net157),
    .A_N(net174));
 sg13g2_xnor2_1 _1441_ (.Y(_0701_),
    .A(_0699_),
    .B(_0700_));
 sg13g2_xnor2_1 _1442_ (.Y(_0702_),
    .A(_0698_),
    .B(_0701_));
 sg13g2_xnor2_1 _1443_ (.Y(_0703_),
    .A(_0683_),
    .B(_0702_));
 sg13g2_xnor2_1 _1444_ (.Y(_0704_),
    .A(_0682_),
    .B(_0703_));
 sg13g2_xnor2_1 _1445_ (.Y(_0705_),
    .A(_0681_),
    .B(_0704_));
 sg13g2_o21ai_1 _1446_ (.B1(_0705_),
    .Y(_0706_),
    .A1(_0673_),
    .A2(_0675_));
 sg13g2_or3_1 _1447_ (.A(_0673_),
    .B(_0675_),
    .C(_0705_),
    .X(_0707_));
 sg13g2_nand3_1 _1448_ (.B(_0706_),
    .C(_0707_),
    .A(net153),
    .Y(_0708_));
 sg13g2_xnor2_1 _1449_ (.Y(_0709_),
    .A(_0116_),
    .B(_0191_));
 sg13g2_a21oi_1 _1450_ (.A1(_0226_),
    .A2(_0709_),
    .Y(_0710_),
    .B1(net141));
 sg13g2_a22oi_1 _1451_ (.Y(_0056_),
    .B1(_0708_),
    .B2(_0710_),
    .A2(net141),
    .A1(_0116_));
 sg13g2_nand2_2 _1452_ (.Y(_0711_),
    .A(net120),
    .B(_0208_));
 sg13g2_nor2_1 _1453_ (.A(_0169_),
    .B(net150),
    .Y(_0712_));
 sg13g2_mux2_1 _1454_ (.A0(net183),
    .A1(net108),
    .S(net148),
    .X(_0057_));
 sg13g2_mux2_1 _1455_ (.A0(net182),
    .A1(net131),
    .S(net148),
    .X(_0058_));
 sg13g2_mux2_1 _1456_ (.A0(net180),
    .A1(net121),
    .S(net149),
    .X(_0059_));
 sg13g2_nor2_1 _1457_ (.A(net179),
    .B(net149),
    .Y(_0713_));
 sg13g2_a21oi_1 _1458_ (.A1(net37),
    .A2(net148),
    .Y(_0060_),
    .B1(_0713_));
 sg13g2_mux2_1 _1459_ (.A0(net178),
    .A1(net205),
    .S(net147),
    .X(_0061_));
 sg13g2_nor2_1 _1460_ (.A(net177),
    .B(net148),
    .Y(_0714_));
 sg13g2_a21oi_1 _1461_ (.A1(net39),
    .A2(net147),
    .Y(_0062_),
    .B1(_0714_));
 sg13g2_nor2_1 _1462_ (.A(net176),
    .B(net147),
    .Y(_0715_));
 sg13g2_a21oi_1 _1463_ (.A1(net57),
    .A2(net147),
    .Y(_0063_),
    .B1(_0715_));
 sg13g2_nor2_1 _1464_ (.A(net175),
    .B(net146),
    .Y(_0716_));
 sg13g2_a21oi_1 _1465_ (.A1(net29),
    .A2(net146),
    .Y(_0064_),
    .B1(_0716_));
 sg13g2_nor2_1 _1466_ (.A(_0006_),
    .B(net148),
    .Y(_0717_));
 sg13g2_a21oi_1 _1467_ (.A1(net25),
    .A2(net148),
    .Y(_0065_),
    .B1(_0717_));
 sg13g2_nor2_1 _1468_ (.A(_0007_),
    .B(net148),
    .Y(_0718_));
 sg13g2_a21oi_1 _1469_ (.A1(net27),
    .A2(net148),
    .Y(_0066_),
    .B1(_0718_));
 sg13g2_mux2_1 _1470_ (.A0(\controller_inst.pulse_width[10] ),
    .A1(net116),
    .S(net147),
    .X(_0067_));
 sg13g2_mux2_1 _1471_ (.A0(\controller_inst.pulse_width[11] ),
    .A1(net112),
    .S(net146),
    .X(_0068_));
 sg13g2_mux2_1 _1472_ (.A0(net111),
    .A1(net109),
    .S(net146),
    .X(_0069_));
 sg13g2_mux2_1 _1473_ (.A0(net114),
    .A1(net185),
    .S(net146),
    .X(_0070_));
 sg13g2_mux2_1 _1474_ (.A0(net106),
    .A1(net184),
    .S(net146),
    .X(_0071_));
 sg13g2_nor2_1 _1475_ (.A(net35),
    .B(net146),
    .Y(_0719_));
 sg13g2_a21oi_1 _1476_ (.A1(_0119_),
    .A2(net146),
    .Y(_0072_),
    .B1(_0719_));
 sg13g2_mux2_1 _1477_ (.A0(net108),
    .A1(net173),
    .S(net150),
    .X(_0073_));
 sg13g2_mux2_1 _1478_ (.A0(net131),
    .A1(net168),
    .S(_0711_),
    .X(_0074_));
 sg13g2_mux2_1 _1479_ (.A0(net121),
    .A1(net165),
    .S(net150),
    .X(_0075_));
 sg13g2_mux2_1 _1480_ (.A0(net37),
    .A1(net164),
    .S(net150),
    .X(_0076_));
 sg13g2_mux2_1 _1481_ (.A0(net205),
    .A1(net162),
    .S(net150),
    .X(_0077_));
 sg13g2_mux2_1 _1482_ (.A0(net39),
    .A1(net159),
    .S(net150),
    .X(_0078_));
 sg13g2_mux2_1 _1483_ (.A0(net57),
    .A1(net158),
    .S(net150),
    .X(_0079_));
 sg13g2_mux2_1 _1484_ (.A0(net29),
    .A1(net157),
    .S(net150),
    .X(_0080_));
 sg13g2_nand2_1 _1485_ (.Y(_0720_),
    .A(\controller_inst.byte_ready ),
    .B(net155));
 sg13g2_nand4_1 _1486_ (.B(net155),
    .C(_0135_),
    .A(\controller_inst.byte_ready ),
    .Y(_0721_),
    .D(_0193_));
 sg13g2_mux2_1 _1487_ (.A0(net108),
    .A1(net129),
    .S(_0721_),
    .X(_0081_));
 sg13g2_mux2_1 _1488_ (.A0(\controller_inst.shift_reg_in[1] ),
    .A1(net126),
    .S(_0721_),
    .X(_0082_));
 sg13g2_mux2_1 _1489_ (.A0(net121),
    .A1(net137),
    .S(_0721_),
    .X(_0083_));
 sg13g2_mux2_1 _1490_ (.A0(net37),
    .A1(net128),
    .S(_0721_),
    .X(_0084_));
 sg13g2_mux2_1 _1491_ (.A0(\controller_inst.shift_reg_in[4] ),
    .A1(net70),
    .S(_0721_),
    .X(_0085_));
 sg13g2_mux2_1 _1492_ (.A0(net39),
    .A1(net52),
    .S(_0721_),
    .X(_0086_));
 sg13g2_mux2_1 _1493_ (.A0(net57),
    .A1(net59),
    .S(_0721_),
    .X(_0087_));
 sg13g2_mux2_1 _1494_ (.A0(net29),
    .A1(net60),
    .S(_0721_),
    .X(_0088_));
 sg13g2_nand2_1 _1495_ (.Y(_0722_),
    .A(net43),
    .B(_0125_));
 sg13g2_nor2b_1 _1496_ (.A(\controller_inst.bit_cnt[2] ),
    .B_N(\controller_inst.shift_reg_out[5] ),
    .Y(_0723_));
 sg13g2_a21oi_1 _1497_ (.A1(\controller_inst.bit_cnt[2] ),
    .A2(net34),
    .Y(_0724_),
    .B1(_0723_));
 sg13g2_a21oi_1 _1498_ (.A1(\controller_inst.bit_cnt[2] ),
    .A2(net31),
    .Y(_0725_),
    .B1(\controller_inst.bit_cnt[1] ));
 sg13g2_a21oi_1 _1499_ (.A1(_0120_),
    .A2(net43),
    .Y(_0726_),
    .B1(\controller_inst.bit_cnt[0] ));
 sg13g2_a22oi_1 _1500_ (.Y(_0727_),
    .B1(_0725_),
    .B2(_0726_),
    .A2(\controller_inst.bit_cnt[0] ),
    .A1(\controller_inst.bit_cnt[1] ));
 sg13g2_nor2b_1 _1501_ (.A(\controller_inst.bit_cnt[2] ),
    .B_N(\controller_inst.shift_reg_out[6] ),
    .Y(_0728_));
 sg13g2_a21oi_1 _1502_ (.A1(\controller_inst.bit_cnt[2] ),
    .A2(net32),
    .Y(_0729_),
    .B1(_0728_));
 sg13g2_a22oi_1 _1503_ (.Y(_0730_),
    .B1(_0729_),
    .B2(\controller_inst.bit_cnt[0] ),
    .A2(_0724_),
    .A1(\controller_inst.bit_cnt[1] ));
 sg13g2_nor2b_1 _1504_ (.A(net22),
    .B_N(\controller_inst.sck_d3 ),
    .Y(_0731_));
 sg13g2_o21ai_1 _1505_ (.B1(_0731_),
    .Y(_0732_),
    .A1(_0124_),
    .A2(_0127_));
 sg13g2_a21oi_1 _1506_ (.A1(_0727_),
    .A2(_0730_),
    .Y(_0733_),
    .B1(_0732_));
 sg13g2_o21ai_1 _1507_ (.B1(net155),
    .Y(_0734_),
    .A1(\controller_inst.spi_miso ),
    .A2(_0731_));
 sg13g2_o21ai_1 _1508_ (.B1(net44),
    .Y(_0089_),
    .A1(_0733_),
    .A2(_0734_));
 sg13g2_nand3b_1 _1509_ (.B(_0137_),
    .C(_0201_),
    .Y(_0735_),
    .A_N(\controller_inst.byte_ready ));
 sg13g2_nand3_1 _1510_ (.B(_0193_),
    .C(_0720_),
    .A(_0135_),
    .Y(_0736_));
 sg13g2_nand3_1 _1511_ (.B(_0735_),
    .C(_0736_),
    .A(_0153_),
    .Y(_0737_));
 sg13g2_nor2_2 _1512_ (.A(_0210_),
    .B(_0737_),
    .Y(_0738_));
 sg13g2_a21oi_1 _1513_ (.A1(_0169_),
    .A2(_0198_),
    .Y(_0739_),
    .B1(\controller_inst.byte_ready ));
 sg13g2_nor4_1 _1514_ (.A(_0102_),
    .B(_0167_),
    .C(_0200_),
    .D(_0739_),
    .Y(_0740_));
 sg13g2_o21ai_1 _1515_ (.B1(_0212_),
    .Y(_0741_),
    .A1(_0136_),
    .A2(_0740_));
 sg13g2_mux2_1 _1516_ (.A0(net156),
    .A1(_0741_),
    .S(_0738_),
    .X(_0090_));
 sg13g2_nor3_1 _1517_ (.A(net219),
    .B(net120),
    .C(_0167_),
    .Y(_0742_));
 sg13g2_nand2_1 _1518_ (.Y(_0743_),
    .A(_0137_),
    .B(_0199_));
 sg13g2_o21ai_1 _1519_ (.B1(_0219_),
    .Y(_0744_),
    .A1(_0742_),
    .A2(_0743_));
 sg13g2_mux2_1 _1520_ (.A0(net219),
    .A1(_0744_),
    .S(_0738_),
    .X(_0091_));
 sg13g2_nand2_1 _1521_ (.Y(_0745_),
    .A(_0212_),
    .B(_0219_));
 sg13g2_a21oi_1 _1522_ (.A1(_0137_),
    .A2(_0168_),
    .Y(_0746_),
    .B1(_0745_));
 sg13g2_nor2_1 _1523_ (.A(net87),
    .B(_0738_),
    .Y(_0747_));
 sg13g2_a21oi_1 _1524_ (.A1(_0738_),
    .A2(_0746_),
    .Y(_0092_),
    .B1(_0747_));
 sg13g2_a21oi_1 _1525_ (.A1(_0137_),
    .A2(_0200_),
    .Y(_0748_),
    .B1(_0147_));
 sg13g2_nand2b_1 _1526_ (.Y(_0749_),
    .B(_0738_),
    .A_N(_0748_));
 sg13g2_nand2_1 _1527_ (.Y(_0093_),
    .A(net203),
    .B(_0749_));
 sg13g2_nor2_1 _1528_ (.A(_0130_),
    .B(_0217_),
    .Y(_0750_));
 sg13g2_nor3_2 _1529_ (.A(_0206_),
    .B(_0211_),
    .C(_0750_),
    .Y(_0751_));
 sg13g2_nor3_1 _1530_ (.A(net51),
    .B(net184),
    .C(net185),
    .Y(_0752_));
 sg13g2_a21oi_1 _1531_ (.A1(\controller_inst.data_reg1[1] ),
    .A2(_0197_),
    .Y(_0753_),
    .B1(_0217_));
 sg13g2_nand2_2 _1532_ (.Y(_0754_),
    .A(_0153_),
    .B(_0753_));
 sg13g2_inv_1 _1533_ (.Y(_0755_),
    .A(_0754_));
 sg13g2_nand2b_2 _1534_ (.Y(_0756_),
    .B(_0197_),
    .A_N(\controller_inst.data_reg1[1] ));
 sg13g2_a22oi_1 _1535_ (.Y(_0757_),
    .B1(_0752_),
    .B2(_0754_),
    .A2(net152),
    .A1(net25));
 sg13g2_o21ai_1 _1536_ (.B1(_0757_),
    .Y(_0758_),
    .A1(_0752_),
    .A2(_0756_));
 sg13g2_mux2_1 _1537_ (.A0(net104),
    .A1(_0758_),
    .S(net140),
    .X(_0094_));
 sg13g2_nor2_1 _1538_ (.A(net72),
    .B(net140),
    .Y(_0759_));
 sg13g2_nor2b_1 _1539_ (.A(net184),
    .B_N(net185),
    .Y(_0760_));
 sg13g2_nand2_1 _1540_ (.Y(_0761_),
    .A(_0119_),
    .B(_0760_));
 sg13g2_or2_1 _1541_ (.X(_0762_),
    .B(_0761_),
    .A(_0754_));
 sg13g2_a21oi_1 _1542_ (.A1(_0756_),
    .A2(_0761_),
    .Y(_0763_),
    .B1(net152));
 sg13g2_a22oi_1 _1543_ (.Y(_0764_),
    .B1(_0762_),
    .B2(_0763_),
    .A2(net152),
    .A1(net27));
 sg13g2_a21oi_1 _1544_ (.A1(net140),
    .A2(_0764_),
    .Y(_0095_),
    .B1(_0759_));
 sg13g2_nor2_1 _1545_ (.A(net88),
    .B(net140),
    .Y(_0765_));
 sg13g2_nor2b_1 _1546_ (.A(net185),
    .B_N(net184),
    .Y(_0766_));
 sg13g2_nand2_1 _1547_ (.Y(_0767_),
    .A(_0119_),
    .B(_0766_));
 sg13g2_or2_1 _1548_ (.X(_0768_),
    .B(_0767_),
    .A(_0754_));
 sg13g2_a21oi_1 _1549_ (.A1(_0756_),
    .A2(_0767_),
    .Y(_0769_),
    .B1(net151));
 sg13g2_a22oi_1 _1550_ (.Y(_0770_),
    .B1(_0768_),
    .B2(_0769_),
    .A2(net151),
    .A1(\controller_inst.data_reg1[2] ));
 sg13g2_a21oi_1 _1551_ (.A1(net140),
    .A2(_0770_),
    .Y(_0096_),
    .B1(_0765_));
 sg13g2_nor2_1 _1552_ (.A(net85),
    .B(net140),
    .Y(_0771_));
 sg13g2_nand3_1 _1553_ (.B(net184),
    .C(net185),
    .A(_0119_),
    .Y(_0772_));
 sg13g2_or2_1 _1554_ (.X(_0773_),
    .B(_0772_),
    .A(_0754_));
 sg13g2_a21oi_1 _1555_ (.A1(_0756_),
    .A2(_0772_),
    .Y(_0774_),
    .B1(net151));
 sg13g2_a22oi_1 _1556_ (.Y(_0775_),
    .B1(_0773_),
    .B2(_0774_),
    .A2(net151),
    .A1(\controller_inst.data_reg1[3] ));
 sg13g2_a21oi_1 _1557_ (.A1(net139),
    .A2(_0775_),
    .Y(_0097_),
    .B1(_0771_));
 sg13g2_nor2_1 _1558_ (.A(net65),
    .B(net139),
    .Y(_0776_));
 sg13g2_nor3_1 _1559_ (.A(_0119_),
    .B(net184),
    .C(net185),
    .Y(_0777_));
 sg13g2_nand2_1 _1560_ (.Y(_0778_),
    .A(_0223_),
    .B(_0777_));
 sg13g2_a22oi_1 _1561_ (.Y(_0779_),
    .B1(_0778_),
    .B2(_0756_),
    .A2(_0777_),
    .A1(_0755_));
 sg13g2_a21oi_1 _1562_ (.A1(\controller_inst.data_reg1[4] ),
    .A2(net151),
    .Y(_0780_),
    .B1(_0779_));
 sg13g2_a21oi_1 _1563_ (.A1(net139),
    .A2(_0780_),
    .Y(_0098_),
    .B1(_0776_));
 sg13g2_nor2_1 _1564_ (.A(net75),
    .B(net140),
    .Y(_0781_));
 sg13g2_nand2_1 _1565_ (.Y(_0782_),
    .A(net51),
    .B(_0760_));
 sg13g2_or2_1 _1566_ (.X(_0783_),
    .B(_0782_),
    .A(_0754_));
 sg13g2_a21oi_1 _1567_ (.A1(_0756_),
    .A2(_0782_),
    .Y(_0784_),
    .B1(net151));
 sg13g2_a22oi_1 _1568_ (.Y(_0785_),
    .B1(_0783_),
    .B2(_0784_),
    .A2(net151),
    .A1(net185));
 sg13g2_a21oi_1 _1569_ (.A1(net139),
    .A2(_0785_),
    .Y(_0099_),
    .B1(_0781_));
 sg13g2_nor2_1 _1570_ (.A(net81),
    .B(net139),
    .Y(_0786_));
 sg13g2_and2_1 _1571_ (.A(net51),
    .B(_0766_),
    .X(_0787_));
 sg13g2_nor2_1 _1572_ (.A(_0756_),
    .B(_0787_),
    .Y(_0788_));
 sg13g2_a221oi_1 _1573_ (.B2(_0787_),
    .C1(_0788_),
    .B1(_0754_),
    .A1(net184),
    .Y(_0789_),
    .A2(net151));
 sg13g2_a21oi_1 _1574_ (.A1(net139),
    .A2(_0789_),
    .Y(_0100_),
    .B1(_0786_));
 sg13g2_and3_1 _1575_ (.X(_0790_),
    .A(net51),
    .B(\controller_inst.data_reg1[6] ),
    .C(\controller_inst.data_reg1[5] ));
 sg13g2_nand2_1 _1576_ (.Y(_0791_),
    .A(net51),
    .B(net152));
 sg13g2_o21ai_1 _1577_ (.B1(_0791_),
    .Y(_0792_),
    .A1(_0756_),
    .A2(_0790_));
 sg13g2_a21oi_1 _1578_ (.A1(_0754_),
    .A2(_0790_),
    .Y(_0793_),
    .B1(_0792_));
 sg13g2_nor2_1 _1579_ (.A(net83),
    .B(net139),
    .Y(_0794_));
 sg13g2_a21oi_1 _1580_ (.A1(net139),
    .A2(_0793_),
    .Y(_0101_),
    .B1(_0794_));
 sg13g2_buf_1 _1581_ (.A(net23),
    .X(_0011_));
 sg13g2_dfrbpq_1 _1582_ (.RESET_B(net198),
    .D(_0012_),
    .Q(\controller_inst.shift_reg_out[0] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_1 _1583_ (.RESET_B(net197),
    .D(_0013_),
    .Q(\controller_inst.shift_reg_out[1] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_1 _1584_ (.RESET_B(net197),
    .D(_0014_),
    .Q(\controller_inst.shift_reg_out[2] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_1 _1585_ (.RESET_B(net197),
    .D(_0015_),
    .Q(\controller_inst.shift_reg_out[3] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_1 _1586_ (.RESET_B(net197),
    .D(net42),
    .Q(\controller_inst.shift_reg_out[5] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_1 _1587_ (.RESET_B(net197),
    .D(net64),
    .Q(\controller_inst.shift_reg_out[6] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_1 _1588_ (.RESET_B(net196),
    .D(_0018_),
    .Q(\controller_inst.shift_reg_out[7] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_1 _1589_ (.RESET_B(net191),
    .D(_0019_),
    .Q(\controller_inst.data_reg1[0] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _1590_ (.RESET_B(net191),
    .D(_0020_),
    .Q(\controller_inst.data_reg1[1] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_1 _1591_ (.RESET_B(net190),
    .D(_0021_),
    .Q(\controller_inst.data_reg1[2] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_1 _1592_ (.RESET_B(net188),
    .D(_0022_),
    .Q(\controller_inst.data_reg1[3] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_2 _1593_ (.RESET_B(net188),
    .D(net110),
    .Q(\controller_inst.data_reg1[4] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_1 _1594_ (.RESET_B(net189),
    .D(_0024_),
    .Q(\controller_inst.data_reg1[5] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_1 _1595_ (.RESET_B(net189),
    .D(_0025_),
    .Q(\controller_inst.data_reg1[6] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_2 _1596_ (.RESET_B(net190),
    .D(_0026_),
    .Q(\controller_inst.data_reg1[7] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_2 _1597_ (.RESET_B(net199),
    .D(net54),
    .Q(\controller_inst.bit_cnt[0] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _1598_ (.RESET_B(net197),
    .D(net50),
    .Q(\controller_inst.bit_cnt[1] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _1599_ (.RESET_B(net198),
    .D(net69),
    .Q(\controller_inst.bit_cnt[2] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_1 _1600_ (.RESET_B(net196),
    .D(net74),
    .Q(\controller_inst.prog_done ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_2 _1601_ (.RESET_B(net199),
    .D(_0031_),
    .Q(\controller_inst.shift_reg_in[0] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _1602_ (.RESET_B(net191),
    .D(_0032_),
    .Q(\controller_inst.shift_reg_in[1] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _1603_ (.RESET_B(net191),
    .D(_0033_),
    .Q(\controller_inst.shift_reg_in[2] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _1604_ (.RESET_B(net191),
    .D(_0034_),
    .Q(\controller_inst.shift_reg_in[3] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_2 _1605_ (.RESET_B(net190),
    .D(_0035_),
    .Q(\controller_inst.shift_reg_in[4] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_2 _1606_ (.RESET_B(net188),
    .D(_0036_),
    .Q(\controller_inst.shift_reg_in[5] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_2 _1607_ (.RESET_B(net189),
    .D(_0037_),
    .Q(\controller_inst.shift_reg_in[6] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_2 _1608_ (.RESET_B(net188),
    .D(_0038_),
    .Q(\controller_inst.shift_reg_in[7] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _1609_ (.RESET_B(net196),
    .D(net24),
    .Q(\controller_inst.error ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_1 _1610_ (.RESET_B(net197),
    .D(net2),
    .Q(\controller_inst.sck_d1 ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_1 _1611_ (.RESET_B(net196),
    .D(net56),
    .Q(_0001_),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _1612_ (.RESET_B(net195),
    .D(net218),
    .Q(\controller_inst.pulse_counter[0] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _1613_ (.RESET_B(net199),
    .D(net91),
    .Q(\controller_inst.pulse_counter[1] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _1614_ (.RESET_B(net199),
    .D(net123),
    .Q(\controller_inst.pulse_counter[2] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _1615_ (.RESET_B(net199),
    .D(net97),
    .Q(\controller_inst.pulse_counter[3] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _1616_ (.RESET_B(net195),
    .D(net47),
    .Q(\controller_inst.pulse_counter[4] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_1 _1617_ (.RESET_B(net195),
    .D(net62),
    .Q(\controller_inst.pulse_counter[5] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _1618_ (.RESET_B(net195),
    .D(net135),
    .Q(\controller_inst.pulse_counter[6] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_1 _1619_ (.RESET_B(net195),
    .D(net78),
    .Q(\controller_inst.pulse_counter[7] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _1620_ (.RESET_B(net194),
    .D(net119),
    .Q(\controller_inst.pulse_counter[8] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_1 _1621_ (.RESET_B(net194),
    .D(net103),
    .Q(\controller_inst.pulse_counter[9] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_2 _1622_ (.RESET_B(net194),
    .D(net99),
    .Q(\controller_inst.pulse_counter[10] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_2 _1623_ (.RESET_B(net194),
    .D(net93),
    .Q(\controller_inst.pulse_counter[11] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _1624_ (.RESET_B(net194),
    .D(net125),
    .Q(\controller_inst.pulse_counter[12] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _1625_ (.RESET_B(net194),
    .D(net101),
    .Q(\controller_inst.pulse_counter[13] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _1626_ (.RESET_B(net194),
    .D(net80),
    .Q(\controller_inst.pulse_counter[14] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _1627_ (.RESET_B(net194),
    .D(net95),
    .Q(\controller_inst.pulse_counter[15] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _1628_ (.RESET_B(net197),
    .D(net21),
    .Q(\controller_inst.sck_d2 ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _1629_ (.RESET_B(net196),
    .D(_0057_),
    .Q(\controller_inst.pulse_width[0] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _1630_ (.RESET_B(net191),
    .D(_0058_),
    .Q(\controller_inst.pulse_width[1] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _1631_ (.RESET_B(net187),
    .D(_0059_),
    .Q(\controller_inst.pulse_width[2] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _1632_ (.RESET_B(net187),
    .D(net38),
    .Q(_0002_),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_2 _1633_ (.RESET_B(net187),
    .D(_0061_),
    .Q(\controller_inst.pulse_width[4] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _1634_ (.RESET_B(net187),
    .D(net40),
    .Q(_0003_),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_1 _1635_ (.RESET_B(net186),
    .D(net58),
    .Q(_0004_),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_1 _1636_ (.RESET_B(net186),
    .D(net30),
    .Q(_0005_),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _1637_ (.RESET_B(net191),
    .D(net26),
    .Q(_0006_),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_2 _1638_ (.RESET_B(net187),
    .D(net28),
    .Q(_0007_),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _1639_ (.RESET_B(net190),
    .D(net117),
    .Q(\controller_inst.pulse_width[10] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_2 _1640_ (.RESET_B(net188),
    .D(net113),
    .Q(\controller_inst.pulse_width[11] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_2 _1641_ (.RESET_B(net186),
    .D(_0069_),
    .Q(\controller_inst.pulse_width[12] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_2 _1642_ (.RESET_B(net186),
    .D(net115),
    .Q(\controller_inst.pulse_width[13] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _1643_ (.RESET_B(net188),
    .D(net107),
    .Q(\controller_inst.pulse_width[14] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _1644_ (.RESET_B(net188),
    .D(net36),
    .Q(\controller_inst.pulse_width[15] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _1645_ (.RESET_B(net196),
    .D(_0073_),
    .Q(\controller_inst.data_reg2[0] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _1646_ (.RESET_B(net193),
    .D(_0074_),
    .Q(\controller_inst.data_reg2[1] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _1647_ (.RESET_B(net187),
    .D(_0075_),
    .Q(\controller_inst.data_reg2[2] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _1648_ (.RESET_B(net186),
    .D(_0076_),
    .Q(\controller_inst.data_reg2[3] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _1649_ (.RESET_B(net186),
    .D(net206),
    .Q(\controller_inst.data_reg2[4] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _1650_ (.RESET_B(net187),
    .D(_0078_),
    .Q(\controller_inst.data_reg2[5] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_2 _1651_ (.RESET_B(net186),
    .D(_0079_),
    .Q(\controller_inst.data_reg2[6] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _1652_ (.RESET_B(net186),
    .D(_0080_),
    .Q(\controller_inst.data_reg2[7] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _1653_ (.RESET_B(net198),
    .D(net22),
    .Q(\controller_inst.sck_d3 ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _1654_ (.RESET_B(net192),
    .D(_0081_),
    .Q(\controller_inst.cmd_reg[0] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _1655_ (.RESET_B(net191),
    .D(net127),
    .Q(\controller_inst.cmd_reg[1] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _1656_ (.RESET_B(net192),
    .D(_0083_),
    .Q(\controller_inst.cmd_reg[2] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_2 _1657_ (.RESET_B(net192),
    .D(_0084_),
    .Q(\controller_inst.cmd_reg[3] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_1 _1658_ (.RESET_B(net188),
    .D(net71),
    .Q(\controller_inst.cmd_reg[4] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_1 _1659_ (.RESET_B(net189),
    .D(_0086_),
    .Q(\controller_inst.cmd_reg[5] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_1 _1660_ (.RESET_B(net189),
    .D(_0087_),
    .Q(\controller_inst.cmd_reg[6] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_1 _1661_ (.RESET_B(net189),
    .D(_0088_),
    .Q(\controller_inst.cmd_reg[7] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_1 _1662_ (.RESET_B(net200),
    .D(net45),
    .Q(\controller_inst.spi_miso ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_2 _1663_ (.RESET_B(net199),
    .D(_0090_),
    .Q(\controller_inst.state[0] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _1664_ (.RESET_B(net196),
    .D(_0091_),
    .Q(\controller_inst.state[1] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _1665_ (.RESET_B(net196),
    .D(_0092_),
    .Q(\controller_inst.state[2] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _1666_ (.RESET_B(net200),
    .D(_0093_),
    .Q(\controller_inst.state[3] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _1667_ (.RESET_B(net198),
    .D(_0010_),
    .Q(_0008_),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_1 _1668_ (.RESET_B(net192),
    .D(net105),
    .Q(uio_out[0]),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_1 _1669_ (.RESET_B(net193),
    .D(_0095_),
    .Q(uio_out[1]),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_1 _1670_ (.RESET_B(net192),
    .D(net89),
    .Q(uio_out[2]),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_1 _1671_ (.RESET_B(net192),
    .D(net86),
    .Q(uio_out[3]),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_1 _1672_ (.RESET_B(net192),
    .D(net66),
    .Q(uio_out[4]),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_1 _1673_ (.RESET_B(net192),
    .D(net76),
    .Q(uio_out[5]),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_1 _1674_ (.RESET_B(net189),
    .D(net82),
    .Q(uio_out[6]),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_1 _1675_ (.RESET_B(net189),
    .D(net84),
    .Q(uio_out[7]),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_2 _1676_ (.RESET_B(net199),
    .D(_0000_),
    .Q(\controller_inst.byte_ready ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _1677_ (.RESET_B(net198),
    .D(_0011_),
    .Q(_0009_),
    .CLK(clknet_4_14_0_clk));
 sg13g2_tiehi tt_um_sujanreddy_synapse_14 (.L_HI(net14));
 sg13g2_tiehi tt_um_sujanreddy_synapse_15 (.L_HI(net15));
 sg13g2_tiehi tt_um_sujanreddy_synapse_16 (.L_HI(net16));
 sg13g2_tiehi tt_um_sujanreddy_synapse_17 (.L_HI(net17));
 sg13g2_tiehi tt_um_sujanreddy_synapse_18 (.L_HI(net18));
 sg13g2_tiehi tt_um_sujanreddy_synapse_19 (.L_HI(net19));
 sg13g2_tiehi tt_um_sujanreddy_synapse_20 (.L_HI(net20));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_sujanreddy_synapse_10 (.L_LO(net10));
 sg13g2_tielo tt_um_sujanreddy_synapse_11 (.L_LO(net11));
 sg13g2_tielo tt_um_sujanreddy_synapse_12 (.L_LO(net12));
 sg13g2_tiehi tt_um_sujanreddy_synapse_13 (.L_HI(net13));
 sg13g2_buf_1 _1690_ (.A(\controller_inst.spi_miso ),
    .X(uo_out[0]));
 sg13g2_buf_1 _1691_ (.A(\controller_inst.ready ),
    .X(uo_out[1]));
 sg13g2_buf_1 _1692_ (.A(\controller_inst.error ),
    .X(uo_out[2]));
 sg13g2_buf_1 _1693_ (.A(\controller_inst.prog_done ),
    .X(uo_out[3]));
 sg13g2_buf_8 fanout138 (.A(_0154_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(net140),
    .X(net139));
 sg13g2_buf_8 fanout140 (.A(_0751_),
    .X(net140));
 sg13g2_buf_8 fanout141 (.A(_0224_),
    .X(net141));
 sg13g2_buf_1 fanout142 (.A(_0224_),
    .X(net142));
 sg13g2_buf_8 fanout143 (.A(net144),
    .X(net143));
 sg13g2_buf_8 fanout144 (.A(_0224_),
    .X(net144));
 sg13g2_buf_8 fanout145 (.A(_0174_),
    .X(net145));
 sg13g2_buf_8 fanout146 (.A(net149),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(net149),
    .X(net147));
 sg13g2_buf_8 fanout148 (.A(net149),
    .X(net148));
 sg13g2_buf_8 fanout149 (.A(_0712_),
    .X(net149));
 sg13g2_buf_8 fanout150 (.A(_0711_),
    .X(net150));
 sg13g2_buf_8 fanout151 (.A(net152),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_0222_),
    .X(net152));
 sg13g2_buf_8 fanout153 (.A(_0220_),
    .X(net153));
 sg13g2_buf_8 fanout154 (.A(_0129_),
    .X(net154));
 sg13g2_buf_8 fanout155 (.A(net67),
    .X(net155));
 sg13g2_buf_8 fanout156 (.A(net220),
    .X(net156));
 sg13g2_buf_8 fanout157 (.A(net133),
    .X(net157));
 sg13g2_buf_8 fanout158 (.A(net214),
    .X(net158));
 sg13g2_buf_8 fanout159 (.A(net210),
    .X(net159));
 sg13g2_buf_1 fanout160 (.A(\controller_inst.data_reg2[5] ),
    .X(net160));
 sg13g2_buf_8 fanout161 (.A(net162),
    .X(net161));
 sg13g2_buf_8 fanout162 (.A(\controller_inst.data_reg2[4] ),
    .X(net162));
 sg13g2_buf_8 fanout163 (.A(net164),
    .X(net163));
 sg13g2_buf_8 fanout164 (.A(net208),
    .X(net164));
 sg13g2_buf_8 fanout165 (.A(net212),
    .X(net165));
 sg13g2_buf_8 fanout166 (.A(\controller_inst.data_reg2[2] ),
    .X(net166));
 sg13g2_buf_8 fanout167 (.A(net170),
    .X(net167));
 sg13g2_buf_8 fanout168 (.A(net170),
    .X(net168));
 sg13g2_buf_1 fanout169 (.A(net170),
    .X(net169));
 sg13g2_buf_8 fanout170 (.A(net132),
    .X(net170));
 sg13g2_buf_8 fanout171 (.A(net172),
    .X(net171));
 sg13g2_buf_8 fanout172 (.A(net216),
    .X(net172));
 sg13g2_buf_1 fanout173 (.A(net216),
    .X(net173));
 sg13g2_buf_8 fanout174 (.A(_0006_),
    .X(net174));
 sg13g2_buf_8 fanout175 (.A(_0005_),
    .X(net175));
 sg13g2_buf_8 fanout176 (.A(_0004_),
    .X(net176));
 sg13g2_buf_8 fanout177 (.A(_0003_),
    .X(net177));
 sg13g2_buf_8 fanout178 (.A(net211),
    .X(net178));
 sg13g2_buf_8 fanout179 (.A(_0002_),
    .X(net179));
 sg13g2_buf_8 fanout180 (.A(net207),
    .X(net180));
 sg13g2_buf_8 fanout181 (.A(\controller_inst.pulse_width[1] ),
    .X(net181));
 sg13g2_buf_1 fanout182 (.A(net136),
    .X(net182));
 sg13g2_buf_8 fanout183 (.A(net215),
    .X(net183));
 sg13g2_buf_8 fanout184 (.A(net209),
    .X(net184));
 sg13g2_buf_8 fanout185 (.A(net204),
    .X(net185));
 sg13g2_buf_8 fanout186 (.A(net187),
    .X(net186));
 sg13g2_buf_8 fanout187 (.A(net201),
    .X(net187));
 sg13g2_buf_8 fanout188 (.A(net190),
    .X(net188));
 sg13g2_buf_8 fanout189 (.A(net190),
    .X(net189));
 sg13g2_buf_8 fanout190 (.A(net201),
    .X(net190));
 sg13g2_buf_8 fanout191 (.A(net193),
    .X(net191));
 sg13g2_buf_8 fanout192 (.A(net193),
    .X(net192));
 sg13g2_buf_8 fanout193 (.A(net201),
    .X(net193));
 sg13g2_buf_8 fanout194 (.A(net201),
    .X(net194));
 sg13g2_buf_8 fanout195 (.A(net201),
    .X(net195));
 sg13g2_buf_8 fanout196 (.A(net200),
    .X(net196));
 sg13g2_buf_8 fanout197 (.A(net200),
    .X(net197));
 sg13g2_buf_8 fanout198 (.A(net199),
    .X(net198));
 sg13g2_buf_8 fanout199 (.A(net200),
    .X(net199));
 sg13g2_buf_8 fanout200 (.A(net201),
    .X(net200));
 sg13g2_buf_8 fanout201 (.A(rst_n),
    .X(net201));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_sujanreddy_synapse_9 (.L_LO(net9));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_4_0_0_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_4_1_0_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_4_2_0_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_4_3_0_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_4_4_0_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_4_5_0_clk));
 sg13g2_buf_1 clkload6 (.A(clknet_4_6_0_clk));
 sg13g2_buf_1 clkload7 (.A(clknet_4_7_0_clk));
 sg13g2_buf_1 clkload8 (.A(clknet_4_8_0_clk));
 sg13g2_buf_1 clkload9 (.A(clknet_4_10_0_clk));
 sg13g2_buf_1 clkload10 (.A(clknet_4_11_0_clk));
 sg13g2_buf_1 clkload11 (.A(clknet_4_12_0_clk));
 sg13g2_buf_1 clkload12 (.A(clknet_4_13_0_clk));
 sg13g2_buf_1 clkload13 (.A(clknet_4_14_0_clk));
 sg13g2_buf_1 clkload14 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\controller_inst.sck_d1 ),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold2 (.A(\controller_inst.sck_d2 ),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0008_),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0039_),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold5 (.A(\controller_inst.data_reg1[0] ),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0065_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold7 (.A(\controller_inst.data_reg1[1] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0066_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold9 (.A(\controller_inst.shift_reg_in[7] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0064_),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold11 (.A(\controller_inst.shift_reg_out[3] ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold12 (.A(\controller_inst.shift_reg_out[2] ),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold13 (.A(\controller_inst.shift_reg_out[0] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold14 (.A(\controller_inst.shift_reg_out[1] ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold15 (.A(\controller_inst.pulse_width[15] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0072_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold17 (.A(\controller_inst.shift_reg_in[3] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0060_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold19 (.A(\controller_inst.shift_reg_in[5] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0062_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold21 (.A(\controller_inst.shift_reg_out[5] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0016_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold23 (.A(\controller_inst.shift_reg_out[7] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0722_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0089_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold26 (.A(\controller_inst.pulse_counter[4] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0045_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold28 (.A(\controller_inst.bit_cnt[1] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0178_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0028_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold31 (.A(\controller_inst.data_reg1[7] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold32 (.A(\controller_inst.cmd_reg[5] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold33 (.A(\controller_inst.bit_cnt[0] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0027_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0001_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0040_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold37 (.A(\controller_inst.shift_reg_in[6] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0063_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold39 (.A(\controller_inst.cmd_reg[6] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold40 (.A(\controller_inst.cmd_reg[7] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold41 (.A(\controller_inst.pulse_counter[5] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0046_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold43 (.A(\controller_inst.shift_reg_out[6] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0017_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold45 (.A(uio_out[4]),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0098_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0009_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0181_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0029_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold50 (.A(\controller_inst.cmd_reg[4] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0085_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold52 (.A(uio_out[1]),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold53 (.A(\controller_inst.prog_done ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0030_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold55 (.A(uio_out[5]),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0099_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold57 (.A(\controller_inst.pulse_counter[7] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0048_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold59 (.A(\controller_inst.pulse_counter[14] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0055_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold61 (.A(uio_out[6]),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0100_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold63 (.A(uio_out[7]),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0101_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold65 (.A(uio_out[3]),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0097_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold67 (.A(\controller_inst.state[2] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold68 (.A(uio_out[2]),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0096_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold70 (.A(\controller_inst.pulse_counter[1] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0042_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold72 (.A(\controller_inst.pulse_counter[11] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0052_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold74 (.A(\controller_inst.pulse_counter[15] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0056_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold76 (.A(\controller_inst.pulse_counter[3] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0044_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold78 (.A(\controller_inst.pulse_counter[10] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0051_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold80 (.A(\controller_inst.pulse_counter[13] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0054_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold82 (.A(\controller_inst.pulse_counter[9] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0050_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold84 (.A(uio_out[0]),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0094_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold86 (.A(\controller_inst.pulse_width[14] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0071_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold88 (.A(\controller_inst.shift_reg_in[0] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold89 (.A(\controller_inst.data_reg1[4] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0023_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold91 (.A(\controller_inst.pulse_width[12] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold92 (.A(\controller_inst.data_reg1[3] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0068_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold94 (.A(\controller_inst.pulse_width[13] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0070_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold96 (.A(\controller_inst.data_reg1[2] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0067_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold98 (.A(\controller_inst.pulse_counter[8] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0049_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold100 (.A(\controller_inst.byte_ready ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold101 (.A(\controller_inst.shift_reg_in[2] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold102 (.A(\controller_inst.pulse_counter[2] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0043_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold104 (.A(\controller_inst.pulse_counter[12] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0053_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold106 (.A(\controller_inst.cmd_reg[1] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0082_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold108 (.A(\controller_inst.cmd_reg[3] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold109 (.A(\controller_inst.cmd_reg[0] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold110 (.A(\controller_inst.sck_d3 ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold111 (.A(\controller_inst.shift_reg_in[1] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold112 (.A(\controller_inst.data_reg2[1] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold113 (.A(\controller_inst.data_reg2[7] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold114 (.A(\controller_inst.pulse_counter[6] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0047_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold116 (.A(\controller_inst.pulse_width[1] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold117 (.A(\controller_inst.cmd_reg[2] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold118 (.A(\controller_inst.state[3] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0207_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold120 (.A(\controller_inst.data_reg1[5] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold121 (.A(\controller_inst.shift_reg_in[4] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0077_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold123 (.A(\controller_inst.pulse_width[2] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold124 (.A(\controller_inst.data_reg2[3] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold125 (.A(\controller_inst.data_reg1[6] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold126 (.A(\controller_inst.data_reg2[5] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold127 (.A(\controller_inst.pulse_width[4] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold128 (.A(\controller_inst.data_reg2[2] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold129 (.A(\controller_inst.bit_cnt[2] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold130 (.A(\controller_inst.data_reg2[6] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold131 (.A(\controller_inst.pulse_width[0] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold132 (.A(\controller_inst.data_reg2[0] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold133 (.A(\controller_inst.pulse_counter[0] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0041_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold135 (.A(\controller_inst.state[1] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold136 (.A(\controller_inst.state[0] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold137 (.A(\controller_inst.state[1] ),
    .X(net221));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_fill_2 FILLER_6_77 ();
 sg13g2_fill_1 FILLER_6_79 ();
 sg13g2_decap_8 FILLER_6_85 ();
 sg13g2_decap_8 FILLER_6_92 ();
 sg13g2_decap_8 FILLER_6_99 ();
 sg13g2_decap_8 FILLER_6_106 ();
 sg13g2_decap_8 FILLER_6_118 ();
 sg13g2_fill_2 FILLER_6_125 ();
 sg13g2_decap_8 FILLER_6_135 ();
 sg13g2_decap_8 FILLER_6_142 ();
 sg13g2_decap_8 FILLER_6_149 ();
 sg13g2_decap_8 FILLER_6_156 ();
 sg13g2_decap_8 FILLER_6_163 ();
 sg13g2_decap_8 FILLER_6_170 ();
 sg13g2_decap_8 FILLER_6_177 ();
 sg13g2_decap_8 FILLER_6_184 ();
 sg13g2_decap_8 FILLER_6_191 ();
 sg13g2_fill_2 FILLER_6_198 ();
 sg13g2_fill_1 FILLER_6_200 ();
 sg13g2_decap_8 FILLER_6_206 ();
 sg13g2_decap_8 FILLER_6_213 ();
 sg13g2_decap_8 FILLER_6_220 ();
 sg13g2_decap_8 FILLER_6_227 ();
 sg13g2_decap_8 FILLER_6_234 ();
 sg13g2_decap_8 FILLER_6_241 ();
 sg13g2_decap_8 FILLER_6_248 ();
 sg13g2_decap_8 FILLER_6_255 ();
 sg13g2_decap_8 FILLER_6_262 ();
 sg13g2_decap_8 FILLER_6_269 ();
 sg13g2_decap_8 FILLER_6_276 ();
 sg13g2_decap_8 FILLER_6_283 ();
 sg13g2_decap_8 FILLER_6_290 ();
 sg13g2_decap_8 FILLER_6_297 ();
 sg13g2_decap_8 FILLER_6_304 ();
 sg13g2_decap_8 FILLER_6_311 ();
 sg13g2_decap_8 FILLER_6_318 ();
 sg13g2_decap_8 FILLER_6_325 ();
 sg13g2_decap_8 FILLER_6_332 ();
 sg13g2_decap_8 FILLER_6_339 ();
 sg13g2_decap_8 FILLER_6_346 ();
 sg13g2_decap_8 FILLER_6_353 ();
 sg13g2_decap_8 FILLER_6_360 ();
 sg13g2_decap_8 FILLER_6_367 ();
 sg13g2_decap_8 FILLER_6_374 ();
 sg13g2_decap_8 FILLER_6_381 ();
 sg13g2_decap_8 FILLER_6_388 ();
 sg13g2_decap_8 FILLER_6_395 ();
 sg13g2_decap_8 FILLER_6_402 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_fill_2 FILLER_7_56 ();
 sg13g2_fill_1 FILLER_7_58 ();
 sg13g2_decap_8 FILLER_7_64 ();
 sg13g2_fill_1 FILLER_7_71 ();
 sg13g2_decap_8 FILLER_7_92 ();
 sg13g2_fill_1 FILLER_7_99 ();
 sg13g2_fill_1 FILLER_7_121 ();
 sg13g2_decap_8 FILLER_7_143 ();
 sg13g2_decap_4 FILLER_7_150 ();
 sg13g2_fill_1 FILLER_7_154 ();
 sg13g2_decap_4 FILLER_7_168 ();
 sg13g2_fill_1 FILLER_7_172 ();
 sg13g2_decap_4 FILLER_7_178 ();
 sg13g2_fill_2 FILLER_7_182 ();
 sg13g2_fill_2 FILLER_7_197 ();
 sg13g2_fill_1 FILLER_7_199 ();
 sg13g2_decap_8 FILLER_7_213 ();
 sg13g2_decap_8 FILLER_7_220 ();
 sg13g2_decap_8 FILLER_7_227 ();
 sg13g2_decap_4 FILLER_7_234 ();
 sg13g2_decap_8 FILLER_7_242 ();
 sg13g2_decap_4 FILLER_7_249 ();
 sg13g2_fill_2 FILLER_7_253 ();
 sg13g2_decap_8 FILLER_7_260 ();
 sg13g2_decap_8 FILLER_7_267 ();
 sg13g2_decap_8 FILLER_7_274 ();
 sg13g2_decap_8 FILLER_7_281 ();
 sg13g2_decap_8 FILLER_7_288 ();
 sg13g2_decap_8 FILLER_7_295 ();
 sg13g2_decap_8 FILLER_7_302 ();
 sg13g2_fill_2 FILLER_7_309 ();
 sg13g2_fill_1 FILLER_7_311 ();
 sg13g2_decap_8 FILLER_7_321 ();
 sg13g2_decap_8 FILLER_7_328 ();
 sg13g2_decap_8 FILLER_7_335 ();
 sg13g2_decap_8 FILLER_7_342 ();
 sg13g2_decap_8 FILLER_7_349 ();
 sg13g2_decap_8 FILLER_7_356 ();
 sg13g2_decap_8 FILLER_7_363 ();
 sg13g2_decap_8 FILLER_7_370 ();
 sg13g2_decap_8 FILLER_7_377 ();
 sg13g2_decap_8 FILLER_7_384 ();
 sg13g2_decap_8 FILLER_7_391 ();
 sg13g2_decap_8 FILLER_7_398 ();
 sg13g2_decap_4 FILLER_7_405 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_4 FILLER_8_35 ();
 sg13g2_fill_1 FILLER_8_39 ();
 sg13g2_fill_2 FILLER_8_45 ();
 sg13g2_fill_1 FILLER_8_47 ();
 sg13g2_decap_8 FILLER_8_68 ();
 sg13g2_fill_2 FILLER_8_75 ();
 sg13g2_decap_8 FILLER_8_90 ();
 sg13g2_decap_8 FILLER_8_97 ();
 sg13g2_fill_2 FILLER_8_104 ();
 sg13g2_decap_8 FILLER_8_123 ();
 sg13g2_decap_8 FILLER_8_130 ();
 sg13g2_decap_4 FILLER_8_137 ();
 sg13g2_fill_2 FILLER_8_154 ();
 sg13g2_fill_2 FILLER_8_172 ();
 sg13g2_decap_4 FILLER_8_182 ();
 sg13g2_fill_2 FILLER_8_198 ();
 sg13g2_decap_8 FILLER_8_204 ();
 sg13g2_fill_2 FILLER_8_211 ();
 sg13g2_fill_2 FILLER_8_218 ();
 sg13g2_fill_1 FILLER_8_220 ();
 sg13g2_fill_2 FILLER_8_234 ();
 sg13g2_fill_1 FILLER_8_236 ();
 sg13g2_fill_2 FILLER_8_263 ();
 sg13g2_decap_8 FILLER_8_275 ();
 sg13g2_fill_2 FILLER_8_282 ();
 sg13g2_fill_2 FILLER_8_287 ();
 sg13g2_fill_1 FILLER_8_289 ();
 sg13g2_decap_8 FILLER_8_300 ();
 sg13g2_fill_2 FILLER_8_340 ();
 sg13g2_fill_1 FILLER_8_347 ();
 sg13g2_decap_8 FILLER_8_363 ();
 sg13g2_decap_8 FILLER_8_370 ();
 sg13g2_decap_8 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_4 FILLER_9_14 ();
 sg13g2_decap_4 FILLER_9_52 ();
 sg13g2_fill_1 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_65 ();
 sg13g2_fill_2 FILLER_9_85 ();
 sg13g2_decap_8 FILLER_9_92 ();
 sg13g2_fill_2 FILLER_9_99 ();
 sg13g2_fill_2 FILLER_9_118 ();
 sg13g2_decap_8 FILLER_9_125 ();
 sg13g2_fill_2 FILLER_9_132 ();
 sg13g2_fill_1 FILLER_9_134 ();
 sg13g2_decap_8 FILLER_9_145 ();
 sg13g2_fill_2 FILLER_9_152 ();
 sg13g2_fill_1 FILLER_9_154 ();
 sg13g2_fill_1 FILLER_9_160 ();
 sg13g2_fill_1 FILLER_9_178 ();
 sg13g2_fill_1 FILLER_9_197 ();
 sg13g2_fill_2 FILLER_9_206 ();
 sg13g2_fill_2 FILLER_9_229 ();
 sg13g2_decap_8 FILLER_9_239 ();
 sg13g2_decap_8 FILLER_9_246 ();
 sg13g2_fill_2 FILLER_9_253 ();
 sg13g2_fill_1 FILLER_9_255 ();
 sg13g2_fill_2 FILLER_9_289 ();
 sg13g2_decap_8 FILLER_9_298 ();
 sg13g2_decap_4 FILLER_9_305 ();
 sg13g2_fill_2 FILLER_9_325 ();
 sg13g2_fill_1 FILLER_9_346 ();
 sg13g2_decap_8 FILLER_9_383 ();
 sg13g2_decap_8 FILLER_9_390 ();
 sg13g2_decap_8 FILLER_9_397 ();
 sg13g2_decap_4 FILLER_9_404 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_4 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_4 ();
 sg13g2_decap_4 FILLER_10_27 ();
 sg13g2_fill_2 FILLER_10_31 ();
 sg13g2_decap_8 FILLER_10_51 ();
 sg13g2_decap_4 FILLER_10_58 ();
 sg13g2_fill_1 FILLER_10_62 ();
 sg13g2_fill_2 FILLER_10_76 ();
 sg13g2_decap_8 FILLER_10_83 ();
 sg13g2_decap_8 FILLER_10_90 ();
 sg13g2_fill_2 FILLER_10_112 ();
 sg13g2_fill_1 FILLER_10_114 ();
 sg13g2_fill_2 FILLER_10_123 ();
 sg13g2_fill_1 FILLER_10_125 ();
 sg13g2_fill_1 FILLER_10_142 ();
 sg13g2_decap_8 FILLER_10_151 ();
 sg13g2_decap_8 FILLER_10_158 ();
 sg13g2_decap_4 FILLER_10_165 ();
 sg13g2_fill_1 FILLER_10_169 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_fill_2 FILLER_10_194 ();
 sg13g2_fill_1 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_202 ();
 sg13g2_decap_8 FILLER_10_209 ();
 sg13g2_fill_1 FILLER_10_216 ();
 sg13g2_decap_8 FILLER_10_226 ();
 sg13g2_decap_4 FILLER_10_233 ();
 sg13g2_fill_2 FILLER_10_237 ();
 sg13g2_decap_8 FILLER_10_256 ();
 sg13g2_decap_8 FILLER_10_263 ();
 sg13g2_fill_2 FILLER_10_270 ();
 sg13g2_decap_8 FILLER_10_276 ();
 sg13g2_decap_8 FILLER_10_297 ();
 sg13g2_fill_1 FILLER_10_327 ();
 sg13g2_decap_4 FILLER_10_343 ();
 sg13g2_fill_2 FILLER_10_347 ();
 sg13g2_decap_8 FILLER_10_360 ();
 sg13g2_fill_2 FILLER_10_367 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_4 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_4 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_fill_1 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_30 ();
 sg13g2_decap_8 FILLER_11_37 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_fill_1 FILLER_11_76 ();
 sg13g2_decap_4 FILLER_11_90 ();
 sg13g2_fill_2 FILLER_11_99 ();
 sg13g2_fill_1 FILLER_11_101 ();
 sg13g2_fill_2 FILLER_11_110 ();
 sg13g2_decap_8 FILLER_11_117 ();
 sg13g2_decap_8 FILLER_11_124 ();
 sg13g2_fill_2 FILLER_11_131 ();
 sg13g2_fill_1 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_144 ();
 sg13g2_decap_4 FILLER_11_151 ();
 sg13g2_fill_1 FILLER_11_155 ();
 sg13g2_decap_4 FILLER_11_181 ();
 sg13g2_fill_2 FILLER_11_185 ();
 sg13g2_decap_8 FILLER_11_199 ();
 sg13g2_fill_2 FILLER_11_206 ();
 sg13g2_fill_1 FILLER_11_221 ();
 sg13g2_decap_4 FILLER_11_230 ();
 sg13g2_decap_4 FILLER_11_247 ();
 sg13g2_fill_2 FILLER_11_259 ();
 sg13g2_fill_2 FILLER_11_279 ();
 sg13g2_fill_1 FILLER_11_298 ();
 sg13g2_decap_8 FILLER_11_304 ();
 sg13g2_fill_2 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_383 ();
 sg13g2_decap_8 FILLER_11_390 ();
 sg13g2_decap_8 FILLER_11_397 ();
 sg13g2_decap_4 FILLER_11_404 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_4 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_4 ();
 sg13g2_decap_4 FILLER_12_13 ();
 sg13g2_decap_4 FILLER_12_30 ();
 sg13g2_fill_2 FILLER_12_47 ();
 sg13g2_fill_1 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_59 ();
 sg13g2_fill_1 FILLER_12_66 ();
 sg13g2_fill_2 FILLER_12_72 ();
 sg13g2_fill_1 FILLER_12_74 ();
 sg13g2_fill_2 FILLER_12_87 ();
 sg13g2_fill_2 FILLER_12_102 ();
 sg13g2_fill_1 FILLER_12_104 ();
 sg13g2_decap_8 FILLER_12_118 ();
 sg13g2_fill_2 FILLER_12_125 ();
 sg13g2_fill_1 FILLER_12_127 ();
 sg13g2_fill_2 FILLER_12_141 ();
 sg13g2_fill_1 FILLER_12_143 ();
 sg13g2_fill_1 FILLER_12_157 ();
 sg13g2_decap_4 FILLER_12_171 ();
 sg13g2_fill_1 FILLER_12_175 ();
 sg13g2_fill_2 FILLER_12_181 ();
 sg13g2_decap_8 FILLER_12_205 ();
 sg13g2_decap_4 FILLER_12_212 ();
 sg13g2_decap_8 FILLER_12_237 ();
 sg13g2_decap_4 FILLER_12_244 ();
 sg13g2_fill_1 FILLER_12_248 ();
 sg13g2_decap_8 FILLER_12_262 ();
 sg13g2_fill_2 FILLER_12_269 ();
 sg13g2_fill_1 FILLER_12_271 ();
 sg13g2_decap_8 FILLER_12_276 ();
 sg13g2_decap_4 FILLER_12_283 ();
 sg13g2_fill_2 FILLER_12_287 ();
 sg13g2_fill_2 FILLER_12_294 ();
 sg13g2_fill_1 FILLER_12_296 ();
 sg13g2_fill_2 FILLER_12_302 ();
 sg13g2_decap_8 FILLER_12_316 ();
 sg13g2_decap_4 FILLER_12_323 ();
 sg13g2_fill_2 FILLER_12_364 ();
 sg13g2_fill_1 FILLER_12_366 ();
 sg13g2_decap_8 FILLER_12_376 ();
 sg13g2_decap_8 FILLER_12_383 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_12 ();
 sg13g2_fill_1 FILLER_13_16 ();
 sg13g2_fill_2 FILLER_13_24 ();
 sg13g2_decap_4 FILLER_13_36 ();
 sg13g2_decap_4 FILLER_13_58 ();
 sg13g2_fill_1 FILLER_13_62 ();
 sg13g2_decap_8 FILLER_13_71 ();
 sg13g2_fill_2 FILLER_13_78 ();
 sg13g2_fill_1 FILLER_13_80 ();
 sg13g2_fill_1 FILLER_13_86 ();
 sg13g2_decap_8 FILLER_13_95 ();
 sg13g2_decap_4 FILLER_13_102 ();
 sg13g2_fill_1 FILLER_13_106 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_4 FILLER_13_133 ();
 sg13g2_fill_1 FILLER_13_137 ();
 sg13g2_fill_2 FILLER_13_155 ();
 sg13g2_fill_1 FILLER_13_157 ();
 sg13g2_decap_4 FILLER_13_180 ();
 sg13g2_decap_8 FILLER_13_193 ();
 sg13g2_fill_2 FILLER_13_200 ();
 sg13g2_fill_1 FILLER_13_202 ();
 sg13g2_decap_8 FILLER_13_208 ();
 sg13g2_decap_8 FILLER_13_215 ();
 sg13g2_fill_1 FILLER_13_222 ();
 sg13g2_fill_1 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_251 ();
 sg13g2_fill_2 FILLER_13_258 ();
 sg13g2_decap_8 FILLER_13_272 ();
 sg13g2_fill_2 FILLER_13_289 ();
 sg13g2_fill_1 FILLER_13_291 ();
 sg13g2_decap_4 FILLER_13_311 ();
 sg13g2_fill_1 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_23 ();
 sg13g2_fill_2 FILLER_14_39 ();
 sg13g2_decap_4 FILLER_14_65 ();
 sg13g2_fill_1 FILLER_14_69 ();
 sg13g2_decap_8 FILLER_14_92 ();
 sg13g2_decap_8 FILLER_14_99 ();
 sg13g2_fill_1 FILLER_14_106 ();
 sg13g2_decap_4 FILLER_14_125 ();
 sg13g2_fill_2 FILLER_14_129 ();
 sg13g2_fill_1 FILLER_14_150 ();
 sg13g2_decap_8 FILLER_14_156 ();
 sg13g2_fill_1 FILLER_14_163 ();
 sg13g2_fill_1 FILLER_14_177 ();
 sg13g2_decap_4 FILLER_14_199 ();
 sg13g2_fill_1 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_225 ();
 sg13g2_fill_1 FILLER_14_236 ();
 sg13g2_fill_2 FILLER_14_245 ();
 sg13g2_fill_2 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_285 ();
 sg13g2_fill_2 FILLER_14_292 ();
 sg13g2_decap_8 FILLER_14_309 ();
 sg13g2_decap_4 FILLER_14_316 ();
 sg13g2_decap_8 FILLER_14_384 ();
 sg13g2_decap_8 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_398 ();
 sg13g2_decap_4 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_4 FILLER_15_7 ();
 sg13g2_fill_2 FILLER_15_11 ();
 sg13g2_fill_2 FILLER_15_21 ();
 sg13g2_fill_1 FILLER_15_23 ();
 sg13g2_decap_4 FILLER_15_38 ();
 sg13g2_fill_2 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_58 ();
 sg13g2_decap_8 FILLER_15_65 ();
 sg13g2_decap_4 FILLER_15_72 ();
 sg13g2_fill_1 FILLER_15_76 ();
 sg13g2_decap_8 FILLER_15_86 ();
 sg13g2_decap_8 FILLER_15_101 ();
 sg13g2_fill_2 FILLER_15_108 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_fill_1 FILLER_15_126 ();
 sg13g2_fill_2 FILLER_15_137 ();
 sg13g2_fill_2 FILLER_15_147 ();
 sg13g2_decap_4 FILLER_15_163 ();
 sg13g2_fill_2 FILLER_15_167 ();
 sg13g2_decap_8 FILLER_15_174 ();
 sg13g2_decap_4 FILLER_15_181 ();
 sg13g2_decap_8 FILLER_15_202 ();
 sg13g2_decap_4 FILLER_15_209 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_fill_2 FILLER_15_224 ();
 sg13g2_fill_1 FILLER_15_226 ();
 sg13g2_fill_1 FILLER_15_231 ();
 sg13g2_decap_4 FILLER_15_241 ();
 sg13g2_fill_1 FILLER_15_245 ();
 sg13g2_fill_2 FILLER_15_251 ();
 sg13g2_fill_1 FILLER_15_253 ();
 sg13g2_decap_4 FILLER_15_270 ();
 sg13g2_fill_2 FILLER_15_274 ();
 sg13g2_decap_4 FILLER_15_284 ();
 sg13g2_fill_2 FILLER_15_288 ();
 sg13g2_decap_4 FILLER_15_298 ();
 sg13g2_decap_8 FILLER_15_314 ();
 sg13g2_fill_1 FILLER_15_321 ();
 sg13g2_fill_1 FILLER_15_338 ();
 sg13g2_fill_1 FILLER_15_347 ();
 sg13g2_decap_8 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_4 ();
 sg13g2_decap_8 FILLER_16_32 ();
 sg13g2_decap_4 FILLER_16_39 ();
 sg13g2_fill_2 FILLER_16_43 ();
 sg13g2_decap_4 FILLER_16_58 ();
 sg13g2_fill_2 FILLER_16_62 ();
 sg13g2_fill_2 FILLER_16_92 ();
 sg13g2_fill_1 FILLER_16_94 ();
 sg13g2_fill_2 FILLER_16_123 ();
 sg13g2_fill_2 FILLER_16_130 ();
 sg13g2_fill_1 FILLER_16_132 ();
 sg13g2_decap_4 FILLER_16_138 ();
 sg13g2_fill_2 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_165 ();
 sg13g2_fill_2 FILLER_16_172 ();
 sg13g2_fill_1 FILLER_16_178 ();
 sg13g2_fill_2 FILLER_16_191 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_fill_2 FILLER_16_203 ();
 sg13g2_fill_1 FILLER_16_205 ();
 sg13g2_fill_2 FILLER_16_210 ();
 sg13g2_fill_2 FILLER_16_220 ();
 sg13g2_fill_2 FILLER_16_235 ();
 sg13g2_fill_2 FILLER_16_245 ();
 sg13g2_fill_1 FILLER_16_247 ();
 sg13g2_decap_8 FILLER_16_256 ();
 sg13g2_decap_8 FILLER_16_263 ();
 sg13g2_fill_1 FILLER_16_283 ();
 sg13g2_decap_8 FILLER_16_293 ();
 sg13g2_fill_1 FILLER_16_300 ();
 sg13g2_fill_2 FILLER_16_311 ();
 sg13g2_fill_2 FILLER_16_340 ();
 sg13g2_decap_8 FILLER_16_388 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_fill_1 FILLER_17_16 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_fill_1 FILLER_17_28 ();
 sg13g2_decap_4 FILLER_17_41 ();
 sg13g2_fill_2 FILLER_17_53 ();
 sg13g2_fill_1 FILLER_17_55 ();
 sg13g2_decap_8 FILLER_17_66 ();
 sg13g2_decap_8 FILLER_17_73 ();
 sg13g2_decap_4 FILLER_17_80 ();
 sg13g2_fill_1 FILLER_17_84 ();
 sg13g2_fill_2 FILLER_17_95 ();
 sg13g2_decap_4 FILLER_17_141 ();
 sg13g2_fill_2 FILLER_17_145 ();
 sg13g2_fill_1 FILLER_17_154 ();
 sg13g2_fill_2 FILLER_17_175 ();
 sg13g2_fill_1 FILLER_17_177 ();
 sg13g2_decap_4 FILLER_17_187 ();
 sg13g2_fill_1 FILLER_17_191 ();
 sg13g2_decap_4 FILLER_17_197 ();
 sg13g2_fill_1 FILLER_17_201 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_4 FILLER_17_231 ();
 sg13g2_fill_2 FILLER_17_244 ();
 sg13g2_fill_2 FILLER_17_255 ();
 sg13g2_fill_1 FILLER_17_257 ();
 sg13g2_fill_1 FILLER_17_276 ();
 sg13g2_fill_2 FILLER_17_281 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_fill_2 FILLER_17_301 ();
 sg13g2_fill_1 FILLER_17_303 ();
 sg13g2_decap_8 FILLER_17_309 ();
 sg13g2_fill_1 FILLER_17_316 ();
 sg13g2_fill_1 FILLER_17_330 ();
 sg13g2_fill_1 FILLER_17_342 ();
 sg13g2_fill_2 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_373 ();
 sg13g2_decap_8 FILLER_17_380 ();
 sg13g2_decap_8 FILLER_17_387 ();
 sg13g2_decap_8 FILLER_17_394 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_7 ();
 sg13g2_fill_2 FILLER_18_16 ();
 sg13g2_decap_4 FILLER_18_22 ();
 sg13g2_fill_1 FILLER_18_26 ();
 sg13g2_fill_2 FILLER_18_43 ();
 sg13g2_decap_8 FILLER_18_57 ();
 sg13g2_decap_8 FILLER_18_64 ();
 sg13g2_decap_8 FILLER_18_71 ();
 sg13g2_fill_2 FILLER_18_78 ();
 sg13g2_fill_1 FILLER_18_93 ();
 sg13g2_decap_4 FILLER_18_126 ();
 sg13g2_fill_1 FILLER_18_156 ();
 sg13g2_fill_1 FILLER_18_170 ();
 sg13g2_decap_4 FILLER_18_199 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_4 FILLER_18_255 ();
 sg13g2_fill_1 FILLER_18_271 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_4 FILLER_18_287 ();
 sg13g2_fill_1 FILLER_18_291 ();
 sg13g2_decap_8 FILLER_18_318 ();
 sg13g2_fill_2 FILLER_18_325 ();
 sg13g2_decap_4 FILLER_18_336 ();
 sg13g2_fill_1 FILLER_18_367 ();
 sg13g2_decap_8 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_2 ();
 sg13g2_fill_2 FILLER_19_25 ();
 sg13g2_fill_2 FILLER_19_31 ();
 sg13g2_fill_2 FILLER_19_49 ();
 sg13g2_fill_1 FILLER_19_51 ();
 sg13g2_fill_2 FILLER_19_84 ();
 sg13g2_fill_1 FILLER_19_86 ();
 sg13g2_fill_1 FILLER_19_101 ();
 sg13g2_decap_4 FILLER_19_111 ();
 sg13g2_decap_8 FILLER_19_137 ();
 sg13g2_decap_4 FILLER_19_144 ();
 sg13g2_fill_2 FILLER_19_148 ();
 sg13g2_decap_8 FILLER_19_155 ();
 sg13g2_fill_2 FILLER_19_180 ();
 sg13g2_fill_2 FILLER_19_187 ();
 sg13g2_fill_1 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_200 ();
 sg13g2_fill_1 FILLER_19_207 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_fill_2 FILLER_19_238 ();
 sg13g2_fill_1 FILLER_19_240 ();
 sg13g2_decap_8 FILLER_19_254 ();
 sg13g2_decap_8 FILLER_19_261 ();
 sg13g2_fill_2 FILLER_19_268 ();
 sg13g2_fill_1 FILLER_19_275 ();
 sg13g2_fill_1 FILLER_19_281 ();
 sg13g2_decap_8 FILLER_19_295 ();
 sg13g2_fill_2 FILLER_19_302 ();
 sg13g2_decap_4 FILLER_19_314 ();
 sg13g2_fill_2 FILLER_19_318 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_34 ();
 sg13g2_fill_1 FILLER_20_41 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_fill_2 FILLER_20_77 ();
 sg13g2_decap_4 FILLER_20_92 ();
 sg13g2_fill_1 FILLER_20_123 ();
 sg13g2_decap_8 FILLER_20_152 ();
 sg13g2_decap_8 FILLER_20_159 ();
 sg13g2_fill_1 FILLER_20_166 ();
 sg13g2_fill_2 FILLER_20_180 ();
 sg13g2_fill_2 FILLER_20_190 ();
 sg13g2_fill_1 FILLER_20_192 ();
 sg13g2_fill_2 FILLER_20_201 ();
 sg13g2_fill_1 FILLER_20_203 ();
 sg13g2_fill_2 FILLER_20_220 ();
 sg13g2_decap_4 FILLER_20_235 ();
 sg13g2_fill_1 FILLER_20_239 ();
 sg13g2_decap_8 FILLER_20_246 ();
 sg13g2_fill_1 FILLER_20_253 ();
 sg13g2_fill_1 FILLER_20_258 ();
 sg13g2_decap_4 FILLER_20_264 ();
 sg13g2_decap_8 FILLER_20_284 ();
 sg13g2_decap_4 FILLER_20_291 ();
 sg13g2_fill_2 FILLER_20_295 ();
 sg13g2_decap_4 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_88 ();
 sg13g2_decap_8 FILLER_21_134 ();
 sg13g2_decap_8 FILLER_21_191 ();
 sg13g2_decap_4 FILLER_21_198 ();
 sg13g2_fill_1 FILLER_21_202 ();
 sg13g2_decap_4 FILLER_21_208 ();
 sg13g2_fill_2 FILLER_21_217 ();
 sg13g2_fill_1 FILLER_21_219 ();
 sg13g2_decap_4 FILLER_21_224 ();
 sg13g2_fill_2 FILLER_21_228 ();
 sg13g2_decap_4 FILLER_21_234 ();
 sg13g2_fill_1 FILLER_21_238 ();
 sg13g2_fill_2 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_268 ();
 sg13g2_decap_8 FILLER_21_275 ();
 sg13g2_fill_2 FILLER_21_282 ();
 sg13g2_fill_1 FILLER_21_284 ();
 sg13g2_decap_8 FILLER_21_298 ();
 sg13g2_decap_8 FILLER_21_305 ();
 sg13g2_fill_2 FILLER_21_312 ();
 sg13g2_fill_2 FILLER_21_340 ();
 sg13g2_fill_1 FILLER_21_353 ();
 sg13g2_decap_8 FILLER_21_391 ();
 sg13g2_decap_8 FILLER_21_398 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_fill_2 FILLER_22_36 ();
 sg13g2_fill_2 FILLER_22_111 ();
 sg13g2_decap_4 FILLER_22_171 ();
 sg13g2_decap_4 FILLER_22_188 ();
 sg13g2_fill_1 FILLER_22_192 ();
 sg13g2_fill_1 FILLER_22_223 ();
 sg13g2_fill_2 FILLER_22_246 ();
 sg13g2_fill_1 FILLER_22_248 ();
 sg13g2_decap_8 FILLER_22_253 ();
 sg13g2_decap_8 FILLER_22_260 ();
 sg13g2_fill_2 FILLER_22_267 ();
 sg13g2_fill_1 FILLER_22_269 ();
 sg13g2_fill_2 FILLER_22_275 ();
 sg13g2_decap_8 FILLER_22_289 ();
 sg13g2_fill_2 FILLER_22_296 ();
 sg13g2_decap_4 FILLER_22_313 ();
 sg13g2_fill_1 FILLER_22_317 ();
 sg13g2_fill_2 FILLER_22_351 ();
 sg13g2_fill_2 FILLER_22_362 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_52 ();
 sg13g2_decap_4 FILLER_23_76 ();
 sg13g2_fill_2 FILLER_23_80 ();
 sg13g2_fill_2 FILLER_23_95 ();
 sg13g2_decap_4 FILLER_23_120 ();
 sg13g2_decap_4 FILLER_23_134 ();
 sg13g2_fill_2 FILLER_23_138 ();
 sg13g2_decap_8 FILLER_23_180 ();
 sg13g2_fill_1 FILLER_23_187 ();
 sg13g2_fill_2 FILLER_23_247 ();
 sg13g2_fill_1 FILLER_23_249 ();
 sg13g2_fill_2 FILLER_23_255 ();
 sg13g2_fill_1 FILLER_23_257 ();
 sg13g2_decap_8 FILLER_23_278 ();
 sg13g2_fill_1 FILLER_23_285 ();
 sg13g2_decap_8 FILLER_23_300 ();
 sg13g2_fill_2 FILLER_23_307 ();
 sg13g2_fill_1 FILLER_23_309 ();
 sg13g2_fill_2 FILLER_23_323 ();
 sg13g2_fill_1 FILLER_23_325 ();
 sg13g2_fill_1 FILLER_23_335 ();
 sg13g2_fill_1 FILLER_23_349 ();
 sg13g2_fill_1 FILLER_23_355 ();
 sg13g2_decap_8 FILLER_23_390 ();
 sg13g2_decap_8 FILLER_23_397 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_fill_2 FILLER_24_14 ();
 sg13g2_decap_4 FILLER_24_26 ();
 sg13g2_fill_2 FILLER_24_86 ();
 sg13g2_fill_1 FILLER_24_88 ();
 sg13g2_fill_1 FILLER_24_122 ();
 sg13g2_fill_1 FILLER_24_136 ();
 sg13g2_fill_1 FILLER_24_150 ();
 sg13g2_decap_4 FILLER_24_169 ();
 sg13g2_decap_4 FILLER_24_196 ();
 sg13g2_fill_1 FILLER_24_200 ();
 sg13g2_decap_8 FILLER_24_205 ();
 sg13g2_decap_8 FILLER_24_212 ();
 sg13g2_fill_2 FILLER_24_219 ();
 sg13g2_decap_8 FILLER_24_230 ();
 sg13g2_fill_2 FILLER_24_237 ();
 sg13g2_fill_1 FILLER_24_251 ();
 sg13g2_decap_8 FILLER_24_260 ();
 sg13g2_fill_2 FILLER_24_267 ();
 sg13g2_fill_1 FILLER_24_269 ();
 sg13g2_fill_2 FILLER_24_285 ();
 sg13g2_fill_1 FILLER_24_287 ();
 sg13g2_decap_4 FILLER_24_301 ();
 sg13g2_fill_1 FILLER_24_305 ();
 sg13g2_decap_4 FILLER_24_322 ();
 sg13g2_fill_1 FILLER_24_352 ();
 sg13g2_decap_8 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_7 ();
 sg13g2_fill_2 FILLER_25_11 ();
 sg13g2_fill_2 FILLER_25_23 ();
 sg13g2_fill_1 FILLER_25_25 ();
 sg13g2_fill_2 FILLER_25_36 ();
 sg13g2_decap_8 FILLER_25_75 ();
 sg13g2_fill_2 FILLER_25_120 ();
 sg13g2_fill_1 FILLER_25_122 ();
 sg13g2_decap_4 FILLER_25_128 ();
 sg13g2_fill_1 FILLER_25_132 ();
 sg13g2_fill_1 FILLER_25_146 ();
 sg13g2_decap_4 FILLER_25_169 ();
 sg13g2_fill_2 FILLER_25_173 ();
 sg13g2_fill_2 FILLER_25_202 ();
 sg13g2_fill_1 FILLER_25_204 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_fill_1 FILLER_25_252 ();
 sg13g2_decap_4 FILLER_25_266 ();
 sg13g2_fill_1 FILLER_25_270 ();
 sg13g2_decap_8 FILLER_25_275 ();
 sg13g2_fill_1 FILLER_25_282 ();
 sg13g2_fill_2 FILLER_25_296 ();
 sg13g2_fill_1 FILLER_25_298 ();
 sg13g2_fill_2 FILLER_25_324 ();
 sg13g2_fill_2 FILLER_25_356 ();
 sg13g2_decap_8 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_29 ();
 sg13g2_fill_1 FILLER_26_33 ();
 sg13g2_fill_2 FILLER_26_141 ();
 sg13g2_fill_1 FILLER_26_180 ();
 sg13g2_decap_8 FILLER_26_191 ();
 sg13g2_decap_8 FILLER_26_198 ();
 sg13g2_fill_1 FILLER_26_205 ();
 sg13g2_fill_2 FILLER_26_233 ();
 sg13g2_fill_1 FILLER_26_235 ();
 sg13g2_fill_2 FILLER_26_246 ();
 sg13g2_decap_8 FILLER_26_296 ();
 sg13g2_fill_2 FILLER_26_303 ();
 sg13g2_decap_8 FILLER_26_377 ();
 sg13g2_decap_8 FILLER_26_384 ();
 sg13g2_decap_8 FILLER_26_391 ();
 sg13g2_decap_8 FILLER_26_398 ();
 sg13g2_decap_4 FILLER_26_405 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_24 ();
 sg13g2_fill_1 FILLER_27_26 ();
 sg13g2_decap_4 FILLER_27_41 ();
 sg13g2_fill_1 FILLER_27_54 ();
 sg13g2_decap_4 FILLER_27_102 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_fill_2 FILLER_27_171 ();
 sg13g2_fill_1 FILLER_27_173 ();
 sg13g2_decap_4 FILLER_27_223 ();
 sg13g2_fill_2 FILLER_27_227 ();
 sg13g2_decap_8 FILLER_27_244 ();
 sg13g2_fill_1 FILLER_27_251 ();
 sg13g2_fill_1 FILLER_27_269 ();
 sg13g2_decap_8 FILLER_27_277 ();
 sg13g2_fill_2 FILLER_27_284 ();
 sg13g2_fill_2 FILLER_27_292 ();
 sg13g2_decap_8 FILLER_27_304 ();
 sg13g2_decap_8 FILLER_27_311 ();
 sg13g2_fill_2 FILLER_27_318 ();
 sg13g2_fill_2 FILLER_27_350 ();
 sg13g2_decap_4 FILLER_27_361 ();
 sg13g2_fill_1 FILLER_27_365 ();
 sg13g2_decap_8 FILLER_27_375 ();
 sg13g2_decap_8 FILLER_27_382 ();
 sg13g2_decap_8 FILLER_27_389 ();
 sg13g2_decap_8 FILLER_27_396 ();
 sg13g2_decap_4 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_4 FILLER_28_27 ();
 sg13g2_fill_1 FILLER_28_31 ();
 sg13g2_fill_2 FILLER_28_87 ();
 sg13g2_fill_1 FILLER_28_149 ();
 sg13g2_decap_8 FILLER_28_188 ();
 sg13g2_decap_8 FILLER_28_195 ();
 sg13g2_decap_4 FILLER_28_202 ();
 sg13g2_fill_2 FILLER_28_239 ();
 sg13g2_fill_1 FILLER_28_241 ();
 sg13g2_fill_1 FILLER_28_249 ();
 sg13g2_fill_1 FILLER_28_266 ();
 sg13g2_fill_2 FILLER_28_302 ();
 sg13g2_decap_8 FILLER_28_383 ();
 sg13g2_decap_8 FILLER_28_390 ();
 sg13g2_decap_8 FILLER_28_397 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_17 ();
 sg13g2_fill_1 FILLER_29_29 ();
 sg13g2_fill_2 FILLER_29_44 ();
 sg13g2_fill_1 FILLER_29_46 ();
 sg13g2_fill_1 FILLER_29_60 ();
 sg13g2_fill_2 FILLER_29_78 ();
 sg13g2_fill_2 FILLER_29_111 ();
 sg13g2_fill_1 FILLER_29_123 ();
 sg13g2_decap_8 FILLER_29_143 ();
 sg13g2_decap_8 FILLER_29_169 ();
 sg13g2_decap_8 FILLER_29_176 ();
 sg13g2_fill_1 FILLER_29_183 ();
 sg13g2_fill_2 FILLER_29_199 ();
 sg13g2_decap_4 FILLER_29_213 ();
 sg13g2_fill_1 FILLER_29_217 ();
 sg13g2_fill_2 FILLER_29_222 ();
 sg13g2_fill_1 FILLER_29_224 ();
 sg13g2_fill_2 FILLER_29_243 ();
 sg13g2_fill_2 FILLER_29_249 ();
 sg13g2_fill_2 FILLER_29_257 ();
 sg13g2_fill_2 FILLER_29_272 ();
 sg13g2_fill_2 FILLER_29_291 ();
 sg13g2_fill_1 FILLER_29_293 ();
 sg13g2_fill_2 FILLER_29_307 ();
 sg13g2_decap_8 FILLER_29_382 ();
 sg13g2_decap_8 FILLER_29_389 ();
 sg13g2_decap_8 FILLER_29_396 ();
 sg13g2_decap_4 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_fill_2 FILLER_30_73 ();
 sg13g2_fill_2 FILLER_30_98 ();
 sg13g2_fill_2 FILLER_30_135 ();
 sg13g2_fill_1 FILLER_30_137 ();
 sg13g2_fill_1 FILLER_30_165 ();
 sg13g2_decap_4 FILLER_30_199 ();
 sg13g2_fill_1 FILLER_30_207 ();
 sg13g2_decap_4 FILLER_30_221 ();
 sg13g2_fill_2 FILLER_30_273 ();
 sg13g2_fill_1 FILLER_30_320 ();
 sg13g2_decap_8 FILLER_30_390 ();
 sg13g2_decap_8 FILLER_30_397 ();
 sg13g2_decap_4 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_24 ();
 sg13g2_fill_1 FILLER_31_26 ();
 sg13g2_fill_2 FILLER_31_80 ();
 sg13g2_fill_1 FILLER_31_82 ();
 sg13g2_fill_2 FILLER_31_94 ();
 sg13g2_fill_1 FILLER_31_96 ();
 sg13g2_decap_4 FILLER_31_106 ();
 sg13g2_decap_8 FILLER_31_115 ();
 sg13g2_decap_4 FILLER_31_122 ();
 sg13g2_decap_4 FILLER_31_137 ();
 sg13g2_fill_2 FILLER_31_141 ();
 sg13g2_fill_1 FILLER_31_156 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_fill_2 FILLER_31_196 ();
 sg13g2_fill_2 FILLER_31_210 ();
 sg13g2_fill_1 FILLER_31_212 ();
 sg13g2_decap_8 FILLER_31_218 ();
 sg13g2_decap_4 FILLER_31_225 ();
 sg13g2_fill_2 FILLER_31_229 ();
 sg13g2_fill_1 FILLER_31_239 ();
 sg13g2_fill_2 FILLER_31_280 ();
 sg13g2_fill_1 FILLER_31_328 ();
 sg13g2_fill_2 FILLER_31_342 ();
 sg13g2_fill_1 FILLER_31_344 ();
 sg13g2_fill_2 FILLER_31_370 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_4 FILLER_32_49 ();
 sg13g2_fill_1 FILLER_32_53 ();
 sg13g2_fill_2 FILLER_32_76 ();
 sg13g2_fill_2 FILLER_32_88 ();
 sg13g2_fill_1 FILLER_32_90 ();
 sg13g2_fill_2 FILLER_32_136 ();
 sg13g2_fill_1 FILLER_32_138 ();
 sg13g2_fill_2 FILLER_32_159 ();
 sg13g2_fill_1 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_184 ();
 sg13g2_decap_4 FILLER_32_191 ();
 sg13g2_fill_1 FILLER_32_195 ();
 sg13g2_fill_1 FILLER_32_201 ();
 sg13g2_decap_4 FILLER_32_210 ();
 sg13g2_fill_2 FILLER_32_249 ();
 sg13g2_fill_1 FILLER_32_251 ();
 sg13g2_fill_2 FILLER_32_333 ();
 sg13g2_fill_1 FILLER_32_335 ();
 sg13g2_fill_2 FILLER_32_341 ();
 sg13g2_fill_1 FILLER_32_356 ();
 sg13g2_fill_2 FILLER_32_380 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_11 ();
 sg13g2_decap_4 FILLER_33_22 ();
 sg13g2_fill_1 FILLER_33_26 ();
 sg13g2_fill_2 FILLER_33_94 ();
 sg13g2_fill_1 FILLER_33_96 ();
 sg13g2_fill_1 FILLER_33_101 ();
 sg13g2_decap_8 FILLER_33_108 ();
 sg13g2_decap_4 FILLER_33_147 ();
 sg13g2_fill_2 FILLER_33_151 ();
 sg13g2_decap_4 FILLER_33_181 ();
 sg13g2_fill_1 FILLER_33_185 ();
 sg13g2_decap_4 FILLER_33_211 ();
 sg13g2_fill_1 FILLER_33_215 ();
 sg13g2_fill_1 FILLER_33_225 ();
 sg13g2_fill_2 FILLER_33_236 ();
 sg13g2_fill_1 FILLER_33_257 ();
 sg13g2_fill_2 FILLER_33_263 ();
 sg13g2_fill_1 FILLER_33_265 ();
 sg13g2_fill_2 FILLER_33_301 ();
 sg13g2_decap_4 FILLER_33_316 ();
 sg13g2_fill_2 FILLER_33_320 ();
 sg13g2_fill_2 FILLER_33_359 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_36 ();
 sg13g2_decap_8 FILLER_34_43 ();
 sg13g2_fill_2 FILLER_34_50 ();
 sg13g2_fill_1 FILLER_34_52 ();
 sg13g2_fill_2 FILLER_34_83 ();
 sg13g2_fill_2 FILLER_34_99 ();
 sg13g2_fill_1 FILLER_34_101 ();
 sg13g2_fill_1 FILLER_34_129 ();
 sg13g2_fill_1 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_4 FILLER_34_182 ();
 sg13g2_fill_1 FILLER_34_191 ();
 sg13g2_decap_8 FILLER_34_212 ();
 sg13g2_decap_4 FILLER_34_219 ();
 sg13g2_fill_1 FILLER_34_223 ();
 sg13g2_fill_2 FILLER_34_253 ();
 sg13g2_fill_1 FILLER_34_255 ();
 sg13g2_fill_2 FILLER_34_265 ();
 sg13g2_fill_1 FILLER_34_267 ();
 sg13g2_fill_1 FILLER_34_298 ();
 sg13g2_fill_1 FILLER_34_322 ();
 sg13g2_fill_1 FILLER_34_388 ();
 sg13g2_decap_4 FILLER_34_396 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_7 ();
 sg13g2_fill_1 FILLER_35_9 ();
 sg13g2_fill_2 FILLER_35_147 ();
 sg13g2_fill_1 FILLER_35_149 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_fill_1 FILLER_35_189 ();
 sg13g2_fill_2 FILLER_35_195 ();
 sg13g2_fill_1 FILLER_35_197 ();
 sg13g2_decap_4 FILLER_35_216 ();
 sg13g2_fill_2 FILLER_35_220 ();
 sg13g2_decap_4 FILLER_35_227 ();
 sg13g2_fill_1 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_273 ();
 sg13g2_decap_4 FILLER_35_280 ();
 sg13g2_fill_1 FILLER_35_284 ();
 sg13g2_fill_2 FILLER_35_322 ();
 sg13g2_fill_2 FILLER_35_349 ();
 sg13g2_fill_1 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_30 ();
 sg13g2_decap_8 FILLER_36_37 ();
 sg13g2_decap_4 FILLER_36_44 ();
 sg13g2_fill_1 FILLER_36_48 ();
 sg13g2_fill_2 FILLER_36_145 ();
 sg13g2_fill_1 FILLER_36_147 ();
 sg13g2_fill_1 FILLER_36_167 ();
 sg13g2_fill_1 FILLER_36_206 ();
 sg13g2_decap_8 FILLER_36_216 ();
 sg13g2_fill_1 FILLER_36_223 ();
 sg13g2_fill_1 FILLER_36_238 ();
 sg13g2_decap_4 FILLER_36_251 ();
 sg13g2_fill_2 FILLER_36_255 ();
 sg13g2_decap_4 FILLER_36_270 ();
 sg13g2_fill_1 FILLER_36_274 ();
 sg13g2_fill_2 FILLER_36_285 ();
 sg13g2_fill_1 FILLER_36_287 ();
 sg13g2_fill_1 FILLER_36_297 ();
 sg13g2_fill_2 FILLER_36_333 ();
 sg13g2_fill_2 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_4 FILLER_37_49 ();
 sg13g2_fill_2 FILLER_37_53 ();
 sg13g2_fill_2 FILLER_37_197 ();
 sg13g2_fill_1 FILLER_37_199 ();
 sg13g2_fill_2 FILLER_37_204 ();
 sg13g2_fill_1 FILLER_37_241 ();
 sg13g2_decap_8 FILLER_37_256 ();
 sg13g2_decap_4 FILLER_37_263 ();
 sg13g2_fill_1 FILLER_37_267 ();
 sg13g2_fill_2 FILLER_37_347 ();
 sg13g2_decap_4 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_4 FILLER_38_42 ();
 sg13g2_fill_2 FILLER_38_46 ();
 sg13g2_fill_2 FILLER_38_73 ();
 sg13g2_fill_1 FILLER_38_75 ();
 sg13g2_fill_1 FILLER_38_81 ();
 sg13g2_fill_2 FILLER_38_91 ();
 sg13g2_fill_2 FILLER_38_142 ();
 sg13g2_decap_8 FILLER_38_153 ();
 sg13g2_decap_4 FILLER_38_160 ();
 sg13g2_fill_2 FILLER_38_164 ();
 sg13g2_fill_2 FILLER_38_175 ();
 sg13g2_fill_1 FILLER_38_177 ();
 sg13g2_fill_2 FILLER_38_206 ();
 sg13g2_decap_8 FILLER_38_212 ();
 sg13g2_decap_8 FILLER_38_219 ();
 sg13g2_decap_4 FILLER_38_226 ();
 sg13g2_fill_2 FILLER_38_230 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_decap_4 FILLER_38_243 ();
 sg13g2_fill_2 FILLER_38_274 ();
 sg13g2_fill_1 FILLER_38_276 ();
 sg13g2_fill_1 FILLER_38_343 ();
 sg13g2_fill_1 FILLER_38_349 ();
 sg13g2_fill_2 FILLER_38_380 ();
 sg13g2_fill_1 FILLER_38_382 ();
 sg13g2_decap_4 FILLER_38_396 ();
 assign uio_oe[0] = net13;
 assign uio_oe[1] = net14;
 assign uio_oe[2] = net15;
 assign uio_oe[3] = net16;
 assign uio_oe[4] = net17;
 assign uio_oe[5] = net18;
 assign uio_oe[6] = net19;
 assign uio_oe[7] = net20;
 assign uo_out[4] = net9;
 assign uo_out[5] = net10;
 assign uo_out[6] = net11;
 assign uo_out[7] = net12;
endmodule
