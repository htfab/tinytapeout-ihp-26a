module tt_um_themightyduckofdoom_bitserial_collatz_checker (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire \bit_counter_q[0] ;
 wire \bit_counter_q[1] ;
 wire \bit_counter_q[2] ;
 wire \bit_counter_q[3] ;
 wire \bit_counter_q[4] ;
 wire \bit_counter_q[5] ;
 wire \bit_counter_q[6] ;
 wire \bit_counter_q[7] ;
 wire \bit_counter_q[8] ;
 wire \bit_counter_q[9] ;
 wire carry_q;
 wire finished_q;
 wire \i_main_reg.data_d[0] ;
 wire \i_main_reg.data_d[100] ;
 wire \i_main_reg.data_d[101] ;
 wire \i_main_reg.data_d[102] ;
 wire \i_main_reg.data_d[103] ;
 wire \i_main_reg.data_d[104] ;
 wire \i_main_reg.data_d[105] ;
 wire \i_main_reg.data_d[106] ;
 wire \i_main_reg.data_d[107] ;
 wire \i_main_reg.data_d[108] ;
 wire \i_main_reg.data_d[109] ;
 wire \i_main_reg.data_d[10] ;
 wire \i_main_reg.data_d[110] ;
 wire \i_main_reg.data_d[111] ;
 wire \i_main_reg.data_d[112] ;
 wire \i_main_reg.data_d[113] ;
 wire \i_main_reg.data_d[114] ;
 wire \i_main_reg.data_d[115] ;
 wire \i_main_reg.data_d[116] ;
 wire \i_main_reg.data_d[117] ;
 wire \i_main_reg.data_d[118] ;
 wire \i_main_reg.data_d[119] ;
 wire \i_main_reg.data_d[11] ;
 wire \i_main_reg.data_d[120] ;
 wire \i_main_reg.data_d[121] ;
 wire \i_main_reg.data_d[122] ;
 wire \i_main_reg.data_d[123] ;
 wire \i_main_reg.data_d[124] ;
 wire \i_main_reg.data_d[125] ;
 wire \i_main_reg.data_d[126] ;
 wire \i_main_reg.data_d[127] ;
 wire \i_main_reg.data_d[128] ;
 wire \i_main_reg.data_d[129] ;
 wire \i_main_reg.data_d[12] ;
 wire \i_main_reg.data_d[130] ;
 wire \i_main_reg.data_d[131] ;
 wire \i_main_reg.data_d[132] ;
 wire \i_main_reg.data_d[133] ;
 wire \i_main_reg.data_d[134] ;
 wire \i_main_reg.data_d[135] ;
 wire \i_main_reg.data_d[136] ;
 wire \i_main_reg.data_d[137] ;
 wire \i_main_reg.data_d[138] ;
 wire \i_main_reg.data_d[139] ;
 wire \i_main_reg.data_d[13] ;
 wire \i_main_reg.data_d[140] ;
 wire \i_main_reg.data_d[141] ;
 wire \i_main_reg.data_d[142] ;
 wire \i_main_reg.data_d[143] ;
 wire \i_main_reg.data_d[144] ;
 wire \i_main_reg.data_d[145] ;
 wire \i_main_reg.data_d[146] ;
 wire \i_main_reg.data_d[147] ;
 wire \i_main_reg.data_d[148] ;
 wire \i_main_reg.data_d[149] ;
 wire \i_main_reg.data_d[14] ;
 wire \i_main_reg.data_d[150] ;
 wire \i_main_reg.data_d[151] ;
 wire \i_main_reg.data_d[152] ;
 wire \i_main_reg.data_d[153] ;
 wire \i_main_reg.data_d[154] ;
 wire \i_main_reg.data_d[155] ;
 wire \i_main_reg.data_d[156] ;
 wire \i_main_reg.data_d[157] ;
 wire \i_main_reg.data_d[158] ;
 wire \i_main_reg.data_d[159] ;
 wire \i_main_reg.data_d[15] ;
 wire \i_main_reg.data_d[160] ;
 wire \i_main_reg.data_d[161] ;
 wire \i_main_reg.data_d[162] ;
 wire \i_main_reg.data_d[163] ;
 wire \i_main_reg.data_d[164] ;
 wire \i_main_reg.data_d[165] ;
 wire \i_main_reg.data_d[166] ;
 wire \i_main_reg.data_d[167] ;
 wire \i_main_reg.data_d[168] ;
 wire \i_main_reg.data_d[169] ;
 wire \i_main_reg.data_d[16] ;
 wire \i_main_reg.data_d[170] ;
 wire \i_main_reg.data_d[171] ;
 wire \i_main_reg.data_d[172] ;
 wire \i_main_reg.data_d[173] ;
 wire \i_main_reg.data_d[174] ;
 wire \i_main_reg.data_d[175] ;
 wire \i_main_reg.data_d[176] ;
 wire \i_main_reg.data_d[177] ;
 wire \i_main_reg.data_d[178] ;
 wire \i_main_reg.data_d[179] ;
 wire \i_main_reg.data_d[17] ;
 wire \i_main_reg.data_d[180] ;
 wire \i_main_reg.data_d[181] ;
 wire \i_main_reg.data_d[182] ;
 wire \i_main_reg.data_d[183] ;
 wire \i_main_reg.data_d[184] ;
 wire \i_main_reg.data_d[185] ;
 wire \i_main_reg.data_d[186] ;
 wire \i_main_reg.data_d[187] ;
 wire \i_main_reg.data_d[188] ;
 wire \i_main_reg.data_d[189] ;
 wire \i_main_reg.data_d[18] ;
 wire \i_main_reg.data_d[190] ;
 wire \i_main_reg.data_d[191] ;
 wire \i_main_reg.data_d[192] ;
 wire \i_main_reg.data_d[193] ;
 wire \i_main_reg.data_d[194] ;
 wire \i_main_reg.data_d[195] ;
 wire \i_main_reg.data_d[196] ;
 wire \i_main_reg.data_d[197] ;
 wire \i_main_reg.data_d[198] ;
 wire \i_main_reg.data_d[199] ;
 wire \i_main_reg.data_d[19] ;
 wire \i_main_reg.data_d[1] ;
 wire \i_main_reg.data_d[200] ;
 wire \i_main_reg.data_d[201] ;
 wire \i_main_reg.data_d[202] ;
 wire \i_main_reg.data_d[203] ;
 wire \i_main_reg.data_d[204] ;
 wire \i_main_reg.data_d[205] ;
 wire \i_main_reg.data_d[206] ;
 wire \i_main_reg.data_d[207] ;
 wire \i_main_reg.data_d[208] ;
 wire \i_main_reg.data_d[209] ;
 wire \i_main_reg.data_d[20] ;
 wire \i_main_reg.data_d[210] ;
 wire \i_main_reg.data_d[211] ;
 wire \i_main_reg.data_d[212] ;
 wire \i_main_reg.data_d[213] ;
 wire \i_main_reg.data_d[214] ;
 wire \i_main_reg.data_d[215] ;
 wire \i_main_reg.data_d[216] ;
 wire \i_main_reg.data_d[217] ;
 wire \i_main_reg.data_d[218] ;
 wire \i_main_reg.data_d[219] ;
 wire \i_main_reg.data_d[21] ;
 wire \i_main_reg.data_d[220] ;
 wire \i_main_reg.data_d[221] ;
 wire \i_main_reg.data_d[222] ;
 wire \i_main_reg.data_d[223] ;
 wire \i_main_reg.data_d[224] ;
 wire \i_main_reg.data_d[225] ;
 wire \i_main_reg.data_d[226] ;
 wire \i_main_reg.data_d[227] ;
 wire \i_main_reg.data_d[228] ;
 wire \i_main_reg.data_d[229] ;
 wire \i_main_reg.data_d[22] ;
 wire \i_main_reg.data_d[230] ;
 wire \i_main_reg.data_d[231] ;
 wire \i_main_reg.data_d[232] ;
 wire \i_main_reg.data_d[233] ;
 wire \i_main_reg.data_d[234] ;
 wire \i_main_reg.data_d[235] ;
 wire \i_main_reg.data_d[236] ;
 wire \i_main_reg.data_d[237] ;
 wire \i_main_reg.data_d[238] ;
 wire \i_main_reg.data_d[239] ;
 wire \i_main_reg.data_d[23] ;
 wire \i_main_reg.data_d[240] ;
 wire \i_main_reg.data_d[241] ;
 wire \i_main_reg.data_d[242] ;
 wire \i_main_reg.data_d[243] ;
 wire \i_main_reg.data_d[244] ;
 wire \i_main_reg.data_d[245] ;
 wire \i_main_reg.data_d[246] ;
 wire \i_main_reg.data_d[247] ;
 wire \i_main_reg.data_d[248] ;
 wire \i_main_reg.data_d[249] ;
 wire \i_main_reg.data_d[24] ;
 wire \i_main_reg.data_d[250] ;
 wire \i_main_reg.data_d[251] ;
 wire \i_main_reg.data_d[252] ;
 wire \i_main_reg.data_d[253] ;
 wire \i_main_reg.data_d[254] ;
 wire \i_main_reg.data_d[255] ;
 wire \i_main_reg.data_d[256] ;
 wire \i_main_reg.data_d[257] ;
 wire \i_main_reg.data_d[258] ;
 wire \i_main_reg.data_d[259] ;
 wire \i_main_reg.data_d[25] ;
 wire \i_main_reg.data_d[260] ;
 wire \i_main_reg.data_d[261] ;
 wire \i_main_reg.data_d[262] ;
 wire \i_main_reg.data_d[263] ;
 wire \i_main_reg.data_d[264] ;
 wire \i_main_reg.data_d[265] ;
 wire \i_main_reg.data_d[266] ;
 wire \i_main_reg.data_d[267] ;
 wire \i_main_reg.data_d[268] ;
 wire \i_main_reg.data_d[269] ;
 wire \i_main_reg.data_d[26] ;
 wire \i_main_reg.data_d[270] ;
 wire \i_main_reg.data_d[271] ;
 wire \i_main_reg.data_d[272] ;
 wire \i_main_reg.data_d[273] ;
 wire \i_main_reg.data_d[274] ;
 wire \i_main_reg.data_d[275] ;
 wire \i_main_reg.data_d[276] ;
 wire \i_main_reg.data_d[277] ;
 wire \i_main_reg.data_d[278] ;
 wire \i_main_reg.data_d[279] ;
 wire \i_main_reg.data_d[27] ;
 wire \i_main_reg.data_d[280] ;
 wire \i_main_reg.data_d[281] ;
 wire \i_main_reg.data_d[282] ;
 wire \i_main_reg.data_d[283] ;
 wire \i_main_reg.data_d[284] ;
 wire \i_main_reg.data_d[285] ;
 wire \i_main_reg.data_d[286] ;
 wire \i_main_reg.data_d[287] ;
 wire \i_main_reg.data_d[288] ;
 wire \i_main_reg.data_d[289] ;
 wire \i_main_reg.data_d[28] ;
 wire \i_main_reg.data_d[290] ;
 wire \i_main_reg.data_d[291] ;
 wire \i_main_reg.data_d[292] ;
 wire \i_main_reg.data_d[293] ;
 wire \i_main_reg.data_d[294] ;
 wire \i_main_reg.data_d[295] ;
 wire \i_main_reg.data_d[296] ;
 wire \i_main_reg.data_d[297] ;
 wire \i_main_reg.data_d[298] ;
 wire \i_main_reg.data_d[299] ;
 wire \i_main_reg.data_d[29] ;
 wire \i_main_reg.data_d[2] ;
 wire \i_main_reg.data_d[300] ;
 wire \i_main_reg.data_d[301] ;
 wire \i_main_reg.data_d[302] ;
 wire \i_main_reg.data_d[303] ;
 wire \i_main_reg.data_d[304] ;
 wire \i_main_reg.data_d[305] ;
 wire \i_main_reg.data_d[306] ;
 wire \i_main_reg.data_d[307] ;
 wire \i_main_reg.data_d[308] ;
 wire \i_main_reg.data_d[309] ;
 wire \i_main_reg.data_d[30] ;
 wire \i_main_reg.data_d[310] ;
 wire \i_main_reg.data_d[311] ;
 wire \i_main_reg.data_d[312] ;
 wire \i_main_reg.data_d[313] ;
 wire \i_main_reg.data_d[314] ;
 wire \i_main_reg.data_d[315] ;
 wire \i_main_reg.data_d[316] ;
 wire \i_main_reg.data_d[317] ;
 wire \i_main_reg.data_d[318] ;
 wire \i_main_reg.data_d[319] ;
 wire \i_main_reg.data_d[31] ;
 wire \i_main_reg.data_d[320] ;
 wire \i_main_reg.data_d[321] ;
 wire \i_main_reg.data_d[322] ;
 wire \i_main_reg.data_d[323] ;
 wire \i_main_reg.data_d[324] ;
 wire \i_main_reg.data_d[325] ;
 wire \i_main_reg.data_d[326] ;
 wire \i_main_reg.data_d[327] ;
 wire \i_main_reg.data_d[328] ;
 wire \i_main_reg.data_d[329] ;
 wire \i_main_reg.data_d[32] ;
 wire \i_main_reg.data_d[330] ;
 wire \i_main_reg.data_d[331] ;
 wire \i_main_reg.data_d[332] ;
 wire \i_main_reg.data_d[333] ;
 wire \i_main_reg.data_d[334] ;
 wire \i_main_reg.data_d[335] ;
 wire \i_main_reg.data_d[336] ;
 wire \i_main_reg.data_d[337] ;
 wire \i_main_reg.data_d[338] ;
 wire \i_main_reg.data_d[339] ;
 wire \i_main_reg.data_d[33] ;
 wire \i_main_reg.data_d[340] ;
 wire \i_main_reg.data_d[341] ;
 wire \i_main_reg.data_d[342] ;
 wire \i_main_reg.data_d[343] ;
 wire \i_main_reg.data_d[344] ;
 wire \i_main_reg.data_d[345] ;
 wire \i_main_reg.data_d[346] ;
 wire \i_main_reg.data_d[347] ;
 wire \i_main_reg.data_d[348] ;
 wire \i_main_reg.data_d[349] ;
 wire \i_main_reg.data_d[34] ;
 wire \i_main_reg.data_d[350] ;
 wire \i_main_reg.data_d[351] ;
 wire \i_main_reg.data_d[352] ;
 wire \i_main_reg.data_d[353] ;
 wire \i_main_reg.data_d[354] ;
 wire \i_main_reg.data_d[355] ;
 wire \i_main_reg.data_d[356] ;
 wire \i_main_reg.data_d[357] ;
 wire \i_main_reg.data_d[358] ;
 wire \i_main_reg.data_d[359] ;
 wire \i_main_reg.data_d[35] ;
 wire \i_main_reg.data_d[360] ;
 wire \i_main_reg.data_d[361] ;
 wire \i_main_reg.data_d[362] ;
 wire \i_main_reg.data_d[363] ;
 wire \i_main_reg.data_d[364] ;
 wire \i_main_reg.data_d[365] ;
 wire \i_main_reg.data_d[366] ;
 wire \i_main_reg.data_d[367] ;
 wire \i_main_reg.data_d[368] ;
 wire \i_main_reg.data_d[369] ;
 wire \i_main_reg.data_d[36] ;
 wire \i_main_reg.data_d[370] ;
 wire \i_main_reg.data_d[371] ;
 wire \i_main_reg.data_d[372] ;
 wire \i_main_reg.data_d[373] ;
 wire \i_main_reg.data_d[374] ;
 wire \i_main_reg.data_d[375] ;
 wire \i_main_reg.data_d[376] ;
 wire \i_main_reg.data_d[377] ;
 wire \i_main_reg.data_d[378] ;
 wire \i_main_reg.data_d[379] ;
 wire \i_main_reg.data_d[37] ;
 wire \i_main_reg.data_d[380] ;
 wire \i_main_reg.data_d[381] ;
 wire \i_main_reg.data_d[382] ;
 wire \i_main_reg.data_d[383] ;
 wire \i_main_reg.data_d[384] ;
 wire \i_main_reg.data_d[385] ;
 wire \i_main_reg.data_d[386] ;
 wire \i_main_reg.data_d[387] ;
 wire \i_main_reg.data_d[388] ;
 wire \i_main_reg.data_d[389] ;
 wire \i_main_reg.data_d[38] ;
 wire \i_main_reg.data_d[390] ;
 wire \i_main_reg.data_d[391] ;
 wire \i_main_reg.data_d[392] ;
 wire \i_main_reg.data_d[393] ;
 wire \i_main_reg.data_d[394] ;
 wire \i_main_reg.data_d[395] ;
 wire \i_main_reg.data_d[396] ;
 wire \i_main_reg.data_d[397] ;
 wire \i_main_reg.data_d[398] ;
 wire \i_main_reg.data_d[399] ;
 wire \i_main_reg.data_d[39] ;
 wire \i_main_reg.data_d[3] ;
 wire \i_main_reg.data_d[400] ;
 wire \i_main_reg.data_d[401] ;
 wire \i_main_reg.data_d[402] ;
 wire \i_main_reg.data_d[403] ;
 wire \i_main_reg.data_d[404] ;
 wire \i_main_reg.data_d[405] ;
 wire \i_main_reg.data_d[406] ;
 wire \i_main_reg.data_d[407] ;
 wire \i_main_reg.data_d[408] ;
 wire \i_main_reg.data_d[409] ;
 wire \i_main_reg.data_d[40] ;
 wire \i_main_reg.data_d[410] ;
 wire \i_main_reg.data_d[411] ;
 wire \i_main_reg.data_d[412] ;
 wire \i_main_reg.data_d[413] ;
 wire \i_main_reg.data_d[414] ;
 wire \i_main_reg.data_d[415] ;
 wire \i_main_reg.data_d[416] ;
 wire \i_main_reg.data_d[417] ;
 wire \i_main_reg.data_d[418] ;
 wire \i_main_reg.data_d[419] ;
 wire \i_main_reg.data_d[41] ;
 wire \i_main_reg.data_d[420] ;
 wire \i_main_reg.data_d[421] ;
 wire \i_main_reg.data_d[422] ;
 wire \i_main_reg.data_d[423] ;
 wire \i_main_reg.data_d[424] ;
 wire \i_main_reg.data_d[425] ;
 wire \i_main_reg.data_d[426] ;
 wire \i_main_reg.data_d[427] ;
 wire \i_main_reg.data_d[428] ;
 wire \i_main_reg.data_d[429] ;
 wire \i_main_reg.data_d[42] ;
 wire \i_main_reg.data_d[430] ;
 wire \i_main_reg.data_d[431] ;
 wire \i_main_reg.data_d[432] ;
 wire \i_main_reg.data_d[433] ;
 wire \i_main_reg.data_d[434] ;
 wire \i_main_reg.data_d[435] ;
 wire \i_main_reg.data_d[436] ;
 wire \i_main_reg.data_d[437] ;
 wire \i_main_reg.data_d[438] ;
 wire \i_main_reg.data_d[439] ;
 wire \i_main_reg.data_d[43] ;
 wire \i_main_reg.data_d[440] ;
 wire \i_main_reg.data_d[441] ;
 wire \i_main_reg.data_d[442] ;
 wire \i_main_reg.data_d[443] ;
 wire \i_main_reg.data_d[444] ;
 wire \i_main_reg.data_d[445] ;
 wire \i_main_reg.data_d[446] ;
 wire \i_main_reg.data_d[44] ;
 wire \i_main_reg.data_d[45] ;
 wire \i_main_reg.data_d[46] ;
 wire \i_main_reg.data_d[47] ;
 wire \i_main_reg.data_d[48] ;
 wire \i_main_reg.data_d[49] ;
 wire \i_main_reg.data_d[4] ;
 wire \i_main_reg.data_d[50] ;
 wire \i_main_reg.data_d[51] ;
 wire \i_main_reg.data_d[52] ;
 wire \i_main_reg.data_d[53] ;
 wire \i_main_reg.data_d[54] ;
 wire \i_main_reg.data_d[55] ;
 wire \i_main_reg.data_d[56] ;
 wire \i_main_reg.data_d[57] ;
 wire \i_main_reg.data_d[58] ;
 wire \i_main_reg.data_d[59] ;
 wire \i_main_reg.data_d[5] ;
 wire \i_main_reg.data_d[60] ;
 wire \i_main_reg.data_d[61] ;
 wire \i_main_reg.data_d[62] ;
 wire \i_main_reg.data_d[63] ;
 wire \i_main_reg.data_d[64] ;
 wire \i_main_reg.data_d[65] ;
 wire \i_main_reg.data_d[66] ;
 wire \i_main_reg.data_d[67] ;
 wire \i_main_reg.data_d[68] ;
 wire \i_main_reg.data_d[69] ;
 wire \i_main_reg.data_d[6] ;
 wire \i_main_reg.data_d[70] ;
 wire \i_main_reg.data_d[71] ;
 wire \i_main_reg.data_d[72] ;
 wire \i_main_reg.data_d[73] ;
 wire \i_main_reg.data_d[74] ;
 wire \i_main_reg.data_d[75] ;
 wire \i_main_reg.data_d[76] ;
 wire \i_main_reg.data_d[77] ;
 wire \i_main_reg.data_d[78] ;
 wire \i_main_reg.data_d[79] ;
 wire \i_main_reg.data_d[7] ;
 wire \i_main_reg.data_d[80] ;
 wire \i_main_reg.data_d[81] ;
 wire \i_main_reg.data_d[82] ;
 wire \i_main_reg.data_d[83] ;
 wire \i_main_reg.data_d[84] ;
 wire \i_main_reg.data_d[85] ;
 wire \i_main_reg.data_d[86] ;
 wire \i_main_reg.data_d[87] ;
 wire \i_main_reg.data_d[88] ;
 wire \i_main_reg.data_d[89] ;
 wire \i_main_reg.data_d[8] ;
 wire \i_main_reg.data_d[90] ;
 wire \i_main_reg.data_d[91] ;
 wire \i_main_reg.data_d[92] ;
 wire \i_main_reg.data_d[93] ;
 wire \i_main_reg.data_d[94] ;
 wire \i_main_reg.data_d[95] ;
 wire \i_main_reg.data_d[96] ;
 wire \i_main_reg.data_d[97] ;
 wire \i_main_reg.data_d[98] ;
 wire \i_main_reg.data_d[99] ;
 wire \i_main_reg.data_d[9] ;
 wire \i_main_reg.data_o ;
 wire \i_step_counter.data_d[0] ;
 wire \i_step_counter.data_d[10] ;
 wire \i_step_counter.data_d[11] ;
 wire \i_step_counter.data_d[12] ;
 wire \i_step_counter.data_d[13] ;
 wire \i_step_counter.data_d[14] ;
 wire \i_step_counter.data_d[1] ;
 wire \i_step_counter.data_d[2] ;
 wire \i_step_counter.data_d[3] ;
 wire \i_step_counter.data_d[4] ;
 wire \i_step_counter.data_d[5] ;
 wire \i_step_counter.data_d[6] ;
 wire \i_step_counter.data_d[7] ;
 wire \i_step_counter.data_d[8] ;
 wire \i_step_counter.data_d[9] ;
 wire \i_step_counter.data_o ;
 wire \one_count_q[0] ;
 wire \one_count_q[1] ;
 wire overflow_q;
 wire previous_bit_q;
 wire \state_q[0] ;
 wire \state_q[1] ;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire clknet_leaf_0_clk;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;

 sg13g2_inv_2 _0628_ (.Y(_0597_),
    .A(net870));
 sg13g2_inv_1 _0629_ (.Y(_0598_),
    .A(net669));
 sg13g2_inv_1 _0630_ (.Y(_0599_),
    .A(net345));
 sg13g2_inv_1 _0631_ (.Y(_0600_),
    .A(net58));
 sg13g2_inv_1 _0632_ (.Y(_0601_),
    .A(net41));
 sg13g2_inv_1 _0633_ (.Y(_0602_),
    .A(net793));
 sg13g2_inv_1 _0634_ (.Y(_0603_),
    .A(net43));
 sg13g2_inv_1 _0635_ (.Y(_0604_),
    .A(net858));
 sg13g2_inv_2 _0636_ (.Y(_0605_),
    .A(net805));
 sg13g2_inv_1 _0637_ (.Y(_0606_),
    .A(net27));
 sg13g2_nor2_1 _0638_ (.A(net437),
    .B(\state_q[0] ),
    .Y(_0607_));
 sg13g2_and2_1 _0639_ (.A(net3),
    .B(_0607_),
    .X(_0608_));
 sg13g2_nand2_1 _0640_ (.Y(_0609_),
    .A(\bit_counter_q[8] ),
    .B(\bit_counter_q[7] ));
 sg13g2_and3_2 _0641_ (.X(_0610_),
    .A(\bit_counter_q[8] ),
    .B(\bit_counter_q[7] ),
    .C(\bit_counter_q[6] ));
 sg13g2_nand3_1 _0642_ (.B(\bit_counter_q[7] ),
    .C(\bit_counter_q[6] ),
    .A(\bit_counter_q[8] ),
    .Y(_0611_));
 sg13g2_nor2_2 _0643_ (.A(net669),
    .B(_0610_),
    .Y(_0612_));
 sg13g2_nor2b_2 _0644_ (.A(net870),
    .B_N(net437),
    .Y(_0613_));
 sg13g2_nand2b_2 _0645_ (.Y(_0614_),
    .B(net436),
    .A_N(\state_q[0] ));
 sg13g2_nand2_1 _0646_ (.Y(_0615_),
    .A(_0612_),
    .B(_0613_));
 sg13g2_nand2b_1 _0647_ (.Y(_0616_),
    .B(net33),
    .A_N(net435));
 sg13g2_nor2_1 _0648_ (.A(net345),
    .B(net33),
    .Y(_0617_));
 sg13g2_nand2_1 _0649_ (.Y(_0618_),
    .A(_0599_),
    .B(_0616_));
 sg13g2_a221oi_1 _0650_ (.B2(_0599_),
    .C1(_0614_),
    .B1(_0616_),
    .A1(_0598_),
    .Y(_0619_),
    .A2(_0611_));
 sg13g2_nand3b_1 _0651_ (.B(_0613_),
    .C(_0618_),
    .Y(_0620_),
    .A_N(_0612_));
 sg13g2_nor3_2 _0652_ (.A(net437),
    .B(\state_q[0] ),
    .C(net4),
    .Y(_0621_));
 sg13g2_nor2_1 _0653_ (.A(net436),
    .B(_0597_),
    .Y(_0622_));
 sg13g2_and2_1 _0654_ (.A(_0612_),
    .B(_0622_),
    .X(_0623_));
 sg13g2_nand2_1 _0655_ (.Y(_0624_),
    .A(_0612_),
    .B(_0622_));
 sg13g2_xnor2_1 _0656_ (.Y(_0625_),
    .A(net436),
    .B(\state_q[0] ));
 sg13g2_nand2b_2 _0657_ (.Y(_0626_),
    .B(_0612_),
    .A_N(_0625_));
 sg13g2_nor3_2 _0658_ (.A(net669),
    .B(_0610_),
    .C(_0625_),
    .Y(_0627_));
 sg13g2_nor2_1 _0659_ (.A(_0621_),
    .B(_0623_),
    .Y(_0482_));
 sg13g2_nor4_2 _0660_ (.A(\state_q[0] ),
    .B(_0619_),
    .C(_0621_),
    .Y(_0483_),
    .D(_0627_));
 sg13g2_a21o_1 _0661_ (.A2(\state_q[0] ),
    .A1(net436),
    .B1(_0621_),
    .X(_0484_));
 sg13g2_a21oi_2 _0662_ (.B1(_0484_),
    .Y(_0485_),
    .A2(_0483_),
    .A1(net436));
 sg13g2_a221oi_1 _0663_ (.B2(net436),
    .C1(_0484_),
    .B1(_0483_),
    .A1(_0612_),
    .Y(_0486_),
    .A2(_0613_));
 sg13g2_a21oi_2 _0664_ (.B1(net434),
    .Y(_0487_),
    .A2(_0486_),
    .A1(_0597_));
 sg13g2_a21o_2 _0665_ (.A2(_0486_),
    .A1(_0597_),
    .B1(net434),
    .X(_0488_));
 sg13g2_a22oi_1 _0666_ (.Y(_0489_),
    .B1(_0487_),
    .B2(net670),
    .A2(_0608_),
    .A1(\i_step_counter.data_d[0] ));
 sg13g2_o21ai_1 _0667_ (.B1(_0489_),
    .Y(_0000_),
    .A1(net670),
    .A2(_0620_));
 sg13g2_xor2_1 _0668_ (.B(net670),
    .A(net877),
    .X(_0490_));
 sg13g2_nand3_1 _0669_ (.B(net352),
    .C(_0490_),
    .A(_0613_),
    .Y(_0491_));
 sg13g2_a22oi_1 _0670_ (.Y(_0492_),
    .B1(_0487_),
    .B2(net877),
    .A2(net434),
    .A1(net864));
 sg13g2_nand2_1 _0671_ (.Y(_0001_),
    .A(_0491_),
    .B(_0492_));
 sg13g2_nand3_1 _0672_ (.B(net670),
    .C(net864),
    .A(\i_step_counter.data_d[0] ),
    .Y(_0493_));
 sg13g2_a21o_1 _0673_ (.A2(net670),
    .A1(\i_step_counter.data_d[0] ),
    .B1(net864),
    .X(_0494_));
 sg13g2_nand2_1 _0674_ (.Y(_0495_),
    .A(_0493_),
    .B(_0494_));
 sg13g2_a22oi_1 _0675_ (.Y(_0496_),
    .B1(net353),
    .B2(net864),
    .A2(net434),
    .A1(\i_step_counter.data_d[2] ));
 sg13g2_o21ai_1 _0676_ (.B1(net865),
    .Y(_0002_),
    .A1(_0620_),
    .A2(_0495_));
 sg13g2_and4_1 _0677_ (.A(\i_step_counter.data_d[0] ),
    .B(\i_step_counter.data_o ),
    .C(\i_step_counter.data_d[1] ),
    .D(\i_step_counter.data_d[2] ),
    .X(_0497_));
 sg13g2_xor2_1 _0678_ (.B(_0493_),
    .A(net871),
    .X(_0498_));
 sg13g2_a22oi_1 _0679_ (.Y(_0499_),
    .B1(_0487_),
    .B2(net871),
    .A2(_0608_),
    .A1(\i_step_counter.data_d[3] ));
 sg13g2_o21ai_1 _0680_ (.B1(net872),
    .Y(_0003_),
    .A1(_0620_),
    .A2(_0498_));
 sg13g2_nand2_1 _0681_ (.Y(_0500_),
    .A(net58),
    .B(net433));
 sg13g2_nand2_1 _0682_ (.Y(_0501_),
    .A(\i_step_counter.data_d[3] ),
    .B(_0497_));
 sg13g2_a21oi_1 _0683_ (.A1(_0613_),
    .A2(_0501_),
    .Y(_0502_),
    .B1(net353));
 sg13g2_a21oi_1 _0684_ (.A1(net352),
    .A2(_0497_),
    .Y(_0503_),
    .B1(\i_step_counter.data_d[3] ));
 sg13g2_o21ai_1 _0685_ (.B1(_0500_),
    .Y(_0004_),
    .A1(_0502_),
    .A2(_0503_));
 sg13g2_nor2_1 _0686_ (.A(net58),
    .B(_0501_),
    .Y(_0504_));
 sg13g2_a22oi_1 _0687_ (.Y(_0505_),
    .B1(_0619_),
    .B2(_0504_),
    .A2(net433),
    .A1(net874));
 sg13g2_o21ai_1 _0688_ (.B1(net875),
    .Y(_0005_),
    .A1(_0600_),
    .A2(_0502_));
 sg13g2_nand2_1 _0689_ (.Y(_0506_),
    .A(net41),
    .B(net433));
 sg13g2_and2_1 _0690_ (.A(\i_step_counter.data_d[3] ),
    .B(\i_step_counter.data_d[4] ),
    .X(_0507_));
 sg13g2_nor2_1 _0691_ (.A(_0600_),
    .B(_0501_),
    .Y(_0508_));
 sg13g2_nand2_1 _0692_ (.Y(_0509_),
    .A(\i_step_counter.data_d[5] ),
    .B(_0508_));
 sg13g2_a21oi_1 _0693_ (.A1(_0613_),
    .A2(_0509_),
    .Y(_0510_),
    .B1(net353));
 sg13g2_a21oi_1 _0694_ (.A1(net352),
    .A2(_0508_),
    .Y(_0511_),
    .B1(\i_step_counter.data_d[5] ));
 sg13g2_o21ai_1 _0695_ (.B1(_0506_),
    .Y(_0006_),
    .A1(_0510_),
    .A2(_0511_));
 sg13g2_nor2_1 _0696_ (.A(net41),
    .B(_0509_),
    .Y(_0512_));
 sg13g2_a22oi_1 _0697_ (.Y(_0513_),
    .B1(_0619_),
    .B2(_0512_),
    .A2(net433),
    .A1(net833));
 sg13g2_o21ai_1 _0698_ (.B1(net834),
    .Y(_0007_),
    .A1(_0601_),
    .A2(_0510_));
 sg13g2_nand2_1 _0699_ (.Y(_0514_),
    .A(net793),
    .B(net433));
 sg13g2_and3_1 _0700_ (.X(_0515_),
    .A(\i_step_counter.data_d[5] ),
    .B(net41),
    .C(_0508_));
 sg13g2_nand4_1 _0701_ (.B(net41),
    .C(_0497_),
    .A(\i_step_counter.data_d[5] ),
    .Y(_0516_),
    .D(_0507_));
 sg13g2_a21oi_1 _0702_ (.A1(net833),
    .A2(_0515_),
    .Y(_0517_),
    .B1(_0614_));
 sg13g2_nor2_1 _0703_ (.A(net353),
    .B(_0517_),
    .Y(_0518_));
 sg13g2_a21oi_1 _0704_ (.A1(net352),
    .A2(_0515_),
    .Y(_0519_),
    .B1(\i_step_counter.data_d[7] ));
 sg13g2_o21ai_1 _0705_ (.B1(_0514_),
    .Y(_0008_),
    .A1(_0518_),
    .A2(_0519_));
 sg13g2_o21ai_1 _0706_ (.B1(net793),
    .Y(_0520_),
    .A1(net353),
    .A2(_0517_));
 sg13g2_nand2_1 _0707_ (.Y(_0521_),
    .A(net867),
    .B(net433));
 sg13g2_nand4_1 _0708_ (.B(_0602_),
    .C(_0619_),
    .A(net833),
    .Y(_0522_),
    .D(_0515_));
 sg13g2_nand3_1 _0709_ (.B(_0521_),
    .C(_0522_),
    .A(_0520_),
    .Y(_0009_));
 sg13g2_nand2_1 _0710_ (.Y(_0523_),
    .A(net43),
    .B(net433));
 sg13g2_nand2_1 _0711_ (.Y(_0524_),
    .A(net833),
    .B(net793));
 sg13g2_nor2_1 _0712_ (.A(_0516_),
    .B(_0524_),
    .Y(_0525_));
 sg13g2_a21oi_1 _0713_ (.A1(\i_step_counter.data_d[9] ),
    .A2(_0525_),
    .Y(_0526_),
    .B1(_0614_));
 sg13g2_nor2_1 _0714_ (.A(net353),
    .B(_0526_),
    .Y(_0527_));
 sg13g2_a21oi_1 _0715_ (.A1(net352),
    .A2(_0525_),
    .Y(_0528_),
    .B1(\i_step_counter.data_d[9] ));
 sg13g2_o21ai_1 _0716_ (.B1(_0523_),
    .Y(_0010_),
    .A1(_0527_),
    .A2(_0528_));
 sg13g2_and4_1 _0717_ (.A(\i_step_counter.data_d[9] ),
    .B(_0603_),
    .C(_0619_),
    .D(_0525_),
    .X(_0529_));
 sg13g2_a21oi_1 _0718_ (.A1(net858),
    .A2(net433),
    .Y(_0530_),
    .B1(_0529_));
 sg13g2_o21ai_1 _0719_ (.B1(net859),
    .Y(_0011_),
    .A1(_0603_),
    .A2(_0527_));
 sg13g2_nand2_1 _0720_ (.Y(_0531_),
    .A(net854),
    .B(net434));
 sg13g2_nand2_1 _0721_ (.Y(_0532_),
    .A(\i_step_counter.data_d[9] ),
    .B(net43));
 sg13g2_nor3_1 _0722_ (.A(_0516_),
    .B(_0524_),
    .C(_0532_),
    .Y(_0533_));
 sg13g2_nor4_1 _0723_ (.A(_0604_),
    .B(_0516_),
    .C(_0524_),
    .D(_0532_),
    .Y(_0534_));
 sg13g2_nor2_1 _0724_ (.A(_0614_),
    .B(_0534_),
    .Y(_0535_));
 sg13g2_nor2_1 _0725_ (.A(net353),
    .B(_0535_),
    .Y(_0536_));
 sg13g2_a21oi_1 _0726_ (.A1(net352),
    .A2(_0533_),
    .Y(_0537_),
    .B1(\i_step_counter.data_d[11] ));
 sg13g2_o21ai_1 _0727_ (.B1(_0531_),
    .Y(_0012_),
    .A1(_0536_),
    .A2(_0537_));
 sg13g2_o21ai_1 _0728_ (.B1(net854),
    .Y(_0538_),
    .A1(net353),
    .A2(_0535_));
 sg13g2_nand2_1 _0729_ (.Y(_0539_),
    .A(net862),
    .B(net434));
 sg13g2_nand3b_1 _0730_ (.B(_0619_),
    .C(_0534_),
    .Y(_0540_),
    .A_N(net854));
 sg13g2_nand3_1 _0731_ (.B(_0539_),
    .C(_0540_),
    .A(_0538_),
    .Y(_0013_));
 sg13g2_nand2_1 _0732_ (.Y(_0541_),
    .A(net805),
    .B(net434));
 sg13g2_and2_1 _0733_ (.A(\i_step_counter.data_d[12] ),
    .B(_0534_),
    .X(_0542_));
 sg13g2_nand3_1 _0734_ (.B(net862),
    .C(_0534_),
    .A(net854),
    .Y(_0543_));
 sg13g2_nand2_1 _0735_ (.Y(_0544_),
    .A(_0613_),
    .B(_0543_));
 sg13g2_and2_1 _0736_ (.A(net352),
    .B(_0544_),
    .X(_0545_));
 sg13g2_a21oi_1 _0737_ (.A1(net352),
    .A2(_0542_),
    .Y(_0546_),
    .B1(\i_step_counter.data_d[13] ));
 sg13g2_o21ai_1 _0738_ (.B1(_0541_),
    .Y(_0014_),
    .A1(_0545_),
    .A2(_0546_));
 sg13g2_o21ai_1 _0739_ (.B1(_0619_),
    .Y(_0547_),
    .A1(_0605_),
    .A2(_0543_));
 sg13g2_a21o_1 _0740_ (.A2(_0543_),
    .A1(_0605_),
    .B1(_0547_),
    .X(_0548_));
 sg13g2_o21ai_1 _0741_ (.B1(_0548_),
    .Y(_0015_),
    .A1(_0605_),
    .A2(_0488_));
 sg13g2_mux2_1 _0742_ (.A0(net98),
    .A1(net437),
    .S(_0483_),
    .X(_0016_));
 sg13g2_and2_1 _0743_ (.A(net25),
    .B(net29),
    .X(_0549_));
 sg13g2_and4_1 _0744_ (.A(net31),
    .B(\bit_counter_q[3] ),
    .C(net753),
    .D(_0549_),
    .X(_0550_));
 sg13g2_and2_1 _0745_ (.A(\bit_counter_q[5] ),
    .B(_0550_),
    .X(_0551_));
 sg13g2_a21o_1 _0746_ (.A2(net824),
    .A1(net435),
    .B1(previous_bit_q),
    .X(_0552_));
 sg13g2_o21ai_1 _0747_ (.B1(_0552_),
    .Y(_0553_),
    .A1(net435),
    .A2(net824));
 sg13g2_nor4_1 _0748_ (.A(\bit_counter_q[9] ),
    .B(\bit_counter_q[6] ),
    .C(_0609_),
    .D(_0553_),
    .Y(_0554_));
 sg13g2_nand2_1 _0749_ (.Y(_0555_),
    .A(_0551_),
    .B(_0554_));
 sg13g2_a22oi_1 _0750_ (.Y(_0556_),
    .B1(_0622_),
    .B2(_0555_),
    .A2(_0613_),
    .A1(_0605_));
 sg13g2_nand3_1 _0751_ (.B(_0544_),
    .C(_0556_),
    .A(_0486_),
    .Y(_0557_));
 sg13g2_a22oi_1 _0752_ (.Y(_0017_),
    .B1(_0557_),
    .B2(_0606_),
    .A2(_0607_),
    .A1(net4));
 sg13g2_nor2_1 _0753_ (.A(net435),
    .B(_0614_),
    .Y(_0558_));
 sg13g2_nor3_1 _0754_ (.A(net435),
    .B(_0614_),
    .C(_0617_),
    .Y(_0559_));
 sg13g2_nand2b_1 _0755_ (.Y(_0560_),
    .B(_0558_),
    .A_N(_0617_));
 sg13g2_a221oi_1 _0756_ (.B2(_0614_),
    .C1(_0559_),
    .B1(_0624_),
    .A1(_0597_),
    .Y(_0030_),
    .A2(_0620_));
 sg13g2_nor2_1 _0757_ (.A(net824),
    .B(_0030_),
    .Y(_0561_));
 sg13g2_a21oi_1 _0758_ (.A1(_0623_),
    .A2(_0553_),
    .Y(_0018_),
    .B1(_0561_));
 sg13g2_nor2b_1 _0759_ (.A(_0030_),
    .B_N(net879),
    .Y(_0562_));
 sg13g2_a21o_1 _0760_ (.A2(_0623_),
    .A1(net435),
    .B1(_0562_),
    .X(_0019_));
 sg13g2_nor2_1 _0761_ (.A(net29),
    .B(_0627_),
    .Y(_0563_));
 sg13g2_a21oi_1 _0762_ (.A1(net29),
    .A2(net354),
    .Y(_0020_),
    .B1(_0563_));
 sg13g2_a21oi_1 _0763_ (.A1(\bit_counter_q[0] ),
    .A2(net354),
    .Y(_0564_),
    .B1(net25));
 sg13g2_o21ai_1 _0764_ (.B1(net354),
    .Y(_0565_),
    .A1(_0626_),
    .A2(_0549_));
 sg13g2_nor2b_1 _0765_ (.A(net26),
    .B_N(_0565_),
    .Y(_0021_));
 sg13g2_nand2_1 _0766_ (.Y(_0566_),
    .A(_0627_),
    .B(_0549_));
 sg13g2_nand2_1 _0767_ (.Y(_0567_),
    .A(net31),
    .B(_0565_));
 sg13g2_o21ai_1 _0768_ (.B1(_0567_),
    .Y(_0022_),
    .A1(net31),
    .A2(_0566_));
 sg13g2_nand3_1 _0769_ (.B(_0485_),
    .C(_0549_),
    .A(net31),
    .Y(_0568_));
 sg13g2_and4_1 _0770_ (.A(net31),
    .B(\bit_counter_q[3] ),
    .C(_0485_),
    .D(_0549_),
    .X(_0569_));
 sg13g2_xor2_1 _0771_ (.B(_0568_),
    .A(net861),
    .X(_0570_));
 sg13g2_a21oi_1 _0772_ (.A1(_0626_),
    .A2(net354),
    .Y(_0023_),
    .B1(_0570_));
 sg13g2_o21ai_1 _0773_ (.B1(_0485_),
    .Y(_0571_),
    .A1(_0626_),
    .A2(_0550_));
 sg13g2_o21ai_1 _0774_ (.B1(_0571_),
    .Y(_0572_),
    .A1(net753),
    .A2(_0569_));
 sg13g2_inv_1 _0775_ (.Y(_0024_),
    .A(net754));
 sg13g2_and2_1 _0776_ (.A(_0627_),
    .B(_0550_),
    .X(_0573_));
 sg13g2_mux2_1 _0777_ (.A0(_0573_),
    .A1(_0571_),
    .S(net850),
    .X(_0025_));
 sg13g2_a21oi_1 _0778_ (.A1(net354),
    .A2(_0551_),
    .Y(_0574_),
    .B1(net39));
 sg13g2_and2_1 _0779_ (.A(net39),
    .B(_0551_),
    .X(_0575_));
 sg13g2_o21ai_1 _0780_ (.B1(net354),
    .Y(_0576_),
    .A1(_0626_),
    .A2(_0575_));
 sg13g2_nor2b_1 _0781_ (.A(net40),
    .B_N(_0576_),
    .Y(_0026_));
 sg13g2_and2_1 _0782_ (.A(_0627_),
    .B(_0575_),
    .X(_0577_));
 sg13g2_mux2_1 _0783_ (.A0(_0577_),
    .A1(_0576_),
    .S(net869),
    .X(_0027_));
 sg13g2_a21oi_1 _0784_ (.A1(\bit_counter_q[7] ),
    .A2(_0577_),
    .Y(_0578_),
    .B1(net47));
 sg13g2_a21oi_1 _0785_ (.A1(_0626_),
    .A2(net354),
    .Y(_0028_),
    .B1(net48));
 sg13g2_nor2_1 _0786_ (.A(_0598_),
    .B(net354),
    .Y(_0029_));
 sg13g2_nand3_1 _0787_ (.B(_0626_),
    .C(_0560_),
    .A(net436),
    .Y(_0579_));
 sg13g2_and2_1 _0788_ (.A(_0482_),
    .B(_0579_),
    .X(_0031_));
 sg13g2_nor2_1 _0789_ (.A(net2),
    .B(_0627_),
    .Y(_0580_));
 sg13g2_nor3_2 _0790_ (.A(net2),
    .B(_0627_),
    .C(_0559_),
    .Y(_0581_));
 sg13g2_nand2_1 _0791_ (.Y(_0582_),
    .A(_0560_),
    .B(_0580_));
 sg13g2_a22oi_1 _0792_ (.Y(_0583_),
    .B1(_0582_),
    .B2(net37),
    .A2(_0580_),
    .A1(\i_main_reg.data_o ));
 sg13g2_inv_1 _0793_ (.Y(_0032_),
    .A(net38));
 sg13g2_mux2_1 _0794_ (.A0(net88),
    .A1(net37),
    .S(net431),
    .X(_0033_));
 sg13g2_mux2_1 _0795_ (.A0(\i_main_reg.data_d[2] ),
    .A1(net88),
    .S(net429),
    .X(_0034_));
 sg13g2_mux2_1 _0796_ (.A0(net596),
    .A1(net702),
    .S(net430),
    .X(_0035_));
 sg13g2_mux2_1 _0797_ (.A0(\i_main_reg.data_d[4] ),
    .A1(net596),
    .S(net430),
    .X(_0036_));
 sg13g2_mux2_1 _0798_ (.A0(\i_main_reg.data_d[5] ),
    .A1(net708),
    .S(net429),
    .X(_0037_));
 sg13g2_mux2_1 _0799_ (.A0(net274),
    .A1(\i_main_reg.data_d[5] ),
    .S(net429),
    .X(_0038_));
 sg13g2_mux2_1 _0800_ (.A0(net602),
    .A1(net274),
    .S(net429),
    .X(_0039_));
 sg13g2_mux2_1 _0801_ (.A0(net737),
    .A1(net602),
    .S(net415),
    .X(_0040_));
 sg13g2_mux2_1 _0802_ (.A0(net755),
    .A1(net737),
    .S(net415),
    .X(_0041_));
 sg13g2_mux2_1 _0803_ (.A0(net569),
    .A1(\i_main_reg.data_d[9] ),
    .S(net415),
    .X(_0042_));
 sg13g2_mux2_1 _0804_ (.A0(net304),
    .A1(net569),
    .S(net414),
    .X(_0043_));
 sg13g2_mux2_1 _0805_ (.A0(\i_main_reg.data_d[12] ),
    .A1(net304),
    .S(net414),
    .X(_0044_));
 sg13g2_mux2_1 _0806_ (.A0(net103),
    .A1(\i_main_reg.data_d[12] ),
    .S(net414),
    .X(_0045_));
 sg13g2_mux2_1 _0807_ (.A0(net80),
    .A1(net103),
    .S(net414),
    .X(_0046_));
 sg13g2_mux2_1 _0808_ (.A0(\i_main_reg.data_d[15] ),
    .A1(net80),
    .S(net410),
    .X(_0047_));
 sg13g2_mux2_1 _0809_ (.A0(\i_main_reg.data_d[16] ),
    .A1(net175),
    .S(net410),
    .X(_0048_));
 sg13g2_mux2_1 _0810_ (.A0(\i_main_reg.data_d[17] ),
    .A1(net676),
    .S(net410),
    .X(_0049_));
 sg13g2_mux2_1 _0811_ (.A0(net545),
    .A1(\i_main_reg.data_d[17] ),
    .S(net409),
    .X(_0050_));
 sg13g2_mux2_1 _0812_ (.A0(net184),
    .A1(net545),
    .S(net409),
    .X(_0051_));
 sg13g2_mux2_1 _0813_ (.A0(\i_main_reg.data_d[20] ),
    .A1(net184),
    .S(net410),
    .X(_0052_));
 sg13g2_mux2_1 _0814_ (.A0(net230),
    .A1(\i_main_reg.data_d[20] ),
    .S(net409),
    .X(_0053_));
 sg13g2_mux2_1 _0815_ (.A0(net549),
    .A1(net230),
    .S(net409),
    .X(_0054_));
 sg13g2_mux2_1 _0816_ (.A0(net265),
    .A1(net549),
    .S(net409),
    .X(_0055_));
 sg13g2_mux2_1 _0817_ (.A0(\i_main_reg.data_d[24] ),
    .A1(net265),
    .S(net409),
    .X(_0056_));
 sg13g2_mux2_1 _0818_ (.A0(\i_main_reg.data_d[25] ),
    .A1(net652),
    .S(net409),
    .X(_0057_));
 sg13g2_mux2_1 _0819_ (.A0(net553),
    .A1(net654),
    .S(net409),
    .X(_0058_));
 sg13g2_mux2_1 _0820_ (.A0(net216),
    .A1(net553),
    .S(net411),
    .X(_0059_));
 sg13g2_mux2_1 _0821_ (.A0(\i_main_reg.data_d[28] ),
    .A1(net216),
    .S(net411),
    .X(_0060_));
 sg13g2_mux2_1 _0822_ (.A0(net234),
    .A1(net254),
    .S(net408),
    .X(_0061_));
 sg13g2_mux2_1 _0823_ (.A0(\i_main_reg.data_d[30] ),
    .A1(net234),
    .S(net412),
    .X(_0062_));
 sg13g2_mux2_1 _0824_ (.A0(\i_main_reg.data_d[31] ),
    .A1(net564),
    .S(net412),
    .X(_0063_));
 sg13g2_mux2_1 _0825_ (.A0(net575),
    .A1(\i_main_reg.data_d[31] ),
    .S(net412),
    .X(_0064_));
 sg13g2_mux2_1 _0826_ (.A0(net149),
    .A1(\i_main_reg.data_d[32] ),
    .S(net413),
    .X(_0065_));
 sg13g2_mux2_1 _0827_ (.A0(net703),
    .A1(net149),
    .S(net413),
    .X(_0066_));
 sg13g2_mux2_1 _0828_ (.A0(net715),
    .A1(net703),
    .S(net413),
    .X(_0067_));
 sg13g2_mux2_1 _0829_ (.A0(net828),
    .A1(net715),
    .S(net413),
    .X(_0068_));
 sg13g2_mux2_1 _0830_ (.A0(\i_main_reg.data_d[37] ),
    .A1(net828),
    .S(net413),
    .X(_0069_));
 sg13g2_mux2_1 _0831_ (.A0(net581),
    .A1(\i_main_reg.data_d[37] ),
    .S(net412),
    .X(_0070_));
 sg13g2_mux2_1 _0832_ (.A0(net123),
    .A1(\i_main_reg.data_d[38] ),
    .S(net412),
    .X(_0071_));
 sg13g2_mux2_1 _0833_ (.A0(net215),
    .A1(net123),
    .S(net412),
    .X(_0072_));
 sg13g2_mux2_1 _0834_ (.A0(net804),
    .A1(net215),
    .S(net430),
    .X(_0073_));
 sg13g2_mux2_1 _0835_ (.A0(net812),
    .A1(net804),
    .S(net430),
    .X(_0074_));
 sg13g2_mux2_1 _0836_ (.A0(net155),
    .A1(\i_main_reg.data_d[42] ),
    .S(net420),
    .X(_0075_));
 sg13g2_mux2_1 _0837_ (.A0(net218),
    .A1(net155),
    .S(net420),
    .X(_0076_));
 sg13g2_mux2_1 _0838_ (.A0(net552),
    .A1(net218),
    .S(net420),
    .X(_0077_));
 sg13g2_mux2_1 _0839_ (.A0(net779),
    .A1(net552),
    .S(net420),
    .X(_0078_));
 sg13g2_mux2_1 _0840_ (.A0(net293),
    .A1(\i_main_reg.data_d[46] ),
    .S(net421),
    .X(_0079_));
 sg13g2_mux2_1 _0841_ (.A0(net342),
    .A1(net293),
    .S(net420),
    .X(_0080_));
 sg13g2_mux2_1 _0842_ (.A0(net598),
    .A1(net342),
    .S(net427),
    .X(_0081_));
 sg13g2_mux2_1 _0843_ (.A0(\i_main_reg.data_d[50] ),
    .A1(net598),
    .S(net425),
    .X(_0082_));
 sg13g2_mux2_1 _0844_ (.A0(net642),
    .A1(net647),
    .S(net425),
    .X(_0083_));
 sg13g2_mux2_1 _0845_ (.A0(\i_main_reg.data_d[52] ),
    .A1(net642),
    .S(net426),
    .X(_0084_));
 sg13g2_mux2_1 _0846_ (.A0(net310),
    .A1(\i_main_reg.data_d[52] ),
    .S(net427),
    .X(_0085_));
 sg13g2_mux2_1 _0847_ (.A0(net520),
    .A1(net310),
    .S(net426),
    .X(_0086_));
 sg13g2_mux2_1 _0848_ (.A0(net146),
    .A1(net520),
    .S(net427),
    .X(_0087_));
 sg13g2_mux2_1 _0849_ (.A0(net84),
    .A1(net146),
    .S(net426),
    .X(_0088_));
 sg13g2_mux2_1 _0850_ (.A0(\i_main_reg.data_d[57] ),
    .A1(net84),
    .S(net427),
    .X(_0089_));
 sg13g2_mux2_1 _0851_ (.A0(net621),
    .A1(net678),
    .S(net426),
    .X(_0090_));
 sg13g2_mux2_1 _0852_ (.A0(\i_main_reg.data_d[59] ),
    .A1(net621),
    .S(net426),
    .X(_0091_));
 sg13g2_mux2_1 _0853_ (.A0(net268),
    .A1(\i_main_reg.data_d[59] ),
    .S(net425),
    .X(_0092_));
 sg13g2_mux2_1 _0854_ (.A0(net716),
    .A1(net268),
    .S(net425),
    .X(_0093_));
 sg13g2_mux2_1 _0855_ (.A0(net725),
    .A1(net716),
    .S(net425),
    .X(_0094_));
 sg13g2_mux2_1 _0856_ (.A0(net732),
    .A1(net725),
    .S(net421),
    .X(_0095_));
 sg13g2_mux2_1 _0857_ (.A0(net762),
    .A1(net732),
    .S(net421),
    .X(_0096_));
 sg13g2_mux2_1 _0858_ (.A0(net704),
    .A1(net762),
    .S(net421),
    .X(_0097_));
 sg13g2_mux2_1 _0859_ (.A0(net686),
    .A1(net704),
    .S(net419),
    .X(_0098_));
 sg13g2_mux2_1 _0860_ (.A0(\i_main_reg.data_d[67] ),
    .A1(net686),
    .S(net418),
    .X(_0099_));
 sg13g2_mux2_1 _0861_ (.A0(net839),
    .A1(\i_main_reg.data_d[67] ),
    .S(net418),
    .X(_0100_));
 sg13g2_mux2_1 _0862_ (.A0(net830),
    .A1(\i_main_reg.data_d[68] ),
    .S(net418),
    .X(_0101_));
 sg13g2_mux2_1 _0863_ (.A0(net843),
    .A1(net830),
    .S(net418),
    .X(_0102_));
 sg13g2_mux2_1 _0864_ (.A0(net785),
    .A1(net843),
    .S(net419),
    .X(_0103_));
 sg13g2_mux2_1 _0865_ (.A0(\i_main_reg.data_d[72] ),
    .A1(net785),
    .S(net419),
    .X(_0104_));
 sg13g2_mux2_1 _0866_ (.A0(net674),
    .A1(\i_main_reg.data_d[72] ),
    .S(net419),
    .X(_0105_));
 sg13g2_mux2_1 _0867_ (.A0(net86),
    .A1(\i_main_reg.data_d[73] ),
    .S(net417),
    .X(_0106_));
 sg13g2_mux2_1 _0868_ (.A0(net561),
    .A1(net86),
    .S(net417),
    .X(_0107_));
 sg13g2_mux2_1 _0869_ (.A0(net333),
    .A1(\i_main_reg.data_d[75] ),
    .S(net417),
    .X(_0108_));
 sg13g2_mux2_1 _0870_ (.A0(net600),
    .A1(net333),
    .S(net417),
    .X(_0109_));
 sg13g2_mux2_1 _0871_ (.A0(net347),
    .A1(\i_main_reg.data_d[77] ),
    .S(net417),
    .X(_0110_));
 sg13g2_mux2_1 _0872_ (.A0(net658),
    .A1(net347),
    .S(net417),
    .X(_0111_));
 sg13g2_mux2_1 _0873_ (.A0(net672),
    .A1(net658),
    .S(net417),
    .X(_0112_));
 sg13g2_mux2_1 _0874_ (.A0(net733),
    .A1(net672),
    .S(net417),
    .X(_0113_));
 sg13g2_mux2_1 _0875_ (.A0(\i_main_reg.data_d[82] ),
    .A1(net733),
    .S(net418),
    .X(_0114_));
 sg13g2_mux2_1 _0876_ (.A0(net728),
    .A1(net846),
    .S(net418),
    .X(_0115_));
 sg13g2_mux2_1 _0877_ (.A0(net705),
    .A1(net728),
    .S(net418),
    .X(_0116_));
 sg13g2_mux2_1 _0878_ (.A0(net662),
    .A1(net705),
    .S(net418),
    .X(_0117_));
 sg13g2_mux2_1 _0879_ (.A0(\i_main_reg.data_d[86] ),
    .A1(net662),
    .S(net424),
    .X(_0118_));
 sg13g2_mux2_1 _0880_ (.A0(\i_main_reg.data_d[87] ),
    .A1(net694),
    .S(net424),
    .X(_0119_));
 sg13g2_mux2_1 _0881_ (.A0(net726),
    .A1(net763),
    .S(net424),
    .X(_0120_));
 sg13g2_mux2_1 _0882_ (.A0(net696),
    .A1(net726),
    .S(net424),
    .X(_0121_));
 sg13g2_mux2_1 _0883_ (.A0(net523),
    .A1(net696),
    .S(net422),
    .X(_0122_));
 sg13g2_mux2_1 _0884_ (.A0(net222),
    .A1(net523),
    .S(net422),
    .X(_0123_));
 sg13g2_mux2_1 _0885_ (.A0(\i_main_reg.data_d[92] ),
    .A1(net222),
    .S(net422),
    .X(_0124_));
 sg13g2_mux2_1 _0886_ (.A0(net153),
    .A1(\i_main_reg.data_d[92] ),
    .S(net422),
    .X(_0125_));
 sg13g2_mux2_1 _0887_ (.A0(net233),
    .A1(net153),
    .S(net423),
    .X(_0126_));
 sg13g2_mux2_1 _0888_ (.A0(net122),
    .A1(net233),
    .S(net422),
    .X(_0127_));
 sg13g2_mux2_1 _0889_ (.A0(net100),
    .A1(net122),
    .S(net422),
    .X(_0128_));
 sg13g2_mux2_1 _0890_ (.A0(net94),
    .A1(net100),
    .S(net422),
    .X(_0129_));
 sg13g2_mux2_1 _0891_ (.A0(\i_main_reg.data_d[98] ),
    .A1(net94),
    .S(net422),
    .X(_0130_));
 sg13g2_mux2_1 _0892_ (.A0(\i_main_reg.data_d[99] ),
    .A1(net135),
    .S(net423),
    .X(_0131_));
 sg13g2_mux2_1 _0893_ (.A0(net226),
    .A1(net263),
    .S(net423),
    .X(_0132_));
 sg13g2_mux2_1 _0894_ (.A0(\i_main_reg.data_d[101] ),
    .A1(net226),
    .S(net423),
    .X(_0133_));
 sg13g2_mux2_1 _0895_ (.A0(\i_main_reg.data_d[102] ),
    .A1(net279),
    .S(net423),
    .X(_0134_));
 sg13g2_mux2_1 _0896_ (.A0(\i_main_reg.data_d[103] ),
    .A1(net649),
    .S(net424),
    .X(_0135_));
 sg13g2_mux2_1 _0897_ (.A0(\i_main_reg.data_d[104] ),
    .A1(net742),
    .S(net423),
    .X(_0136_));
 sg13g2_mux2_1 _0898_ (.A0(net588),
    .A1(\i_main_reg.data_d[104] ),
    .S(net423),
    .X(_0137_));
 sg13g2_mux2_1 _0899_ (.A0(net554),
    .A1(\i_main_reg.data_d[105] ),
    .S(net426),
    .X(_0138_));
 sg13g2_mux2_1 _0900_ (.A0(net623),
    .A1(net554),
    .S(net426),
    .X(_0139_));
 sg13g2_mux2_1 _0901_ (.A0(net673),
    .A1(net623),
    .S(net426),
    .X(_0140_));
 sg13g2_mux2_1 _0902_ (.A0(net745),
    .A1(net673),
    .S(net425),
    .X(_0141_));
 sg13g2_mux2_1 _0903_ (.A0(\i_main_reg.data_d[110] ),
    .A1(net745),
    .S(net425),
    .X(_0142_));
 sg13g2_mux2_1 _0904_ (.A0(\i_main_reg.data_d[111] ),
    .A1(net807),
    .S(net425),
    .X(_0143_));
 sg13g2_mux2_1 _0905_ (.A0(net204),
    .A1(\i_main_reg.data_d[111] ),
    .S(net421),
    .X(_0144_));
 sg13g2_mux2_1 _0906_ (.A0(net219),
    .A1(net204),
    .S(net421),
    .X(_0145_));
 sg13g2_mux2_1 _0907_ (.A0(net132),
    .A1(\i_main_reg.data_d[113] ),
    .S(net420),
    .X(_0146_));
 sg13g2_mux2_1 _0908_ (.A0(net281),
    .A1(net132),
    .S(net420),
    .X(_0147_));
 sg13g2_mux2_1 _0909_ (.A0(\i_main_reg.data_d[116] ),
    .A1(net281),
    .S(net420),
    .X(_0148_));
 sg13g2_mux2_1 _0910_ (.A0(net76),
    .A1(\i_main_reg.data_d[116] ),
    .S(net405),
    .X(_0149_));
 sg13g2_mux2_1 _0911_ (.A0(net113),
    .A1(net76),
    .S(net405),
    .X(_0150_));
 sg13g2_mux2_1 _0912_ (.A0(net191),
    .A1(net113),
    .S(net405),
    .X(_0151_));
 sg13g2_mux2_1 _0913_ (.A0(\i_main_reg.data_d[120] ),
    .A1(net191),
    .S(net405),
    .X(_0152_));
 sg13g2_mux2_1 _0914_ (.A0(\i_main_reg.data_d[121] ),
    .A1(net800),
    .S(net403),
    .X(_0153_));
 sg13g2_mux2_1 _0915_ (.A0(net766),
    .A1(net852),
    .S(net403),
    .X(_0154_));
 sg13g2_mux2_1 _0916_ (.A0(net727),
    .A1(net766),
    .S(net403),
    .X(_0155_));
 sg13g2_mux2_1 _0917_ (.A0(net682),
    .A1(net727),
    .S(net403),
    .X(_0156_));
 sg13g2_mux2_1 _0918_ (.A0(net594),
    .A1(net682),
    .S(net398),
    .X(_0157_));
 sg13g2_mux2_1 _0919_ (.A0(\i_main_reg.data_d[126] ),
    .A1(net594),
    .S(net398),
    .X(_0158_));
 sg13g2_mux2_1 _0920_ (.A0(net655),
    .A1(\i_main_reg.data_d[126] ),
    .S(net401),
    .X(_0159_));
 sg13g2_mux2_1 _0921_ (.A0(net62),
    .A1(\i_main_reg.data_d[127] ),
    .S(net400),
    .X(_0160_));
 sg13g2_mux2_1 _0922_ (.A0(net134),
    .A1(net62),
    .S(net400),
    .X(_0161_));
 sg13g2_mux2_1 _0923_ (.A0(net255),
    .A1(net134),
    .S(net400),
    .X(_0162_));
 sg13g2_mux2_1 _0924_ (.A0(\i_main_reg.data_d[131] ),
    .A1(net255),
    .S(net385),
    .X(_0163_));
 sg13g2_mux2_1 _0925_ (.A0(\i_main_reg.data_d[132] ),
    .A1(net257),
    .S(net386),
    .X(_0164_));
 sg13g2_mux2_1 _0926_ (.A0(\i_main_reg.data_d[133] ),
    .A1(net628),
    .S(net385),
    .X(_0165_));
 sg13g2_mux2_1 _0927_ (.A0(\i_main_reg.data_d[134] ),
    .A1(net722),
    .S(net385),
    .X(_0166_));
 sg13g2_mux2_1 _0928_ (.A0(net797),
    .A1(net845),
    .S(net383),
    .X(_0167_));
 sg13g2_mux2_1 _0929_ (.A0(\i_main_reg.data_d[136] ),
    .A1(net797),
    .S(net383),
    .X(_0168_));
 sg13g2_mux2_1 _0930_ (.A0(net144),
    .A1(\i_main_reg.data_d[136] ),
    .S(net383),
    .X(_0169_));
 sg13g2_mux2_1 _0931_ (.A0(net232),
    .A1(net144),
    .S(net383),
    .X(_0170_));
 sg13g2_mux2_1 _0932_ (.A0(net731),
    .A1(net232),
    .S(net384),
    .X(_0171_));
 sg13g2_mux2_1 _0933_ (.A0(net639),
    .A1(\i_main_reg.data_d[139] ),
    .S(net384),
    .X(_0172_));
 sg13g2_mux2_1 _0934_ (.A0(net767),
    .A1(net639),
    .S(net384),
    .X(_0173_));
 sg13g2_mux2_1 _0935_ (.A0(net527),
    .A1(\i_main_reg.data_d[141] ),
    .S(net384),
    .X(_0174_));
 sg13g2_mux2_1 _0936_ (.A0(net541),
    .A1(net527),
    .S(net392),
    .X(_0175_));
 sg13g2_mux2_1 _0937_ (.A0(net116),
    .A1(net541),
    .S(net392),
    .X(_0176_));
 sg13g2_mux2_1 _0938_ (.A0(\i_main_reg.data_d[145] ),
    .A1(net116),
    .S(net392),
    .X(_0177_));
 sg13g2_mux2_1 _0939_ (.A0(\i_main_reg.data_d[146] ),
    .A1(net557),
    .S(net392),
    .X(_0178_));
 sg13g2_mux2_1 _0940_ (.A0(net313),
    .A1(\i_main_reg.data_d[146] ),
    .S(net392),
    .X(_0179_));
 sg13g2_mux2_1 _0941_ (.A0(net186),
    .A1(net313),
    .S(net393),
    .X(_0180_));
 sg13g2_mux2_1 _0942_ (.A0(net180),
    .A1(net186),
    .S(net393),
    .X(_0181_));
 sg13g2_mux2_1 _0943_ (.A0(\i_main_reg.data_d[150] ),
    .A1(net180),
    .S(net393),
    .X(_0182_));
 sg13g2_mux2_1 _0944_ (.A0(net712),
    .A1(\i_main_reg.data_d[150] ),
    .S(net393),
    .X(_0183_));
 sg13g2_mux2_1 _0945_ (.A0(net788),
    .A1(net712),
    .S(net393),
    .X(_0184_));
 sg13g2_mux2_1 _0946_ (.A0(net729),
    .A1(\i_main_reg.data_d[152] ),
    .S(net396),
    .X(_0185_));
 sg13g2_mux2_1 _0947_ (.A0(net52),
    .A1(\i_main_reg.data_d[153] ),
    .S(net393),
    .X(_0186_));
 sg13g2_mux2_1 _0948_ (.A0(net112),
    .A1(net52),
    .S(net392),
    .X(_0187_));
 sg13g2_mux2_1 _0949_ (.A0(net157),
    .A1(net112),
    .S(net392),
    .X(_0188_));
 sg13g2_mux2_1 _0950_ (.A0(\i_main_reg.data_d[157] ),
    .A1(net157),
    .S(net392),
    .X(_0189_));
 sg13g2_mux2_1 _0951_ (.A0(\i_main_reg.data_d[158] ),
    .A1(net349),
    .S(net393),
    .X(_0190_));
 sg13g2_mux2_1 _0952_ (.A0(net343),
    .A1(\i_main_reg.data_d[158] ),
    .S(net387),
    .X(_0191_));
 sg13g2_mux2_1 _0953_ (.A0(net535),
    .A1(net343),
    .S(net388),
    .X(_0192_));
 sg13g2_mux2_1 _0954_ (.A0(net106),
    .A1(net535),
    .S(net388),
    .X(_0193_));
 sg13g2_mux2_1 _0955_ (.A0(\i_main_reg.data_d[162] ),
    .A1(net106),
    .S(net388),
    .X(_0194_));
 sg13g2_mux2_1 _0956_ (.A0(net114),
    .A1(net168),
    .S(net387),
    .X(_0195_));
 sg13g2_mux2_1 _0957_ (.A0(\i_main_reg.data_d[164] ),
    .A1(net114),
    .S(net387),
    .X(_0196_));
 sg13g2_mux2_1 _0958_ (.A0(\i_main_reg.data_d[165] ),
    .A1(net571),
    .S(net387),
    .X(_0197_));
 sg13g2_mux2_1 _0959_ (.A0(\i_main_reg.data_d[166] ),
    .A1(net614),
    .S(net372),
    .X(_0198_));
 sg13g2_mux2_1 _0960_ (.A0(\i_main_reg.data_d[167] ),
    .A1(net802),
    .S(net372),
    .X(_0199_));
 sg13g2_mux2_1 _0961_ (.A0(net760),
    .A1(\i_main_reg.data_d[167] ),
    .S(net372),
    .X(_0200_));
 sg13g2_mux2_1 _0962_ (.A0(net826),
    .A1(net760),
    .S(net372),
    .X(_0201_));
 sg13g2_mux2_1 _0963_ (.A0(net847),
    .A1(net826),
    .S(net372),
    .X(_0202_));
 sg13g2_mux2_1 _0964_ (.A0(net771),
    .A1(\i_main_reg.data_d[170] ),
    .S(net372),
    .X(_0203_));
 sg13g2_mux2_1 _0965_ (.A0(net603),
    .A1(\i_main_reg.data_d[171] ),
    .S(net368),
    .X(_0204_));
 sg13g2_mux2_1 _0966_ (.A0(net608),
    .A1(net603),
    .S(net368),
    .X(_0205_));
 sg13g2_mux2_1 _0967_ (.A0(net101),
    .A1(net608),
    .S(net368),
    .X(_0206_));
 sg13g2_mux2_1 _0968_ (.A0(\i_main_reg.data_d[175] ),
    .A1(net101),
    .S(net368),
    .X(_0207_));
 sg13g2_mux2_1 _0969_ (.A0(net328),
    .A1(net532),
    .S(net366),
    .X(_0208_));
 sg13g2_mux2_1 _0970_ (.A0(net209),
    .A1(net328),
    .S(net366),
    .X(_0209_));
 sg13g2_mux2_1 _0971_ (.A0(net142),
    .A1(net209),
    .S(net366),
    .X(_0210_));
 sg13g2_mux2_1 _0972_ (.A0(\i_main_reg.data_d[179] ),
    .A1(net142),
    .S(net367),
    .X(_0211_));
 sg13g2_mux2_1 _0973_ (.A0(net303),
    .A1(net559),
    .S(net367),
    .X(_0212_));
 sg13g2_mux2_1 _0974_ (.A0(net285),
    .A1(net303),
    .S(net367),
    .X(_0213_));
 sg13g2_mux2_1 _0975_ (.A0(\i_main_reg.data_d[182] ),
    .A1(net285),
    .S(net367),
    .X(_0214_));
 sg13g2_mux2_1 _0976_ (.A0(\i_main_reg.data_d[183] ),
    .A1(net777),
    .S(net370),
    .X(_0215_));
 sg13g2_mux2_1 _0977_ (.A0(\i_main_reg.data_d[184] ),
    .A1(net782),
    .S(net370),
    .X(_0216_));
 sg13g2_mux2_1 _0978_ (.A0(net818),
    .A1(\i_main_reg.data_d[184] ),
    .S(net370),
    .X(_0217_));
 sg13g2_mux2_1 _0979_ (.A0(net751),
    .A1(\i_main_reg.data_d[185] ),
    .S(net370),
    .X(_0218_));
 sg13g2_mux2_1 _0980_ (.A0(net340),
    .A1(\i_main_reg.data_d[186] ),
    .S(net370),
    .X(_0219_));
 sg13g2_mux2_1 _0981_ (.A0(net538),
    .A1(net340),
    .S(net370),
    .X(_0220_));
 sg13g2_mux2_1 _0982_ (.A0(net182),
    .A1(\i_main_reg.data_d[188] ),
    .S(net370),
    .X(_0221_));
 sg13g2_mux2_1 _0983_ (.A0(net315),
    .A1(net182),
    .S(net370),
    .X(_0222_));
 sg13g2_mux2_1 _0984_ (.A0(net125),
    .A1(net315),
    .S(net369),
    .X(_0223_));
 sg13g2_mux2_1 _0985_ (.A0(\i_main_reg.data_d[192] ),
    .A1(net125),
    .S(net369),
    .X(_0224_));
 sg13g2_mux2_1 _0986_ (.A0(net200),
    .A1(\i_main_reg.data_d[192] ),
    .S(net369),
    .X(_0225_));
 sg13g2_mux2_1 _0987_ (.A0(net236),
    .A1(net200),
    .S(net369),
    .X(_0226_));
 sg13g2_mux2_1 _0988_ (.A0(net272),
    .A1(net236),
    .S(net369),
    .X(_0227_));
 sg13g2_mux2_1 _0989_ (.A0(net224),
    .A1(net272),
    .S(net369),
    .X(_0228_));
 sg13g2_mux2_1 _0990_ (.A0(net206),
    .A1(net224),
    .S(net369),
    .X(_0229_));
 sg13g2_mux2_1 _0991_ (.A0(\i_main_reg.data_d[198] ),
    .A1(net206),
    .S(net369),
    .X(_0230_));
 sg13g2_mux2_1 _0992_ (.A0(\i_main_reg.data_d[199] ),
    .A1(net717),
    .S(net371),
    .X(_0231_));
 sg13g2_mux2_1 _0993_ (.A0(\i_main_reg.data_d[200] ),
    .A1(net856),
    .S(net371),
    .X(_0232_));
 sg13g2_mux2_1 _0994_ (.A0(net259),
    .A1(\i_main_reg.data_d[200] ),
    .S(net371),
    .X(_0233_));
 sg13g2_mux2_1 _0995_ (.A0(net165),
    .A1(\i_main_reg.data_d[201] ),
    .S(net371),
    .X(_0234_));
 sg13g2_mux2_1 _0996_ (.A0(net567),
    .A1(net165),
    .S(net371),
    .X(_0235_));
 sg13g2_mux2_1 _0997_ (.A0(net264),
    .A1(net567),
    .S(net374),
    .X(_0236_));
 sg13g2_mux2_1 _0998_ (.A0(net195),
    .A1(net264),
    .S(net375),
    .X(_0237_));
 sg13g2_mux2_1 _0999_ (.A0(\i_main_reg.data_d[206] ),
    .A1(net195),
    .S(net375),
    .X(_0238_));
 sg13g2_mux2_1 _1000_ (.A0(net542),
    .A1(\i_main_reg.data_d[206] ),
    .S(net375),
    .X(_0239_));
 sg13g2_mux2_1 _1001_ (.A0(net267),
    .A1(net542),
    .S(net375),
    .X(_0240_));
 sg13g2_mux2_1 _1002_ (.A0(net248),
    .A1(net267),
    .S(net375),
    .X(_0241_));
 sg13g2_mux2_1 _1003_ (.A0(\i_main_reg.data_d[210] ),
    .A1(net248),
    .S(net375),
    .X(_0242_));
 sg13g2_mux2_1 _1004_ (.A0(\i_main_reg.data_d[211] ),
    .A1(net331),
    .S(net375),
    .X(_0243_));
 sg13g2_mux2_1 _1005_ (.A0(\i_main_reg.data_d[212] ),
    .A1(net530),
    .S(net389),
    .X(_0244_));
 sg13g2_mux2_1 _1006_ (.A0(net562),
    .A1(net648),
    .S(net389),
    .X(_0245_));
 sg13g2_mux2_1 _1007_ (.A0(\i_main_reg.data_d[214] ),
    .A1(net562),
    .S(net389),
    .X(_0246_));
 sg13g2_mux2_1 _1008_ (.A0(net692),
    .A1(net699),
    .S(net389),
    .X(_0247_));
 sg13g2_mux2_1 _1009_ (.A0(net633),
    .A1(net692),
    .S(net389),
    .X(_0248_));
 sg13g2_mux2_1 _1010_ (.A0(\i_main_reg.data_d[217] ),
    .A1(net633),
    .S(net390),
    .X(_0249_));
 sg13g2_mux2_1 _1011_ (.A0(\i_main_reg.data_d[218] ),
    .A1(net735),
    .S(net390),
    .X(_0250_));
 sg13g2_mux2_1 _1012_ (.A0(net590),
    .A1(net849),
    .S(net390),
    .X(_0251_));
 sg13g2_mux2_1 _1013_ (.A0(net189),
    .A1(net590),
    .S(net389),
    .X(_0252_));
 sg13g2_mux2_1 _1014_ (.A0(\i_main_reg.data_d[221] ),
    .A1(net189),
    .S(net394),
    .X(_0253_));
 sg13g2_mux2_1 _1015_ (.A0(\i_main_reg.data_d[222] ),
    .A1(net637),
    .S(net394),
    .X(_0254_));
 sg13g2_mux2_1 _1016_ (.A0(net307),
    .A1(net657),
    .S(net394),
    .X(_0255_));
 sg13g2_mux2_1 _1017_ (.A0(net127),
    .A1(net307),
    .S(net394),
    .X(_0256_));
 sg13g2_mux2_1 _1018_ (.A0(net105),
    .A1(net127),
    .S(net394),
    .X(_0257_));
 sg13g2_mux2_1 _1019_ (.A0(net78),
    .A1(net105),
    .S(net394),
    .X(_0258_));
 sg13g2_mux2_1 _1020_ (.A0(\i_main_reg.data_d[227] ),
    .A1(net78),
    .S(net394),
    .X(_0259_));
 sg13g2_mux2_1 _1021_ (.A0(net147),
    .A1(\i_main_reg.data_d[227] ),
    .S(net394),
    .X(_0260_));
 sg13g2_mux2_1 _1022_ (.A0(net194),
    .A1(net147),
    .S(net395),
    .X(_0261_));
 sg13g2_mux2_1 _1023_ (.A0(net550),
    .A1(net194),
    .S(net395),
    .X(_0262_));
 sg13g2_mux2_1 _1024_ (.A0(\i_main_reg.data_d[231] ),
    .A1(net550),
    .S(net395),
    .X(_0263_));
 sg13g2_mux2_1 _1025_ (.A0(\i_main_reg.data_d[232] ),
    .A1(net836),
    .S(net390),
    .X(_0264_));
 sg13g2_mux2_1 _1026_ (.A0(net816),
    .A1(\i_main_reg.data_d[232] ),
    .S(net390),
    .X(_0265_));
 sg13g2_mux2_1 _1027_ (.A0(net832),
    .A1(net816),
    .S(net390),
    .X(_0266_));
 sg13g2_mux2_1 _1028_ (.A0(net764),
    .A1(\i_main_reg.data_d[234] ),
    .S(net389),
    .X(_0267_));
 sg13g2_mux2_1 _1029_ (.A0(net630),
    .A1(net764),
    .S(net389),
    .X(_0268_));
 sg13g2_mux2_1 _1030_ (.A0(net619),
    .A1(net630),
    .S(net376),
    .X(_0269_));
 sg13g2_mux2_1 _1031_ (.A0(\i_main_reg.data_d[238] ),
    .A1(net619),
    .S(net376),
    .X(_0270_));
 sg13g2_mux2_1 _1032_ (.A0(net601),
    .A1(net714),
    .S(net376),
    .X(_0271_));
 sg13g2_mux2_1 _1033_ (.A0(net539),
    .A1(net601),
    .S(net374),
    .X(_0272_));
 sg13g2_mux2_1 _1034_ (.A0(\i_main_reg.data_d[241] ),
    .A1(net539),
    .S(net374),
    .X(_0273_));
 sg13g2_mux2_1 _1035_ (.A0(\i_main_reg.data_d[242] ),
    .A1(net688),
    .S(net374),
    .X(_0274_));
 sg13g2_mux2_1 _1036_ (.A0(net616),
    .A1(net739),
    .S(net374),
    .X(_0275_));
 sg13g2_mux2_1 _1037_ (.A0(net237),
    .A1(net616),
    .S(net374),
    .X(_0276_));
 sg13g2_mux2_1 _1038_ (.A0(\i_main_reg.data_d[245] ),
    .A1(net237),
    .S(net374),
    .X(_0277_));
 sg13g2_mux2_1 _1039_ (.A0(\i_main_reg.data_d[246] ),
    .A1(net684),
    .S(net374),
    .X(_0278_));
 sg13g2_mux2_1 _1040_ (.A0(\i_main_reg.data_d[247] ),
    .A1(net740),
    .S(net372),
    .X(_0279_));
 sg13g2_mux2_1 _1041_ (.A0(net710),
    .A1(net770),
    .S(net372),
    .X(_0280_));
 sg13g2_mux2_1 _1042_ (.A0(\i_main_reg.data_d[249] ),
    .A1(net710),
    .S(net373),
    .X(_0281_));
 sg13g2_mux2_1 _1043_ (.A0(net706),
    .A1(net744),
    .S(net373),
    .X(_0282_));
 sg13g2_mux2_1 _1044_ (.A0(\i_main_reg.data_d[251] ),
    .A1(net706),
    .S(net373),
    .X(_0283_));
 sg13g2_mux2_1 _1045_ (.A0(net790),
    .A1(\i_main_reg.data_d[251] ),
    .S(net373),
    .X(_0284_));
 sg13g2_mux2_1 _1046_ (.A0(net635),
    .A1(\i_main_reg.data_d[252] ),
    .S(net387),
    .X(_0285_));
 sg13g2_mux2_1 _1047_ (.A0(net681),
    .A1(net635),
    .S(net387),
    .X(_0286_));
 sg13g2_mux2_1 _1048_ (.A0(net667),
    .A1(\i_main_reg.data_d[254] ),
    .S(net387),
    .X(_0287_));
 sg13g2_mux2_1 _1049_ (.A0(net261),
    .A1(\i_main_reg.data_d[255] ),
    .S(net387),
    .X(_0288_));
 sg13g2_mux2_1 _1050_ (.A0(net296),
    .A1(net261),
    .S(net388),
    .X(_0289_));
 sg13g2_mux2_1 _1051_ (.A0(net120),
    .A1(net296),
    .S(net388),
    .X(_0290_));
 sg13g2_mux2_1 _1052_ (.A0(\i_main_reg.data_d[259] ),
    .A1(net120),
    .S(net380),
    .X(_0291_));
 sg13g2_mux2_1 _1053_ (.A0(net70),
    .A1(net225),
    .S(net380),
    .X(_0292_));
 sg13g2_mux2_1 _1054_ (.A0(\i_main_reg.data_d[261] ),
    .A1(net70),
    .S(net380),
    .X(_0293_));
 sg13g2_mux2_1 _1055_ (.A0(\i_main_reg.data_d[262] ),
    .A1(net586),
    .S(net380),
    .X(_0294_));
 sg13g2_mux2_1 _1056_ (.A0(\i_main_reg.data_d[263] ),
    .A1(net822),
    .S(net380),
    .X(_0295_));
 sg13g2_mux2_1 _1057_ (.A0(net841),
    .A1(\i_main_reg.data_d[263] ),
    .S(net380),
    .X(_0296_));
 sg13g2_mux2_1 _1058_ (.A0(net773),
    .A1(\i_main_reg.data_d[264] ),
    .S(net363),
    .X(_0297_));
 sg13g2_mux2_1 _1059_ (.A0(net848),
    .A1(net773),
    .S(net363),
    .X(_0298_));
 sg13g2_mux2_1 _1060_ (.A0(net853),
    .A1(net848),
    .S(net365),
    .X(_0299_));
 sg13g2_mux2_1 _1061_ (.A0(net820),
    .A1(\i_main_reg.data_d[267] ),
    .S(net363),
    .X(_0300_));
 sg13g2_mux2_1 _1062_ (.A0(net838),
    .A1(net820),
    .S(net363),
    .X(_0301_));
 sg13g2_mux2_1 _1063_ (.A0(net198),
    .A1(\i_main_reg.data_d[269] ),
    .S(net364),
    .X(_0302_));
 sg13g2_mux2_1 _1064_ (.A0(net210),
    .A1(net198),
    .S(net364),
    .X(_0303_));
 sg13g2_mux2_1 _1065_ (.A0(net68),
    .A1(net210),
    .S(net364),
    .X(_0304_));
 sg13g2_mux2_1 _1066_ (.A0(\i_main_reg.data_d[273] ),
    .A1(net68),
    .S(net364),
    .X(_0305_));
 sg13g2_mux2_1 _1067_ (.A0(\i_main_reg.data_d[274] ),
    .A1(net611),
    .S(net360),
    .X(_0306_));
 sg13g2_mux2_1 _1068_ (.A0(net645),
    .A1(net698),
    .S(net368),
    .X(_0307_));
 sg13g2_mux2_1 _1069_ (.A0(net613),
    .A1(net645),
    .S(net368),
    .X(_0308_));
 sg13g2_mux2_1 _1070_ (.A0(net607),
    .A1(net613),
    .S(net366),
    .X(_0309_));
 sg13g2_mux2_1 _1071_ (.A0(net544),
    .A1(net607),
    .S(net366),
    .X(_0310_));
 sg13g2_mux2_1 _1072_ (.A0(net529),
    .A1(net544),
    .S(net366),
    .X(_0311_));
 sg13g2_mux2_1 _1073_ (.A0(net299),
    .A1(net529),
    .S(net366),
    .X(_0312_));
 sg13g2_mux2_1 _1074_ (.A0(net173),
    .A1(net299),
    .S(net366),
    .X(_0313_));
 sg13g2_mux2_1 _1075_ (.A0(\i_main_reg.data_d[282] ),
    .A1(net173),
    .S(net358),
    .X(_0314_));
 sg13g2_mux2_1 _1076_ (.A0(net337),
    .A1(net625),
    .S(net359),
    .X(_0315_));
 sg13g2_mux2_1 _1077_ (.A0(\i_main_reg.data_d[284] ),
    .A1(net337),
    .S(net359),
    .X(_0316_));
 sg13g2_mux2_1 _1078_ (.A0(net54),
    .A1(\i_main_reg.data_d[284] ),
    .S(net359),
    .X(_0317_));
 sg13g2_mux2_1 _1079_ (.A0(net247),
    .A1(net54),
    .S(net359),
    .X(_0318_));
 sg13g2_mux2_1 _1080_ (.A0(net243),
    .A1(\i_main_reg.data_d[286] ),
    .S(net359),
    .X(_0319_));
 sg13g2_mux2_1 _1081_ (.A0(net45),
    .A1(\i_main_reg.data_d[287] ),
    .S(net359),
    .X(_0320_));
 sg13g2_mux2_1 _1082_ (.A0(net188),
    .A1(net45),
    .S(net358),
    .X(_0321_));
 sg13g2_mux2_1 _1083_ (.A0(net252),
    .A1(net188),
    .S(net358),
    .X(_0322_));
 sg13g2_mux2_1 _1084_ (.A0(\i_main_reg.data_d[291] ),
    .A1(net252),
    .S(net358),
    .X(_0323_));
 sg13g2_mux2_1 _1085_ (.A0(net250),
    .A1(net295),
    .S(net358),
    .X(_0324_));
 sg13g2_mux2_1 _1086_ (.A0(\i_main_reg.data_d[293] ),
    .A1(net250),
    .S(net358),
    .X(_0325_));
 sg13g2_mux2_1 _1087_ (.A0(net679),
    .A1(net756),
    .S(net358),
    .X(_0326_));
 sg13g2_mux2_1 _1088_ (.A0(\i_main_reg.data_d[295] ),
    .A1(net679),
    .S(net355),
    .X(_0327_));
 sg13g2_mux2_1 _1089_ (.A0(net665),
    .A1(\i_main_reg.data_d[295] ),
    .S(net356),
    .X(_0328_));
 sg13g2_mux2_1 _1090_ (.A0(net775),
    .A1(net665),
    .S(net358),
    .X(_0329_));
 sg13g2_mux2_1 _1091_ (.A0(net644),
    .A1(net775),
    .S(net360),
    .X(_0330_));
 sg13g2_mux2_1 _1092_ (.A0(net606),
    .A1(net644),
    .S(net360),
    .X(_0331_));
 sg13g2_mux2_1 _1093_ (.A0(net521),
    .A1(net606),
    .S(net360),
    .X(_0332_));
 sg13g2_mux2_1 _1094_ (.A0(\i_main_reg.data_d[301] ),
    .A1(net521),
    .S(net360),
    .X(_0333_));
 sg13g2_mux2_1 _1095_ (.A0(net118),
    .A1(\i_main_reg.data_d[301] ),
    .S(net364),
    .X(_0334_));
 sg13g2_mux2_1 _1096_ (.A0(net187),
    .A1(net118),
    .S(net364),
    .X(_0335_));
 sg13g2_mux2_1 _1097_ (.A0(net631),
    .A1(net187),
    .S(net364),
    .X(_0336_));
 sg13g2_mux2_1 _1098_ (.A0(\i_main_reg.data_d[305] ),
    .A1(net631),
    .S(net364),
    .X(_0337_));
 sg13g2_mux2_1 _1099_ (.A0(net720),
    .A1(net799),
    .S(net363),
    .X(_0338_));
 sg13g2_mux2_1 _1100_ (.A0(\i_main_reg.data_d[307] ),
    .A1(net720),
    .S(net363),
    .X(_0339_));
 sg13g2_mux2_1 _1101_ (.A0(net690),
    .A1(\i_main_reg.data_d[307] ),
    .S(net363),
    .X(_0340_));
 sg13g2_mux2_1 _1102_ (.A0(net697),
    .A1(net690),
    .S(net363),
    .X(_0341_));
 sg13g2_mux2_1 _1103_ (.A0(net309),
    .A1(net697),
    .S(net397),
    .X(_0342_));
 sg13g2_mux2_1 _1104_ (.A0(net240),
    .A1(net309),
    .S(net378),
    .X(_0343_));
 sg13g2_mux2_1 _1105_ (.A0(net213),
    .A1(net240),
    .S(net378),
    .X(_0344_));
 sg13g2_mux2_1 _1106_ (.A0(\i_main_reg.data_d[313] ),
    .A1(net213),
    .S(net362),
    .X(_0345_));
 sg13g2_mux2_1 _1107_ (.A0(net202),
    .A1(\i_main_reg.data_d[313] ),
    .S(net362),
    .X(_0346_));
 sg13g2_mux2_1 _1108_ (.A0(net241),
    .A1(net202),
    .S(net362),
    .X(_0347_));
 sg13g2_mux2_1 _1109_ (.A0(\i_main_reg.data_d[316] ),
    .A1(net241),
    .S(net362),
    .X(_0348_));
 sg13g2_mux2_1 _1110_ (.A0(net329),
    .A1(\i_main_reg.data_d[316] ),
    .S(net361),
    .X(_0349_));
 sg13g2_mux2_1 _1111_ (.A0(net556),
    .A1(net329),
    .S(net361),
    .X(_0350_));
 sg13g2_mux2_1 _1112_ (.A0(net792),
    .A1(net556),
    .S(net361),
    .X(_0351_));
 sg13g2_mux2_1 _1113_ (.A0(net809),
    .A1(net792),
    .S(net361),
    .X(_0352_));
 sg13g2_mux2_1 _1114_ (.A0(net776),
    .A1(net809),
    .S(net357),
    .X(_0353_));
 sg13g2_mux2_1 _1115_ (.A0(net768),
    .A1(net776),
    .S(net357),
    .X(_0354_));
 sg13g2_mux2_1 _1116_ (.A0(net547),
    .A1(net768),
    .S(net357),
    .X(_0355_));
 sg13g2_mux2_1 _1117_ (.A0(\i_main_reg.data_d[324] ),
    .A1(net547),
    .S(net356),
    .X(_0356_));
 sg13g2_mux2_1 _1118_ (.A0(net749),
    .A1(net769),
    .S(net356),
    .X(_0357_));
 sg13g2_mux2_1 _1119_ (.A0(\i_main_reg.data_d[326] ),
    .A1(net749),
    .S(net356),
    .X(_0358_));
 sg13g2_mux2_1 _1120_ (.A0(\i_main_reg.data_d[327] ),
    .A1(net758),
    .S(net355),
    .X(_0359_));
 sg13g2_mux2_1 _1121_ (.A0(net700),
    .A1(\i_main_reg.data_d[327] ),
    .S(net355),
    .X(_0360_));
 sg13g2_mux2_1 _1122_ (.A0(net318),
    .A1(\i_main_reg.data_d[328] ),
    .S(net355),
    .X(_0361_));
 sg13g2_mux2_1 _1123_ (.A0(net297),
    .A1(\i_main_reg.data_d[329] ),
    .S(net355),
    .X(_0362_));
 sg13g2_mux2_1 _1124_ (.A0(net308),
    .A1(net297),
    .S(net355),
    .X(_0363_));
 sg13g2_mux2_1 _1125_ (.A0(net151),
    .A1(net308),
    .S(net355),
    .X(_0364_));
 sg13g2_mux2_1 _1126_ (.A0(\i_main_reg.data_d[333] ),
    .A1(net151),
    .S(net355),
    .X(_0365_));
 sg13g2_mux2_1 _1127_ (.A0(\i_main_reg.data_d[334] ),
    .A1(net321),
    .S(net357),
    .X(_0366_));
 sg13g2_mux2_1 _1128_ (.A0(net291),
    .A1(\i_main_reg.data_d[334] ),
    .S(net357),
    .X(_0367_));
 sg13g2_mux2_1 _1129_ (.A0(net108),
    .A1(\i_main_reg.data_d[335] ),
    .S(net357),
    .X(_0368_));
 sg13g2_mux2_1 _1130_ (.A0(net609),
    .A1(net108),
    .S(net361),
    .X(_0369_));
 sg13g2_mux2_1 _1131_ (.A0(net110),
    .A1(\i_main_reg.data_d[337] ),
    .S(net361),
    .X(_0370_));
 sg13g2_mux2_1 _1132_ (.A0(net193),
    .A1(net110),
    .S(net361),
    .X(_0371_));
 sg13g2_mux2_1 _1133_ (.A0(net312),
    .A1(net193),
    .S(net361),
    .X(_0372_));
 sg13g2_mux2_1 _1134_ (.A0(net66),
    .A1(\i_main_reg.data_d[340] ),
    .S(net362),
    .X(_0373_));
 sg13g2_mux2_1 _1135_ (.A0(net137),
    .A1(net66),
    .S(net362),
    .X(_0374_));
 sg13g2_mux2_1 _1136_ (.A0(net579),
    .A1(net137),
    .S(net362),
    .X(_0375_));
 sg13g2_mux2_1 _1137_ (.A0(net814),
    .A1(net579),
    .S(net362),
    .X(_0376_));
 sg13g2_mux2_1 _1138_ (.A0(net827),
    .A1(net814),
    .S(net378),
    .X(_0377_));
 sg13g2_mux2_1 _1139_ (.A0(net789),
    .A1(net827),
    .S(net378),
    .X(_0378_));
 sg13g2_mux2_1 _1140_ (.A0(net784),
    .A1(net789),
    .S(net378),
    .X(_0379_));
 sg13g2_mux2_1 _1141_ (.A0(net592),
    .A1(net784),
    .S(net378),
    .X(_0380_));
 sg13g2_mux2_1 _1142_ (.A0(\i_main_reg.data_d[349] ),
    .A1(net592),
    .S(net378),
    .X(_0381_));
 sg13g2_mux2_1 _1143_ (.A0(net283),
    .A1(\i_main_reg.data_d[349] ),
    .S(net379),
    .X(_0382_));
 sg13g2_mux2_1 _1144_ (.A0(net316),
    .A1(net283),
    .S(net379),
    .X(_0383_));
 sg13g2_mux2_1 _1145_ (.A0(\i_main_reg.data_d[352] ),
    .A1(net316),
    .S(net378),
    .X(_0384_));
 sg13g2_mux2_1 _1146_ (.A0(net323),
    .A1(net560),
    .S(net379),
    .X(_0385_));
 sg13g2_mux2_1 _1147_ (.A0(\i_main_reg.data_d[354] ),
    .A1(net323),
    .S(net379),
    .X(_0386_));
 sg13g2_mux2_1 _1148_ (.A0(net169),
    .A1(\i_main_reg.data_d[354] ),
    .S(net381),
    .X(_0387_));
 sg13g2_mux2_1 _1149_ (.A0(net239),
    .A1(net169),
    .S(net381),
    .X(_0388_));
 sg13g2_mux2_1 _1150_ (.A0(net60),
    .A1(\i_main_reg.data_d[356] ),
    .S(net381),
    .X(_0389_));
 sg13g2_mux2_1 _1151_ (.A0(net320),
    .A1(net60),
    .S(net381),
    .X(_0390_));
 sg13g2_mux2_1 _1152_ (.A0(net270),
    .A1(\i_main_reg.data_d[358] ),
    .S(net382),
    .X(_0391_));
 sg13g2_mux2_1 _1153_ (.A0(net273),
    .A1(net270),
    .S(net382),
    .X(_0392_));
 sg13g2_mux2_1 _1154_ (.A0(net56),
    .A1(\i_main_reg.data_d[360] ),
    .S(net382),
    .X(_0393_));
 sg13g2_mux2_1 _1155_ (.A0(net178),
    .A1(net56),
    .S(net382),
    .X(_0394_));
 sg13g2_mux2_1 _1156_ (.A0(net301),
    .A1(net178),
    .S(net399),
    .X(_0395_));
 sg13g2_mux2_1 _1157_ (.A0(net171),
    .A1(net301),
    .S(net399),
    .X(_0396_));
 sg13g2_mux2_1 _1158_ (.A0(\i_main_reg.data_d[365] ),
    .A1(net171),
    .S(net399),
    .X(_0397_));
 sg13g2_mux2_1 _1159_ (.A0(net90),
    .A1(net278),
    .S(net398),
    .X(_0398_));
 sg13g2_mux2_1 _1160_ (.A0(\i_main_reg.data_d[367] ),
    .A1(net90),
    .S(net398),
    .X(_0399_));
 sg13g2_mux2_1 _1161_ (.A0(net211),
    .A1(net306),
    .S(net398),
    .X(_0400_));
 sg13g2_mux2_1 _1162_ (.A0(\i_main_reg.data_d[369] ),
    .A1(net211),
    .S(net398),
    .X(_0401_));
 sg13g2_mux2_1 _1163_ (.A0(net74),
    .A1(\i_main_reg.data_d[369] ),
    .S(net402),
    .X(_0402_));
 sg13g2_mux2_1 _1164_ (.A0(net208),
    .A1(net74),
    .S(net402),
    .X(_0403_));
 sg13g2_mux2_1 _1165_ (.A0(net177),
    .A1(net208),
    .S(net402),
    .X(_0404_));
 sg13g2_mux2_1 _1166_ (.A0(net130),
    .A1(net177),
    .S(net402),
    .X(_0405_));
 sg13g2_mux2_1 _1167_ (.A0(\i_main_reg.data_d[374] ),
    .A1(net130),
    .S(net402),
    .X(_0406_));
 sg13g2_mux2_1 _1168_ (.A0(net566),
    .A1(net605),
    .S(net402),
    .X(_0407_));
 sg13g2_mux2_1 _1169_ (.A0(net536),
    .A1(net566),
    .S(net403),
    .X(_0408_));
 sg13g2_mux2_1 _1170_ (.A0(\i_main_reg.data_d[377] ),
    .A1(net536),
    .S(net402),
    .X(_0409_));
 sg13g2_mux2_1 _1171_ (.A0(\i_main_reg.data_d[378] ),
    .A1(net584),
    .S(net402),
    .X(_0410_));
 sg13g2_mux2_1 _1172_ (.A0(\i_main_reg.data_d[379] ),
    .A1(net795),
    .S(net398),
    .X(_0411_));
 sg13g2_mux2_1 _1173_ (.A0(net325),
    .A1(\i_main_reg.data_d[379] ),
    .S(net398),
    .X(_0412_));
 sg13g2_mux2_1 _1174_ (.A0(net82),
    .A1(\i_main_reg.data_d[380] ),
    .S(net399),
    .X(_0413_));
 sg13g2_mux2_1 _1175_ (.A0(net179),
    .A1(net82),
    .S(net399),
    .X(_0414_));
 sg13g2_mux2_1 _1176_ (.A0(net159),
    .A1(net179),
    .S(net399),
    .X(_0415_));
 sg13g2_mux2_1 _1177_ (.A0(\i_main_reg.data_d[384] ),
    .A1(net159),
    .S(net399),
    .X(_0416_));
 sg13g2_mux2_1 _1178_ (.A0(\i_main_reg.data_d[385] ),
    .A1(net162),
    .S(net382),
    .X(_0417_));
 sg13g2_mux2_1 _1179_ (.A0(net339),
    .A1(net646),
    .S(net382),
    .X(_0418_));
 sg13g2_mux2_1 _1180_ (.A0(net64),
    .A1(net339),
    .S(net382),
    .X(_0419_));
 sg13g2_mux2_1 _1181_ (.A0(\i_main_reg.data_d[388] ),
    .A1(net64),
    .S(net381),
    .X(_0420_));
 sg13g2_mux2_1 _1182_ (.A0(net624),
    .A1(net738),
    .S(net381),
    .X(_0421_));
 sg13g2_mux2_1 _1183_ (.A0(net583),
    .A1(net624),
    .S(net381),
    .X(_0422_));
 sg13g2_mux2_1 _1184_ (.A0(net524),
    .A1(net583),
    .S(net381),
    .X(_0423_));
 sg13g2_mux2_1 _1185_ (.A0(\i_main_reg.data_d[392] ),
    .A1(net524),
    .S(net383),
    .X(_0424_));
 sg13g2_mux2_1 _1186_ (.A0(net573),
    .A1(\i_main_reg.data_d[392] ),
    .S(net383),
    .X(_0425_));
 sg13g2_mux2_1 _1187_ (.A0(net641),
    .A1(net573),
    .S(net383),
    .X(_0426_));
 sg13g2_mux2_1 _1188_ (.A0(net757),
    .A1(net641),
    .S(net383),
    .X(_0427_));
 sg13g2_mux2_1 _1189_ (.A0(net626),
    .A1(\i_main_reg.data_d[395] ),
    .S(net385),
    .X(_0428_));
 sg13g2_mux2_1 _1190_ (.A0(net50),
    .A1(\i_main_reg.data_d[396] ),
    .S(net385),
    .X(_0429_));
 sg13g2_mux2_1 _1191_ (.A0(net164),
    .A1(net50),
    .S(net385),
    .X(_0430_));
 sg13g2_mux2_1 _1192_ (.A0(net140),
    .A1(net164),
    .S(net400),
    .X(_0431_));
 sg13g2_mux2_1 _1193_ (.A0(\i_main_reg.data_d[400] ),
    .A1(net140),
    .S(net400),
    .X(_0432_));
 sg13g2_mux2_1 _1194_ (.A0(net568),
    .A1(net693),
    .S(net400),
    .X(_0433_));
 sg13g2_mux2_1 _1195_ (.A0(net526),
    .A1(net568),
    .S(net400),
    .X(_0434_));
 sg13g2_mux2_1 _1196_ (.A0(net245),
    .A1(net526),
    .S(net400),
    .X(_0435_));
 sg13g2_mux2_1 _1197_ (.A0(\i_main_reg.data_d[404] ),
    .A1(net245),
    .S(net401),
    .X(_0436_));
 sg13g2_mux2_1 _1198_ (.A0(\i_main_reg.data_d[405] ),
    .A1(net780),
    .S(net401),
    .X(_0437_));
 sg13g2_mux2_1 _1199_ (.A0(net810),
    .A1(\i_main_reg.data_d[405] ),
    .S(net401),
    .X(_0438_));
 sg13g2_mux2_1 _1200_ (.A0(net813),
    .A1(net810),
    .S(net401),
    .X(_0439_));
 sg13g2_mux2_1 _1201_ (.A0(net844),
    .A1(net813),
    .S(net404),
    .X(_0440_));
 sg13g2_mux2_1 _1202_ (.A0(net228),
    .A1(\i_main_reg.data_d[408] ),
    .S(net404),
    .X(_0441_));
 sg13g2_mux2_1 _1203_ (.A0(net220),
    .A1(net228),
    .S(net404),
    .X(_0442_));
 sg13g2_mux2_1 _1204_ (.A0(\i_main_reg.data_d[411] ),
    .A1(net220),
    .S(net404),
    .X(_0443_));
 sg13g2_mux2_1 _1205_ (.A0(\i_main_reg.data_d[412] ),
    .A1(net659),
    .S(net404),
    .X(_0444_));
 sg13g2_mux2_1 _1206_ (.A0(net351),
    .A1(net787),
    .S(net404),
    .X(_0445_));
 sg13g2_mux2_1 _1207_ (.A0(net276),
    .A1(net351),
    .S(net404),
    .X(_0446_));
 sg13g2_mux2_1 _1208_ (.A0(\i_main_reg.data_d[415] ),
    .A1(net276),
    .S(net404),
    .X(_0447_));
 sg13g2_mux2_1 _1209_ (.A0(net287),
    .A1(\i_main_reg.data_d[415] ),
    .S(net412),
    .X(_0448_));
 sg13g2_mux2_1 _1210_ (.A0(net591),
    .A1(net287),
    .S(net412),
    .X(_0449_));
 sg13g2_mux2_1 _1211_ (.A0(net719),
    .A1(net591),
    .S(net407),
    .X(_0450_));
 sg13g2_mux2_1 _1212_ (.A0(net724),
    .A1(net719),
    .S(net407),
    .X(_0451_));
 sg13g2_mux2_1 _1213_ (.A0(net161),
    .A1(net724),
    .S(net407),
    .X(_0452_));
 sg13g2_mux2_1 _1214_ (.A0(net72),
    .A1(net161),
    .S(net407),
    .X(_0453_));
 sg13g2_mux2_1 _1215_ (.A0(\i_main_reg.data_d[422] ),
    .A1(net72),
    .S(net407),
    .X(_0454_));
 sg13g2_mux2_1 _1216_ (.A0(\i_main_reg.data_d[423] ),
    .A1(net617),
    .S(net408),
    .X(_0455_));
 sg13g2_mux2_1 _1217_ (.A0(net747),
    .A1(\i_main_reg.data_d[423] ),
    .S(net408),
    .X(_0456_));
 sg13g2_mux2_1 _1218_ (.A0(net577),
    .A1(\i_main_reg.data_d[424] ),
    .S(net408),
    .X(_0457_));
 sg13g2_mux2_1 _1219_ (.A0(net128),
    .A1(net577),
    .S(net408),
    .X(_0458_));
 sg13g2_mux2_1 _1220_ (.A0(\i_main_reg.data_d[427] ),
    .A1(net128),
    .S(net408),
    .X(_0459_));
 sg13g2_mux2_1 _1221_ (.A0(\i_main_reg.data_d[428] ),
    .A1(net335),
    .S(net408),
    .X(_0460_));
 sg13g2_mux2_1 _1222_ (.A0(net651),
    .A1(net815),
    .S(net407),
    .X(_0461_));
 sg13g2_mux2_1 _1223_ (.A0(net580),
    .A1(net651),
    .S(net407),
    .X(_0462_));
 sg13g2_mux2_1 _1224_ (.A0(net300),
    .A1(net580),
    .S(net407),
    .X(_0463_));
 sg13g2_mux2_1 _1225_ (.A0(net167),
    .A1(net300),
    .S(net410),
    .X(_0464_));
 sg13g2_mux2_1 _1226_ (.A0(net96),
    .A1(net167),
    .S(net410),
    .X(_0465_));
 sg13g2_mux2_1 _1227_ (.A0(\i_main_reg.data_d[434] ),
    .A1(net96),
    .S(net414),
    .X(_0466_));
 sg13g2_mux2_1 _1228_ (.A0(net610),
    .A1(net683),
    .S(net414),
    .X(_0467_));
 sg13g2_mux2_1 _1229_ (.A0(net533),
    .A1(net610),
    .S(net414),
    .X(_0468_));
 sg13g2_mux2_1 _1230_ (.A0(\i_main_reg.data_d[437] ),
    .A1(net533),
    .S(net414),
    .X(_0469_));
 sg13g2_mux2_1 _1231_ (.A0(net92),
    .A1(\i_main_reg.data_d[437] ),
    .S(net415),
    .X(_0470_));
 sg13g2_mux2_1 _1232_ (.A0(net302),
    .A1(net92),
    .S(net415),
    .X(_0471_));
 sg13g2_mux2_1 _1233_ (.A0(net138),
    .A1(\i_main_reg.data_d[439] ),
    .S(net415),
    .X(_0472_));
 sg13g2_mux2_1 _1234_ (.A0(net197),
    .A1(net138),
    .S(net415),
    .X(_0473_));
 sg13g2_mux2_1 _1235_ (.A0(net327),
    .A1(net197),
    .S(net429),
    .X(_0474_));
 sg13g2_mux2_1 _1236_ (.A0(net664),
    .A1(net327),
    .S(net429),
    .X(_0475_));
 sg13g2_mux2_1 _1237_ (.A0(net289),
    .A1(net664),
    .S(net429),
    .X(_0476_));
 sg13g2_mux2_1 _1238_ (.A0(\i_main_reg.data_d[445] ),
    .A1(net289),
    .S(net430),
    .X(_0477_));
 sg13g2_mux2_1 _1239_ (.A0(net35),
    .A1(net661),
    .S(net429),
    .X(_0478_));
 sg13g2_nand2_1 _1240_ (.Y(_0584_),
    .A(net35),
    .B(net431));
 sg13g2_xnor2_1 _1241_ (.Y(_0585_),
    .A(net435),
    .B(carry_q));
 sg13g2_xnor2_1 _1242_ (.Y(_0586_),
    .A(previous_bit_q),
    .B(_0585_));
 sg13g2_nor2_1 _1243_ (.A(_0623_),
    .B(_0558_),
    .Y(_0587_));
 sg13g2_a221oi_1 _1244_ (.B2(_0622_),
    .C1(_0587_),
    .B1(_0586_),
    .A1(net436),
    .Y(_0588_),
    .A2(_0483_));
 sg13g2_o21ai_1 _1245_ (.B1(_0582_),
    .Y(_0589_),
    .A1(net1),
    .A2(_0627_));
 sg13g2_o21ai_1 _1246_ (.B1(_0584_),
    .Y(_0479_),
    .A1(_0588_),
    .A2(_0589_));
 sg13g2_nand2_1 _1247_ (.Y(_0590_),
    .A(net345),
    .B(net33));
 sg13g2_a21o_1 _1248_ (.A2(_0590_),
    .A1(net435),
    .B1(_0615_),
    .X(_0591_));
 sg13g2_nand3_1 _1249_ (.B(_0579_),
    .C(_0591_),
    .A(_0482_),
    .Y(_0592_));
 sg13g2_or2_1 _1250_ (.X(_0593_),
    .B(_0592_),
    .A(_0615_));
 sg13g2_nand2_1 _1251_ (.Y(_0594_),
    .A(net33),
    .B(_0592_));
 sg13g2_o21ai_1 _1252_ (.B1(_0594_),
    .Y(_0480_),
    .A1(net33),
    .A2(_0593_));
 sg13g2_nand2_1 _1253_ (.Y(_0595_),
    .A(net345),
    .B(_0592_));
 sg13g2_nand2b_1 _1254_ (.Y(_0596_),
    .B(_0590_),
    .A_N(_0617_));
 sg13g2_o21ai_1 _1255_ (.B1(_0595_),
    .Y(_0481_),
    .A1(_0593_),
    .A2(_0596_));
 sg13g2_dfrbpq_2 _1256_ (.RESET_B(net515),
    .D(net671),
    .Q(\i_step_counter.data_o ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _1257_ (.RESET_B(net515),
    .D(net878),
    .Q(\i_step_counter.data_d[0] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _1258_ (.RESET_B(net515),
    .D(net866),
    .Q(\i_step_counter.data_d[1] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _1259_ (.RESET_B(net515),
    .D(net873),
    .Q(\i_step_counter.data_d[2] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _1260_ (.RESET_B(net514),
    .D(net59),
    .Q(\i_step_counter.data_d[3] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _1261_ (.RESET_B(net514),
    .D(net876),
    .Q(\i_step_counter.data_d[4] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _1262_ (.RESET_B(net514),
    .D(net42),
    .Q(\i_step_counter.data_d[5] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _1263_ (.RESET_B(net514),
    .D(net835),
    .Q(\i_step_counter.data_d[6] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _1264_ (.RESET_B(net514),
    .D(net794),
    .Q(\i_step_counter.data_d[7] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _1265_ (.RESET_B(net513),
    .D(net868),
    .Q(\i_step_counter.data_d[8] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _1266_ (.RESET_B(net513),
    .D(net44),
    .Q(\i_step_counter.data_d[9] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _1267_ (.RESET_B(net513),
    .D(net860),
    .Q(\i_step_counter.data_d[10] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _1268_ (.RESET_B(net513),
    .D(net855),
    .Q(\i_step_counter.data_d[11] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _1269_ (.RESET_B(net514),
    .D(net863),
    .Q(\i_step_counter.data_d[12] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _1270_ (.RESET_B(net514),
    .D(net806),
    .Q(\i_step_counter.data_d[13] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _1271_ (.RESET_B(net514),
    .D(_0015_),
    .Q(\i_step_counter.data_d[14] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _1272_ (.RESET_B(net515),
    .D(net99),
    .Q(finished_q),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _1273_ (.RESET_B(net515),
    .D(net28),
    .Q(overflow_q),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _1274_ (.RESET_B(net516),
    .D(net825),
    .Q(carry_q),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _1275_ (.RESET_B(net516),
    .D(net880),
    .Q(previous_bit_q),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _1276_ (.RESET_B(net516),
    .D(net30),
    .Q(\bit_counter_q[0] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _1277_ (.RESET_B(net516),
    .D(_0021_),
    .Q(\bit_counter_q[1] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _1278_ (.RESET_B(net516),
    .D(net32),
    .Q(\bit_counter_q[2] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _1279_ (.RESET_B(net518),
    .D(_0023_),
    .Q(\bit_counter_q[3] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _1280_ (.RESET_B(net518),
    .D(_0024_),
    .Q(\bit_counter_q[4] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _1281_ (.RESET_B(net516),
    .D(net851),
    .Q(\bit_counter_q[5] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _1282_ (.RESET_B(net517),
    .D(_0026_),
    .Q(\bit_counter_q[6] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _1283_ (.RESET_B(net517),
    .D(_0027_),
    .Q(\bit_counter_q[7] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _1284_ (.RESET_B(net517),
    .D(net49),
    .Q(\bit_counter_q[8] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _1285_ (.RESET_B(net517),
    .D(_0029_),
    .Q(\bit_counter_q[9] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _1286_ (.RESET_B(net516),
    .D(_0030_),
    .Q(\state_q[0] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _1287_ (.RESET_B(net516),
    .D(_0031_),
    .Q(\state_q[1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _1288_ (.RESET_B(net517),
    .D(_0032_),
    .Q(\i_main_reg.data_o ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _1289_ (.RESET_B(net512),
    .D(_0033_),
    .Q(\i_main_reg.data_d[0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _1290_ (.RESET_B(net512),
    .D(net89),
    .Q(\i_main_reg.data_d[1] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _1291_ (.RESET_B(net513),
    .D(_0035_),
    .Q(\i_main_reg.data_d[2] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _1292_ (.RESET_B(net512),
    .D(net597),
    .Q(\i_main_reg.data_d[3] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _1293_ (.RESET_B(net512),
    .D(net709),
    .Q(\i_main_reg.data_d[4] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _1294_ (.RESET_B(net512),
    .D(net275),
    .Q(\i_main_reg.data_d[5] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _1295_ (.RESET_B(net497),
    .D(_0039_),
    .Q(\i_main_reg.data_d[6] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _1296_ (.RESET_B(net497),
    .D(_0040_),
    .Q(\i_main_reg.data_d[7] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _1297_ (.RESET_B(net497),
    .D(_0041_),
    .Q(\i_main_reg.data_d[8] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _1298_ (.RESET_B(net496),
    .D(net570),
    .Q(\i_main_reg.data_d[9] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _1299_ (.RESET_B(net496),
    .D(_0043_),
    .Q(\i_main_reg.data_d[10] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _1300_ (.RESET_B(net496),
    .D(net305),
    .Q(\i_main_reg.data_d[11] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _1301_ (.RESET_B(net496),
    .D(net104),
    .Q(\i_main_reg.data_d[12] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _1302_ (.RESET_B(net493),
    .D(_0046_),
    .Q(\i_main_reg.data_d[13] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _1303_ (.RESET_B(net493),
    .D(net81),
    .Q(\i_main_reg.data_d[14] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _1304_ (.RESET_B(net493),
    .D(net176),
    .Q(\i_main_reg.data_d[15] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _1305_ (.RESET_B(net493),
    .D(net677),
    .Q(\i_main_reg.data_d[16] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _1306_ (.RESET_B(net493),
    .D(net546),
    .Q(\i_main_reg.data_d[17] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _1307_ (.RESET_B(net492),
    .D(_0051_),
    .Q(\i_main_reg.data_d[18] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _1308_ (.RESET_B(net492),
    .D(net185),
    .Q(\i_main_reg.data_d[19] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _1309_ (.RESET_B(net492),
    .D(net231),
    .Q(\i_main_reg.data_d[20] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _1310_ (.RESET_B(net492),
    .D(_0054_),
    .Q(\i_main_reg.data_d[21] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _1311_ (.RESET_B(net492),
    .D(_0055_),
    .Q(\i_main_reg.data_d[22] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _1312_ (.RESET_B(net492),
    .D(net266),
    .Q(\i_main_reg.data_d[23] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _1313_ (.RESET_B(net492),
    .D(net653),
    .Q(\i_main_reg.data_d[24] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _1314_ (.RESET_B(net492),
    .D(_0058_),
    .Q(\i_main_reg.data_d[25] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _1315_ (.RESET_B(net489),
    .D(_0059_),
    .Q(\i_main_reg.data_d[26] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1316_ (.RESET_B(net490),
    .D(net217),
    .Q(\i_main_reg.data_d[27] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _1317_ (.RESET_B(net490),
    .D(_0061_),
    .Q(\i_main_reg.data_d[28] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _1318_ (.RESET_B(net490),
    .D(net235),
    .Q(\i_main_reg.data_d[29] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _1319_ (.RESET_B(net494),
    .D(net565),
    .Q(\i_main_reg.data_d[30] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _1320_ (.RESET_B(net494),
    .D(net576),
    .Q(\i_main_reg.data_d[31] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _1321_ (.RESET_B(net494),
    .D(net150),
    .Q(\i_main_reg.data_d[32] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _1322_ (.RESET_B(net494),
    .D(_0066_),
    .Q(\i_main_reg.data_d[33] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _1323_ (.RESET_B(net495),
    .D(_0067_),
    .Q(\i_main_reg.data_d[34] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _1324_ (.RESET_B(net495),
    .D(_0068_),
    .Q(\i_main_reg.data_d[35] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _1325_ (.RESET_B(net495),
    .D(net829),
    .Q(\i_main_reg.data_d[36] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _1326_ (.RESET_B(net495),
    .D(net582),
    .Q(\i_main_reg.data_d[37] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _1327_ (.RESET_B(net494),
    .D(net124),
    .Q(\i_main_reg.data_d[38] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _1328_ (.RESET_B(net494),
    .D(_0072_),
    .Q(\i_main_reg.data_d[39] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _1329_ (.RESET_B(net495),
    .D(_0073_),
    .Q(\i_main_reg.data_d[40] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _1330_ (.RESET_B(net494),
    .D(_0074_),
    .Q(\i_main_reg.data_d[41] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _1331_ (.RESET_B(net504),
    .D(net156),
    .Q(\i_main_reg.data_d[42] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _1332_ (.RESET_B(net504),
    .D(_0076_),
    .Q(\i_main_reg.data_d[43] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1333_ (.RESET_B(net504),
    .D(_0077_),
    .Q(\i_main_reg.data_d[44] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _1334_ (.RESET_B(net504),
    .D(_0078_),
    .Q(\i_main_reg.data_d[45] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _1335_ (.RESET_B(net504),
    .D(net294),
    .Q(\i_main_reg.data_d[46] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1336_ (.RESET_B(net505),
    .D(_0080_),
    .Q(\i_main_reg.data_d[47] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1337_ (.RESET_B(net503),
    .D(_0081_),
    .Q(\i_main_reg.data_d[48] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _1338_ (.RESET_B(net503),
    .D(net599),
    .Q(\i_main_reg.data_d[49] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _1339_ (.RESET_B(net509),
    .D(_0083_),
    .Q(\i_main_reg.data_d[50] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _1340_ (.RESET_B(net509),
    .D(net643),
    .Q(\i_main_reg.data_d[51] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _1341_ (.RESET_B(net510),
    .D(net311),
    .Q(\i_main_reg.data_d[52] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _1342_ (.RESET_B(net510),
    .D(_0086_),
    .Q(\i_main_reg.data_d[53] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _1343_ (.RESET_B(net510),
    .D(_0087_),
    .Q(\i_main_reg.data_d[54] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _1344_ (.RESET_B(net510),
    .D(_0088_),
    .Q(\i_main_reg.data_d[55] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _1345_ (.RESET_B(net510),
    .D(net85),
    .Q(\i_main_reg.data_d[56] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _1346_ (.RESET_B(net511),
    .D(_0090_),
    .Q(\i_main_reg.data_d[57] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1347_ (.RESET_B(net509),
    .D(net622),
    .Q(\i_main_reg.data_d[58] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1348_ (.RESET_B(net509),
    .D(net269),
    .Q(\i_main_reg.data_d[59] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1349_ (.RESET_B(net509),
    .D(_0093_),
    .Q(\i_main_reg.data_d[60] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1350_ (.RESET_B(net503),
    .D(_0094_),
    .Q(\i_main_reg.data_d[61] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _1351_ (.RESET_B(net503),
    .D(_0095_),
    .Q(\i_main_reg.data_d[62] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _1352_ (.RESET_B(net503),
    .D(_0096_),
    .Q(\i_main_reg.data_d[63] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1353_ (.RESET_B(net503),
    .D(_0097_),
    .Q(\i_main_reg.data_d[64] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1354_ (.RESET_B(net502),
    .D(_0098_),
    .Q(\i_main_reg.data_d[65] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _1355_ (.RESET_B(net502),
    .D(net687),
    .Q(\i_main_reg.data_d[66] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _1356_ (.RESET_B(net502),
    .D(net840),
    .Q(\i_main_reg.data_d[67] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _1357_ (.RESET_B(net502),
    .D(net831),
    .Q(\i_main_reg.data_d[68] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _1358_ (.RESET_B(net501),
    .D(_0102_),
    .Q(\i_main_reg.data_d[69] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1359_ (.RESET_B(net501),
    .D(_0103_),
    .Q(\i_main_reg.data_d[70] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1360_ (.RESET_B(net501),
    .D(net786),
    .Q(\i_main_reg.data_d[71] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1361_ (.RESET_B(net486),
    .D(net675),
    .Q(\i_main_reg.data_d[72] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1362_ (.RESET_B(net486),
    .D(net87),
    .Q(\i_main_reg.data_d[73] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1363_ (.RESET_B(net486),
    .D(_0107_),
    .Q(\i_main_reg.data_d[74] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1364_ (.RESET_B(net486),
    .D(net334),
    .Q(\i_main_reg.data_d[75] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1365_ (.RESET_B(net486),
    .D(_0109_),
    .Q(\i_main_reg.data_d[76] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1366_ (.RESET_B(net486),
    .D(net348),
    .Q(\i_main_reg.data_d[77] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1367_ (.RESET_B(net501),
    .D(_0111_),
    .Q(\i_main_reg.data_d[78] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1368_ (.RESET_B(net501),
    .D(_0112_),
    .Q(\i_main_reg.data_d[79] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1369_ (.RESET_B(net501),
    .D(_0113_),
    .Q(\i_main_reg.data_d[80] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1370_ (.RESET_B(net501),
    .D(net734),
    .Q(\i_main_reg.data_d[81] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1371_ (.RESET_B(net501),
    .D(_0115_),
    .Q(\i_main_reg.data_d[82] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1372_ (.RESET_B(net502),
    .D(_0116_),
    .Q(\i_main_reg.data_d[83] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _1373_ (.RESET_B(net502),
    .D(_0117_),
    .Q(\i_main_reg.data_d[84] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1374_ (.RESET_B(net502),
    .D(net663),
    .Q(\i_main_reg.data_d[85] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1375_ (.RESET_B(net502),
    .D(net695),
    .Q(\i_main_reg.data_d[86] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1376_ (.RESET_B(net508),
    .D(_0120_),
    .Q(\i_main_reg.data_d[87] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _1377_ (.RESET_B(net508),
    .D(_0121_),
    .Q(\i_main_reg.data_d[88] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1378_ (.RESET_B(net508),
    .D(_0122_),
    .Q(\i_main_reg.data_d[89] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _1379_ (.RESET_B(net508),
    .D(_0123_),
    .Q(\i_main_reg.data_d[90] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _1380_ (.RESET_B(net506),
    .D(net223),
    .Q(\i_main_reg.data_d[91] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1381_ (.RESET_B(net506),
    .D(net154),
    .Q(\i_main_reg.data_d[92] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1382_ (.RESET_B(net506),
    .D(_0126_),
    .Q(\i_main_reg.data_d[93] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1383_ (.RESET_B(net506),
    .D(_0127_),
    .Q(\i_main_reg.data_d[94] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1384_ (.RESET_B(net506),
    .D(_0128_),
    .Q(\i_main_reg.data_d[95] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1385_ (.RESET_B(net506),
    .D(_0129_),
    .Q(\i_main_reg.data_d[96] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1386_ (.RESET_B(net506),
    .D(net95),
    .Q(\i_main_reg.data_d[97] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1387_ (.RESET_B(net506),
    .D(net136),
    .Q(\i_main_reg.data_d[98] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1388_ (.RESET_B(net507),
    .D(_0132_),
    .Q(\i_main_reg.data_d[99] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _1389_ (.RESET_B(net507),
    .D(net227),
    .Q(\i_main_reg.data_d[100] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _1390_ (.RESET_B(net507),
    .D(net280),
    .Q(\i_main_reg.data_d[101] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _1391_ (.RESET_B(net507),
    .D(net650),
    .Q(\i_main_reg.data_d[102] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1392_ (.RESET_B(net507),
    .D(net743),
    .Q(\i_main_reg.data_d[103] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _1393_ (.RESET_B(net507),
    .D(net589),
    .Q(\i_main_reg.data_d[104] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _1394_ (.RESET_B(net510),
    .D(net555),
    .Q(\i_main_reg.data_d[105] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1395_ (.RESET_B(net510),
    .D(_0139_),
    .Q(\i_main_reg.data_d[106] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1396_ (.RESET_B(net509),
    .D(_0140_),
    .Q(\i_main_reg.data_d[107] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1397_ (.RESET_B(net509),
    .D(_0141_),
    .Q(\i_main_reg.data_d[108] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1398_ (.RESET_B(net509),
    .D(net746),
    .Q(\i_main_reg.data_d[109] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1399_ (.RESET_B(net503),
    .D(net808),
    .Q(\i_main_reg.data_d[110] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1400_ (.RESET_B(net503),
    .D(net205),
    .Q(\i_main_reg.data_d[111] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1401_ (.RESET_B(net504),
    .D(_0145_),
    .Q(\i_main_reg.data_d[112] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1402_ (.RESET_B(net504),
    .D(net133),
    .Q(\i_main_reg.data_d[113] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1403_ (.RESET_B(net504),
    .D(_0147_),
    .Q(\i_main_reg.data_d[114] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1404_ (.RESET_B(net488),
    .D(net282),
    .Q(\i_main_reg.data_d[115] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1405_ (.RESET_B(net488),
    .D(net77),
    .Q(\i_main_reg.data_d[116] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1406_ (.RESET_B(net488),
    .D(_0150_),
    .Q(\i_main_reg.data_d[117] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1407_ (.RESET_B(net488),
    .D(_0151_),
    .Q(\i_main_reg.data_d[118] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _1408_ (.RESET_B(net487),
    .D(net192),
    .Q(\i_main_reg.data_d[119] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1409_ (.RESET_B(net487),
    .D(net801),
    .Q(\i_main_reg.data_d[120] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1410_ (.RESET_B(net485),
    .D(_0154_),
    .Q(\i_main_reg.data_d[121] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1411_ (.RESET_B(net486),
    .D(_0155_),
    .Q(\i_main_reg.data_d[122] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1412_ (.RESET_B(net481),
    .D(_0156_),
    .Q(\i_main_reg.data_d[123] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1413_ (.RESET_B(net481),
    .D(_0157_),
    .Q(\i_main_reg.data_d[124] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1414_ (.RESET_B(net481),
    .D(net595),
    .Q(\i_main_reg.data_d[125] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1415_ (.RESET_B(net482),
    .D(net656),
    .Q(\i_main_reg.data_d[126] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1416_ (.RESET_B(net483),
    .D(net63),
    .Q(\i_main_reg.data_d[127] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1417_ (.RESET_B(net483),
    .D(_0161_),
    .Q(\i_main_reg.data_d[128] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1418_ (.RESET_B(net483),
    .D(_0162_),
    .Q(\i_main_reg.data_d[129] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1419_ (.RESET_B(net469),
    .D(net256),
    .Q(\i_main_reg.data_d[130] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1420_ (.RESET_B(net470),
    .D(net258),
    .Q(\i_main_reg.data_d[131] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1421_ (.RESET_B(net470),
    .D(net629),
    .Q(\i_main_reg.data_d[132] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1422_ (.RESET_B(net468),
    .D(net723),
    .Q(\i_main_reg.data_d[133] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1423_ (.RESET_B(net468),
    .D(_0167_),
    .Q(\i_main_reg.data_d[134] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1424_ (.RESET_B(net468),
    .D(net798),
    .Q(\i_main_reg.data_d[135] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1425_ (.RESET_B(net464),
    .D(net145),
    .Q(\i_main_reg.data_d[136] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _1426_ (.RESET_B(net465),
    .D(_0170_),
    .Q(\i_main_reg.data_d[137] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1427_ (.RESET_B(net465),
    .D(_0171_),
    .Q(\i_main_reg.data_d[138] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1428_ (.RESET_B(net469),
    .D(net640),
    .Q(\i_main_reg.data_d[139] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1429_ (.RESET_B(net468),
    .D(_0173_),
    .Q(\i_main_reg.data_d[140] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1430_ (.RESET_B(net468),
    .D(net528),
    .Q(\i_main_reg.data_d[141] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _1431_ (.RESET_B(net475),
    .D(_0175_),
    .Q(\i_main_reg.data_d[142] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _1432_ (.RESET_B(net475),
    .D(_0176_),
    .Q(\i_main_reg.data_d[143] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _1433_ (.RESET_B(net475),
    .D(net117),
    .Q(\i_main_reg.data_d[144] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _1434_ (.RESET_B(net475),
    .D(net558),
    .Q(\i_main_reg.data_d[145] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _1435_ (.RESET_B(net475),
    .D(net314),
    .Q(\i_main_reg.data_d[146] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _1436_ (.RESET_B(net475),
    .D(_0180_),
    .Q(\i_main_reg.data_d[147] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _1437_ (.RESET_B(net476),
    .D(_0181_),
    .Q(\i_main_reg.data_d[148] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _1438_ (.RESET_B(net476),
    .D(net181),
    .Q(\i_main_reg.data_d[149] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _1439_ (.RESET_B(net476),
    .D(net713),
    .Q(\i_main_reg.data_d[150] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _1440_ (.RESET_B(net476),
    .D(_0184_),
    .Q(\i_main_reg.data_d[151] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _1441_ (.RESET_B(net476),
    .D(net730),
    .Q(\i_main_reg.data_d[152] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _1442_ (.RESET_B(net475),
    .D(net53),
    .Q(\i_main_reg.data_d[153] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _1443_ (.RESET_B(net475),
    .D(_0187_),
    .Q(\i_main_reg.data_d[154] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _1444_ (.RESET_B(net476),
    .D(_0188_),
    .Q(\i_main_reg.data_d[155] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _1445_ (.RESET_B(net476),
    .D(net158),
    .Q(\i_main_reg.data_d[156] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _1446_ (.RESET_B(net472),
    .D(net350),
    .Q(\i_main_reg.data_d[157] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _1447_ (.RESET_B(net472),
    .D(net344),
    .Q(\i_main_reg.data_d[158] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _1448_ (.RESET_B(net472),
    .D(_0192_),
    .Q(\i_main_reg.data_d[159] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _1449_ (.RESET_B(net472),
    .D(_0193_),
    .Q(\i_main_reg.data_d[160] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _1450_ (.RESET_B(net472),
    .D(net107),
    .Q(\i_main_reg.data_d[161] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _1451_ (.RESET_B(net471),
    .D(_0195_),
    .Q(\i_main_reg.data_d[162] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _1452_ (.RESET_B(net471),
    .D(net115),
    .Q(\i_main_reg.data_d[163] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _1453_ (.RESET_B(net471),
    .D(net572),
    .Q(\i_main_reg.data_d[164] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _1454_ (.RESET_B(net456),
    .D(net615),
    .Q(\i_main_reg.data_d[165] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _1455_ (.RESET_B(net456),
    .D(net803),
    .Q(\i_main_reg.data_d[166] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _1456_ (.RESET_B(net457),
    .D(net761),
    .Q(\i_main_reg.data_d[167] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _1457_ (.RESET_B(net456),
    .D(_0201_),
    .Q(\i_main_reg.data_d[168] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _1458_ (.RESET_B(net456),
    .D(_0202_),
    .Q(\i_main_reg.data_d[169] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _1459_ (.RESET_B(net456),
    .D(net772),
    .Q(\i_main_reg.data_d[170] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _1460_ (.RESET_B(net452),
    .D(net604),
    .Q(\i_main_reg.data_d[171] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _1461_ (.RESET_B(net452),
    .D(_0205_),
    .Q(\i_main_reg.data_d[172] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _1462_ (.RESET_B(net452),
    .D(_0206_),
    .Q(\i_main_reg.data_d[173] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _1463_ (.RESET_B(net452),
    .D(net102),
    .Q(\i_main_reg.data_d[174] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _1464_ (.RESET_B(net450),
    .D(_0208_),
    .Q(\i_main_reg.data_d[175] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _1465_ (.RESET_B(net450),
    .D(_0209_),
    .Q(\i_main_reg.data_d[176] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _1466_ (.RESET_B(net450),
    .D(_0210_),
    .Q(\i_main_reg.data_d[177] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _1467_ (.RESET_B(net451),
    .D(net143),
    .Q(\i_main_reg.data_d[178] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _1468_ (.RESET_B(net451),
    .D(_0212_),
    .Q(\i_main_reg.data_d[179] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _1469_ (.RESET_B(net451),
    .D(_0213_),
    .Q(\i_main_reg.data_d[180] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _1470_ (.RESET_B(net451),
    .D(net286),
    .Q(\i_main_reg.data_d[181] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _1471_ (.RESET_B(net450),
    .D(net778),
    .Q(\i_main_reg.data_d[182] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _1472_ (.RESET_B(net454),
    .D(net783),
    .Q(\i_main_reg.data_d[183] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _1473_ (.RESET_B(net454),
    .D(net819),
    .Q(\i_main_reg.data_d[184] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _1474_ (.RESET_B(net454),
    .D(net752),
    .Q(\i_main_reg.data_d[185] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _1475_ (.RESET_B(net454),
    .D(net341),
    .Q(\i_main_reg.data_d[186] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _1476_ (.RESET_B(net454),
    .D(_0220_),
    .Q(\i_main_reg.data_d[187] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _1477_ (.RESET_B(net454),
    .D(net183),
    .Q(\i_main_reg.data_d[188] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _1478_ (.RESET_B(net454),
    .D(_0222_),
    .Q(\i_main_reg.data_d[189] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _1479_ (.RESET_B(net453),
    .D(_0223_),
    .Q(\i_main_reg.data_d[190] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _1480_ (.RESET_B(net453),
    .D(net126),
    .Q(\i_main_reg.data_d[191] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _1481_ (.RESET_B(net453),
    .D(net201),
    .Q(\i_main_reg.data_d[192] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _1482_ (.RESET_B(net453),
    .D(_0226_),
    .Q(\i_main_reg.data_d[193] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _1483_ (.RESET_B(net453),
    .D(_0227_),
    .Q(\i_main_reg.data_d[194] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _1484_ (.RESET_B(net453),
    .D(_0228_),
    .Q(\i_main_reg.data_d[195] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _1485_ (.RESET_B(net453),
    .D(_0229_),
    .Q(\i_main_reg.data_d[196] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _1486_ (.RESET_B(net453),
    .D(net207),
    .Q(\i_main_reg.data_d[197] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _1487_ (.RESET_B(net455),
    .D(net718),
    .Q(\i_main_reg.data_d[198] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _1488_ (.RESET_B(net455),
    .D(net857),
    .Q(\i_main_reg.data_d[199] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _1489_ (.RESET_B(net455),
    .D(net260),
    .Q(\i_main_reg.data_d[200] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _1490_ (.RESET_B(net455),
    .D(net166),
    .Q(\i_main_reg.data_d[201] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _1491_ (.RESET_B(net455),
    .D(_0235_),
    .Q(\i_main_reg.data_d[202] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _1492_ (.RESET_B(net455),
    .D(_0236_),
    .Q(\i_main_reg.data_d[203] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _1493_ (.RESET_B(net459),
    .D(_0237_),
    .Q(\i_main_reg.data_d[204] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _1494_ (.RESET_B(net458),
    .D(net196),
    .Q(\i_main_reg.data_d[205] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _1495_ (.RESET_B(net459),
    .D(net543),
    .Q(\i_main_reg.data_d[206] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _1496_ (.RESET_B(net459),
    .D(_0240_),
    .Q(\i_main_reg.data_d[207] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _1497_ (.RESET_B(net459),
    .D(_0241_),
    .Q(\i_main_reg.data_d[208] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _1498_ (.RESET_B(net459),
    .D(net249),
    .Q(\i_main_reg.data_d[209] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _1499_ (.RESET_B(net459),
    .D(net332),
    .Q(\i_main_reg.data_d[210] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _1500_ (.RESET_B(net459),
    .D(net531),
    .Q(\i_main_reg.data_d[211] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _1501_ (.RESET_B(net473),
    .D(_0245_),
    .Q(\i_main_reg.data_d[212] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _1502_ (.RESET_B(net473),
    .D(net563),
    .Q(\i_main_reg.data_d[213] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _1503_ (.RESET_B(net473),
    .D(_0247_),
    .Q(\i_main_reg.data_d[214] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _1504_ (.RESET_B(net473),
    .D(_0248_),
    .Q(\i_main_reg.data_d[215] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _1505_ (.RESET_B(net473),
    .D(net634),
    .Q(\i_main_reg.data_d[216] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _1506_ (.RESET_B(net473),
    .D(net736),
    .Q(\i_main_reg.data_d[217] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _1507_ (.RESET_B(net474),
    .D(_0251_),
    .Q(\i_main_reg.data_d[218] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _1508_ (.RESET_B(net474),
    .D(_0252_),
    .Q(\i_main_reg.data_d[219] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _1509_ (.RESET_B(net477),
    .D(net190),
    .Q(\i_main_reg.data_d[220] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _1510_ (.RESET_B(net477),
    .D(net638),
    .Q(\i_main_reg.data_d[221] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _1511_ (.RESET_B(net477),
    .D(_0255_),
    .Q(\i_main_reg.data_d[222] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _1512_ (.RESET_B(net477),
    .D(_0256_),
    .Q(\i_main_reg.data_d[223] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _1513_ (.RESET_B(net477),
    .D(_0257_),
    .Q(\i_main_reg.data_d[224] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _1514_ (.RESET_B(net478),
    .D(_0258_),
    .Q(\i_main_reg.data_d[225] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _1515_ (.RESET_B(net478),
    .D(net79),
    .Q(\i_main_reg.data_d[226] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _1516_ (.RESET_B(net478),
    .D(net148),
    .Q(\i_main_reg.data_d[227] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _1517_ (.RESET_B(net477),
    .D(_0261_),
    .Q(\i_main_reg.data_d[228] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _1518_ (.RESET_B(net477),
    .D(_0262_),
    .Q(\i_main_reg.data_d[229] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _1519_ (.RESET_B(net477),
    .D(net551),
    .Q(\i_main_reg.data_d[230] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _1520_ (.RESET_B(net474),
    .D(net837),
    .Q(\i_main_reg.data_d[231] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _1521_ (.RESET_B(net474),
    .D(net817),
    .Q(\i_main_reg.data_d[232] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _1522_ (.RESET_B(net474),
    .D(_0266_),
    .Q(\i_main_reg.data_d[233] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _1523_ (.RESET_B(net473),
    .D(net765),
    .Q(\i_main_reg.data_d[234] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _1524_ (.RESET_B(net473),
    .D(_0268_),
    .Q(\i_main_reg.data_d[235] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _1525_ (.RESET_B(net460),
    .D(_0269_),
    .Q(\i_main_reg.data_d[236] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _1526_ (.RESET_B(net460),
    .D(net620),
    .Q(\i_main_reg.data_d[237] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _1527_ (.RESET_B(net460),
    .D(_0271_),
    .Q(\i_main_reg.data_d[238] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _1528_ (.RESET_B(net458),
    .D(_0272_),
    .Q(\i_main_reg.data_d[239] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _1529_ (.RESET_B(net458),
    .D(net540),
    .Q(\i_main_reg.data_d[240] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _1530_ (.RESET_B(net458),
    .D(net689),
    .Q(\i_main_reg.data_d[241] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _1531_ (.RESET_B(net458),
    .D(_0275_),
    .Q(\i_main_reg.data_d[242] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _1532_ (.RESET_B(net458),
    .D(_0276_),
    .Q(\i_main_reg.data_d[243] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _1533_ (.RESET_B(net458),
    .D(net238),
    .Q(\i_main_reg.data_d[244] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _1534_ (.RESET_B(net458),
    .D(net685),
    .Q(\i_main_reg.data_d[245] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _1535_ (.RESET_B(net456),
    .D(net741),
    .Q(\i_main_reg.data_d[246] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _1536_ (.RESET_B(net456),
    .D(_0280_),
    .Q(\i_main_reg.data_d[247] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _1537_ (.RESET_B(net456),
    .D(net711),
    .Q(\i_main_reg.data_d[248] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _1538_ (.RESET_B(net457),
    .D(_0282_),
    .Q(\i_main_reg.data_d[249] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _1539_ (.RESET_B(net457),
    .D(net707),
    .Q(\i_main_reg.data_d[250] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _1540_ (.RESET_B(net457),
    .D(net791),
    .Q(\i_main_reg.data_d[251] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _1541_ (.RESET_B(net471),
    .D(net636),
    .Q(\i_main_reg.data_d[252] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _1542_ (.RESET_B(net471),
    .D(_0286_),
    .Q(\i_main_reg.data_d[253] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _1543_ (.RESET_B(net471),
    .D(net668),
    .Q(\i_main_reg.data_d[254] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _1544_ (.RESET_B(net471),
    .D(net262),
    .Q(\i_main_reg.data_d[255] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _1545_ (.RESET_B(net471),
    .D(_0289_),
    .Q(\i_main_reg.data_d[256] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _1546_ (.RESET_B(net472),
    .D(_0290_),
    .Q(\i_main_reg.data_d[257] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _1547_ (.RESET_B(net464),
    .D(net121),
    .Q(\i_main_reg.data_d[258] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _1548_ (.RESET_B(net464),
    .D(_0292_),
    .Q(\i_main_reg.data_d[259] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _1549_ (.RESET_B(net464),
    .D(net71),
    .Q(\i_main_reg.data_d[260] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _1550_ (.RESET_B(net464),
    .D(net587),
    .Q(\i_main_reg.data_d[261] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _1551_ (.RESET_B(net464),
    .D(net823),
    .Q(\i_main_reg.data_d[262] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _1552_ (.RESET_B(net464),
    .D(net842),
    .Q(\i_main_reg.data_d[263] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _1553_ (.RESET_B(net446),
    .D(net774),
    .Q(\i_main_reg.data_d[264] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _1554_ (.RESET_B(net446),
    .D(_0298_),
    .Q(\i_main_reg.data_d[265] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _1555_ (.RESET_B(net446),
    .D(_0299_),
    .Q(\i_main_reg.data_d[266] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _1556_ (.RESET_B(net448),
    .D(net821),
    .Q(\i_main_reg.data_d[267] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _1557_ (.RESET_B(net446),
    .D(_0301_),
    .Q(\i_main_reg.data_d[268] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _1558_ (.RESET_B(net447),
    .D(net199),
    .Q(\i_main_reg.data_d[269] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _1559_ (.RESET_B(net447),
    .D(_0303_),
    .Q(\i_main_reg.data_d[270] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _1560_ (.RESET_B(net447),
    .D(_0304_),
    .Q(\i_main_reg.data_d[271] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _1561_ (.RESET_B(net447),
    .D(net69),
    .Q(\i_main_reg.data_d[272] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _1562_ (.RESET_B(net443),
    .D(net612),
    .Q(\i_main_reg.data_d[273] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _1563_ (.RESET_B(net452),
    .D(_0307_),
    .Q(\i_main_reg.data_d[274] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _1564_ (.RESET_B(net452),
    .D(_0308_),
    .Q(\i_main_reg.data_d[275] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _1565_ (.RESET_B(net461),
    .D(_0309_),
    .Q(\i_main_reg.data_d[276] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _1566_ (.RESET_B(net450),
    .D(_0310_),
    .Q(\i_main_reg.data_d[277] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _1567_ (.RESET_B(net450),
    .D(_0311_),
    .Q(\i_main_reg.data_d[278] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _1568_ (.RESET_B(net450),
    .D(_0312_),
    .Q(\i_main_reg.data_d[279] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _1569_ (.RESET_B(net450),
    .D(_0313_),
    .Q(\i_main_reg.data_d[280] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _1570_ (.RESET_B(net442),
    .D(net174),
    .Q(\i_main_reg.data_d[281] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _1571_ (.RESET_B(net442),
    .D(_0315_),
    .Q(\i_main_reg.data_d[282] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _1572_ (.RESET_B(net442),
    .D(net338),
    .Q(\i_main_reg.data_d[283] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _1573_ (.RESET_B(net442),
    .D(net55),
    .Q(\i_main_reg.data_d[284] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _1574_ (.RESET_B(net441),
    .D(_0318_),
    .Q(\i_main_reg.data_d[285] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _1575_ (.RESET_B(net442),
    .D(net244),
    .Q(\i_main_reg.data_d[286] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _1576_ (.RESET_B(net442),
    .D(net46),
    .Q(\i_main_reg.data_d[287] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _1577_ (.RESET_B(net441),
    .D(_0321_),
    .Q(\i_main_reg.data_d[288] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _1578_ (.RESET_B(net441),
    .D(_0322_),
    .Q(\i_main_reg.data_d[289] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _1579_ (.RESET_B(net441),
    .D(net253),
    .Q(\i_main_reg.data_d[290] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _1580_ (.RESET_B(net441),
    .D(_0324_),
    .Q(\i_main_reg.data_d[291] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _1581_ (.RESET_B(net441),
    .D(net251),
    .Q(\i_main_reg.data_d[292] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _1582_ (.RESET_B(net441),
    .D(_0326_),
    .Q(\i_main_reg.data_d[293] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _1583_ (.RESET_B(net438),
    .D(net680),
    .Q(\i_main_reg.data_d[294] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _1584_ (.RESET_B(net439),
    .D(net666),
    .Q(\i_main_reg.data_d[295] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _1585_ (.RESET_B(net441),
    .D(_0329_),
    .Q(\i_main_reg.data_d[296] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _1586_ (.RESET_B(net443),
    .D(_0330_),
    .Q(\i_main_reg.data_d[297] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _1587_ (.RESET_B(net443),
    .D(_0331_),
    .Q(\i_main_reg.data_d[298] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _1588_ (.RESET_B(net443),
    .D(_0332_),
    .Q(\i_main_reg.data_d[299] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _1589_ (.RESET_B(net443),
    .D(net522),
    .Q(\i_main_reg.data_d[300] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _1590_ (.RESET_B(net447),
    .D(net119),
    .Q(\i_main_reg.data_d[301] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _1591_ (.RESET_B(net447),
    .D(_0335_),
    .Q(\i_main_reg.data_d[302] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _1592_ (.RESET_B(net447),
    .D(_0336_),
    .Q(\i_main_reg.data_d[303] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _1593_ (.RESET_B(net447),
    .D(net632),
    .Q(\i_main_reg.data_d[304] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _1594_ (.RESET_B(net446),
    .D(_0338_),
    .Q(\i_main_reg.data_d[305] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _1595_ (.RESET_B(net446),
    .D(net721),
    .Q(\i_main_reg.data_d[306] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _1596_ (.RESET_B(net446),
    .D(net691),
    .Q(\i_main_reg.data_d[307] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _1597_ (.RESET_B(net446),
    .D(_0341_),
    .Q(\i_main_reg.data_d[308] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _1598_ (.RESET_B(net464),
    .D(_0342_),
    .Q(\i_main_reg.data_d[309] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _1599_ (.RESET_B(net462),
    .D(_0343_),
    .Q(\i_main_reg.data_d[310] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1600_ (.RESET_B(net462),
    .D(_0344_),
    .Q(\i_main_reg.data_d[311] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _1601_ (.RESET_B(net445),
    .D(net214),
    .Q(\i_main_reg.data_d[312] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _1602_ (.RESET_B(net445),
    .D(net203),
    .Q(\i_main_reg.data_d[313] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1603_ (.RESET_B(net445),
    .D(_0347_),
    .Q(\i_main_reg.data_d[314] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _1604_ (.RESET_B(net445),
    .D(net242),
    .Q(\i_main_reg.data_d[315] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1605_ (.RESET_B(net444),
    .D(net330),
    .Q(\i_main_reg.data_d[316] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1606_ (.RESET_B(net444),
    .D(_0350_),
    .Q(\i_main_reg.data_d[317] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _1607_ (.RESET_B(net444),
    .D(_0351_),
    .Q(\i_main_reg.data_d[318] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1608_ (.RESET_B(net444),
    .D(_0352_),
    .Q(\i_main_reg.data_d[319] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _1609_ (.RESET_B(net440),
    .D(_0353_),
    .Q(\i_main_reg.data_d[320] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _1610_ (.RESET_B(net440),
    .D(_0354_),
    .Q(\i_main_reg.data_d[321] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _1611_ (.RESET_B(net449),
    .D(_0355_),
    .Q(\i_main_reg.data_d[322] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _1612_ (.RESET_B(net439),
    .D(net548),
    .Q(\i_main_reg.data_d[323] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _1613_ (.RESET_B(net439),
    .D(_0357_),
    .Q(\i_main_reg.data_d[324] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _1614_ (.RESET_B(net439),
    .D(net750),
    .Q(\i_main_reg.data_d[325] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _1615_ (.RESET_B(net438),
    .D(net759),
    .Q(\i_main_reg.data_d[326] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _1616_ (.RESET_B(net438),
    .D(net701),
    .Q(\i_main_reg.data_d[327] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _1617_ (.RESET_B(net438),
    .D(net319),
    .Q(\i_main_reg.data_d[328] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _1618_ (.RESET_B(net438),
    .D(net298),
    .Q(\i_main_reg.data_d[329] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _1619_ (.RESET_B(net438),
    .D(_0363_),
    .Q(\i_main_reg.data_d[330] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _1620_ (.RESET_B(net438),
    .D(_0364_),
    .Q(\i_main_reg.data_d[331] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _1621_ (.RESET_B(net438),
    .D(net152),
    .Q(\i_main_reg.data_d[332] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _1622_ (.RESET_B(net440),
    .D(net322),
    .Q(\i_main_reg.data_d[333] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _1623_ (.RESET_B(net440),
    .D(net292),
    .Q(\i_main_reg.data_d[334] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _1624_ (.RESET_B(net440),
    .D(net109),
    .Q(\i_main_reg.data_d[335] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _1625_ (.RESET_B(net440),
    .D(_0369_),
    .Q(\i_main_reg.data_d[336] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _1626_ (.RESET_B(net444),
    .D(net111),
    .Q(\i_main_reg.data_d[337] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _1627_ (.RESET_B(net444),
    .D(_0371_),
    .Q(\i_main_reg.data_d[338] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _1628_ (.RESET_B(net444),
    .D(_0372_),
    .Q(\i_main_reg.data_d[339] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _1629_ (.RESET_B(net444),
    .D(net67),
    .Q(\i_main_reg.data_d[340] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1630_ (.RESET_B(net445),
    .D(_0374_),
    .Q(\i_main_reg.data_d[341] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1631_ (.RESET_B(net445),
    .D(_0375_),
    .Q(\i_main_reg.data_d[342] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1632_ (.RESET_B(net445),
    .D(_0376_),
    .Q(\i_main_reg.data_d[343] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1633_ (.RESET_B(net462),
    .D(_0377_),
    .Q(\i_main_reg.data_d[344] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _1634_ (.RESET_B(net462),
    .D(_0378_),
    .Q(\i_main_reg.data_d[345] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _1635_ (.RESET_B(net462),
    .D(_0379_),
    .Q(\i_main_reg.data_d[346] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _1636_ (.RESET_B(net462),
    .D(_0380_),
    .Q(\i_main_reg.data_d[347] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _1637_ (.RESET_B(net462),
    .D(net593),
    .Q(\i_main_reg.data_d[348] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _1638_ (.RESET_B(net462),
    .D(net284),
    .Q(\i_main_reg.data_d[349] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1639_ (.RESET_B(net463),
    .D(_0383_),
    .Q(\i_main_reg.data_d[350] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _1640_ (.RESET_B(net463),
    .D(net317),
    .Q(\i_main_reg.data_d[351] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _1641_ (.RESET_B(net463),
    .D(_0385_),
    .Q(\i_main_reg.data_d[352] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _1642_ (.RESET_B(net463),
    .D(net324),
    .Q(\i_main_reg.data_d[353] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _1643_ (.RESET_B(net463),
    .D(net170),
    .Q(\i_main_reg.data_d[354] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _1644_ (.RESET_B(net466),
    .D(_0388_),
    .Q(\i_main_reg.data_d[355] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1645_ (.RESET_B(net466),
    .D(net61),
    .Q(\i_main_reg.data_d[356] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1646_ (.RESET_B(net466),
    .D(_0390_),
    .Q(\i_main_reg.data_d[357] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1647_ (.RESET_B(net466),
    .D(net271),
    .Q(\i_main_reg.data_d[358] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1648_ (.RESET_B(net467),
    .D(_0392_),
    .Q(\i_main_reg.data_d[359] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1649_ (.RESET_B(net467),
    .D(net57),
    .Q(\i_main_reg.data_d[360] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1650_ (.RESET_B(net467),
    .D(_0394_),
    .Q(\i_main_reg.data_d[361] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1651_ (.RESET_B(net467),
    .D(_0395_),
    .Q(\i_main_reg.data_d[362] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1652_ (.RESET_B(net482),
    .D(_0396_),
    .Q(\i_main_reg.data_d[363] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1653_ (.RESET_B(net482),
    .D(net172),
    .Q(\i_main_reg.data_d[364] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1654_ (.RESET_B(net482),
    .D(_0398_),
    .Q(\i_main_reg.data_d[365] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1655_ (.RESET_B(net482),
    .D(net91),
    .Q(\i_main_reg.data_d[366] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1656_ (.RESET_B(net481),
    .D(_0400_),
    .Q(\i_main_reg.data_d[367] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1657_ (.RESET_B(net481),
    .D(net212),
    .Q(\i_main_reg.data_d[368] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1658_ (.RESET_B(net481),
    .D(net75),
    .Q(\i_main_reg.data_d[369] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1659_ (.RESET_B(net485),
    .D(_0403_),
    .Q(\i_main_reg.data_d[370] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1660_ (.RESET_B(net485),
    .D(_0404_),
    .Q(\i_main_reg.data_d[371] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1661_ (.RESET_B(net485),
    .D(_0405_),
    .Q(\i_main_reg.data_d[372] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1662_ (.RESET_B(net485),
    .D(net131),
    .Q(\i_main_reg.data_d[373] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1663_ (.RESET_B(net485),
    .D(_0407_),
    .Q(\i_main_reg.data_d[374] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1664_ (.RESET_B(net485),
    .D(_0408_),
    .Q(\i_main_reg.data_d[375] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1665_ (.RESET_B(net485),
    .D(net537),
    .Q(\i_main_reg.data_d[376] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1666_ (.RESET_B(net481),
    .D(net585),
    .Q(\i_main_reg.data_d[377] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1667_ (.RESET_B(net481),
    .D(net796),
    .Q(\i_main_reg.data_d[378] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1668_ (.RESET_B(net484),
    .D(net326),
    .Q(\i_main_reg.data_d[379] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1669_ (.RESET_B(net482),
    .D(net83),
    .Q(\i_main_reg.data_d[380] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1670_ (.RESET_B(net482),
    .D(_0414_),
    .Q(\i_main_reg.data_d[381] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1671_ (.RESET_B(net482),
    .D(_0415_),
    .Q(\i_main_reg.data_d[382] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1672_ (.RESET_B(net467),
    .D(net160),
    .Q(\i_main_reg.data_d[383] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1673_ (.RESET_B(net467),
    .D(net163),
    .Q(\i_main_reg.data_d[384] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1674_ (.RESET_B(net466),
    .D(_0418_),
    .Q(\i_main_reg.data_d[385] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1675_ (.RESET_B(net467),
    .D(_0419_),
    .Q(\i_main_reg.data_d[386] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1676_ (.RESET_B(net466),
    .D(net65),
    .Q(\i_main_reg.data_d[387] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1677_ (.RESET_B(net466),
    .D(_0421_),
    .Q(\i_main_reg.data_d[388] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1678_ (.RESET_B(net466),
    .D(_0422_),
    .Q(\i_main_reg.data_d[389] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1679_ (.RESET_B(net463),
    .D(_0423_),
    .Q(\i_main_reg.data_d[390] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1680_ (.RESET_B(net463),
    .D(net525),
    .Q(\i_main_reg.data_d[391] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1681_ (.RESET_B(net468),
    .D(net574),
    .Q(\i_main_reg.data_d[392] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1682_ (.RESET_B(net468),
    .D(_0426_),
    .Q(\i_main_reg.data_d[393] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1683_ (.RESET_B(net468),
    .D(_0427_),
    .Q(\i_main_reg.data_d[394] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1684_ (.RESET_B(net469),
    .D(net627),
    .Q(\i_main_reg.data_d[395] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1685_ (.RESET_B(net469),
    .D(net51),
    .Q(\i_main_reg.data_d[396] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1686_ (.RESET_B(net469),
    .D(_0430_),
    .Q(\i_main_reg.data_d[397] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1687_ (.RESET_B(net469),
    .D(_0431_),
    .Q(\i_main_reg.data_d[398] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1688_ (.RESET_B(net469),
    .D(net141),
    .Q(\i_main_reg.data_d[399] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1689_ (.RESET_B(net483),
    .D(_0433_),
    .Q(\i_main_reg.data_d[400] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1690_ (.RESET_B(net483),
    .D(_0434_),
    .Q(\i_main_reg.data_d[401] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1691_ (.RESET_B(net483),
    .D(_0435_),
    .Q(\i_main_reg.data_d[402] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1692_ (.RESET_B(net483),
    .D(net246),
    .Q(\i_main_reg.data_d[403] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1693_ (.RESET_B(net483),
    .D(net781),
    .Q(\i_main_reg.data_d[404] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1694_ (.RESET_B(net484),
    .D(net811),
    .Q(\i_main_reg.data_d[405] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1695_ (.RESET_B(net484),
    .D(_0439_),
    .Q(\i_main_reg.data_d[406] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1696_ (.RESET_B(net484),
    .D(_0440_),
    .Q(\i_main_reg.data_d[407] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1697_ (.RESET_B(net487),
    .D(net229),
    .Q(\i_main_reg.data_d[408] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1698_ (.RESET_B(net487),
    .D(_0442_),
    .Q(\i_main_reg.data_d[409] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1699_ (.RESET_B(net487),
    .D(net221),
    .Q(\i_main_reg.data_d[410] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1700_ (.RESET_B(net487),
    .D(net660),
    .Q(\i_main_reg.data_d[411] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1701_ (.RESET_B(net487),
    .D(_0445_),
    .Q(\i_main_reg.data_d[412] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1702_ (.RESET_B(net487),
    .D(_0446_),
    .Q(\i_main_reg.data_d[413] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1703_ (.RESET_B(net488),
    .D(net277),
    .Q(\i_main_reg.data_d[414] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1704_ (.RESET_B(net494),
    .D(net288),
    .Q(\i_main_reg.data_d[415] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _1705_ (.RESET_B(net490),
    .D(_0449_),
    .Q(\i_main_reg.data_d[416] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1706_ (.RESET_B(net490),
    .D(_0450_),
    .Q(\i_main_reg.data_d[417] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1707_ (.RESET_B(net490),
    .D(_0451_),
    .Q(\i_main_reg.data_d[418] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1708_ (.RESET_B(net490),
    .D(_0452_),
    .Q(\i_main_reg.data_d[419] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1709_ (.RESET_B(net490),
    .D(_0453_),
    .Q(\i_main_reg.data_d[420] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1710_ (.RESET_B(net489),
    .D(net73),
    .Q(\i_main_reg.data_d[421] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1711_ (.RESET_B(net489),
    .D(net618),
    .Q(\i_main_reg.data_d[422] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1712_ (.RESET_B(net489),
    .D(net748),
    .Q(\i_main_reg.data_d[423] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1713_ (.RESET_B(net489),
    .D(net578),
    .Q(\i_main_reg.data_d[424] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1714_ (.RESET_B(net489),
    .D(_0458_),
    .Q(\i_main_reg.data_d[425] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1715_ (.RESET_B(net489),
    .D(net129),
    .Q(\i_main_reg.data_d[426] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _1716_ (.RESET_B(net489),
    .D(net336),
    .Q(\i_main_reg.data_d[427] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _1717_ (.RESET_B(net491),
    .D(_0461_),
    .Q(\i_main_reg.data_d[428] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1718_ (.RESET_B(net491),
    .D(_0462_),
    .Q(\i_main_reg.data_d[429] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1719_ (.RESET_B(net491),
    .D(_0463_),
    .Q(\i_main_reg.data_d[430] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1720_ (.RESET_B(net493),
    .D(_0464_),
    .Q(\i_main_reg.data_d[431] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _1721_ (.RESET_B(net499),
    .D(_0465_),
    .Q(\i_main_reg.data_d[432] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _1722_ (.RESET_B(net493),
    .D(net97),
    .Q(\i_main_reg.data_d[433] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _1723_ (.RESET_B(net496),
    .D(_0467_),
    .Q(\i_main_reg.data_d[434] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _1724_ (.RESET_B(net496),
    .D(_0468_),
    .Q(\i_main_reg.data_d[435] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _1725_ (.RESET_B(net496),
    .D(net534),
    .Q(\i_main_reg.data_d[436] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _1726_ (.RESET_B(net496),
    .D(net93),
    .Q(\i_main_reg.data_d[437] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _1727_ (.RESET_B(net497),
    .D(_0471_),
    .Q(\i_main_reg.data_d[438] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _1728_ (.RESET_B(net497),
    .D(net139),
    .Q(\i_main_reg.data_d[439] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _1729_ (.RESET_B(net497),
    .D(_0473_),
    .Q(\i_main_reg.data_d[440] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _1730_ (.RESET_B(net497),
    .D(_0474_),
    .Q(\i_main_reg.data_d[441] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _1731_ (.RESET_B(net512),
    .D(_0475_),
    .Q(\i_main_reg.data_d[442] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _1732_ (.RESET_B(net512),
    .D(_0476_),
    .Q(\i_main_reg.data_d[443] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _1733_ (.RESET_B(net512),
    .D(net290),
    .Q(\i_main_reg.data_d[444] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _1734_ (.RESET_B(net513),
    .D(_0478_),
    .Q(\i_main_reg.data_d[445] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _1735_ (.RESET_B(net513),
    .D(net36),
    .Q(\i_main_reg.data_d[446] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _1736_ (.RESET_B(net517),
    .D(net34),
    .Q(\one_count_q[0] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _1737_ (.RESET_B(net517),
    .D(net346),
    .Q(\one_count_q[1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_6 (.L_LO(net6));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_7 (.L_LO(net7));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_8 (.L_LO(net8));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_9 (.L_LO(net9));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_10 (.L_LO(net10));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_11 (.L_LO(net11));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_12 (.L_LO(net12));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_13 (.L_LO(net13));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_14 (.L_LO(net14));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_15 (.L_LO(net15));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_16 (.L_LO(net16));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_17 (.L_LO(net17));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_18 (.L_LO(net18));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_19 (.L_LO(net19));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_20 (.L_LO(net20));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_21 (.L_LO(net21));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_22 (.L_LO(net22));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_23 (.L_LO(net23));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_24 (.L_LO(net24));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _1758_ (.A(\i_main_reg.data_o ),
    .X(uo_out[0]));
 sg13g2_buf_1 _1759_ (.A(\i_step_counter.data_o ),
    .X(uo_out[1]));
 sg13g2_buf_1 _1760_ (.A(finished_q),
    .X(uo_out[2]));
 sg13g2_buf_1 _1761_ (.A(overflow_q),
    .X(uo_out[3]));
 sg13g2_buf_8 fanout352 (.A(_0488_),
    .X(net352));
 sg13g2_buf_8 fanout353 (.A(_0487_),
    .X(net353));
 sg13g2_buf_8 fanout354 (.A(_0485_),
    .X(net354));
 sg13g2_buf_8 fanout355 (.A(net357),
    .X(net355));
 sg13g2_buf_1 fanout356 (.A(net357),
    .X(net356));
 sg13g2_buf_8 fanout357 (.A(net377),
    .X(net357));
 sg13g2_buf_8 fanout358 (.A(net360),
    .X(net358));
 sg13g2_buf_8 fanout359 (.A(net360),
    .X(net359));
 sg13g2_buf_8 fanout360 (.A(net377),
    .X(net360));
 sg13g2_buf_8 fanout361 (.A(net365),
    .X(net361));
 sg13g2_buf_8 fanout362 (.A(net365),
    .X(net362));
 sg13g2_buf_8 fanout363 (.A(net365),
    .X(net363));
 sg13g2_buf_8 fanout364 (.A(net365),
    .X(net364));
 sg13g2_buf_8 fanout365 (.A(net377),
    .X(net365));
 sg13g2_buf_8 fanout366 (.A(net368),
    .X(net366));
 sg13g2_buf_1 fanout367 (.A(net368),
    .X(net367));
 sg13g2_buf_8 fanout368 (.A(net377),
    .X(net368));
 sg13g2_buf_8 fanout369 (.A(net371),
    .X(net369));
 sg13g2_buf_8 fanout370 (.A(net371),
    .X(net370));
 sg13g2_buf_8 fanout371 (.A(net377),
    .X(net371));
 sg13g2_buf_8 fanout372 (.A(net376),
    .X(net372));
 sg13g2_buf_1 fanout373 (.A(net376),
    .X(net373));
 sg13g2_buf_8 fanout374 (.A(net375),
    .X(net374));
 sg13g2_buf_8 fanout375 (.A(net376),
    .X(net375));
 sg13g2_buf_8 fanout376 (.A(net377),
    .X(net376));
 sg13g2_buf_8 fanout377 (.A(_0581_),
    .X(net377));
 sg13g2_buf_8 fanout378 (.A(net380),
    .X(net378));
 sg13g2_buf_1 fanout379 (.A(net380),
    .X(net379));
 sg13g2_buf_8 fanout380 (.A(net397),
    .X(net380));
 sg13g2_buf_8 fanout381 (.A(net386),
    .X(net381));
 sg13g2_buf_8 fanout382 (.A(net386),
    .X(net382));
 sg13g2_buf_8 fanout383 (.A(net385),
    .X(net383));
 sg13g2_buf_1 fanout384 (.A(net385),
    .X(net384));
 sg13g2_buf_8 fanout385 (.A(net386),
    .X(net385));
 sg13g2_buf_8 fanout386 (.A(net397),
    .X(net386));
 sg13g2_buf_8 fanout387 (.A(net391),
    .X(net387));
 sg13g2_buf_8 fanout388 (.A(net391),
    .X(net388));
 sg13g2_buf_8 fanout389 (.A(net391),
    .X(net389));
 sg13g2_buf_8 fanout390 (.A(net391),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(net396),
    .X(net391));
 sg13g2_buf_8 fanout392 (.A(net393),
    .X(net392));
 sg13g2_buf_8 fanout393 (.A(net396),
    .X(net393));
 sg13g2_buf_8 fanout394 (.A(net395),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(net396),
    .X(net395));
 sg13g2_buf_1 fanout396 (.A(net397),
    .X(net396));
 sg13g2_buf_8 fanout397 (.A(_0581_),
    .X(net397));
 sg13g2_buf_8 fanout398 (.A(net399),
    .X(net398));
 sg13g2_buf_8 fanout399 (.A(net406),
    .X(net399));
 sg13g2_buf_8 fanout400 (.A(net406),
    .X(net400));
 sg13g2_buf_8 fanout401 (.A(net406),
    .X(net401));
 sg13g2_buf_8 fanout402 (.A(net403),
    .X(net402));
 sg13g2_buf_8 fanout403 (.A(net406),
    .X(net403));
 sg13g2_buf_8 fanout404 (.A(net406),
    .X(net404));
 sg13g2_buf_1 fanout405 (.A(net406),
    .X(net405));
 sg13g2_buf_8 fanout406 (.A(net432),
    .X(net406));
 sg13g2_buf_8 fanout407 (.A(net408),
    .X(net407));
 sg13g2_buf_8 fanout408 (.A(net411),
    .X(net408));
 sg13g2_buf_8 fanout409 (.A(net410),
    .X(net409));
 sg13g2_buf_8 fanout410 (.A(net411),
    .X(net410));
 sg13g2_buf_8 fanout411 (.A(net432),
    .X(net411));
 sg13g2_buf_8 fanout412 (.A(net416),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(net416),
    .X(net413));
 sg13g2_buf_8 fanout414 (.A(net416),
    .X(net414));
 sg13g2_buf_8 fanout415 (.A(net416),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(net432),
    .X(net416));
 sg13g2_buf_8 fanout417 (.A(net419),
    .X(net417));
 sg13g2_buf_8 fanout418 (.A(net419),
    .X(net418));
 sg13g2_buf_8 fanout419 (.A(net428),
    .X(net419));
 sg13g2_buf_8 fanout420 (.A(net428),
    .X(net420));
 sg13g2_buf_8 fanout421 (.A(net428),
    .X(net421));
 sg13g2_buf_8 fanout422 (.A(net423),
    .X(net422));
 sg13g2_buf_8 fanout423 (.A(net424),
    .X(net423));
 sg13g2_buf_8 fanout424 (.A(net428),
    .X(net424));
 sg13g2_buf_8 fanout425 (.A(net427),
    .X(net425));
 sg13g2_buf_8 fanout426 (.A(net427),
    .X(net426));
 sg13g2_buf_8 fanout427 (.A(net428),
    .X(net427));
 sg13g2_buf_8 fanout428 (.A(net431),
    .X(net428));
 sg13g2_buf_8 fanout429 (.A(net430),
    .X(net429));
 sg13g2_buf_8 fanout430 (.A(net431),
    .X(net430));
 sg13g2_buf_8 fanout431 (.A(net432),
    .X(net431));
 sg13g2_buf_8 fanout432 (.A(_0581_),
    .X(net432));
 sg13g2_buf_8 fanout433 (.A(net434),
    .X(net433));
 sg13g2_buf_8 fanout434 (.A(_0608_),
    .X(net434));
 sg13g2_buf_8 fanout435 (.A(\i_main_reg.data_o ),
    .X(net435));
 sg13g2_buf_8 fanout436 (.A(net437),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(\state_q[1] ),
    .X(net437));
 sg13g2_buf_8 fanout438 (.A(net440),
    .X(net438));
 sg13g2_buf_1 fanout439 (.A(net440),
    .X(net439));
 sg13g2_buf_8 fanout440 (.A(net449),
    .X(net440));
 sg13g2_buf_8 fanout441 (.A(net443),
    .X(net441));
 sg13g2_buf_8 fanout442 (.A(net443),
    .X(net442));
 sg13g2_buf_8 fanout443 (.A(net449),
    .X(net443));
 sg13g2_buf_8 fanout444 (.A(net448),
    .X(net444));
 sg13g2_buf_8 fanout445 (.A(net448),
    .X(net445));
 sg13g2_buf_8 fanout446 (.A(net448),
    .X(net446));
 sg13g2_buf_8 fanout447 (.A(net448),
    .X(net447));
 sg13g2_buf_8 fanout448 (.A(net449),
    .X(net448));
 sg13g2_buf_8 fanout449 (.A(net480),
    .X(net449));
 sg13g2_buf_8 fanout450 (.A(net452),
    .X(net450));
 sg13g2_buf_1 fanout451 (.A(net452),
    .X(net451));
 sg13g2_buf_8 fanout452 (.A(net461),
    .X(net452));
 sg13g2_buf_8 fanout453 (.A(net454),
    .X(net453));
 sg13g2_buf_8 fanout454 (.A(net455),
    .X(net454));
 sg13g2_buf_8 fanout455 (.A(net461),
    .X(net455));
 sg13g2_buf_8 fanout456 (.A(net460),
    .X(net456));
 sg13g2_buf_1 fanout457 (.A(net460),
    .X(net457));
 sg13g2_buf_8 fanout458 (.A(net459),
    .X(net458));
 sg13g2_buf_8 fanout459 (.A(net460),
    .X(net459));
 sg13g2_buf_8 fanout460 (.A(net461),
    .X(net460));
 sg13g2_buf_8 fanout461 (.A(net480),
    .X(net461));
 sg13g2_buf_8 fanout462 (.A(net465),
    .X(net462));
 sg13g2_buf_8 fanout463 (.A(net465),
    .X(net463));
 sg13g2_buf_8 fanout464 (.A(net465),
    .X(net464));
 sg13g2_buf_8 fanout465 (.A(net480),
    .X(net465));
 sg13g2_buf_8 fanout466 (.A(net470),
    .X(net466));
 sg13g2_buf_8 fanout467 (.A(net470),
    .X(net467));
 sg13g2_buf_8 fanout468 (.A(net469),
    .X(net468));
 sg13g2_buf_8 fanout469 (.A(net470),
    .X(net469));
 sg13g2_buf_8 fanout470 (.A(net480),
    .X(net470));
 sg13g2_buf_8 fanout471 (.A(net472),
    .X(net471));
 sg13g2_buf_8 fanout472 (.A(net479),
    .X(net472));
 sg13g2_buf_8 fanout473 (.A(net479),
    .X(net473));
 sg13g2_buf_8 fanout474 (.A(net479),
    .X(net474));
 sg13g2_buf_8 fanout475 (.A(net476),
    .X(net475));
 sg13g2_buf_8 fanout476 (.A(net479),
    .X(net476));
 sg13g2_buf_8 fanout477 (.A(net478),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(net479),
    .X(net478));
 sg13g2_buf_8 fanout479 (.A(net480),
    .X(net479));
 sg13g2_buf_8 fanout480 (.A(rst_n),
    .X(net480));
 sg13g2_buf_8 fanout481 (.A(net484),
    .X(net481));
 sg13g2_buf_8 fanout482 (.A(net484),
    .X(net482));
 sg13g2_buf_8 fanout483 (.A(net484),
    .X(net483));
 sg13g2_buf_8 fanout484 (.A(net500),
    .X(net484));
 sg13g2_buf_8 fanout485 (.A(net486),
    .X(net485));
 sg13g2_buf_8 fanout486 (.A(net500),
    .X(net486));
 sg13g2_buf_8 fanout487 (.A(net488),
    .X(net487));
 sg13g2_buf_8 fanout488 (.A(net500),
    .X(net488));
 sg13g2_buf_8 fanout489 (.A(net491),
    .X(net489));
 sg13g2_buf_8 fanout490 (.A(net491),
    .X(net490));
 sg13g2_buf_8 fanout491 (.A(net499),
    .X(net491));
 sg13g2_buf_8 fanout492 (.A(net493),
    .X(net492));
 sg13g2_buf_8 fanout493 (.A(net499),
    .X(net493));
 sg13g2_buf_8 fanout494 (.A(net498),
    .X(net494));
 sg13g2_buf_8 fanout495 (.A(net498),
    .X(net495));
 sg13g2_buf_8 fanout496 (.A(net498),
    .X(net496));
 sg13g2_buf_8 fanout497 (.A(net498),
    .X(net497));
 sg13g2_buf_8 fanout498 (.A(net499),
    .X(net498));
 sg13g2_buf_8 fanout499 (.A(net500),
    .X(net499));
 sg13g2_buf_8 fanout500 (.A(net519),
    .X(net500));
 sg13g2_buf_8 fanout501 (.A(net505),
    .X(net501));
 sg13g2_buf_8 fanout502 (.A(net505),
    .X(net502));
 sg13g2_buf_8 fanout503 (.A(net505),
    .X(net503));
 sg13g2_buf_8 fanout504 (.A(net505),
    .X(net504));
 sg13g2_buf_8 fanout505 (.A(net511),
    .X(net505));
 sg13g2_buf_8 fanout506 (.A(net508),
    .X(net506));
 sg13g2_buf_8 fanout507 (.A(net508),
    .X(net507));
 sg13g2_buf_8 fanout508 (.A(net511),
    .X(net508));
 sg13g2_buf_8 fanout509 (.A(net510),
    .X(net509));
 sg13g2_buf_8 fanout510 (.A(net511),
    .X(net510));
 sg13g2_buf_8 fanout511 (.A(net519),
    .X(net511));
 sg13g2_buf_8 fanout512 (.A(net513),
    .X(net512));
 sg13g2_buf_8 fanout513 (.A(net519),
    .X(net513));
 sg13g2_buf_8 fanout514 (.A(net518),
    .X(net514));
 sg13g2_buf_8 fanout515 (.A(net518),
    .X(net515));
 sg13g2_buf_8 fanout516 (.A(net517),
    .X(net516));
 sg13g2_buf_8 fanout517 (.A(net518),
    .X(net517));
 sg13g2_buf_8 fanout518 (.A(net519),
    .X(net518));
 sg13g2_buf_8 fanout519 (.A(rst_n),
    .X(net519));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_5 (.L_LO(net5));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_4_7_0_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_4_11_0_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_4_15_0_clk));
 sg13g2_inv_8 clkload3 (.A(clknet_leaf_15_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\bit_counter_q[1] ),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0564_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold3 (.A(overflow_q),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0017_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold5 (.A(\bit_counter_q[0] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0020_),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold7 (.A(\bit_counter_q[2] ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0022_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold9 (.A(\one_count_q[0] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0480_),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold11 (.A(\i_main_reg.data_d[446] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0479_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold13 (.A(\i_main_reg.data_d[0] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0583_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold15 (.A(\bit_counter_q[6] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0574_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold17 (.A(\i_step_counter.data_d[6] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0006_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold19 (.A(\i_step_counter.data_d[10] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0010_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold21 (.A(\i_main_reg.data_d[288] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0320_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold23 (.A(\bit_counter_q[8] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0578_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0028_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold26 (.A(\i_main_reg.data_d[397] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0429_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold28 (.A(\i_main_reg.data_d[154] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0186_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold30 (.A(\i_main_reg.data_d[285] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0317_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold32 (.A(\i_main_reg.data_d[361] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0393_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold34 (.A(\i_step_counter.data_d[4] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0004_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold36 (.A(\i_main_reg.data_d[357] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0389_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold38 (.A(\i_main_reg.data_d[128] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0160_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold40 (.A(\i_main_reg.data_d[387] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0420_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold42 (.A(\i_main_reg.data_d[341] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0373_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold44 (.A(\i_main_reg.data_d[272] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0305_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold46 (.A(\i_main_reg.data_d[260] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0293_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold48 (.A(\i_main_reg.data_d[421] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0454_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold50 (.A(\i_main_reg.data_d[370] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0402_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold52 (.A(\i_main_reg.data_d[117] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0149_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold54 (.A(\i_main_reg.data_d[226] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0259_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold56 (.A(\i_main_reg.data_d[14] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0047_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold58 (.A(\i_main_reg.data_d[381] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0413_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold60 (.A(\i_main_reg.data_d[56] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0089_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold62 (.A(\i_main_reg.data_d[74] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0106_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold64 (.A(\i_main_reg.data_d[1] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0034_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold66 (.A(\i_main_reg.data_d[366] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0399_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold68 (.A(\i_main_reg.data_d[438] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0470_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold70 (.A(\i_main_reg.data_d[97] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0130_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold72 (.A(\i_main_reg.data_d[433] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0466_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold74 (.A(finished_q),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0016_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold76 (.A(\i_main_reg.data_d[96] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold77 (.A(\i_main_reg.data_d[174] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0207_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold79 (.A(\i_main_reg.data_d[13] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0045_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold81 (.A(\i_main_reg.data_d[225] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold82 (.A(\i_main_reg.data_d[161] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0194_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold84 (.A(\i_main_reg.data_d[336] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0368_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold86 (.A(\i_main_reg.data_d[338] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0370_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold88 (.A(\i_main_reg.data_d[155] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold89 (.A(\i_main_reg.data_d[118] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold90 (.A(\i_main_reg.data_d[163] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0196_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold92 (.A(\i_main_reg.data_d[144] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0177_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold94 (.A(\i_main_reg.data_d[302] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0334_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold96 (.A(\i_main_reg.data_d[258] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0291_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold98 (.A(\i_main_reg.data_d[95] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold99 (.A(\i_main_reg.data_d[39] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0071_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold101 (.A(\i_main_reg.data_d[191] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0224_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold103 (.A(\i_main_reg.data_d[224] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold104 (.A(\i_main_reg.data_d[426] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0459_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold106 (.A(\i_main_reg.data_d[373] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0406_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold108 (.A(\i_main_reg.data_d[114] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0146_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold110 (.A(\i_main_reg.data_d[129] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold111 (.A(\i_main_reg.data_d[98] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0131_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold113 (.A(\i_main_reg.data_d[342] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold114 (.A(\i_main_reg.data_d[440] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0472_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold116 (.A(\i_main_reg.data_d[399] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0432_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold118 (.A(\i_main_reg.data_d[178] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0211_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold120 (.A(\i_main_reg.data_d[137] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0169_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold122 (.A(\i_main_reg.data_d[55] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold123 (.A(\i_main_reg.data_d[228] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0260_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold125 (.A(\i_main_reg.data_d[33] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0065_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold127 (.A(\i_main_reg.data_d[332] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0365_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold129 (.A(\i_main_reg.data_d[93] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0125_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold131 (.A(\i_main_reg.data_d[43] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0075_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold133 (.A(\i_main_reg.data_d[156] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0189_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold135 (.A(\i_main_reg.data_d[383] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0416_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold137 (.A(\i_main_reg.data_d[420] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold138 (.A(\i_main_reg.data_d[384] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0417_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold140 (.A(\i_main_reg.data_d[398] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold141 (.A(\i_main_reg.data_d[202] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0234_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold143 (.A(\i_main_reg.data_d[432] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold144 (.A(\i_main_reg.data_d[162] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold145 (.A(\i_main_reg.data_d[355] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0387_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold147 (.A(\i_main_reg.data_d[364] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0397_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold149 (.A(\i_main_reg.data_d[281] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0314_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold151 (.A(\i_main_reg.data_d[15] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0048_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold153 (.A(\i_main_reg.data_d[372] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold154 (.A(\i_main_reg.data_d[362] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold155 (.A(\i_main_reg.data_d[382] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold156 (.A(\i_main_reg.data_d[149] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0182_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold158 (.A(\i_main_reg.data_d[189] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0221_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold160 (.A(\i_main_reg.data_d[19] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0052_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold162 (.A(\i_main_reg.data_d[148] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold163 (.A(\i_main_reg.data_d[303] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold164 (.A(\i_main_reg.data_d[289] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold165 (.A(\i_main_reg.data_d[220] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0253_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold167 (.A(\i_main_reg.data_d[119] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0152_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold169 (.A(\i_main_reg.data_d[339] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold170 (.A(\i_main_reg.data_d[229] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold171 (.A(\i_main_reg.data_d[205] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0238_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold173 (.A(\i_main_reg.data_d[441] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold174 (.A(\i_main_reg.data_d[270] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0302_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold176 (.A(\i_main_reg.data_d[193] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0225_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold178 (.A(\i_main_reg.data_d[314] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0346_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold180 (.A(\i_main_reg.data_d[112] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0144_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold182 (.A(\i_main_reg.data_d[197] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0230_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold184 (.A(\i_main_reg.data_d[371] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold185 (.A(\i_main_reg.data_d[177] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold186 (.A(\i_main_reg.data_d[271] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold187 (.A(\i_main_reg.data_d[368] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0401_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold189 (.A(\i_main_reg.data_d[312] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0345_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold191 (.A(\i_main_reg.data_d[40] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold192 (.A(\i_main_reg.data_d[27] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0060_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold194 (.A(\i_main_reg.data_d[44] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold195 (.A(\i_main_reg.data_d[113] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold196 (.A(\i_main_reg.data_d[410] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0443_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold198 (.A(\i_main_reg.data_d[91] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0124_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold200 (.A(\i_main_reg.data_d[196] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold201 (.A(\i_main_reg.data_d[259] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold202 (.A(\i_main_reg.data_d[100] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0133_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold204 (.A(\i_main_reg.data_d[409] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0441_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold206 (.A(\i_main_reg.data_d[21] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0053_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold208 (.A(\i_main_reg.data_d[138] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold209 (.A(\i_main_reg.data_d[94] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold210 (.A(\i_main_reg.data_d[29] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0062_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold212 (.A(\i_main_reg.data_d[194] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold213 (.A(\i_main_reg.data_d[244] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0277_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold215 (.A(\i_main_reg.data_d[356] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold216 (.A(\i_main_reg.data_d[311] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold217 (.A(\i_main_reg.data_d[315] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0348_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold219 (.A(\i_main_reg.data_d[287] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0319_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold221 (.A(\i_main_reg.data_d[403] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0436_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold223 (.A(\i_main_reg.data_d[286] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold224 (.A(\i_main_reg.data_d[209] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0242_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold226 (.A(\i_main_reg.data_d[292] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0325_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold228 (.A(\i_main_reg.data_d[290] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0323_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold230 (.A(\i_main_reg.data_d[28] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold231 (.A(\i_main_reg.data_d[130] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0163_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold233 (.A(\i_main_reg.data_d[131] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0164_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold235 (.A(\i_main_reg.data_d[201] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0233_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold237 (.A(\i_main_reg.data_d[256] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0288_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold239 (.A(\i_main_reg.data_d[99] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold240 (.A(\i_main_reg.data_d[204] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold241 (.A(\i_main_reg.data_d[23] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0056_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold243 (.A(\i_main_reg.data_d[208] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold244 (.A(\i_main_reg.data_d[60] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0092_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold246 (.A(\i_main_reg.data_d[359] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0391_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold248 (.A(\i_main_reg.data_d[195] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold249 (.A(\i_main_reg.data_d[360] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold250 (.A(\i_main_reg.data_d[6] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0038_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold252 (.A(\i_main_reg.data_d[414] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0447_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold254 (.A(\i_main_reg.data_d[365] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold255 (.A(\i_main_reg.data_d[101] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0134_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold257 (.A(\i_main_reg.data_d[115] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0148_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold259 (.A(\i_main_reg.data_d[350] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0382_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold261 (.A(\i_main_reg.data_d[181] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0214_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold263 (.A(\i_main_reg.data_d[416] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0448_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold265 (.A(\i_main_reg.data_d[444] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0477_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold267 (.A(\i_main_reg.data_d[335] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0367_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold269 (.A(\i_main_reg.data_d[47] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0079_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold271 (.A(\i_main_reg.data_d[291] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold272 (.A(\i_main_reg.data_d[257] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold273 (.A(\i_main_reg.data_d[330] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold274 (.A(_0362_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold275 (.A(\i_main_reg.data_d[280] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold276 (.A(\i_main_reg.data_d[431] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold277 (.A(\i_main_reg.data_d[363] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold278 (.A(\i_main_reg.data_d[439] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold279 (.A(\i_main_reg.data_d[180] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold280 (.A(\i_main_reg.data_d[11] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold281 (.A(_0044_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold282 (.A(\i_main_reg.data_d[367] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold283 (.A(\i_main_reg.data_d[223] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold284 (.A(\i_main_reg.data_d[331] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold285 (.A(\i_main_reg.data_d[310] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold286 (.A(\i_main_reg.data_d[53] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0085_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold288 (.A(\i_main_reg.data_d[340] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold289 (.A(\i_main_reg.data_d[147] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0179_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold291 (.A(\i_main_reg.data_d[190] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold292 (.A(\i_main_reg.data_d[351] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0384_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold294 (.A(\i_main_reg.data_d[329] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0361_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold296 (.A(\i_main_reg.data_d[358] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold297 (.A(\i_main_reg.data_d[333] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0366_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold299 (.A(\i_main_reg.data_d[353] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0386_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold301 (.A(\i_main_reg.data_d[380] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0412_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold303 (.A(\i_main_reg.data_d[442] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold304 (.A(\i_main_reg.data_d[176] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold305 (.A(\i_main_reg.data_d[317] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold306 (.A(_0349_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold307 (.A(\i_main_reg.data_d[210] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0243_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold309 (.A(\i_main_reg.data_d[76] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold310 (.A(_0108_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold311 (.A(\i_main_reg.data_d[427] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold312 (.A(_0460_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold313 (.A(\i_main_reg.data_d[283] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0316_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold315 (.A(\i_main_reg.data_d[386] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold316 (.A(\i_main_reg.data_d[187] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0219_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold318 (.A(\i_main_reg.data_d[48] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold319 (.A(\i_main_reg.data_d[159] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0191_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold321 (.A(\one_count_q[1] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold322 (.A(_0481_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold323 (.A(\i_main_reg.data_d[78] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold324 (.A(_0110_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold325 (.A(\i_main_reg.data_d[157] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold326 (.A(_0190_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold327 (.A(\i_main_reg.data_d[413] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold328 (.A(\i_main_reg.data_d[54] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold329 (.A(\i_main_reg.data_d[300] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold330 (.A(_0333_),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold331 (.A(\i_main_reg.data_d[90] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold332 (.A(\i_main_reg.data_d[391] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold333 (.A(_0424_),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold334 (.A(\i_main_reg.data_d[402] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold335 (.A(\i_main_reg.data_d[142] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold336 (.A(_0174_),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold337 (.A(\i_main_reg.data_d[279] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold338 (.A(\i_main_reg.data_d[211] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold339 (.A(_0244_),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold340 (.A(\i_main_reg.data_d[175] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold341 (.A(\i_main_reg.data_d[436] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold342 (.A(_0469_),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold343 (.A(\i_main_reg.data_d[160] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold344 (.A(\i_main_reg.data_d[376] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold345 (.A(_0409_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold346 (.A(\i_main_reg.data_d[188] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold347 (.A(\i_main_reg.data_d[240] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0273_),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold349 (.A(\i_main_reg.data_d[143] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold350 (.A(\i_main_reg.data_d[207] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold351 (.A(_0239_),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold352 (.A(\i_main_reg.data_d[278] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold353 (.A(\i_main_reg.data_d[18] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold354 (.A(_0050_),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold355 (.A(\i_main_reg.data_d[323] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold356 (.A(_0356_),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold357 (.A(\i_main_reg.data_d[22] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold358 (.A(\i_main_reg.data_d[230] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold359 (.A(_0263_),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold360 (.A(\i_main_reg.data_d[45] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold361 (.A(\i_main_reg.data_d[26] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold362 (.A(\i_main_reg.data_d[106] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold363 (.A(_0138_),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold364 (.A(\i_main_reg.data_d[318] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold365 (.A(\i_main_reg.data_d[145] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold366 (.A(_0178_),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold367 (.A(\i_main_reg.data_d[179] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold368 (.A(\i_main_reg.data_d[352] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold369 (.A(\i_main_reg.data_d[75] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold370 (.A(\i_main_reg.data_d[213] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold371 (.A(_0246_),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold372 (.A(\i_main_reg.data_d[30] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0063_),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold374 (.A(\i_main_reg.data_d[375] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold375 (.A(\i_main_reg.data_d[203] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold376 (.A(\i_main_reg.data_d[401] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold377 (.A(\i_main_reg.data_d[10] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold378 (.A(_0042_),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold379 (.A(\i_main_reg.data_d[164] ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold380 (.A(_0197_),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold381 (.A(\i_main_reg.data_d[393] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold382 (.A(_0425_),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold383 (.A(\i_main_reg.data_d[32] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold384 (.A(_0064_),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold385 (.A(\i_main_reg.data_d[425] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold386 (.A(_0457_),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold387 (.A(\i_main_reg.data_d[343] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold388 (.A(\i_main_reg.data_d[430] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold389 (.A(\i_main_reg.data_d[38] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold390 (.A(_0070_),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold391 (.A(\i_main_reg.data_d[390] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold392 (.A(\i_main_reg.data_d[377] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold393 (.A(_0410_),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold394 (.A(\i_main_reg.data_d[261] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold395 (.A(_0294_),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold396 (.A(\i_main_reg.data_d[105] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold397 (.A(_0137_),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold398 (.A(\i_main_reg.data_d[219] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold399 (.A(\i_main_reg.data_d[417] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold400 (.A(\i_main_reg.data_d[348] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0381_),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold402 (.A(\i_main_reg.data_d[125] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold403 (.A(_0158_),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold404 (.A(\i_main_reg.data_d[3] ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold405 (.A(_0036_),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold406 (.A(\i_main_reg.data_d[49] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold407 (.A(_0082_),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold408 (.A(\i_main_reg.data_d[77] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold409 (.A(\i_main_reg.data_d[239] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold410 (.A(\i_main_reg.data_d[7] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold411 (.A(\i_main_reg.data_d[172] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold412 (.A(_0204_),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold413 (.A(\i_main_reg.data_d[374] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold414 (.A(\i_main_reg.data_d[299] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold415 (.A(\i_main_reg.data_d[277] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold416 (.A(\i_main_reg.data_d[173] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold417 (.A(\i_main_reg.data_d[337] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold418 (.A(\i_main_reg.data_d[435] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold419 (.A(\i_main_reg.data_d[273] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold420 (.A(_0306_),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold421 (.A(\i_main_reg.data_d[276] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold422 (.A(\i_main_reg.data_d[165] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0198_),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold424 (.A(\i_main_reg.data_d[243] ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold425 (.A(\i_main_reg.data_d[422] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold426 (.A(_0455_),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold427 (.A(\i_main_reg.data_d[237] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold428 (.A(_0270_),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold429 (.A(\i_main_reg.data_d[58] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold430 (.A(_0091_),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold431 (.A(\i_main_reg.data_d[107] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold432 (.A(\i_main_reg.data_d[389] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold433 (.A(\i_main_reg.data_d[282] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold434 (.A(\i_main_reg.data_d[396] ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold435 (.A(_0428_),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold436 (.A(\i_main_reg.data_d[132] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold437 (.A(_0165_),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold438 (.A(\i_main_reg.data_d[236] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold439 (.A(\i_main_reg.data_d[304] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold440 (.A(_0337_),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold441 (.A(\i_main_reg.data_d[216] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold442 (.A(_0249_),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold443 (.A(\i_main_reg.data_d[253] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold444 (.A(_0285_),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold445 (.A(\i_main_reg.data_d[221] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold446 (.A(_0254_),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold447 (.A(\i_main_reg.data_d[140] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold448 (.A(_0172_),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold449 (.A(\i_main_reg.data_d[394] ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold450 (.A(\i_main_reg.data_d[51] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold451 (.A(_0084_),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold452 (.A(\i_main_reg.data_d[298] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold453 (.A(\i_main_reg.data_d[275] ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold454 (.A(\i_main_reg.data_d[385] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold455 (.A(\i_main_reg.data_d[50] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold456 (.A(\i_main_reg.data_d[212] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold457 (.A(\i_main_reg.data_d[102] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold458 (.A(_0135_),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold459 (.A(\i_main_reg.data_d[429] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold460 (.A(\i_main_reg.data_d[24] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold461 (.A(_0057_),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold462 (.A(\i_main_reg.data_d[25] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold463 (.A(\i_main_reg.data_d[127] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold464 (.A(_0159_),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold465 (.A(\i_main_reg.data_d[222] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold466 (.A(\i_main_reg.data_d[79] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold467 (.A(\i_main_reg.data_d[411] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold468 (.A(_0444_),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold469 (.A(\i_main_reg.data_d[445] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold470 (.A(\i_main_reg.data_d[85] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold471 (.A(_0118_),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold472 (.A(\i_main_reg.data_d[443] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold473 (.A(\i_main_reg.data_d[296] ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold474 (.A(_0328_),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold475 (.A(\i_main_reg.data_d[255] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold476 (.A(_0287_),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold477 (.A(\bit_counter_q[9] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold478 (.A(\i_step_counter.data_o ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold479 (.A(_0000_),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold480 (.A(\i_main_reg.data_d[80] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold481 (.A(\i_main_reg.data_d[108] ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold482 (.A(\i_main_reg.data_d[73] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold483 (.A(_0105_),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold484 (.A(\i_main_reg.data_d[16] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold485 (.A(_0049_),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold486 (.A(\i_main_reg.data_d[57] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold487 (.A(\i_main_reg.data_d[294] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold488 (.A(_0327_),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold489 (.A(\i_main_reg.data_d[254] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold490 (.A(\i_main_reg.data_d[124] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold491 (.A(\i_main_reg.data_d[434] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold492 (.A(\i_main_reg.data_d[245] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold493 (.A(_0278_),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold494 (.A(\i_main_reg.data_d[66] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold495 (.A(_0099_),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold496 (.A(\i_main_reg.data_d[241] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold497 (.A(_0274_),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold498 (.A(\i_main_reg.data_d[308] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold499 (.A(_0340_),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold500 (.A(\i_main_reg.data_d[215] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold501 (.A(\i_main_reg.data_d[400] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold502 (.A(\i_main_reg.data_d[86] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold503 (.A(_0119_),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold504 (.A(\i_main_reg.data_d[89] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold505 (.A(\i_main_reg.data_d[309] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold506 (.A(\i_main_reg.data_d[274] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold507 (.A(\i_main_reg.data_d[214] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold508 (.A(\i_main_reg.data_d[328] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold509 (.A(_0360_),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold510 (.A(\i_main_reg.data_d[2] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold511 (.A(\i_main_reg.data_d[34] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold512 (.A(\i_main_reg.data_d[65] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold513 (.A(\i_main_reg.data_d[84] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold514 (.A(\i_main_reg.data_d[250] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold515 (.A(_0283_),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold516 (.A(\i_main_reg.data_d[4] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold517 (.A(_0037_),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold518 (.A(\i_main_reg.data_d[248] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold519 (.A(_0281_),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold520 (.A(\i_main_reg.data_d[151] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold521 (.A(_0183_),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold522 (.A(\i_main_reg.data_d[238] ),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold523 (.A(\i_main_reg.data_d[35] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold524 (.A(\i_main_reg.data_d[61] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold525 (.A(\i_main_reg.data_d[198] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold526 (.A(_0231_),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold527 (.A(\i_main_reg.data_d[418] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold528 (.A(\i_main_reg.data_d[306] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold529 (.A(_0339_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold530 (.A(\i_main_reg.data_d[133] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold531 (.A(_0166_),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold532 (.A(\i_main_reg.data_d[419] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold533 (.A(\i_main_reg.data_d[62] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold534 (.A(\i_main_reg.data_d[88] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold535 (.A(\i_main_reg.data_d[123] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold536 (.A(\i_main_reg.data_d[83] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold537 (.A(\i_main_reg.data_d[153] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold538 (.A(_0185_),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold539 (.A(\i_main_reg.data_d[139] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold540 (.A(\i_main_reg.data_d[63] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold541 (.A(\i_main_reg.data_d[81] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold542 (.A(_0114_),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold543 (.A(\i_main_reg.data_d[217] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold544 (.A(_0250_),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold545 (.A(\i_main_reg.data_d[8] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold546 (.A(\i_main_reg.data_d[388] ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold547 (.A(\i_main_reg.data_d[242] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold548 (.A(\i_main_reg.data_d[246] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold549 (.A(_0279_),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold550 (.A(\i_main_reg.data_d[103] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold551 (.A(_0136_),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold552 (.A(\i_main_reg.data_d[249] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold553 (.A(\i_main_reg.data_d[109] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold554 (.A(_0142_),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold555 (.A(\i_main_reg.data_d[424] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold556 (.A(_0456_),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold557 (.A(\i_main_reg.data_d[325] ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold558 (.A(_0358_),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold559 (.A(\i_main_reg.data_d[186] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold560 (.A(_0218_),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold561 (.A(\bit_counter_q[4] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold562 (.A(_0572_),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold563 (.A(\i_main_reg.data_d[9] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold564 (.A(\i_main_reg.data_d[293] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold565 (.A(\i_main_reg.data_d[395] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold566 (.A(\i_main_reg.data_d[326] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold567 (.A(_0359_),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold568 (.A(\i_main_reg.data_d[168] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold569 (.A(_0200_),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold570 (.A(\i_main_reg.data_d[64] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold571 (.A(\i_main_reg.data_d[87] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold572 (.A(\i_main_reg.data_d[235] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold573 (.A(_0267_),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold574 (.A(\i_main_reg.data_d[122] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold575 (.A(\i_main_reg.data_d[141] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold576 (.A(\i_main_reg.data_d[322] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold577 (.A(\i_main_reg.data_d[324] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold578 (.A(\i_main_reg.data_d[247] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold579 (.A(\i_main_reg.data_d[171] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold580 (.A(_0203_),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold581 (.A(\i_main_reg.data_d[265] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold582 (.A(_0297_),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold583 (.A(\i_main_reg.data_d[297] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold584 (.A(\i_main_reg.data_d[321] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold585 (.A(\i_main_reg.data_d[182] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold586 (.A(_0215_),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold587 (.A(\i_main_reg.data_d[46] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold588 (.A(\i_main_reg.data_d[404] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold589 (.A(_0437_),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold590 (.A(\i_main_reg.data_d[183] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold591 (.A(_0216_),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold592 (.A(\i_main_reg.data_d[347] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold593 (.A(\i_main_reg.data_d[71] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold594 (.A(_0104_),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold595 (.A(\i_main_reg.data_d[412] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold596 (.A(\i_main_reg.data_d[152] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold597 (.A(\i_main_reg.data_d[346] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold598 (.A(\i_main_reg.data_d[252] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold599 (.A(_0284_),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold600 (.A(\i_main_reg.data_d[319] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold601 (.A(\i_step_counter.data_d[8] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold602 (.A(_0008_),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold603 (.A(\i_main_reg.data_d[378] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold604 (.A(_0411_),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold605 (.A(\i_main_reg.data_d[135] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold606 (.A(_0168_),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold607 (.A(\i_main_reg.data_d[305] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold608 (.A(\i_main_reg.data_d[120] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold609 (.A(_0153_),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold610 (.A(\i_main_reg.data_d[166] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold611 (.A(_0199_),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold612 (.A(\i_main_reg.data_d[41] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold613 (.A(\i_step_counter.data_d[14] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold614 (.A(_0014_),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold615 (.A(\i_main_reg.data_d[110] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold616 (.A(_0143_),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold617 (.A(\i_main_reg.data_d[320] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold618 (.A(\i_main_reg.data_d[406] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold619 (.A(_0438_),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold620 (.A(\i_main_reg.data_d[42] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold621 (.A(\i_main_reg.data_d[407] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold622 (.A(\i_main_reg.data_d[344] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold623 (.A(\i_main_reg.data_d[428] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold624 (.A(\i_main_reg.data_d[233] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold625 (.A(_0265_),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold626 (.A(\i_main_reg.data_d[185] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold627 (.A(_0217_),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold628 (.A(\i_main_reg.data_d[268] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold629 (.A(_0300_),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold630 (.A(\i_main_reg.data_d[262] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold631 (.A(_0295_),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold632 (.A(carry_q),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold633 (.A(_0018_),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold634 (.A(\i_main_reg.data_d[169] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold635 (.A(\i_main_reg.data_d[345] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold636 (.A(\i_main_reg.data_d[36] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold637 (.A(_0069_),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold638 (.A(\i_main_reg.data_d[69] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold639 (.A(_0101_),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold640 (.A(\i_main_reg.data_d[234] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold641 (.A(\i_step_counter.data_d[7] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold642 (.A(_0513_),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold643 (.A(_0007_),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold644 (.A(\i_main_reg.data_d[231] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold645 (.A(_0264_),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold646 (.A(\i_main_reg.data_d[269] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold647 (.A(\i_main_reg.data_d[68] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold648 (.A(_0100_),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold649 (.A(\i_main_reg.data_d[264] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold650 (.A(_0296_),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold651 (.A(\i_main_reg.data_d[70] ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold652 (.A(\i_main_reg.data_d[408] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold653 (.A(\i_main_reg.data_d[134] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold654 (.A(\i_main_reg.data_d[82] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold655 (.A(\i_main_reg.data_d[170] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold656 (.A(\i_main_reg.data_d[266] ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold657 (.A(\i_main_reg.data_d[218] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold658 (.A(\bit_counter_q[5] ),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold659 (.A(_0025_),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold660 (.A(\i_main_reg.data_d[121] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold661 (.A(\i_main_reg.data_d[267] ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold662 (.A(\i_step_counter.data_d[12] ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold663 (.A(_0012_),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold664 (.A(\i_main_reg.data_d[199] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold665 (.A(_0232_),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold666 (.A(\i_step_counter.data_d[11] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold667 (.A(_0530_),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold668 (.A(_0011_),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold669 (.A(\bit_counter_q[3] ),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold670 (.A(\i_step_counter.data_d[13] ),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold671 (.A(_0013_),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold672 (.A(\i_step_counter.data_d[1] ),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold673 (.A(_0496_),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold674 (.A(_0002_),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold675 (.A(\i_step_counter.data_d[9] ),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold676 (.A(_0009_),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold677 (.A(\bit_counter_q[7] ),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold678 (.A(\state_q[0] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold679 (.A(\i_step_counter.data_d[2] ),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold680 (.A(_0499_),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold681 (.A(_0003_),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold682 (.A(\i_step_counter.data_d[5] ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold683 (.A(_0505_),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold684 (.A(_0005_),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold685 (.A(\i_step_counter.data_d[0] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold686 (.A(_0001_),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold687 (.A(previous_bit_q),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold688 (.A(_0019_),
    .X(net880));
 sg13g2_antennanp ANTENNA_1 (.A(_0203_));
 sg13g2_antennanp ANTENNA_2 (.A(_0234_));
 sg13g2_antennanp ANTENNA_3 (.A(_0319_));
 sg13g2_antennanp ANTENNA_4 (.A(_0319_));
 sg13g2_antennanp ANTENNA_5 (.A(_0325_));
 sg13g2_antennanp ANTENNA_6 (.A(_0339_));
 sg13g2_antennanp ANTENNA_7 (.A(_0339_));
 sg13g2_antennanp ANTENNA_8 (.A(_0381_));
 sg13g2_antennanp ANTENNA_9 (.A(_0381_));
 sg13g2_antennanp ANTENNA_10 (.A(\i_main_reg.data_d[166] ));
 sg13g2_antennanp ANTENNA_11 (.A(\i_main_reg.data_d[183] ));
 sg13g2_antennanp ANTENNA_12 (.A(\i_main_reg.data_d[183] ));
 sg13g2_antennanp ANTENNA_13 (.A(\i_main_reg.data_d[185] ));
 sg13g2_antennanp ANTENNA_14 (.A(\i_main_reg.data_d[186] ));
 sg13g2_antennanp ANTENNA_15 (.A(\i_main_reg.data_d[201] ));
 sg13g2_antennanp ANTENNA_16 (.A(\i_main_reg.data_d[261] ));
 sg13g2_antennanp ANTENNA_17 (.A(\i_main_reg.data_d[342] ));
 sg13g2_antennanp ANTENNA_18 (.A(\i_main_reg.data_d[342] ));
 sg13g2_antennanp ANTENNA_19 (.A(\i_main_reg.data_d[344] ));
 sg13g2_antennanp ANTENNA_20 (.A(net689));
 sg13g2_antennanp ANTENNA_21 (.A(_0207_));
 sg13g2_antennanp ANTENNA_22 (.A(_0214_));
 sg13g2_antennanp ANTENNA_23 (.A(_0232_));
 sg13g2_antennanp ANTENNA_24 (.A(_0232_));
 sg13g2_antennanp ANTENNA_25 (.A(\i_main_reg.data_d[171] ));
 sg13g2_antennanp ANTENNA_26 (.A(\i_main_reg.data_d[171] ));
 sg13g2_antennanp ANTENNA_27 (.A(\i_main_reg.data_d[174] ));
 sg13g2_antennanp ANTENNA_28 (.A(\i_main_reg.data_d[178] ));
 sg13g2_antennanp ANTENNA_29 (.A(\i_main_reg.data_d[187] ));
 sg13g2_antennanp ANTENNA_30 (.A(\i_main_reg.data_d[191] ));
 sg13g2_antennanp ANTENNA_31 (.A(\i_main_reg.data_d[194] ));
 sg13g2_antennanp ANTENNA_32 (.A(\i_main_reg.data_d[276] ));
 sg13g2_antennanp ANTENNA_33 (.A(\i_main_reg.data_d[325] ));
 sg13g2_antennanp ANTENNA_34 (.A(\i_main_reg.data_d[325] ));
 sg13g2_antennanp ANTENNA_35 (.A(net207));
 sg13g2_antennanp ANTENNA_36 (.A(\i_main_reg.data_d[197] ));
 sg13g2_antennanp ANTENNA_37 (.A(\i_main_reg.data_d[197] ));
 sg13g2_antennanp ANTENNA_38 (.A(\i_main_reg.data_d[330] ));
 sg13g2_antennanp ANTENNA_39 (.A(\i_main_reg.data_d[331] ));
 sg13g2_antennanp ANTENNA_40 (.A(\i_main_reg.data_d[331] ));
 sg13g2_decap_4 FILLER_0_163 ();
 sg13g2_decap_4 FILLER_0_216 ();
 sg13g2_fill_2 FILLER_0_230 ();
 sg13g2_fill_1 FILLER_0_232 ();
 sg13g2_decap_4 FILLER_0_296 ();
 sg13g2_fill_2 FILLER_0_300 ();
 sg13g2_fill_1 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_402 ();
 sg13g2_fill_2 FILLER_1_0 ();
 sg13g2_fill_1 FILLER_1_11 ();
 sg13g2_decap_4 FILLER_1_24 ();
 sg13g2_fill_1 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_fill_1 FILLER_1_140 ();
 sg13g2_decap_4 FILLER_1_205 ();
 sg13g2_fill_2 FILLER_1_209 ();
 sg13g2_decap_8 FILLER_1_284 ();
 sg13g2_fill_1 FILLER_1_291 ();
 sg13g2_fill_1 FILLER_1_311 ();
 sg13g2_decap_4 FILLER_1_405 ();
 sg13g2_fill_2 FILLER_2_0 ();
 sg13g2_decap_4 FILLER_2_5 ();
 sg13g2_decap_8 FILLER_2_48 ();
 sg13g2_fill_1 FILLER_2_55 ();
 sg13g2_fill_2 FILLER_2_138 ();
 sg13g2_fill_1 FILLER_2_140 ();
 sg13g2_decap_4 FILLER_2_249 ();
 sg13g2_decap_4 FILLER_2_271 ();
 sg13g2_fill_1 FILLER_2_275 ();
 sg13g2_decap_8 FILLER_2_402 ();
 sg13g2_fill_2 FILLER_3_0 ();
 sg13g2_fill_1 FILLER_3_2 ();
 sg13g2_decap_4 FILLER_3_27 ();
 sg13g2_fill_2 FILLER_3_31 ();
 sg13g2_fill_2 FILLER_3_81 ();
 sg13g2_fill_1 FILLER_3_83 ();
 sg13g2_fill_2 FILLER_3_138 ();
 sg13g2_fill_2 FILLER_3_224 ();
 sg13g2_fill_1 FILLER_3_255 ();
 sg13g2_fill_2 FILLER_3_276 ();
 sg13g2_fill_1 FILLER_3_278 ();
 sg13g2_fill_2 FILLER_3_347 ();
 sg13g2_fill_1 FILLER_3_349 ();
 sg13g2_decap_4 FILLER_3_404 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_4 FILLER_4_131 ();
 sg13g2_fill_1 FILLER_4_135 ();
 sg13g2_decap_4 FILLER_4_183 ();
 sg13g2_fill_2 FILLER_4_187 ();
 sg13g2_fill_1 FILLER_4_255 ();
 sg13g2_fill_2 FILLER_4_279 ();
 sg13g2_fill_1 FILLER_4_281 ();
 sg13g2_decap_4 FILLER_4_319 ();
 sg13g2_fill_2 FILLER_4_323 ();
 sg13g2_decap_4 FILLER_4_335 ();
 sg13g2_decap_4 FILLER_4_352 ();
 sg13g2_fill_2 FILLER_4_356 ();
 sg13g2_decap_4 FILLER_4_405 ();
 sg13g2_fill_1 FILLER_5_0 ();
 sg13g2_fill_2 FILLER_5_10 ();
 sg13g2_fill_1 FILLER_5_12 ();
 sg13g2_fill_2 FILLER_5_25 ();
 sg13g2_decap_4 FILLER_5_81 ();
 sg13g2_fill_2 FILLER_5_85 ();
 sg13g2_fill_2 FILLER_5_164 ();
 sg13g2_fill_2 FILLER_5_179 ();
 sg13g2_fill_1 FILLER_5_314 ();
 sg13g2_fill_2 FILLER_5_335 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_fill_2 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_11 ();
 sg13g2_fill_2 FILLER_6_16 ();
 sg13g2_fill_1 FILLER_6_48 ();
 sg13g2_fill_2 FILLER_6_79 ();
 sg13g2_decap_4 FILLER_6_147 ();
 sg13g2_fill_1 FILLER_6_151 ();
 sg13g2_decap_8 FILLER_6_172 ();
 sg13g2_decap_4 FILLER_6_216 ();
 sg13g2_fill_2 FILLER_6_220 ();
 sg13g2_fill_2 FILLER_6_397 ();
 sg13g2_fill_1 FILLER_7_9 ();
 sg13g2_fill_2 FILLER_7_22 ();
 sg13g2_fill_1 FILLER_7_24 ();
 sg13g2_decap_4 FILLER_7_55 ();
 sg13g2_fill_1 FILLER_7_59 ();
 sg13g2_fill_1 FILLER_7_78 ();
 sg13g2_fill_2 FILLER_7_148 ();
 sg13g2_fill_1 FILLER_7_150 ();
 sg13g2_decap_4 FILLER_7_178 ();
 sg13g2_fill_2 FILLER_7_182 ();
 sg13g2_fill_2 FILLER_7_197 ();
 sg13g2_fill_1 FILLER_7_286 ();
 sg13g2_fill_2 FILLER_7_318 ();
 sg13g2_fill_1 FILLER_7_320 ();
 sg13g2_decap_4 FILLER_7_348 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_4 FILLER_8_46 ();
 sg13g2_fill_1 FILLER_8_77 ();
 sg13g2_decap_4 FILLER_8_259 ();
 sg13g2_fill_1 FILLER_8_263 ();
 sg13g2_decap_8 FILLER_8_314 ();
 sg13g2_fill_1 FILLER_8_321 ();
 sg13g2_decap_4 FILLER_8_403 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_fill_2 FILLER_9_27 ();
 sg13g2_decap_4 FILLER_9_50 ();
 sg13g2_fill_1 FILLER_9_54 ();
 sg13g2_decap_4 FILLER_9_73 ();
 sg13g2_fill_2 FILLER_9_124 ();
 sg13g2_fill_1 FILLER_9_149 ();
 sg13g2_decap_4 FILLER_9_214 ();
 sg13g2_fill_1 FILLER_9_218 ();
 sg13g2_decap_8 FILLER_9_242 ();
 sg13g2_fill_1 FILLER_9_249 ();
 sg13g2_fill_2 FILLER_9_280 ();
 sg13g2_fill_1 FILLER_9_295 ();
 sg13g2_decap_4 FILLER_9_309 ();
 sg13g2_decap_8 FILLER_9_333 ();
 sg13g2_decap_4 FILLER_9_379 ();
 sg13g2_decap_4 FILLER_9_403 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_4 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_4 ();
 sg13g2_fill_2 FILLER_10_15 ();
 sg13g2_fill_1 FILLER_10_17 ();
 sg13g2_fill_1 FILLER_10_72 ();
 sg13g2_decap_4 FILLER_10_109 ();
 sg13g2_fill_2 FILLER_10_130 ();
 sg13g2_fill_1 FILLER_10_132 ();
 sg13g2_fill_1 FILLER_10_237 ();
 sg13g2_decap_4 FILLER_10_381 ();
 sg13g2_fill_1 FILLER_10_385 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_2 ();
 sg13g2_decap_4 FILLER_11_66 ();
 sg13g2_fill_2 FILLER_11_70 ();
 sg13g2_fill_2 FILLER_11_119 ();
 sg13g2_fill_1 FILLER_11_121 ();
 sg13g2_fill_2 FILLER_11_185 ();
 sg13g2_decap_4 FILLER_11_200 ();
 sg13g2_decap_8 FILLER_11_267 ();
 sg13g2_fill_1 FILLER_11_274 ();
 sg13g2_decap_4 FILLER_11_302 ();
 sg13g2_fill_2 FILLER_11_306 ();
 sg13g2_decap_8 FILLER_11_335 ();
 sg13g2_decap_4 FILLER_11_369 ();
 sg13g2_decap_8 FILLER_11_386 ();
 sg13g2_decap_4 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_4 FILLER_12_34 ();
 sg13g2_fill_1 FILLER_12_38 ();
 sg13g2_decap_8 FILLER_12_190 ();
 sg13g2_fill_1 FILLER_12_197 ();
 sg13g2_decap_8 FILLER_12_211 ();
 sg13g2_fill_2 FILLER_12_272 ();
 sg13g2_fill_1 FILLER_12_274 ();
 sg13g2_decap_4 FILLER_12_393 ();
 sg13g2_fill_2 FILLER_12_397 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_43 ();
 sg13g2_decap_4 FILLER_13_76 ();
 sg13g2_decap_4 FILLER_13_107 ();
 sg13g2_decap_8 FILLER_13_173 ();
 sg13g2_fill_1 FILLER_13_236 ();
 sg13g2_fill_2 FILLER_13_317 ();
 sg13g2_decap_8 FILLER_13_346 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_2 ();
 sg13g2_fill_2 FILLER_14_12 ();
 sg13g2_fill_2 FILLER_14_32 ();
 sg13g2_fill_1 FILLER_14_34 ();
 sg13g2_fill_2 FILLER_14_47 ();
 sg13g2_fill_2 FILLER_14_106 ();
 sg13g2_fill_1 FILLER_14_184 ();
 sg13g2_fill_1 FILLER_14_225 ();
 sg13g2_fill_2 FILLER_14_273 ();
 sg13g2_fill_1 FILLER_14_275 ();
 sg13g2_fill_2 FILLER_14_289 ();
 sg13g2_decap_4 FILLER_14_304 ();
 sg13g2_fill_2 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_333 ();
 sg13g2_fill_1 FILLER_14_340 ();
 sg13g2_decap_8 FILLER_14_367 ();
 sg13g2_fill_1 FILLER_14_374 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_decap_4 FILLER_15_27 ();
 sg13g2_fill_1 FILLER_15_31 ();
 sg13g2_fill_1 FILLER_15_115 ();
 sg13g2_decap_4 FILLER_15_129 ();
 sg13g2_fill_2 FILLER_15_133 ();
 sg13g2_fill_2 FILLER_15_162 ();
 sg13g2_decap_8 FILLER_15_191 ();
 sg13g2_fill_1 FILLER_15_198 ();
 sg13g2_decap_4 FILLER_15_253 ();
 sg13g2_fill_2 FILLER_15_257 ();
 sg13g2_fill_1 FILLER_15_279 ();
 sg13g2_fill_1 FILLER_15_310 ();
 sg13g2_decap_4 FILLER_15_371 ();
 sg13g2_fill_1 FILLER_15_375 ();
 sg13g2_decap_4 FILLER_15_403 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_20 ();
 sg13g2_decap_4 FILLER_16_72 ();
 sg13g2_fill_1 FILLER_16_76 ();
 sg13g2_decap_4 FILLER_16_131 ();
 sg13g2_fill_1 FILLER_16_135 ();
 sg13g2_fill_2 FILLER_16_163 ();
 sg13g2_fill_1 FILLER_16_165 ();
 sg13g2_fill_2 FILLER_16_179 ();
 sg13g2_fill_2 FILLER_16_194 ();
 sg13g2_fill_1 FILLER_16_196 ();
 sg13g2_decap_4 FILLER_16_251 ();
 sg13g2_fill_1 FILLER_16_255 ();
 sg13g2_fill_2 FILLER_16_283 ();
 sg13g2_fill_2 FILLER_16_343 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_14 ();
 sg13g2_fill_2 FILLER_17_18 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_fill_1 FILLER_17_209 ();
 sg13g2_fill_1 FILLER_17_223 ();
 sg13g2_fill_2 FILLER_17_278 ();
 sg13g2_fill_1 FILLER_17_334 ();
 sg13g2_fill_2 FILLER_17_339 ();
 sg13g2_fill_1 FILLER_17_341 ();
 sg13g2_decap_8 FILLER_17_369 ();
 sg13g2_decap_4 FILLER_17_403 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_2 ();
 sg13g2_fill_1 FILLER_18_15 ();
 sg13g2_fill_2 FILLER_18_28 ();
 sg13g2_decap_4 FILLER_18_69 ();
 sg13g2_fill_1 FILLER_18_73 ();
 sg13g2_fill_1 FILLER_18_110 ();
 sg13g2_decap_4 FILLER_18_168 ();
 sg13g2_fill_1 FILLER_18_172 ();
 sg13g2_decap_8 FILLER_18_240 ();
 sg13g2_fill_2 FILLER_18_334 ();
 sg13g2_fill_1 FILLER_18_336 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_fill_1 FILLER_19_12 ();
 sg13g2_fill_2 FILLER_19_61 ();
 sg13g2_decap_4 FILLER_19_121 ();
 sg13g2_fill_1 FILLER_19_125 ();
 sg13g2_fill_2 FILLER_19_182 ();
 sg13g2_fill_1 FILLER_19_184 ();
 sg13g2_decap_4 FILLER_19_212 ();
 sg13g2_decap_4 FILLER_19_226 ();
 sg13g2_decap_4 FILLER_19_240 ();
 sg13g2_fill_2 FILLER_19_244 ();
 sg13g2_fill_2 FILLER_19_299 ();
 sg13g2_fill_1 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_312 ();
 sg13g2_fill_1 FILLER_19_319 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_20 ();
 sg13g2_decap_8 FILLER_20_27 ();
 sg13g2_decap_4 FILLER_20_34 ();
 sg13g2_fill_2 FILLER_20_59 ();
 sg13g2_fill_1 FILLER_20_217 ();
 sg13g2_fill_1 FILLER_20_245 ();
 sg13g2_fill_2 FILLER_20_273 ();
 sg13g2_fill_2 FILLER_20_369 ();
 sg13g2_fill_1 FILLER_20_371 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_11 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_65 ();
 sg13g2_fill_1 FILLER_21_72 ();
 sg13g2_decap_8 FILLER_21_86 ();
 sg13g2_decap_4 FILLER_21_123 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_fill_1 FILLER_21_161 ();
 sg13g2_decap_4 FILLER_21_189 ();
 sg13g2_decap_4 FILLER_21_203 ();
 sg13g2_fill_2 FILLER_21_207 ();
 sg13g2_decap_8 FILLER_21_236 ();
 sg13g2_fill_1 FILLER_21_243 ();
 sg13g2_fill_1 FILLER_21_398 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_4 FILLER_22_42 ();
 sg13g2_fill_1 FILLER_22_46 ();
 sg13g2_fill_1 FILLER_22_256 ();
 sg13g2_decap_4 FILLER_22_267 ();
 sg13g2_fill_2 FILLER_22_284 ();
 sg13g2_fill_2 FILLER_22_313 ();
 sg13g2_fill_1 FILLER_22_315 ();
 sg13g2_fill_2 FILLER_22_343 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_fill_2 FILLER_23_49 ();
 sg13g2_fill_1 FILLER_23_51 ();
 sg13g2_fill_2 FILLER_23_130 ();
 sg13g2_fill_1 FILLER_23_132 ();
 sg13g2_fill_1 FILLER_23_233 ();
 sg13g2_fill_2 FILLER_23_271 ();
 sg13g2_fill_1 FILLER_23_273 ();
 sg13g2_fill_1 FILLER_23_287 ();
 sg13g2_fill_2 FILLER_23_380 ();
 sg13g2_fill_1 FILLER_23_382 ();
 sg13g2_decap_4 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_4 FILLER_24_42 ();
 sg13g2_fill_2 FILLER_24_46 ();
 sg13g2_fill_1 FILLER_24_129 ();
 sg13g2_fill_2 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_186 ();
 sg13g2_decap_4 FILLER_24_230 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_fill_1 FILLER_24_308 ();
 sg13g2_decap_4 FILLER_24_332 ();
 sg13g2_decap_4 FILLER_24_363 ();
 sg13g2_decap_4 FILLER_24_403 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_fill_1 FILLER_25_42 ();
 sg13g2_fill_2 FILLER_25_179 ();
 sg13g2_fill_2 FILLER_25_321 ();
 sg13g2_fill_1 FILLER_25_323 ();
 sg13g2_fill_1 FILLER_25_351 ();
 sg13g2_decap_8 FILLER_25_365 ();
 sg13g2_fill_1 FILLER_25_372 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_4 FILLER_26_42 ();
 sg13g2_fill_2 FILLER_26_140 ();
 sg13g2_fill_2 FILLER_26_195 ();
 sg13g2_fill_1 FILLER_26_197 ();
 sg13g2_fill_1 FILLER_26_221 ();
 sg13g2_fill_2 FILLER_26_367 ();
 sg13g2_fill_1 FILLER_26_369 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_4 FILLER_27_35 ();
 sg13g2_fill_1 FILLER_27_39 ();
 sg13g2_decap_8 FILLER_27_123 ();
 sg13g2_fill_1 FILLER_27_130 ();
 sg13g2_fill_2 FILLER_27_157 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_fill_1 FILLER_27_223 ();
 sg13g2_fill_1 FILLER_27_325 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_4 FILLER_28_35 ();
 sg13g2_fill_2 FILLER_28_39 ();
 sg13g2_decap_4 FILLER_28_183 ();
 sg13g2_decap_4 FILLER_28_259 ();
 sg13g2_fill_2 FILLER_28_263 ();
 sg13g2_decap_4 FILLER_28_354 ();
 sg13g2_fill_1 FILLER_28_358 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_fill_1 FILLER_29_35 ();
 sg13g2_decap_4 FILLER_29_100 ();
 sg13g2_decap_4 FILLER_29_127 ();
 sg13g2_fill_1 FILLER_29_131 ();
 sg13g2_decap_4 FILLER_29_159 ();
 sg13g2_decap_8 FILLER_29_248 ();
 sg13g2_fill_2 FILLER_29_292 ();
 sg13g2_fill_1 FILLER_29_294 ();
 sg13g2_decap_8 FILLER_29_402 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_4 FILLER_30_28 ();
 sg13g2_fill_2 FILLER_30_149 ();
 sg13g2_decap_4 FILLER_30_205 ();
 sg13g2_fill_2 FILLER_30_209 ();
 sg13g2_decap_4 FILLER_30_238 ();
 sg13g2_fill_2 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_358 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_4 FILLER_31_28 ();
 sg13g2_fill_2 FILLER_31_105 ();
 sg13g2_fill_1 FILLER_31_144 ();
 sg13g2_fill_2 FILLER_31_158 ();
 sg13g2_decap_4 FILLER_31_193 ();
 sg13g2_fill_2 FILLER_31_197 ();
 sg13g2_decap_4 FILLER_31_226 ();
 sg13g2_decap_4 FILLER_31_287 ();
 sg13g2_decap_4 FILLER_31_318 ();
 sg13g2_fill_1 FILLER_31_332 ();
 sg13g2_decap_4 FILLER_31_360 ();
 sg13g2_fill_1 FILLER_31_364 ();
 sg13g2_decap_8 FILLER_31_401 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_4 FILLER_32_28 ();
 sg13g2_fill_1 FILLER_32_128 ();
 sg13g2_fill_1 FILLER_32_192 ();
 sg13g2_fill_2 FILLER_32_256 ();
 sg13g2_decap_4 FILLER_32_300 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_fill_2 FILLER_33_35 ();
 sg13g2_fill_1 FILLER_33_122 ();
 sg13g2_decap_8 FILLER_33_159 ();
 sg13g2_fill_2 FILLER_33_193 ();
 sg13g2_fill_1 FILLER_33_224 ();
 sg13g2_fill_2 FILLER_33_349 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_4 FILLER_34_94 ();
 sg13g2_fill_2 FILLER_34_98 ();
 sg13g2_decap_4 FILLER_34_127 ();
 sg13g2_fill_1 FILLER_34_131 ();
 sg13g2_decap_4 FILLER_34_159 ();
 sg13g2_fill_1 FILLER_34_163 ();
 sg13g2_decap_4 FILLER_34_201 ();
 sg13g2_fill_1 FILLER_34_205 ();
 sg13g2_fill_2 FILLER_34_233 ();
 sg13g2_decap_4 FILLER_34_282 ();
 sg13g2_fill_2 FILLER_34_286 ();
 sg13g2_fill_2 FILLER_34_311 ();
 sg13g2_fill_1 FILLER_34_313 ();
 sg13g2_decap_4 FILLER_34_341 ();
 sg13g2_fill_2 FILLER_34_345 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_fill_2 FILLER_35_28 ();
 sg13g2_fill_2 FILLER_35_93 ();
 sg13g2_decap_4 FILLER_35_149 ();
 sg13g2_fill_2 FILLER_35_176 ();
 sg13g2_decap_8 FILLER_35_309 ();
 sg13g2_decap_8 FILLER_35_401 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_4 FILLER_36_28 ();
 sg13g2_fill_1 FILLER_36_32 ();
 sg13g2_fill_1 FILLER_36_120 ();
 sg13g2_decap_4 FILLER_36_148 ();
 sg13g2_fill_2 FILLER_36_152 ();
 sg13g2_decap_4 FILLER_36_217 ();
 sg13g2_decap_4 FILLER_36_248 ();
 sg13g2_fill_1 FILLER_36_252 ();
 sg13g2_decap_8 FILLER_36_263 ();
 sg13g2_fill_2 FILLER_36_315 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_fill_2 FILLER_37_28 ();
 sg13g2_decap_4 FILLER_37_93 ();
 sg13g2_fill_2 FILLER_37_97 ();
 sg13g2_decap_4 FILLER_37_126 ();
 sg13g2_fill_2 FILLER_37_130 ();
 sg13g2_decap_8 FILLER_37_142 ();
 sg13g2_decap_4 FILLER_37_223 ();
 sg13g2_fill_2 FILLER_37_227 ();
 sg13g2_fill_1 FILLER_37_242 ();
 sg13g2_fill_1 FILLER_37_275 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_4 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_117 ();
 sg13g2_fill_1 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_181 ();
 sg13g2_fill_2 FILLER_38_185 ();
 sg13g2_decap_8 FILLER_38_219 ();
 sg13g2_fill_1 FILLER_38_226 ();
 sg13g2_decap_4 FILLER_38_237 ();
 sg13g2_fill_2 FILLER_38_241 ();
 sg13g2_decap_8 FILLER_38_253 ();
 sg13g2_fill_2 FILLER_38_386 ();
 sg13g2_fill_1 FILLER_38_388 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_fill_2 FILLER_39_28 ();
 sg13g2_fill_1 FILLER_39_30 ();
 sg13g2_fill_2 FILLER_39_94 ();
 sg13g2_fill_1 FILLER_39_96 ();
 sg13g2_fill_2 FILLER_39_124 ();
 sg13g2_fill_1 FILLER_39_227 ();
 sg13g2_fill_2 FILLER_39_292 ();
 sg13g2_decap_4 FILLER_39_405 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_fill_2 FILLER_40_42 ();
 sg13g2_fill_1 FILLER_40_89 ();
 sg13g2_fill_2 FILLER_40_117 ();
 sg13g2_fill_1 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_157 ();
 sg13g2_fill_2 FILLER_40_200 ();
 sg13g2_fill_2 FILLER_40_310 ();
 sg13g2_fill_1 FILLER_40_312 ();
 sg13g2_decap_4 FILLER_40_404 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_fill_2 FILLER_41_42 ();
 sg13g2_fill_1 FILLER_41_89 ();
 sg13g2_fill_2 FILLER_41_117 ();
 sg13g2_decap_4 FILLER_41_166 ();
 sg13g2_fill_1 FILLER_41_170 ();
 sg13g2_decap_4 FILLER_41_264 ();
 sg13g2_fill_1 FILLER_41_268 ();
 sg13g2_decap_4 FILLER_41_405 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_4 FILLER_42_35 ();
 sg13g2_decap_4 FILLER_42_85 ();
 sg13g2_fill_1 FILLER_42_89 ();
 sg13g2_fill_1 FILLER_42_183 ();
 sg13g2_fill_2 FILLER_42_194 ();
 sg13g2_fill_2 FILLER_42_249 ();
 sg13g2_decap_8 FILLER_42_264 ();
 sg13g2_fill_2 FILLER_42_377 ();
 sg13g2_fill_2 FILLER_42_406 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_4 FILLER_43_35 ();
 sg13g2_fill_1 FILLER_43_39 ();
 sg13g2_decap_4 FILLER_43_100 ();
 sg13g2_fill_2 FILLER_43_104 ();
 sg13g2_fill_2 FILLER_43_182 ();
 sg13g2_fill_1 FILLER_43_385 ();
 sg13g2_decap_4 FILLER_43_395 ();
 sg13g2_fill_1 FILLER_43_399 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_4 FILLER_44_28 ();
 sg13g2_fill_2 FILLER_44_32 ();
 sg13g2_decap_4 FILLER_44_107 ();
 sg13g2_fill_2 FILLER_44_111 ();
 sg13g2_decap_4 FILLER_44_167 ();
 sg13g2_fill_2 FILLER_44_171 ();
 sg13g2_decap_4 FILLER_44_200 ();
 sg13g2_fill_2 FILLER_44_204 ();
 sg13g2_decap_4 FILLER_44_233 ();
 sg13g2_fill_1 FILLER_44_237 ();
 sg13g2_fill_2 FILLER_44_347 ();
 sg13g2_fill_1 FILLER_44_349 ();
 sg13g2_decap_8 FILLER_44_377 ();
 sg13g2_fill_1 FILLER_44_384 ();
 sg13g2_fill_1 FILLER_44_394 ();
 sg13g2_decap_4 FILLER_44_404 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_4 FILLER_45_35 ();
 sg13g2_fill_1 FILLER_45_39 ();
 sg13g2_decap_8 FILLER_45_166 ();
 sg13g2_decap_4 FILLER_45_200 ();
 sg13g2_fill_2 FILLER_45_204 ();
 sg13g2_decap_4 FILLER_45_293 ();
 sg13g2_fill_2 FILLER_45_297 ();
 sg13g2_decap_8 FILLER_45_353 ();
 sg13g2_decap_8 FILLER_45_360 ();
 sg13g2_decap_8 FILLER_45_367 ();
 sg13g2_decap_8 FILLER_45_374 ();
 sg13g2_decap_8 FILLER_45_381 ();
 sg13g2_fill_2 FILLER_45_388 ();
 sg13g2_fill_1 FILLER_45_390 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_4 FILLER_46_21 ();
 sg13g2_decap_4 FILLER_46_89 ();
 sg13g2_fill_1 FILLER_46_93 ();
 sg13g2_fill_1 FILLER_46_121 ();
 sg13g2_fill_2 FILLER_46_159 ();
 sg13g2_fill_1 FILLER_46_161 ();
 sg13g2_fill_2 FILLER_46_202 ();
 sg13g2_fill_2 FILLER_46_270 ();
 sg13g2_decap_8 FILLER_46_344 ();
 sg13g2_decap_8 FILLER_46_351 ();
 sg13g2_decap_8 FILLER_46_358 ();
 sg13g2_decap_8 FILLER_46_365 ();
 sg13g2_decap_8 FILLER_46_372 ();
 sg13g2_decap_8 FILLER_46_379 ();
 sg13g2_decap_8 FILLER_46_386 ();
 sg13g2_fill_2 FILLER_46_393 ();
 sg13g2_fill_1 FILLER_46_395 ();
 sg13g2_decap_4 FILLER_46_405 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_4 FILLER_47_28 ();
 sg13g2_fill_1 FILLER_47_32 ();
 sg13g2_decap_4 FILLER_47_92 ();
 sg13g2_fill_1 FILLER_47_96 ();
 sg13g2_decap_4 FILLER_47_110 ();
 sg13g2_fill_1 FILLER_47_114 ();
 sg13g2_decap_8 FILLER_47_141 ();
 sg13g2_fill_1 FILLER_47_148 ();
 sg13g2_fill_2 FILLER_47_175 ();
 sg13g2_fill_1 FILLER_47_177 ();
 sg13g2_fill_1 FILLER_47_228 ();
 sg13g2_fill_2 FILLER_47_274 ();
 sg13g2_decap_8 FILLER_47_353 ();
 sg13g2_decap_8 FILLER_47_360 ();
 sg13g2_decap_8 FILLER_47_367 ();
 sg13g2_decap_8 FILLER_47_374 ();
 sg13g2_decap_8 FILLER_47_381 ();
 sg13g2_decap_8 FILLER_47_388 ();
 sg13g2_decap_8 FILLER_47_395 ();
 sg13g2_decap_8 FILLER_47_402 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_fill_1 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_135 ();
 sg13g2_fill_1 FILLER_48_152 ();
 sg13g2_fill_1 FILLER_48_193 ();
 sg13g2_decap_4 FILLER_48_221 ();
 sg13g2_fill_2 FILLER_48_277 ();
 sg13g2_decap_8 FILLER_48_355 ();
 sg13g2_decap_8 FILLER_48_362 ();
 sg13g2_decap_8 FILLER_48_369 ();
 sg13g2_decap_8 FILLER_48_376 ();
 sg13g2_decap_8 FILLER_48_383 ();
 sg13g2_decap_8 FILLER_48_390 ();
 sg13g2_decap_8 FILLER_48_397 ();
 sg13g2_decap_4 FILLER_48_404 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_fill_2 FILLER_49_21 ();
 sg13g2_fill_1 FILLER_49_23 ();
 sg13g2_fill_2 FILLER_49_144 ();
 sg13g2_decap_8 FILLER_49_193 ();
 sg13g2_fill_2 FILLER_49_250 ();
 sg13g2_fill_2 FILLER_49_279 ();
 sg13g2_decap_8 FILLER_49_364 ();
 sg13g2_decap_8 FILLER_49_371 ();
 sg13g2_decap_8 FILLER_49_378 ();
 sg13g2_decap_8 FILLER_49_385 ();
 sg13g2_decap_8 FILLER_49_392 ();
 sg13g2_decap_8 FILLER_49_399 ();
 sg13g2_fill_2 FILLER_49_406 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_fill_2 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_89 ();
 sg13g2_fill_1 FILLER_50_96 ();
 sg13g2_fill_2 FILLER_50_110 ();
 sg13g2_fill_2 FILLER_50_316 ();
 sg13g2_decap_8 FILLER_50_359 ();
 sg13g2_decap_8 FILLER_50_366 ();
 sg13g2_decap_8 FILLER_50_373 ();
 sg13g2_decap_8 FILLER_50_380 ();
 sg13g2_decap_8 FILLER_50_387 ();
 sg13g2_decap_8 FILLER_50_394 ();
 sg13g2_decap_8 FILLER_50_401 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_fill_2 FILLER_51_14 ();
 sg13g2_fill_1 FILLER_51_16 ();
 sg13g2_fill_1 FILLER_51_89 ();
 sg13g2_fill_1 FILLER_51_117 ();
 sg13g2_fill_1 FILLER_51_158 ();
 sg13g2_fill_1 FILLER_51_249 ();
 sg13g2_decap_8 FILLER_51_367 ();
 sg13g2_decap_8 FILLER_51_374 ();
 sg13g2_decap_8 FILLER_51_381 ();
 sg13g2_decap_8 FILLER_51_388 ();
 sg13g2_decap_8 FILLER_51_395 ();
 sg13g2_decap_8 FILLER_51_402 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_4 FILLER_52_21 ();
 sg13g2_fill_2 FILLER_52_25 ();
 sg13g2_decap_4 FILLER_52_97 ();
 sg13g2_decap_8 FILLER_52_171 ();
 sg13g2_fill_1 FILLER_52_178 ();
 sg13g2_decap_4 FILLER_52_202 ();
 sg13g2_fill_1 FILLER_52_206 ();
 sg13g2_decap_8 FILLER_52_365 ();
 sg13g2_decap_8 FILLER_52_372 ();
 sg13g2_decap_8 FILLER_52_379 ();
 sg13g2_decap_8 FILLER_52_386 ();
 sg13g2_decap_8 FILLER_52_393 ();
 sg13g2_decap_8 FILLER_52_400 ();
 sg13g2_fill_2 FILLER_52_407 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_4 FILLER_53_28 ();
 sg13g2_fill_2 FILLER_53_32 ();
 sg13g2_decap_4 FILLER_53_89 ();
 sg13g2_fill_1 FILLER_53_120 ();
 sg13g2_decap_8 FILLER_53_158 ();
 sg13g2_decap_8 FILLER_53_185 ();
 sg13g2_fill_1 FILLER_53_192 ();
 sg13g2_decap_4 FILLER_53_240 ();
 sg13g2_fill_2 FILLER_53_271 ();
 sg13g2_fill_1 FILLER_53_273 ();
 sg13g2_decap_8 FILLER_53_364 ();
 sg13g2_decap_8 FILLER_53_371 ();
 sg13g2_decap_8 FILLER_53_378 ();
 sg13g2_decap_8 FILLER_53_385 ();
 sg13g2_decap_8 FILLER_53_392 ();
 sg13g2_decap_8 FILLER_53_399 ();
 sg13g2_fill_2 FILLER_53_406 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_4 FILLER_54_21 ();
 sg13g2_fill_2 FILLER_54_99 ();
 sg13g2_fill_2 FILLER_54_154 ();
 sg13g2_fill_2 FILLER_54_160 ();
 sg13g2_fill_2 FILLER_54_175 ();
 sg13g2_fill_1 FILLER_54_177 ();
 sg13g2_fill_2 FILLER_54_215 ();
 sg13g2_decap_4 FILLER_54_240 ();
 sg13g2_fill_2 FILLER_54_244 ();
 sg13g2_decap_8 FILLER_54_363 ();
 sg13g2_decap_8 FILLER_54_370 ();
 sg13g2_decap_8 FILLER_54_377 ();
 sg13g2_decap_8 FILLER_54_384 ();
 sg13g2_decap_8 FILLER_54_391 ();
 sg13g2_decap_8 FILLER_54_398 ();
 sg13g2_decap_4 FILLER_54_405 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_4 FILLER_55_21 ();
 sg13g2_fill_1 FILLER_55_25 ();
 sg13g2_decap_4 FILLER_55_89 ();
 sg13g2_fill_2 FILLER_55_106 ();
 sg13g2_fill_1 FILLER_55_108 ();
 sg13g2_decap_4 FILLER_55_163 ();
 sg13g2_fill_1 FILLER_55_167 ();
 sg13g2_fill_2 FILLER_55_241 ();
 sg13g2_fill_1 FILLER_55_243 ();
 sg13g2_decap_8 FILLER_55_368 ();
 sg13g2_decap_8 FILLER_55_375 ();
 sg13g2_decap_8 FILLER_55_382 ();
 sg13g2_decap_8 FILLER_55_389 ();
 sg13g2_decap_8 FILLER_55_396 ();
 sg13g2_decap_4 FILLER_55_403 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_fill_1 FILLER_56_28 ();
 sg13g2_decap_4 FILLER_56_130 ();
 sg13g2_fill_2 FILLER_56_134 ();
 sg13g2_fill_2 FILLER_56_193 ();
 sg13g2_fill_1 FILLER_56_195 ();
 sg13g2_decap_4 FILLER_56_223 ();
 sg13g2_fill_2 FILLER_56_227 ();
 sg13g2_fill_1 FILLER_56_298 ();
 sg13g2_decap_8 FILLER_56_375 ();
 sg13g2_decap_8 FILLER_56_382 ();
 sg13g2_decap_8 FILLER_56_389 ();
 sg13g2_decap_8 FILLER_56_396 ();
 sg13g2_decap_4 FILLER_56_403 ();
 sg13g2_fill_2 FILLER_56_407 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_fill_2 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_113 ();
 sg13g2_fill_2 FILLER_57_187 ();
 sg13g2_fill_1 FILLER_57_189 ();
 sg13g2_decap_8 FILLER_57_213 ();
 sg13g2_fill_1 FILLER_57_220 ();
 sg13g2_fill_2 FILLER_57_302 ();
 sg13g2_decap_8 FILLER_57_384 ();
 sg13g2_decap_8 FILLER_57_391 ();
 sg13g2_decap_8 FILLER_57_398 ();
 sg13g2_decap_4 FILLER_57_405 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_4 FILLER_58_89 ();
 sg13g2_fill_2 FILLER_58_93 ();
 sg13g2_fill_2 FILLER_58_122 ();
 sg13g2_fill_1 FILLER_58_124 ();
 sg13g2_fill_1 FILLER_58_152 ();
 sg13g2_fill_1 FILLER_58_271 ();
 sg13g2_decap_8 FILLER_58_392 ();
 sg13g2_decap_8 FILLER_58_399 ();
 sg13g2_fill_2 FILLER_58_406 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_fill_2 FILLER_59_116 ();
 sg13g2_fill_2 FILLER_59_219 ();
 sg13g2_fill_2 FILLER_59_329 ();
 sg13g2_decap_8 FILLER_59_400 ();
 sg13g2_fill_2 FILLER_59_407 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_fill_1 FILLER_60_35 ();
 sg13g2_fill_2 FILLER_60_100 ();
 sg13g2_decap_4 FILLER_60_115 ();
 sg13g2_fill_2 FILLER_60_119 ();
 sg13g2_decap_8 FILLER_60_161 ();
 sg13g2_fill_2 FILLER_60_232 ();
 sg13g2_fill_1 FILLER_60_234 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_4 FILLER_61_35 ();
 sg13g2_fill_2 FILLER_61_39 ();
 sg13g2_decap_4 FILLER_61_134 ();
 sg13g2_fill_1 FILLER_61_191 ();
 sg13g2_fill_1 FILLER_61_215 ();
 sg13g2_fill_2 FILLER_61_406 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_4 FILLER_62_35 ();
 sg13g2_fill_2 FILLER_62_39 ();
 sg13g2_fill_2 FILLER_62_97 ();
 sg13g2_fill_1 FILLER_62_99 ();
 sg13g2_decap_4 FILLER_62_140 ();
 sg13g2_fill_1 FILLER_62_144 ();
 sg13g2_fill_2 FILLER_62_208 ();
 sg13g2_fill_2 FILLER_62_284 ();
 sg13g2_fill_2 FILLER_62_407 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_fill_2 FILLER_63_49 ();
 sg13g2_fill_1 FILLER_63_51 ();
 sg13g2_fill_2 FILLER_63_126 ();
 sg13g2_fill_1 FILLER_63_128 ();
 sg13g2_fill_2 FILLER_63_209 ();
 sg13g2_fill_1 FILLER_63_211 ();
 sg13g2_fill_1 FILLER_63_252 ();
 sg13g2_fill_2 FILLER_63_406 ();
 sg13g2_fill_1 FILLER_63_408 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_fill_2 FILLER_64_49 ();
 sg13g2_fill_1 FILLER_64_51 ();
 sg13g2_fill_2 FILLER_64_112 ();
 sg13g2_fill_1 FILLER_64_114 ();
 sg13g2_decap_4 FILLER_64_152 ();
 sg13g2_fill_1 FILLER_64_156 ();
 sg13g2_fill_2 FILLER_64_246 ();
 sg13g2_fill_1 FILLER_64_359 ();
 sg13g2_fill_2 FILLER_64_406 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_fill_2 FILLER_65_63 ();
 sg13g2_decap_4 FILLER_65_136 ();
 sg13g2_fill_1 FILLER_65_140 ();
 sg13g2_fill_2 FILLER_65_181 ();
 sg13g2_fill_1 FILLER_65_183 ();
 sg13g2_fill_2 FILLER_65_210 ();
 sg13g2_fill_1 FILLER_65_212 ();
 sg13g2_fill_2 FILLER_65_231 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_fill_2 FILLER_66_125 ();
 sg13g2_fill_1 FILLER_66_127 ();
 sg13g2_decap_4 FILLER_66_155 ();
 sg13g2_fill_2 FILLER_66_172 ();
 sg13g2_fill_1 FILLER_66_174 ();
 sg13g2_fill_2 FILLER_66_198 ();
 sg13g2_fill_1 FILLER_66_200 ();
 sg13g2_fill_1 FILLER_66_224 ();
 sg13g2_fill_2 FILLER_66_407 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_fill_2 FILLER_67_124 ();
 sg13g2_fill_1 FILLER_67_126 ();
 sg13g2_fill_2 FILLER_67_154 ();
 sg13g2_fill_2 FILLER_67_210 ();
 sg13g2_fill_1 FILLER_67_212 ();
 sg13g2_fill_2 FILLER_67_280 ();
 sg13g2_fill_2 FILLER_67_406 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_fill_1 FILLER_68_70 ();
 sg13g2_fill_1 FILLER_68_125 ();
 sg13g2_fill_2 FILLER_68_370 ();
 sg13g2_fill_2 FILLER_68_407 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_fill_2 FILLER_69_247 ();
 sg13g2_fill_1 FILLER_69_344 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_fill_2 FILLER_70_151 ();
 sg13g2_fill_1 FILLER_70_153 ();
 sg13g2_fill_2 FILLER_70_286 ();
 sg13g2_fill_1 FILLER_70_360 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_fill_2 FILLER_71_84 ();
 sg13g2_fill_1 FILLER_71_86 ();
 sg13g2_fill_2 FILLER_71_124 ();
 sg13g2_fill_1 FILLER_71_180 ();
 sg13g2_fill_2 FILLER_71_376 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_4 FILLER_72_84 ();
 sg13g2_fill_2 FILLER_72_249 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_fill_2 FILLER_73_84 ();
 sg13g2_fill_1 FILLER_73_183 ();
 sg13g2_fill_2 FILLER_73_202 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_fill_1 FILLER_74_98 ();
 sg13g2_fill_1 FILLER_74_153 ();
 sg13g2_fill_1 FILLER_74_198 ();
 sg13g2_fill_1 FILLER_74_209 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_fill_2 FILLER_75_98 ();
 sg13g2_fill_1 FILLER_75_162 ();
 sg13g2_fill_2 FILLER_75_341 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_4 FILLER_76_91 ();
 sg13g2_fill_1 FILLER_76_95 ();
 sg13g2_fill_2 FILLER_76_164 ();
 sg13g2_fill_1 FILLER_76_166 ();
 sg13g2_fill_2 FILLER_76_257 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_4 FILLER_77_84 ();
 sg13g2_fill_1 FILLER_77_152 ();
 sg13g2_fill_2 FILLER_77_200 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_fill_2 FILLER_78_77 ();
 sg13g2_fill_1 FILLER_78_79 ();
 sg13g2_fill_1 FILLER_78_152 ();
 sg13g2_fill_2 FILLER_78_190 ();
 sg13g2_fill_1 FILLER_78_192 ();
 sg13g2_fill_2 FILLER_78_310 ();
 sg13g2_fill_2 FILLER_78_407 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_fill_2 FILLER_79_70 ();
 sg13g2_fill_2 FILLER_79_160 ();
 sg13g2_fill_2 FILLER_79_189 ();
 sg13g2_fill_1 FILLER_79_284 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_4 FILLER_80_49 ();
 sg13g2_fill_1 FILLER_80_53 ();
 sg13g2_fill_2 FILLER_80_187 ();
 sg13g2_fill_1 FILLER_80_228 ();
 assign uio_oe[0] = net5;
 assign uio_oe[1] = net6;
 assign uio_oe[2] = net7;
 assign uio_oe[3] = net8;
 assign uio_oe[4] = net9;
 assign uio_oe[5] = net10;
 assign uio_oe[6] = net11;
 assign uio_oe[7] = net12;
 assign uio_out[0] = net13;
 assign uio_out[1] = net14;
 assign uio_out[2] = net15;
 assign uio_out[3] = net16;
 assign uio_out[4] = net17;
 assign uio_out[5] = net18;
 assign uio_out[6] = net19;
 assign uio_out[7] = net20;
 assign uo_out[4] = net21;
 assign uo_out[5] = net22;
 assign uo_out[6] = net23;
 assign uo_out[7] = net24;
endmodule
