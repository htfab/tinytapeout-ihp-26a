module tt_um_algofoogle_fomo (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire clknet_0_clk;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire \h[0] ;
 wire \h[1] ;
 wire \h[2] ;
 wire \h[3] ;
 wire \h[4] ;
 wire \h[5] ;
 wire \h[6] ;
 wire \h[7] ;
 wire \h[8] ;
 wire \h[9] ;
 wire hsync;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire \pix_y[0] ;
 wire \pix_y[1] ;
 wire \pix_y[2] ;
 wire \pix_y[3] ;
 wire \pix_y[4] ;
 wire \pix_y[5] ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire \vx[0] ;
 wire \vx[10] ;
 wire \vx[11] ;
 wire \vx[12] ;
 wire \vx[13] ;
 wire \vx[14] ;
 wire \vx[15] ;
 wire \vx[16] ;
 wire \vx[17] ;
 wire \vx[1] ;
 wire \vx[2] ;
 wire \vx[3] ;
 wire \vx[4] ;
 wire \vx[5] ;
 wire \vx[6] ;
 wire \vx[7] ;
 wire \vx[8] ;
 wire \vx[9] ;
 wire \vy[0] ;
 wire \vy[1] ;
 wire \vy[2] ;
 wire \vy[3] ;
 wire \vy[4] ;
 wire \vy[5] ;
 wire \vy[6] ;
 wire \vy[7] ;
 wire \vy[8] ;
 wire \vy[9] ;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net1;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net39;
 wire net40;
 wire net41;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;

 sg13g2_inv_1 _364_ (.Y(_066_),
    .A(net135));
 sg13g2_inv_1 _365_ (.Y(_067_),
    .A(net145));
 sg13g2_inv_1 _366_ (.Y(_068_),
    .A(net123));
 sg13g2_inv_1 _367_ (.Y(_069_),
    .A(net138));
 sg13g2_inv_1 _368_ (.Y(_070_),
    .A(net51));
 sg13g2_inv_1 _369_ (.Y(_071_),
    .A(\counter[3] ));
 sg13g2_inv_1 _370_ (.Y(_002_),
    .A(\counter[0] ));
 sg13g2_inv_1 _371_ (.Y(_072_),
    .A(net62));
 sg13g2_inv_1 _372_ (.Y(_073_),
    .A(net113));
 sg13g2_inv_1 _373_ (.Y(_074_),
    .A(\counter[7] ));
 sg13g2_inv_1 _374_ (.Y(_075_),
    .A(net149));
 sg13g2_inv_1 _375_ (.Y(_076_),
    .A(net63));
 sg13g2_inv_1 _376_ (.Y(_077_),
    .A(net132));
 sg13g2_nor2_1 _377_ (.A(\counter[2] ),
    .B(\vx[12] ),
    .Y(_078_));
 sg13g2_nor2_1 _378_ (.A(\counter[1] ),
    .B(\vx[11] ),
    .Y(_079_));
 sg13g2_a22oi_1 _379_ (.Y(_080_),
    .B1(\vx[10] ),
    .B2(\counter[0] ),
    .A2(\vx[11] ),
    .A1(\counter[1] ));
 sg13g2_or3_1 _380_ (.A(_078_),
    .B(_079_),
    .C(_080_),
    .X(_081_));
 sg13g2_a22oi_1 _381_ (.Y(_082_),
    .B1(\counter[2] ),
    .B2(\vx[12] ),
    .A2(\vx[13] ),
    .A1(\counter[3] ));
 sg13g2_or2_1 _382_ (.X(_083_),
    .B(\vx[13] ),
    .A(\counter[3] ));
 sg13g2_a22oi_1 _383_ (.Y(_084_),
    .B1(_081_),
    .B2(_082_),
    .A2(_070_),
    .A1(_069_));
 sg13g2_a22oi_1 _384_ (.Y(_085_),
    .B1(_083_),
    .B2(_084_),
    .A2(net51),
    .A1(\vx[14] ));
 sg13g2_nand2_1 _385_ (.Y(_086_),
    .A(net50),
    .B(\vx[15] ));
 sg13g2_nor2_1 _386_ (.A(net50),
    .B(\vx[15] ),
    .Y(_087_));
 sg13g2_xnor2_1 _387_ (.Y(_088_),
    .A(net50),
    .B(\vx[15] ));
 sg13g2_nand4_1 _388_ (.B(net104),
    .C(net115),
    .A(net82),
    .Y(_089_),
    .D(net140));
 sg13g2_nand2_1 _389_ (.Y(_090_),
    .A(\h[7] ),
    .B(net77));
 sg13g2_o21ai_1 _390_ (.B1(net77),
    .Y(_091_),
    .A1(\h[7] ),
    .A2(\h[8] ));
 sg13g2_and3_2 _391_ (.X(_092_),
    .A(_067_),
    .B(_089_),
    .C(_091_));
 sg13g2_nand3_1 _392_ (.B(_089_),
    .C(_091_),
    .A(_067_),
    .Y(_093_));
 sg13g2_o21ai_1 _393_ (.B1(_092_),
    .Y(_094_),
    .A1(_085_),
    .A2(_088_));
 sg13g2_a21oi_1 _394_ (.A1(_085_),
    .A2(_088_),
    .Y(uo_out[0]),
    .B1(_094_));
 sg13g2_nor2_1 _395_ (.A(_072_),
    .B(net49),
    .Y(uo_out[5]));
 sg13g2_and2_1 _396_ (.A(\vx[16] ),
    .B(\counter[6] ),
    .X(_095_));
 sg13g2_xnor2_1 _397_ (.Y(_096_),
    .A(\vx[16] ),
    .B(\counter[6] ));
 sg13g2_a21oi_1 _398_ (.A1(_085_),
    .A2(_086_),
    .Y(_097_),
    .B1(_087_));
 sg13g2_nor2b_1 _399_ (.A(_097_),
    .B_N(_096_),
    .Y(_098_));
 sg13g2_nor2b_1 _400_ (.A(_096_),
    .B_N(_097_),
    .Y(_099_));
 sg13g2_nor3_1 _401_ (.A(net49),
    .B(_098_),
    .C(_099_),
    .Y(uo_out[1]));
 sg13g2_nor2_1 _402_ (.A(_073_),
    .B(net49),
    .Y(uo_out[6]));
 sg13g2_xor2_1 _403_ (.B(\counter[7] ),
    .A(\vx[17] ),
    .X(_100_));
 sg13g2_o21ai_1 _404_ (.B1(_100_),
    .Y(_101_),
    .A1(_095_),
    .A2(_099_));
 sg13g2_or3_1 _405_ (.A(_095_),
    .B(_099_),
    .C(_100_),
    .X(_102_));
 sg13g2_and3_1 _406_ (.X(uo_out[2]),
    .A(_092_),
    .B(_101_),
    .C(_102_));
 sg13g2_nor2_1 _407_ (.A(net145),
    .B(_089_),
    .Y(_103_));
 sg13g2_nor2b_1 _408_ (.A(\hvsync_gen.vpos[2] ),
    .B_N(\hvsync_gen.vpos[3] ),
    .Y(_104_));
 sg13g2_nand4_1 _409_ (.B(_068_),
    .C(_103_),
    .A(net128),
    .Y(_001_),
    .D(_104_));
 sg13g2_nand3_1 _410_ (.B(net135),
    .C(net120),
    .A(net67),
    .Y(_105_));
 sg13g2_nor3_1 _411_ (.A(net67),
    .B(net135),
    .C(net120),
    .Y(_106_));
 sg13g2_nor3_1 _412_ (.A(net125),
    .B(_090_),
    .C(_106_),
    .Y(_107_));
 sg13g2_nand2_1 _413_ (.Y(_000_),
    .A(_105_),
    .B(_107_));
 sg13g2_xor2_1 _414_ (.B(\counter[0] ),
    .A(\counter[1] ),
    .X(_003_));
 sg13g2_nand3_1 _415_ (.B(\counter[1] ),
    .C(\counter[0] ),
    .A(\counter[2] ),
    .Y(_108_));
 sg13g2_a21o_1 _416_ (.A2(\counter[0] ),
    .A1(\counter[1] ),
    .B1(\counter[2] ),
    .X(_109_));
 sg13g2_and2_1 _417_ (.A(_108_),
    .B(_109_),
    .X(_004_));
 sg13g2_nor2_2 _418_ (.A(_071_),
    .B(_108_),
    .Y(_110_));
 sg13g2_xnor2_1 _419_ (.Y(_005_),
    .A(\counter[3] ),
    .B(_108_));
 sg13g2_xnor2_1 _420_ (.Y(_006_),
    .A(_070_),
    .B(_110_));
 sg13g2_nand3_1 _421_ (.B(net51),
    .C(_110_),
    .A(net50),
    .Y(_111_));
 sg13g2_a21o_1 _422_ (.A2(_110_),
    .A1(net51),
    .B1(net50),
    .X(_112_));
 sg13g2_and2_1 _423_ (.A(_111_),
    .B(_112_),
    .X(_007_));
 sg13g2_nand4_1 _424_ (.B(net51),
    .C(\counter[6] ),
    .A(net50),
    .Y(_113_),
    .D(_110_));
 sg13g2_xnor2_1 _425_ (.Y(_008_),
    .A(\counter[6] ),
    .B(_111_));
 sg13g2_nor2_1 _426_ (.A(_074_),
    .B(_113_),
    .Y(_114_));
 sg13g2_xnor2_1 _427_ (.Y(_009_),
    .A(\counter[7] ),
    .B(_113_));
 sg13g2_nand2_1 _428_ (.Y(_115_),
    .A(\counter[8] ),
    .B(_114_));
 sg13g2_xor2_1 _429_ (.B(_114_),
    .A(\counter[8] ),
    .X(_010_));
 sg13g2_xnor2_1 _430_ (.Y(_011_),
    .A(\counter[9] ),
    .B(_115_));
 sg13g2_and3_2 _431_ (.X(_116_),
    .A(net40),
    .B(net79),
    .C(net70));
 sg13g2_nand2_2 _432_ (.Y(_117_),
    .A(net147),
    .B(_116_));
 sg13g2_nor2_2 _433_ (.A(_066_),
    .B(_117_),
    .Y(_118_));
 sg13g2_nor3_1 _434_ (.A(net67),
    .B(\h[7] ),
    .C(net120),
    .Y(_119_));
 sg13g2_nand4_1 _435_ (.B(net125),
    .C(_118_),
    .A(net77),
    .Y(_120_),
    .D(_119_));
 sg13g2_and2_1 _436_ (.A(net55),
    .B(_120_),
    .X(_121_));
 sg13g2_nand2_2 _437_ (.Y(_122_),
    .A(net55),
    .B(_120_));
 sg13g2_nor2_1 _438_ (.A(net40),
    .B(_122_),
    .Y(_012_));
 sg13g2_o21ai_1 _439_ (.B1(_121_),
    .Y(_123_),
    .A1(net40),
    .A2(net79));
 sg13g2_a21oi_1 _440_ (.A1(net40),
    .A2(net79),
    .Y(_013_),
    .B1(_123_));
 sg13g2_a21oi_1 _441_ (.A1(net40),
    .A2(\h[1] ),
    .Y(_124_),
    .B1(net70));
 sg13g2_nor3_1 _442_ (.A(_116_),
    .B(_122_),
    .C(net71),
    .Y(_014_));
 sg13g2_o21ai_1 _443_ (.B1(net55),
    .Y(_125_),
    .A1(net147),
    .A2(_116_));
 sg13g2_nor2b_1 _444_ (.A(_125_),
    .B_N(_117_),
    .Y(_015_));
 sg13g2_o21ai_1 _445_ (.B1(net55),
    .Y(_126_),
    .A1(_066_),
    .A2(_117_));
 sg13g2_a21oi_1 _446_ (.A1(_066_),
    .A2(_117_),
    .Y(_016_),
    .B1(_126_));
 sg13g2_o21ai_1 _447_ (.B1(_121_),
    .Y(_127_),
    .A1(net67),
    .A2(_118_));
 sg13g2_a21oi_1 _448_ (.A1(net67),
    .A2(_118_),
    .Y(_017_),
    .B1(_127_));
 sg13g2_a21oi_1 _449_ (.A1(net67),
    .A2(_118_),
    .Y(_128_),
    .B1(net120));
 sg13g2_nor2_2 _450_ (.A(_105_),
    .B(_117_),
    .Y(_129_));
 sg13g2_nor3_1 _451_ (.A(_122_),
    .B(net121),
    .C(_129_),
    .Y(_018_));
 sg13g2_xnor2_1 _452_ (.Y(_130_),
    .A(net148),
    .B(_129_));
 sg13g2_nor2_1 _453_ (.A(_122_),
    .B(_130_),
    .Y(_019_));
 sg13g2_a21oi_1 _454_ (.A1(\h[7] ),
    .A2(_129_),
    .Y(_131_),
    .B1(net125));
 sg13g2_and3_1 _455_ (.X(_132_),
    .A(\h[7] ),
    .B(net125),
    .C(_129_));
 sg13g2_nor3_1 _456_ (.A(_122_),
    .B(net126),
    .C(_132_),
    .Y(_020_));
 sg13g2_o21ai_1 _457_ (.B1(_121_),
    .Y(_133_),
    .A1(net77),
    .A2(_132_));
 sg13g2_a21oi_1 _458_ (.A1(net77),
    .A2(_132_),
    .Y(_021_),
    .B1(_133_));
 sg13g2_nand2_1 _459_ (.Y(_134_),
    .A(\counter[2] ),
    .B(_092_));
 sg13g2_xnor2_1 _460_ (.Y(_022_),
    .A(net61),
    .B(_134_));
 sg13g2_nand2_1 _461_ (.Y(_135_),
    .A(net91),
    .B(net49));
 sg13g2_and2_1 _462_ (.A(\counter[2] ),
    .B(net61),
    .X(_136_));
 sg13g2_and2_1 _463_ (.A(\counter[3] ),
    .B(net91),
    .X(_137_));
 sg13g2_xor2_1 _464_ (.B(net91),
    .A(\counter[3] ),
    .X(_138_));
 sg13g2_xnor2_1 _465_ (.Y(_139_),
    .A(_136_),
    .B(_138_));
 sg13g2_o21ai_1 _466_ (.B1(_135_),
    .Y(_023_),
    .A1(net49),
    .A2(_139_));
 sg13g2_a21oi_1 _467_ (.A1(_136_),
    .A2(_138_),
    .Y(_140_),
    .B1(_137_));
 sg13g2_nor2_1 _468_ (.A(net51),
    .B(\vx[2] ),
    .Y(_141_));
 sg13g2_xnor2_1 _469_ (.Y(_142_),
    .A(\counter[4] ),
    .B(net101));
 sg13g2_nand2_1 _470_ (.Y(_143_),
    .A(net101),
    .B(net49));
 sg13g2_xnor2_1 _471_ (.Y(_144_),
    .A(_140_),
    .B(_142_));
 sg13g2_o21ai_1 _472_ (.B1(_143_),
    .Y(_024_),
    .A1(net49),
    .A2(_144_));
 sg13g2_nand2_1 _473_ (.Y(_145_),
    .A(\counter[5] ),
    .B(\vx[3] ));
 sg13g2_xor2_1 _474_ (.B(net89),
    .A(\counter[5] ),
    .X(_146_));
 sg13g2_a221oi_1 _475_ (.B2(_138_),
    .C1(_137_),
    .B1(_136_),
    .A1(\counter[4] ),
    .Y(_147_),
    .A2(\vx[2] ));
 sg13g2_nor2_1 _476_ (.A(_141_),
    .B(_147_),
    .Y(_148_));
 sg13g2_nor2_1 _477_ (.A(_146_),
    .B(_148_),
    .Y(_149_));
 sg13g2_nand2b_1 _478_ (.Y(_150_),
    .B(_146_),
    .A_N(_141_));
 sg13g2_or2_1 _479_ (.X(_151_),
    .B(_150_),
    .A(_147_));
 sg13g2_nand2_1 _480_ (.Y(_152_),
    .A(_092_),
    .B(_151_));
 sg13g2_nand2_1 _481_ (.Y(_153_),
    .A(net89),
    .B(net48));
 sg13g2_o21ai_1 _482_ (.B1(_153_),
    .Y(_025_),
    .A1(_149_),
    .A2(_152_));
 sg13g2_nand2_1 _483_ (.Y(_154_),
    .A(\counter[6] ),
    .B(\vx[4] ));
 sg13g2_xnor2_1 _484_ (.Y(_155_),
    .A(\counter[6] ),
    .B(\vx[4] ));
 sg13g2_xnor2_1 _485_ (.Y(_156_),
    .A(_145_),
    .B(_155_));
 sg13g2_o21ai_1 _486_ (.B1(_092_),
    .Y(_157_),
    .A1(_151_),
    .A2(_155_));
 sg13g2_a21oi_1 _487_ (.A1(_151_),
    .A2(_156_),
    .Y(_158_),
    .B1(_157_));
 sg13g2_a21o_1 _488_ (.A2(net48),
    .A1(net133),
    .B1(_158_),
    .X(_026_));
 sg13g2_a21oi_1 _489_ (.A1(_145_),
    .A2(_151_),
    .Y(_159_),
    .B1(_155_));
 sg13g2_nand2_1 _490_ (.Y(_160_),
    .A(\counter[7] ),
    .B(\vx[5] ));
 sg13g2_xor2_1 _491_ (.B(\vx[5] ),
    .A(\counter[7] ),
    .X(_161_));
 sg13g2_xor2_1 _492_ (.B(_161_),
    .A(_154_),
    .X(_162_));
 sg13g2_xnor2_1 _493_ (.Y(_163_),
    .A(_159_),
    .B(_162_));
 sg13g2_mux2_1 _494_ (.A0(net141),
    .A1(_163_),
    .S(_092_),
    .X(_027_));
 sg13g2_nor2_1 _495_ (.A(\counter[8] ),
    .B(\vx[6] ),
    .Y(_164_));
 sg13g2_xnor2_1 _496_ (.Y(_165_),
    .A(\counter[8] ),
    .B(\vx[6] ));
 sg13g2_nor2b_1 _497_ (.A(_160_),
    .B_N(_165_),
    .Y(_166_));
 sg13g2_nand2b_1 _498_ (.Y(_167_),
    .B(_165_),
    .A_N(_160_));
 sg13g2_nand2b_1 _499_ (.Y(_168_),
    .B(_160_),
    .A_N(_165_));
 sg13g2_nand2_1 _500_ (.Y(_169_),
    .A(_167_),
    .B(_168_));
 sg13g2_or4_1 _501_ (.A(_147_),
    .B(_150_),
    .C(_156_),
    .D(_162_),
    .X(_170_));
 sg13g2_o21ai_1 _502_ (.B1(_154_),
    .Y(_171_),
    .A1(_145_),
    .A2(_155_));
 sg13g2_nand2_1 _503_ (.Y(_172_),
    .A(_161_),
    .B(_171_));
 sg13g2_and2_1 _504_ (.A(_170_),
    .B(_172_),
    .X(_173_));
 sg13g2_xnor2_1 _505_ (.Y(_174_),
    .A(_169_),
    .B(_173_));
 sg13g2_nand2_1 _506_ (.Y(_175_),
    .A(net103),
    .B(net48));
 sg13g2_o21ai_1 _507_ (.B1(_175_),
    .Y(_028_),
    .A1(net48),
    .A2(_174_));
 sg13g2_or2_1 _508_ (.X(_176_),
    .B(\vx[7] ),
    .A(\counter[9] ));
 sg13g2_nand2_1 _509_ (.Y(_177_),
    .A(\counter[9] ),
    .B(\vx[7] ));
 sg13g2_a21oi_1 _510_ (.A1(_176_),
    .A2(_177_),
    .Y(_178_),
    .B1(_164_));
 sg13g2_a21o_1 _511_ (.A2(_177_),
    .A1(_176_),
    .B1(_164_),
    .X(_179_));
 sg13g2_nand3_1 _512_ (.B(_176_),
    .C(_177_),
    .A(_164_),
    .Y(_180_));
 sg13g2_nand2_1 _513_ (.Y(_181_),
    .A(_179_),
    .B(_180_));
 sg13g2_o21ai_1 _514_ (.B1(_167_),
    .Y(_182_),
    .A1(_169_),
    .A2(_173_));
 sg13g2_xor2_1 _515_ (.B(_182_),
    .A(_181_),
    .X(_183_));
 sg13g2_nand2_1 _516_ (.Y(_184_),
    .A(net80),
    .B(net48));
 sg13g2_o21ai_1 _517_ (.B1(_184_),
    .Y(_029_),
    .A1(_093_),
    .A2(_183_));
 sg13g2_a221oi_1 _518_ (.B2(_166_),
    .C1(_178_),
    .B1(_180_),
    .A1(_161_),
    .Y(_185_),
    .A2(_171_));
 sg13g2_nand2_1 _519_ (.Y(_186_),
    .A(_168_),
    .B(_180_));
 sg13g2_a22oi_1 _520_ (.Y(_187_),
    .B1(_186_),
    .B2(_179_),
    .A2(_185_),
    .A1(_170_));
 sg13g2_nand2_1 _521_ (.Y(_188_),
    .A(\vx[8] ),
    .B(_176_));
 sg13g2_xnor2_1 _522_ (.Y(_189_),
    .A(_077_),
    .B(_176_));
 sg13g2_a21oi_1 _523_ (.A1(_187_),
    .A2(_189_),
    .Y(_190_),
    .B1(_093_));
 sg13g2_o21ai_1 _524_ (.B1(_190_),
    .Y(_191_),
    .A1(_187_),
    .A2(_189_));
 sg13g2_o21ai_1 _525_ (.B1(_191_),
    .Y(_030_),
    .A1(_077_),
    .A2(_092_));
 sg13g2_nand2_1 _526_ (.Y(_192_),
    .A(_188_),
    .B(_190_));
 sg13g2_xnor2_1 _527_ (.Y(_031_),
    .A(net106),
    .B(_192_));
 sg13g2_nand2_1 _528_ (.Y(_193_),
    .A(net130),
    .B(net48));
 sg13g2_and2_1 _529_ (.A(\vx[10] ),
    .B(net106),
    .X(_194_));
 sg13g2_xnor2_1 _530_ (.Y(_195_),
    .A(net130),
    .B(net106));
 sg13g2_inv_1 _531_ (.Y(_196_),
    .A(_195_));
 sg13g2_nor2b_1 _532_ (.A(\vx[9] ),
    .B_N(_189_),
    .Y(_197_));
 sg13g2_nand2_1 _533_ (.Y(_198_),
    .A(_187_),
    .B(_197_));
 sg13g2_or2_1 _534_ (.X(_199_),
    .B(_188_),
    .A(\vx[9] ));
 sg13g2_nand2_1 _535_ (.Y(_200_),
    .A(_198_),
    .B(_199_));
 sg13g2_a21oi_1 _536_ (.A1(_198_),
    .A2(_199_),
    .Y(_201_),
    .B1(_195_));
 sg13g2_xnor2_1 _537_ (.Y(_202_),
    .A(_196_),
    .B(_200_));
 sg13g2_o21ai_1 _538_ (.B1(_193_),
    .Y(_032_),
    .A1(net48),
    .A2(_202_));
 sg13g2_o21ai_1 _539_ (.B1(_092_),
    .Y(_203_),
    .A1(_194_),
    .A2(_201_));
 sg13g2_nand4_1 _540_ (.B(_187_),
    .C(_196_),
    .A(\vx[11] ),
    .Y(_204_),
    .D(_197_));
 sg13g2_nand2b_1 _541_ (.Y(_205_),
    .B(_188_),
    .A_N(\vx[9] ));
 sg13g2_nand3_1 _542_ (.B(\vx[10] ),
    .C(_205_),
    .A(\vx[11] ),
    .Y(_206_));
 sg13g2_a21oi_2 _543_ (.B1(net48),
    .Y(_207_),
    .A2(_206_),
    .A1(_204_));
 sg13g2_xnor2_1 _544_ (.Y(_033_),
    .A(net117),
    .B(_203_));
 sg13g2_xor2_1 _545_ (.B(net42),
    .A(net73),
    .X(_034_));
 sg13g2_and2_1 _546_ (.A(net88),
    .B(net73),
    .X(_208_));
 sg13g2_nand2_1 _547_ (.Y(_209_),
    .A(net42),
    .B(_208_));
 sg13g2_a21oi_1 _548_ (.A1(net73),
    .A2(net42),
    .Y(_210_),
    .B1(net88));
 sg13g2_a21oi_1 _549_ (.A1(net42),
    .A2(_208_),
    .Y(_035_),
    .B1(_210_));
 sg13g2_and2_1 _550_ (.A(net138),
    .B(_208_),
    .X(_211_));
 sg13g2_a22oi_1 _551_ (.Y(_036_),
    .B1(_211_),
    .B2(net42),
    .A2(_209_),
    .A1(_069_));
 sg13g2_and2_1 _552_ (.A(net110),
    .B(_211_),
    .X(_212_));
 sg13g2_a21oi_1 _553_ (.A1(net42),
    .A2(_211_),
    .Y(_213_),
    .B1(net110));
 sg13g2_a21oi_1 _554_ (.A1(net42),
    .A2(_212_),
    .Y(_037_),
    .B1(net111));
 sg13g2_and2_1 _555_ (.A(net85),
    .B(_212_),
    .X(_214_));
 sg13g2_nand2_1 _556_ (.Y(_215_),
    .A(net42),
    .B(_214_));
 sg13g2_a21oi_1 _557_ (.A1(_207_),
    .A2(_212_),
    .Y(_216_),
    .B1(net85));
 sg13g2_a21oi_1 _558_ (.A1(_207_),
    .A2(_214_),
    .Y(_038_),
    .B1(net86));
 sg13g2_xnor2_1 _559_ (.Y(_039_),
    .A(net75),
    .B(_215_));
 sg13g2_nor3_1 _560_ (.A(\h[7] ),
    .B(\h[9] ),
    .C(\h[8] ),
    .Y(_217_));
 sg13g2_nor4_1 _561_ (.A(\h[0] ),
    .B(\h[1] ),
    .C(\h[3] ),
    .D(\h[2] ),
    .Y(_218_));
 sg13g2_nand3_1 _562_ (.B(_217_),
    .C(_218_),
    .A(_106_),
    .Y(_219_));
 sg13g2_inv_2 _563_ (.Y(_220_),
    .A(net46));
 sg13g2_nor2_1 _564_ (.A(_002_),
    .B(net47),
    .Y(_221_));
 sg13g2_xor2_1 _565_ (.B(_221_),
    .A(net39),
    .X(_040_));
 sg13g2_nand2_1 _566_ (.Y(_222_),
    .A(\counter[0] ),
    .B(net39));
 sg13g2_nand2_1 _567_ (.Y(_223_),
    .A(\counter[1] ),
    .B(\vy[1] ));
 sg13g2_xnor2_1 _568_ (.Y(_224_),
    .A(\counter[1] ),
    .B(net108));
 sg13g2_xnor2_1 _569_ (.Y(_225_),
    .A(_222_),
    .B(_224_));
 sg13g2_nand2_1 _570_ (.Y(_226_),
    .A(net108),
    .B(net47));
 sg13g2_o21ai_1 _571_ (.B1(_226_),
    .Y(_041_),
    .A1(net47),
    .A2(_225_));
 sg13g2_and2_1 _572_ (.A(\counter[2] ),
    .B(\vy[2] ),
    .X(_227_));
 sg13g2_xor2_1 _573_ (.B(net93),
    .A(\counter[2] ),
    .X(_228_));
 sg13g2_o21ai_1 _574_ (.B1(_223_),
    .Y(_229_),
    .A1(_222_),
    .A2(_224_));
 sg13g2_xnor2_1 _575_ (.Y(_230_),
    .A(_228_),
    .B(_229_));
 sg13g2_nand2_1 _576_ (.Y(_231_),
    .A(net93),
    .B(net47));
 sg13g2_o21ai_1 _577_ (.B1(_231_),
    .Y(_042_),
    .A1(net47),
    .A2(_230_));
 sg13g2_nand2_1 _578_ (.Y(_232_),
    .A(\counter[3] ),
    .B(\vy[3] ));
 sg13g2_xor2_1 _579_ (.B(\vy[3] ),
    .A(\counter[3] ),
    .X(_233_));
 sg13g2_a21o_2 _580_ (.A2(_229_),
    .A1(_228_),
    .B1(_227_),
    .X(_234_));
 sg13g2_nand2_1 _581_ (.Y(_235_),
    .A(_233_),
    .B(_234_));
 sg13g2_xor2_1 _582_ (.B(_234_),
    .A(_233_),
    .X(_236_));
 sg13g2_mux2_1 _583_ (.A0(net139),
    .A1(_236_),
    .S(_220_),
    .X(_043_));
 sg13g2_or2_1 _584_ (.X(_237_),
    .B(\vy[4] ),
    .A(net51));
 sg13g2_xnor2_1 _585_ (.Y(_238_),
    .A(net51),
    .B(\vy[4] ));
 sg13g2_nand2b_1 _586_ (.Y(_239_),
    .B(_238_),
    .A_N(_232_));
 sg13g2_xor2_1 _587_ (.B(_238_),
    .A(_232_),
    .X(_240_));
 sg13g2_nand3_1 _588_ (.B(_234_),
    .C(_238_),
    .A(_233_),
    .Y(_241_));
 sg13g2_a21oi_1 _589_ (.A1(_235_),
    .A2(_240_),
    .Y(_242_),
    .B1(net47));
 sg13g2_a22oi_1 _590_ (.Y(_243_),
    .B1(_241_),
    .B2(_242_),
    .A2(net47),
    .A1(net137));
 sg13g2_inv_1 _591_ (.Y(_044_),
    .A(_243_));
 sg13g2_nand2_1 _592_ (.Y(_244_),
    .A(net50),
    .B(\vy[5] ));
 sg13g2_xor2_1 _593_ (.B(\vy[5] ),
    .A(net50),
    .X(_245_));
 sg13g2_nor2_1 _594_ (.A(_237_),
    .B(_245_),
    .Y(_246_));
 sg13g2_nand2_1 _595_ (.Y(_247_),
    .A(_237_),
    .B(_245_));
 sg13g2_nor2b_2 _596_ (.A(_246_),
    .B_N(_247_),
    .Y(_248_));
 sg13g2_nand2_1 _597_ (.Y(_249_),
    .A(_239_),
    .B(_241_));
 sg13g2_xnor2_1 _598_ (.Y(_250_),
    .A(_248_),
    .B(_249_));
 sg13g2_nand2_1 _599_ (.Y(_251_),
    .A(net99),
    .B(net45));
 sg13g2_o21ai_1 _600_ (.B1(_251_),
    .Y(_045_),
    .A1(net45),
    .A2(_250_));
 sg13g2_nand2_1 _601_ (.Y(_252_),
    .A(net92),
    .B(net45));
 sg13g2_nor2_1 _602_ (.A(\counter[6] ),
    .B(\vy[6] ),
    .Y(_253_));
 sg13g2_xnor2_1 _603_ (.Y(_254_),
    .A(\counter[6] ),
    .B(\vy[6] ));
 sg13g2_nor2b_1 _604_ (.A(_244_),
    .B_N(_254_),
    .Y(_255_));
 sg13g2_xor2_1 _605_ (.B(_254_),
    .A(_244_),
    .X(_256_));
 sg13g2_nor2_1 _606_ (.A(_239_),
    .B(_246_),
    .Y(_257_));
 sg13g2_a21oi_1 _607_ (.A1(_237_),
    .A2(_245_),
    .Y(_258_),
    .B1(_257_));
 sg13g2_o21ai_1 _608_ (.B1(_247_),
    .Y(_259_),
    .A1(_239_),
    .A2(_246_));
 sg13g2_nand4_1 _609_ (.B(_234_),
    .C(_238_),
    .A(_233_),
    .Y(_260_),
    .D(_248_));
 sg13g2_nand3_1 _610_ (.B(_258_),
    .C(_260_),
    .A(_256_),
    .Y(_261_));
 sg13g2_a21oi_1 _611_ (.A1(_258_),
    .A2(_260_),
    .Y(_262_),
    .B1(_256_));
 sg13g2_nand2_1 _612_ (.Y(_263_),
    .A(_220_),
    .B(_261_));
 sg13g2_o21ai_1 _613_ (.B1(_252_),
    .Y(_046_),
    .A1(_262_),
    .A2(_263_));
 sg13g2_nor2_1 _614_ (.A(\counter[7] ),
    .B(net95),
    .Y(_264_));
 sg13g2_xor2_1 _615_ (.B(\vy[7] ),
    .A(\counter[7] ),
    .X(_265_));
 sg13g2_nor2_1 _616_ (.A(_253_),
    .B(_265_),
    .Y(_266_));
 sg13g2_nand2_1 _617_ (.Y(_267_),
    .A(_253_),
    .B(_265_));
 sg13g2_xnor2_1 _618_ (.Y(_268_),
    .A(_253_),
    .B(_265_));
 sg13g2_nor2_1 _619_ (.A(_255_),
    .B(_262_),
    .Y(_269_));
 sg13g2_xnor2_1 _620_ (.Y(_270_),
    .A(_268_),
    .B(_269_));
 sg13g2_nand2_1 _621_ (.Y(_271_),
    .A(net95),
    .B(net45));
 sg13g2_o21ai_1 _622_ (.B1(_271_),
    .Y(_047_),
    .A1(net45),
    .A2(_270_));
 sg13g2_nor2_1 _623_ (.A(_256_),
    .B(_268_),
    .Y(_272_));
 sg13g2_nor3_1 _624_ (.A(_240_),
    .B(_256_),
    .C(_268_),
    .Y(_273_));
 sg13g2_nand4_1 _625_ (.B(_234_),
    .C(_248_),
    .A(_233_),
    .Y(_274_),
    .D(_273_));
 sg13g2_or2_1 _626_ (.X(_275_),
    .B(_266_),
    .A(_255_));
 sg13g2_a22oi_1 _627_ (.Y(_276_),
    .B1(_275_),
    .B2(_267_),
    .A2(_272_),
    .A1(_259_));
 sg13g2_nand2_1 _628_ (.Y(_277_),
    .A(_274_),
    .B(_276_));
 sg13g2_nand2_1 _629_ (.Y(_278_),
    .A(net97),
    .B(\counter[8] ));
 sg13g2_xor2_1 _630_ (.B(\counter[8] ),
    .A(\vy[8] ),
    .X(_279_));
 sg13g2_nor2b_1 _631_ (.A(_264_),
    .B_N(_279_),
    .Y(_280_));
 sg13g2_nand2b_1 _632_ (.Y(_281_),
    .B(_279_),
    .A_N(_264_));
 sg13g2_xnor2_1 _633_ (.Y(_282_),
    .A(_264_),
    .B(_279_));
 sg13g2_xnor2_1 _634_ (.Y(_283_),
    .A(_277_),
    .B(_282_));
 sg13g2_nand2_1 _635_ (.Y(_284_),
    .A(net97),
    .B(net45));
 sg13g2_o21ai_1 _636_ (.B1(_284_),
    .Y(_048_),
    .A1(net45),
    .A2(_283_));
 sg13g2_a21oi_1 _637_ (.A1(_277_),
    .A2(_282_),
    .Y(_285_),
    .B1(_280_));
 sg13g2_xor2_1 _638_ (.B(\counter[9] ),
    .A(\vy[9] ),
    .X(_286_));
 sg13g2_xnor2_1 _639_ (.Y(_287_),
    .A(_278_),
    .B(_286_));
 sg13g2_xnor2_1 _640_ (.Y(_288_),
    .A(_285_),
    .B(_287_));
 sg13g2_nand2_1 _641_ (.Y(_289_),
    .A(net102),
    .B(net45));
 sg13g2_o21ai_1 _642_ (.B1(_289_),
    .Y(_049_),
    .A1(net46),
    .A2(_288_));
 sg13g2_o21ai_1 _643_ (.B1(\pix_y[0] ),
    .Y(_290_),
    .A1(\vy[9] ),
    .A2(\counter[9] ));
 sg13g2_inv_1 _644_ (.Y(_291_),
    .A(_290_));
 sg13g2_or3_1 _645_ (.A(\vy[9] ),
    .B(\counter[9] ),
    .C(\pix_y[0] ),
    .X(_292_));
 sg13g2_and2_1 _646_ (.A(_290_),
    .B(_292_),
    .X(_293_));
 sg13g2_nor2b_1 _647_ (.A(_287_),
    .B_N(_282_),
    .Y(_294_));
 sg13g2_inv_1 _648_ (.Y(_295_),
    .A(_294_));
 sg13g2_a21oi_1 _649_ (.A1(_274_),
    .A2(_276_),
    .Y(_296_),
    .B1(_295_));
 sg13g2_a21oi_1 _650_ (.A1(_278_),
    .A2(_281_),
    .Y(_297_),
    .B1(_286_));
 sg13g2_nor3_1 _651_ (.A(_293_),
    .B(_296_),
    .C(_297_),
    .Y(_298_));
 sg13g2_o21ai_1 _652_ (.B1(_293_),
    .Y(_299_),
    .A1(_296_),
    .A2(_297_));
 sg13g2_nand2_1 _653_ (.Y(_300_),
    .A(_220_),
    .B(_299_));
 sg13g2_nand2_1 _654_ (.Y(_301_),
    .A(net69),
    .B(net46));
 sg13g2_o21ai_1 _655_ (.B1(_301_),
    .Y(_050_),
    .A1(_298_),
    .A2(_300_));
 sg13g2_a21oi_1 _656_ (.A1(_290_),
    .A2(_299_),
    .Y(_302_),
    .B1(net46));
 sg13g2_nand3_1 _657_ (.B(_293_),
    .C(_294_),
    .A(\pix_y[1] ),
    .Y(_303_));
 sg13g2_a21oi_1 _658_ (.A1(_274_),
    .A2(_276_),
    .Y(_304_),
    .B1(_303_));
 sg13g2_o21ai_1 _659_ (.B1(\pix_y[1] ),
    .Y(_305_),
    .A1(_291_),
    .A2(_297_));
 sg13g2_nor2b_1 _660_ (.A(_305_),
    .B_N(_292_),
    .Y(_306_));
 sg13g2_o21ai_1 _661_ (.B1(_220_),
    .Y(_307_),
    .A1(_304_),
    .A2(_306_));
 sg13g2_xor2_1 _662_ (.B(_302_),
    .A(net65),
    .X(_051_));
 sg13g2_xnor2_1 _663_ (.Y(_052_),
    .A(net62),
    .B(_307_));
 sg13g2_or3_1 _664_ (.A(_072_),
    .B(_075_),
    .C(_307_),
    .X(_308_));
 sg13g2_o21ai_1 _665_ (.B1(_075_),
    .Y(_309_),
    .A1(_072_),
    .A2(_307_));
 sg13g2_and2_1 _666_ (.A(_308_),
    .B(_309_),
    .X(_053_));
 sg13g2_nor4_1 _667_ (.A(_072_),
    .B(_075_),
    .C(_076_),
    .D(_307_),
    .Y(_310_));
 sg13g2_xnor2_1 _668_ (.Y(_054_),
    .A(net63),
    .B(_308_));
 sg13g2_xnor2_1 _669_ (.Y(_055_),
    .A(_073_),
    .B(_310_));
 sg13g2_or4_1 _670_ (.A(\hvsync_gen.vpos[0] ),
    .B(\hvsync_gen.vpos[8] ),
    .C(\hvsync_gen.vpos[5] ),
    .D(\hvsync_gen.vpos[1] ),
    .X(_311_));
 sg13g2_nand4_1 _671_ (.B(\hvsync_gen.vpos[3] ),
    .C(\hvsync_gen.vpos[2] ),
    .A(\hvsync_gen.vpos[9] ),
    .Y(_312_),
    .D(_068_));
 sg13g2_nor4_1 _672_ (.A(\hvsync_gen.vpos[7] ),
    .B(\hvsync_gen.vpos[6] ),
    .C(_311_),
    .D(_312_),
    .Y(_313_));
 sg13g2_nand2b_1 _673_ (.Y(_314_),
    .B(net55),
    .A_N(_313_));
 sg13g2_nor2_2 _674_ (.A(_120_),
    .B(_314_),
    .Y(_315_));
 sg13g2_nor2_1 _675_ (.A(net119),
    .B(net43),
    .Y(_316_));
 sg13g2_a21oi_1 _676_ (.A1(net119),
    .A2(_122_),
    .Y(_056_),
    .B1(_316_));
 sg13g2_xor2_1 _677_ (.B(net128),
    .A(net119),
    .X(_317_));
 sg13g2_a22oi_1 _678_ (.Y(_318_),
    .B1(net43),
    .B2(_317_),
    .A2(net44),
    .A1(net128));
 sg13g2_inv_1 _679_ (.Y(_057_),
    .A(_318_));
 sg13g2_a21oi_1 _680_ (.A1(net119),
    .A2(net128),
    .Y(_319_),
    .B1(net144));
 sg13g2_nand3_1 _681_ (.B(net128),
    .C(net144),
    .A(net119),
    .Y(_320_));
 sg13g2_nor2b_1 _682_ (.A(_319_),
    .B_N(_320_),
    .Y(_321_));
 sg13g2_a22oi_1 _683_ (.Y(_322_),
    .B1(net43),
    .B2(_321_),
    .A2(net44),
    .A1(net144));
 sg13g2_inv_1 _684_ (.Y(_058_),
    .A(_322_));
 sg13g2_and4_1 _685_ (.A(net119),
    .B(\hvsync_gen.vpos[1] ),
    .C(\hvsync_gen.vpos[3] ),
    .D(\hvsync_gen.vpos[2] ),
    .X(_323_));
 sg13g2_xnor2_1 _686_ (.Y(_324_),
    .A(net142),
    .B(_320_));
 sg13g2_a22oi_1 _687_ (.Y(_325_),
    .B1(net43),
    .B2(_324_),
    .A2(net44),
    .A1(net142));
 sg13g2_inv_1 _688_ (.Y(_059_),
    .A(net143));
 sg13g2_and2_1 _689_ (.A(net123),
    .B(_323_),
    .X(_326_));
 sg13g2_xnor2_1 _690_ (.Y(_327_),
    .A(_068_),
    .B(_323_));
 sg13g2_a22oi_1 _691_ (.Y(_328_),
    .B1(net43),
    .B2(_327_),
    .A2(net44),
    .A1(net123));
 sg13g2_inv_1 _692_ (.Y(_060_),
    .A(net124));
 sg13g2_and2_1 _693_ (.A(\hvsync_gen.vpos[5] ),
    .B(_326_),
    .X(_329_));
 sg13g2_xor2_1 _694_ (.B(_326_),
    .A(net140),
    .X(_330_));
 sg13g2_a22oi_1 _695_ (.Y(_331_),
    .B1(net43),
    .B2(_330_),
    .A2(net44),
    .A1(net140));
 sg13g2_inv_1 _696_ (.Y(_061_),
    .A(_331_));
 sg13g2_nand2_1 _697_ (.Y(_332_),
    .A(net115),
    .B(net44));
 sg13g2_and2_1 _698_ (.A(net115),
    .B(_329_),
    .X(_333_));
 sg13g2_o21ai_1 _699_ (.B1(net43),
    .Y(_334_),
    .A1(net115),
    .A2(_329_));
 sg13g2_o21ai_1 _700_ (.B1(_332_),
    .Y(_062_),
    .A1(_333_),
    .A2(_334_));
 sg13g2_nand2_1 _701_ (.Y(_335_),
    .A(net104),
    .B(net44));
 sg13g2_and2_1 _702_ (.A(net104),
    .B(_333_),
    .X(_336_));
 sg13g2_o21ai_1 _703_ (.B1(net43),
    .Y(_337_),
    .A1(net104),
    .A2(_333_));
 sg13g2_o21ai_1 _704_ (.B1(_335_),
    .Y(_063_),
    .A1(_336_),
    .A2(_337_));
 sg13g2_a21oi_1 _705_ (.A1(net82),
    .A2(_336_),
    .Y(_338_),
    .B1(_314_));
 sg13g2_nor2_1 _706_ (.A(net44),
    .B(_338_),
    .Y(_339_));
 sg13g2_a21oi_1 _707_ (.A1(_315_),
    .A2(_336_),
    .Y(_340_),
    .B1(net82));
 sg13g2_nor2_1 _708_ (.A(_339_),
    .B(net83),
    .Y(_064_));
 sg13g2_nand3_1 _709_ (.B(_315_),
    .C(_326_),
    .A(_103_),
    .Y(_341_));
 sg13g2_o21ai_1 _710_ (.B1(_341_),
    .Y(_065_),
    .A1(_067_),
    .A2(_339_));
 sg13g2_dfrbpq_2 _711_ (.RESET_B(net22),
    .D(net41),
    .Q(\h[0] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _712_ (.RESET_B(net31),
    .D(_013_),
    .Q(\h[1] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _713_ (.RESET_B(net30),
    .D(net72),
    .Q(\h[2] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _714_ (.RESET_B(net29),
    .D(_015_),
    .Q(\h[3] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _715_ (.RESET_B(net28),
    .D(_016_),
    .Q(\h[4] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _716_ (.RESET_B(net27),
    .D(net68),
    .Q(\h[5] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _717_ (.RESET_B(net26),
    .D(net122),
    .Q(\h[6] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_2 _718_ (.RESET_B(net25),
    .D(_019_),
    .Q(\h[7] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _719_ (.RESET_B(net24),
    .D(net127),
    .Q(\h[8] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _720_ (.RESET_B(net23),
    .D(net78),
    .Q(\h[9] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _721_ (.RESET_B(net54),
    .D(_022_),
    .Q(\vx[0] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _722_ (.RESET_B(net57),
    .D(_023_),
    .Q(\vx[1] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_2 _723_ (.RESET_B(net57),
    .D(_024_),
    .Q(\vx[2] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_1 _724_ (.RESET_B(net56),
    .D(net90),
    .Q(\vx[3] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_1 _725_ (.RESET_B(net57),
    .D(net134),
    .Q(\vx[4] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_1 _726_ (.RESET_B(net59),
    .D(_027_),
    .Q(\vx[5] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_1 _727_ (.RESET_B(net59),
    .D(_028_),
    .Q(\vx[6] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_1 _728_ (.RESET_B(net59),
    .D(net81),
    .Q(\vx[7] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_1 _729_ (.RESET_B(net59),
    .D(_030_),
    .Q(\vx[8] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_2 _730_ (.RESET_B(net59),
    .D(net107),
    .Q(\vx[9] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_2 _731_ (.RESET_B(net59),
    .D(net131),
    .Q(\vx[10] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_2 _732_ (.RESET_B(net57),
    .D(net118),
    .Q(\vx[11] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_2 _733_ (.RESET_B(net54),
    .D(net74),
    .Q(\vx[12] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _734_ (.RESET_B(net54),
    .D(_035_),
    .Q(\vx[13] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _735_ (.RESET_B(net53),
    .D(_036_),
    .Q(\vx[14] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _736_ (.RESET_B(net54),
    .D(net112),
    .Q(\vx[15] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_2 _737_ (.RESET_B(net57),
    .D(net87),
    .Q(\vx[16] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _738_ (.RESET_B(net57),
    .D(net76),
    .Q(\vx[17] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_2 _739_ (.RESET_B(net53),
    .D(_002_),
    .Q(\counter[0] ),
    .CLK(net52));
 sg13g2_dfrbpq_2 _740_ (.RESET_B(net53),
    .D(_003_),
    .Q(\counter[1] ),
    .CLK(net52));
 sg13g2_dfrbpq_2 _741_ (.RESET_B(net53),
    .D(_004_),
    .Q(\counter[2] ),
    .CLK(net52));
 sg13g2_dfrbpq_2 _742_ (.RESET_B(net53),
    .D(_005_),
    .Q(\counter[3] ),
    .CLK(net52));
 sg13g2_dfrbpq_2 _743_ (.RESET_B(net56),
    .D(_006_),
    .Q(\counter[4] ),
    .CLK(net52));
 sg13g2_dfrbpq_2 _744_ (.RESET_B(net56),
    .D(_007_),
    .Q(\counter[5] ),
    .CLK(net52));
 sg13g2_dfrbpq_2 _745_ (.RESET_B(net56),
    .D(_008_),
    .Q(\counter[6] ),
    .CLK(net52));
 sg13g2_dfrbpq_2 _746_ (.RESET_B(net58),
    .D(_009_),
    .Q(\counter[7] ),
    .CLK(\hvsync_gen.vsync ));
 sg13g2_dfrbpq_2 _747_ (.RESET_B(net58),
    .D(_010_),
    .Q(\counter[8] ),
    .CLK(\hvsync_gen.vsync ));
 sg13g2_dfrbpq_2 _748_ (.RESET_B(net58),
    .D(_011_),
    .Q(\counter[9] ),
    .CLK(\hvsync_gen.vsync ));
 sg13g2_dfrbpq_1 _749_ (.RESET_B(net53),
    .D(_040_),
    .Q(\vy[0] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_1 _750_ (.RESET_B(net53),
    .D(net109),
    .Q(\vy[1] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_1 _751_ (.RESET_B(net53),
    .D(net94),
    .Q(\vy[2] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_1 _752_ (.RESET_B(net56),
    .D(_043_),
    .Q(\vy[3] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_1 _753_ (.RESET_B(net56),
    .D(_044_),
    .Q(\vy[4] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_1 _754_ (.RESET_B(net56),
    .D(net100),
    .Q(\vy[5] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_1 _755_ (.RESET_B(net56),
    .D(_046_),
    .Q(\vy[6] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_1 _756_ (.RESET_B(net58),
    .D(net96),
    .Q(\vy[7] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_1 _757_ (.RESET_B(net58),
    .D(net98),
    .Q(\vy[8] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_2 _758_ (.RESET_B(net58),
    .D(_049_),
    .Q(\vy[9] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_1 _759_ (.RESET_B(net58),
    .D(_050_),
    .Q(\pix_y[0] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_1 _760_ (.RESET_B(net58),
    .D(net66),
    .Q(\pix_y[1] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_1 _761_ (.RESET_B(net54),
    .D(_052_),
    .Q(\pix_y[2] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _762_ (.RESET_B(net54),
    .D(_053_),
    .Q(\pix_y[3] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _763_ (.RESET_B(net55),
    .D(net64),
    .Q(\pix_y[4] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _764_ (.RESET_B(net54),
    .D(net114),
    .Q(\pix_y[5] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _765_ (.RESET_B(net21),
    .D(net136),
    .Q(hsync),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_2 _766_ (.RESET_B(net20),
    .D(_056_),
    .Q(\hvsync_gen.vpos[0] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _767_ (.RESET_B(net18),
    .D(_057_),
    .Q(\hvsync_gen.vpos[1] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _768_ (.RESET_B(net38),
    .D(_058_),
    .Q(\hvsync_gen.vpos[2] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _769_ (.RESET_B(net36),
    .D(_059_),
    .Q(\hvsync_gen.vpos[3] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_1 _770_ (.RESET_B(net34),
    .D(_060_),
    .Q(\hvsync_gen.vpos[4] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _771_ (.RESET_B(net32),
    .D(_061_),
    .Q(\hvsync_gen.vpos[5] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _772_ (.RESET_B(net17),
    .D(net116),
    .Q(\hvsync_gen.vpos[6] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _773_ (.RESET_B(net35),
    .D(net105),
    .Q(\hvsync_gen.vpos[7] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_2 _774_ (.RESET_B(net19),
    .D(net84),
    .Q(\hvsync_gen.vpos[8] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_1 _775_ (.RESET_B(net37),
    .D(net146),
    .Q(\hvsync_gen.vpos[9] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_2 _776_ (.RESET_B(net33),
    .D(net129),
    .Q(\hvsync_gen.vsync ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_tiehi _767__18 (.L_HI(net18));
 sg13g2_tiehi _774__19 (.L_HI(net19));
 sg13g2_tiehi _766__20 (.L_HI(net20));
 sg13g2_tiehi _765__21 (.L_HI(net21));
 sg13g2_tiehi _711__22 (.L_HI(net22));
 sg13g2_tiehi _720__23 (.L_HI(net23));
 sg13g2_tiehi _719__24 (.L_HI(net24));
 sg13g2_tiehi _718__25 (.L_HI(net25));
 sg13g2_tiehi _717__26 (.L_HI(net26));
 sg13g2_tiehi _716__27 (.L_HI(net27));
 sg13g2_tiehi _715__28 (.L_HI(net28));
 sg13g2_tiehi _714__29 (.L_HI(net29));
 sg13g2_tiehi _713__30 (.L_HI(net30));
 sg13g2_tiehi _712__31 (.L_HI(net31));
 sg13g2_tiehi _771__32 (.L_HI(net32));
 sg13g2_tiehi _776__33 (.L_HI(net33));
 sg13g2_tiehi _770__34 (.L_HI(net34));
 sg13g2_tiehi _773__35 (.L_HI(net35));
 sg13g2_tiehi _769__36 (.L_HI(net36));
 sg13g2_tiehi _775__37 (.L_HI(net37));
 sg13g2_tiehi _768__38 (.L_HI(net38));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_algofoogle_fomo_2 (.L_LO(net2));
 sg13g2_tielo tt_um_algofoogle_fomo_3 (.L_LO(net3));
 sg13g2_tielo tt_um_algofoogle_fomo_4 (.L_LO(net4));
 sg13g2_tielo tt_um_algofoogle_fomo_5 (.L_LO(net5));
 sg13g2_tielo tt_um_algofoogle_fomo_6 (.L_LO(net6));
 sg13g2_tielo tt_um_algofoogle_fomo_7 (.L_LO(net7));
 sg13g2_tielo tt_um_algofoogle_fomo_8 (.L_LO(net8));
 sg13g2_tielo tt_um_algofoogle_fomo_9 (.L_LO(net9));
 sg13g2_tielo tt_um_algofoogle_fomo_10 (.L_LO(net10));
 sg13g2_tielo tt_um_algofoogle_fomo_11 (.L_LO(net11));
 sg13g2_tielo tt_um_algofoogle_fomo_12 (.L_LO(net12));
 sg13g2_tielo tt_um_algofoogle_fomo_13 (.L_LO(net13));
 sg13g2_tielo tt_um_algofoogle_fomo_14 (.L_LO(net14));
 sg13g2_tielo tt_um_algofoogle_fomo_15 (.L_LO(net15));
 sg13g2_tielo tt_um_algofoogle_fomo_16 (.L_LO(net16));
 sg13g2_tiehi _772__17 (.L_HI(net17));
 sg13g2_buf_1 _815_ (.A(net52),
    .X(uo_out[3]));
 sg13g2_buf_1 _816_ (.A(uo_out[5]),
    .X(uo_out[4]));
 sg13g2_buf_1 _817_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout42 (.A(_207_),
    .X(net42));
 sg13g2_buf_8 fanout43 (.A(_315_),
    .X(net43));
 sg13g2_buf_8 fanout44 (.A(_121_),
    .X(net44));
 sg13g2_buf_8 fanout45 (.A(_219_),
    .X(net45));
 sg13g2_buf_1 fanout46 (.A(net47),
    .X(net46));
 sg13g2_buf_8 fanout47 (.A(_219_),
    .X(net47));
 sg13g2_buf_8 fanout48 (.A(net49),
    .X(net48));
 sg13g2_buf_8 fanout49 (.A(_093_),
    .X(net49));
 sg13g2_buf_8 fanout50 (.A(\counter[5] ),
    .X(net50));
 sg13g2_buf_8 fanout51 (.A(\counter[4] ),
    .X(net51));
 sg13g2_buf_8 fanout52 (.A(\hvsync_gen.vsync ),
    .X(net52));
 sg13g2_buf_8 fanout53 (.A(net55),
    .X(net53));
 sg13g2_buf_8 fanout54 (.A(net55),
    .X(net54));
 sg13g2_buf_8 fanout55 (.A(rst_n),
    .X(net55));
 sg13g2_buf_8 fanout56 (.A(net60),
    .X(net56));
 sg13g2_buf_8 fanout57 (.A(net60),
    .X(net57));
 sg13g2_buf_8 fanout58 (.A(net60),
    .X(net58));
 sg13g2_buf_8 fanout59 (.A(net60),
    .X(net59));
 sg13g2_buf_8 fanout60 (.A(rst_n),
    .X(net60));
 sg13g2_tielo tt_um_algofoogle_fomo_1 (.L_LO(net1));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_3_6__leaf_clk));
 sg13g2_buf_1 clkload6 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\vy[0] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold2 (.A(\h[0] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold3 (.A(_012_),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold4 (.A(\vx[0] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold5 (.A(\pix_y[2] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold6 (.A(\pix_y[4] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold7 (.A(_054_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold8 (.A(\pix_y[1] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold9 (.A(_051_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold10 (.A(\h[5] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold11 (.A(_017_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold12 (.A(\pix_y[0] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold13 (.A(\h[2] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold14 (.A(_124_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold15 (.A(_014_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold16 (.A(\vx[12] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold17 (.A(_034_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold18 (.A(\vx[17] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold19 (.A(_039_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold20 (.A(\h[9] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold21 (.A(_021_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold22 (.A(\h[1] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold23 (.A(\vx[7] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold24 (.A(_029_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold25 (.A(\hvsync_gen.vpos[8] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold26 (.A(_340_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold27 (.A(_064_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold28 (.A(\vx[16] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold29 (.A(_216_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold30 (.A(_038_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold31 (.A(\vx[13] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold32 (.A(\vx[3] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold33 (.A(_025_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold34 (.A(\vx[1] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold35 (.A(\vy[6] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold36 (.A(\vy[2] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold37 (.A(_042_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold38 (.A(\vy[7] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold39 (.A(_047_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold40 (.A(\vy[8] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold41 (.A(_048_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold42 (.A(\vy[5] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold43 (.A(_045_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold44 (.A(\vx[2] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold45 (.A(\vy[9] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold46 (.A(\vx[6] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold47 (.A(\hvsync_gen.vpos[7] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold48 (.A(_063_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold49 (.A(\vx[9] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold50 (.A(_031_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold51 (.A(\vy[1] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold52 (.A(_041_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold53 (.A(\vx[15] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold54 (.A(_213_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold55 (.A(_037_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold56 (.A(\pix_y[5] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold57 (.A(_055_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold58 (.A(\hvsync_gen.vpos[6] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold59 (.A(_062_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold60 (.A(\vx[11] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold61 (.A(_033_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold62 (.A(\hvsync_gen.vpos[0] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold63 (.A(\h[6] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold64 (.A(_128_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold65 (.A(_018_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold66 (.A(\hvsync_gen.vpos[4] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold67 (.A(_328_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold68 (.A(\h[8] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold69 (.A(_131_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold70 (.A(_020_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold71 (.A(\hvsync_gen.vpos[1] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold72 (.A(_001_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold73 (.A(\vx[10] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold74 (.A(_032_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold75 (.A(\vx[8] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold76 (.A(\vx[4] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold77 (.A(_026_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold78 (.A(\h[4] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold79 (.A(_000_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold80 (.A(\vy[4] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold81 (.A(\vx[14] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold82 (.A(\vy[3] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold83 (.A(\hvsync_gen.vpos[5] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold84 (.A(\vx[5] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold85 (.A(\hvsync_gen.vpos[3] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold86 (.A(_325_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold87 (.A(\hvsync_gen.vpos[2] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold88 (.A(\hvsync_gen.vpos[9] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold89 (.A(_065_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold90 (.A(\h[3] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold91 (.A(\h[7] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold92 (.A(\pix_y[3] ),
    .X(net149));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_fill_2 FILLER_17_322 ();
 sg13g2_fill_1 FILLER_17_324 ();
 sg13g2_decap_8 FILLER_17_333 ();
 sg13g2_decap_8 FILLER_17_340 ();
 sg13g2_decap_8 FILLER_17_347 ();
 sg13g2_decap_8 FILLER_17_354 ();
 sg13g2_decap_8 FILLER_17_361 ();
 sg13g2_decap_8 FILLER_17_368 ();
 sg13g2_decap_8 FILLER_17_375 ();
 sg13g2_decap_8 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_4 FILLER_17_403 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_fill_2 FILLER_18_294 ();
 sg13g2_fill_1 FILLER_18_296 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_317 ();
 sg13g2_fill_1 FILLER_18_324 ();
 sg13g2_decap_8 FILLER_18_334 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_4 FILLER_19_280 ();
 sg13g2_fill_1 FILLER_19_284 ();
 sg13g2_decap_4 FILLER_19_317 ();
 sg13g2_fill_2 FILLER_19_321 ();
 sg13g2_decap_8 FILLER_19_377 ();
 sg13g2_decap_8 FILLER_19_384 ();
 sg13g2_decap_8 FILLER_19_391 ();
 sg13g2_decap_8 FILLER_19_398 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_4 FILLER_20_203 ();
 sg13g2_fill_1 FILLER_20_207 ();
 sg13g2_fill_1 FILLER_20_221 ();
 sg13g2_decap_8 FILLER_20_254 ();
 sg13g2_decap_8 FILLER_20_261 ();
 sg13g2_fill_1 FILLER_20_268 ();
 sg13g2_fill_1 FILLER_20_273 ();
 sg13g2_fill_2 FILLER_20_282 ();
 sg13g2_fill_1 FILLER_20_284 ();
 sg13g2_decap_8 FILLER_20_299 ();
 sg13g2_decap_8 FILLER_20_306 ();
 sg13g2_decap_8 FILLER_20_313 ();
 sg13g2_decap_8 FILLER_20_320 ();
 sg13g2_decap_4 FILLER_20_327 ();
 sg13g2_fill_1 FILLER_20_331 ();
 sg13g2_fill_2 FILLER_20_337 ();
 sg13g2_decap_4 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_352 ();
 sg13g2_fill_1 FILLER_20_359 ();
 sg13g2_decap_4 FILLER_20_364 ();
 sg13g2_fill_2 FILLER_20_368 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_4 FILLER_21_168 ();
 sg13g2_fill_1 FILLER_21_172 ();
 sg13g2_fill_1 FILLER_21_194 ();
 sg13g2_fill_2 FILLER_21_230 ();
 sg13g2_decap_8 FILLER_21_235 ();
 sg13g2_decap_4 FILLER_21_242 ();
 sg13g2_decap_4 FILLER_21_271 ();
 sg13g2_fill_1 FILLER_21_275 ();
 sg13g2_fill_2 FILLER_21_300 ();
 sg13g2_fill_1 FILLER_21_302 ();
 sg13g2_decap_4 FILLER_21_323 ();
 sg13g2_fill_2 FILLER_21_327 ();
 sg13g2_decap_8 FILLER_21_352 ();
 sg13g2_decap_4 FILLER_21_359 ();
 sg13g2_fill_2 FILLER_21_384 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_fill_2 FILLER_22_154 ();
 sg13g2_decap_4 FILLER_22_183 ();
 sg13g2_fill_2 FILLER_22_187 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_4 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_4 FILLER_22_238 ();
 sg13g2_fill_2 FILLER_22_242 ();
 sg13g2_decap_4 FILLER_22_274 ();
 sg13g2_fill_1 FILLER_22_278 ();
 sg13g2_fill_2 FILLER_22_285 ();
 sg13g2_decap_8 FILLER_22_292 ();
 sg13g2_fill_1 FILLER_22_299 ();
 sg13g2_decap_8 FILLER_22_313 ();
 sg13g2_decap_8 FILLER_22_320 ();
 sg13g2_decap_4 FILLER_22_327 ();
 sg13g2_fill_2 FILLER_22_331 ();
 sg13g2_decap_8 FILLER_22_351 ();
 sg13g2_decap_4 FILLER_22_358 ();
 sg13g2_fill_1 FILLER_22_362 ();
 sg13g2_decap_4 FILLER_22_376 ();
 sg13g2_fill_1 FILLER_22_393 ();
 sg13g2_decap_8 FILLER_22_402 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_fill_2 FILLER_23_98 ();
 sg13g2_fill_1 FILLER_23_100 ();
 sg13g2_decap_8 FILLER_23_109 ();
 sg13g2_decap_8 FILLER_23_116 ();
 sg13g2_decap_8 FILLER_23_123 ();
 sg13g2_decap_8 FILLER_23_130 ();
 sg13g2_decap_8 FILLER_23_137 ();
 sg13g2_decap_8 FILLER_23_144 ();
 sg13g2_decap_8 FILLER_23_151 ();
 sg13g2_decap_8 FILLER_23_158 ();
 sg13g2_decap_4 FILLER_23_165 ();
 sg13g2_fill_1 FILLER_23_169 ();
 sg13g2_fill_2 FILLER_23_179 ();
 sg13g2_decap_8 FILLER_23_198 ();
 sg13g2_decap_8 FILLER_23_205 ();
 sg13g2_fill_2 FILLER_23_225 ();
 sg13g2_fill_2 FILLER_23_254 ();
 sg13g2_decap_8 FILLER_23_270 ();
 sg13g2_decap_4 FILLER_23_277 ();
 sg13g2_fill_1 FILLER_23_281 ();
 sg13g2_fill_2 FILLER_23_302 ();
 sg13g2_decap_8 FILLER_23_323 ();
 sg13g2_decap_4 FILLER_23_330 ();
 sg13g2_fill_1 FILLER_23_334 ();
 sg13g2_decap_8 FILLER_23_349 ();
 sg13g2_fill_1 FILLER_23_356 ();
 sg13g2_fill_2 FILLER_23_378 ();
 sg13g2_fill_1 FILLER_23_380 ();
 sg13g2_fill_1 FILLER_23_390 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_4 FILLER_24_35 ();
 sg13g2_fill_1 FILLER_24_39 ();
 sg13g2_decap_8 FILLER_24_44 ();
 sg13g2_decap_8 FILLER_24_51 ();
 sg13g2_decap_8 FILLER_24_58 ();
 sg13g2_fill_1 FILLER_24_65 ();
 sg13g2_fill_2 FILLER_24_93 ();
 sg13g2_fill_1 FILLER_24_95 ();
 sg13g2_fill_2 FILLER_24_124 ();
 sg13g2_decap_8 FILLER_24_130 ();
 sg13g2_fill_2 FILLER_24_141 ();
 sg13g2_fill_1 FILLER_24_143 ();
 sg13g2_fill_2 FILLER_24_188 ();
 sg13g2_decap_8 FILLER_24_198 ();
 sg13g2_decap_4 FILLER_24_205 ();
 sg13g2_fill_2 FILLER_24_209 ();
 sg13g2_decap_8 FILLER_24_237 ();
 sg13g2_decap_8 FILLER_24_244 ();
 sg13g2_decap_8 FILLER_24_276 ();
 sg13g2_decap_8 FILLER_24_283 ();
 sg13g2_fill_1 FILLER_24_290 ();
 sg13g2_decap_8 FILLER_24_296 ();
 sg13g2_decap_4 FILLER_24_303 ();
 sg13g2_fill_2 FILLER_24_307 ();
 sg13g2_decap_4 FILLER_24_347 ();
 sg13g2_fill_1 FILLER_24_351 ();
 sg13g2_fill_1 FILLER_24_365 ();
 sg13g2_fill_1 FILLER_24_371 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_4 FILLER_25_28 ();
 sg13g2_fill_2 FILLER_25_69 ();
 sg13g2_decap_4 FILLER_25_78 ();
 sg13g2_fill_1 FILLER_25_82 ();
 sg13g2_fill_2 FILLER_25_98 ();
 sg13g2_decap_4 FILLER_25_123 ();
 sg13g2_decap_8 FILLER_25_160 ();
 sg13g2_decap_8 FILLER_25_167 ();
 sg13g2_decap_8 FILLER_25_174 ();
 sg13g2_decap_4 FILLER_25_212 ();
 sg13g2_fill_2 FILLER_25_292 ();
 sg13g2_fill_1 FILLER_25_294 ();
 sg13g2_fill_2 FILLER_25_307 ();
 sg13g2_decap_4 FILLER_25_326 ();
 sg13g2_decap_8 FILLER_25_365 ();
 sg13g2_decap_8 FILLER_25_372 ();
 sg13g2_decap_8 FILLER_25_379 ();
 sg13g2_decap_8 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_4 FILLER_26_28 ();
 sg13g2_fill_2 FILLER_26_32 ();
 sg13g2_decap_8 FILLER_26_38 ();
 sg13g2_fill_1 FILLER_26_73 ();
 sg13g2_fill_1 FILLER_26_105 ();
 sg13g2_fill_2 FILLER_26_116 ();
 sg13g2_fill_1 FILLER_26_118 ();
 sg13g2_fill_2 FILLER_26_129 ();
 sg13g2_fill_1 FILLER_26_131 ();
 sg13g2_fill_1 FILLER_26_141 ();
 sg13g2_decap_8 FILLER_26_146 ();
 sg13g2_decap_8 FILLER_26_174 ();
 sg13g2_decap_8 FILLER_26_181 ();
 sg13g2_decap_8 FILLER_26_188 ();
 sg13g2_decap_4 FILLER_26_195 ();
 sg13g2_fill_2 FILLER_26_199 ();
 sg13g2_decap_8 FILLER_26_213 ();
 sg13g2_decap_8 FILLER_26_220 ();
 sg13g2_decap_4 FILLER_26_227 ();
 sg13g2_decap_8 FILLER_26_240 ();
 sg13g2_decap_8 FILLER_26_247 ();
 sg13g2_decap_4 FILLER_26_254 ();
 sg13g2_decap_8 FILLER_26_263 ();
 sg13g2_decap_4 FILLER_26_270 ();
 sg13g2_fill_2 FILLER_26_274 ();
 sg13g2_fill_1 FILLER_26_293 ();
 sg13g2_decap_8 FILLER_26_355 ();
 sg13g2_fill_2 FILLER_26_362 ();
 sg13g2_fill_1 FILLER_26_364 ();
 sg13g2_fill_1 FILLER_26_377 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_4 FILLER_27_21 ();
 sg13g2_fill_1 FILLER_27_25 ();
 sg13g2_fill_2 FILLER_27_57 ();
 sg13g2_decap_4 FILLER_27_94 ();
 sg13g2_decap_8 FILLER_27_125 ();
 sg13g2_decap_4 FILLER_27_231 ();
 sg13g2_fill_1 FILLER_27_235 ();
 sg13g2_decap_8 FILLER_27_249 ();
 sg13g2_decap_4 FILLER_27_256 ();
 sg13g2_decap_8 FILLER_27_272 ();
 sg13g2_decap_8 FILLER_27_285 ();
 sg13g2_decap_4 FILLER_27_292 ();
 sg13g2_fill_2 FILLER_27_296 ();
 sg13g2_decap_8 FILLER_27_311 ();
 sg13g2_decap_8 FILLER_27_318 ();
 sg13g2_decap_4 FILLER_27_325 ();
 sg13g2_fill_2 FILLER_27_329 ();
 sg13g2_fill_1 FILLER_27_366 ();
 sg13g2_fill_2 FILLER_27_375 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_fill_2 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_37 ();
 sg13g2_decap_4 FILLER_28_44 ();
 sg13g2_fill_2 FILLER_28_48 ();
 sg13g2_fill_2 FILLER_28_87 ();
 sg13g2_fill_1 FILLER_28_89 ();
 sg13g2_decap_4 FILLER_28_111 ();
 sg13g2_fill_2 FILLER_28_115 ();
 sg13g2_decap_8 FILLER_28_159 ();
 sg13g2_decap_8 FILLER_28_192 ();
 sg13g2_fill_2 FILLER_28_199 ();
 sg13g2_fill_1 FILLER_28_201 ();
 sg13g2_decap_8 FILLER_28_207 ();
 sg13g2_decap_4 FILLER_28_214 ();
 sg13g2_fill_1 FILLER_28_231 ();
 sg13g2_fill_2 FILLER_28_335 ();
 sg13g2_decap_4 FILLER_28_341 ();
 sg13g2_fill_1 FILLER_28_345 ();
 sg13g2_decap_8 FILLER_28_355 ();
 sg13g2_decap_4 FILLER_28_362 ();
 sg13g2_fill_2 FILLER_28_366 ();
 sg13g2_decap_8 FILLER_28_377 ();
 sg13g2_decap_8 FILLER_28_384 ();
 sg13g2_decap_8 FILLER_28_391 ();
 sg13g2_decap_8 FILLER_28_398 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_fill_1 FILLER_29_75 ();
 sg13g2_decap_8 FILLER_29_104 ();
 sg13g2_fill_1 FILLER_29_111 ();
 sg13g2_fill_1 FILLER_29_131 ();
 sg13g2_fill_1 FILLER_29_169 ();
 sg13g2_fill_1 FILLER_29_211 ();
 sg13g2_decap_8 FILLER_29_242 ();
 sg13g2_decap_8 FILLER_29_249 ();
 sg13g2_decap_4 FILLER_29_256 ();
 sg13g2_fill_2 FILLER_29_260 ();
 sg13g2_decap_4 FILLER_29_280 ();
 sg13g2_fill_1 FILLER_29_284 ();
 sg13g2_decap_4 FILLER_29_289 ();
 sg13g2_fill_1 FILLER_29_293 ();
 sg13g2_fill_1 FILLER_29_302 ();
 sg13g2_decap_4 FILLER_29_317 ();
 sg13g2_fill_1 FILLER_29_321 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_4 FILLER_30_28 ();
 sg13g2_fill_1 FILLER_30_32 ();
 sg13g2_fill_2 FILLER_30_66 ();
 sg13g2_decap_4 FILLER_30_85 ();
 sg13g2_fill_1 FILLER_30_89 ();
 sg13g2_fill_2 FILLER_30_110 ();
 sg13g2_fill_2 FILLER_30_121 ();
 sg13g2_fill_1 FILLER_30_123 ();
 sg13g2_decap_8 FILLER_30_162 ();
 sg13g2_decap_8 FILLER_30_169 ();
 sg13g2_decap_8 FILLER_30_176 ();
 sg13g2_fill_1 FILLER_30_183 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_4 FILLER_30_203 ();
 sg13g2_fill_2 FILLER_30_207 ();
 sg13g2_decap_8 FILLER_30_219 ();
 sg13g2_decap_4 FILLER_30_226 ();
 sg13g2_decap_8 FILLER_30_244 ();
 sg13g2_fill_2 FILLER_30_293 ();
 sg13g2_fill_1 FILLER_30_295 ();
 sg13g2_fill_2 FILLER_30_306 ();
 sg13g2_fill_1 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_317 ();
 sg13g2_decap_8 FILLER_30_324 ();
 sg13g2_decap_8 FILLER_30_331 ();
 sg13g2_decap_4 FILLER_30_338 ();
 sg13g2_fill_1 FILLER_30_342 ();
 sg13g2_fill_2 FILLER_30_347 ();
 sg13g2_decap_4 FILLER_30_354 ();
 sg13g2_fill_1 FILLER_30_362 ();
 sg13g2_fill_1 FILLER_30_375 ();
 sg13g2_decap_8 FILLER_30_381 ();
 sg13g2_fill_2 FILLER_30_388 ();
 sg13g2_fill_1 FILLER_30_390 ();
 sg13g2_decap_8 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_fill_2 FILLER_31_35 ();
 sg13g2_fill_1 FILLER_31_37 ();
 sg13g2_decap_4 FILLER_31_42 ();
 sg13g2_fill_2 FILLER_31_55 ();
 sg13g2_fill_1 FILLER_31_57 ();
 sg13g2_fill_2 FILLER_31_67 ();
 sg13g2_fill_1 FILLER_31_69 ();
 sg13g2_decap_4 FILLER_31_77 ();
 sg13g2_fill_1 FILLER_31_103 ();
 sg13g2_fill_2 FILLER_31_132 ();
 sg13g2_fill_2 FILLER_31_139 ();
 sg13g2_fill_1 FILLER_31_141 ();
 sg13g2_decap_8 FILLER_31_202 ();
 sg13g2_fill_2 FILLER_31_209 ();
 sg13g2_fill_1 FILLER_31_211 ();
 sg13g2_fill_2 FILLER_31_223 ();
 sg13g2_fill_2 FILLER_31_237 ();
 sg13g2_decap_8 FILLER_31_256 ();
 sg13g2_decap_4 FILLER_31_263 ();
 sg13g2_decap_8 FILLER_31_275 ();
 sg13g2_decap_8 FILLER_31_282 ();
 sg13g2_decap_4 FILLER_31_289 ();
 sg13g2_fill_2 FILLER_31_293 ();
 sg13g2_fill_2 FILLER_31_311 ();
 sg13g2_fill_2 FILLER_31_318 ();
 sg13g2_fill_1 FILLER_31_320 ();
 sg13g2_fill_2 FILLER_31_337 ();
 sg13g2_fill_1 FILLER_31_358 ();
 sg13g2_decap_4 FILLER_31_367 ();
 sg13g2_fill_1 FILLER_31_371 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_4 FILLER_32_28 ();
 sg13g2_fill_1 FILLER_32_64 ();
 sg13g2_fill_2 FILLER_32_93 ();
 sg13g2_fill_2 FILLER_32_120 ();
 sg13g2_fill_2 FILLER_32_150 ();
 sg13g2_fill_1 FILLER_32_152 ();
 sg13g2_fill_2 FILLER_32_166 ();
 sg13g2_fill_2 FILLER_32_193 ();
 sg13g2_fill_1 FILLER_32_195 ();
 sg13g2_decap_8 FILLER_32_209 ();
 sg13g2_decap_8 FILLER_32_216 ();
 sg13g2_fill_1 FILLER_32_223 ();
 sg13g2_fill_1 FILLER_32_244 ();
 sg13g2_decap_4 FILLER_32_280 ();
 sg13g2_fill_2 FILLER_32_284 ();
 sg13g2_fill_1 FILLER_32_295 ();
 sg13g2_decap_8 FILLER_32_333 ();
 sg13g2_decap_8 FILLER_32_340 ();
 sg13g2_decap_8 FILLER_32_351 ();
 sg13g2_decap_8 FILLER_32_358 ();
 sg13g2_fill_1 FILLER_32_365 ();
 sg13g2_decap_4 FILLER_32_384 ();
 sg13g2_fill_1 FILLER_32_388 ();
 sg13g2_decap_8 FILLER_32_398 ();
 sg13g2_decap_4 FILLER_32_405 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_fill_2 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_41 ();
 sg13g2_decap_8 FILLER_33_48 ();
 sg13g2_decap_4 FILLER_33_55 ();
 sg13g2_fill_1 FILLER_33_59 ();
 sg13g2_decap_8 FILLER_33_69 ();
 sg13g2_fill_1 FILLER_33_95 ();
 sg13g2_fill_2 FILLER_33_133 ();
 sg13g2_fill_1 FILLER_33_135 ();
 sg13g2_fill_2 FILLER_33_149 ();
 sg13g2_fill_1 FILLER_33_151 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_fill_2 FILLER_33_175 ();
 sg13g2_fill_1 FILLER_33_177 ();
 sg13g2_fill_2 FILLER_33_221 ();
 sg13g2_fill_1 FILLER_33_223 ();
 sg13g2_fill_1 FILLER_33_320 ();
 sg13g2_decap_8 FILLER_33_358 ();
 sg13g2_fill_2 FILLER_33_365 ();
 sg13g2_fill_1 FILLER_33_367 ();
 sg13g2_decap_8 FILLER_33_376 ();
 sg13g2_decap_4 FILLER_33_383 ();
 sg13g2_fill_2 FILLER_33_387 ();
 sg13g2_decap_8 FILLER_33_398 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_fill_2 FILLER_34_60 ();
 sg13g2_fill_1 FILLER_34_62 ();
 sg13g2_decap_4 FILLER_34_76 ();
 sg13g2_fill_2 FILLER_34_80 ();
 sg13g2_fill_2 FILLER_34_128 ();
 sg13g2_decap_4 FILLER_34_195 ();
 sg13g2_fill_2 FILLER_34_199 ();
 sg13g2_fill_1 FILLER_34_256 ();
 sg13g2_fill_2 FILLER_34_272 ();
 sg13g2_fill_1 FILLER_34_274 ();
 sg13g2_fill_2 FILLER_34_292 ();
 sg13g2_decap_8 FILLER_34_321 ();
 sg13g2_decap_4 FILLER_34_328 ();
 sg13g2_decap_4 FILLER_34_350 ();
 sg13g2_fill_2 FILLER_34_354 ();
 sg13g2_fill_2 FILLER_34_374 ();
 sg13g2_decap_4 FILLER_34_403 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_4 FILLER_35_28 ();
 sg13g2_fill_2 FILLER_35_32 ();
 sg13g2_fill_1 FILLER_35_75 ();
 sg13g2_decap_4 FILLER_35_81 ();
 sg13g2_fill_2 FILLER_35_85 ();
 sg13g2_decap_4 FILLER_35_91 ();
 sg13g2_fill_2 FILLER_35_118 ();
 sg13g2_fill_1 FILLER_35_120 ();
 sg13g2_fill_2 FILLER_35_139 ();
 sg13g2_fill_2 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_206 ();
 sg13g2_fill_2 FILLER_35_213 ();
 sg13g2_fill_1 FILLER_35_215 ();
 sg13g2_fill_2 FILLER_35_225 ();
 sg13g2_fill_1 FILLER_35_227 ();
 sg13g2_fill_2 FILLER_35_289 ();
 sg13g2_fill_1 FILLER_35_291 ();
 sg13g2_fill_1 FILLER_35_300 ();
 sg13g2_fill_2 FILLER_35_352 ();
 sg13g2_fill_1 FILLER_35_354 ();
 sg13g2_fill_2 FILLER_35_373 ();
 sg13g2_decap_8 FILLER_35_388 ();
 sg13g2_decap_8 FILLER_35_395 ();
 sg13g2_decap_8 FILLER_35_402 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_4 FILLER_36_35 ();
 sg13g2_decap_4 FILLER_36_43 ();
 sg13g2_fill_2 FILLER_36_47 ();
 sg13g2_fill_1 FILLER_36_58 ();
 sg13g2_fill_2 FILLER_36_174 ();
 sg13g2_fill_2 FILLER_36_198 ();
 sg13g2_fill_1 FILLER_36_200 ();
 sg13g2_fill_1 FILLER_36_233 ();
 sg13g2_fill_1 FILLER_36_261 ();
 sg13g2_fill_2 FILLER_36_271 ();
 sg13g2_fill_1 FILLER_36_273 ();
 sg13g2_decap_4 FILLER_36_301 ();
 sg13g2_fill_2 FILLER_36_305 ();
 sg13g2_fill_2 FILLER_36_353 ();
 sg13g2_fill_1 FILLER_36_355 ();
 sg13g2_decap_8 FILLER_36_392 ();
 sg13g2_decap_8 FILLER_36_399 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_fill_2 FILLER_37_56 ();
 sg13g2_fill_1 FILLER_37_58 ();
 sg13g2_fill_2 FILLER_37_95 ();
 sg13g2_fill_1 FILLER_37_97 ();
 sg13g2_fill_2 FILLER_37_102 ();
 sg13g2_fill_1 FILLER_37_108 ();
 sg13g2_fill_2 FILLER_37_116 ();
 sg13g2_decap_8 FILLER_37_131 ();
 sg13g2_decap_8 FILLER_37_138 ();
 sg13g2_decap_8 FILLER_37_145 ();
 sg13g2_decap_8 FILLER_37_152 ();
 sg13g2_decap_8 FILLER_37_159 ();
 sg13g2_fill_2 FILLER_37_166 ();
 sg13g2_fill_2 FILLER_37_172 ();
 sg13g2_decap_4 FILLER_37_183 ();
 sg13g2_fill_2 FILLER_37_190 ();
 sg13g2_decap_8 FILLER_37_209 ();
 sg13g2_decap_8 FILLER_37_216 ();
 sg13g2_fill_1 FILLER_37_235 ();
 sg13g2_fill_2 FILLER_37_286 ();
 sg13g2_fill_1 FILLER_37_342 ();
 sg13g2_fill_2 FILLER_37_352 ();
 sg13g2_fill_1 FILLER_37_354 ();
 sg13g2_decap_8 FILLER_37_368 ();
 sg13g2_decap_8 FILLER_37_375 ();
 sg13g2_decap_8 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_37_396 ();
 sg13g2_decap_4 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_4 FILLER_38_49 ();
 sg13g2_fill_1 FILLER_38_53 ();
 sg13g2_fill_1 FILLER_38_71 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_fill_1 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_fill_2 FILLER_38_156 ();
 sg13g2_fill_2 FILLER_38_198 ();
 sg13g2_fill_2 FILLER_38_236 ();
 sg13g2_fill_1 FILLER_38_243 ();
 sg13g2_fill_1 FILLER_38_249 ();
 sg13g2_fill_1 FILLER_38_268 ();
 sg13g2_decap_8 FILLER_38_277 ();
 sg13g2_fill_2 FILLER_38_284 ();
 sg13g2_fill_1 FILLER_38_286 ();
 sg13g2_decap_8 FILLER_38_296 ();
 sg13g2_decap_8 FILLER_38_303 ();
 sg13g2_decap_8 FILLER_38_310 ();
 sg13g2_decap_8 FILLER_38_317 ();
 sg13g2_decap_8 FILLER_38_324 ();
 sg13g2_decap_4 FILLER_38_331 ();
 sg13g2_fill_2 FILLER_38_335 ();
 sg13g2_decap_8 FILLER_38_365 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_379 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net1;
 assign uio_oe[1] = net2;
 assign uio_oe[2] = net3;
 assign uio_oe[3] = net4;
 assign uio_oe[4] = net5;
 assign uio_oe[5] = net6;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net8;
 assign uio_out[0] = net9;
 assign uio_out[1] = net10;
 assign uio_out[2] = net11;
 assign uio_out[3] = net12;
 assign uio_out[4] = net13;
 assign uio_out[5] = net14;
 assign uio_out[6] = net15;
 assign uio_out[7] = net16;
endmodule
