module tt_um_vga_tetris (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire clknet_leaf_0_clk;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire vga_hs;
 wire \vga_tetris._inputs_io_downButtonActive ;
 wire \vga_tetris._inputs_io_leftButtonActive ;
 wire \vga_tetris._inputs_io_rightButtonActive ;
 wire \vga_tetris._inputs_io_rotateButtonActive ;
 wire \vga_tetris._tetrisDisplay_io_boardYCoord[0] ;
 wire \vga_tetris._tetrisDisplay_io_boardYCoord[1] ;
 wire \vga_tetris._tetrisLogic_io_gameOver ;
 wire \vga_tetris._tetrisLogic_io_score_0[0] ;
 wire \vga_tetris._tetrisLogic_io_score_0[1] ;
 wire \vga_tetris._tetrisLogic_io_score_0[2] ;
 wire \vga_tetris._tetrisLogic_io_score_0[3] ;
 wire \vga_tetris._tetrisLogic_io_score_1[0] ;
 wire \vga_tetris._tetrisLogic_io_score_1[1] ;
 wire \vga_tetris._tetrisLogic_io_score_1[2] ;
 wire \vga_tetris._tetrisLogic_io_score_1[3] ;
 wire \vga_tetris._tetrisLogic_io_score_2[0] ;
 wire \vga_tetris._tetrisLogic_io_score_2[1] ;
 wire \vga_tetris._tetrisLogic_io_score_2[2] ;
 wire \vga_tetris._tetrisLogic_io_score_2[3] ;
 wire \vga_tetris._tetrisLogic_io_score_3[0] ;
 wire \vga_tetris._tetrisLogic_io_score_3[1] ;
 wire \vga_tetris._tetrisLogic_io_score_3[2] ;
 wire \vga_tetris._tetrisLogic_io_score_3[3] ;
 wire \vga_tetris._vgaController_io_pixelPosX[0] ;
 wire \vga_tetris._vgaController_io_pixelPosX[1] ;
 wire \vga_tetris._vgaController_io_pixelPosX[2] ;
 wire \vga_tetris._vgaController_io_pixelPosX[3] ;
 wire \vga_tetris._vgaController_io_pixelPosX[4] ;
 wire \vga_tetris._vgaController_io_pixelPosX[5] ;
 wire \vga_tetris._vgaController_io_pixelPosX[6] ;
 wire \vga_tetris._vgaController_io_pixelPosX[7] ;
 wire \vga_tetris._vgaController_io_pixelPosX[8] ;
 wire \vga_tetris._vgaController_io_pixelPosX[9] ;
 wire \vga_tetris._vgaController_io_pixelPosY[0] ;
 wire \vga_tetris._vgaController_io_pixelPosY[1] ;
 wire \vga_tetris._vgaController_io_pixelPosY[2] ;
 wire \vga_tetris._vgaController_io_pixelPosY[3] ;
 wire \vga_tetris._vgaController_io_pixelPosY[6] ;
 wire \vga_tetris._vgaController_io_pixelPosY[7] ;
 wire \vga_tetris._vgaController_io_pixelPosY[8] ;
 wire \vga_tetris._vgaController_io_pixelPosY[9] ;
 wire \vga_tetris._vgaController_io_vSync ;
 wire \vga_tetris.boardMem.board_0[0] ;
 wire \vga_tetris.boardMem.board_0[10] ;
 wire \vga_tetris.boardMem.board_0[11] ;
 wire \vga_tetris.boardMem.board_0[12] ;
 wire \vga_tetris.boardMem.board_0[13] ;
 wire \vga_tetris.boardMem.board_0[14] ;
 wire \vga_tetris.boardMem.board_0[15] ;
 wire \vga_tetris.boardMem.board_0[16] ;
 wire \vga_tetris.boardMem.board_0[17] ;
 wire \vga_tetris.boardMem.board_0[18] ;
 wire \vga_tetris.boardMem.board_0[19] ;
 wire \vga_tetris.boardMem.board_0[1] ;
 wire \vga_tetris.boardMem.board_0[2] ;
 wire \vga_tetris.boardMem.board_0[3] ;
 wire \vga_tetris.boardMem.board_0[4] ;
 wire \vga_tetris.boardMem.board_0[5] ;
 wire \vga_tetris.boardMem.board_0[6] ;
 wire \vga_tetris.boardMem.board_0[7] ;
 wire \vga_tetris.boardMem.board_0[8] ;
 wire \vga_tetris.boardMem.board_0[9] ;
 wire \vga_tetris.boardMem.board_10[0] ;
 wire \vga_tetris.boardMem.board_10[10] ;
 wire \vga_tetris.boardMem.board_10[11] ;
 wire \vga_tetris.boardMem.board_10[12] ;
 wire \vga_tetris.boardMem.board_10[13] ;
 wire \vga_tetris.boardMem.board_10[14] ;
 wire \vga_tetris.boardMem.board_10[15] ;
 wire \vga_tetris.boardMem.board_10[16] ;
 wire \vga_tetris.boardMem.board_10[17] ;
 wire \vga_tetris.boardMem.board_10[18] ;
 wire \vga_tetris.boardMem.board_10[19] ;
 wire \vga_tetris.boardMem.board_10[1] ;
 wire \vga_tetris.boardMem.board_10[2] ;
 wire \vga_tetris.boardMem.board_10[3] ;
 wire \vga_tetris.boardMem.board_10[4] ;
 wire \vga_tetris.boardMem.board_10[5] ;
 wire \vga_tetris.boardMem.board_10[6] ;
 wire \vga_tetris.boardMem.board_10[7] ;
 wire \vga_tetris.boardMem.board_10[8] ;
 wire \vga_tetris.boardMem.board_10[9] ;
 wire \vga_tetris.boardMem.board_11[0] ;
 wire \vga_tetris.boardMem.board_11[10] ;
 wire \vga_tetris.boardMem.board_11[11] ;
 wire \vga_tetris.boardMem.board_11[12] ;
 wire \vga_tetris.boardMem.board_11[13] ;
 wire \vga_tetris.boardMem.board_11[14] ;
 wire \vga_tetris.boardMem.board_11[15] ;
 wire \vga_tetris.boardMem.board_11[16] ;
 wire \vga_tetris.boardMem.board_11[17] ;
 wire \vga_tetris.boardMem.board_11[18] ;
 wire \vga_tetris.boardMem.board_11[19] ;
 wire \vga_tetris.boardMem.board_11[1] ;
 wire \vga_tetris.boardMem.board_11[2] ;
 wire \vga_tetris.boardMem.board_11[3] ;
 wire \vga_tetris.boardMem.board_11[4] ;
 wire \vga_tetris.boardMem.board_11[5] ;
 wire \vga_tetris.boardMem.board_11[6] ;
 wire \vga_tetris.boardMem.board_11[7] ;
 wire \vga_tetris.boardMem.board_11[8] ;
 wire \vga_tetris.boardMem.board_11[9] ;
 wire \vga_tetris.boardMem.board_12[0] ;
 wire \vga_tetris.boardMem.board_12[10] ;
 wire \vga_tetris.boardMem.board_12[11] ;
 wire \vga_tetris.boardMem.board_12[12] ;
 wire \vga_tetris.boardMem.board_12[13] ;
 wire \vga_tetris.boardMem.board_12[14] ;
 wire \vga_tetris.boardMem.board_12[15] ;
 wire \vga_tetris.boardMem.board_12[16] ;
 wire \vga_tetris.boardMem.board_12[17] ;
 wire \vga_tetris.boardMem.board_12[18] ;
 wire \vga_tetris.boardMem.board_12[19] ;
 wire \vga_tetris.boardMem.board_12[1] ;
 wire \vga_tetris.boardMem.board_12[2] ;
 wire \vga_tetris.boardMem.board_12[3] ;
 wire \vga_tetris.boardMem.board_12[4] ;
 wire \vga_tetris.boardMem.board_12[5] ;
 wire \vga_tetris.boardMem.board_12[6] ;
 wire \vga_tetris.boardMem.board_12[7] ;
 wire \vga_tetris.boardMem.board_12[8] ;
 wire \vga_tetris.boardMem.board_12[9] ;
 wire \vga_tetris.boardMem.board_13[0] ;
 wire \vga_tetris.boardMem.board_13[10] ;
 wire \vga_tetris.boardMem.board_13[11] ;
 wire \vga_tetris.boardMem.board_13[12] ;
 wire \vga_tetris.boardMem.board_13[13] ;
 wire \vga_tetris.boardMem.board_13[14] ;
 wire \vga_tetris.boardMem.board_13[15] ;
 wire \vga_tetris.boardMem.board_13[16] ;
 wire \vga_tetris.boardMem.board_13[17] ;
 wire \vga_tetris.boardMem.board_13[18] ;
 wire \vga_tetris.boardMem.board_13[19] ;
 wire \vga_tetris.boardMem.board_13[1] ;
 wire \vga_tetris.boardMem.board_13[2] ;
 wire \vga_tetris.boardMem.board_13[3] ;
 wire \vga_tetris.boardMem.board_13[4] ;
 wire \vga_tetris.boardMem.board_13[5] ;
 wire \vga_tetris.boardMem.board_13[6] ;
 wire \vga_tetris.boardMem.board_13[7] ;
 wire \vga_tetris.boardMem.board_13[8] ;
 wire \vga_tetris.boardMem.board_13[9] ;
 wire \vga_tetris.boardMem.board_14[0] ;
 wire \vga_tetris.boardMem.board_14[10] ;
 wire \vga_tetris.boardMem.board_14[11] ;
 wire \vga_tetris.boardMem.board_14[12] ;
 wire \vga_tetris.boardMem.board_14[13] ;
 wire \vga_tetris.boardMem.board_14[14] ;
 wire \vga_tetris.boardMem.board_14[15] ;
 wire \vga_tetris.boardMem.board_14[16] ;
 wire \vga_tetris.boardMem.board_14[17] ;
 wire \vga_tetris.boardMem.board_14[18] ;
 wire \vga_tetris.boardMem.board_14[19] ;
 wire \vga_tetris.boardMem.board_14[1] ;
 wire \vga_tetris.boardMem.board_14[2] ;
 wire \vga_tetris.boardMem.board_14[3] ;
 wire \vga_tetris.boardMem.board_14[4] ;
 wire \vga_tetris.boardMem.board_14[5] ;
 wire \vga_tetris.boardMem.board_14[6] ;
 wire \vga_tetris.boardMem.board_14[7] ;
 wire \vga_tetris.boardMem.board_14[8] ;
 wire \vga_tetris.boardMem.board_14[9] ;
 wire \vga_tetris.boardMem.board_15[0] ;
 wire \vga_tetris.boardMem.board_15[10] ;
 wire \vga_tetris.boardMem.board_15[11] ;
 wire \vga_tetris.boardMem.board_15[12] ;
 wire \vga_tetris.boardMem.board_15[13] ;
 wire \vga_tetris.boardMem.board_15[14] ;
 wire \vga_tetris.boardMem.board_15[15] ;
 wire \vga_tetris.boardMem.board_15[16] ;
 wire \vga_tetris.boardMem.board_15[17] ;
 wire \vga_tetris.boardMem.board_15[18] ;
 wire \vga_tetris.boardMem.board_15[19] ;
 wire \vga_tetris.boardMem.board_15[1] ;
 wire \vga_tetris.boardMem.board_15[2] ;
 wire \vga_tetris.boardMem.board_15[3] ;
 wire \vga_tetris.boardMem.board_15[4] ;
 wire \vga_tetris.boardMem.board_15[5] ;
 wire \vga_tetris.boardMem.board_15[6] ;
 wire \vga_tetris.boardMem.board_15[7] ;
 wire \vga_tetris.boardMem.board_15[8] ;
 wire \vga_tetris.boardMem.board_15[9] ;
 wire \vga_tetris.boardMem.board_16[0] ;
 wire \vga_tetris.boardMem.board_16[10] ;
 wire \vga_tetris.boardMem.board_16[11] ;
 wire \vga_tetris.boardMem.board_16[12] ;
 wire \vga_tetris.boardMem.board_16[13] ;
 wire \vga_tetris.boardMem.board_16[14] ;
 wire \vga_tetris.boardMem.board_16[15] ;
 wire \vga_tetris.boardMem.board_16[16] ;
 wire \vga_tetris.boardMem.board_16[17] ;
 wire \vga_tetris.boardMem.board_16[18] ;
 wire \vga_tetris.boardMem.board_16[19] ;
 wire \vga_tetris.boardMem.board_16[1] ;
 wire \vga_tetris.boardMem.board_16[2] ;
 wire \vga_tetris.boardMem.board_16[3] ;
 wire \vga_tetris.boardMem.board_16[4] ;
 wire \vga_tetris.boardMem.board_16[5] ;
 wire \vga_tetris.boardMem.board_16[6] ;
 wire \vga_tetris.boardMem.board_16[7] ;
 wire \vga_tetris.boardMem.board_16[8] ;
 wire \vga_tetris.boardMem.board_16[9] ;
 wire \vga_tetris.boardMem.board_17[0] ;
 wire \vga_tetris.boardMem.board_17[10] ;
 wire \vga_tetris.boardMem.board_17[11] ;
 wire \vga_tetris.boardMem.board_17[12] ;
 wire \vga_tetris.boardMem.board_17[13] ;
 wire \vga_tetris.boardMem.board_17[14] ;
 wire \vga_tetris.boardMem.board_17[15] ;
 wire \vga_tetris.boardMem.board_17[16] ;
 wire \vga_tetris.boardMem.board_17[17] ;
 wire \vga_tetris.boardMem.board_17[18] ;
 wire \vga_tetris.boardMem.board_17[19] ;
 wire \vga_tetris.boardMem.board_17[1] ;
 wire \vga_tetris.boardMem.board_17[2] ;
 wire \vga_tetris.boardMem.board_17[3] ;
 wire \vga_tetris.boardMem.board_17[4] ;
 wire \vga_tetris.boardMem.board_17[5] ;
 wire \vga_tetris.boardMem.board_17[6] ;
 wire \vga_tetris.boardMem.board_17[7] ;
 wire \vga_tetris.boardMem.board_17[8] ;
 wire \vga_tetris.boardMem.board_17[9] ;
 wire \vga_tetris.boardMem.board_18[0] ;
 wire \vga_tetris.boardMem.board_18[10] ;
 wire \vga_tetris.boardMem.board_18[11] ;
 wire \vga_tetris.boardMem.board_18[12] ;
 wire \vga_tetris.boardMem.board_18[13] ;
 wire \vga_tetris.boardMem.board_18[14] ;
 wire \vga_tetris.boardMem.board_18[15] ;
 wire \vga_tetris.boardMem.board_18[16] ;
 wire \vga_tetris.boardMem.board_18[17] ;
 wire \vga_tetris.boardMem.board_18[18] ;
 wire \vga_tetris.boardMem.board_18[19] ;
 wire \vga_tetris.boardMem.board_18[1] ;
 wire \vga_tetris.boardMem.board_18[2] ;
 wire \vga_tetris.boardMem.board_18[3] ;
 wire \vga_tetris.boardMem.board_18[4] ;
 wire \vga_tetris.boardMem.board_18[5] ;
 wire \vga_tetris.boardMem.board_18[6] ;
 wire \vga_tetris.boardMem.board_18[7] ;
 wire \vga_tetris.boardMem.board_18[8] ;
 wire \vga_tetris.boardMem.board_18[9] ;
 wire \vga_tetris.boardMem.board_19[0] ;
 wire \vga_tetris.boardMem.board_19[10] ;
 wire \vga_tetris.boardMem.board_19[11] ;
 wire \vga_tetris.boardMem.board_19[12] ;
 wire \vga_tetris.boardMem.board_19[13] ;
 wire \vga_tetris.boardMem.board_19[14] ;
 wire \vga_tetris.boardMem.board_19[15] ;
 wire \vga_tetris.boardMem.board_19[16] ;
 wire \vga_tetris.boardMem.board_19[17] ;
 wire \vga_tetris.boardMem.board_19[18] ;
 wire \vga_tetris.boardMem.board_19[19] ;
 wire \vga_tetris.boardMem.board_19[1] ;
 wire \vga_tetris.boardMem.board_19[2] ;
 wire \vga_tetris.boardMem.board_19[3] ;
 wire \vga_tetris.boardMem.board_19[4] ;
 wire \vga_tetris.boardMem.board_19[5] ;
 wire \vga_tetris.boardMem.board_19[6] ;
 wire \vga_tetris.boardMem.board_19[7] ;
 wire \vga_tetris.boardMem.board_19[8] ;
 wire \vga_tetris.boardMem.board_19[9] ;
 wire \vga_tetris.boardMem.board_1[0] ;
 wire \vga_tetris.boardMem.board_1[10] ;
 wire \vga_tetris.boardMem.board_1[11] ;
 wire \vga_tetris.boardMem.board_1[12] ;
 wire \vga_tetris.boardMem.board_1[13] ;
 wire \vga_tetris.boardMem.board_1[14] ;
 wire \vga_tetris.boardMem.board_1[15] ;
 wire \vga_tetris.boardMem.board_1[16] ;
 wire \vga_tetris.boardMem.board_1[17] ;
 wire \vga_tetris.boardMem.board_1[18] ;
 wire \vga_tetris.boardMem.board_1[19] ;
 wire \vga_tetris.boardMem.board_1[1] ;
 wire \vga_tetris.boardMem.board_1[2] ;
 wire \vga_tetris.boardMem.board_1[3] ;
 wire \vga_tetris.boardMem.board_1[4] ;
 wire \vga_tetris.boardMem.board_1[5] ;
 wire \vga_tetris.boardMem.board_1[6] ;
 wire \vga_tetris.boardMem.board_1[7] ;
 wire \vga_tetris.boardMem.board_1[8] ;
 wire \vga_tetris.boardMem.board_1[9] ;
 wire \vga_tetris.boardMem.board_2[0] ;
 wire \vga_tetris.boardMem.board_2[10] ;
 wire \vga_tetris.boardMem.board_2[11] ;
 wire \vga_tetris.boardMem.board_2[12] ;
 wire \vga_tetris.boardMem.board_2[13] ;
 wire \vga_tetris.boardMem.board_2[14] ;
 wire \vga_tetris.boardMem.board_2[15] ;
 wire \vga_tetris.boardMem.board_2[16] ;
 wire \vga_tetris.boardMem.board_2[17] ;
 wire \vga_tetris.boardMem.board_2[18] ;
 wire \vga_tetris.boardMem.board_2[19] ;
 wire \vga_tetris.boardMem.board_2[1] ;
 wire \vga_tetris.boardMem.board_2[2] ;
 wire \vga_tetris.boardMem.board_2[3] ;
 wire \vga_tetris.boardMem.board_2[4] ;
 wire \vga_tetris.boardMem.board_2[5] ;
 wire \vga_tetris.boardMem.board_2[6] ;
 wire \vga_tetris.boardMem.board_2[7] ;
 wire \vga_tetris.boardMem.board_2[8] ;
 wire \vga_tetris.boardMem.board_2[9] ;
 wire \vga_tetris.boardMem.board_3[0] ;
 wire \vga_tetris.boardMem.board_3[10] ;
 wire \vga_tetris.boardMem.board_3[11] ;
 wire \vga_tetris.boardMem.board_3[12] ;
 wire \vga_tetris.boardMem.board_3[13] ;
 wire \vga_tetris.boardMem.board_3[14] ;
 wire \vga_tetris.boardMem.board_3[15] ;
 wire \vga_tetris.boardMem.board_3[16] ;
 wire \vga_tetris.boardMem.board_3[17] ;
 wire \vga_tetris.boardMem.board_3[18] ;
 wire \vga_tetris.boardMem.board_3[19] ;
 wire \vga_tetris.boardMem.board_3[1] ;
 wire \vga_tetris.boardMem.board_3[2] ;
 wire \vga_tetris.boardMem.board_3[3] ;
 wire \vga_tetris.boardMem.board_3[4] ;
 wire \vga_tetris.boardMem.board_3[5] ;
 wire \vga_tetris.boardMem.board_3[6] ;
 wire \vga_tetris.boardMem.board_3[7] ;
 wire \vga_tetris.boardMem.board_3[8] ;
 wire \vga_tetris.boardMem.board_3[9] ;
 wire \vga_tetris.boardMem.board_4[0] ;
 wire \vga_tetris.boardMem.board_4[10] ;
 wire \vga_tetris.boardMem.board_4[11] ;
 wire \vga_tetris.boardMem.board_4[12] ;
 wire \vga_tetris.boardMem.board_4[13] ;
 wire \vga_tetris.boardMem.board_4[14] ;
 wire \vga_tetris.boardMem.board_4[15] ;
 wire \vga_tetris.boardMem.board_4[16] ;
 wire \vga_tetris.boardMem.board_4[17] ;
 wire \vga_tetris.boardMem.board_4[18] ;
 wire \vga_tetris.boardMem.board_4[19] ;
 wire \vga_tetris.boardMem.board_4[1] ;
 wire \vga_tetris.boardMem.board_4[2] ;
 wire \vga_tetris.boardMem.board_4[3] ;
 wire \vga_tetris.boardMem.board_4[4] ;
 wire \vga_tetris.boardMem.board_4[5] ;
 wire \vga_tetris.boardMem.board_4[6] ;
 wire \vga_tetris.boardMem.board_4[7] ;
 wire \vga_tetris.boardMem.board_4[8] ;
 wire \vga_tetris.boardMem.board_4[9] ;
 wire \vga_tetris.boardMem.board_5[0] ;
 wire \vga_tetris.boardMem.board_5[10] ;
 wire \vga_tetris.boardMem.board_5[11] ;
 wire \vga_tetris.boardMem.board_5[12] ;
 wire \vga_tetris.boardMem.board_5[13] ;
 wire \vga_tetris.boardMem.board_5[14] ;
 wire \vga_tetris.boardMem.board_5[15] ;
 wire \vga_tetris.boardMem.board_5[16] ;
 wire \vga_tetris.boardMem.board_5[17] ;
 wire \vga_tetris.boardMem.board_5[18] ;
 wire \vga_tetris.boardMem.board_5[19] ;
 wire \vga_tetris.boardMem.board_5[1] ;
 wire \vga_tetris.boardMem.board_5[2] ;
 wire \vga_tetris.boardMem.board_5[3] ;
 wire \vga_tetris.boardMem.board_5[4] ;
 wire \vga_tetris.boardMem.board_5[5] ;
 wire \vga_tetris.boardMem.board_5[6] ;
 wire \vga_tetris.boardMem.board_5[7] ;
 wire \vga_tetris.boardMem.board_5[8] ;
 wire \vga_tetris.boardMem.board_5[9] ;
 wire \vga_tetris.boardMem.board_6[0] ;
 wire \vga_tetris.boardMem.board_6[10] ;
 wire \vga_tetris.boardMem.board_6[11] ;
 wire \vga_tetris.boardMem.board_6[12] ;
 wire \vga_tetris.boardMem.board_6[13] ;
 wire \vga_tetris.boardMem.board_6[14] ;
 wire \vga_tetris.boardMem.board_6[15] ;
 wire \vga_tetris.boardMem.board_6[16] ;
 wire \vga_tetris.boardMem.board_6[17] ;
 wire \vga_tetris.boardMem.board_6[18] ;
 wire \vga_tetris.boardMem.board_6[19] ;
 wire \vga_tetris.boardMem.board_6[1] ;
 wire \vga_tetris.boardMem.board_6[2] ;
 wire \vga_tetris.boardMem.board_6[3] ;
 wire \vga_tetris.boardMem.board_6[4] ;
 wire \vga_tetris.boardMem.board_6[5] ;
 wire \vga_tetris.boardMem.board_6[6] ;
 wire \vga_tetris.boardMem.board_6[7] ;
 wire \vga_tetris.boardMem.board_6[8] ;
 wire \vga_tetris.boardMem.board_6[9] ;
 wire \vga_tetris.boardMem.board_7[0] ;
 wire \vga_tetris.boardMem.board_7[10] ;
 wire \vga_tetris.boardMem.board_7[11] ;
 wire \vga_tetris.boardMem.board_7[12] ;
 wire \vga_tetris.boardMem.board_7[13] ;
 wire \vga_tetris.boardMem.board_7[14] ;
 wire \vga_tetris.boardMem.board_7[15] ;
 wire \vga_tetris.boardMem.board_7[16] ;
 wire \vga_tetris.boardMem.board_7[17] ;
 wire \vga_tetris.boardMem.board_7[18] ;
 wire \vga_tetris.boardMem.board_7[19] ;
 wire \vga_tetris.boardMem.board_7[1] ;
 wire \vga_tetris.boardMem.board_7[2] ;
 wire \vga_tetris.boardMem.board_7[3] ;
 wire \vga_tetris.boardMem.board_7[4] ;
 wire \vga_tetris.boardMem.board_7[5] ;
 wire \vga_tetris.boardMem.board_7[6] ;
 wire \vga_tetris.boardMem.board_7[7] ;
 wire \vga_tetris.boardMem.board_7[8] ;
 wire \vga_tetris.boardMem.board_7[9] ;
 wire \vga_tetris.boardMem.board_8[0] ;
 wire \vga_tetris.boardMem.board_8[10] ;
 wire \vga_tetris.boardMem.board_8[11] ;
 wire \vga_tetris.boardMem.board_8[12] ;
 wire \vga_tetris.boardMem.board_8[13] ;
 wire \vga_tetris.boardMem.board_8[14] ;
 wire \vga_tetris.boardMem.board_8[15] ;
 wire \vga_tetris.boardMem.board_8[16] ;
 wire \vga_tetris.boardMem.board_8[17] ;
 wire \vga_tetris.boardMem.board_8[18] ;
 wire \vga_tetris.boardMem.board_8[19] ;
 wire \vga_tetris.boardMem.board_8[1] ;
 wire \vga_tetris.boardMem.board_8[2] ;
 wire \vga_tetris.boardMem.board_8[3] ;
 wire \vga_tetris.boardMem.board_8[4] ;
 wire \vga_tetris.boardMem.board_8[5] ;
 wire \vga_tetris.boardMem.board_8[6] ;
 wire \vga_tetris.boardMem.board_8[7] ;
 wire \vga_tetris.boardMem.board_8[8] ;
 wire \vga_tetris.boardMem.board_8[9] ;
 wire \vga_tetris.boardMem.board_9[0] ;
 wire \vga_tetris.boardMem.board_9[10] ;
 wire \vga_tetris.boardMem.board_9[11] ;
 wire \vga_tetris.boardMem.board_9[12] ;
 wire \vga_tetris.boardMem.board_9[13] ;
 wire \vga_tetris.boardMem.board_9[14] ;
 wire \vga_tetris.boardMem.board_9[15] ;
 wire \vga_tetris.boardMem.board_9[16] ;
 wire \vga_tetris.boardMem.board_9[17] ;
 wire \vga_tetris.boardMem.board_9[18] ;
 wire \vga_tetris.boardMem.board_9[19] ;
 wire \vga_tetris.boardMem.board_9[1] ;
 wire \vga_tetris.boardMem.board_9[2] ;
 wire \vga_tetris.boardMem.board_9[3] ;
 wire \vga_tetris.boardMem.board_9[4] ;
 wire \vga_tetris.boardMem.board_9[5] ;
 wire \vga_tetris.boardMem.board_9[6] ;
 wire \vga_tetris.boardMem.board_9[7] ;
 wire \vga_tetris.boardMem.board_9[8] ;
 wire \vga_tetris.boardMem.board_9[9] ;
 wire \vga_tetris.inputs.buttonTimerQ_0[0] ;
 wire \vga_tetris.inputs.buttonTimerQ_0[1] ;
 wire \vga_tetris.inputs.buttonTimerQ_0[2] ;
 wire \vga_tetris.inputs.buttonTimerQ_0[3] ;
 wire \vga_tetris.inputs.buttonTimerQ_0[4] ;
 wire \vga_tetris.inputs.buttonTimerQ_0[5] ;
 wire \vga_tetris.inputs.buttonTimerQ_0[6] ;
 wire \vga_tetris.inputs.buttonTimerQ_0[7] ;
 wire \vga_tetris.inputs.buttonTimerQ_1[0] ;
 wire \vga_tetris.inputs.buttonTimerQ_1[1] ;
 wire \vga_tetris.inputs.buttonTimerQ_1[2] ;
 wire \vga_tetris.inputs.buttonTimerQ_1[3] ;
 wire \vga_tetris.inputs.buttonTimerQ_1[4] ;
 wire \vga_tetris.inputs.buttonTimerQ_1[5] ;
 wire \vga_tetris.inputs.buttonTimerQ_1[6] ;
 wire \vga_tetris.inputs.buttonTimerQ_1[7] ;
 wire \vga_tetris.inputs.buttonTimerQ_2[0] ;
 wire \vga_tetris.inputs.buttonTimerQ_2[1] ;
 wire \vga_tetris.inputs.buttonTimerQ_2[2] ;
 wire \vga_tetris.inputs.buttonTimerQ_2[3] ;
 wire \vga_tetris.inputs.buttonTimerQ_2[4] ;
 wire \vga_tetris.inputs.buttonTimerQ_2[5] ;
 wire \vga_tetris.inputs.buttonTimerQ_2[6] ;
 wire \vga_tetris.inputs.buttonTimerQ_2[7] ;
 wire \vga_tetris.inputs.buttonTimerQ_3[0] ;
 wire \vga_tetris.inputs.buttonTimerQ_3[1] ;
 wire \vga_tetris.inputs.buttonTimerQ_3[2] ;
 wire \vga_tetris.inputs.buttonTimerQ_3[3] ;
 wire \vga_tetris.inputs.buttonTimerQ_3[4] ;
 wire \vga_tetris.inputs.buttonTimerQ_3[5] ;
 wire \vga_tetris.inputs.buttonTimerQ_3[6] ;
 wire \vga_tetris.inputs.buttonTimerQ_3[7] ;
 wire \vga_tetris.msTimer.msTimerQ[0] ;
 wire \vga_tetris.msTimer.msTimerQ[10] ;
 wire \vga_tetris.msTimer.msTimerQ[11] ;
 wire \vga_tetris.msTimer.msTimerQ[12] ;
 wire \vga_tetris.msTimer.msTimerQ[13] ;
 wire \vga_tetris.msTimer.msTimerQ[14] ;
 wire \vga_tetris.msTimer.msTimerQ[1] ;
 wire \vga_tetris.msTimer.msTimerQ[2] ;
 wire \vga_tetris.msTimer.msTimerQ[3] ;
 wire \vga_tetris.msTimer.msTimerQ[4] ;
 wire \vga_tetris.msTimer.msTimerQ[5] ;
 wire \vga_tetris.msTimer.msTimerQ[6] ;
 wire \vga_tetris.msTimer.msTimerQ[7] ;
 wire \vga_tetris.msTimer.msTimerQ[8] ;
 wire \vga_tetris.msTimer.msTimerQ[9] ;
 wire \vga_tetris.runningTetrisLogicQ ;
 wire \vga_tetris.startTetrisLogicQ ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[0] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[10] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[11] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[12] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[13] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[14] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[15] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[16] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[17] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[18] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[19] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[1] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[2] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[3] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[4] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[5] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[6] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[7] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[8] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[9] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_done ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_rowIndex[0] ;
 wire \vga_tetris.tetrisLogic._addOrRemoveShape_io_rowIndex[1] ;
 wire \vga_tetris.tetrisLogic._checkMoveAllowed_io_checkDone ;
 wire \vga_tetris.tetrisLogic._checkMoveAllowed_io_rowIndex[0] ;
 wire \vga_tetris.tetrisLogic._checkMoveAllowed_io_rowIndex[1] ;
 wire \vga_tetris.tetrisLogic.addOrRemoveShape.clearingQ ;
 wire \vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[0] ;
 wire \vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[1] ;
 wire \vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[2] ;
 wire \vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[3] ;
 wire \vga_tetris.tetrisLogic.addOrRemoveShape.stateQ[0] ;
 wire \vga_tetris.tetrisLogic.addOrRemoveShape.stateQ[1] ;
 wire \vga_tetris.tetrisLogic.adderSubtracter.io_a[0] ;
 wire \vga_tetris.tetrisLogic.adderSubtracter.io_a[1] ;
 wire \vga_tetris.tetrisLogic.adderSubtracter.io_a[2] ;
 wire \vga_tetris.tetrisLogic.adderSubtracter.io_a[3] ;
 wire \vga_tetris.tetrisLogic.adderSubtracter.io_a[4] ;
 wire \vga_tetris.tetrisLogic.checkMoveAllowed.checkIsRunningQ ;
 wire \vga_tetris.tetrisLogic.gameOverLogic.buttonPressesCounterQ[0] ;
 wire \vga_tetris.tetrisLogic.gameOverLogic.buttonPressesCounterQ[1] ;
 wire \vga_tetris.tetrisLogic.gameOverResetHappenedQ ;
 wire \vga_tetris.tetrisLogic.rotationQ[0] ;
 wire \vga_tetris.tetrisLogic.rotationQ[1] ;
 wire \vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[0] ;
 wire \vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[1] ;
 wire \vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[2] ;
 wire \vga_tetris.tetrisLogic.shapeDropTimerQ[0] ;
 wire \vga_tetris.tetrisLogic.shapeDropTimerQ[1] ;
 wire \vga_tetris.tetrisLogic.shapeDropTimerQ[2] ;
 wire \vga_tetris.tetrisLogic.shapeDropTimerQ[3] ;
 wire \vga_tetris.tetrisLogic.shapeDropTimerQ[4] ;
 wire \vga_tetris.tetrisLogic.shapeDropTimerQ[5] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[0] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[10] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[11] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[12] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[13] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[14] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[15] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[16] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[17] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[18] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[19] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[1] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[2] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[3] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[4] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[5] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[6] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[7] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[8] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[9] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.internalStartTriggerQ ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[0] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[1] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[2] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[3] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[4] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.operationIsRunningQ ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[0] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[1] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[2] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[3] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[4] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[0] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[1] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[2] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[3] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[4] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.stateQ[0] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.stateQ[1] ;
 wire \vga_tetris.tetrisLogic.shiftTheBoard.stateQ[2] ;
 wire \vga_tetris.tetrisLogic.stateQ[0] ;
 wire \vga_tetris.tetrisLogic.stateQ[1] ;
 wire \vga_tetris.tetrisLogic.stateQ[2] ;
 wire \vga_tetris.tetrisLogic.stateQ[3] ;
 wire \vga_tetris.tetrisLogic.stateQ[4] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[0] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[10] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[11] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[12] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[13] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[14] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[15] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[1] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[2] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[3] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[4] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[5] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[6] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[7] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[8] ;
 wire \vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[9] ;
 wire \vga_tetris.vgaController.horizontalCounterQ[0] ;
 wire \vga_tetris.vgaController.horizontalCounterQ[1] ;
 wire \vga_tetris.vgaController.horizontalCounterQ[2] ;
 wire \vga_tetris.vgaController.horizontalCounterQ[3] ;
 wire \vga_tetris.vgaController.horizontalCounterQ[4] ;
 wire \vga_tetris.vgaController.horizontalCounterQ[5] ;
 wire \vga_tetris.vgaController.horizontalCounterQ[6] ;
 wire \vga_tetris.vgaController.horizontalCounterQ[7] ;
 wire \vga_tetris.vgaController.horizontalCounterQ[8] ;
 wire \vga_tetris.vgaController.horizontalCounterQ[9] ;
 wire \vga_tetris.vgaController.verticalCounterQ[0] ;
 wire \vga_tetris.vgaController.verticalCounterQ[1] ;
 wire \vga_tetris.vgaController.verticalCounterQ[2] ;
 wire \vga_tetris.vgaController.verticalCounterQ[3] ;
 wire \vga_tetris.vgaController.verticalCounterQ[4] ;
 wire \vga_tetris.vgaController.verticalCounterQ[5] ;
 wire \vga_tetris.vgaController.verticalCounterQ[6] ;
 wire \vga_tetris.vgaController.verticalCounterQ[7] ;
 wire \vga_tetris.vgaController.verticalCounterQ[8] ;
 wire \vga_tetris.vgaController.verticalCounterQ[9] ;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;

 sg13g2_inv_2 _3561_ (.Y(_0624_),
    .A(net1667));
 sg13g2_inv_1 _3562_ (.Y(_0625_),
    .A(net1703));
 sg13g2_inv_1 _3563_ (.Y(_0626_),
    .A(\vga_tetris._vgaController_io_pixelPosX[9] ));
 sg13g2_inv_2 _3564_ (.Y(_0627_),
    .A(\vga_tetris._vgaController_io_pixelPosX[3] ));
 sg13g2_inv_2 _3565_ (.Y(_0628_),
    .A(net1198));
 sg13g2_inv_1 _3566_ (.Y(_0629_),
    .A(net1826));
 sg13g2_inv_1 _3567_ (.Y(_0630_),
    .A(net1602));
 sg13g2_inv_1 _3568_ (.Y(_0631_),
    .A(net1593));
 sg13g2_inv_1 _3569_ (.Y(_0632_),
    .A(net1411));
 sg13g2_inv_1 _3570_ (.Y(_0633_),
    .A(net1327));
 sg13g2_inv_1 _3571_ (.Y(_0634_),
    .A(net1273));
 sg13g2_inv_1 _3572_ (.Y(_0635_),
    .A(net831));
 sg13g2_inv_1 _3573_ (.Y(_0636_),
    .A(net1404));
 sg13g2_inv_1 _3574_ (.Y(_0637_),
    .A(net1706));
 sg13g2_inv_2 _3575_ (.Y(_0638_),
    .A(net1604));
 sg13g2_inv_1 _3576_ (.Y(_0639_),
    .A(net1552));
 sg13g2_inv_1 _3577_ (.Y(_0640_),
    .A(net1651));
 sg13g2_inv_1 _3578_ (.Y(_0641_),
    .A(net1287));
 sg13g2_inv_1 _3579_ (.Y(_0642_),
    .A(net1357));
 sg13g2_inv_1 _3580_ (.Y(_0643_),
    .A(net1626));
 sg13g2_inv_1 _3581_ (.Y(_0644_),
    .A(net1401));
 sg13g2_inv_1 _3582_ (.Y(_0645_),
    .A(net1349));
 sg13g2_inv_1 _3583_ (.Y(_0646_),
    .A(net1305));
 sg13g2_inv_1 _3584_ (.Y(_0647_),
    .A(net1382));
 sg13g2_inv_1 _3585_ (.Y(_0648_),
    .A(net1483));
 sg13g2_inv_1 _3586_ (.Y(_0649_),
    .A(net1365));
 sg13g2_inv_1 _3587_ (.Y(_0650_),
    .A(net1295));
 sg13g2_inv_1 _3588_ (.Y(_0651_),
    .A(net1595));
 sg13g2_inv_1 _3589_ (.Y(_0652_),
    .A(net1583));
 sg13g2_inv_1 _3590_ (.Y(_0653_),
    .A(net1206));
 sg13g2_inv_2 _3591_ (.Y(_0654_),
    .A(net1209));
 sg13g2_inv_2 _3592_ (.Y(_0655_),
    .A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[3] ));
 sg13g2_inv_1 _3593_ (.Y(_0656_),
    .A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[2] ));
 sg13g2_inv_1 _3594_ (.Y(_0657_),
    .A(net1400));
 sg13g2_inv_4 _3595_ (.A(net1217),
    .Y(_0658_));
 sg13g2_inv_2 _3596_ (.Y(_0659_),
    .A(net1202));
 sg13g2_inv_1 _3597_ (.Y(_0660_),
    .A(net1806));
 sg13g2_inv_2 _3598_ (.Y(_0661_),
    .A(net1810));
 sg13g2_inv_2 _3599_ (.Y(_0662_),
    .A(net1177));
 sg13g2_inv_1 _3600_ (.Y(_0663_),
    .A(net1539));
 sg13g2_inv_1 _3601_ (.Y(_0664_),
    .A(net648));
 sg13g2_inv_1 _3602_ (.Y(_0665_),
    .A(net1433));
 sg13g2_inv_1 _3603_ (.Y(_0666_),
    .A(net1470));
 sg13g2_inv_1 _3604_ (.Y(_0667_),
    .A(\vga_tetris.boardMem.board_0[9] ));
 sg13g2_inv_1 _3605_ (.Y(_0668_),
    .A(net1530));
 sg13g2_inv_1 _3606_ (.Y(_0669_),
    .A(net1490));
 sg13g2_inv_1 _3607_ (.Y(_0670_),
    .A(\vga_tetris.boardMem.board_0[12] ));
 sg13g2_inv_1 _3608_ (.Y(_0671_),
    .A(\vga_tetris.boardMem.board_0[13] ));
 sg13g2_inv_1 _3609_ (.Y(_0672_),
    .A(net1510));
 sg13g2_inv_1 _3610_ (.Y(_0673_),
    .A(net1398));
 sg13g2_inv_1 _3611_ (.Y(_0674_),
    .A(net1555));
 sg13g2_inv_1 _3612_ (.Y(_0675_),
    .A(\vga_tetris.msTimer.msTimerQ[2] ));
 sg13g2_inv_1 _3613_ (.Y(_0676_),
    .A(\vga_tetris.msTimer.msTimerQ[5] ));
 sg13g2_inv_1 _3614_ (.Y(_0677_),
    .A(\vga_tetris._inputs_io_rightButtonActive ));
 sg13g2_inv_1 _3615_ (.Y(_0678_),
    .A(net804));
 sg13g2_inv_2 _3616_ (.Y(_0679_),
    .A(net1589));
 sg13g2_inv_1 _3617_ (.Y(_0680_),
    .A(net1842));
 sg13g2_inv_1 _3618_ (.Y(_0681_),
    .A(net1836));
 sg13g2_inv_4 _3619_ (.A(net1213),
    .Y(_0682_));
 sg13g2_inv_1 _3620_ (.Y(_0683_),
    .A(net1684));
 sg13g2_inv_4 _3621_ (.A(net1235),
    .Y(_0684_));
 sg13g2_inv_1 _3622_ (.Y(_0685_),
    .A(net1770));
 sg13g2_inv_1 _3623_ (.Y(_0686_),
    .A(net1829));
 sg13g2_inv_1 _3624_ (.Y(_0687_),
    .A(net1846));
 sg13g2_inv_1 _3625_ (.Y(_0688_),
    .A(net1660));
 sg13g2_inv_2 _3626_ (.Y(_0689_),
    .A(net1804));
 sg13g2_inv_1 _3627_ (.Y(_0690_),
    .A(net1813));
 sg13g2_inv_1 _3628_ (.Y(_0691_),
    .A(net1759));
 sg13g2_inv_1 _3629_ (.Y(_0692_),
    .A(net1753));
 sg13g2_inv_1 _3630_ (.Y(_0693_),
    .A(\vga_tetris._tetrisLogic_io_score_0[2] ));
 sg13g2_inv_1 _3631_ (.Y(_0694_),
    .A(net1686));
 sg13g2_inv_1 _3632_ (.Y(_0695_),
    .A(net1820));
 sg13g2_inv_1 _3633_ (.Y(_0696_),
    .A(net1816));
 sg13g2_nor2b_2 _3634_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[0] ),
    .B_N(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[2] ),
    .Y(_0697_));
 sg13g2_nor2b_2 _3635_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[1] ),
    .B_N(_0697_),
    .Y(_0698_));
 sg13g2_nand2b_1 _3636_ (.Y(_0699_),
    .B(_0697_),
    .A_N(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[1] ));
 sg13g2_nor2b_1 _3637_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[2] ),
    .B_N(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[1] ),
    .Y(_0700_));
 sg13g2_nand2b_1 _3638_ (.Y(_0701_),
    .B(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[1] ),
    .A_N(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[2] ));
 sg13g2_and2_1 _3639_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[0] ),
    .B(_0700_),
    .X(_0702_));
 sg13g2_nand2_1 _3640_ (.Y(_0703_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[0] ),
    .B(_0700_));
 sg13g2_nand2_1 _3641_ (.Y(_0704_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[4] ),
    .B(net1168));
 sg13g2_o21ai_1 _3642_ (.B1(_0704_),
    .Y(_0705_),
    .A1(_0660_),
    .A2(net1168));
 sg13g2_nor2b_1 _3643_ (.A(net1206),
    .B_N(\vga_tetris.tetrisLogic.stateQ[3] ),
    .Y(_0706_));
 sg13g2_nand3b_1 _3644_ (.B(\vga_tetris.tetrisLogic.stateQ[2] ),
    .C(\vga_tetris.tetrisLogic.stateQ[3] ),
    .Y(_0707_),
    .A_N(net1206));
 sg13g2_nand2_2 _3645_ (.Y(_0708_),
    .A(net1215),
    .B(_0658_));
 sg13g2_nor2_2 _3646_ (.A(_0707_),
    .B(_0708_),
    .Y(_0709_));
 sg13g2_or2_1 _3647_ (.X(_0710_),
    .B(_0708_),
    .A(_0707_));
 sg13g2_o21ai_1 _3648_ (.B1(_0709_),
    .Y(_0711_),
    .A1(_0637_),
    .A2(net1173));
 sg13g2_a21oi_1 _3649_ (.A1(net1173),
    .A2(_0705_),
    .Y(_0712_),
    .B1(_0711_));
 sg13g2_nor2_2 _3650_ (.A(net1216),
    .B(net1217),
    .Y(_0713_));
 sg13g2_inv_1 _3651_ (.Y(_0714_),
    .A(_0713_));
 sg13g2_nor2_1 _3652_ (.A(\vga_tetris.tetrisLogic.stateQ[2] ),
    .B(\vga_tetris.tetrisLogic.stateQ[3] ),
    .Y(_0715_));
 sg13g2_and2_1 _3653_ (.A(net1205),
    .B(_0715_),
    .X(_0716_));
 sg13g2_nand2_1 _3654_ (.Y(_0717_),
    .A(net1205),
    .B(_0715_));
 sg13g2_nand3_1 _3655_ (.B(_0713_),
    .C(_0715_),
    .A(net1205),
    .Y(_0718_));
 sg13g2_nor2b_1 _3656_ (.A(\vga_tetris.tetrisLogic.stateQ[2] ),
    .B_N(_0706_),
    .Y(_0719_));
 sg13g2_nand2b_2 _3657_ (.Y(_0720_),
    .B(_0706_),
    .A_N(\vga_tetris.tetrisLogic.stateQ[2] ));
 sg13g2_nor2b_2 _3658_ (.A(net1215),
    .B_N(net1217),
    .Y(_0721_));
 sg13g2_and2_1 _3659_ (.A(_0719_),
    .B(_0721_),
    .X(_0722_));
 sg13g2_nand3_1 _3660_ (.B(_0715_),
    .C(_0721_),
    .A(net1205),
    .Y(_0723_));
 sg13g2_nand2_2 _3661_ (.Y(_0724_),
    .A(net1215),
    .B(\vga_tetris.tetrisLogic.stateQ[0] ));
 sg13g2_o21ai_1 _3662_ (.B1(_0723_),
    .Y(_0725_),
    .A1(_0720_),
    .A2(_0724_));
 sg13g2_nor2b_1 _3663_ (.A(\vga_tetris.tetrisLogic.stateQ[3] ),
    .B_N(\vga_tetris.tetrisLogic.stateQ[2] ),
    .Y(_0726_));
 sg13g2_nand2b_1 _3664_ (.Y(_0727_),
    .B(\vga_tetris.tetrisLogic.stateQ[2] ),
    .A_N(\vga_tetris.tetrisLogic.stateQ[3] ));
 sg13g2_nor2_1 _3665_ (.A(net1205),
    .B(_0727_),
    .Y(_0728_));
 sg13g2_nand3_1 _3666_ (.B(net1216),
    .C(_0726_),
    .A(_0653_),
    .Y(_0729_));
 sg13g2_o21ai_1 _3667_ (.B1(_0729_),
    .Y(_0730_),
    .A1(_0714_),
    .A2(_0720_));
 sg13g2_and4_1 _3668_ (.A(_0718_),
    .B(_0720_),
    .C(_0723_),
    .D(_0729_),
    .X(_0731_));
 sg13g2_nor4_2 _3669_ (.A(net1205),
    .B(net1215),
    .C(net1217),
    .Y(_0732_),
    .D(_0727_));
 sg13g2_nand3_1 _3670_ (.B(_0713_),
    .C(_0726_),
    .A(_0653_),
    .Y(_0733_));
 sg13g2_nor2_2 _3671_ (.A(net1215),
    .B(_0707_),
    .Y(_0734_));
 sg13g2_or2_1 _3672_ (.X(_0735_),
    .B(_0707_),
    .A(net1216));
 sg13g2_nor2_2 _3673_ (.A(_0732_),
    .B(_0734_),
    .Y(_0736_));
 sg13g2_nand3_1 _3674_ (.B(_0733_),
    .C(_0735_),
    .A(\vga_tetris.tetrisLogic._checkMoveAllowed_io_rowIndex[1] ),
    .Y(_0737_));
 sg13g2_o21ai_1 _3675_ (.B1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_rowIndex[1] ),
    .Y(_0738_),
    .A1(_0732_),
    .A2(_0734_));
 sg13g2_o21ai_1 _3676_ (.B1(_0738_),
    .Y(_0739_),
    .A1(_0731_),
    .A2(_0737_));
 sg13g2_and2_1 _3677_ (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[1] ),
    .B(_0739_),
    .X(_0740_));
 sg13g2_nand3_1 _3678_ (.B(_0733_),
    .C(_0735_),
    .A(\vga_tetris.tetrisLogic._checkMoveAllowed_io_rowIndex[0] ),
    .Y(_0741_));
 sg13g2_o21ai_1 _3679_ (.B1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_rowIndex[0] ),
    .Y(_0742_),
    .A1(_0732_),
    .A2(_0734_));
 sg13g2_o21ai_1 _3680_ (.B1(_0742_),
    .Y(_0743_),
    .A1(_0731_),
    .A2(_0741_));
 sg13g2_and2_1 _3681_ (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[0] ),
    .B(_0743_),
    .X(_0744_));
 sg13g2_xor2_1 _3682_ (.B(_0739_),
    .A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[1] ),
    .X(_0745_));
 sg13g2_a21oi_2 _3683_ (.B1(_0740_),
    .Y(_0746_),
    .A2(_0745_),
    .A1(_0744_));
 sg13g2_nand3b_1 _3684_ (.B(\vga_tetris.tetrisLogic.adderSubtracter.io_a[2] ),
    .C(\vga_tetris.tetrisLogic.adderSubtracter.io_a[3] ),
    .Y(_0747_),
    .A_N(_0746_));
 sg13g2_xor2_1 _3685_ (.B(_0747_),
    .A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[4] ),
    .X(_0748_));
 sg13g2_a21oi_2 _3686_ (.B1(_0712_),
    .Y(_0749_),
    .A2(_0748_),
    .A1(net1150));
 sg13g2_a21o_2 _3687_ (.A2(_0748_),
    .A1(net1150),
    .B1(_0712_),
    .X(_0750_));
 sg13g2_mux2_1 _3688_ (.A0(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[3] ),
    .A1(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[3] ),
    .S(net1168),
    .X(_0751_));
 sg13g2_a21oi_1 _3689_ (.A1(_0638_),
    .A2(_0698_),
    .Y(_0752_),
    .B1(net1150));
 sg13g2_o21ai_1 _3690_ (.B1(_0752_),
    .Y(_0753_),
    .A1(net1174),
    .A2(_0751_));
 sg13g2_o21ai_1 _3691_ (.B1(_0655_),
    .Y(_0754_),
    .A1(_0656_),
    .A2(_0746_));
 sg13g2_nand3_1 _3692_ (.B(_0747_),
    .C(_0754_),
    .A(net1150),
    .Y(_0755_));
 sg13g2_xnor2_1 _3693_ (.Y(_0756_),
    .A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[2] ),
    .B(_0746_));
 sg13g2_nor2_1 _3694_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[2] ),
    .B(_0703_),
    .Y(_0757_));
 sg13g2_o21ai_1 _3695_ (.B1(net1173),
    .Y(_0758_),
    .A1(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[2] ),
    .A2(net1168));
 sg13g2_a21oi_1 _3696_ (.A1(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[2] ),
    .A2(net1174),
    .Y(_0759_),
    .B1(net1150));
 sg13g2_o21ai_1 _3697_ (.B1(_0759_),
    .Y(_0760_),
    .A1(_0757_),
    .A2(_0758_));
 sg13g2_o21ai_1 _3698_ (.B1(_0760_),
    .Y(_0761_),
    .A1(_0709_),
    .A2(_0756_));
 sg13g2_and3_2 _3699_ (.X(_0762_),
    .A(_0753_),
    .B(_0755_),
    .C(_0761_));
 sg13g2_nand3_1 _3700_ (.B(_0755_),
    .C(_0761_),
    .A(_0753_),
    .Y(_0763_));
 sg13g2_nand2_1 _3701_ (.Y(_0764_),
    .A(_0749_),
    .B(_0763_));
 sg13g2_nand3_1 _3702_ (.B(_0749_),
    .C(_0763_),
    .A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[2] ),
    .Y(_0765_));
 sg13g2_nand2b_2 _3703_ (.Y(_0766_),
    .B(_0750_),
    .A_N(_0761_));
 sg13g2_nand2_2 _3704_ (.Y(_0767_),
    .A(_0765_),
    .B(_0766_));
 sg13g2_nand3_1 _3705_ (.B(_0765_),
    .C(_0766_),
    .A(net1177),
    .Y(_0768_));
 sg13g2_nand2_2 _3706_ (.Y(_0769_),
    .A(net1179),
    .B(net1175));
 sg13g2_or2_1 _3707_ (.X(_0770_),
    .B(net1177),
    .A(net1179));
 sg13g2_a21o_1 _3708_ (.A2(_0766_),
    .A1(_0765_),
    .B1(net1175),
    .X(_0771_));
 sg13g2_o21ai_1 _3709_ (.B1(_0749_),
    .Y(_0772_),
    .A1(\vga_tetris.tetrisLogic.adderSubtracter.io_a[4] ),
    .A2(_0762_));
 sg13g2_inv_1 _3710_ (.Y(_0773_),
    .A(_0772_));
 sg13g2_or2_1 _3711_ (.X(_0774_),
    .B(net1179),
    .A(\vga_tetris._vgaController_io_pixelPosY[7] ));
 sg13g2_nor2_2 _3712_ (.A(\vga_tetris._vgaController_io_pixelPosY[8] ),
    .B(_0774_),
    .Y(_0775_));
 sg13g2_and2_1 _3713_ (.A(\vga_tetris._vgaController_io_pixelPosY[8] ),
    .B(\vga_tetris._vgaController_io_pixelPosY[6] ),
    .X(_0776_));
 sg13g2_and2_1 _3714_ (.A(\vga_tetris._vgaController_io_pixelPosY[8] ),
    .B(\vga_tetris._vgaController_io_pixelPosY[7] ),
    .X(_0777_));
 sg13g2_nor4_1 _3715_ (.A(net1177),
    .B(_0775_),
    .C(_0776_),
    .D(_0777_),
    .Y(_0778_));
 sg13g2_a21oi_2 _3716_ (.B1(_0778_),
    .Y(_0779_),
    .A2(_0772_),
    .A1(net1177));
 sg13g2_a21o_1 _3717_ (.A2(_0772_),
    .A1(net1177),
    .B1(_0778_),
    .X(_0780_));
 sg13g2_nand2_2 _3718_ (.Y(_0781_),
    .A(net1703),
    .B(net1179));
 sg13g2_a21o_1 _3719_ (.A2(_0781_),
    .A1(_0774_),
    .B1(net1177),
    .X(_0782_));
 sg13g2_a21oi_1 _3720_ (.A1(_0753_),
    .A2(_0755_),
    .Y(_0783_),
    .B1(_0749_));
 sg13g2_nor3_1 _3721_ (.A(_0655_),
    .B(_0750_),
    .C(_0762_),
    .Y(_0784_));
 sg13g2_or2_1 _3722_ (.X(_0785_),
    .B(_0784_),
    .A(_0783_));
 sg13g2_o21ai_1 _3723_ (.B1(net1178),
    .Y(_0786_),
    .A1(_0783_),
    .A2(_0784_));
 sg13g2_nand3_1 _3724_ (.B(_0774_),
    .C(_0781_),
    .A(net1175),
    .Y(_0787_));
 sg13g2_or3_1 _3725_ (.A(net1175),
    .B(_0783_),
    .C(_0784_),
    .X(_0788_));
 sg13g2_a221oi_1 _3726_ (.B2(_0786_),
    .C1(_0779_),
    .B1(_0782_),
    .A1(_0768_),
    .Y(_0789_),
    .A2(_0769_));
 sg13g2_xnor2_1 _3727_ (.Y(_0790_),
    .A(_0657_),
    .B(_0743_));
 sg13g2_a21oi_1 _3728_ (.A1(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[0] ),
    .A2(net1174),
    .Y(_0791_),
    .B1(net1150));
 sg13g2_nand2_1 _3729_ (.Y(_0792_),
    .A(_0661_),
    .B(net1168));
 sg13g2_o21ai_1 _3730_ (.B1(_0792_),
    .Y(_0793_),
    .A1(net1201),
    .A2(net1168));
 sg13g2_o21ai_1 _3731_ (.B1(_0791_),
    .Y(_0794_),
    .A1(net1174),
    .A2(_0793_));
 sg13g2_o21ai_1 _3732_ (.B1(_0794_),
    .Y(_0795_),
    .A1(_0709_),
    .A2(_0790_));
 sg13g2_inv_1 _3733_ (.Y(_0796_),
    .A(_0795_));
 sg13g2_nand3_1 _3734_ (.B(_0749_),
    .C(_0763_),
    .A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[0] ),
    .Y(_0797_));
 sg13g2_o21ai_1 _3735_ (.B1(_0796_),
    .Y(_0798_),
    .A1(_0750_),
    .A2(_0762_));
 sg13g2_nand2_2 _3736_ (.Y(_0799_),
    .A(_0797_),
    .B(_0798_));
 sg13g2_and2_1 _3737_ (.A(_0797_),
    .B(_0798_),
    .X(_0800_));
 sg13g2_nand3_1 _3738_ (.B(_0797_),
    .C(_0798_),
    .A(net1178),
    .Y(_0801_));
 sg13g2_nor2_1 _3739_ (.A(net1184),
    .B(net1178),
    .Y(_0802_));
 sg13g2_or2_1 _3740_ (.X(_0803_),
    .B(net1178),
    .A(net1184));
 sg13g2_xor2_1 _3741_ (.B(_0745_),
    .A(_0744_),
    .X(_0804_));
 sg13g2_nor2_1 _3742_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[1] ),
    .B(_0703_),
    .Y(_0805_));
 sg13g2_nor2_1 _3743_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[1] ),
    .B(net1169),
    .Y(_0806_));
 sg13g2_a21oi_1 _3744_ (.A1(_0640_),
    .A2(net1174),
    .Y(_0807_),
    .B1(net1150));
 sg13g2_o21ai_1 _3745_ (.B1(net1173),
    .Y(_0808_),
    .A1(_0805_),
    .A2(_0806_));
 sg13g2_a22oi_1 _3746_ (.Y(_0809_),
    .B1(_0807_),
    .B2(_0808_),
    .A2(_0804_),
    .A1(net1150));
 sg13g2_inv_1 _3747_ (.Y(_0810_),
    .A(_0809_));
 sg13g2_a21oi_2 _3748_ (.B1(_0810_),
    .Y(_0811_),
    .A2(_0763_),
    .A1(_0749_));
 sg13g2_nor3_2 _3749_ (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[1] ),
    .B(_0750_),
    .C(_0762_),
    .Y(_0812_));
 sg13g2_nor2_2 _3750_ (.A(_0811_),
    .B(_0812_),
    .Y(_0813_));
 sg13g2_nand2_1 _3751_ (.Y(_0814_),
    .A(net1181),
    .B(net1175));
 sg13g2_nor3_1 _3752_ (.A(_0662_),
    .B(_0811_),
    .C(_0812_),
    .Y(_0815_));
 sg13g2_or3_1 _3753_ (.A(_0662_),
    .B(_0811_),
    .C(_0812_),
    .X(_0816_));
 sg13g2_a221oi_1 _3754_ (.B2(_0816_),
    .C1(_0802_),
    .B1(_0814_),
    .A1(net1178),
    .Y(_0817_),
    .A2(_0800_));
 sg13g2_and2_1 _3755_ (.A(net1054),
    .B(net1048),
    .X(_0818_));
 sg13g2_a22oi_1 _3756_ (.Y(_0819_),
    .B1(_0787_),
    .B2(_0788_),
    .A2(_0769_),
    .A1(_0768_));
 sg13g2_a221oi_1 _3757_ (.B2(_0788_),
    .C1(_0779_),
    .B1(_0787_),
    .A1(_0768_),
    .Y(_0820_),
    .A2(_0769_));
 sg13g2_and2_1 _3758_ (.A(net1050),
    .B(net1044),
    .X(_0821_));
 sg13g2_nand3_1 _3759_ (.B(net1048),
    .C(net1042),
    .A(\vga_tetris.boardMem.board_3[16] ),
    .Y(_0822_));
 sg13g2_and4_1 _3760_ (.A(_0801_),
    .B(_0803_),
    .C(_0814_),
    .D(_0816_),
    .X(_0823_));
 sg13g2_a221oi_1 _3761_ (.B2(_0786_),
    .C1(_0779_),
    .B1(_0782_),
    .A1(_0770_),
    .Y(_0824_),
    .A2(_0771_));
 sg13g2_and2_1 _3762_ (.A(net1035),
    .B(net1030),
    .X(_0825_));
 sg13g2_nand3_1 _3763_ (.B(net1035),
    .C(net1029),
    .A(\vga_tetris.boardMem.board_13[16] ),
    .Y(_0826_));
 sg13g2_and2_1 _3764_ (.A(net1055),
    .B(net1036),
    .X(_0827_));
 sg13g2_a221oi_1 _3765_ (.B2(_0788_),
    .C1(_0780_),
    .B1(_0787_),
    .A1(_0768_),
    .Y(_0828_),
    .A2(_0769_));
 sg13g2_nand2_1 _3766_ (.Y(_0829_),
    .A(_0779_),
    .B(_0819_));
 sg13g2_a221oi_1 _3767_ (.B2(_0803_),
    .C1(_0815_),
    .B1(_0801_),
    .A1(net1181),
    .Y(_0830_),
    .A2(_0662_));
 sg13g2_a21o_1 _3768_ (.A2(net1019),
    .A1(_0819_),
    .B1(_0779_),
    .X(_0831_));
 sg13g2_and2_1 _3769_ (.A(net995),
    .B(net993),
    .X(_0832_));
 sg13g2_nand2_1 _3770_ (.Y(_0833_),
    .A(net995),
    .B(net994));
 sg13g2_and2_1 _3771_ (.A(net1030),
    .B(net1019),
    .X(_0834_));
 sg13g2_nand3_1 _3772_ (.B(net1029),
    .C(net1018),
    .A(\vga_tetris.boardMem.board_12[16] ),
    .Y(_0835_));
 sg13g2_a22oi_1 _3773_ (.Y(_0836_),
    .B1(_0814_),
    .B2(_0816_),
    .A2(_0803_),
    .A1(_0801_));
 sg13g2_and2_1 _3774_ (.A(net1026),
    .B(net1013),
    .X(_0837_));
 sg13g2_nand3_1 _3775_ (.B(net1024),
    .C(net1011),
    .A(\vga_tetris.boardMem.board_18[16] ),
    .Y(_0838_));
 sg13g2_and2_1 _3776_ (.A(net1049),
    .B(net1030),
    .X(_0839_));
 sg13g2_nand3_1 _3777_ (.B(net1048),
    .C(net1029),
    .A(\vga_tetris.boardMem.board_15[16] ),
    .Y(_0840_));
 sg13g2_and2_1 _3778_ (.A(net1055),
    .B(net1012),
    .X(_0841_));
 sg13g2_and2_1 _3779_ (.A(net1049),
    .B(net1025),
    .X(_0842_));
 sg13g2_and2_1 _3780_ (.A(net1023),
    .B(net1017),
    .X(_0843_));
 sg13g2_a221oi_1 _3781_ (.B2(_0788_),
    .C1(_0779_),
    .B1(_0787_),
    .A1(_0770_),
    .Y(_0844_),
    .A2(_0771_));
 sg13g2_and2_1 _3782_ (.A(net1012),
    .B(net1004),
    .X(_0845_));
 sg13g2_and2_1 _3783_ (.A(net1018),
    .B(net1004),
    .X(_0846_));
 sg13g2_and3_1 _3784_ (.X(_0847_),
    .A(\vga_tetris.boardMem.board_4[16] ),
    .B(net1018),
    .C(net1004));
 sg13g2_and2_1 _3785_ (.A(net1053),
    .B(net1019),
    .X(_0848_));
 sg13g2_nand3_1 _3786_ (.B(net1054),
    .C(net1018),
    .A(\vga_tetris.boardMem.board_8[16] ),
    .Y(_0849_));
 sg13g2_and2_1 _3787_ (.A(net1042),
    .B(net1011),
    .X(_0850_));
 sg13g2_and2_1 _3788_ (.A(net1048),
    .B(net1004),
    .X(_0851_));
 sg13g2_nand3_1 _3789_ (.B(net1049),
    .C(net1004),
    .A(\vga_tetris.boardMem.board_7[16] ),
    .Y(_0852_));
 sg13g2_and2_1 _3790_ (.A(net1035),
    .B(net1004),
    .X(_0853_));
 sg13g2_and2_1 _3791_ (.A(net1043),
    .B(net1036),
    .X(_0854_));
 sg13g2_nand3_1 _3792_ (.B(net1042),
    .C(net1035),
    .A(\vga_tetris.boardMem.board_1[16] ),
    .Y(_0855_));
 sg13g2_and2_1 _3793_ (.A(net1028),
    .B(net1009),
    .X(_0856_));
 sg13g2_and2_1 _3794_ (.A(net1035),
    .B(net1024),
    .X(_0857_));
 sg13g2_a22oi_1 _3795_ (.Y(_0858_),
    .B1(net983),
    .B2(\vga_tetris.boardMem.board_16[16] ),
    .A2(net985),
    .A1(\vga_tetris.boardMem.board_19[16] ));
 sg13g2_a22oi_1 _3796_ (.Y(_0859_),
    .B1(net969),
    .B2(\vga_tetris.boardMem.board_17[16] ),
    .A2(net978),
    .A1(\vga_tetris.boardMem.board_2[16] ));
 sg13g2_a22oi_1 _3797_ (.Y(_0860_),
    .B1(net974),
    .B2(\vga_tetris.boardMem.board_5[16] ),
    .A2(net1003),
    .A1(\vga_tetris.boardMem.board_11[16] ));
 sg13g2_a22oi_1 _3798_ (.Y(_0861_),
    .B1(net981),
    .B2(\vga_tetris.boardMem.board_6[16] ),
    .A2(net997),
    .A1(\vga_tetris.boardMem.board_9[16] ));
 sg13g2_a221oi_1 _3799_ (.B2(\vga_tetris.boardMem.board_14[16] ),
    .C1(_0847_),
    .B1(net971),
    .A1(\vga_tetris.boardMem.board_10[16] ),
    .Y(_0862_),
    .A2(net987));
 sg13g2_and4_1 _3800_ (.A(_0826_),
    .B(_0835_),
    .C(_0838_),
    .D(_0849_),
    .X(_0863_));
 sg13g2_nand4_1 _3801_ (.B(_0859_),
    .C(_0862_),
    .A(_0858_),
    .Y(_0864_),
    .D(_0863_));
 sg13g2_and4_1 _3802_ (.A(_0822_),
    .B(_0840_),
    .C(_0852_),
    .D(_0855_),
    .X(_0865_));
 sg13g2_nand4_1 _3803_ (.B(_0860_),
    .C(_0861_),
    .A(net964),
    .Y(_0866_),
    .D(_0865_));
 sg13g2_nand2_1 _3804_ (.Y(_0867_),
    .A(_0626_),
    .B(\vga_tetris._vgaController_io_pixelPosX[8] ));
 sg13g2_a21o_1 _3805_ (.A2(net1191),
    .A1(net1190),
    .B1(_0867_),
    .X(_0868_));
 sg13g2_a21o_1 _3806_ (.A2(net1193),
    .A1(net1190),
    .B1(_0868_),
    .X(_0869_));
 sg13g2_nor4_1 _3807_ (.A(\vga_tetris._vgaController_io_pixelPosY[9] ),
    .B(_0775_),
    .C(_0777_),
    .D(_0869_),
    .Y(_0870_));
 sg13g2_or4_1 _3808_ (.A(net1187),
    .B(net1188),
    .C(\vga_tetris._vgaController_io_pixelPosY[1] ),
    .D(\vga_tetris._vgaController_io_pixelPosY[0] ),
    .X(_0871_));
 sg13g2_nand2_2 _3809_ (.Y(_0872_),
    .A(net1599),
    .B(net1723));
 sg13g2_nand2_2 _3810_ (.Y(_0873_),
    .A(net1782),
    .B(net1198));
 sg13g2_nor2_1 _3811_ (.A(_0628_),
    .B(_0872_),
    .Y(_0874_));
 sg13g2_nor2_2 _3812_ (.A(_0872_),
    .B(_0873_),
    .Y(_0875_));
 sg13g2_nand2_2 _3813_ (.Y(_0876_),
    .A(net1782),
    .B(_0874_));
 sg13g2_nand3_1 _3814_ (.B(net1779),
    .C(net1610),
    .A(net1188),
    .Y(_0877_));
 sg13g2_nand4_1 _3815_ (.B(net1188),
    .C(net1779),
    .A(net1187),
    .Y(_0878_),
    .D(net1892));
 sg13g2_inv_1 _3816_ (.Y(_0879_),
    .A(_0878_));
 sg13g2_nand4_1 _3817_ (.B(_0871_),
    .C(_0876_),
    .A(_0870_),
    .Y(_0880_),
    .D(_0878_));
 sg13g2_inv_1 _3818_ (.Y(_0881_),
    .A(_0880_));
 sg13g2_nor2_1 _3819_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[0] ),
    .B(_0701_),
    .Y(_0882_));
 sg13g2_nor2b_1 _3820_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[1] ),
    .B_N(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[0] ),
    .Y(_0883_));
 sg13g2_nor2b_2 _3821_ (.A(net1611),
    .B_N(_0883_),
    .Y(_0884_));
 sg13g2_inv_1 _3822_ (.Y(_0885_),
    .A(_0884_));
 sg13g2_o21ai_1 _3823_ (.B1(net1149),
    .Y(_0886_),
    .A1(_0882_),
    .A2(_0884_));
 sg13g2_nand2_1 _3824_ (.Y(_0887_),
    .A(\vga_tetris.tetrisLogic.addOrRemoveShape.stateQ[0] ),
    .B(_0664_));
 sg13g2_o21ai_1 _3825_ (.B1(_0886_),
    .Y(_0888_),
    .A1(net1149),
    .A2(net1164));
 sg13g2_nor2_1 _3826_ (.A(net1175),
    .B(_0888_),
    .Y(_0889_));
 sg13g2_nand2_1 _3827_ (.Y(_0890_),
    .A(_0731_),
    .B(_0889_));
 sg13g2_a22oi_1 _3828_ (.Y(_0891_),
    .B1(_0889_),
    .B2(_0731_),
    .A2(_0880_),
    .A1(net1175));
 sg13g2_o21ai_1 _3829_ (.B1(_0890_),
    .Y(_0892_),
    .A1(net1178),
    .A2(_0881_));
 sg13g2_nand3b_1 _3830_ (.B(net995),
    .C(net993),
    .Y(_0893_),
    .A_N(\vga_tetris.boardMem.board_0[16] ));
 sg13g2_and2_1 _3831_ (.A(net1068),
    .B(_0893_),
    .X(_0894_));
 sg13g2_o21ai_1 _3832_ (.B1(_0893_),
    .Y(_0895_),
    .A1(_0864_),
    .A2(_0866_));
 sg13g2_nor2_1 _3833_ (.A(net1065),
    .B(_0895_),
    .Y(_0896_));
 sg13g2_o21ai_1 _3834_ (.B1(_0894_),
    .Y(_0897_),
    .A1(_0864_),
    .A2(_0866_));
 sg13g2_nor2b_2 _3835_ (.A(net1191),
    .B_N(net1190),
    .Y(_0898_));
 sg13g2_nor2_1 _3836_ (.A(net1193),
    .B(net1197),
    .Y(_0899_));
 sg13g2_nand2_1 _3837_ (.Y(_0900_),
    .A(_0898_),
    .B(_0899_));
 sg13g2_nor2_2 _3838_ (.A(net1190),
    .B(net1191),
    .Y(_0901_));
 sg13g2_and2_1 _3839_ (.A(_0899_),
    .B(_0901_),
    .X(_0902_));
 sg13g2_nand2_1 _3840_ (.Y(_0903_),
    .A(_0899_),
    .B(_0901_));
 sg13g2_nand3_1 _3841_ (.B(net1031),
    .C(net1012),
    .A(\vga_tetris.boardMem.board_14[0] ),
    .Y(_0904_));
 sg13g2_nand3_1 _3842_ (.B(net1037),
    .C(net1005),
    .A(\vga_tetris.boardMem.board_5[0] ),
    .Y(_0905_));
 sg13g2_nand3_1 _3843_ (.B(net1047),
    .C(net1023),
    .A(\vga_tetris.boardMem.board_19[0] ),
    .Y(_0906_));
 sg13g2_nand3_1 _3844_ (.B(net1047),
    .C(net1041),
    .A(\vga_tetris.boardMem.board_3[0] ),
    .Y(_0907_));
 sg13g2_nand3_1 _3845_ (.B(net1037),
    .C(net1023),
    .A(\vga_tetris.boardMem.board_17[0] ),
    .Y(_0908_));
 sg13g2_nand3_1 _3846_ (.B(net1053),
    .C(net1047),
    .A(\vga_tetris.boardMem.board_11[0] ),
    .Y(_0909_));
 sg13g2_and3_1 _3847_ (.X(_0910_),
    .A(\vga_tetris.boardMem.board_10[0] ),
    .B(net1056),
    .C(net1015));
 sg13g2_nand3_1 _3848_ (.B(net1047),
    .C(net1028),
    .A(\vga_tetris.boardMem.board_15[0] ),
    .Y(_0911_));
 sg13g2_nand3_1 _3849_ (.B(net1043),
    .C(net1012),
    .A(\vga_tetris.boardMem.board_2[0] ),
    .Y(_0912_));
 sg13g2_nand2_1 _3850_ (.Y(_0913_),
    .A(\vga_tetris.boardMem.board_1[0] ),
    .B(net972));
 sg13g2_a221oi_1 _3851_ (.B2(\vga_tetris.boardMem.board_4[0] ),
    .C1(_0910_),
    .B1(net980),
    .A1(\vga_tetris.boardMem.board_16[0] ),
    .Y(_0914_),
    .A2(net983));
 sg13g2_a22oi_1 _3852_ (.Y(_0915_),
    .B1(net991),
    .B2(\vga_tetris.boardMem.board_18[0] ),
    .A2(net999),
    .A1(\vga_tetris.boardMem.board_13[0] ));
 sg13g2_a22oi_1 _3853_ (.Y(_0916_),
    .B1(net977),
    .B2(\vga_tetris.boardMem.board_7[0] ),
    .A2(net981),
    .A1(\vga_tetris.boardMem.board_6[0] ));
 sg13g2_nand4_1 _3854_ (.B(_0914_),
    .C(_0915_),
    .A(_0913_),
    .Y(_0917_),
    .D(_0916_));
 sg13g2_and4_1 _3855_ (.A(_0904_),
    .B(_0907_),
    .C(_0908_),
    .D(_0909_),
    .X(_0918_));
 sg13g2_a22oi_1 _3856_ (.Y(_0919_),
    .B1(_0848_),
    .B2(\vga_tetris.boardMem.board_8[0] ),
    .A2(net997),
    .A1(\vga_tetris.boardMem.board_9[0] ));
 sg13g2_a22oi_1 _3857_ (.Y(_0920_),
    .B1(net992),
    .B2(\vga_tetris.boardMem.board_12[0] ),
    .A2(net993),
    .A1(net995));
 sg13g2_and4_1 _3858_ (.A(_0905_),
    .B(_0906_),
    .C(_0911_),
    .D(_0912_),
    .X(_0921_));
 sg13g2_nand4_1 _3859_ (.B(_0919_),
    .C(_0920_),
    .A(_0918_),
    .Y(_0922_),
    .D(_0921_));
 sg13g2_a21oi_1 _3860_ (.A1(_0663_),
    .A2(net967),
    .Y(_0923_),
    .B1(net1065));
 sg13g2_o21ai_1 _3861_ (.B1(_0923_),
    .Y(_0924_),
    .A1(_0917_),
    .A2(_0922_));
 sg13g2_nand3_1 _3862_ (.B(net1017),
    .C(net1005),
    .A(\vga_tetris.boardMem.board_4[10] ),
    .Y(_0925_));
 sg13g2_nand2_1 _3863_ (.Y(_0926_),
    .A(\vga_tetris.boardMem.board_7[10] ),
    .B(net977));
 sg13g2_nand3_1 _3864_ (.B(net1052),
    .C(net1037),
    .A(\vga_tetris.boardMem.board_9[10] ),
    .Y(_0927_));
 sg13g2_nand3_1 _3865_ (.B(net1041),
    .C(net1008),
    .A(\vga_tetris.boardMem.board_2[10] ),
    .Y(_0928_));
 sg13g2_nand3_1 _3866_ (.B(net1023),
    .C(net1008),
    .A(\vga_tetris.boardMem.board_18[10] ),
    .Y(_0929_));
 sg13g2_nand3_1 _3867_ (.B(net1028),
    .C(net1017),
    .A(\vga_tetris.boardMem.board_12[10] ),
    .Y(_0930_));
 sg13g2_nand3_1 _3868_ (.B(net1028),
    .C(net1009),
    .A(\vga_tetris.boardMem.board_14[10] ),
    .Y(_0931_));
 sg13g2_nand3_1 _3869_ (.B(net1052),
    .C(net1046),
    .A(\vga_tetris.boardMem.board_11[10] ),
    .Y(_0932_));
 sg13g2_nand3_1 _3870_ (.B(net1046),
    .C(net1041),
    .A(\vga_tetris.boardMem.board_3[10] ),
    .Y(_0933_));
 sg13g2_and3_1 _3871_ (.X(_0934_),
    .A(\vga_tetris.boardMem.board_6[10] ),
    .B(net1009),
    .C(net1005));
 sg13g2_a22oi_1 _3872_ (.Y(_0935_),
    .B1(net969),
    .B2(\vga_tetris.boardMem.board_17[10] ),
    .A2(net987),
    .A1(\vga_tetris.boardMem.board_10[10] ));
 sg13g2_a22oi_1 _3873_ (.Y(_0936_),
    .B1(_0848_),
    .B2(\vga_tetris.boardMem.board_8[10] ),
    .A2(net993),
    .A1(net995));
 sg13g2_a22oi_1 _3874_ (.Y(_0937_),
    .B1(net974),
    .B2(\vga_tetris.boardMem.board_5[10] ),
    .A2(net983),
    .A1(\vga_tetris.boardMem.board_16[10] ));
 sg13g2_a22oi_1 _3875_ (.Y(_0938_),
    .B1(net990),
    .B2(\vga_tetris.boardMem.board_15[10] ),
    .A2(net999),
    .A1(\vga_tetris.boardMem.board_13[10] ));
 sg13g2_nand4_1 _3876_ (.B(_0936_),
    .C(_0937_),
    .A(_0935_),
    .Y(_0939_),
    .D(_0938_));
 sg13g2_and4_1 _3877_ (.A(_0925_),
    .B(_0927_),
    .C(_0930_),
    .D(_0931_),
    .X(_0940_));
 sg13g2_a221oi_1 _3878_ (.B2(\vga_tetris.boardMem.board_1[10] ),
    .C1(_0934_),
    .B1(net972),
    .A1(\vga_tetris.boardMem.board_19[10] ),
    .Y(_0941_),
    .A2(net985));
 sg13g2_and4_1 _3879_ (.A(_0928_),
    .B(_0929_),
    .C(_0932_),
    .D(_0933_),
    .X(_0942_));
 sg13g2_nand4_1 _3880_ (.B(_0940_),
    .C(_0941_),
    .A(_0926_),
    .Y(_0943_),
    .D(_0942_));
 sg13g2_a21oi_1 _3881_ (.A1(_0668_),
    .A2(net967),
    .Y(_0944_),
    .B1(net1065));
 sg13g2_o21ai_1 _3882_ (.B1(_0944_),
    .Y(_0945_),
    .A1(_0939_),
    .A2(_0943_));
 sg13g2_nand2b_2 _3883_ (.Y(_0946_),
    .B(net1191),
    .A_N(net1190));
 sg13g2_nor2b_2 _3884_ (.A(net1193),
    .B_N(net1197),
    .Y(_0947_));
 sg13g2_nand2b_1 _3885_ (.Y(_0948_),
    .B(_0947_),
    .A_N(_0946_));
 sg13g2_or2_1 _3886_ (.X(_0949_),
    .B(_0948_),
    .A(_0945_));
 sg13g2_nand2_2 _3887_ (.Y(_0950_),
    .A(net1193),
    .B(net1196));
 sg13g2_or2_1 _3888_ (.X(_0951_),
    .B(_0950_),
    .A(_0946_));
 sg13g2_nand3_1 _3889_ (.B(net1052),
    .C(net1046),
    .A(\vga_tetris.boardMem.board_11[14] ),
    .Y(_0952_));
 sg13g2_and3_1 _3890_ (.X(_0953_),
    .A(\vga_tetris.boardMem.board_10[14] ),
    .B(net1052),
    .C(net1009));
 sg13g2_nand3_1 _3891_ (.B(net1023),
    .C(net1017),
    .A(\vga_tetris.boardMem.board_16[14] ),
    .Y(_0954_));
 sg13g2_nand2_1 _3892_ (.Y(_0955_),
    .A(\vga_tetris.boardMem.board_1[14] ),
    .B(net972));
 sg13g2_nand3_1 _3893_ (.B(net1052),
    .C(net1017),
    .A(\vga_tetris.boardMem.board_8[14] ),
    .Y(_0956_));
 sg13g2_nand3_1 _3894_ (.B(net1028),
    .C(net1008),
    .A(\vga_tetris.boardMem.board_14[14] ),
    .Y(_0957_));
 sg13g2_nand3_1 _3895_ (.B(net1046),
    .C(net1041),
    .A(\vga_tetris.boardMem.board_3[14] ),
    .Y(_0958_));
 sg13g2_nand3_1 _3896_ (.B(net1041),
    .C(net1008),
    .A(\vga_tetris.boardMem.board_2[14] ),
    .Y(_0959_));
 sg13g2_nand3_1 _3897_ (.B(net1052),
    .C(net1037),
    .A(\vga_tetris.boardMem.board_9[14] ),
    .Y(_0960_));
 sg13g2_nand3_1 _3898_ (.B(net1023),
    .C(net1008),
    .A(\vga_tetris.boardMem.board_18[14] ),
    .Y(_0961_));
 sg13g2_a22oi_1 _3899_ (.Y(_0962_),
    .B1(net969),
    .B2(\vga_tetris.boardMem.board_17[14] ),
    .A2(net977),
    .A1(\vga_tetris.boardMem.board_7[14] ));
 sg13g2_a22oi_1 _3900_ (.Y(_0963_),
    .B1(net992),
    .B2(\vga_tetris.boardMem.board_12[14] ),
    .A2(net993),
    .A1(net995));
 sg13g2_a22oi_1 _3901_ (.Y(_0964_),
    .B1(net985),
    .B2(\vga_tetris.boardMem.board_19[14] ),
    .A2(net990),
    .A1(\vga_tetris.boardMem.board_15[14] ));
 sg13g2_a22oi_1 _3902_ (.Y(_0965_),
    .B1(net974),
    .B2(\vga_tetris.boardMem.board_5[14] ),
    .A2(net999),
    .A1(\vga_tetris.boardMem.board_13[14] ));
 sg13g2_nand4_1 _3903_ (.B(_0963_),
    .C(_0964_),
    .A(_0962_),
    .Y(_0966_),
    .D(_0965_));
 sg13g2_and4_1 _3904_ (.A(_0956_),
    .B(_0957_),
    .C(_0958_),
    .D(_0959_),
    .X(_0967_));
 sg13g2_a221oi_1 _3905_ (.B2(\vga_tetris.boardMem.board_4[14] ),
    .C1(_0953_),
    .B1(net980),
    .A1(\vga_tetris.boardMem.board_6[14] ),
    .Y(_0968_),
    .A2(net981));
 sg13g2_and4_1 _3906_ (.A(_0952_),
    .B(_0954_),
    .C(_0960_),
    .D(_0961_),
    .X(_0969_));
 sg13g2_nand4_1 _3907_ (.B(_0967_),
    .C(_0968_),
    .A(_0955_),
    .Y(_0970_),
    .D(_0969_));
 sg13g2_a21oi_1 _3908_ (.A1(_0672_),
    .A2(net967),
    .Y(_0971_),
    .B1(net1065));
 sg13g2_o21ai_1 _3909_ (.B1(_0971_),
    .Y(_0972_),
    .A1(_0966_),
    .A2(_0970_));
 sg13g2_nor2_1 _3910_ (.A(_0951_),
    .B(_0972_),
    .Y(_0973_));
 sg13g2_nand2_1 _3911_ (.Y(_0974_),
    .A(\vga_tetris.boardMem.board_18[18] ),
    .B(net991));
 sg13g2_a22oi_1 _3912_ (.Y(_0975_),
    .B1(net974),
    .B2(\vga_tetris.boardMem.board_5[18] ),
    .A2(net987),
    .A1(\vga_tetris.boardMem.board_10[18] ));
 sg13g2_a22oi_1 _3913_ (.Y(_0976_),
    .B1(net970),
    .B2(\vga_tetris.boardMem.board_17[18] ),
    .A2(net1001),
    .A1(\vga_tetris.boardMem.board_3[18] ));
 sg13g2_a22oi_1 _3914_ (.Y(_0977_),
    .B1(net972),
    .B2(\vga_tetris.boardMem.board_1[18] ),
    .A2(net999),
    .A1(\vga_tetris.boardMem.board_13[18] ));
 sg13g2_a22oi_1 _3915_ (.Y(_0978_),
    .B1(_0848_),
    .B2(\vga_tetris.boardMem.board_8[18] ),
    .A2(net989),
    .A1(\vga_tetris.boardMem.board_15[18] ));
 sg13g2_nand4_1 _3916_ (.B(_0976_),
    .C(_0977_),
    .A(_0975_),
    .Y(_0979_),
    .D(_0978_));
 sg13g2_a22oi_1 _3917_ (.Y(_0980_),
    .B1(net981),
    .B2(\vga_tetris.boardMem.board_6[18] ),
    .A2(net985),
    .A1(\vga_tetris.boardMem.board_19[18] ));
 sg13g2_a22oi_1 _3918_ (.Y(_0981_),
    .B1(net978),
    .B2(\vga_tetris.boardMem.board_2[18] ),
    .A2(net1002),
    .A1(\vga_tetris.boardMem.board_11[18] ));
 sg13g2_a22oi_1 _3919_ (.Y(_0982_),
    .B1(net976),
    .B2(\vga_tetris.boardMem.board_7[18] ),
    .A2(net984),
    .A1(\vga_tetris.boardMem.board_16[18] ));
 sg13g2_a22oi_1 _3920_ (.Y(_0983_),
    .B1(net971),
    .B2(\vga_tetris.boardMem.board_14[18] ),
    .A2(net979),
    .A1(\vga_tetris.boardMem.board_4[18] ));
 sg13g2_nand4_1 _3921_ (.B(_0981_),
    .C(_0982_),
    .A(_0980_),
    .Y(_0984_),
    .D(_0983_));
 sg13g2_a22oi_1 _3922_ (.Y(_0985_),
    .B1(net992),
    .B2(\vga_tetris.boardMem.board_12[18] ),
    .A2(net997),
    .A1(\vga_tetris.boardMem.board_9[18] ));
 sg13g2_nand3_1 _3923_ (.B(_0974_),
    .C(_0985_),
    .A(net965),
    .Y(_0986_));
 sg13g2_nor3_2 _3924_ (.A(_0979_),
    .B(_0984_),
    .C(_0986_),
    .Y(_0987_));
 sg13g2_o21ai_1 _3925_ (.B1(net1068),
    .Y(_0988_),
    .A1(\vga_tetris.boardMem.board_0[18] ),
    .A2(net965));
 sg13g2_nor2_2 _3926_ (.A(_0987_),
    .B(_0988_),
    .Y(_0989_));
 sg13g2_nand2_1 _3927_ (.Y(_0990_),
    .A(_0898_),
    .B(_0947_));
 sg13g2_nand3_1 _3928_ (.B(_0947_),
    .C(_0989_),
    .A(_0898_),
    .Y(_0991_));
 sg13g2_a22oi_1 _3929_ (.Y(_0992_),
    .B1(_0848_),
    .B2(\vga_tetris.boardMem.board_8[4] ),
    .A2(net1002),
    .A1(\vga_tetris.boardMem.board_11[4] ));
 sg13g2_nand2_1 _3930_ (.Y(_0993_),
    .A(\vga_tetris.boardMem.board_18[4] ),
    .B(net991));
 sg13g2_a22oi_1 _3931_ (.Y(_0994_),
    .B1(net976),
    .B2(\vga_tetris.boardMem.board_7[4] ),
    .A2(net1001),
    .A1(\vga_tetris.boardMem.board_3[4] ));
 sg13g2_a22oi_1 _3932_ (.Y(_0995_),
    .B1(net978),
    .B2(\vga_tetris.boardMem.board_2[4] ),
    .A2(net1000),
    .A1(\vga_tetris.boardMem.board_13[4] ));
 sg13g2_a22oi_1 _3933_ (.Y(_0996_),
    .B1(net985),
    .B2(\vga_tetris.boardMem.board_19[4] ),
    .A2(net989),
    .A1(\vga_tetris.boardMem.board_15[4] ));
 sg13g2_a22oi_1 _3934_ (.Y(_0997_),
    .B1(net970),
    .B2(\vga_tetris.boardMem.board_17[4] ),
    .A2(net981),
    .A1(\vga_tetris.boardMem.board_6[4] ));
 sg13g2_nand4_1 _3935_ (.B(_0995_),
    .C(_0996_),
    .A(_0994_),
    .Y(_0998_),
    .D(_0997_));
 sg13g2_a22oi_1 _3936_ (.Y(_0999_),
    .B1(net979),
    .B2(\vga_tetris.boardMem.board_4[4] ),
    .A2(net987),
    .A1(\vga_tetris.boardMem.board_10[4] ));
 sg13g2_a22oi_1 _3937_ (.Y(_1000_),
    .B1(net973),
    .B2(\vga_tetris.boardMem.board_1[4] ),
    .A2(net997),
    .A1(\vga_tetris.boardMem.board_9[4] ));
 sg13g2_a22oi_1 _3938_ (.Y(_1001_),
    .B1(net975),
    .B2(\vga_tetris.boardMem.board_5[4] ),
    .A2(net983),
    .A1(\vga_tetris.boardMem.board_16[4] ));
 sg13g2_a22oi_1 _3939_ (.Y(_1002_),
    .B1(net971),
    .B2(\vga_tetris.boardMem.board_14[4] ),
    .A2(net992),
    .A1(\vga_tetris.boardMem.board_12[4] ));
 sg13g2_nand2_1 _3940_ (.Y(_1003_),
    .A(_0993_),
    .B(_1001_));
 sg13g2_nand4_1 _3941_ (.B(_0999_),
    .C(_1000_),
    .A(_0992_),
    .Y(_1004_),
    .D(_1002_));
 sg13g2_or4_1 _3942_ (.A(net968),
    .B(_0998_),
    .C(_1003_),
    .D(_1004_),
    .X(_1005_));
 sg13g2_a21oi_1 _3943_ (.A1(_0666_),
    .A2(net967),
    .Y(_1006_),
    .B1(net1065));
 sg13g2_nand2_2 _3944_ (.Y(_1007_),
    .A(_1005_),
    .B(_1006_));
 sg13g2_nor2b_2 _3945_ (.A(net1197),
    .B_N(net1193),
    .Y(_1008_));
 sg13g2_nand2_1 _3946_ (.Y(_1009_),
    .A(_0901_),
    .B(_1008_));
 sg13g2_o21ai_1 _3947_ (.B1(_0991_),
    .Y(_1010_),
    .A1(_1007_),
    .A2(_1009_));
 sg13g2_nand3_1 _3948_ (.B(net1050),
    .C(net1027),
    .A(\vga_tetris.boardMem.board_19[6] ),
    .Y(_1011_));
 sg13g2_nand3_1 _3949_ (.B(net1040),
    .C(net1034),
    .A(\vga_tetris.boardMem.board_13[6] ),
    .Y(_1012_));
 sg13g2_nand3_1 _3950_ (.B(net1014),
    .C(net1007),
    .A(\vga_tetris.boardMem.board_6[6] ),
    .Y(_1013_));
 sg13g2_nand3_1 _3951_ (.B(net1051),
    .C(net1045),
    .A(\vga_tetris.boardMem.board_3[6] ),
    .Y(_1014_));
 sg13g2_and3_1 _3952_ (.X(_1015_),
    .A(\vga_tetris.boardMem.board_18[6] ),
    .B(net1027),
    .C(net1014));
 sg13g2_nand3_1 _3953_ (.B(net1032),
    .C(net1015),
    .A(\vga_tetris.boardMem.board_14[6] ),
    .Y(_1016_));
 sg13g2_nand3_1 _3954_ (.B(net1044),
    .C(net1040),
    .A(\vga_tetris.boardMem.board_1[6] ),
    .Y(_1017_));
 sg13g2_nand3_1 _3955_ (.B(net1058),
    .C(net1021),
    .A(\vga_tetris.boardMem.board_8[6] ),
    .Y(_1018_));
 sg13g2_nand3_1 _3956_ (.B(net1034),
    .C(net1021),
    .A(\vga_tetris.boardMem.board_12[6] ),
    .Y(_1019_));
 sg13g2_a22oi_1 _3957_ (.Y(_1020_),
    .B1(net970),
    .B2(\vga_tetris.boardMem.board_17[6] ),
    .A2(net990),
    .A1(\vga_tetris.boardMem.board_15[6] ));
 sg13g2_a22oi_1 _3958_ (.Y(_1021_),
    .B1(net976),
    .B2(\vga_tetris.boardMem.board_7[6] ),
    .A2(net978),
    .A1(\vga_tetris.boardMem.board_2[6] ));
 sg13g2_a22oi_1 _3959_ (.Y(_1022_),
    .B1(net974),
    .B2(\vga_tetris.boardMem.board_5[6] ),
    .A2(net997),
    .A1(\vga_tetris.boardMem.board_9[6] ));
 sg13g2_a22oi_1 _3960_ (.Y(_1023_),
    .B1(net980),
    .B2(\vga_tetris.boardMem.board_4[6] ),
    .A2(net987),
    .A1(\vga_tetris.boardMem.board_10[6] ));
 sg13g2_a221oi_1 _3961_ (.B2(\vga_tetris.boardMem.board_16[6] ),
    .C1(_1015_),
    .B1(net984),
    .A1(\vga_tetris.boardMem.board_11[6] ),
    .Y(_1024_),
    .A2(net1002));
 sg13g2_and4_1 _3962_ (.A(_1012_),
    .B(_1013_),
    .C(_1014_),
    .D(_1018_),
    .X(_1025_));
 sg13g2_and4_1 _3963_ (.A(_1020_),
    .B(_1021_),
    .C(_1024_),
    .D(_1025_),
    .X(_1026_));
 sg13g2_and4_1 _3964_ (.A(_1011_),
    .B(_1016_),
    .C(_1017_),
    .D(_1019_),
    .X(_1027_));
 sg13g2_and4_1 _3965_ (.A(net964),
    .B(_1022_),
    .C(_1023_),
    .D(_1027_),
    .X(_1028_));
 sg13g2_o21ai_1 _3966_ (.B1(net1068),
    .Y(_1029_),
    .A1(net1467),
    .A2(net964));
 sg13g2_a21oi_2 _3967_ (.B1(_1029_),
    .Y(_1030_),
    .A2(_1028_),
    .A1(_1026_));
 sg13g2_a21o_1 _3968_ (.A2(_1028_),
    .A1(_1026_),
    .B1(_1029_),
    .X(_1031_));
 sg13g2_nor3_1 _3969_ (.A(net1190),
    .B(net1191),
    .C(_0950_),
    .Y(_1032_));
 sg13g2_nand2_1 _3970_ (.Y(_1033_),
    .A(_1030_),
    .B(_1032_));
 sg13g2_a22oi_1 _3971_ (.Y(_1034_),
    .B1(net970),
    .B2(\vga_tetris.boardMem.board_17[2] ),
    .A2(_0848_),
    .A1(\vga_tetris.boardMem.board_8[2] ));
 sg13g2_nand2_1 _3972_ (.Y(_1035_),
    .A(\vga_tetris.boardMem.board_5[2] ),
    .B(net975));
 sg13g2_a22oi_1 _3973_ (.Y(_1036_),
    .B1(net991),
    .B2(\vga_tetris.boardMem.board_18[2] ),
    .A2(net1001),
    .A1(\vga_tetris.boardMem.board_3[2] ));
 sg13g2_a22oi_1 _3974_ (.Y(_1037_),
    .B1(net971),
    .B2(\vga_tetris.boardMem.board_14[2] ),
    .A2(net984),
    .A1(\vga_tetris.boardMem.board_16[2] ));
 sg13g2_a22oi_1 _3975_ (.Y(_1038_),
    .B1(net982),
    .B2(\vga_tetris.boardMem.board_6[2] ),
    .A2(net992),
    .A1(\vga_tetris.boardMem.board_12[2] ));
 sg13g2_a22oi_1 _3976_ (.Y(_1039_),
    .B1(net976),
    .B2(\vga_tetris.boardMem.board_7[2] ),
    .A2(net997),
    .A1(\vga_tetris.boardMem.board_9[2] ));
 sg13g2_a22oi_1 _3977_ (.Y(_1040_),
    .B1(net988),
    .B2(\vga_tetris.boardMem.board_10[2] ),
    .A2(net989),
    .A1(\vga_tetris.boardMem.board_15[2] ));
 sg13g2_a22oi_1 _3978_ (.Y(_1041_),
    .B1(net1000),
    .B2(\vga_tetris.boardMem.board_13[2] ),
    .A2(net1002),
    .A1(\vga_tetris.boardMem.board_11[2] ));
 sg13g2_nand2_1 _3979_ (.Y(_1042_),
    .A(_1035_),
    .B(_1039_));
 sg13g2_a22oi_1 _3980_ (.Y(_1043_),
    .B1(net973),
    .B2(\vga_tetris.boardMem.board_1[2] ),
    .A2(net979),
    .A1(\vga_tetris.boardMem.board_4[2] ));
 sg13g2_nand4_1 _3981_ (.B(_1040_),
    .C(_1041_),
    .A(_1034_),
    .Y(_1044_),
    .D(_1043_));
 sg13g2_a22oi_1 _3982_ (.Y(_1045_),
    .B1(net978),
    .B2(\vga_tetris.boardMem.board_2[2] ),
    .A2(net985),
    .A1(\vga_tetris.boardMem.board_19[2] ));
 sg13g2_nand4_1 _3983_ (.B(_1037_),
    .C(_1038_),
    .A(_1036_),
    .Y(_1046_),
    .D(_1045_));
 sg13g2_or4_1 _3984_ (.A(net968),
    .B(_1042_),
    .C(_1044_),
    .D(_1046_),
    .X(_1047_));
 sg13g2_a21oi_2 _3985_ (.B1(net1066),
    .Y(_1048_),
    .A2(net968),
    .A1(_0665_));
 sg13g2_nand2_1 _3986_ (.Y(_1049_),
    .A(_1047_),
    .B(_1048_));
 sg13g2_and4_1 _3987_ (.A(_0901_),
    .B(_0947_),
    .C(_1047_),
    .D(_1048_),
    .X(_1050_));
 sg13g2_nand3_1 _3988_ (.B(net1038),
    .C(net1026),
    .A(\vga_tetris.boardMem.board_17[12] ),
    .Y(_1051_));
 sg13g2_nand3_1 _3989_ (.B(net1032),
    .C(net1013),
    .A(\vga_tetris.boardMem.board_14[12] ),
    .Y(_1052_));
 sg13g2_nand3_1 _3990_ (.B(net1038),
    .C(net1006),
    .A(\vga_tetris.boardMem.board_5[12] ),
    .Y(_1053_));
 sg13g2_nand3_1 _3991_ (.B(net1056),
    .C(net1038),
    .A(\vga_tetris.boardMem.board_9[12] ),
    .Y(_1054_));
 sg13g2_nand3_1 _3992_ (.B(net1057),
    .C(net1013),
    .A(\vga_tetris.boardMem.board_10[12] ),
    .Y(_1055_));
 sg13g2_nand3_1 _3993_ (.B(net1033),
    .C(net1020),
    .A(\vga_tetris.boardMem.board_12[12] ),
    .Y(_1056_));
 sg13g2_and3_1 _3994_ (.X(_1057_),
    .A(\vga_tetris.boardMem.board_2[12] ),
    .B(net1044),
    .C(net1013));
 sg13g2_nand3_1 _3995_ (.B(net1050),
    .C(net1033),
    .A(\vga_tetris.boardMem.board_15[12] ),
    .Y(_1058_));
 sg13g2_nand3_1 _3996_ (.B(net1057),
    .C(net1021),
    .A(\vga_tetris.boardMem.board_8[12] ),
    .Y(_1059_));
 sg13g2_and4_1 _3997_ (.A(_1054_),
    .B(_1055_),
    .C(_1056_),
    .D(_1058_),
    .X(_1060_));
 sg13g2_a22oi_1 _3998_ (.Y(_1061_),
    .B1(_0851_),
    .B2(\vga_tetris.boardMem.board_7[12] ),
    .A2(net1001),
    .A1(\vga_tetris.boardMem.board_3[12] ));
 sg13g2_a22oi_1 _3999_ (.Y(_1062_),
    .B1(net973),
    .B2(\vga_tetris.boardMem.board_1[12] ),
    .A2(net991),
    .A1(\vga_tetris.boardMem.board_18[12] ));
 sg13g2_a22oi_1 _4000_ (.Y(_1063_),
    .B1(net982),
    .B2(\vga_tetris.boardMem.board_6[12] ),
    .A2(net1003),
    .A1(\vga_tetris.boardMem.board_11[12] ));
 sg13g2_a22oi_1 _4001_ (.Y(_1064_),
    .B1(net979),
    .B2(\vga_tetris.boardMem.board_4[12] ),
    .A2(net1000),
    .A1(\vga_tetris.boardMem.board_13[12] ));
 sg13g2_and4_1 _4002_ (.A(_1051_),
    .B(_1052_),
    .C(_1053_),
    .D(_1059_),
    .X(_1065_));
 sg13g2_a221oi_1 _4003_ (.B2(\vga_tetris.boardMem.board_16[12] ),
    .C1(_1057_),
    .B1(net984),
    .A1(\vga_tetris.boardMem.board_19[12] ),
    .Y(_1066_),
    .A2(net986));
 sg13g2_nand4_1 _4004_ (.B(_1064_),
    .C(_1065_),
    .A(_1063_),
    .Y(_1067_),
    .D(_1066_));
 sg13g2_nand4_1 _4005_ (.B(_1060_),
    .C(_1061_),
    .A(net965),
    .Y(_1068_),
    .D(_1062_));
 sg13g2_a21oi_1 _4006_ (.A1(_0670_),
    .A2(net968),
    .Y(_1069_),
    .B1(net1066));
 sg13g2_o21ai_1 _4007_ (.B1(_1069_),
    .Y(_1070_),
    .A1(_1067_),
    .A2(_1068_));
 sg13g2_nand2b_1 _4008_ (.Y(_1071_),
    .B(_1008_),
    .A_N(_0946_));
 sg13g2_a22oi_1 _4009_ (.Y(_1072_),
    .B1(net971),
    .B2(\vga_tetris.boardMem.board_14[8] ),
    .A2(net998),
    .A1(\vga_tetris.boardMem.board_9[8] ));
 sg13g2_a22oi_1 _4010_ (.Y(_1073_),
    .B1(net973),
    .B2(\vga_tetris.boardMem.board_1[8] ),
    .A2(net989),
    .A1(\vga_tetris.boardMem.board_15[8] ));
 sg13g2_a22oi_1 _4011_ (.Y(_1074_),
    .B1(net996),
    .B2(net994),
    .A2(net1002),
    .A1(\vga_tetris.boardMem.board_11[8] ));
 sg13g2_a22oi_1 _4012_ (.Y(_1075_),
    .B1(net984),
    .B2(\vga_tetris.boardMem.board_16[8] ),
    .A2(net986),
    .A1(\vga_tetris.boardMem.board_19[8] ));
 sg13g2_and4_1 _4013_ (.A(_1072_),
    .B(_1073_),
    .C(_1074_),
    .D(_1075_),
    .X(_1076_));
 sg13g2_a22oi_1 _4014_ (.Y(_1077_),
    .B1(_0837_),
    .B2(\vga_tetris.boardMem.board_18[8] ),
    .A2(net1001),
    .A1(\vga_tetris.boardMem.board_3[8] ));
 sg13g2_a22oi_1 _4015_ (.Y(_1078_),
    .B1(net976),
    .B2(\vga_tetris.boardMem.board_7[8] ),
    .A2(_0846_),
    .A1(\vga_tetris.boardMem.board_4[8] ));
 sg13g2_nand3_1 _4016_ (.B(net1057),
    .C(net1013),
    .A(\vga_tetris.boardMem.board_10[8] ),
    .Y(_1079_));
 sg13g2_nand3_1 _4017_ (.B(net1038),
    .C(net1033),
    .A(\vga_tetris.boardMem.board_13[8] ),
    .Y(_1080_));
 sg13g2_nand3_1 _4018_ (.B(net1014),
    .C(net1006),
    .A(\vga_tetris.boardMem.board_6[8] ),
    .Y(_1081_));
 sg13g2_nand3_1 _4019_ (.B(net1057),
    .C(net1021),
    .A(\vga_tetris.boardMem.board_8[8] ),
    .Y(_1082_));
 sg13g2_and4_1 _4020_ (.A(_1079_),
    .B(_1080_),
    .C(_1081_),
    .D(_1082_),
    .X(_1083_));
 sg13g2_nand3_1 _4021_ (.B(net1044),
    .C(net1013),
    .A(\vga_tetris.boardMem.board_2[8] ),
    .Y(_1084_));
 sg13g2_nand3_1 _4022_ (.B(net1038),
    .C(net1026),
    .A(\vga_tetris.boardMem.board_17[8] ),
    .Y(_1085_));
 sg13g2_nand3_1 _4023_ (.B(net1038),
    .C(net1006),
    .A(\vga_tetris.boardMem.board_5[8] ),
    .Y(_1086_));
 sg13g2_nand3_1 _4024_ (.B(net1033),
    .C(net1021),
    .A(\vga_tetris.boardMem.board_12[8] ),
    .Y(_1087_));
 sg13g2_and4_1 _4025_ (.A(_1084_),
    .B(_1085_),
    .C(_1086_),
    .D(_1087_),
    .X(_1088_));
 sg13g2_and4_1 _4026_ (.A(_1077_),
    .B(_1078_),
    .C(_1083_),
    .D(_1088_),
    .X(_1089_));
 sg13g2_o21ai_1 _4027_ (.B1(net1068),
    .Y(_1090_),
    .A1(net1572),
    .A2(net965));
 sg13g2_a21o_2 _4028_ (.A2(_1089_),
    .A1(_1076_),
    .B1(_1090_),
    .X(_1091_));
 sg13g2_or4_1 _4029_ (.A(net1193),
    .B(net1197),
    .C(_0946_),
    .D(_1091_),
    .X(_1092_));
 sg13g2_o21ai_1 _4030_ (.B1(_0949_),
    .Y(_1093_),
    .A1(_1070_),
    .A2(_1071_));
 sg13g2_o21ai_1 _4031_ (.B1(_1033_),
    .Y(_1094_),
    .A1(_0897_),
    .A2(_0900_));
 sg13g2_o21ai_1 _4032_ (.B1(_1092_),
    .Y(_1095_),
    .A1(_0903_),
    .A2(_0924_));
 sg13g2_or4_1 _4033_ (.A(_0973_),
    .B(_1010_),
    .C(_1050_),
    .D(_1095_),
    .X(_1096_));
 sg13g2_nor3_1 _4034_ (.A(_1093_),
    .B(_1094_),
    .C(_1096_),
    .Y(_1097_));
 sg13g2_nand4_1 _4035_ (.B(net1809),
    .C(net1853),
    .A(net1602),
    .Y(_1098_),
    .D(\vga_tetris.vgaController.verticalCounterQ[5] ));
 sg13g2_inv_1 _4036_ (.Y(_1099_),
    .A(_1098_));
 sg13g2_nand2_1 _4037_ (.Y(_1100_),
    .A(\vga_tetris.vgaController.horizontalCounterQ[7] ),
    .B(\vga_tetris.vgaController.horizontalCounterQ[9] ));
 sg13g2_nand2_1 _4038_ (.Y(_1101_),
    .A(\vga_tetris.vgaController.horizontalCounterQ[8] ),
    .B(\vga_tetris.vgaController.horizontalCounterQ[9] ));
 sg13g2_nor2_1 _4039_ (.A(\vga_tetris.vgaController.verticalCounterQ[9] ),
    .B(net1223),
    .Y(_1102_));
 sg13g2_nand4_1 _4040_ (.B(_1100_),
    .C(_1101_),
    .A(_1098_),
    .Y(_1103_),
    .D(_1102_));
 sg13g2_or2_1 _4041_ (.X(_1104_),
    .B(_1103_),
    .A(_0880_));
 sg13g2_nor2_1 _4042_ (.A(_1097_),
    .B(_1104_),
    .Y(_1105_));
 sg13g2_nand2b_1 _4043_ (.Y(_1106_),
    .B(net1188),
    .A_N(net1183));
 sg13g2_xnor2_1 _4044_ (.Y(_1107_),
    .A(net1183),
    .B(net1188));
 sg13g2_nor2b_1 _4045_ (.A(\vga_tetris._vgaController_io_pixelPosY[1] ),
    .B_N(net1187),
    .Y(_1108_));
 sg13g2_nand2b_1 _4046_ (.Y(_1109_),
    .B(\vga_tetris._vgaController_io_pixelPosY[1] ),
    .A_N(net1187));
 sg13g2_nor2b_1 _4047_ (.A(\vga_tetris._vgaController_io_pixelPosY[0] ),
    .B_N(net1188),
    .Y(_1110_));
 sg13g2_a21oi_1 _4048_ (.A1(_1109_),
    .A2(_1110_),
    .Y(_1111_),
    .B1(_1108_));
 sg13g2_nand2_1 _4049_ (.Y(_1112_),
    .A(_1107_),
    .B(_1111_));
 sg13g2_nand2_1 _4050_ (.Y(_1113_),
    .A(_1106_),
    .B(_1112_));
 sg13g2_xor2_1 _4051_ (.B(_1113_),
    .A(net1185),
    .X(_1114_));
 sg13g2_xnor2_1 _4052_ (.Y(_1115_),
    .A(_1107_),
    .B(_1111_));
 sg13g2_nor2b_1 _4053_ (.A(net1182),
    .B_N(_1115_),
    .Y(_1116_));
 sg13g2_nor2b_1 _4054_ (.A(_1114_),
    .B_N(_1116_),
    .Y(_1117_));
 sg13g2_nand2_1 _4055_ (.Y(_1118_),
    .A(_1114_),
    .B(_1115_));
 sg13g2_inv_1 _4056_ (.Y(_1119_),
    .A(_1118_));
 sg13g2_nor2_2 _4057_ (.A(_1114_),
    .B(_1115_),
    .Y(_1120_));
 sg13g2_nand3b_1 _4058_ (.B(net1184),
    .C(_1118_),
    .Y(_1121_),
    .A_N(_1120_));
 sg13g2_nor2_1 _4059_ (.A(\vga_tetris._vgaController_io_pixelPosX[3] ),
    .B(\vga_tetris._vgaController_io_pixelPosX[2] ),
    .Y(_1122_));
 sg13g2_nand2_2 _4060_ (.Y(_1123_),
    .A(_0627_),
    .B(_0628_));
 sg13g2_a21oi_2 _4061_ (.B1(net1193),
    .Y(_1124_),
    .A2(_1123_),
    .A1(net1196));
 sg13g2_mux2_1 _4062_ (.A0(_0898_),
    .A1(_0901_),
    .S(_1124_),
    .X(_1125_));
 sg13g2_nand3_1 _4063_ (.B(net1180),
    .C(_0775_),
    .A(_0624_),
    .Y(_1126_));
 sg13g2_and2_1 _4064_ (.A(_0873_),
    .B(_1123_),
    .X(_1127_));
 sg13g2_nand2_1 _4065_ (.Y(_1128_),
    .A(_0873_),
    .B(_1123_));
 sg13g2_nor2_1 _4066_ (.A(net1195),
    .B(_1123_),
    .Y(_1129_));
 sg13g2_xnor2_1 _4067_ (.Y(_1130_),
    .A(net1195),
    .B(_1122_));
 sg13g2_nand2_1 _4068_ (.Y(_1131_),
    .A(_1128_),
    .B(_1130_));
 sg13g2_nor3_1 _4069_ (.A(_0868_),
    .B(_1125_),
    .C(_1126_),
    .Y(_1132_));
 sg13g2_nand3_1 _4070_ (.B(_1131_),
    .C(_1132_),
    .A(_1121_),
    .Y(_1133_));
 sg13g2_nor2_1 _4071_ (.A(_0950_),
    .B(_1122_),
    .Y(_1134_));
 sg13g2_nor2_2 _4072_ (.A(_1124_),
    .B(_1134_),
    .Y(_1135_));
 sg13g2_xnor2_1 _4073_ (.Y(_1136_),
    .A(net1192),
    .B(_1124_));
 sg13g2_nor2_1 _4074_ (.A(_1135_),
    .B(_1136_),
    .Y(_1137_));
 sg13g2_and2_1 _4075_ (.A(net1192),
    .B(_1135_),
    .X(_1138_));
 sg13g2_nand2b_1 _4076_ (.Y(_1139_),
    .B(_1138_),
    .A_N(\vga_tetris._tetrisLogic_io_score_1[2] ));
 sg13g2_a21o_1 _4077_ (.A2(_1136_),
    .A1(\vga_tetris._tetrisLogic_io_score_2[2] ),
    .B1(_1135_),
    .X(_1140_));
 sg13g2_nand2b_2 _4078_ (.Y(_1141_),
    .B(_1135_),
    .A_N(net1192));
 sg13g2_a22oi_1 _4079_ (.Y(_1142_),
    .B1(_1139_),
    .B2(_1140_),
    .A2(_1137_),
    .A1(\vga_tetris._tetrisLogic_io_score_0[2] ));
 sg13g2_nor2_1 _4080_ (.A(\vga_tetris._tetrisLogic_io_score_3[2] ),
    .B(_1141_),
    .Y(_1143_));
 sg13g2_nor3_2 _4081_ (.A(_1133_),
    .B(_1142_),
    .C(_1143_),
    .Y(_1144_));
 sg13g2_inv_2 _4082_ (.Y(_1145_),
    .A(_1144_));
 sg13g2_nor2_1 _4083_ (.A(\vga_tetris._tetrisLogic_io_score_3[1] ),
    .B(_1141_),
    .Y(_1146_));
 sg13g2_nand2_1 _4084_ (.Y(_1147_),
    .A(\vga_tetris._tetrisLogic_io_score_0[1] ),
    .B(_1137_));
 sg13g2_or2_1 _4085_ (.X(_1148_),
    .B(_1135_),
    .A(\vga_tetris._tetrisLogic_io_score_2[1] ));
 sg13g2_a22oi_1 _4086_ (.Y(_1149_),
    .B1(_1148_),
    .B2(_1136_),
    .A2(_1138_),
    .A1(\vga_tetris._tetrisLogic_io_score_1[1] ));
 sg13g2_a21oi_2 _4087_ (.B1(_1146_),
    .Y(_1150_),
    .A2(_1149_),
    .A1(_1147_));
 sg13g2_inv_1 _4088_ (.Y(_1151_),
    .A(_1150_));
 sg13g2_nand2b_1 _4089_ (.Y(_1152_),
    .B(_1150_),
    .A_N(_1133_));
 sg13g2_nor2b_1 _4090_ (.A(_1144_),
    .B_N(_1152_),
    .Y(_1153_));
 sg13g2_nand2_1 _4091_ (.Y(_1154_),
    .A(\vga_tetris._tetrisLogic_io_score_0[3] ),
    .B(_1137_));
 sg13g2_o21ai_1 _4092_ (.B1(_0689_),
    .Y(_1155_),
    .A1(_1124_),
    .A2(_1134_));
 sg13g2_a22oi_1 _4093_ (.Y(_1156_),
    .B1(_1155_),
    .B2(_1136_),
    .A2(_1138_),
    .A1(\vga_tetris._tetrisLogic_io_score_1[3] ));
 sg13g2_a21oi_1 _4094_ (.A1(_1154_),
    .A2(_1156_),
    .Y(_1157_),
    .B1(_1133_));
 sg13g2_o21ai_1 _4095_ (.B1(_1157_),
    .Y(_1158_),
    .A1(\vga_tetris._tetrisLogic_io_score_3[3] ),
    .A2(_1141_));
 sg13g2_o21ai_1 _4096_ (.B1(_1136_),
    .Y(_1159_),
    .A1(\vga_tetris._tetrisLogic_io_score_2[0] ),
    .A2(_1135_));
 sg13g2_a22oi_1 _4097_ (.Y(_1160_),
    .B1(_1138_),
    .B2(\vga_tetris._tetrisLogic_io_score_1[0] ),
    .A2(_1137_),
    .A1(\vga_tetris._tetrisLogic_io_score_0[0] ));
 sg13g2_nor2_1 _4098_ (.A(\vga_tetris._tetrisLogic_io_score_3[0] ),
    .B(_1141_),
    .Y(_1161_));
 sg13g2_a21oi_1 _4099_ (.A1(_1159_),
    .A2(_1160_),
    .Y(_1162_),
    .B1(_1161_));
 sg13g2_nand2b_2 _4100_ (.Y(_1163_),
    .B(_1162_),
    .A_N(_1133_));
 sg13g2_nor2_1 _4101_ (.A(_1150_),
    .B(_1163_),
    .Y(_1164_));
 sg13g2_nor2_1 _4102_ (.A(_1144_),
    .B(_1164_),
    .Y(_1165_));
 sg13g2_nor2_1 _4103_ (.A(_1151_),
    .B(_1163_),
    .Y(_1166_));
 sg13g2_nor2_1 _4104_ (.A(_1145_),
    .B(_1166_),
    .Y(_1167_));
 sg13g2_o21ai_1 _4105_ (.B1(_1158_),
    .Y(_1168_),
    .A1(_1165_),
    .A2(_1167_));
 sg13g2_xnor2_1 _4106_ (.Y(_1169_),
    .A(_1153_),
    .B(_1168_));
 sg13g2_nor2_1 _4107_ (.A(net1183),
    .B(_1115_),
    .Y(_1170_));
 sg13g2_nor2_1 _4108_ (.A(_1120_),
    .B(_1170_),
    .Y(_1171_));
 sg13g2_nand3_1 _4109_ (.B(_1158_),
    .C(_1164_),
    .A(_1145_),
    .Y(_1172_));
 sg13g2_o21ai_1 _4110_ (.B1(_1128_),
    .Y(_1173_),
    .A1(_1171_),
    .A2(_1172_));
 sg13g2_a21oi_1 _4111_ (.A1(_1117_),
    .A2(_1169_),
    .Y(_1174_),
    .B1(_1173_));
 sg13g2_o21ai_1 _4112_ (.B1(_1158_),
    .Y(_1175_),
    .A1(_1145_),
    .A2(_1166_));
 sg13g2_o21ai_1 _4113_ (.B1(_1117_),
    .Y(_1176_),
    .A1(_1165_),
    .A2(_1175_));
 sg13g2_and2_1 _4114_ (.A(_1114_),
    .B(_1170_),
    .X(_1177_));
 sg13g2_and2_1 _4115_ (.A(_1152_),
    .B(_1163_),
    .X(_1178_));
 sg13g2_or2_1 _4116_ (.X(_1179_),
    .B(_1178_),
    .A(_1175_));
 sg13g2_o21ai_1 _4117_ (.B1(_1163_),
    .Y(_1180_),
    .A1(_1145_),
    .A2(_1150_));
 sg13g2_and2_1 _4118_ (.A(_1144_),
    .B(_1158_),
    .X(_1181_));
 sg13g2_a22oi_1 _4119_ (.Y(_1182_),
    .B1(_1180_),
    .B2(_1158_),
    .A2(_1164_),
    .A1(_1145_));
 sg13g2_nand2_1 _4120_ (.Y(_1183_),
    .A(net1195),
    .B(_1127_));
 sg13g2_a221oi_1 _4121_ (.B2(_1120_),
    .C1(_1183_),
    .B1(_1182_),
    .A1(_1177_),
    .Y(_1184_),
    .A2(_1179_));
 sg13g2_a21oi_1 _4122_ (.A1(_1176_),
    .A2(_1184_),
    .Y(_1185_),
    .B1(_1174_));
 sg13g2_nand2_1 _4123_ (.Y(_1186_),
    .A(net1184),
    .B(_1119_));
 sg13g2_or2_1 _4124_ (.X(_1187_),
    .B(_1178_),
    .A(_1166_));
 sg13g2_a21oi_1 _4125_ (.A1(_1181_),
    .A2(_1187_),
    .Y(_1188_),
    .B1(_1186_));
 sg13g2_o21ai_1 _4126_ (.B1(_1121_),
    .Y(_1189_),
    .A1(net1184),
    .A2(_1118_));
 sg13g2_nor3_1 _4127_ (.A(_1185_),
    .B(_1188_),
    .C(_1189_),
    .Y(_1190_));
 sg13g2_nand2b_1 _4128_ (.Y(_1191_),
    .B(_1121_),
    .A_N(_1116_));
 sg13g2_nor2b_1 _4129_ (.A(_1187_),
    .B_N(_1158_),
    .Y(_1192_));
 sg13g2_a221oi_1 _4130_ (.B2(_1144_),
    .C1(net1195),
    .B1(_1120_),
    .A1(net1184),
    .Y(_1193_),
    .A2(_1119_));
 sg13g2_nand2_1 _4131_ (.Y(_1194_),
    .A(_1127_),
    .B(_1193_));
 sg13g2_a21oi_1 _4132_ (.A1(_1165_),
    .A2(_1177_),
    .Y(_1195_),
    .B1(_1194_));
 sg13g2_o21ai_1 _4133_ (.B1(_1195_),
    .Y(_1196_),
    .A1(_1171_),
    .A2(_1192_));
 sg13g2_a21oi_1 _4134_ (.A1(_1172_),
    .A2(_1191_),
    .Y(_1197_),
    .B1(_1196_));
 sg13g2_and4_1 _4135_ (.A(_1128_),
    .B(_1178_),
    .C(_1181_),
    .D(_1189_),
    .X(_1198_));
 sg13g2_nor2_1 _4136_ (.A(net1887),
    .B(net1579),
    .Y(_1199_));
 sg13g2_nor2_1 _4137_ (.A(net1180),
    .B(net1182),
    .Y(_1200_));
 sg13g2_nand2b_1 _4138_ (.Y(_1201_),
    .B(_1200_),
    .A_N(_0871_));
 sg13g2_nand2_1 _4139_ (.Y(_1202_),
    .A(_0777_),
    .B(_1201_));
 sg13g2_and3_1 _4140_ (.X(_1203_),
    .A(_0624_),
    .B(net1179),
    .C(_0777_));
 sg13g2_inv_1 _4141_ (.Y(_1204_),
    .A(_1203_));
 sg13g2_nor4_1 _4142_ (.A(\vga_tetris._vgaController_io_pixelPosY[9] ),
    .B(_0775_),
    .C(_0867_),
    .D(_1203_),
    .Y(_1205_));
 sg13g2_a22oi_1 _4143_ (.Y(_1206_),
    .B1(_1202_),
    .B2(_1205_),
    .A2(_1199_),
    .A1(_0902_));
 sg13g2_or2_1 _4144_ (.X(_1207_),
    .B(\vga_tetris._vgaController_io_pixelPosX[0] ),
    .A(net1599));
 sg13g2_a21oi_1 _4145_ (.A1(_0898_),
    .A2(_1008_),
    .Y(_1208_),
    .B1(_0902_));
 sg13g2_nor4_1 _4146_ (.A(_1123_),
    .B(_1206_),
    .C(_1207_),
    .D(_1208_),
    .Y(_1209_));
 sg13g2_nor2_1 _4147_ (.A(net1640),
    .B(_0625_),
    .Y(_1210_));
 sg13g2_nor4_1 _4148_ (.A(\vga_tetris._vgaController_io_pixelPosY[9] ),
    .B(_0776_),
    .C(_0869_),
    .D(_1210_),
    .Y(_1211_));
 sg13g2_a22oi_1 _4149_ (.Y(_1212_),
    .B1(_1211_),
    .B2(_0774_),
    .A2(_0775_),
    .A1(_0624_));
 sg13g2_nor2_1 _4150_ (.A(_1201_),
    .B(_1212_),
    .Y(_1213_));
 sg13g2_nand2_1 _4151_ (.Y(_1214_),
    .A(net1182),
    .B(_0879_));
 sg13g2_nor3_1 _4152_ (.A(net1180),
    .B(_1204_),
    .C(_1214_),
    .Y(_1215_));
 sg13g2_nor4_1 _4153_ (.A(_0626_),
    .B(\vga_tetris._vgaController_io_pixelPosX[8] ),
    .C(_0876_),
    .D(_0951_),
    .Y(_1216_));
 sg13g2_nor4_1 _4154_ (.A(_1209_),
    .B(_1213_),
    .C(_1215_),
    .D(_1216_),
    .Y(_1217_));
 sg13g2_nor2_1 _4155_ (.A(_0870_),
    .B(_1103_),
    .Y(_1218_));
 sg13g2_nand3_1 _4156_ (.B(_1217_),
    .C(_1218_),
    .A(_1131_),
    .Y(_1219_));
 sg13g2_nor4_1 _4157_ (.A(_1133_),
    .B(_1197_),
    .C(_1198_),
    .D(_1219_),
    .Y(_1220_));
 sg13g2_nand2b_2 _4158_ (.Y(_1221_),
    .B(_1220_),
    .A_N(_1190_));
 sg13g2_a21oi_1 _4159_ (.A1(net1185),
    .A2(net1189),
    .Y(_1222_),
    .B1(net1183));
 sg13g2_nand2b_1 _4160_ (.Y(_1223_),
    .B(net1180),
    .A_N(_1222_));
 sg13g2_nand2b_1 _4161_ (.Y(_1224_),
    .B(_1222_),
    .A_N(net1180));
 sg13g2_and2_1 _4162_ (.A(_1223_),
    .B(_1224_),
    .X(_1225_));
 sg13g2_nand2b_1 _4163_ (.Y(_1226_),
    .B(_1225_),
    .A_N(net1189));
 sg13g2_or2_1 _4164_ (.X(_1227_),
    .B(_1226_),
    .A(net1183));
 sg13g2_or2_1 _4165_ (.X(_1228_),
    .B(_1226_),
    .A(net1186));
 sg13g2_nor2_1 _4166_ (.A(net1185),
    .B(_1227_),
    .Y(_1229_));
 sg13g2_nand2_2 _4167_ (.Y(_1230_),
    .A(net1180),
    .B(net1182));
 sg13g2_o21ai_1 _4168_ (.B1(_1226_),
    .Y(_1231_),
    .A1(net1186),
    .A2(_1230_));
 sg13g2_nand2b_2 _4169_ (.Y(_1232_),
    .B(net1189),
    .A_N(net1185));
 sg13g2_a21oi_1 _4170_ (.A1(net1185),
    .A2(_1106_),
    .Y(_1233_),
    .B1(_1223_));
 sg13g2_nand2_2 _4171_ (.Y(_1234_),
    .A(_1232_),
    .B(_1233_));
 sg13g2_nand4_1 _4172_ (.B(\vga_tetris._vgaController_io_pixelPosX[2] ),
    .C(_1227_),
    .A(_0627_),
    .Y(_1235_),
    .D(_1234_));
 sg13g2_a221oi_1 _4173_ (.B2(_0627_),
    .C1(_1229_),
    .B1(_1231_),
    .A1(_0873_),
    .Y(_1236_),
    .A2(_1123_));
 sg13g2_nor2b_1 _4174_ (.A(_1236_),
    .B_N(_1130_),
    .Y(_1237_));
 sg13g2_o21ai_1 _4175_ (.B1(_1231_),
    .Y(_1238_),
    .A1(_0627_),
    .A2(_1234_));
 sg13g2_a21oi_1 _4176_ (.A1(net1185),
    .A2(net1189),
    .Y(_1239_),
    .B1(_1200_));
 sg13g2_o21ai_1 _4177_ (.B1(net1181),
    .Y(_1240_),
    .A1(net1185),
    .A2(net1189));
 sg13g2_a21o_1 _4178_ (.A2(_1240_),
    .A1(_1239_),
    .B1(_0873_),
    .X(_1241_));
 sg13g2_a21oi_1 _4179_ (.A1(_1127_),
    .A2(_1238_),
    .Y(_1242_),
    .B1(_1130_));
 sg13g2_a22oi_1 _4180_ (.Y(_1243_),
    .B1(_1241_),
    .B2(_1242_),
    .A2(_1237_),
    .A1(_1235_));
 sg13g2_o21ai_1 _4181_ (.B1(net1194),
    .Y(_1244_),
    .A1(net1195),
    .A2(_1123_));
 sg13g2_xor2_1 _4182_ (.B(_1244_),
    .A(net1192),
    .X(_1245_));
 sg13g2_nand2b_1 _4183_ (.Y(_1246_),
    .B(_1245_),
    .A_N(_1243_));
 sg13g2_xnor2_1 _4184_ (.Y(_1247_),
    .A(net1194),
    .B(_1129_));
 sg13g2_nor2_1 _4185_ (.A(_1230_),
    .B(_1232_),
    .Y(_1248_));
 sg13g2_a21oi_1 _4186_ (.A1(net1182),
    .A2(_1232_),
    .Y(_1249_),
    .B1(_1222_));
 sg13g2_nor2b_1 _4187_ (.A(_1249_),
    .B_N(_1225_),
    .Y(_1250_));
 sg13g2_nor3_1 _4188_ (.A(_0873_),
    .B(_1229_),
    .C(_1233_),
    .Y(_1251_));
 sg13g2_nand3_1 _4189_ (.B(_1127_),
    .C(_1228_),
    .A(net1198),
    .Y(_1252_));
 sg13g2_nand2_1 _4190_ (.Y(_1253_),
    .A(_1127_),
    .B(_1229_));
 sg13g2_a21oi_1 _4191_ (.A1(_0628_),
    .A2(_1232_),
    .Y(_1254_),
    .B1(\vga_tetris._vgaController_io_pixelPosX[3] ));
 sg13g2_nand3_1 _4192_ (.B(_1230_),
    .C(_1239_),
    .A(_1106_),
    .Y(_1255_));
 sg13g2_a21oi_1 _4193_ (.A1(_1234_),
    .A2(_1255_),
    .Y(_1256_),
    .B1(_1254_));
 sg13g2_nor3_1 _4194_ (.A(net1195),
    .B(_1248_),
    .C(_1250_),
    .Y(_1257_));
 sg13g2_nor2_1 _4195_ (.A(_1251_),
    .B(_1257_),
    .Y(_1258_));
 sg13g2_a21oi_1 _4196_ (.A1(_1252_),
    .A2(_1258_),
    .Y(_1259_),
    .B1(_1130_));
 sg13g2_nand2_1 _4197_ (.Y(_1260_),
    .A(_1130_),
    .B(_1253_));
 sg13g2_nor3_1 _4198_ (.A(_1245_),
    .B(_1247_),
    .C(_1259_),
    .Y(_1261_));
 sg13g2_o21ai_1 _4199_ (.B1(_1261_),
    .Y(_1262_),
    .A1(_1256_),
    .A2(_1260_));
 sg13g2_a21oi_1 _4200_ (.A1(net1198),
    .A2(_1127_),
    .Y(_1263_),
    .B1(_1249_));
 sg13g2_o21ai_1 _4201_ (.B1(_0628_),
    .Y(_1264_),
    .A1(net1186),
    .A2(_1107_));
 sg13g2_nand2b_1 _4202_ (.Y(_1265_),
    .B(_1232_),
    .A_N(_0873_));
 sg13g2_nand3_1 _4203_ (.B(_1264_),
    .C(_1265_),
    .A(_1225_),
    .Y(_1266_));
 sg13g2_o21ai_1 _4204_ (.B1(_1266_),
    .Y(_1267_),
    .A1(_1225_),
    .A2(_1263_));
 sg13g2_a21oi_1 _4205_ (.A1(_1253_),
    .A2(_1267_),
    .Y(_1268_),
    .B1(_1130_));
 sg13g2_nor2_1 _4206_ (.A(net1198),
    .B(_1248_),
    .Y(_1269_));
 sg13g2_a21oi_1 _4207_ (.A1(net1198),
    .A2(_1234_),
    .Y(_1270_),
    .B1(_1269_));
 sg13g2_nand2b_1 _4208_ (.Y(_1271_),
    .B(_1127_),
    .A_N(_1250_));
 sg13g2_o21ai_1 _4209_ (.B1(_1130_),
    .Y(_1272_),
    .A1(_1270_),
    .A2(_1271_));
 sg13g2_o21ai_1 _4210_ (.B1(net1192),
    .Y(_1273_),
    .A1(_1251_),
    .A2(_1272_));
 sg13g2_o21ai_1 _4211_ (.B1(_1247_),
    .Y(_1274_),
    .A1(_1268_),
    .A2(_1273_));
 sg13g2_nor3_1 _4212_ (.A(\vga_tetris._vgaController_io_pixelPosY[9] ),
    .B(\vga_tetris._vgaController_io_pixelPosY[8] ),
    .C(_0781_),
    .Y(_1275_));
 sg13g2_nand3_1 _4213_ (.B(net1182),
    .C(net1185),
    .A(net1180),
    .Y(_1276_));
 sg13g2_nand4_1 _4214_ (.B(_1224_),
    .C(_1275_),
    .A(\vga_tetris._tetrisLogic_io_gameOver ),
    .Y(_1277_),
    .D(_1276_));
 sg13g2_nor3_1 _4215_ (.A(_0869_),
    .B(_1103_),
    .C(_1277_),
    .Y(_1278_));
 sg13g2_nand4_1 _4216_ (.B(_1262_),
    .C(_1274_),
    .A(_1246_),
    .Y(_1279_),
    .D(_1278_));
 sg13g2_and2_1 _4217_ (.A(_1217_),
    .B(_1279_),
    .X(_1280_));
 sg13g2_inv_1 _4218_ (.Y(_1281_),
    .A(_1280_));
 sg13g2_o21ai_1 _4219_ (.B1(_1221_),
    .Y(_1282_),
    .A1(_1103_),
    .A2(_1280_));
 sg13g2_or2_1 _4220_ (.X(uo_out[4]),
    .B(_1282_),
    .A(_1105_));
 sg13g2_nand3_1 _4221_ (.B(net1056),
    .C(net1020),
    .A(\vga_tetris.boardMem.board_8[9] ),
    .Y(_1283_));
 sg13g2_nand3_1 _4222_ (.B(net1032),
    .C(net1015),
    .A(\vga_tetris.boardMem.board_14[9] ),
    .Y(_1284_));
 sg13g2_nand3_1 _4223_ (.B(net1032),
    .C(net1020),
    .A(\vga_tetris.boardMem.board_12[9] ),
    .Y(_1285_));
 sg13g2_nand3_1 _4224_ (.B(net1039),
    .C(net1032),
    .A(\vga_tetris.boardMem.board_13[9] ),
    .Y(_1286_));
 sg13g2_nand3_1 _4225_ (.B(net1044),
    .C(net1039),
    .A(\vga_tetris.boardMem.board_1[9] ),
    .Y(_1287_));
 sg13g2_nand3_1 _4226_ (.B(net1056),
    .C(net1015),
    .A(\vga_tetris.boardMem.board_10[9] ),
    .Y(_1288_));
 sg13g2_nand3_1 _4227_ (.B(net1039),
    .C(net1026),
    .A(\vga_tetris.boardMem.board_17[9] ),
    .Y(_1289_));
 sg13g2_nand3_1 _4228_ (.B(net1015),
    .C(net1006),
    .A(\vga_tetris.boardMem.board_6[9] ),
    .Y(_1290_));
 sg13g2_and3_1 _4229_ (.X(_1291_),
    .A(\vga_tetris.boardMem.board_5[9] ),
    .B(net1039),
    .C(net1007));
 sg13g2_and4_1 _4230_ (.A(_1284_),
    .B(_1286_),
    .C(_1287_),
    .D(_1290_),
    .X(_1292_));
 sg13g2_a22oi_1 _4231_ (.Y(_1293_),
    .B1(net976),
    .B2(\vga_tetris.boardMem.board_7[9] ),
    .A2(net979),
    .A1(\vga_tetris.boardMem.board_4[9] ));
 sg13g2_a22oi_1 _4232_ (.Y(_1294_),
    .B1(_0850_),
    .B2(\vga_tetris.boardMem.board_2[9] ),
    .A2(net1001),
    .A1(\vga_tetris.boardMem.board_3[9] ));
 sg13g2_a22oi_1 _4233_ (.Y(_1295_),
    .B1(net989),
    .B2(\vga_tetris.boardMem.board_15[9] ),
    .A2(net998),
    .A1(\vga_tetris.boardMem.board_9[9] ));
 sg13g2_a221oi_1 _4234_ (.B2(\vga_tetris.boardMem.board_19[9] ),
    .C1(_1291_),
    .B1(net985),
    .A1(\vga_tetris.boardMem.board_11[9] ),
    .Y(_1296_),
    .A2(net1002));
 sg13g2_and4_1 _4235_ (.A(_1283_),
    .B(_1285_),
    .C(_1288_),
    .D(_1289_),
    .X(_1297_));
 sg13g2_nand4_1 _4236_ (.B(_1294_),
    .C(_1296_),
    .A(_1293_),
    .Y(_1298_),
    .D(_1297_));
 sg13g2_a22oi_1 _4237_ (.Y(_1299_),
    .B1(net983),
    .B2(\vga_tetris.boardMem.board_16[9] ),
    .A2(net991),
    .A1(\vga_tetris.boardMem.board_18[9] ));
 sg13g2_nand4_1 _4238_ (.B(_1292_),
    .C(_1295_),
    .A(net965),
    .Y(_1300_),
    .D(_1299_));
 sg13g2_a21oi_1 _4239_ (.A1(_0667_),
    .A2(net967),
    .Y(_1301_),
    .B1(net1066));
 sg13g2_o21ai_1 _4240_ (.B1(_1301_),
    .Y(_1302_),
    .A1(_1298_),
    .A2(_1300_));
 sg13g2_nor4_1 _4241_ (.A(net1193),
    .B(net1197),
    .C(_0946_),
    .D(_1302_),
    .Y(_1303_));
 sg13g2_nand3_1 _4242_ (.B(net1056),
    .C(net1039),
    .A(\vga_tetris.boardMem.board_9[19] ),
    .Y(_1304_));
 sg13g2_nand3_1 _4243_ (.B(net1050),
    .C(net1006),
    .A(\vga_tetris.boardMem.board_7[19] ),
    .Y(_1305_));
 sg13g2_nand3_1 _4244_ (.B(net1044),
    .C(net1015),
    .A(\vga_tetris.boardMem.board_2[19] ),
    .Y(_1306_));
 sg13g2_nand3_1 _4245_ (.B(net1050),
    .C(net1026),
    .A(\vga_tetris.boardMem.board_19[19] ),
    .Y(_1307_));
 sg13g2_nand3_1 _4246_ (.B(net1056),
    .C(net1020),
    .A(\vga_tetris.boardMem.board_8[19] ),
    .Y(_1308_));
 sg13g2_nand3_1 _4247_ (.B(net1020),
    .C(net1006),
    .A(\vga_tetris.boardMem.board_4[19] ),
    .Y(_1309_));
 sg13g2_nand3_1 _4248_ (.B(net1026),
    .C(net1020),
    .A(\vga_tetris.boardMem.board_16[19] ),
    .Y(_1310_));
 sg13g2_and3_1 _4249_ (.X(_1311_),
    .A(\vga_tetris.boardMem.board_14[19] ),
    .B(net1032),
    .C(net1015));
 sg13g2_nand3_1 _4250_ (.B(net1015),
    .C(net1006),
    .A(\vga_tetris.boardMem.board_6[19] ),
    .Y(_1312_));
 sg13g2_nand2_1 _4251_ (.Y(_1313_),
    .A(\vga_tetris.boardMem.board_3[19] ),
    .B(net1001));
 sg13g2_a221oi_1 _4252_ (.B2(\vga_tetris.boardMem.board_5[19] ),
    .C1(_1311_),
    .B1(net975),
    .A1(\vga_tetris.boardMem.board_12[19] ),
    .Y(_1314_),
    .A2(net992));
 sg13g2_a22oi_1 _4253_ (.Y(_1315_),
    .B1(net988),
    .B2(\vga_tetris.boardMem.board_10[19] ),
    .A2(net991),
    .A1(\vga_tetris.boardMem.board_18[19] ));
 sg13g2_a22oi_1 _4254_ (.Y(_1316_),
    .B1(net989),
    .B2(\vga_tetris.boardMem.board_15[19] ),
    .A2(net1002),
    .A1(\vga_tetris.boardMem.board_11[19] ));
 sg13g2_nand4_1 _4255_ (.B(_1314_),
    .C(_1315_),
    .A(_1313_),
    .Y(_1317_),
    .D(_1316_));
 sg13g2_and4_1 _4256_ (.A(_1304_),
    .B(_1307_),
    .C(_1308_),
    .D(_1309_),
    .X(_1318_));
 sg13g2_a22oi_1 _4257_ (.Y(_1319_),
    .B1(net969),
    .B2(\vga_tetris.boardMem.board_17[19] ),
    .A2(net999),
    .A1(\vga_tetris.boardMem.board_13[19] ));
 sg13g2_a22oi_1 _4258_ (.Y(_1320_),
    .B1(net972),
    .B2(\vga_tetris.boardMem.board_1[19] ),
    .A2(net993),
    .A1(net996));
 sg13g2_and4_1 _4259_ (.A(_1305_),
    .B(_1306_),
    .C(_1310_),
    .D(_1312_),
    .X(_1321_));
 sg13g2_nand4_1 _4260_ (.B(_1319_),
    .C(_1320_),
    .A(_1318_),
    .Y(_1322_),
    .D(_1321_));
 sg13g2_a21oi_1 _4261_ (.A1(_0674_),
    .A2(net967),
    .Y(_1323_),
    .B1(net1066));
 sg13g2_o21ai_1 _4262_ (.B1(_1323_),
    .Y(_1324_),
    .A1(_1317_),
    .A2(_1322_));
 sg13g2_or2_1 _4263_ (.X(_1325_),
    .B(_1324_),
    .A(_0990_));
 sg13g2_nand3_1 _4264_ (.B(net1038),
    .C(net1033),
    .A(\vga_tetris.boardMem.board_13[13] ),
    .Y(_1326_));
 sg13g2_and3_1 _4265_ (.X(_1327_),
    .A(\vga_tetris.boardMem.board_18[13] ),
    .B(net1026),
    .C(net1013));
 sg13g2_nand3_1 _4266_ (.B(net1050),
    .C(net1007),
    .A(\vga_tetris.boardMem.board_7[13] ),
    .Y(_1328_));
 sg13g2_nand3_1 _4267_ (.B(net1038),
    .C(net1006),
    .A(\vga_tetris.boardMem.board_5[13] ),
    .Y(_1329_));
 sg13g2_nand3_1 _4268_ (.B(net1056),
    .C(net1013),
    .A(\vga_tetris.boardMem.board_10[13] ),
    .Y(_1330_));
 sg13g2_nand3_1 _4269_ (.B(net1050),
    .C(net1026),
    .A(\vga_tetris.boardMem.board_19[13] ),
    .Y(_1331_));
 sg13g2_a22oi_1 _4270_ (.Y(_1332_),
    .B1(net984),
    .B2(\vga_tetris.boardMem.board_16[13] ),
    .A2(net1003),
    .A1(\vga_tetris.boardMem.board_11[13] ));
 sg13g2_nand3_1 _4271_ (.B(net1032),
    .C(net1020),
    .A(\vga_tetris.boardMem.board_12[13] ),
    .Y(_1333_));
 sg13g2_nand3_1 _4272_ (.B(net1045),
    .C(net1039),
    .A(\vga_tetris.boardMem.board_1[13] ),
    .Y(_1334_));
 sg13g2_nand3_1 _4273_ (.B(net1056),
    .C(net1020),
    .A(\vga_tetris.boardMem.board_8[13] ),
    .Y(_1335_));
 sg13g2_and4_1 _4274_ (.A(_1328_),
    .B(_1329_),
    .C(_1331_),
    .D(_1334_),
    .X(_1336_));
 sg13g2_a22oi_1 _4275_ (.Y(_1337_),
    .B1(_0850_),
    .B2(\vga_tetris.boardMem.board_2[13] ),
    .A2(net982),
    .A1(\vga_tetris.boardMem.board_6[13] ));
 sg13g2_a22oi_1 _4276_ (.Y(_1338_),
    .B1(net979),
    .B2(\vga_tetris.boardMem.board_4[13] ),
    .A2(net1001),
    .A1(\vga_tetris.boardMem.board_3[13] ));
 sg13g2_a221oi_1 _4277_ (.B2(\vga_tetris.boardMem.board_14[13] ),
    .C1(_1327_),
    .B1(net971),
    .A1(\vga_tetris.boardMem.board_15[13] ),
    .Y(_1339_),
    .A2(net989));
 sg13g2_and4_1 _4278_ (.A(_1326_),
    .B(_1330_),
    .C(_1333_),
    .D(_1335_),
    .X(_1340_));
 sg13g2_nand4_1 _4279_ (.B(_1338_),
    .C(_1339_),
    .A(_1337_),
    .Y(_1341_),
    .D(_1340_));
 sg13g2_a22oi_1 _4280_ (.Y(_1342_),
    .B1(net970),
    .B2(\vga_tetris.boardMem.board_17[13] ),
    .A2(net998),
    .A1(\vga_tetris.boardMem.board_9[13] ));
 sg13g2_nand4_1 _4281_ (.B(_1332_),
    .C(_1336_),
    .A(net966),
    .Y(_1343_),
    .D(_1342_));
 sg13g2_a21oi_1 _4282_ (.A1(_0671_),
    .A2(net968),
    .Y(_1344_),
    .B1(net1066));
 sg13g2_o21ai_1 _4283_ (.B1(_1344_),
    .Y(_1345_),
    .A1(_1341_),
    .A2(_1343_));
 sg13g2_or2_1 _4284_ (.X(_1346_),
    .B(_1345_),
    .A(_1071_));
 sg13g2_nand3_1 _4285_ (.B(net1028),
    .C(net1017),
    .A(\vga_tetris.boardMem.board_12[15] ),
    .Y(_1347_));
 sg13g2_nand3_1 _4286_ (.B(net1041),
    .C(net1037),
    .A(\vga_tetris.boardMem.board_1[15] ),
    .Y(_1348_));
 sg13g2_and3_1 _4287_ (.X(_1349_),
    .A(\vga_tetris.boardMem.board_18[15] ),
    .B(net1023),
    .C(net1008));
 sg13g2_nand3_1 _4288_ (.B(net1037),
    .C(net1028),
    .A(\vga_tetris.boardMem.board_13[15] ),
    .Y(_1350_));
 sg13g2_nand3_1 _4289_ (.B(net1046),
    .C(net1023),
    .A(\vga_tetris.boardMem.board_19[15] ),
    .Y(_1351_));
 sg13g2_nand3_1 _4290_ (.B(net1028),
    .C(net1008),
    .A(\vga_tetris.boardMem.board_14[15] ),
    .Y(_1352_));
 sg13g2_nand3_1 _4291_ (.B(net1008),
    .C(net1005),
    .A(\vga_tetris.boardMem.board_6[15] ),
    .Y(_1353_));
 sg13g2_nand3_1 _4292_ (.B(net1046),
    .C(net1041),
    .A(\vga_tetris.boardMem.board_3[15] ),
    .Y(_1354_));
 sg13g2_nand3_1 _4293_ (.B(net1052),
    .C(net1017),
    .A(\vga_tetris.boardMem.board_8[15] ),
    .Y(_1355_));
 sg13g2_a22oi_1 _4294_ (.Y(_1356_),
    .B1(net977),
    .B2(\vga_tetris.boardMem.board_7[15] ),
    .A2(net978),
    .A1(\vga_tetris.boardMem.board_2[15] ));
 sg13g2_a22oi_1 _4295_ (.Y(_1357_),
    .B1(net969),
    .B2(\vga_tetris.boardMem.board_17[15] ),
    .A2(net983),
    .A1(\vga_tetris.boardMem.board_16[15] ));
 sg13g2_a22oi_1 _4296_ (.Y(_1358_),
    .B1(net974),
    .B2(\vga_tetris.boardMem.board_5[15] ),
    .A2(net997),
    .A1(\vga_tetris.boardMem.board_9[15] ));
 sg13g2_a22oi_1 _4297_ (.Y(_1359_),
    .B1(net980),
    .B2(\vga_tetris.boardMem.board_4[15] ),
    .A2(net987),
    .A1(\vga_tetris.boardMem.board_10[15] ));
 sg13g2_a221oi_1 _4298_ (.B2(\vga_tetris.boardMem.board_15[15] ),
    .C1(_1349_),
    .B1(net990),
    .A1(\vga_tetris.boardMem.board_11[15] ),
    .Y(_1360_),
    .A2(net1003));
 sg13g2_and4_1 _4299_ (.A(_1347_),
    .B(_1353_),
    .C(_1354_),
    .D(_1355_),
    .X(_1361_));
 sg13g2_nand4_1 _4300_ (.B(_1357_),
    .C(_1360_),
    .A(_1356_),
    .Y(_1362_),
    .D(_1361_));
 sg13g2_and4_1 _4301_ (.A(_1348_),
    .B(_1350_),
    .C(_1351_),
    .D(_1352_),
    .X(_1363_));
 sg13g2_nand4_1 _4302_ (.B(_1358_),
    .C(_1359_),
    .A(net964),
    .Y(_1364_),
    .D(_1363_));
 sg13g2_a21oi_1 _4303_ (.A1(_0673_),
    .A2(net967),
    .Y(_1365_),
    .B1(net1065));
 sg13g2_o21ai_1 _4304_ (.B1(_1365_),
    .Y(_1366_),
    .A1(_1362_),
    .A2(_1364_));
 sg13g2_nand3_1 _4305_ (.B(net1042),
    .C(net1036),
    .A(\vga_tetris.boardMem.board_1[7] ),
    .Y(_1367_));
 sg13g2_nand3_1 _4306_ (.B(net1029),
    .C(net1011),
    .A(\vga_tetris.boardMem.board_14[7] ),
    .Y(_1368_));
 sg13g2_nand3_1 _4307_ (.B(net1029),
    .C(net1019),
    .A(\vga_tetris.boardMem.board_12[7] ),
    .Y(_1369_));
 sg13g2_nand3_1 _4308_ (.B(net1010),
    .C(net1004),
    .A(\vga_tetris.boardMem.board_6[7] ),
    .Y(_1370_));
 sg13g2_and3_1 _4309_ (.X(_1371_),
    .A(\vga_tetris.boardMem.board_18[7] ),
    .B(net1024),
    .C(net1010));
 sg13g2_nand3_1 _4310_ (.B(net1049),
    .C(net1042),
    .A(\vga_tetris.boardMem.board_3[7] ),
    .Y(_1372_));
 sg13g2_nand3_1 _4311_ (.B(net1049),
    .C(net1024),
    .A(\vga_tetris.boardMem.board_19[7] ),
    .Y(_1373_));
 sg13g2_nand3_1 _4312_ (.B(net1054),
    .C(net1019),
    .A(\vga_tetris.boardMem.board_8[7] ),
    .Y(_1374_));
 sg13g2_nand3_1 _4313_ (.B(net1036),
    .C(net1030),
    .A(\vga_tetris.boardMem.board_13[7] ),
    .Y(_1375_));
 sg13g2_a22oi_1 _4314_ (.Y(_1376_),
    .B1(net969),
    .B2(\vga_tetris.boardMem.board_17[7] ),
    .A2(net990),
    .A1(\vga_tetris.boardMem.board_15[7] ));
 sg13g2_a22oi_1 _4315_ (.Y(_1377_),
    .B1(net977),
    .B2(\vga_tetris.boardMem.board_7[7] ),
    .A2(net978),
    .A1(\vga_tetris.boardMem.board_2[7] ));
 sg13g2_a22oi_1 _4316_ (.Y(_1378_),
    .B1(net974),
    .B2(\vga_tetris.boardMem.board_5[7] ),
    .A2(net997),
    .A1(\vga_tetris.boardMem.board_9[7] ));
 sg13g2_a22oi_1 _4317_ (.Y(_1379_),
    .B1(net980),
    .B2(\vga_tetris.boardMem.board_4[7] ),
    .A2(net987),
    .A1(\vga_tetris.boardMem.board_10[7] ));
 sg13g2_a221oi_1 _4318_ (.B2(\vga_tetris.boardMem.board_16[7] ),
    .C1(_1371_),
    .B1(net983),
    .A1(\vga_tetris.boardMem.board_11[7] ),
    .Y(_1380_),
    .A2(net1003));
 sg13g2_and4_1 _4319_ (.A(_1369_),
    .B(_1370_),
    .C(_1372_),
    .D(_1374_),
    .X(_1381_));
 sg13g2_and4_1 _4320_ (.A(_1376_),
    .B(_1377_),
    .C(_1380_),
    .D(_1381_),
    .X(_1382_));
 sg13g2_and4_1 _4321_ (.A(_1367_),
    .B(_1368_),
    .C(_1373_),
    .D(_1375_),
    .X(_1383_));
 sg13g2_and4_1 _4322_ (.A(net964),
    .B(_1378_),
    .C(_1379_),
    .D(_1383_),
    .X(_1384_));
 sg13g2_o21ai_1 _4323_ (.B1(net1068),
    .Y(_1385_),
    .A1(net1556),
    .A2(net964));
 sg13g2_a21oi_2 _4324_ (.B1(_1385_),
    .Y(_1386_),
    .A2(_1384_),
    .A1(_1382_));
 sg13g2_a21o_2 _4325_ (.A2(_1384_),
    .A1(_1382_),
    .B1(_1385_),
    .X(_1387_));
 sg13g2_nand3_1 _4326_ (.B(net1046),
    .C(net1043),
    .A(\vga_tetris.boardMem.board_3[11] ),
    .Y(_1388_));
 sg13g2_nand3_1 _4327_ (.B(net1047),
    .C(net1025),
    .A(\vga_tetris.boardMem.board_19[11] ),
    .Y(_1389_));
 sg13g2_nand3_1 _4328_ (.B(net1025),
    .C(net1016),
    .A(\vga_tetris.boardMem.board_18[11] ),
    .Y(_1390_));
 sg13g2_nand3_1 _4329_ (.B(net1031),
    .C(net1012),
    .A(\vga_tetris.boardMem.board_14[11] ),
    .Y(_1391_));
 sg13g2_nand3_1 _4330_ (.B(net1053),
    .C(net1022),
    .A(\vga_tetris.boardMem.board_8[11] ),
    .Y(_1392_));
 sg13g2_nand3_1 _4331_ (.B(net1053),
    .C(net1037),
    .A(\vga_tetris.boardMem.board_9[11] ),
    .Y(_1393_));
 sg13g2_and3_1 _4332_ (.X(_1394_),
    .A(\vga_tetris.boardMem.board_16[11] ),
    .B(net1025),
    .C(net1017));
 sg13g2_nand3_1 _4333_ (.B(net1037),
    .C(net1005),
    .A(\vga_tetris.boardMem.board_5[11] ),
    .Y(_1395_));
 sg13g2_nand3_1 _4334_ (.B(net1047),
    .C(net1031),
    .A(\vga_tetris.boardMem.board_15[11] ),
    .Y(_1396_));
 sg13g2_a22oi_1 _4335_ (.Y(_1397_),
    .B1(net972),
    .B2(\vga_tetris.boardMem.board_1[11] ),
    .A2(net980),
    .A1(\vga_tetris.boardMem.board_4[11] ));
 sg13g2_a22oi_1 _4336_ (.Y(_1398_),
    .B1(net977),
    .B2(\vga_tetris.boardMem.board_7[11] ),
    .A2(net987),
    .A1(\vga_tetris.boardMem.board_10[11] ));
 sg13g2_a22oi_1 _4337_ (.Y(_1399_),
    .B1(net969),
    .B2(\vga_tetris.boardMem.board_17[11] ),
    .A2(net981),
    .A1(\vga_tetris.boardMem.board_6[11] ));
 sg13g2_a22oi_1 _4338_ (.Y(_1400_),
    .B1(net978),
    .B2(\vga_tetris.boardMem.board_2[11] ),
    .A2(net999),
    .A1(\vga_tetris.boardMem.board_13[11] ));
 sg13g2_nand4_1 _4339_ (.B(_1398_),
    .C(_1399_),
    .A(_1397_),
    .Y(_1401_),
    .D(_1400_));
 sg13g2_a221oi_1 _4340_ (.B2(\vga_tetris.boardMem.board_12[11] ),
    .C1(_1394_),
    .B1(net992),
    .A1(\vga_tetris.boardMem.board_11[11] ),
    .Y(_1402_),
    .A2(net1003));
 sg13g2_and4_1 _4341_ (.A(_1388_),
    .B(_1390_),
    .C(_1392_),
    .D(_1395_),
    .X(_1403_));
 sg13g2_and4_1 _4342_ (.A(_1389_),
    .B(_1391_),
    .C(_1393_),
    .D(_1396_),
    .X(_1404_));
 sg13g2_nand4_1 _4343_ (.B(_1402_),
    .C(_1403_),
    .A(net966),
    .Y(_1405_),
    .D(_1404_));
 sg13g2_a21oi_1 _4344_ (.A1(_0669_),
    .A2(net967),
    .Y(_1406_),
    .B1(net1065));
 sg13g2_o21ai_1 _4345_ (.B1(_1406_),
    .Y(_1407_),
    .A1(_1401_),
    .A2(_1405_));
 sg13g2_nand2_1 _4346_ (.Y(_1408_),
    .A(\vga_tetris.boardMem.board_12[1] ),
    .B(net992));
 sg13g2_a22oi_1 _4347_ (.Y(_1409_),
    .B1(net975),
    .B2(\vga_tetris.boardMem.board_5[1] ),
    .A2(_0821_),
    .A1(\vga_tetris.boardMem.board_3[1] ));
 sg13g2_a22oi_1 _4348_ (.Y(_1410_),
    .B1(net982),
    .B2(\vga_tetris.boardMem.board_6[1] ),
    .A2(net984),
    .A1(\vga_tetris.boardMem.board_16[1] ));
 sg13g2_a22oi_1 _4349_ (.Y(_1411_),
    .B1(_0848_),
    .B2(\vga_tetris.boardMem.board_8[1] ),
    .A2(net1002),
    .A1(\vga_tetris.boardMem.board_11[1] ));
 sg13g2_a22oi_1 _4350_ (.Y(_1412_),
    .B1(net979),
    .B2(\vga_tetris.boardMem.board_4[1] ),
    .A2(net986),
    .A1(\vga_tetris.boardMem.board_19[1] ));
 sg13g2_nand4_1 _4351_ (.B(_1410_),
    .C(_1411_),
    .A(_1409_),
    .Y(_1413_),
    .D(_1412_));
 sg13g2_a22oi_1 _4352_ (.Y(_1414_),
    .B1(net973),
    .B2(\vga_tetris.boardMem.board_1[1] ),
    .A2(_0850_),
    .A1(\vga_tetris.boardMem.board_2[1] ));
 sg13g2_a22oi_1 _4353_ (.Y(_1415_),
    .B1(net970),
    .B2(\vga_tetris.boardMem.board_17[1] ),
    .A2(net988),
    .A1(\vga_tetris.boardMem.board_10[1] ));
 sg13g2_a22oi_1 _4354_ (.Y(_1416_),
    .B1(net991),
    .B2(\vga_tetris.boardMem.board_18[1] ),
    .A2(net998),
    .A1(\vga_tetris.boardMem.board_9[1] ));
 sg13g2_a22oi_1 _4355_ (.Y(_1417_),
    .B1(net976),
    .B2(\vga_tetris.boardMem.board_7[1] ),
    .A2(net989),
    .A1(\vga_tetris.boardMem.board_15[1] ));
 sg13g2_nand4_1 _4356_ (.B(_1415_),
    .C(_1416_),
    .A(_1414_),
    .Y(_1418_),
    .D(_1417_));
 sg13g2_a22oi_1 _4357_ (.Y(_1419_),
    .B1(net971),
    .B2(\vga_tetris.boardMem.board_14[1] ),
    .A2(net1000),
    .A1(\vga_tetris.boardMem.board_13[1] ));
 sg13g2_nand3_1 _4358_ (.B(_1408_),
    .C(_1419_),
    .A(net965),
    .Y(_1420_));
 sg13g2_nor3_2 _4359_ (.A(_1413_),
    .B(_1418_),
    .C(_1420_),
    .Y(_1421_));
 sg13g2_o21ai_1 _4360_ (.B1(net1068),
    .Y(_1422_),
    .A1(\vga_tetris.boardMem.board_0[1] ),
    .A2(net965));
 sg13g2_nor2_2 _4361_ (.A(_1421_),
    .B(_1422_),
    .Y(_1423_));
 sg13g2_a22oi_1 _4362_ (.Y(_1424_),
    .B1(_0856_),
    .B2(\vga_tetris.boardMem.board_14[3] ),
    .A2(net1000),
    .A1(\vga_tetris.boardMem.board_13[3] ));
 sg13g2_a22oi_1 _4363_ (.Y(_1425_),
    .B1(net979),
    .B2(\vga_tetris.boardMem.board_4[3] ),
    .A2(_0834_),
    .A1(\vga_tetris.boardMem.board_12[3] ));
 sg13g2_a22oi_1 _4364_ (.Y(_1426_),
    .B1(net988),
    .B2(\vga_tetris.boardMem.board_10[3] ),
    .A2(net994),
    .A1(net996));
 sg13g2_a22oi_1 _4365_ (.Y(_1427_),
    .B1(net976),
    .B2(\vga_tetris.boardMem.board_7[3] ),
    .A2(net982),
    .A1(\vga_tetris.boardMem.board_6[3] ));
 sg13g2_and4_1 _4366_ (.A(_1424_),
    .B(_1425_),
    .C(_1426_),
    .D(_1427_),
    .X(_1428_));
 sg13g2_a22oi_1 _4367_ (.Y(_1429_),
    .B1(_0848_),
    .B2(\vga_tetris.boardMem.board_8[3] ),
    .A2(_0837_),
    .A1(\vga_tetris.boardMem.board_18[3] ));
 sg13g2_a22oi_1 _4368_ (.Y(_1430_),
    .B1(net975),
    .B2(\vga_tetris.boardMem.board_5[3] ),
    .A2(net986),
    .A1(\vga_tetris.boardMem.board_19[3] ));
 sg13g2_nand3_1 _4369_ (.B(net1051),
    .C(net1045),
    .A(\vga_tetris.boardMem.board_3[3] ),
    .Y(_1431_));
 sg13g2_nand3_1 _4370_ (.B(net1040),
    .C(net1027),
    .A(\vga_tetris.boardMem.board_17[3] ),
    .Y(_1432_));
 sg13g2_nand3_1 _4371_ (.B(net1058),
    .C(net1040),
    .A(\vga_tetris.boardMem.board_9[3] ),
    .Y(_1433_));
 sg13g2_nand3_1 _4372_ (.B(net1058),
    .C(net1051),
    .A(\vga_tetris.boardMem.board_11[3] ),
    .Y(_1434_));
 sg13g2_and4_1 _4373_ (.A(_1431_),
    .B(_1432_),
    .C(_1433_),
    .D(_1434_),
    .X(_1435_));
 sg13g2_nand3_1 _4374_ (.B(net1050),
    .C(net1032),
    .A(\vga_tetris.boardMem.board_15[3] ),
    .Y(_1436_));
 sg13g2_nand3_1 _4375_ (.B(net1044),
    .C(net1040),
    .A(\vga_tetris.boardMem.board_1[3] ),
    .Y(_1437_));
 sg13g2_nand3_1 _4376_ (.B(net1044),
    .C(net1014),
    .A(\vga_tetris.boardMem.board_2[3] ),
    .Y(_1438_));
 sg13g2_nand3_1 _4377_ (.B(net1027),
    .C(net1021),
    .A(\vga_tetris.boardMem.board_16[3] ),
    .Y(_1439_));
 sg13g2_and4_1 _4378_ (.A(_1436_),
    .B(_1437_),
    .C(_1438_),
    .D(_1439_),
    .X(_1440_));
 sg13g2_and4_1 _4379_ (.A(_1429_),
    .B(_1430_),
    .C(_1435_),
    .D(_1440_),
    .X(_1441_));
 sg13g2_o21ai_1 _4380_ (.B1(_0891_),
    .Y(_1442_),
    .A1(\vga_tetris.boardMem.board_0[3] ),
    .A2(net965));
 sg13g2_a21oi_2 _4381_ (.B1(_1442_),
    .Y(_1443_),
    .A2(_1441_),
    .A1(_1428_));
 sg13g2_nand3_1 _4382_ (.B(_0947_),
    .C(_1443_),
    .A(_0901_),
    .Y(_1444_));
 sg13g2_nand3_1 _4383_ (.B(net1054),
    .C(net1010),
    .A(\vga_tetris.boardMem.board_10[17] ),
    .Y(_1445_));
 sg13g2_nand3_1 _4384_ (.B(net1054),
    .C(net1035),
    .A(\vga_tetris.boardMem.board_9[17] ),
    .Y(_1446_));
 sg13g2_nand3_1 _4385_ (.B(net1024),
    .C(net1010),
    .A(\vga_tetris.boardMem.board_18[17] ),
    .Y(_1447_));
 sg13g2_nand3_1 _4386_ (.B(net1029),
    .C(net1018),
    .A(\vga_tetris.boardMem.board_12[17] ),
    .Y(_1448_));
 sg13g2_nand3_1 _4387_ (.B(net1035),
    .C(net1004),
    .A(\vga_tetris.boardMem.board_5[17] ),
    .Y(_1449_));
 sg13g2_and3_1 _4388_ (.X(_1450_),
    .A(\vga_tetris.boardMem.board_4[17] ),
    .B(net1019),
    .C(net1005));
 sg13g2_nand3_1 _4389_ (.B(net1042),
    .C(net1011),
    .A(\vga_tetris.boardMem.board_2[17] ),
    .Y(_1451_));
 sg13g2_nand3_1 _4390_ (.B(net1029),
    .C(net1010),
    .A(\vga_tetris.boardMem.board_14[17] ),
    .Y(_1452_));
 sg13g2_nand3_1 _4391_ (.B(net1048),
    .C(net1042),
    .A(\vga_tetris.boardMem.board_3[17] ),
    .Y(_1453_));
 sg13g2_a22oi_1 _4392_ (.Y(_1454_),
    .B1(net977),
    .B2(\vga_tetris.boardMem.board_7[17] ),
    .A2(_0848_),
    .A1(\vga_tetris.boardMem.board_8[17] ));
 sg13g2_a22oi_1 _4393_ (.Y(_1455_),
    .B1(net999),
    .B2(\vga_tetris.boardMem.board_13[17] ),
    .A2(net1003),
    .A1(\vga_tetris.boardMem.board_11[17] ));
 sg13g2_a22oi_1 _4394_ (.Y(_1456_),
    .B1(net985),
    .B2(\vga_tetris.boardMem.board_19[17] ),
    .A2(net990),
    .A1(\vga_tetris.boardMem.board_15[17] ));
 sg13g2_a22oi_1 _4395_ (.Y(_1457_),
    .B1(net969),
    .B2(\vga_tetris.boardMem.board_17[17] ),
    .A2(net981),
    .A1(\vga_tetris.boardMem.board_6[17] ));
 sg13g2_a221oi_1 _4396_ (.B2(\vga_tetris.boardMem.board_1[17] ),
    .C1(_1450_),
    .B1(net972),
    .A1(\vga_tetris.boardMem.board_16[17] ),
    .Y(_1458_),
    .A2(net983));
 sg13g2_and4_1 _4397_ (.A(_1446_),
    .B(_1447_),
    .C(_1448_),
    .D(_1449_),
    .X(_1459_));
 sg13g2_nand4_1 _4398_ (.B(_1455_),
    .C(_1458_),
    .A(_1454_),
    .Y(_1460_),
    .D(_1459_));
 sg13g2_and4_1 _4399_ (.A(_1445_),
    .B(_1451_),
    .C(_1452_),
    .D(_1453_),
    .X(_1461_));
 sg13g2_nand4_1 _4400_ (.B(_1456_),
    .C(_1457_),
    .A(net964),
    .Y(_1462_),
    .D(_1461_));
 sg13g2_nand3b_1 _4401_ (.B(net995),
    .C(net993),
    .Y(_1463_),
    .A_N(\vga_tetris.boardMem.board_0[17] ));
 sg13g2_and2_1 _4402_ (.A(net1068),
    .B(_1463_),
    .X(_1464_));
 sg13g2_o21ai_1 _4403_ (.B1(_1463_),
    .Y(_1465_),
    .A1(_1460_),
    .A2(_1462_));
 sg13g2_nor2_1 _4404_ (.A(net1065),
    .B(_1465_),
    .Y(_1466_));
 sg13g2_o21ai_1 _4405_ (.B1(_1464_),
    .Y(_1467_),
    .A1(_1460_),
    .A2(_1462_));
 sg13g2_and3_1 _4406_ (.X(_1468_),
    .A(_0898_),
    .B(_0899_),
    .C(_1466_));
 sg13g2_nand3_1 _4407_ (.B(net1052),
    .C(net1010),
    .A(\vga_tetris.boardMem.board_10[5] ),
    .Y(_1469_));
 sg13g2_nand3_1 _4408_ (.B(net1024),
    .C(net1010),
    .A(\vga_tetris.boardMem.board_18[5] ),
    .Y(_1470_));
 sg13g2_nand3_1 _4409_ (.B(net1041),
    .C(net1010),
    .A(\vga_tetris.boardMem.board_2[5] ),
    .Y(_1471_));
 sg13g2_nand2_1 _4410_ (.Y(_1472_),
    .A(\vga_tetris.boardMem.board_1[5] ),
    .B(net972));
 sg13g2_and3_1 _4411_ (.X(_1473_),
    .A(\vga_tetris.boardMem.board_7[5] ),
    .B(net1046),
    .C(net1005));
 sg13g2_nand3_1 _4412_ (.B(net1054),
    .C(net1018),
    .A(\vga_tetris.boardMem.board_8[5] ),
    .Y(_1474_));
 sg13g2_nand3_1 _4413_ (.B(net1029),
    .C(net1018),
    .A(\vga_tetris.boardMem.board_12[5] ),
    .Y(_1475_));
 sg13g2_nand3_1 _4414_ (.B(net1024),
    .C(net1018),
    .A(\vga_tetris.boardMem.board_16[5] ),
    .Y(_1476_));
 sg13g2_nand3_1 _4415_ (.B(net1054),
    .C(net1048),
    .A(\vga_tetris.boardMem.board_11[5] ),
    .Y(_1477_));
 sg13g2_and3_1 _4416_ (.X(_1478_),
    .A(\vga_tetris.boardMem.board_17[5] ),
    .B(net1036),
    .C(net1025));
 sg13g2_and3_1 _4417_ (.X(_1479_),
    .A(\vga_tetris.boardMem.board_3[5] ),
    .B(net1048),
    .C(net1042));
 sg13g2_nand3_1 _4418_ (.B(net1054),
    .C(net1035),
    .A(\vga_tetris.boardMem.board_9[5] ),
    .Y(_1480_));
 sg13g2_nand3_1 _4419_ (.B(net1048),
    .C(net1024),
    .A(\vga_tetris.boardMem.board_19[5] ),
    .Y(_1481_));
 sg13g2_a221oi_1 _4420_ (.B2(\vga_tetris.boardMem.board_5[5] ),
    .C1(_1479_),
    .B1(net974),
    .A1(\vga_tetris.boardMem.board_15[5] ),
    .Y(_1482_),
    .A2(net990));
 sg13g2_a221oi_1 _4421_ (.B2(\vga_tetris.boardMem.board_14[5] ),
    .C1(_1473_),
    .B1(net971),
    .A1(\vga_tetris.boardMem.board_13[5] ),
    .Y(_1483_),
    .A2(net999));
 sg13g2_a22oi_1 _4422_ (.Y(_1484_),
    .B1(net980),
    .B2(\vga_tetris.boardMem.board_4[5] ),
    .A2(net981),
    .A1(\vga_tetris.boardMem.board_6[5] ));
 sg13g2_and4_1 _4423_ (.A(_1472_),
    .B(_1482_),
    .C(_1483_),
    .D(_1484_),
    .X(_1485_));
 sg13g2_nand4_1 _4424_ (.B(_1474_),
    .C(_1475_),
    .A(_1470_),
    .Y(_1486_),
    .D(_1480_));
 sg13g2_nand2_1 _4425_ (.Y(_1487_),
    .A(_1469_),
    .B(_1471_));
 sg13g2_a21o_1 _4426_ (.A2(net993),
    .A1(net995),
    .B1(_1478_),
    .X(_1488_));
 sg13g2_nand3_1 _4427_ (.B(_1477_),
    .C(_1481_),
    .A(_1476_),
    .Y(_1489_));
 sg13g2_nor4_1 _4428_ (.A(_1486_),
    .B(_1487_),
    .C(_1488_),
    .D(_1489_),
    .Y(_1490_));
 sg13g2_o21ai_1 _4429_ (.B1(net1068),
    .Y(_1491_),
    .A1(\vga_tetris.boardMem.board_0[5] ),
    .A2(net964));
 sg13g2_a21oi_2 _4430_ (.B1(_1491_),
    .Y(_1492_),
    .A2(_1490_),
    .A1(_1485_));
 sg13g2_nand3_1 _4431_ (.B(_1008_),
    .C(_1492_),
    .A(_0901_),
    .Y(_1493_));
 sg13g2_a221oi_1 _4432_ (.B2(_0902_),
    .C1(_1303_),
    .B1(_1423_),
    .A1(_1032_),
    .Y(_1494_),
    .A2(_1386_));
 sg13g2_o21ai_1 _4433_ (.B1(_1494_),
    .Y(_1495_),
    .A1(_0951_),
    .A2(_1366_));
 sg13g2_nand3_1 _4434_ (.B(_1444_),
    .C(_1493_),
    .A(_1346_),
    .Y(_1496_));
 sg13g2_o21ai_1 _4435_ (.B1(_1325_),
    .Y(_1497_),
    .A1(_0948_),
    .A2(_1407_));
 sg13g2_nor4_2 _4436_ (.A(_1468_),
    .B(_1495_),
    .C(_1496_),
    .Y(_1498_),
    .D(_1497_));
 sg13g2_a21o_2 _4437_ (.A2(_1498_),
    .A1(_1105_),
    .B1(_1282_),
    .X(uo_out[0]));
 sg13g2_nor3_2 _4438_ (.A(_1104_),
    .B(_1281_),
    .C(_1498_),
    .Y(uo_out[6]));
 sg13g2_nand2_1 _4439_ (.Y(_1499_),
    .A(_1097_),
    .B(uo_out[6]));
 sg13g2_nand2_2 _4440_ (.Y(uo_out[1]),
    .A(_1221_),
    .B(_1499_));
 sg13g2_nand3_1 _4441_ (.B(_1280_),
    .C(_1498_),
    .A(_1105_),
    .Y(_1500_));
 sg13g2_nand3_1 _4442_ (.B(_1499_),
    .C(_1500_),
    .A(_1221_),
    .Y(uo_out[5]));
 sg13g2_nor2b_2 _4443_ (.A(_1097_),
    .B_N(uo_out[6]),
    .Y(uo_out[2]));
 sg13g2_nand3_1 _4444_ (.B(\vga_tetris.vgaController.horizontalCounterQ[4] ),
    .C(net1678),
    .A(net1647),
    .Y(_1501_));
 sg13g2_nor3_1 _4445_ (.A(\vga_tetris.vgaController.horizontalCounterQ[5] ),
    .B(\vga_tetris.vgaController.horizontalCounterQ[4] ),
    .C(\vga_tetris.vgaController.horizontalCounterQ[6] ),
    .Y(_1502_));
 sg13g2_nor3_1 _4446_ (.A(\vga_tetris.vgaController.horizontalCounterQ[8] ),
    .B(_1100_),
    .C(_1502_),
    .Y(_1503_));
 sg13g2_nand2_1 _4447_ (.Y(vga_hs),
    .A(_1501_),
    .B(_1503_));
 sg13g2_nand3b_1 _4448_ (.B(net1582),
    .C(net1593),
    .Y(_1504_),
    .A_N(net1606));
 sg13g2_or4_1 _4449_ (.A(net1826),
    .B(net1591),
    .C(_1098_),
    .D(_1504_),
    .X(\vga_tetris._vgaController_io_vSync ));
 sg13g2_nor3_2 _4450_ (.A(net1205),
    .B(\vga_tetris.tetrisLogic.stateQ[2] ),
    .C(net1680),
    .Y(_1505_));
 sg13g2_nand2_1 _4451_ (.Y(_1506_),
    .A(_0721_),
    .B(_1505_));
 sg13g2_o21ai_1 _4452_ (.B1(_1506_),
    .Y(_1507_),
    .A1(_0708_),
    .A2(_0717_));
 sg13g2_and3_1 _4453_ (.X(_1508_),
    .A(_0796_),
    .B(_0810_),
    .C(net1140));
 sg13g2_and3_2 _4454_ (.X(_1509_),
    .A(_0749_),
    .B(_0762_),
    .C(_1508_));
 sg13g2_nand3_1 _4455_ (.B(_0762_),
    .C(_1508_),
    .A(_0749_),
    .Y(_1510_));
 sg13g2_or2_1 _4456_ (.X(_1511_),
    .B(_0724_),
    .A(_0717_));
 sg13g2_nand2_1 _4457_ (.Y(_1512_),
    .A(_1510_),
    .B(_1511_));
 sg13g2_nand4_1 _4458_ (.B(net1217),
    .C(\vga_tetris.tetrisLogic._checkMoveAllowed_io_checkDone ),
    .A(net1215),
    .Y(_1513_),
    .D(_0719_));
 sg13g2_inv_1 _4459_ (.Y(_1514_),
    .A(_1513_));
 sg13g2_nor2_1 _4460_ (.A(net1207),
    .B(net1212),
    .Y(_1515_));
 sg13g2_and3_1 _4461_ (.X(_1516_),
    .A(net1211),
    .B(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[0] ),
    .C(_1515_));
 sg13g2_nor2_2 _4462_ (.A(net1211),
    .B(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[0] ),
    .Y(_1517_));
 sg13g2_nor2_2 _4463_ (.A(net1212),
    .B(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[0] ),
    .Y(_1518_));
 sg13g2_and2_1 _4464_ (.A(_1515_),
    .B(_1517_),
    .X(_1519_));
 sg13g2_nor2_1 _4465_ (.A(net1211),
    .B(_1518_),
    .Y(_1520_));
 sg13g2_inv_1 _4466_ (.Y(_1521_),
    .A(_1520_));
 sg13g2_nor3_1 _4467_ (.A(_1516_),
    .B(_1519_),
    .C(_1520_),
    .Y(_1522_));
 sg13g2_nand2b_2 _4468_ (.Y(_1523_),
    .B(_0743_),
    .A_N(_0739_));
 sg13g2_nor3_1 _4469_ (.A(net1209),
    .B(_1522_),
    .C(_1523_),
    .Y(_1524_));
 sg13g2_or2_1 _4470_ (.X(_1525_),
    .B(_0743_),
    .A(_0739_));
 sg13g2_inv_1 _4471_ (.Y(_1526_),
    .A(_1525_));
 sg13g2_nand2_2 _4472_ (.Y(_1527_),
    .A(net1212),
    .B(_1517_));
 sg13g2_nand2_2 _4473_ (.Y(_1528_),
    .A(net1207),
    .B(_0654_));
 sg13g2_nor2_1 _4474_ (.A(_1527_),
    .B(_1528_),
    .Y(_1529_));
 sg13g2_nor2b_1 _4475_ (.A(_0743_),
    .B_N(_0739_),
    .Y(_1530_));
 sg13g2_nand2b_1 _4476_ (.Y(_1531_),
    .B(_0739_),
    .A_N(_0743_));
 sg13g2_nand2_1 _4477_ (.Y(_1532_),
    .A(net1211),
    .B(_1518_));
 sg13g2_nor2_1 _4478_ (.A(net1208),
    .B(net1210),
    .Y(_1533_));
 sg13g2_nand3_1 _4479_ (.B(_1518_),
    .C(_1533_),
    .A(net1211),
    .Y(_1534_));
 sg13g2_nor2b_2 _4480_ (.A(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[2] ),
    .B_N(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[0] ),
    .Y(_1535_));
 sg13g2_nand2_2 _4481_ (.Y(_1536_),
    .A(net1212),
    .B(_1535_));
 sg13g2_o21ai_1 _4482_ (.B1(_1534_),
    .Y(_1537_),
    .A1(_1528_),
    .A2(_1536_));
 sg13g2_a22oi_1 _4483_ (.Y(_1538_),
    .B1(_1530_),
    .B2(_1537_),
    .A2(_1529_),
    .A1(_1526_));
 sg13g2_nand2b_2 _4484_ (.Y(_1539_),
    .B(_1538_),
    .A_N(_1524_));
 sg13g2_nand2_2 _4485_ (.Y(_1540_),
    .A(_0897_),
    .B(_1467_));
 sg13g2_nand2b_2 _4486_ (.Y(_1541_),
    .B(net1204),
    .A_N(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[0] ));
 sg13g2_nand2_2 _4487_ (.Y(_1542_),
    .A(_0682_),
    .B(net1214));
 sg13g2_nor2_2 _4488_ (.A(_1541_),
    .B(_1542_),
    .Y(_1543_));
 sg13g2_nand2_1 _4489_ (.Y(_1544_),
    .A(_1540_),
    .B(_1543_));
 sg13g2_nand2_1 _4490_ (.Y(_1545_),
    .A(net1204),
    .B(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[0] ));
 sg13g2_nand2b_2 _4491_ (.Y(_1546_),
    .B(_1545_),
    .A_N(net1214));
 sg13g2_nor2_2 _4492_ (.A(net1204),
    .B(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[0] ),
    .Y(_1547_));
 sg13g2_nor2_1 _4493_ (.A(net1214),
    .B(net1204),
    .Y(_1548_));
 sg13g2_nand2b_2 _4494_ (.Y(_1549_),
    .B(_1547_),
    .A_N(net1214));
 sg13g2_nor2_2 _4495_ (.A(net1213),
    .B(_1549_),
    .Y(_1550_));
 sg13g2_a21o_2 _4496_ (.A2(_1546_),
    .A1(net1213),
    .B1(_1550_),
    .X(_1551_));
 sg13g2_a21o_2 _4497_ (.A2(_1006_),
    .A1(_1005_),
    .B1(_1492_),
    .X(_1552_));
 sg13g2_nand2_2 _4498_ (.Y(_1553_),
    .A(_1070_),
    .B(_1345_));
 sg13g2_nor2b_2 _4499_ (.A(_1542_),
    .B_N(_1547_),
    .Y(_1554_));
 sg13g2_a22oi_1 _4500_ (.Y(_1555_),
    .B1(_1553_),
    .B2(_1554_),
    .A2(_1552_),
    .A1(_1551_));
 sg13g2_nor3_2 _4501_ (.A(net1213),
    .B(net1214),
    .C(_1541_),
    .Y(_1556_));
 sg13g2_nand2_2 _4502_ (.Y(_1557_),
    .A(_1091_),
    .B(_1302_));
 sg13g2_nor3_2 _4503_ (.A(net1213),
    .B(net1214),
    .C(_1545_),
    .Y(_1558_));
 sg13g2_nand2_2 _4504_ (.Y(_1559_),
    .A(_0945_),
    .B(_1407_));
 sg13g2_nand2_1 _4505_ (.Y(_1560_),
    .A(_1558_),
    .B(_1559_));
 sg13g2_nor2_1 _4506_ (.A(_1030_),
    .B(_1386_),
    .Y(_1561_));
 sg13g2_inv_2 _4507_ (.Y(_1562_),
    .A(_1561_));
 sg13g2_nand2b_2 _4508_ (.Y(_1563_),
    .B(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[0] ),
    .A_N(net1204));
 sg13g2_nor3_2 _4509_ (.A(net1213),
    .B(net1214),
    .C(_1563_),
    .Y(_1564_));
 sg13g2_nand2_1 _4510_ (.Y(_1565_),
    .A(_1562_),
    .B(_1564_));
 sg13g2_nor2_2 _4511_ (.A(_1542_),
    .B(_1563_),
    .Y(_1566_));
 sg13g2_nand2_2 _4512_ (.Y(_1567_),
    .A(_0972_),
    .B(_1366_));
 sg13g2_a22oi_1 _4513_ (.Y(_1568_),
    .B1(_1566_),
    .B2(_1567_),
    .A2(_1557_),
    .A1(_1556_));
 sg13g2_inv_1 _4514_ (.Y(_1569_),
    .A(_1568_));
 sg13g2_nand4_1 _4515_ (.B(_1555_),
    .C(_1560_),
    .A(_1544_),
    .Y(_1570_),
    .D(_1565_));
 sg13g2_o21ai_1 _4516_ (.B1(_1539_),
    .Y(_1571_),
    .A1(_1569_),
    .A2(_1570_));
 sg13g2_o21ai_1 _4517_ (.B1(_1324_),
    .Y(_1572_),
    .A1(_0987_),
    .A2(_0988_));
 sg13g2_nand3_1 _4518_ (.B(net1204),
    .C(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[0] ),
    .A(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[2] ),
    .Y(_1573_));
 sg13g2_nor2_2 _4519_ (.A(net1213),
    .B(_1573_),
    .Y(_1574_));
 sg13g2_nand2_1 _4520_ (.Y(_1575_),
    .A(_0654_),
    .B(_1519_));
 sg13g2_nor2_1 _4521_ (.A(_1523_),
    .B(_1575_),
    .Y(_1576_));
 sg13g2_and2_1 _4522_ (.A(_1543_),
    .B(net1069),
    .X(_1577_));
 sg13g2_a21o_1 _4523_ (.A2(_1574_),
    .A1(net1064),
    .B1(_1577_),
    .X(_1578_));
 sg13g2_nor2_1 _4524_ (.A(\vga_tetris.tetrisLogic.checkMoveAllowed.checkIsRunningQ ),
    .B(\vga_tetris.tetrisLogic._checkMoveAllowed_io_checkDone ),
    .Y(_1579_));
 sg13g2_nor2_1 _4525_ (.A(net1204),
    .B(net1064),
    .Y(_1580_));
 sg13g2_nor3_1 _4526_ (.A(_0682_),
    .B(_1546_),
    .C(_1580_),
    .Y(_1581_));
 sg13g2_nor2_1 _4527_ (.A(_1579_),
    .B(_1581_),
    .Y(_1582_));
 sg13g2_nand2_2 _4528_ (.Y(_1583_),
    .A(net1211),
    .B(net1212));
 sg13g2_nor3_1 _4529_ (.A(net1207),
    .B(net1209),
    .C(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[0] ),
    .Y(_1584_));
 sg13g2_or2_1 _4530_ (.X(_1585_),
    .B(_1584_),
    .A(_1583_));
 sg13g2_nand3_1 _4531_ (.B(net1212),
    .C(_1517_),
    .A(net1209),
    .Y(_1586_));
 sg13g2_and2_1 _4532_ (.A(net1208),
    .B(net1210),
    .X(_1587_));
 sg13g2_nand2_1 _4533_ (.Y(_1588_),
    .A(net1207),
    .B(net1209));
 sg13g2_nand2b_2 _4534_ (.Y(_1589_),
    .B(_1535_),
    .A_N(net1212));
 sg13g2_nor2_1 _4535_ (.A(_1588_),
    .B(_1589_),
    .Y(_1590_));
 sg13g2_a21oi_1 _4536_ (.A1(net1209),
    .A2(_1519_),
    .Y(_1591_),
    .B1(_1590_));
 sg13g2_and2_1 _4537_ (.A(net1209),
    .B(_1516_),
    .X(_1592_));
 sg13g2_nand3_1 _4538_ (.B(_1586_),
    .C(_1591_),
    .A(_1583_),
    .Y(_1593_));
 sg13g2_nor2_1 _4539_ (.A(_1592_),
    .B(_1593_),
    .Y(_1594_));
 sg13g2_o21ai_1 _4540_ (.B1(_1594_),
    .Y(_1595_),
    .A1(net1207),
    .A2(_1536_));
 sg13g2_nand2_1 _4541_ (.Y(_1596_),
    .A(_1526_),
    .B(_1595_));
 sg13g2_o21ai_1 _4542_ (.B1(_1536_),
    .Y(_1597_),
    .A1(net1207),
    .A2(_1532_));
 sg13g2_nand2_1 _4543_ (.Y(_1598_),
    .A(_1588_),
    .B(_1597_));
 sg13g2_nand2_1 _4544_ (.Y(_1599_),
    .A(_1583_),
    .B(_1589_));
 sg13g2_nor2_1 _4545_ (.A(net1207),
    .B(_0654_),
    .Y(_1600_));
 sg13g2_nand2b_1 _4546_ (.Y(_1601_),
    .B(net1210),
    .A_N(net1208));
 sg13g2_o21ai_1 _4547_ (.B1(_1598_),
    .Y(_1602_),
    .A1(_1527_),
    .A2(_1600_));
 sg13g2_nor4_1 _4548_ (.A(_1519_),
    .B(_1592_),
    .C(_1599_),
    .D(_1602_),
    .Y(_1603_));
 sg13g2_o21ai_1 _4549_ (.B1(_1596_),
    .Y(_1604_),
    .A1(_1523_),
    .A2(_1603_));
 sg13g2_nand2b_1 _4550_ (.Y(_1605_),
    .B(_1527_),
    .A_N(_1516_));
 sg13g2_nand3_1 _4551_ (.B(_1601_),
    .C(_1605_),
    .A(_1528_),
    .Y(_1606_));
 sg13g2_nand2_1 _4552_ (.Y(_1607_),
    .A(net1210),
    .B(_1597_));
 sg13g2_and3_1 _4553_ (.X(_1608_),
    .A(_1591_),
    .B(_1606_),
    .C(_1607_));
 sg13g2_a22oi_1 _4554_ (.Y(_1609_),
    .B1(_1585_),
    .B2(_1604_),
    .A2(_1519_),
    .A1(net1209));
 sg13g2_o21ai_1 _4555_ (.B1(_1609_),
    .Y(_1610_),
    .A1(_1531_),
    .A2(_1608_));
 sg13g2_o21ai_1 _4556_ (.B1(_1586_),
    .Y(_1611_),
    .A1(_1536_),
    .A2(_1588_));
 sg13g2_a21oi_1 _4557_ (.A1(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[0] ),
    .A2(_1515_),
    .Y(_1612_),
    .B1(_1611_));
 sg13g2_a21oi_1 _4558_ (.A1(_1534_),
    .A2(_1612_),
    .Y(_1613_),
    .B1(_1531_));
 sg13g2_a22oi_1 _4559_ (.Y(_1614_),
    .B1(_1601_),
    .B2(_1528_),
    .A2(_1589_),
    .A1(_1586_));
 sg13g2_nand2_1 _4560_ (.Y(_1615_),
    .A(_1583_),
    .B(_1607_));
 sg13g2_o21ai_1 _4561_ (.B1(_1526_),
    .Y(_1616_),
    .A1(_1614_),
    .A2(_1615_));
 sg13g2_nor2_1 _4562_ (.A(_1527_),
    .B(_1587_),
    .Y(_1617_));
 sg13g2_or2_1 _4563_ (.X(_1618_),
    .B(_1517_),
    .A(net1212));
 sg13g2_nor2_1 _4564_ (.A(net1207),
    .B(_1618_),
    .Y(_1619_));
 sg13g2_a21oi_1 _4565_ (.A1(_1536_),
    .A2(_1575_),
    .Y(_1620_),
    .B1(_1600_));
 sg13g2_nor4_1 _4566_ (.A(_1599_),
    .B(_1617_),
    .C(_1619_),
    .D(_1620_),
    .Y(_1621_));
 sg13g2_o21ai_1 _4567_ (.B1(_1616_),
    .Y(_1622_),
    .A1(_1523_),
    .A2(_1621_));
 sg13g2_a21o_2 _4568_ (.A2(_1622_),
    .A1(_1585_),
    .B1(_1613_),
    .X(_1623_));
 sg13g2_nor3_1 _4569_ (.A(_1539_),
    .B(net1059),
    .C(net1062),
    .Y(_1624_));
 sg13g2_a21oi_1 _4570_ (.A1(_0764_),
    .A2(_1582_),
    .Y(_1625_),
    .B1(_1624_));
 sg13g2_a221oi_1 _4571_ (.B2(net1069),
    .C1(_1579_),
    .B1(_1574_),
    .A1(net1213),
    .Y(_1626_),
    .A2(_1546_));
 sg13g2_nand2b_1 _4572_ (.Y(_1627_),
    .B(_1626_),
    .A_N(_1625_));
 sg13g2_a21oi_1 _4573_ (.A1(_1572_),
    .A2(_1578_),
    .Y(_1628_),
    .B1(_1627_));
 sg13g2_nand2_1 _4574_ (.Y(_1629_),
    .A(_1551_),
    .B(_1562_));
 sg13g2_nand2_1 _4575_ (.Y(_1630_),
    .A(_1557_),
    .B(_1564_));
 sg13g2_nand2_1 _4576_ (.Y(_1631_),
    .A(_1556_),
    .B(_1559_));
 sg13g2_nand2_1 _4577_ (.Y(_1632_),
    .A(_1540_),
    .B(_1566_));
 sg13g2_nand4_1 _4578_ (.B(_1630_),
    .C(_1631_),
    .A(_1629_),
    .Y(_1633_),
    .D(_1632_));
 sg13g2_a221oi_1 _4579_ (.B2(_1554_),
    .C1(_1633_),
    .B1(_1567_),
    .A1(_1553_),
    .Y(_1634_),
    .A2(_1558_));
 sg13g2_nand2b_1 _4580_ (.Y(_1635_),
    .B(net1069),
    .A_N(_1634_));
 sg13g2_nor2_2 _4581_ (.A(_0682_),
    .B(_1549_),
    .Y(_1636_));
 sg13g2_a21o_1 _4582_ (.A2(_1048_),
    .A1(_1047_),
    .B1(_1443_),
    .X(_1637_));
 sg13g2_or3_1 _4583_ (.A(_0682_),
    .B(net1214),
    .C(_1563_),
    .X(_1638_));
 sg13g2_inv_2 _4584_ (.Y(_1639_),
    .A(_1638_));
 sg13g2_a21oi_1 _4585_ (.A1(_1551_),
    .A2(_1637_),
    .Y(_1640_),
    .B1(_1639_));
 sg13g2_a22oi_1 _4586_ (.Y(_1641_),
    .B1(_1566_),
    .B2(_1553_),
    .A2(_1562_),
    .A1(_1556_));
 sg13g2_a22oi_1 _4587_ (.Y(_1642_),
    .B1(_1567_),
    .B2(_1543_),
    .A2(_1558_),
    .A1(_1557_));
 sg13g2_a22oi_1 _4588_ (.Y(_1643_),
    .B1(_1564_),
    .B2(_1552_),
    .A2(_1559_),
    .A1(_1554_));
 sg13g2_a22oi_1 _4589_ (.Y(_1644_),
    .B1(_1636_),
    .B2(_1572_),
    .A2(_1574_),
    .A1(_1540_));
 sg13g2_nand2_1 _4590_ (.Y(_1645_),
    .A(_1641_),
    .B(_1644_));
 sg13g2_nand3_1 _4591_ (.B(_1642_),
    .C(_1643_),
    .A(_1640_),
    .Y(_1646_));
 sg13g2_o21ai_1 _4592_ (.B1(net1062),
    .Y(_1647_),
    .A1(_1645_),
    .A2(_1646_));
 sg13g2_o21ai_1 _4593_ (.B1(_0924_),
    .Y(_1648_),
    .A1(_1421_),
    .A2(_1422_));
 sg13g2_a22oi_1 _4594_ (.Y(_1649_),
    .B1(_1648_),
    .B2(_1551_),
    .A2(_1574_),
    .A1(_1567_));
 sg13g2_a22oi_1 _4595_ (.Y(_1650_),
    .B1(_1564_),
    .B2(_1637_),
    .A2(_1553_),
    .A1(_1543_));
 sg13g2_a22oi_1 _4596_ (.Y(_1651_),
    .B1(_1572_),
    .B2(_1639_),
    .A2(_1566_),
    .A1(_1559_));
 sg13g2_nand2_1 _4597_ (.Y(_1652_),
    .A(_1650_),
    .B(_1651_));
 sg13g2_a22oi_1 _4598_ (.Y(_1653_),
    .B1(_1636_),
    .B2(_1540_),
    .A2(_1557_),
    .A1(_1554_));
 sg13g2_a22oi_1 _4599_ (.Y(_1654_),
    .B1(_1558_),
    .B2(_1562_),
    .A2(_1556_),
    .A1(_1552_));
 sg13g2_nand3_1 _4600_ (.B(_1653_),
    .C(_1654_),
    .A(_1649_),
    .Y(_1655_));
 sg13g2_o21ai_1 _4601_ (.B1(net1059),
    .Y(_1656_),
    .A1(_1652_),
    .A2(_1655_));
 sg13g2_and2_1 _4602_ (.A(_1647_),
    .B(_1656_),
    .X(_1657_));
 sg13g2_nand4_1 _4603_ (.B(_1628_),
    .C(_1635_),
    .A(_1571_),
    .Y(_1658_),
    .D(_1657_));
 sg13g2_inv_1 _4604_ (.Y(_1659_),
    .A(_1658_));
 sg13g2_nand4_1 _4605_ (.B(\vga_tetris.tetrisLogic.shapeDropTimerQ[4] ),
    .C(\vga_tetris.tetrisLogic.shapeDropTimerQ[3] ),
    .A(\vga_tetris.tetrisLogic.shapeDropTimerQ[5] ),
    .Y(_1660_),
    .D(\vga_tetris.tetrisLogic.shapeDropTimerQ[2] ));
 sg13g2_o21ai_1 _4606_ (.B1(\vga_tetris.tetrisLogic.shapeDropTimerQ[2] ),
    .Y(_1661_),
    .A1(\vga_tetris.tetrisLogic.shapeDropTimerQ[1] ),
    .A2(\vga_tetris.tetrisLogic.shapeDropTimerQ[0] ));
 sg13g2_nor3_1 _4607_ (.A(\vga_tetris.tetrisLogic.shapeDropTimerQ[5] ),
    .B(\vga_tetris.tetrisLogic.shapeDropTimerQ[4] ),
    .C(\vga_tetris.tetrisLogic.shapeDropTimerQ[3] ),
    .Y(_1662_));
 sg13g2_a22oi_1 _4608_ (.Y(_1663_),
    .B1(_1661_),
    .B2(_1662_),
    .A2(_1660_),
    .A1(_0683_));
 sg13g2_nand2_1 _4609_ (.Y(_1664_),
    .A(_0722_),
    .B(_1663_));
 sg13g2_nand2_1 _4610_ (.Y(_1665_),
    .A(_1513_),
    .B(_1664_));
 sg13g2_and2_1 _4611_ (.A(_0721_),
    .B(_0728_),
    .X(_1666_));
 sg13g2_nand2_2 _4612_ (.Y(_1667_),
    .A(_0721_),
    .B(_0728_));
 sg13g2_nand2_1 _4613_ (.Y(_1668_),
    .A(\vga_tetris.startTetrisLogicQ ),
    .B(_1505_));
 sg13g2_and2_1 _4614_ (.A(net1215),
    .B(_1505_),
    .X(_1669_));
 sg13g2_nand2_1 _4615_ (.Y(_1670_),
    .A(net1199),
    .B(_1669_));
 sg13g2_inv_1 _4616_ (.Y(_1671_),
    .A(_1670_));
 sg13g2_nor2_1 _4617_ (.A(net1200),
    .B(_1670_),
    .Y(_1672_));
 sg13g2_or2_1 _4618_ (.X(_1673_),
    .B(_1670_),
    .A(net1200));
 sg13g2_o21ai_1 _4619_ (.B1(\vga_tetris._inputs_io_leftButtonActive ),
    .Y(_1674_),
    .A1(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[3] ),
    .A2(_1549_));
 sg13g2_nand2_1 _4620_ (.Y(_1675_),
    .A(\vga_tetris._inputs_io_rightButtonActive ),
    .B(_1638_));
 sg13g2_nand2b_2 _4621_ (.Y(_1676_),
    .B(_1674_),
    .A_N(_1675_));
 sg13g2_nor2_2 _4622_ (.A(net1848),
    .B(_1667_),
    .Y(_1677_));
 sg13g2_a22oi_1 _4623_ (.Y(_1678_),
    .B1(_1676_),
    .B2(_1677_),
    .A2(_1673_),
    .A1(_1667_));
 sg13g2_or2_1 _4624_ (.X(_1679_),
    .B(_1678_),
    .A(_1665_));
 sg13g2_o21ai_1 _4625_ (.B1(_1679_),
    .Y(_1680_),
    .A1(_1513_),
    .A2(net837));
 sg13g2_nor2_2 _4626_ (.A(_0707_),
    .B(_0724_),
    .Y(_1681_));
 sg13g2_or2_1 _4627_ (.X(_1682_),
    .B(_0724_),
    .A(_0707_));
 sg13g2_nand2_2 _4628_ (.Y(_1683_),
    .A(net1901),
    .B(_0734_));
 sg13g2_nor2_2 _4629_ (.A(net1217),
    .B(_1683_),
    .Y(_1684_));
 sg13g2_nand3_1 _4630_ (.B(net1794),
    .C(_0734_),
    .A(_0658_),
    .Y(_1685_));
 sg13g2_nor3_1 _4631_ (.A(_1509_),
    .B(_1681_),
    .C(_1684_),
    .Y(_1686_));
 sg13g2_a22oi_1 _4632_ (.Y(_1687_),
    .B1(_1680_),
    .B2(_1686_),
    .A2(_1512_),
    .A1(_1506_));
 sg13g2_nand3_1 _4633_ (.B(_0713_),
    .C(_0716_),
    .A(\vga_tetris.tetrisLogic._checkMoveAllowed_io_checkDone ),
    .Y(_1688_));
 sg13g2_nand4_1 _4634_ (.B(_1670_),
    .C(_1683_),
    .A(_1667_),
    .Y(_1689_),
    .D(_1688_));
 sg13g2_nand4_1 _4635_ (.B(_0658_),
    .C(\vga_tetris.tetrisLogic._checkMoveAllowed_io_checkDone ),
    .A(net1215),
    .Y(_1690_),
    .D(_0719_));
 sg13g2_nand2_1 _4636_ (.Y(_1691_),
    .A(_1682_),
    .B(_1690_));
 sg13g2_nor4_1 _4637_ (.A(_0722_),
    .B(_1514_),
    .C(_1689_),
    .D(_1691_),
    .Y(_1692_));
 sg13g2_nand2_1 _4638_ (.Y(_1693_),
    .A(\vga_tetris.tetrisLogic._checkMoveAllowed_io_checkDone ),
    .B(_0730_));
 sg13g2_nand3_1 _4639_ (.B(_0716_),
    .C(_0721_),
    .A(\vga_tetris.tetrisLogic._checkMoveAllowed_io_checkDone ),
    .Y(_1694_));
 sg13g2_nand3_1 _4640_ (.B(_0713_),
    .C(_1505_),
    .A(\vga_tetris.startTetrisLogicQ ),
    .Y(_1695_));
 sg13g2_nand2_2 _4641_ (.Y(_1696_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[1] ),
    .B(_0697_));
 sg13g2_or2_1 _4642_ (.X(_1697_),
    .B(_1696_),
    .A(_0710_));
 sg13g2_nand3_1 _4643_ (.B(_1695_),
    .C(_1697_),
    .A(_1694_),
    .Y(_1698_));
 sg13g2_a21oi_1 _4644_ (.A1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_done ),
    .A2(_0732_),
    .Y(_1699_),
    .B1(_1698_));
 sg13g2_and3_2 _4645_ (.X(_1700_),
    .A(_1692_),
    .B(_1693_),
    .C(_1699_));
 sg13g2_nand2_2 _4646_ (.Y(_1701_),
    .A(_1510_),
    .B(_1700_));
 sg13g2_inv_1 _4647_ (.Y(_1702_),
    .A(_1701_));
 sg13g2_o21ai_1 _4648_ (.B1(net1242),
    .Y(_1703_),
    .A1(net1217),
    .A2(_1701_));
 sg13g2_nand2_1 _4649_ (.Y(_1704_),
    .A(net1206),
    .B(_0726_));
 sg13g2_o21ai_1 _4650_ (.B1(_1511_),
    .Y(_1705_),
    .A1(net1216),
    .A2(_1704_));
 sg13g2_nor2_1 _4651_ (.A(_1687_),
    .B(_1703_),
    .Y(_0000_));
 sg13g2_and2_1 _4652_ (.A(_1674_),
    .B(_1677_),
    .X(_1706_));
 sg13g2_nand2b_1 _4653_ (.Y(_1707_),
    .B(\vga_tetris.tetrisLogic.gameOverResetHappenedQ ),
    .A_N(net1200));
 sg13g2_a21oi_1 _4654_ (.A1(\vga_tetris.tetrisLogic.gameOverResetHappenedQ ),
    .A2(_1672_),
    .Y(_1708_),
    .B1(_1666_));
 sg13g2_nand3_1 _4655_ (.B(_1690_),
    .C(_1697_),
    .A(_1685_),
    .Y(_1709_));
 sg13g2_nand2_2 _4656_ (.Y(_1710_),
    .A(_1688_),
    .B(_1694_));
 sg13g2_o21ai_1 _4657_ (.B1(_1664_),
    .Y(_1711_),
    .A1(_1706_),
    .A2(_1708_));
 sg13g2_nor3_1 _4658_ (.A(_1709_),
    .B(_1710_),
    .C(_1711_),
    .Y(_1712_));
 sg13g2_nor2_1 _4659_ (.A(net837),
    .B(_1694_),
    .Y(_1713_));
 sg13g2_nor2_1 _4660_ (.A(net837),
    .B(_1688_),
    .Y(_1714_));
 sg13g2_nand2_1 _4661_ (.Y(_1715_),
    .A(net837),
    .B(_1710_));
 sg13g2_nand2_2 _4662_ (.Y(_1716_),
    .A(_1659_),
    .B(_1710_));
 sg13g2_nand2b_1 _4663_ (.Y(_1717_),
    .B(_1716_),
    .A_N(_1712_));
 sg13g2_a21oi_1 _4664_ (.A1(net1216),
    .A2(_1702_),
    .Y(_1718_),
    .B1(net1138));
 sg13g2_a21oi_1 _4665_ (.A1(_1717_),
    .A2(_1718_),
    .Y(_0001_),
    .B1(net1228));
 sg13g2_or2_1 _4666_ (.X(_1719_),
    .B(net1138),
    .A(net1228));
 sg13g2_nand2_1 _4667_ (.Y(_1720_),
    .A(net1680),
    .B(_1692_));
 sg13g2_nand3b_1 _4668_ (.B(_1513_),
    .C(_1693_),
    .Y(_1721_),
    .A_N(_0722_));
 sg13g2_nor3_1 _4669_ (.A(_1706_),
    .B(_1709_),
    .C(_1721_),
    .Y(_1722_));
 sg13g2_a21oi_1 _4670_ (.A1(net1681),
    .A2(_1722_),
    .Y(_0002_),
    .B1(_1719_));
 sg13g2_nand2_1 _4671_ (.Y(_1723_),
    .A(net1242),
    .B(_1682_));
 sg13g2_nand2_1 _4672_ (.Y(_1724_),
    .A(net1243),
    .B(_1715_));
 sg13g2_nand2b_1 _4673_ (.Y(_1725_),
    .B(_1715_),
    .A_N(_1723_));
 sg13g2_nand2_2 _4674_ (.Y(_1726_),
    .A(\vga_tetris.tetrisLogic._checkMoveAllowed_io_checkDone ),
    .B(net837));
 sg13g2_nor3_2 _4675_ (.A(_0658_),
    .B(_0729_),
    .C(_1726_),
    .Y(_1727_));
 sg13g2_nor3_2 _4676_ (.A(_0714_),
    .B(_0720_),
    .C(_1726_),
    .Y(_1728_));
 sg13g2_xnor2_1 _4677_ (.Y(_1729_),
    .A(net1867),
    .B(_1547_));
 sg13g2_nand3b_1 _4678_ (.B(_1573_),
    .C(_1546_),
    .Y(_1730_),
    .A_N(_1676_));
 sg13g2_o21ai_1 _4679_ (.B1(_1730_),
    .Y(_1731_),
    .A1(_1674_),
    .A2(_1729_));
 sg13g2_nor4_2 _4680_ (.A(net1200),
    .B(net1720),
    .C(_0708_),
    .Y(_1732_),
    .D(_1668_));
 sg13g2_a21o_1 _4681_ (.A2(_1675_),
    .A1(_1674_),
    .B1(_1667_),
    .X(_1733_));
 sg13g2_nor2_1 _4682_ (.A(net1848),
    .B(_1733_),
    .Y(_1734_));
 sg13g2_nor2_1 _4683_ (.A(_1732_),
    .B(_1734_),
    .Y(_1735_));
 sg13g2_a22oi_1 _4684_ (.Y(_1736_),
    .B1(_1735_),
    .B2(net1867),
    .A2(_1731_),
    .A1(_1677_));
 sg13g2_nor2_1 _4685_ (.A(_1727_),
    .B(_1736_),
    .Y(_1737_));
 sg13g2_nand3_1 _4686_ (.B(_1573_),
    .C(_1727_),
    .A(_1546_),
    .Y(_1738_));
 sg13g2_nor2_1 _4687_ (.A(_1728_),
    .B(_1737_),
    .Y(_1739_));
 sg13g2_a221oi_1 _4688_ (.B2(_1739_),
    .C1(_1725_),
    .B1(_1738_),
    .A1(_1728_),
    .Y(_0003_),
    .A2(net1868));
 sg13g2_xnor2_1 _4689_ (.Y(_1740_),
    .A(_0682_),
    .B(_1573_));
 sg13g2_and2_1 _4690_ (.A(_1727_),
    .B(_1740_),
    .X(_1741_));
 sg13g2_and2_1 _4691_ (.A(net1884),
    .B(_1549_),
    .X(_1742_));
 sg13g2_nand2_1 _4692_ (.Y(_1743_),
    .A(\vga_tetris._inputs_io_leftButtonActive ),
    .B(_1742_));
 sg13g2_o21ai_1 _4693_ (.B1(_1743_),
    .Y(_1744_),
    .A1(_1676_),
    .A2(_1740_));
 sg13g2_a221oi_1 _4694_ (.B2(_1677_),
    .C1(_1727_),
    .B1(_1744_),
    .A1(net1884),
    .Y(_1745_),
    .A2(_1735_));
 sg13g2_or3_1 _4695_ (.A(_1728_),
    .B(_1741_),
    .C(_1745_),
    .X(_1746_));
 sg13g2_o21ai_1 _4696_ (.B1(_1728_),
    .Y(_1747_),
    .A1(_1550_),
    .A2(_1742_));
 sg13g2_a21oi_1 _4697_ (.A1(_1746_),
    .A2(net1885),
    .Y(_0004_),
    .B1(_1725_));
 sg13g2_and3_1 _4698_ (.X(_1748_),
    .A(net645),
    .B(net650),
    .C(net678));
 sg13g2_and2_1 _4699_ (.A(net1523),
    .B(_1748_),
    .X(_1749_));
 sg13g2_and2_1 _4700_ (.A(net1781),
    .B(_1749_),
    .X(_1750_));
 sg13g2_nor4_1 _4701_ (.A(net1897),
    .B(\vga_tetris.vgaController.horizontalCounterQ[7] ),
    .C(\vga_tetris.vgaController.horizontalCounterQ[6] ),
    .D(_1101_),
    .Y(_1751_));
 sg13g2_nand2_2 _4702_ (.Y(_1752_),
    .A(_1750_),
    .B(net1898));
 sg13g2_nand2_1 _4703_ (.Y(_1753_),
    .A(net1195),
    .B(_0875_));
 sg13g2_nor2_2 _4704_ (.A(_0876_),
    .B(_0950_),
    .Y(_1754_));
 sg13g2_inv_1 _4705_ (.Y(_1755_),
    .A(_1754_));
 sg13g2_nand2_1 _4706_ (.Y(_1756_),
    .A(net1191),
    .B(_1754_));
 sg13g2_nand2b_1 _4707_ (.Y(_1757_),
    .B(_1756_),
    .A_N(net1190));
 sg13g2_nor2_1 _4708_ (.A(net1579),
    .B(_1757_),
    .Y(_1758_));
 sg13g2_o21ai_1 _4709_ (.B1(net1887),
    .Y(_1759_),
    .A1(\vga_tetris._vgaController_io_pixelPosX[8] ),
    .A2(_1757_));
 sg13g2_nor2_2 _4710_ (.A(_1752_),
    .B(net1067),
    .Y(_1760_));
 sg13g2_nor2_2 _4711_ (.A(net1219),
    .B(_1760_),
    .Y(_1761_));
 sg13g2_o21ai_1 _4712_ (.B1(net1234),
    .Y(_1762_),
    .A1(_1752_),
    .A2(net1067));
 sg13g2_nor2_1 _4713_ (.A(net645),
    .B(net1063),
    .Y(_0005_));
 sg13g2_o21ai_1 _4714_ (.B1(_1761_),
    .Y(_1763_),
    .A1(net645),
    .A2(net650));
 sg13g2_a21oi_1 _4715_ (.A1(net645),
    .A2(net650),
    .Y(_0006_),
    .B1(_1763_));
 sg13g2_a21oi_1 _4716_ (.A1(net645),
    .A2(net650),
    .Y(_1764_),
    .B1(net678));
 sg13g2_nor3_1 _4717_ (.A(_1748_),
    .B(net1063),
    .C(_1764_),
    .Y(_0007_));
 sg13g2_nor2_1 _4718_ (.A(net1523),
    .B(_1748_),
    .Y(_1765_));
 sg13g2_nor3_1 _4719_ (.A(net1223),
    .B(_1749_),
    .C(_1765_),
    .Y(_0008_));
 sg13g2_o21ai_1 _4720_ (.B1(net1234),
    .Y(_1766_),
    .A1(net1781),
    .A2(_1749_));
 sg13g2_nor2_1 _4721_ (.A(_1750_),
    .B(_1766_),
    .Y(_0009_));
 sg13g2_and2_1 _4722_ (.A(net1647),
    .B(_1750_),
    .X(_1767_));
 sg13g2_nor2_1 _4723_ (.A(net1647),
    .B(_1750_),
    .Y(_1768_));
 sg13g2_nor3_1 _4724_ (.A(net1063),
    .B(_1767_),
    .C(net1648),
    .Y(_0010_));
 sg13g2_nor2_1 _4725_ (.A(net1678),
    .B(_1767_),
    .Y(_1769_));
 sg13g2_nor2b_1 _4726_ (.A(_1501_),
    .B_N(_1749_),
    .Y(_1770_));
 sg13g2_nor3_1 _4727_ (.A(net1063),
    .B(_1769_),
    .C(_1770_),
    .Y(_0011_));
 sg13g2_and2_1 _4728_ (.A(net1665),
    .B(_1770_),
    .X(_1771_));
 sg13g2_nor2_1 _4729_ (.A(net1665),
    .B(_1770_),
    .Y(_1772_));
 sg13g2_nor3_1 _4730_ (.A(_1762_),
    .B(_1771_),
    .C(net1666),
    .Y(_0012_));
 sg13g2_nand2_1 _4731_ (.Y(_1773_),
    .A(net1766),
    .B(_1771_));
 sg13g2_o21ai_1 _4732_ (.B1(_1761_),
    .Y(_1774_),
    .A1(net1766),
    .A2(_1771_));
 sg13g2_nor2b_1 _4733_ (.A(_1774_),
    .B_N(_1773_),
    .Y(_0013_));
 sg13g2_xor2_1 _4734_ (.B(_1773_),
    .A(net1751),
    .X(_1775_));
 sg13g2_nor2_1 _4735_ (.A(_1762_),
    .B(net1752),
    .Y(_0014_));
 sg13g2_nor4_1 _4736_ (.A(\vga_tetris.msTimer.msTimerQ[9] ),
    .B(\vga_tetris.msTimer.msTimerQ[11] ),
    .C(\vga_tetris.msTimer.msTimerQ[10] ),
    .D(\vga_tetris.msTimer.msTimerQ[12] ),
    .Y(_1776_));
 sg13g2_o21ai_1 _4737_ (.B1(\vga_tetris.msTimer.msTimerQ[5] ),
    .Y(_1777_),
    .A1(\vga_tetris.msTimer.msTimerQ[3] ),
    .A2(\vga_tetris.msTimer.msTimerQ[4] ));
 sg13g2_nor2b_1 _4738_ (.A(\vga_tetris.msTimer.msTimerQ[6] ),
    .B_N(_1777_),
    .Y(_1778_));
 sg13g2_nand2_1 _4739_ (.Y(_1779_),
    .A(net1653),
    .B(net1698));
 sg13g2_o21ai_1 _4740_ (.B1(_1776_),
    .Y(_1780_),
    .A1(_1778_),
    .A2(_1779_));
 sg13g2_nand3_1 _4741_ (.B(net1373),
    .C(_1780_),
    .A(net1353),
    .Y(_1781_));
 sg13g2_nand2_2 _4742_ (.Y(_1782_),
    .A(net1245),
    .B(_1781_));
 sg13g2_inv_2 _4743_ (.Y(_1783_),
    .A(net1135));
 sg13g2_nor2_1 _4744_ (.A(net646),
    .B(net1135),
    .Y(_0015_));
 sg13g2_xnor2_1 _4745_ (.Y(_1784_),
    .A(net1707),
    .B(net646));
 sg13g2_nor2_1 _4746_ (.A(net1135),
    .B(_1784_),
    .Y(_0016_));
 sg13g2_and3_1 _4747_ (.X(_1785_),
    .A(\vga_tetris.msTimer.msTimerQ[1] ),
    .B(net646),
    .C(net1384));
 sg13g2_a21oi_1 _4748_ (.A1(\vga_tetris.msTimer.msTimerQ[1] ),
    .A2(net646),
    .Y(_1786_),
    .B1(net1384));
 sg13g2_nor3_1 _4749_ (.A(net1135),
    .B(_1785_),
    .C(net1385),
    .Y(_0017_));
 sg13g2_and2_1 _4750_ (.A(net1634),
    .B(_1785_),
    .X(_1787_));
 sg13g2_nor2_1 _4751_ (.A(net1634),
    .B(_1785_),
    .Y(_1788_));
 sg13g2_nor3_1 _4752_ (.A(net1135),
    .B(_1787_),
    .C(net1635),
    .Y(_0018_));
 sg13g2_and2_1 _4753_ (.A(net1644),
    .B(_1787_),
    .X(_1789_));
 sg13g2_nor2_1 _4754_ (.A(net1644),
    .B(_1787_),
    .Y(_1790_));
 sg13g2_nor3_1 _4755_ (.A(_1782_),
    .B(_1789_),
    .C(net1645),
    .Y(_0019_));
 sg13g2_and2_1 _4756_ (.A(net1658),
    .B(_1789_),
    .X(_1791_));
 sg13g2_nor2_1 _4757_ (.A(net1658),
    .B(_1789_),
    .Y(_1792_));
 sg13g2_nor3_1 _4758_ (.A(_1782_),
    .B(_1791_),
    .C(_1792_),
    .Y(_0020_));
 sg13g2_and2_1 _4759_ (.A(net1697),
    .B(_1791_),
    .X(_1793_));
 sg13g2_nor2_1 _4760_ (.A(net1697),
    .B(_1791_),
    .Y(_1794_));
 sg13g2_nor3_1 _4761_ (.A(net1135),
    .B(_1793_),
    .C(_1794_),
    .Y(_0021_));
 sg13g2_nor2_1 _4762_ (.A(net1653),
    .B(_1793_),
    .Y(_1795_));
 sg13g2_and2_1 _4763_ (.A(net1653),
    .B(_1793_),
    .X(_1796_));
 sg13g2_nor3_1 _4764_ (.A(net1135),
    .B(net1654),
    .C(_1796_),
    .Y(_0022_));
 sg13g2_nor2b_1 _4765_ (.A(_1779_),
    .B_N(_1793_),
    .Y(_1797_));
 sg13g2_o21ai_1 _4766_ (.B1(_1783_),
    .Y(_1798_),
    .A1(net1698),
    .A2(_1796_));
 sg13g2_nor2_1 _4767_ (.A(_1797_),
    .B(_1798_),
    .Y(_0023_));
 sg13g2_and2_1 _4768_ (.A(net1744),
    .B(_1797_),
    .X(_1799_));
 sg13g2_o21ai_1 _4769_ (.B1(_1783_),
    .Y(_1800_),
    .A1(net1744),
    .A2(_1797_));
 sg13g2_nor2_1 _4770_ (.A(_1799_),
    .B(_1800_),
    .Y(_0024_));
 sg13g2_and2_1 _4771_ (.A(net1733),
    .B(_1799_),
    .X(_1801_));
 sg13g2_o21ai_1 _4772_ (.B1(_1783_),
    .Y(_1802_),
    .A1(net1733),
    .A2(_1799_));
 sg13g2_nor2_1 _4773_ (.A(_1801_),
    .B(net1734),
    .Y(_0025_));
 sg13g2_and2_1 _4774_ (.A(net1780),
    .B(_1801_),
    .X(_1803_));
 sg13g2_o21ai_1 _4775_ (.B1(_1783_),
    .Y(_1804_),
    .A1(net1780),
    .A2(_1801_));
 sg13g2_nor2_1 _4776_ (.A(_1803_),
    .B(_1804_),
    .Y(_0026_));
 sg13g2_and2_1 _4777_ (.A(net1730),
    .B(_1803_),
    .X(_1805_));
 sg13g2_o21ai_1 _4778_ (.B1(_1783_),
    .Y(_1806_),
    .A1(net1730),
    .A2(_1803_));
 sg13g2_nor2_1 _4779_ (.A(_1805_),
    .B(net1731),
    .Y(_0027_));
 sg13g2_o21ai_1 _4780_ (.B1(_1783_),
    .Y(_1807_),
    .A1(net1353),
    .A2(_1805_));
 sg13g2_a21oi_1 _4781_ (.A1(net1353),
    .A2(_1805_),
    .Y(_0028_),
    .B1(_1807_));
 sg13g2_a21oi_1 _4782_ (.A1(net1353),
    .A2(_1805_),
    .Y(_1808_),
    .B1(net1373));
 sg13g2_nor2_1 _4783_ (.A(net1135),
    .B(net1374),
    .Y(_0029_));
 sg13g2_nor2_1 _4784_ (.A(net837),
    .B(_1690_),
    .Y(_1809_));
 sg13g2_nor3_1 _4785_ (.A(net1142),
    .B(_1665_),
    .C(_1809_),
    .Y(_1810_));
 sg13g2_a21oi_2 _4786_ (.B1(_1509_),
    .Y(_1811_),
    .A2(_1810_),
    .A1(_1716_));
 sg13g2_a21oi_1 _4787_ (.A1(_0658_),
    .A2(_1669_),
    .Y(_1812_),
    .B1(\vga_tetris.tetrisLogic.gameOverResetHappenedQ ));
 sg13g2_nor2_1 _4788_ (.A(_1673_),
    .B(_1812_),
    .Y(_1813_));
 sg13g2_nor3_1 _4789_ (.A(_1681_),
    .B(_1710_),
    .C(_1813_),
    .Y(_1814_));
 sg13g2_and2_1 _4790_ (.A(_1810_),
    .B(_1814_),
    .X(_1815_));
 sg13g2_inv_1 _4791_ (.Y(_1816_),
    .A(_1815_));
 sg13g2_o21ai_1 _4792_ (.B1(net1236),
    .Y(_1817_),
    .A1(net1400),
    .A2(_1811_));
 sg13g2_a21oi_1 _4793_ (.A1(net1400),
    .A2(_1816_),
    .Y(_0030_),
    .B1(_1817_));
 sg13g2_and2_1 _4794_ (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[1] ),
    .B(_0725_),
    .X(_1818_));
 sg13g2_xor2_1 _4795_ (.B(_0725_),
    .A(net1792),
    .X(_1819_));
 sg13g2_xnor2_1 _4796_ (.Y(_1820_),
    .A(_0657_),
    .B(_1819_));
 sg13g2_a22oi_1 _4797_ (.Y(_1821_),
    .B1(_1820_),
    .B2(_1811_),
    .A2(_1815_),
    .A1(net1792));
 sg13g2_nor2_1 _4798_ (.A(net1218),
    .B(_1821_),
    .Y(_0031_));
 sg13g2_nand2_1 _4799_ (.Y(_1822_),
    .A(net1904),
    .B(_0725_));
 sg13g2_nor2_1 _4800_ (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[2] ),
    .B(_0725_),
    .Y(_1823_));
 sg13g2_xnor2_1 _4801_ (.Y(_1824_),
    .A(_0656_),
    .B(_0725_));
 sg13g2_a21oi_1 _4802_ (.A1(net1400),
    .A2(_1819_),
    .Y(_1825_),
    .B1(_1818_));
 sg13g2_xnor2_1 _4803_ (.Y(_1826_),
    .A(_1824_),
    .B(_1825_));
 sg13g2_a22oi_1 _4804_ (.Y(_1827_),
    .B1(_1826_),
    .B2(_1811_),
    .A2(_1815_),
    .A1(net1785));
 sg13g2_nor2_1 _4805_ (.A(net1220),
    .B(_1827_),
    .Y(_0032_));
 sg13g2_and2_1 _4806_ (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[3] ),
    .B(_0725_),
    .X(_1828_));
 sg13g2_xnor2_1 _4807_ (.Y(_1829_),
    .A(_0655_),
    .B(_0725_));
 sg13g2_o21ai_1 _4808_ (.B1(_1822_),
    .Y(_1830_),
    .A1(_1823_),
    .A2(_1825_));
 sg13g2_xor2_1 _4809_ (.B(_1830_),
    .A(_1829_),
    .X(_1831_));
 sg13g2_a22oi_1 _4810_ (.Y(_1832_),
    .B1(_1831_),
    .B2(_1811_),
    .A2(_1815_),
    .A1(net1743));
 sg13g2_nor2_1 _4811_ (.A(net1220),
    .B(_1832_),
    .Y(_0033_));
 sg13g2_a21oi_1 _4812_ (.A1(_1829_),
    .A2(_1830_),
    .Y(_1833_),
    .B1(_1828_));
 sg13g2_xor2_1 _4813_ (.B(_0725_),
    .A(net1762),
    .X(_1834_));
 sg13g2_xnor2_1 _4814_ (.Y(_1835_),
    .A(_1833_),
    .B(_1834_));
 sg13g2_a22oi_1 _4815_ (.Y(_1836_),
    .B1(_1835_),
    .B2(_1811_),
    .A2(_1815_),
    .A1(net1762));
 sg13g2_nor2_1 _4816_ (.A(net1220),
    .B(_1836_),
    .Y(_0034_));
 sg13g2_nor2_1 _4817_ (.A(_1681_),
    .B(_1732_),
    .Y(_1837_));
 sg13g2_a21oi_1 _4818_ (.A1(net1595),
    .A2(net1583),
    .Y(_1838_),
    .B1(_1682_));
 sg13g2_a22oi_1 _4819_ (.Y(_1839_),
    .B1(_1838_),
    .B2(net1614),
    .A2(_1837_),
    .A1(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[0] ));
 sg13g2_nor2_1 _4820_ (.A(_1724_),
    .B(net1615),
    .Y(_0035_));
 sg13g2_a22oi_1 _4821_ (.Y(_1840_),
    .B1(_1837_),
    .B2(net1642),
    .A2(_1681_),
    .A1(net1583));
 sg13g2_nor2_1 _4822_ (.A(_1724_),
    .B(net1643),
    .Y(_0036_));
 sg13g2_a22oi_1 _4823_ (.Y(_1841_),
    .B1(_1837_),
    .B2(net1211),
    .A2(_1681_),
    .A1(net1595));
 sg13g2_nor2_1 _4824_ (.A(_1724_),
    .B(net1737),
    .Y(_0037_));
 sg13g2_nor3_2 _4825_ (.A(net1217),
    .B(_0729_),
    .C(_1726_),
    .Y(_1842_));
 sg13g2_nor2_2 _4826_ (.A(_0679_),
    .B(_1667_),
    .Y(_1843_));
 sg13g2_nor2_1 _4827_ (.A(_1842_),
    .B(_1843_),
    .Y(_1844_));
 sg13g2_o21ai_1 _4828_ (.B1(_0654_),
    .Y(_1845_),
    .A1(net1208),
    .A2(_1583_));
 sg13g2_nor2b_1 _4829_ (.A(_1845_),
    .B_N(_1842_),
    .Y(_1846_));
 sg13g2_a21oi_1 _4830_ (.A1(_1533_),
    .A2(_1583_),
    .Y(_1847_),
    .B1(_1520_));
 sg13g2_nor2_1 _4831_ (.A(net1210),
    .B(_1847_),
    .Y(_1848_));
 sg13g2_a221oi_1 _4832_ (.B2(_1843_),
    .C1(_1846_),
    .B1(_1848_),
    .A1(net1210),
    .Y(_1849_),
    .A2(_1844_));
 sg13g2_nor2_1 _4833_ (.A(_1723_),
    .B(net1876),
    .Y(_0038_));
 sg13g2_a21oi_1 _4834_ (.A1(_1520_),
    .A2(_1533_),
    .Y(_1850_),
    .B1(_1587_));
 sg13g2_o21ai_1 _4835_ (.B1(_1850_),
    .Y(_1851_),
    .A1(_1521_),
    .A2(_1842_));
 sg13g2_a21o_1 _4836_ (.A2(_1850_),
    .A1(_1843_),
    .B1(_1842_),
    .X(_1852_));
 sg13g2_a22oi_1 _4837_ (.Y(_1853_),
    .B1(_1851_),
    .B2(_1852_),
    .A2(_1844_),
    .A1(net1208));
 sg13g2_nor2_1 _4838_ (.A(_1723_),
    .B(net1852),
    .Y(_0039_));
 sg13g2_a221oi_1 _4839_ (.B2(_1707_),
    .C1(_1666_),
    .B1(_1671_),
    .A1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_done ),
    .Y(_1854_),
    .A2(_0732_));
 sg13g2_nor3_1 _4840_ (.A(_0722_),
    .B(_1706_),
    .C(_1854_),
    .Y(_1855_));
 sg13g2_nor2b_1 _4841_ (.A(_1663_),
    .B_N(_0722_),
    .Y(_1856_));
 sg13g2_nor2_2 _4842_ (.A(_1514_),
    .B(_1856_),
    .Y(_1857_));
 sg13g2_nand3_1 _4843_ (.B(_1697_),
    .C(_1857_),
    .A(_1683_),
    .Y(_1858_));
 sg13g2_nor4_1 _4844_ (.A(_1700_),
    .B(_1713_),
    .C(_1855_),
    .D(_1858_),
    .Y(_1859_));
 sg13g2_nor2_1 _4845_ (.A(net1761),
    .B(_1701_),
    .Y(_1860_));
 sg13g2_nor3_1 _4846_ (.A(_1719_),
    .B(_1859_),
    .C(_1860_),
    .Y(_0040_));
 sg13g2_nor2_1 _4847_ (.A(net1205),
    .B(_1701_),
    .Y(_1861_));
 sg13g2_o21ai_1 _4848_ (.B1(_1671_),
    .Y(_1862_),
    .A1(net1200),
    .A2(\vga_tetris.tetrisLogic.gameOverResetHappenedQ ));
 sg13g2_a21oi_1 _4849_ (.A1(_1683_),
    .A2(_1862_),
    .Y(_1863_),
    .B1(_1684_));
 sg13g2_nor4_1 _4850_ (.A(_1681_),
    .B(_1700_),
    .C(_1710_),
    .D(_1863_),
    .Y(_1864_));
 sg13g2_nor3_1 _4851_ (.A(_1719_),
    .B(_1861_),
    .C(_1864_),
    .Y(_0041_));
 sg13g2_nor3_1 _4852_ (.A(_1727_),
    .B(_1728_),
    .C(_1734_),
    .Y(_1865_));
 sg13g2_nor2_1 _4853_ (.A(net1880),
    .B(_1732_),
    .Y(_1866_));
 sg13g2_nand2_1 _4854_ (.Y(_1867_),
    .A(_1682_),
    .B(_1715_));
 sg13g2_inv_1 _4855_ (.Y(_1868_),
    .A(_1867_));
 sg13g2_xnor2_1 _4856_ (.Y(_1869_),
    .A(_1865_),
    .B(_1866_));
 sg13g2_a21oi_1 _4857_ (.A1(_1868_),
    .A2(_1869_),
    .Y(_0042_),
    .B1(net1226));
 sg13g2_xnor2_1 _4858_ (.Y(_1870_),
    .A(net1204),
    .B(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[0] ));
 sg13g2_nor2_1 _4859_ (.A(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[1] ),
    .B(_1732_),
    .Y(_1871_));
 sg13g2_nor2_1 _4860_ (.A(_1734_),
    .B(_1871_),
    .Y(_1872_));
 sg13g2_nor2b_1 _4861_ (.A(_1870_),
    .B_N(_1676_),
    .Y(_1873_));
 sg13g2_a21oi_1 _4862_ (.A1(_1674_),
    .A2(_1870_),
    .Y(_1874_),
    .B1(_1873_));
 sg13g2_a21oi_1 _4863_ (.A1(_1677_),
    .A2(_1874_),
    .Y(_1875_),
    .B1(_1872_));
 sg13g2_nand2b_1 _4864_ (.Y(_1876_),
    .B(_1875_),
    .A_N(_1727_));
 sg13g2_a21oi_1 _4865_ (.A1(_1727_),
    .A2(_1870_),
    .Y(_1877_),
    .B1(_1728_));
 sg13g2_a221oi_1 _4866_ (.B2(_1877_),
    .C1(_1867_),
    .B1(_1876_),
    .A1(_1728_),
    .Y(_1878_),
    .A2(_1870_));
 sg13g2_nor2_1 _4867_ (.A(net1226),
    .B(_1878_),
    .Y(_0043_));
 sg13g2_a21o_2 _4868_ (.A2(net1138),
    .A1(_1663_),
    .B1(net1229),
    .X(_1879_));
 sg13g2_xnor2_1 _4869_ (.Y(_1880_),
    .A(net1709),
    .B(net1199));
 sg13g2_nor2_1 _4870_ (.A(_1879_),
    .B(net1710),
    .Y(_0044_));
 sg13g2_a21oi_1 _4871_ (.A1(\vga_tetris.tetrisLogic.shapeDropTimerQ[0] ),
    .A2(net1199),
    .Y(_1881_),
    .B1(net1533));
 sg13g2_and3_1 _4872_ (.X(_1882_),
    .A(net1533),
    .B(net1899),
    .C(\vga_tetris.startTetrisLogicQ ));
 sg13g2_nor3_1 _4873_ (.A(_1879_),
    .B(net1534),
    .C(_1882_),
    .Y(_0045_));
 sg13g2_nor2_1 _4874_ (.A(net1701),
    .B(_1882_),
    .Y(_1883_));
 sg13g2_and2_1 _4875_ (.A(net1701),
    .B(_1882_),
    .X(_1884_));
 sg13g2_nor3_1 _4876_ (.A(_1879_),
    .B(net1702),
    .C(_1884_),
    .Y(_0046_));
 sg13g2_nor2_1 _4877_ (.A(net1692),
    .B(_1884_),
    .Y(_1885_));
 sg13g2_and2_1 _4878_ (.A(net1692),
    .B(_1884_),
    .X(_1886_));
 sg13g2_nor3_1 _4879_ (.A(_1879_),
    .B(net1693),
    .C(_1886_),
    .Y(_0047_));
 sg13g2_nor2_1 _4880_ (.A(net1718),
    .B(_1886_),
    .Y(_1887_));
 sg13g2_and2_1 _4881_ (.A(net1718),
    .B(_1886_),
    .X(_1888_));
 sg13g2_nor3_1 _4882_ (.A(_1879_),
    .B(_1887_),
    .C(_1888_),
    .Y(_0048_));
 sg13g2_xnor2_1 _4883_ (.Y(_1889_),
    .A(net1738),
    .B(_1888_));
 sg13g2_nor2_1 _4884_ (.A(_1879_),
    .B(_1889_),
    .Y(_0049_));
 sg13g2_xnor2_1 _4885_ (.Y(_1890_),
    .A(net1561),
    .B(net1663));
 sg13g2_xnor2_1 _4886_ (.Y(_1891_),
    .A(net1626),
    .B(net1401));
 sg13g2_xnor2_1 _4887_ (.Y(_1892_),
    .A(_1890_),
    .B(_1891_));
 sg13g2_a21oi_1 _4888_ (.A1(net1614),
    .A2(net1156),
    .Y(_1893_),
    .B1(net1227));
 sg13g2_o21ai_1 _4889_ (.B1(_1893_),
    .Y(_0050_),
    .A1(net1157),
    .A2(_1892_));
 sg13g2_o21ai_1 _4890_ (.B1(net1245),
    .Y(_1894_),
    .A1(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[0] ),
    .A2(net1157));
 sg13g2_a21oi_1 _4891_ (.A1(_0652_),
    .A2(net1157),
    .Y(_0051_),
    .B1(_1894_));
 sg13g2_o21ai_1 _4892_ (.B1(net1243),
    .Y(_1895_),
    .A1(net1583),
    .A2(net1160));
 sg13g2_a21oi_1 _4893_ (.A1(_0651_),
    .A2(net1160),
    .Y(_0052_),
    .B1(_1895_));
 sg13g2_o21ai_1 _4894_ (.B1(net1243),
    .Y(_1896_),
    .A1(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[2] ),
    .A2(net1160));
 sg13g2_a21oi_1 _4895_ (.A1(_0650_),
    .A2(net1157),
    .Y(_0053_),
    .B1(_1896_));
 sg13g2_o21ai_1 _4896_ (.B1(net1243),
    .Y(_1897_),
    .A1(net1295),
    .A2(net1157));
 sg13g2_a21oi_1 _4897_ (.A1(_0649_),
    .A2(net1159),
    .Y(_0054_),
    .B1(_1897_));
 sg13g2_a21oi_1 _4898_ (.A1(net1483),
    .A2(net1158),
    .Y(_1898_),
    .B1(net1229));
 sg13g2_o21ai_1 _4899_ (.B1(_1898_),
    .Y(_0055_),
    .A1(_0649_),
    .A2(net1159));
 sg13g2_a21oi_1 _4900_ (.A1(net1382),
    .A2(net1158),
    .Y(_1899_),
    .B1(net1229));
 sg13g2_o21ai_1 _4901_ (.B1(_1899_),
    .Y(_0056_),
    .A1(_0648_),
    .A2(net1159));
 sg13g2_a21oi_1 _4902_ (.A1(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[7] ),
    .A2(net1159),
    .Y(_1900_),
    .B1(net1229));
 sg13g2_o21ai_1 _4903_ (.B1(_1900_),
    .Y(_0057_),
    .A1(_0647_),
    .A2(net1158));
 sg13g2_o21ai_1 _4904_ (.B1(net1243),
    .Y(_1901_),
    .A1(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[7] ),
    .A2(net1159));
 sg13g2_a21oi_1 _4905_ (.A1(_0646_),
    .A2(net1158),
    .Y(_0058_),
    .B1(_1901_));
 sg13g2_o21ai_1 _4906_ (.B1(net1243),
    .Y(_1902_),
    .A1(net1305),
    .A2(net1158));
 sg13g2_a21oi_1 _4907_ (.A1(_0645_),
    .A2(net1158),
    .Y(_0059_),
    .B1(_1902_));
 sg13g2_a21oi_1 _4908_ (.A1(net1401),
    .A2(net1158),
    .Y(_1903_),
    .B1(net1229));
 sg13g2_o21ai_1 _4909_ (.B1(_1903_),
    .Y(_0060_),
    .A1(_0645_),
    .A2(net1158));
 sg13g2_a21oi_1 _4910_ (.A1(net1628),
    .A2(net1160),
    .Y(_1904_),
    .B1(net1229));
 sg13g2_o21ai_1 _4911_ (.B1(_1904_),
    .Y(_0061_),
    .A1(_0644_),
    .A2(net1157));
 sg13g2_o21ai_1 _4912_ (.B1(net1245),
    .Y(_1905_),
    .A1(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[11] ),
    .A2(net1156));
 sg13g2_a21oi_1 _4913_ (.A1(_0643_),
    .A2(net1157),
    .Y(_0062_),
    .B1(_1905_));
 sg13g2_a21oi_1 _4914_ (.A1(net1663),
    .A2(net1156),
    .Y(_1906_),
    .B1(net1227));
 sg13g2_o21ai_1 _4915_ (.B1(_1906_),
    .Y(_0063_),
    .A1(_0643_),
    .A2(net1156));
 sg13g2_o21ai_1 _4916_ (.B1(net1245),
    .Y(_1907_),
    .A1(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[13] ),
    .A2(net1156));
 sg13g2_a21oi_1 _4917_ (.A1(_0642_),
    .A2(net1156),
    .Y(_0064_),
    .B1(_1907_));
 sg13g2_a21oi_1 _4918_ (.A1(net1561),
    .A2(net1156),
    .Y(_1908_),
    .B1(net1227));
 sg13g2_o21ai_1 _4919_ (.B1(_1908_),
    .Y(_0065_),
    .A1(_0642_),
    .A2(net1156));
 sg13g2_nor2_1 _4920_ (.A(net1776),
    .B(_0664_),
    .Y(_1909_));
 sg13g2_nand2b_1 _4921_ (.Y(_1910_),
    .B(net648),
    .A_N(\vga_tetris.tetrisLogic.addOrRemoveShape.stateQ[0] ));
 sg13g2_nand3_1 _4922_ (.B(\vga_tetris.tetrisLogic._addOrRemoveShape_io_rowIndex[0] ),
    .C(_1909_),
    .A(net1623),
    .Y(_1911_));
 sg13g2_nor2_1 _4923_ (.A(net1228),
    .B(net1624),
    .Y(_0066_));
 sg13g2_nor2b_1 _4924_ (.A(net1199),
    .B_N(_1857_),
    .Y(_1912_));
 sg13g2_nand2b_1 _4925_ (.Y(_1913_),
    .B(_1857_),
    .A_N(net1199));
 sg13g2_nand3_1 _4926_ (.B(net1164),
    .C(net1624),
    .A(net1242),
    .Y(_1914_));
 sg13g2_a21oi_1 _4927_ (.A1(_0664_),
    .A2(_1912_),
    .Y(_0067_),
    .B1(_1914_));
 sg13g2_nand2_1 _4928_ (.Y(_1915_),
    .A(\vga_tetris.tetrisLogic.addOrRemoveShape.stateQ[0] ),
    .B(net1239));
 sg13g2_a21oi_1 _4929_ (.A1(net648),
    .A2(_1913_),
    .Y(_0068_),
    .B1(_1915_));
 sg13g2_a21oi_1 _4930_ (.A1(net1623),
    .A2(net1711),
    .Y(_1916_),
    .B1(_1910_));
 sg13g2_o21ai_1 _4931_ (.B1(net1711),
    .Y(_1917_),
    .A1(_1913_),
    .A2(_1916_));
 sg13g2_o21ai_1 _4932_ (.B1(_1917_),
    .Y(_1918_),
    .A1(net1711),
    .A2(_1909_));
 sg13g2_nor2_1 _4933_ (.A(net1226),
    .B(net1777),
    .Y(_0069_));
 sg13g2_nor2_1 _4934_ (.A(net1623),
    .B(net1711),
    .Y(_1919_));
 sg13g2_a21oi_1 _4935_ (.A1(net1623),
    .A2(_1912_),
    .Y(_1920_),
    .B1(_1916_));
 sg13g2_nor3_1 _4936_ (.A(net1228),
    .B(_1919_),
    .C(_1920_),
    .Y(_0070_));
 sg13g2_nand2_1 _4937_ (.Y(_1921_),
    .A(net1387),
    .B(net1163));
 sg13g2_nand2_2 _4938_ (.Y(_1922_),
    .A(_1550_),
    .B(net1059));
 sg13g2_a21oi_1 _4939_ (.A1(net1211),
    .A2(_1518_),
    .Y(_1923_),
    .B1(\vga_tetris.tetrisLogic.addOrRemoveShape.clearingQ ));
 sg13g2_and2_1 _4940_ (.A(_1589_),
    .B(_1923_),
    .X(_1924_));
 sg13g2_nand2_2 _4941_ (.Y(_1925_),
    .A(_1589_),
    .B(_1923_));
 sg13g2_nor2_1 _4942_ (.A(_1922_),
    .B(_1924_),
    .Y(_1926_));
 sg13g2_a21oi_1 _4943_ (.A1(_0924_),
    .A2(_1922_),
    .Y(_1927_),
    .B1(_1926_));
 sg13g2_nand2b_1 _4944_ (.Y(_1928_),
    .B(_1927_),
    .A_N(net1163));
 sg13g2_a21oi_1 _4945_ (.A1(_1921_),
    .A2(_1928_),
    .Y(_0071_),
    .B1(net1225));
 sg13g2_nand2_1 _4946_ (.Y(_1929_),
    .A(net1347),
    .B(net1165));
 sg13g2_a21oi_2 _4947_ (.B1(\vga_tetris.tetrisLogic.addOrRemoveShape.clearingQ ),
    .Y(_1930_),
    .A2(_1618_),
    .A1(_1527_));
 sg13g2_inv_2 _4948_ (.Y(_1931_),
    .A(_1930_));
 sg13g2_mux2_1 _4949_ (.A0(_1930_),
    .A1(_1423_),
    .S(_1922_),
    .X(_1932_));
 sg13g2_nand2b_1 _4950_ (.Y(_1933_),
    .B(_1932_),
    .A_N(net1166));
 sg13g2_a21oi_1 _4951_ (.A1(_1929_),
    .A2(_1933_),
    .Y(_0072_),
    .B1(net1225));
 sg13g2_a22oi_1 _4952_ (.Y(_1934_),
    .B1(_1623_),
    .B2(_1550_),
    .A2(net1060),
    .A1(_1564_));
 sg13g2_nand2_1 _4953_ (.Y(_1935_),
    .A(_1049_),
    .B(_1934_));
 sg13g2_nor2_1 _4954_ (.A(_1924_),
    .B(_1934_),
    .Y(_1936_));
 sg13g2_nor2_1 _4955_ (.A(net1167),
    .B(_1936_),
    .Y(_1937_));
 sg13g2_a22oi_1 _4956_ (.Y(_1938_),
    .B1(_1935_),
    .B2(_1937_),
    .A2(net1167),
    .A1(net1719));
 sg13g2_nor2_1 _4957_ (.A(net1226),
    .B(_1938_),
    .Y(_0073_));
 sg13g2_nand2_1 _4958_ (.Y(_1939_),
    .A(net1379),
    .B(net1165));
 sg13g2_mux2_1 _4959_ (.A0(_1930_),
    .A1(_1443_),
    .S(_1934_),
    .X(_1940_));
 sg13g2_nand2b_1 _4960_ (.Y(_1941_),
    .B(_1940_),
    .A_N(net1167));
 sg13g2_a21oi_1 _4961_ (.A1(_1939_),
    .A2(_1941_),
    .Y(_0074_),
    .B1(net1226));
 sg13g2_nand2_1 _4962_ (.Y(_1942_),
    .A(_1556_),
    .B(net1059));
 sg13g2_a22oi_1 _4963_ (.Y(_1943_),
    .B1(_1564_),
    .B2(net1062),
    .A2(_1550_),
    .A1(net1064));
 sg13g2_nand2_2 _4964_ (.Y(_1944_),
    .A(_1942_),
    .B(_1943_));
 sg13g2_nand2b_1 _4965_ (.Y(_1945_),
    .B(_1007_),
    .A_N(_1944_));
 sg13g2_a21oi_1 _4966_ (.A1(_1925_),
    .A2(_1944_),
    .Y(_1946_),
    .B1(net1163));
 sg13g2_a22oi_1 _4967_ (.Y(_1947_),
    .B1(_1945_),
    .B2(_1946_),
    .A2(net1163),
    .A1(net1619));
 sg13g2_nor2_1 _4968_ (.A(net1225),
    .B(net1620),
    .Y(_0075_));
 sg13g2_nand2_1 _4969_ (.Y(_1948_),
    .A(net1376),
    .B(net1163));
 sg13g2_a21oi_1 _4970_ (.A1(_1931_),
    .A2(_1944_),
    .Y(_1949_),
    .B1(net1163));
 sg13g2_o21ai_1 _4971_ (.B1(_1949_),
    .Y(_1950_),
    .A1(_1492_),
    .A2(_1944_));
 sg13g2_a21oi_1 _4972_ (.A1(_1948_),
    .A2(_1950_),
    .Y(_0076_),
    .B1(net1218));
 sg13g2_nand2_1 _4973_ (.Y(_1951_),
    .A(net1388),
    .B(net1164));
 sg13g2_nand2_1 _4974_ (.Y(_1952_),
    .A(_1556_),
    .B(net1062));
 sg13g2_nand2_1 _4975_ (.Y(_1953_),
    .A(_1558_),
    .B(net1060));
 sg13g2_a22oi_1 _4976_ (.Y(_1954_),
    .B1(_1576_),
    .B2(_1550_),
    .A2(_1564_),
    .A1(_1539_));
 sg13g2_nand3_1 _4977_ (.B(_1953_),
    .C(_1954_),
    .A(_1952_),
    .Y(_1955_));
 sg13g2_a21oi_1 _4978_ (.A1(_1925_),
    .A2(_1955_),
    .Y(_1956_),
    .B1(net1164));
 sg13g2_o21ai_1 _4979_ (.B1(_1956_),
    .Y(_1957_),
    .A1(_1030_),
    .A2(_1955_));
 sg13g2_a21oi_1 _4980_ (.A1(net1389),
    .A2(_1957_),
    .Y(_0077_),
    .B1(net1218));
 sg13g2_nand2_1 _4981_ (.Y(_1958_),
    .A(net1367),
    .B(net1164));
 sg13g2_a21oi_1 _4982_ (.A1(_1931_),
    .A2(_1955_),
    .Y(_1959_),
    .B1(net1164));
 sg13g2_o21ai_1 _4983_ (.B1(_1959_),
    .Y(_1960_),
    .A1(_1386_),
    .A2(_1955_));
 sg13g2_a21oi_1 _4984_ (.A1(net1368),
    .A2(_1960_),
    .Y(_0078_),
    .B1(net1218));
 sg13g2_nand2_1 _4985_ (.Y(_1961_),
    .A(net1506),
    .B(net1166));
 sg13g2_a22oi_1 _4986_ (.Y(_1962_),
    .B1(_1564_),
    .B2(net1069),
    .A2(_1556_),
    .A1(net1064));
 sg13g2_a22oi_1 _4987_ (.Y(_1963_),
    .B1(net1062),
    .B2(_1558_),
    .A2(net1059),
    .A1(_1554_));
 sg13g2_nand2_1 _4988_ (.Y(_1964_),
    .A(_1962_),
    .B(_1963_));
 sg13g2_nand2b_1 _4989_ (.Y(_1965_),
    .B(_1091_),
    .A_N(_1964_));
 sg13g2_a21oi_1 _4990_ (.A1(_1925_),
    .A2(_1964_),
    .Y(_1966_),
    .B1(net1166));
 sg13g2_nand2_1 _4991_ (.Y(_1967_),
    .A(_1965_),
    .B(_1966_));
 sg13g2_a21oi_1 _4992_ (.A1(_1961_),
    .A2(_1967_),
    .Y(_0079_),
    .B1(net1225));
 sg13g2_nand2b_1 _4993_ (.Y(_1968_),
    .B(_1302_),
    .A_N(_1964_));
 sg13g2_a21oi_1 _4994_ (.A1(_1931_),
    .A2(_1964_),
    .Y(_1969_),
    .B1(net1166));
 sg13g2_a22oi_1 _4995_ (.Y(_1970_),
    .B1(_1968_),
    .B2(_1969_),
    .A2(net1166),
    .A1(net1629));
 sg13g2_nor2_1 _4996_ (.A(net1225),
    .B(_1970_),
    .Y(_0080_));
 sg13g2_nand2_1 _4997_ (.Y(_1971_),
    .A(net1518),
    .B(net1161));
 sg13g2_a22oi_1 _4998_ (.Y(_1972_),
    .B1(net1069),
    .B2(_1556_),
    .A2(_1558_),
    .A1(net1064));
 sg13g2_a21oi_2 _4999_ (.B1(_1548_),
    .Y(_1973_),
    .A2(_1563_),
    .A1(_0682_));
 sg13g2_a22oi_1 _5000_ (.Y(_1974_),
    .B1(_1973_),
    .B2(net1059),
    .A2(net1062),
    .A1(_1554_));
 sg13g2_and2_1 _5001_ (.A(_1972_),
    .B(_1974_),
    .X(_1975_));
 sg13g2_nor2_1 _5002_ (.A(_1924_),
    .B(_1975_),
    .Y(_1976_));
 sg13g2_a21oi_1 _5003_ (.A1(_0945_),
    .A2(_1975_),
    .Y(_1977_),
    .B1(_1976_));
 sg13g2_nand2b_1 _5004_ (.Y(_1978_),
    .B(_1977_),
    .A_N(net1161));
 sg13g2_a21oi_1 _5005_ (.A1(_1971_),
    .A2(_1978_),
    .Y(_0081_),
    .B1(net1218));
 sg13g2_nand2_1 _5006_ (.Y(_1979_),
    .A(net1351),
    .B(net1161));
 sg13g2_nor2_1 _5007_ (.A(_1930_),
    .B(_1975_),
    .Y(_1980_));
 sg13g2_a21oi_1 _5008_ (.A1(_1407_),
    .A2(_1975_),
    .Y(_1981_),
    .B1(_1980_));
 sg13g2_nand2b_1 _5009_ (.Y(_1982_),
    .B(_1981_),
    .A_N(net1161));
 sg13g2_a21oi_1 _5010_ (.A1(_1979_),
    .A2(_1982_),
    .Y(_0082_),
    .B1(net1224));
 sg13g2_nand2_1 _5011_ (.Y(_1983_),
    .A(net1370),
    .B(net1165));
 sg13g2_a22oi_1 _5012_ (.Y(_1984_),
    .B1(_1558_),
    .B2(net1069),
    .A2(_1554_),
    .A1(net1064));
 sg13g2_a22oi_1 _5013_ (.Y(_1985_),
    .B1(_1623_),
    .B2(_1973_),
    .A2(net1060),
    .A1(_1543_));
 sg13g2_and2_1 _5014_ (.A(_1984_),
    .B(_1985_),
    .X(_1986_));
 sg13g2_nor2_1 _5015_ (.A(_1924_),
    .B(_1986_),
    .Y(_1987_));
 sg13g2_a21oi_1 _5016_ (.A1(_1070_),
    .A2(_1986_),
    .Y(_1988_),
    .B1(_1987_));
 sg13g2_nand2b_1 _5017_ (.Y(_1989_),
    .B(_1988_),
    .A_N(net1165));
 sg13g2_a21oi_1 _5018_ (.A1(_1983_),
    .A2(_1989_),
    .Y(_0083_),
    .B1(net1225));
 sg13g2_nand2_1 _5019_ (.Y(_1990_),
    .A(net1345),
    .B(net1165));
 sg13g2_nor2_1 _5020_ (.A(_1930_),
    .B(_1986_),
    .Y(_1991_));
 sg13g2_a21oi_1 _5021_ (.A1(_1345_),
    .A2(_1986_),
    .Y(_1992_),
    .B1(_1991_));
 sg13g2_nand2b_1 _5022_ (.Y(_1993_),
    .B(_1992_),
    .A_N(net1165));
 sg13g2_a21oi_1 _5023_ (.A1(_1990_),
    .A2(_1993_),
    .Y(_0084_),
    .B1(net1225));
 sg13g2_a22oi_1 _5024_ (.Y(_1994_),
    .B1(_1973_),
    .B2(net1064),
    .A2(net1059),
    .A1(_1574_));
 sg13g2_a22oi_1 _5025_ (.Y(_1995_),
    .B1(net1062),
    .B2(_1543_),
    .A2(net1069),
    .A1(_1554_));
 sg13g2_and2_1 _5026_ (.A(_1994_),
    .B(_1995_),
    .X(_1996_));
 sg13g2_nand2_1 _5027_ (.Y(_1997_),
    .A(_0972_),
    .B(_1996_));
 sg13g2_nor2_1 _5028_ (.A(_1924_),
    .B(_1996_),
    .Y(_1998_));
 sg13g2_nor2_1 _5029_ (.A(net1161),
    .B(_1998_),
    .Y(_1999_));
 sg13g2_a22oi_1 _5030_ (.Y(_2000_),
    .B1(_1997_),
    .B2(_1999_),
    .A2(net1161),
    .A1(net1625));
 sg13g2_nor2_1 _5031_ (.A(net1224),
    .B(_2000_),
    .Y(_0085_));
 sg13g2_nand2_1 _5032_ (.Y(_2001_),
    .A(_1366_),
    .B(_1996_));
 sg13g2_nor2_1 _5033_ (.A(_1930_),
    .B(_1996_),
    .Y(_2002_));
 sg13g2_nor2_1 _5034_ (.A(net1161),
    .B(_2002_),
    .Y(_2003_));
 sg13g2_a22oi_1 _5035_ (.Y(_2004_),
    .B1(_2001_),
    .B2(_2003_),
    .A2(net1161),
    .A1(net1608));
 sg13g2_nor2_1 _5036_ (.A(net1224),
    .B(net1609),
    .Y(_0086_));
 sg13g2_nand2_1 _5037_ (.Y(_2005_),
    .A(net1778),
    .B(net1162));
 sg13g2_nand2_1 _5038_ (.Y(_2006_),
    .A(_1574_),
    .B(net1062));
 sg13g2_nand2_1 _5039_ (.Y(_2007_),
    .A(net1059),
    .B(_1636_));
 sg13g2_a22oi_1 _5040_ (.Y(_2008_),
    .B1(net1069),
    .B2(_1973_),
    .A2(_1543_),
    .A1(net1064));
 sg13g2_nand3_1 _5041_ (.B(_2007_),
    .C(_2008_),
    .A(_2006_),
    .Y(_2009_));
 sg13g2_nand2_1 _5042_ (.Y(_2010_),
    .A(_1925_),
    .B(_2009_));
 sg13g2_o21ai_1 _5043_ (.B1(_2010_),
    .Y(_2011_),
    .A1(_0896_),
    .A2(_2009_));
 sg13g2_o21ai_1 _5044_ (.B1(_2005_),
    .Y(_2012_),
    .A1(net1162),
    .A2(_2011_));
 sg13g2_and2_1 _5045_ (.A(net1231),
    .B(_2012_),
    .X(_0087_));
 sg13g2_nand2_1 _5046_ (.Y(_2013_),
    .A(net1784),
    .B(net1162));
 sg13g2_nand2_1 _5047_ (.Y(_2014_),
    .A(_1931_),
    .B(_2009_));
 sg13g2_o21ai_1 _5048_ (.B1(_2014_),
    .Y(_2015_),
    .A1(_1466_),
    .A2(_2009_));
 sg13g2_o21ai_1 _5049_ (.B1(_2013_),
    .Y(_2016_),
    .A1(net1162),
    .A2(_2015_));
 sg13g2_and2_1 _5050_ (.A(net1231),
    .B(_2016_),
    .X(_0088_));
 sg13g2_nand2_1 _5051_ (.Y(_2017_),
    .A(net1377),
    .B(net1165));
 sg13g2_a221oi_1 _5052_ (.B2(net1060),
    .C1(_1578_),
    .B1(_1639_),
    .A1(_1623_),
    .Y(_2018_),
    .A2(_1636_));
 sg13g2_mux2_1 _5053_ (.A0(_1924_),
    .A1(_0989_),
    .S(_2018_),
    .X(_2019_));
 sg13g2_nand2b_1 _5054_ (.Y(_2020_),
    .B(_2019_),
    .A_N(net1165));
 sg13g2_a21oi_1 _5055_ (.A1(_2017_),
    .A2(_2020_),
    .Y(_0089_),
    .B1(net1226));
 sg13g2_nand2_1 _5056_ (.Y(_2021_),
    .A(_1324_),
    .B(_2018_));
 sg13g2_nor2_1 _5057_ (.A(_1930_),
    .B(_2018_),
    .Y(_2022_));
 sg13g2_nor2_1 _5058_ (.A(net1166),
    .B(_2022_),
    .Y(_2023_));
 sg13g2_a22oi_1 _5059_ (.Y(_2024_),
    .B1(_2021_),
    .B2(_2023_),
    .A2(net1166),
    .A1(net1621));
 sg13g2_nor2_1 _5060_ (.A(net1225),
    .B(net1622),
    .Y(_0090_));
 sg13g2_o21ai_1 _5061_ (.B1(net1200),
    .Y(_2025_),
    .A1(net1790),
    .A2(_0632_));
 sg13g2_nand3_1 _5062_ (.B(_1511_),
    .C(_2025_),
    .A(net1200),
    .Y(_2026_));
 sg13g2_nand2_1 _5063_ (.Y(_2027_),
    .A(net1720),
    .B(_1673_));
 sg13g2_a21oi_1 _5064_ (.A1(_2026_),
    .A2(_2027_),
    .Y(_0091_),
    .B1(net1228));
 sg13g2_nand2_1 _5065_ (.Y(_2028_),
    .A(_1664_),
    .B(_1733_));
 sg13g2_nor4_1 _5066_ (.A(_1691_),
    .B(_1714_),
    .C(_1843_),
    .D(_2028_),
    .Y(_2029_));
 sg13g2_a21oi_1 _5067_ (.A1(net1380),
    .A2(net1287),
    .Y(_2030_),
    .B1(net837));
 sg13g2_nand2_1 _5068_ (.Y(_2031_),
    .A(net1562),
    .B(net1242));
 sg13g2_nand2_1 _5069_ (.Y(_2032_),
    .A(net1562),
    .B(_2030_));
 sg13g2_a21oi_1 _5070_ (.A1(_2029_),
    .A2(_2032_),
    .Y(_0092_),
    .B1(net1228));
 sg13g2_nor2b_1 _5071_ (.A(net1794),
    .B_N(\vga_tetris.tetrisLogic.addOrRemoveShape.clearingQ ),
    .Y(_2033_));
 sg13g2_a21oi_1 _5072_ (.A1(_1857_),
    .A2(net1795),
    .Y(_2034_),
    .B1(net1199));
 sg13g2_nor2_1 _5073_ (.A(net1228),
    .B(_2034_),
    .Y(_0093_));
 sg13g2_a21o_1 _5074_ (.A2(net837),
    .A1(_0641_),
    .B1(_2031_),
    .X(_2035_));
 sg13g2_a21oi_1 _5075_ (.A1(net1287),
    .A2(_2030_),
    .Y(_0094_),
    .B1(_2035_));
 sg13g2_a21oi_1 _5076_ (.A1(net1287),
    .A2(_1659_),
    .Y(_2036_),
    .B1(net1380));
 sg13g2_nor2_1 _5077_ (.A(_2031_),
    .B(_2036_),
    .Y(_0095_));
 sg13g2_nand2_1 _5078_ (.Y(_2037_),
    .A(net1202),
    .B(_1696_));
 sg13g2_a21oi_1 _5079_ (.A1(_1685_),
    .A2(net1864),
    .Y(_0096_),
    .B1(net1220));
 sg13g2_nand4_1 _5080_ (.B(_1572_),
    .C(_1637_),
    .A(_1557_),
    .Y(_2038_),
    .D(_1648_));
 sg13g2_a22oi_1 _5081_ (.Y(_2039_),
    .B1(_1387_),
    .B2(_1031_),
    .A2(_1345_),
    .A1(_1070_));
 sg13g2_a22oi_1 _5082_ (.Y(_2040_),
    .B1(_1467_),
    .B2(_0897_),
    .A2(_1407_),
    .A1(_0945_));
 sg13g2_nand4_1 _5083_ (.B(_1567_),
    .C(_2039_),
    .A(_1552_),
    .Y(_2041_),
    .D(_2040_));
 sg13g2_nor2_1 _5084_ (.A(_2038_),
    .B(_2041_),
    .Y(_2042_));
 sg13g2_and2_1 _5085_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[0] ),
    .B(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[1] ),
    .X(_2043_));
 sg13g2_and4_1 _5086_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[4] ),
    .B(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[3] ),
    .C(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[2] ),
    .D(_2043_),
    .X(_2044_));
 sg13g2_inv_1 _5087_ (.Y(_2045_),
    .A(_2044_));
 sg13g2_nor2_1 _5088_ (.A(_0885_),
    .B(_2045_),
    .Y(_2046_));
 sg13g2_and2_1 _5089_ (.A(_2042_),
    .B(_2046_),
    .X(_2047_));
 sg13g2_nand2b_1 _5090_ (.Y(_2048_),
    .B(_2047_),
    .A_N(net1201));
 sg13g2_nor3_1 _5091_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[1] ),
    .B(net1201),
    .C(net1763),
    .Y(_2049_));
 sg13g2_nand2b_2 _5092_ (.Y(_2050_),
    .B(_2049_),
    .A_N(net1745));
 sg13g2_nor2_2 _5093_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[4] ),
    .B(_2050_),
    .Y(_2051_));
 sg13g2_inv_1 _5094_ (.Y(_2052_),
    .A(_2051_));
 sg13g2_nor2_1 _5095_ (.A(_0703_),
    .B(_2051_),
    .Y(_2053_));
 sg13g2_nand2_1 _5096_ (.Y(_2054_),
    .A(net1168),
    .B(_2052_));
 sg13g2_nor2_2 _5097_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.internalStartTriggerQ ),
    .B(_1684_),
    .Y(_2055_));
 sg13g2_nand2b_2 _5098_ (.Y(_2056_),
    .B(_1685_),
    .A_N(\vga_tetris.tetrisLogic.shiftTheBoard.internalStartTriggerQ ));
 sg13g2_a21oi_1 _5099_ (.A1(_0661_),
    .A2(_2055_),
    .Y(_2057_),
    .B1(net1137));
 sg13g2_a221oi_1 _5100_ (.B2(_2048_),
    .C1(net1176),
    .B1(_2057_),
    .A1(_0661_),
    .Y(_2058_),
    .A2(net1137));
 sg13g2_nor3_1 _5101_ (.A(net1203),
    .B(net1810),
    .C(net1136),
    .Y(_2059_));
 sg13g2_nor3_1 _5102_ (.A(net1221),
    .B(_2058_),
    .C(net1811),
    .Y(_0097_));
 sg13g2_nor2_1 _5103_ (.A(net1871),
    .B(net1136),
    .Y(_2060_));
 sg13g2_nor2_1 _5104_ (.A(net1203),
    .B(_2060_),
    .Y(_2061_));
 sg13g2_a21oi_1 _5105_ (.A1(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[1] ),
    .A2(_2047_),
    .Y(_2062_),
    .B1(net1137));
 sg13g2_o21ai_1 _5106_ (.B1(_2062_),
    .Y(_2063_),
    .A1(_2047_),
    .A2(_2060_));
 sg13g2_nor2_1 _5107_ (.A(net1810),
    .B(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[1] ),
    .Y(_2064_));
 sg13g2_nor2_1 _5108_ (.A(_2043_),
    .B(_2064_),
    .Y(_2065_));
 sg13g2_a21oi_1 _5109_ (.A1(net1137),
    .A2(_2065_),
    .Y(_2066_),
    .B1(net1176));
 sg13g2_a21oi_1 _5110_ (.A1(_2063_),
    .A2(_2066_),
    .Y(_2067_),
    .B1(_2061_));
 sg13g2_nor2_1 _5111_ (.A(net1221),
    .B(net1872),
    .Y(_0098_));
 sg13g2_or2_1 _5112_ (.X(_2068_),
    .B(net1136),
    .A(net1888));
 sg13g2_nand2_1 _5113_ (.Y(_2069_),
    .A(net1176),
    .B(_2068_));
 sg13g2_mux2_1 _5114_ (.A0(_2068_),
    .A1(net1763),
    .S(_2047_),
    .X(_2070_));
 sg13g2_nor3_1 _5115_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[0] ),
    .B(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[2] ),
    .C(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[1] ),
    .Y(_2071_));
 sg13g2_xnor2_1 _5116_ (.Y(_2072_),
    .A(net1888),
    .B(_2064_));
 sg13g2_a21oi_1 _5117_ (.A1(net1137),
    .A2(_2072_),
    .Y(_2073_),
    .B1(net1176));
 sg13g2_o21ai_1 _5118_ (.B1(_2073_),
    .Y(_2074_),
    .A1(net1137),
    .A2(_2070_));
 sg13g2_a21oi_1 _5119_ (.A1(_2069_),
    .A2(_2074_),
    .Y(_0099_),
    .B1(net1222));
 sg13g2_nor2_1 _5120_ (.A(net1883),
    .B(net1136),
    .Y(_2075_));
 sg13g2_nor2_1 _5121_ (.A(net1203),
    .B(_2075_),
    .Y(_2076_));
 sg13g2_a21oi_1 _5122_ (.A1(net1745),
    .A2(_2047_),
    .Y(_2077_),
    .B1(net1137));
 sg13g2_o21ai_1 _5123_ (.B1(_2077_),
    .Y(_2078_),
    .A1(_2047_),
    .A2(_2075_));
 sg13g2_nor2b_1 _5124_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[3] ),
    .B_N(_2071_),
    .Y(_2079_));
 sg13g2_xnor2_1 _5125_ (.Y(_2080_),
    .A(net1883),
    .B(_2071_));
 sg13g2_a21oi_1 _5126_ (.A1(_2053_),
    .A2(_2080_),
    .Y(_2081_),
    .B1(net1176));
 sg13g2_a21oi_1 _5127_ (.A1(_2078_),
    .A2(_2081_),
    .Y(_2082_),
    .B1(_2076_));
 sg13g2_nor2_1 _5128_ (.A(net1222),
    .B(_2082_),
    .Y(_0100_));
 sg13g2_o21ai_1 _5129_ (.B1(_2054_),
    .Y(_2083_),
    .A1(net1838),
    .A2(net1136));
 sg13g2_a21oi_1 _5130_ (.A1(_0660_),
    .A2(_2047_),
    .Y(_2084_),
    .B1(_2083_));
 sg13g2_xnor2_1 _5131_ (.Y(_2085_),
    .A(net1838),
    .B(_2079_));
 sg13g2_o21ai_1 _5132_ (.B1(net1203),
    .Y(_2086_),
    .A1(_2054_),
    .A2(_2085_));
 sg13g2_nor2_1 _5133_ (.A(_2084_),
    .B(_2086_),
    .Y(_2087_));
 sg13g2_nor3_1 _5134_ (.A(net1203),
    .B(net1838),
    .C(net1136),
    .Y(_2088_));
 sg13g2_nor3_1 _5135_ (.A(net1221),
    .B(_2087_),
    .C(net1839),
    .Y(_0101_));
 sg13g2_or2_1 _5136_ (.X(_2089_),
    .B(net1136),
    .A(net1894));
 sg13g2_nand2_1 _5137_ (.Y(_2090_),
    .A(net1611),
    .B(_0883_));
 sg13g2_nand3_1 _5138_ (.B(_1696_),
    .C(_2090_),
    .A(net1202),
    .Y(_2091_));
 sg13g2_inv_1 _5139_ (.Y(_2092_),
    .A(_2091_));
 sg13g2_o21ai_1 _5140_ (.B1(_2045_),
    .Y(_2093_),
    .A1(_2038_),
    .A2(_2041_));
 sg13g2_a21oi_1 _5141_ (.A1(_2052_),
    .A2(_2093_),
    .Y(_2094_),
    .B1(_0885_));
 sg13g2_nor2_1 _5142_ (.A(_0700_),
    .B(_2094_),
    .Y(_2095_));
 sg13g2_nor3_1 _5143_ (.A(net1552),
    .B(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[1] ),
    .C(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[0] ),
    .Y(_2096_));
 sg13g2_and2_1 _5144_ (.A(_0638_),
    .B(_2096_),
    .X(_2097_));
 sg13g2_and2_1 _5145_ (.A(_0637_),
    .B(_2097_),
    .X(_2098_));
 sg13g2_a21o_1 _5146_ (.A2(_2098_),
    .A1(net1174),
    .B1(_0882_),
    .X(_2099_));
 sg13g2_a21o_1 _5147_ (.A2(_2095_),
    .A1(_2089_),
    .B1(_2099_),
    .X(_2100_));
 sg13g2_a22oi_1 _5148_ (.Y(_2101_),
    .B1(_2092_),
    .B2(_2100_),
    .A2(_2089_),
    .A1(net1176));
 sg13g2_a22oi_1 _5149_ (.Y(_2102_),
    .B1(_2098_),
    .B2(net1174),
    .A2(_2051_),
    .A1(net1169));
 sg13g2_nand2_1 _5150_ (.Y(_2103_),
    .A(_2046_),
    .B(_2051_));
 sg13g2_a21oi_1 _5151_ (.A1(_2102_),
    .A2(_2103_),
    .Y(_2104_),
    .B1(_2091_));
 sg13g2_a21oi_1 _5152_ (.A1(net1202),
    .A2(_2091_),
    .Y(_2105_),
    .B1(net1136));
 sg13g2_a21o_1 _5153_ (.A2(_2105_),
    .A1(net1611),
    .B1(_2104_),
    .X(_2106_));
 sg13g2_nand2_1 _5154_ (.Y(_2107_),
    .A(net1873),
    .B(_2055_));
 sg13g2_nor2_1 _5155_ (.A(net1202),
    .B(net1874),
    .Y(_2108_));
 sg13g2_inv_1 _5156_ (.Y(_2109_),
    .A(_2108_));
 sg13g2_nand2_1 _5157_ (.Y(_2110_),
    .A(_2092_),
    .B(_2102_));
 sg13g2_a21o_1 _5158_ (.A2(net1874),
    .A1(_2095_),
    .B1(_2110_),
    .X(_2111_));
 sg13g2_a21oi_1 _5159_ (.A1(_2109_),
    .A2(_2111_),
    .Y(_2112_),
    .B1(_2106_));
 sg13g2_a21oi_1 _5160_ (.A1(_2101_),
    .A2(_2112_),
    .Y(_2113_),
    .B1(_0885_));
 sg13g2_a21o_1 _5161_ (.A2(_2113_),
    .A1(_2052_),
    .B1(net1137),
    .X(_2114_));
 sg13g2_nand2_2 _5162_ (.Y(_2115_),
    .A(net1203),
    .B(_2114_));
 sg13g2_or2_1 _5163_ (.X(_2116_),
    .B(_2115_),
    .A(net1201));
 sg13g2_o21ai_1 _5164_ (.B1(_2115_),
    .Y(_2117_),
    .A1(net1201),
    .A2(_2056_));
 sg13g2_a21oi_1 _5165_ (.A1(_2116_),
    .A2(_2117_),
    .Y(_0102_),
    .B1(net1221));
 sg13g2_xor2_1 _5166_ (.B(net1201),
    .A(net1886),
    .X(_2118_));
 sg13g2_nor2_1 _5167_ (.A(net1886),
    .B(_2056_),
    .Y(_2119_));
 sg13g2_mux2_1 _5168_ (.A0(_2118_),
    .A1(_2119_),
    .S(_2115_),
    .X(_2120_));
 sg13g2_nor2_1 _5169_ (.A(net1221),
    .B(_2120_),
    .Y(_0103_));
 sg13g2_o21ai_1 _5170_ (.B1(net1763),
    .Y(_2121_),
    .A1(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[1] ),
    .A2(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[0] ));
 sg13g2_nor2b_1 _5171_ (.A(_2049_),
    .B_N(_2121_),
    .Y(_2122_));
 sg13g2_or2_1 _5172_ (.X(_2123_),
    .B(_2122_),
    .A(_2115_));
 sg13g2_nand3_1 _5173_ (.B(_2055_),
    .C(_2115_),
    .A(net1763),
    .Y(_2124_));
 sg13g2_a21oi_1 _5174_ (.A1(_2123_),
    .A2(net1764),
    .Y(_0104_),
    .B1(net1221));
 sg13g2_nand2b_1 _5175_ (.Y(_2125_),
    .B(net1745),
    .A_N(_2049_));
 sg13g2_a21o_1 _5176_ (.A2(_2125_),
    .A1(_2050_),
    .B1(_2115_),
    .X(_2126_));
 sg13g2_nand3_1 _5177_ (.B(_2055_),
    .C(_2115_),
    .A(net1745),
    .Y(_2127_));
 sg13g2_a21oi_1 _5178_ (.A1(_2126_),
    .A2(net1746),
    .Y(_0105_),
    .B1(net1221));
 sg13g2_nor2_1 _5179_ (.A(net1806),
    .B(_2056_),
    .Y(_2128_));
 sg13g2_or2_1 _5180_ (.X(_2129_),
    .B(_2128_),
    .A(_2114_));
 sg13g2_a21oi_1 _5181_ (.A1(net1806),
    .A2(_2050_),
    .Y(_2130_),
    .B1(_0659_));
 sg13g2_a221oi_1 _5182_ (.B2(net1807),
    .C1(net1221),
    .B1(_2129_),
    .A1(_0659_),
    .Y(_0106_),
    .A2(_2128_));
 sg13g2_nor2_1 _5183_ (.A(net1173),
    .B(_2098_),
    .Y(_2131_));
 sg13g2_a21oi_2 _5184_ (.B1(_2131_),
    .Y(_2132_),
    .A2(_2051_),
    .A1(net1169));
 sg13g2_a21o_2 _5185_ (.A2(_2051_),
    .A1(net1168),
    .B1(_2131_),
    .X(_2133_));
 sg13g2_o21ai_1 _5186_ (.B1(net1202),
    .Y(_2134_),
    .A1(_2094_),
    .A2(_2133_));
 sg13g2_nand2_1 _5187_ (.Y(_2135_),
    .A(net1201),
    .B(_0661_));
 sg13g2_nand2b_1 _5188_ (.Y(_2136_),
    .B(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[0] ),
    .A_N(net1201));
 sg13g2_a21o_1 _5189_ (.A2(_2136_),
    .A1(_2135_),
    .B1(_2133_),
    .X(_2137_));
 sg13g2_o21ai_1 _5190_ (.B1(_2137_),
    .Y(_2138_),
    .A1(net1866),
    .A2(_2132_));
 sg13g2_mux2_1 _5191_ (.A0(_2138_),
    .A1(net1866),
    .S(net838),
    .X(_2139_));
 sg13g2_and2_1 _5192_ (.A(net1240),
    .B(_2139_),
    .X(_0107_));
 sg13g2_xnor2_1 _5193_ (.Y(_2140_),
    .A(net1651),
    .B(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[0] ));
 sg13g2_nor2b_1 _5194_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[1] ),
    .B_N(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[1] ),
    .Y(_2141_));
 sg13g2_xnor2_1 _5195_ (.Y(_2142_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[1] ),
    .B(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[1] ));
 sg13g2_xnor2_1 _5196_ (.Y(_2143_),
    .A(_2135_),
    .B(_2142_));
 sg13g2_nand2_1 _5197_ (.Y(_2144_),
    .A(_2133_),
    .B(_2140_));
 sg13g2_o21ai_1 _5198_ (.B1(_2144_),
    .Y(_2145_),
    .A1(_2133_),
    .A2(_2143_));
 sg13g2_o21ai_1 _5199_ (.B1(net1236),
    .Y(_2146_),
    .A1(net838),
    .A2(_2145_));
 sg13g2_a21oi_1 _5200_ (.A1(_0640_),
    .A2(net838),
    .Y(_0108_),
    .B1(_2146_));
 sg13g2_o21ai_1 _5201_ (.B1(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[2] ),
    .Y(_2147_),
    .A1(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[1] ),
    .A2(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[0] ));
 sg13g2_nor2b_1 _5202_ (.A(_2096_),
    .B_N(_2147_),
    .Y(_2148_));
 sg13g2_nand2b_1 _5203_ (.Y(_2149_),
    .B(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[2] ),
    .A_N(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[2] ));
 sg13g2_xor2_1 _5204_ (.B(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[2] ),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[2] ),
    .X(_2150_));
 sg13g2_a21oi_1 _5205_ (.A1(_2135_),
    .A2(_2142_),
    .Y(_2151_),
    .B1(_2141_));
 sg13g2_xor2_1 _5206_ (.B(_2151_),
    .A(_2150_),
    .X(_2152_));
 sg13g2_nand2_1 _5207_ (.Y(_2153_),
    .A(_2132_),
    .B(_2152_));
 sg13g2_o21ai_1 _5208_ (.B1(_2153_),
    .Y(_2154_),
    .A1(_2132_),
    .A2(_2148_));
 sg13g2_o21ai_1 _5209_ (.B1(net1240),
    .Y(_2155_),
    .A1(net838),
    .A2(_2154_));
 sg13g2_a21oi_1 _5210_ (.A1(_0639_),
    .A2(net838),
    .Y(_0109_),
    .B1(_2155_));
 sg13g2_nor2_1 _5211_ (.A(_0638_),
    .B(_2096_),
    .Y(_2156_));
 sg13g2_o21ai_1 _5212_ (.B1(_2133_),
    .Y(_2157_),
    .A1(_2097_),
    .A2(_2156_));
 sg13g2_nor2b_1 _5213_ (.A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[3] ),
    .B_N(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[3] ),
    .Y(_2158_));
 sg13g2_xnor2_1 _5214_ (.Y(_2159_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[3] ),
    .B(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[3] ));
 sg13g2_o21ai_1 _5215_ (.B1(_2149_),
    .Y(_2160_),
    .A1(_2150_),
    .A2(_2151_));
 sg13g2_xor2_1 _5216_ (.B(_2160_),
    .A(_2159_),
    .X(_2161_));
 sg13g2_a21oi_1 _5217_ (.A1(_2132_),
    .A2(_2161_),
    .Y(_2162_),
    .B1(net838));
 sg13g2_a221oi_1 _5218_ (.B2(_2162_),
    .C1(net1230),
    .B1(_2157_),
    .A1(_0638_),
    .Y(_0110_),
    .A2(_2134_));
 sg13g2_a21o_1 _5219_ (.A2(_2160_),
    .A1(_2159_),
    .B1(_2158_),
    .X(_2163_));
 sg13g2_xor2_1 _5220_ (.B(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[4] ),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[4] ),
    .X(_2164_));
 sg13g2_or2_1 _5221_ (.X(_2165_),
    .B(_2164_),
    .A(_2163_));
 sg13g2_a21oi_1 _5222_ (.A1(_2163_),
    .A2(_2164_),
    .Y(_2166_),
    .B1(_2133_));
 sg13g2_xnor2_1 _5223_ (.Y(_2167_),
    .A(net1706),
    .B(_2097_));
 sg13g2_a22oi_1 _5224_ (.Y(_2168_),
    .B1(_2167_),
    .B2(_2133_),
    .A2(_2166_),
    .A1(_2165_));
 sg13g2_o21ai_1 _5225_ (.B1(net1236),
    .Y(_2169_),
    .A1(net838),
    .A2(_2168_));
 sg13g2_a21oi_1 _5226_ (.A1(_0637_),
    .A2(net838),
    .Y(_0111_),
    .B1(_2169_));
 sg13g2_nor2_1 _5227_ (.A(net1220),
    .B(_2101_),
    .Y(_0112_));
 sg13g2_a21oi_1 _5228_ (.A1(_2109_),
    .A2(_2111_),
    .Y(_0113_),
    .B1(net1222));
 sg13g2_and2_1 _5229_ (.A(net1236),
    .B(_2106_),
    .X(_0114_));
 sg13g2_nor3_1 _5230_ (.A(net1176),
    .B(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[0] ),
    .C(_0701_),
    .Y(_2170_));
 sg13g2_nand2_2 _5231_ (.Y(_2171_),
    .A(net1202),
    .B(_0882_));
 sg13g2_o21ai_1 _5232_ (.B1(net1231),
    .Y(_2172_),
    .A1(net1699),
    .A2(net1152));
 sg13g2_a21oi_1 _5233_ (.A1(_0924_),
    .A2(net1152),
    .Y(_0115_),
    .B1(_2172_));
 sg13g2_o21ai_1 _5234_ (.B1(net1239),
    .Y(_2173_),
    .A1(_1423_),
    .A2(_2171_));
 sg13g2_a21oi_1 _5235_ (.A1(_0636_),
    .A2(_2171_),
    .Y(_0116_),
    .B1(_2173_));
 sg13g2_o21ai_1 _5236_ (.B1(net1239),
    .Y(_2174_),
    .A1(net1670),
    .A2(net1155));
 sg13g2_a21oi_1 _5237_ (.A1(_1049_),
    .A2(net1155),
    .Y(_0117_),
    .B1(net1671));
 sg13g2_o21ai_1 _5238_ (.B1(net1238),
    .Y(_2175_),
    .A1(_1443_),
    .A2(_2171_));
 sg13g2_a21oi_1 _5239_ (.A1(_0635_),
    .A2(_2171_),
    .Y(_0118_),
    .B1(_2175_));
 sg13g2_o21ai_1 _5240_ (.B1(net1238),
    .Y(_2176_),
    .A1(net1674),
    .A2(net1152));
 sg13g2_a21oi_1 _5241_ (.A1(_1007_),
    .A2(net1153),
    .Y(_0119_),
    .B1(_2176_));
 sg13g2_o21ai_1 _5242_ (.B1(net1231),
    .Y(_2177_),
    .A1(_1492_),
    .A2(_2171_));
 sg13g2_a21oi_1 _5243_ (.A1(_0634_),
    .A2(_2171_),
    .Y(_0120_),
    .B1(_2177_));
 sg13g2_o21ai_1 _5244_ (.B1(net1232),
    .Y(_2178_),
    .A1(net1669),
    .A2(net1153));
 sg13g2_a21oi_1 _5245_ (.A1(_1031_),
    .A2(net1153),
    .Y(_0121_),
    .B1(_2178_));
 sg13g2_o21ai_1 _5246_ (.B1(net1232),
    .Y(_2179_),
    .A1(net1722),
    .A2(net1153));
 sg13g2_a21oi_1 _5247_ (.A1(_1387_),
    .A2(net1153),
    .Y(_0122_),
    .B1(_2179_));
 sg13g2_o21ai_1 _5248_ (.B1(net1238),
    .Y(_2180_),
    .A1(net1664),
    .A2(net1154));
 sg13g2_a21oi_1 _5249_ (.A1(_1091_),
    .A2(net1154),
    .Y(_0123_),
    .B1(_2180_));
 sg13g2_o21ai_1 _5250_ (.B1(net1238),
    .Y(_2181_),
    .A1(net1700),
    .A2(net1152));
 sg13g2_a21oi_1 _5251_ (.A1(_1302_),
    .A2(net1152),
    .Y(_0124_),
    .B1(_2181_));
 sg13g2_o21ai_1 _5252_ (.B1(net1231),
    .Y(_2182_),
    .A1(net1650),
    .A2(net1151));
 sg13g2_a21oi_1 _5253_ (.A1(_0945_),
    .A2(net1151),
    .Y(_0125_),
    .B1(_2182_));
 sg13g2_o21ai_1 _5254_ (.B1(net1231),
    .Y(_2183_),
    .A1(net1668),
    .A2(net1151));
 sg13g2_a21oi_1 _5255_ (.A1(_1407_),
    .A2(net1151),
    .Y(_0126_),
    .B1(_2183_));
 sg13g2_o21ai_1 _5256_ (.B1(net1238),
    .Y(_2184_),
    .A1(net1683),
    .A2(net1154));
 sg13g2_a21oi_1 _5257_ (.A1(_1070_),
    .A2(net1154),
    .Y(_0127_),
    .B1(_2184_));
 sg13g2_o21ai_1 _5258_ (.B1(net1238),
    .Y(_2185_),
    .A1(net1657),
    .A2(net1154));
 sg13g2_a21oi_1 _5259_ (.A1(_1345_),
    .A2(net1154),
    .Y(_0128_),
    .B1(_2185_));
 sg13g2_o21ai_1 _5260_ (.B1(net1231),
    .Y(_2186_),
    .A1(net1656),
    .A2(net1151));
 sg13g2_a21oi_1 _5261_ (.A1(_0972_),
    .A2(net1151),
    .Y(_0129_),
    .B1(_2186_));
 sg13g2_o21ai_1 _5262_ (.B1(net1232),
    .Y(_2187_),
    .A1(net1673),
    .A2(net1151));
 sg13g2_a21oi_1 _5263_ (.A1(_1366_),
    .A2(net1151),
    .Y(_0130_),
    .B1(_2187_));
 sg13g2_o21ai_1 _5264_ (.B1(net1232),
    .Y(_2188_),
    .A1(net1708),
    .A2(net1153));
 sg13g2_a21oi_1 _5265_ (.A1(_0897_),
    .A2(net1153),
    .Y(_0131_),
    .B1(_2188_));
 sg13g2_o21ai_1 _5266_ (.B1(net1231),
    .Y(_2189_),
    .A1(net1713),
    .A2(net1152));
 sg13g2_a21oi_1 _5267_ (.A1(_1467_),
    .A2(net1152),
    .Y(_0132_),
    .B1(_2189_));
 sg13g2_o21ai_1 _5268_ (.B1(net1238),
    .Y(_2190_),
    .A1(_0989_),
    .A2(_2171_));
 sg13g2_a21oi_1 _5269_ (.A1(_0633_),
    .A2(_2171_),
    .Y(_0133_),
    .B1(_2190_));
 sg13g2_o21ai_1 _5270_ (.B1(net1238),
    .Y(_2191_),
    .A1(net1714),
    .A2(net1154));
 sg13g2_a21oi_1 _5271_ (.A1(_1324_),
    .A2(net1154),
    .Y(_0134_),
    .B1(_2191_));
 sg13g2_or4_1 _5272_ (.A(\vga_tetris._tetrisLogic_io_score_3[1] ),
    .B(_0688_),
    .C(\vga_tetris._tetrisLogic_io_score_3[2] ),
    .D(_0694_),
    .X(_2192_));
 sg13g2_nand3_1 _5273_ (.B(_0884_),
    .C(_2192_),
    .A(net1202),
    .Y(_2193_));
 sg13g2_nand4_1 _5274_ (.B(_0884_),
    .C(_2042_),
    .A(net1203),
    .Y(_2194_),
    .D(_2192_));
 sg13g2_nor4_2 _5275_ (.A(_0695_),
    .B(_2038_),
    .C(_2041_),
    .Y(_2195_),
    .D(_2193_));
 sg13g2_nor3_1 _5276_ (.A(net1756),
    .B(\vga_tetris._tetrisLogic_io_score_0[1] ),
    .C(_2195_),
    .Y(_2196_));
 sg13g2_nand2b_1 _5277_ (.Y(_2197_),
    .B(net1753),
    .A_N(_2196_));
 sg13g2_nor3_2 _5278_ (.A(_0692_),
    .B(_0696_),
    .C(_2196_),
    .Y(_2198_));
 sg13g2_nor3_1 _5279_ (.A(net1596),
    .B(net1789),
    .C(_2198_),
    .Y(_2199_));
 sg13g2_nand2b_2 _5280_ (.Y(_2200_),
    .B(net1759),
    .A_N(_2199_));
 sg13g2_nor3_2 _5281_ (.A(_0690_),
    .B(_0691_),
    .C(_2199_),
    .Y(_2201_));
 sg13g2_nor3_1 _5282_ (.A(net1585),
    .B(net1870),
    .C(_2201_),
    .Y(_2202_));
 sg13g2_nor2_1 _5283_ (.A(_0689_),
    .B(_2202_),
    .Y(_2203_));
 sg13g2_nor2_1 _5284_ (.A(net1660),
    .B(_2203_),
    .Y(_2204_));
 sg13g2_and2_1 _5285_ (.A(net1236),
    .B(_2026_),
    .X(_2205_));
 sg13g2_nand2_1 _5286_ (.Y(_2206_),
    .A(net1236),
    .B(_2026_));
 sg13g2_nor3_1 _5287_ (.A(_0688_),
    .B(_0689_),
    .C(_2202_),
    .Y(_2207_));
 sg13g2_nor3_1 _5288_ (.A(net1661),
    .B(net1133),
    .C(_2207_),
    .Y(_0135_));
 sg13g2_nor4_2 _5289_ (.A(_0687_),
    .B(_0688_),
    .C(_0689_),
    .Y(_2208_),
    .D(_2202_));
 sg13g2_or2_1 _5290_ (.X(_2209_),
    .B(_2208_),
    .A(net1740));
 sg13g2_xnor2_1 _5291_ (.Y(_2210_),
    .A(net1846),
    .B(_2207_));
 sg13g2_nand3_1 _5292_ (.B(_2209_),
    .C(_2210_),
    .A(net1686),
    .Y(_2211_));
 sg13g2_nand2b_1 _5293_ (.Y(_2212_),
    .B(_0694_),
    .A_N(_2210_));
 sg13g2_a21oi_1 _5294_ (.A1(net1687),
    .A2(_2212_),
    .Y(_0136_),
    .B1(net1133));
 sg13g2_nand2_1 _5295_ (.Y(_2213_),
    .A(net1740),
    .B(_2208_));
 sg13g2_nand3_1 _5296_ (.B(net1686),
    .C(_2208_),
    .A(net1740),
    .Y(_2214_));
 sg13g2_xnor2_1 _5297_ (.Y(_2215_),
    .A(net1740),
    .B(_2208_));
 sg13g2_a21o_1 _5298_ (.A2(_2210_),
    .A1(net1686),
    .B1(_2215_),
    .X(_2216_));
 sg13g2_a21oi_1 _5299_ (.A1(net1741),
    .A2(_2216_),
    .Y(_0137_),
    .B1(net1133));
 sg13g2_o21ai_1 _5300_ (.B1(_2213_),
    .Y(_2217_),
    .A1(_0694_),
    .A2(_2209_));
 sg13g2_and4_1 _5301_ (.A(_2205_),
    .B(_2210_),
    .C(_2214_),
    .D(_2217_),
    .X(_0138_));
 sg13g2_a21oi_1 _5302_ (.A1(net1200),
    .A2(\vga_tetris._inputs_io_downButtonActive ),
    .Y(_2218_),
    .B1(net1411));
 sg13g2_nand3_1 _5303_ (.B(net1411),
    .C(net1684),
    .A(\vga_tetris._tetrisLogic_io_gameOver ),
    .Y(_2219_));
 sg13g2_nand3_1 _5304_ (.B(_1511_),
    .C(_2219_),
    .A(net1243),
    .Y(_2220_));
 sg13g2_nor2_1 _5305_ (.A(net1412),
    .B(_2220_),
    .Y(_0139_));
 sg13g2_xnor2_1 _5306_ (.Y(_2221_),
    .A(net1790),
    .B(_2219_));
 sg13g2_and3_1 _5307_ (.X(_0140_),
    .A(net1243),
    .B(_1511_),
    .C(net1791));
 sg13g2_nor2_1 _5308_ (.A(_2030_),
    .B(_2031_),
    .Y(_0141_));
 sg13g2_a21oi_1 _5309_ (.A1(_0690_),
    .A2(_2200_),
    .Y(_2222_),
    .B1(net1133));
 sg13g2_nor2b_1 _5310_ (.A(_2201_),
    .B_N(_2222_),
    .Y(_0142_));
 sg13g2_xnor2_1 _5311_ (.Y(_2223_),
    .A(\vga_tetris._tetrisLogic_io_score_2[1] ),
    .B(_2201_));
 sg13g2_nand2_1 _5312_ (.Y(_2224_),
    .A(_2203_),
    .B(_2223_));
 sg13g2_o21ai_1 _5313_ (.B1(_2224_),
    .Y(_2225_),
    .A1(net1804),
    .A2(_2223_));
 sg13g2_and2_1 _5314_ (.A(_2205_),
    .B(net1805),
    .X(_0143_));
 sg13g2_nand3_1 _5315_ (.B(net1870),
    .C(_2201_),
    .A(net1585),
    .Y(_2226_));
 sg13g2_nand3_1 _5316_ (.B(_2223_),
    .C(_2226_),
    .A(_2203_),
    .Y(_2227_));
 sg13g2_a21oi_1 _5317_ (.A1(\vga_tetris._tetrisLogic_io_score_2[1] ),
    .A2(_2201_),
    .Y(_2228_),
    .B1(net1585));
 sg13g2_o21ai_1 _5318_ (.B1(_2227_),
    .Y(_2229_),
    .A1(\vga_tetris._tetrisLogic_io_score_2[3] ),
    .A2(_2226_));
 sg13g2_nor3_1 _5319_ (.A(net1133),
    .B(net1586),
    .C(_2229_),
    .Y(_0144_));
 sg13g2_a21oi_1 _5320_ (.A1(_0689_),
    .A2(_2226_),
    .Y(_2230_),
    .B1(net1133));
 sg13g2_nor2b_1 _5321_ (.A(_2203_),
    .B_N(_2230_),
    .Y(_0145_));
 sg13g2_a21oi_1 _5322_ (.A1(_0696_),
    .A2(_2197_),
    .Y(_2231_),
    .B1(net1133));
 sg13g2_nor2b_1 _5323_ (.A(_2198_),
    .B_N(_2231_),
    .Y(_0146_));
 sg13g2_xnor2_1 _5324_ (.Y(_2232_),
    .A(net1789),
    .B(_2198_));
 sg13g2_mux2_1 _5325_ (.A0(net1759),
    .A1(_2200_),
    .S(_2232_),
    .X(_2233_));
 sg13g2_nor2_1 _5326_ (.A(net1134),
    .B(_2233_),
    .Y(_0147_));
 sg13g2_nand3_1 _5327_ (.B(\vga_tetris._tetrisLogic_io_score_1[1] ),
    .C(_2198_),
    .A(net1596),
    .Y(_2234_));
 sg13g2_nand3b_1 _5328_ (.B(_2232_),
    .C(_2234_),
    .Y(_2235_),
    .A_N(_2200_));
 sg13g2_a21oi_1 _5329_ (.A1(\vga_tetris._tetrisLogic_io_score_1[1] ),
    .A2(_2198_),
    .Y(_2236_),
    .B1(net1596));
 sg13g2_o21ai_1 _5330_ (.B1(_2235_),
    .Y(_2237_),
    .A1(\vga_tetris._tetrisLogic_io_score_1[3] ),
    .A2(_2234_));
 sg13g2_nor3_1 _5331_ (.A(net1134),
    .B(net1597),
    .C(_2237_),
    .Y(_0148_));
 sg13g2_nand2_1 _5332_ (.Y(_2238_),
    .A(_2200_),
    .B(_2205_));
 sg13g2_a21oi_1 _5333_ (.A1(_0691_),
    .A2(_2234_),
    .Y(_0149_),
    .B1(_2238_));
 sg13g2_a21oi_1 _5334_ (.A1(_0695_),
    .A2(_2194_),
    .Y(_2239_),
    .B1(net1133));
 sg13g2_nor2b_1 _5335_ (.A(_2195_),
    .B_N(net1821),
    .Y(_0150_));
 sg13g2_nand2_1 _5336_ (.Y(_2240_),
    .A(\vga_tetris._tetrisLogic_io_score_0[1] ),
    .B(_2195_));
 sg13g2_xor2_1 _5337_ (.B(_2195_),
    .A(net1825),
    .X(_2241_));
 sg13g2_nor2_1 _5338_ (.A(_2197_),
    .B(_2241_),
    .Y(_2242_));
 sg13g2_a21oi_1 _5339_ (.A1(_0692_),
    .A2(_2241_),
    .Y(_2243_),
    .B1(_2242_));
 sg13g2_nor2_1 _5340_ (.A(net1134),
    .B(_2243_),
    .Y(_0151_));
 sg13g2_nand3_1 _5341_ (.B(\vga_tetris._tetrisLogic_io_score_0[1] ),
    .C(_2195_),
    .A(net1756),
    .Y(_2244_));
 sg13g2_a21oi_1 _5342_ (.A1(_0693_),
    .A2(_2240_),
    .Y(_2245_),
    .B1(net1134));
 sg13g2_o21ai_1 _5343_ (.B1(_2245_),
    .Y(_2246_),
    .A1(net1753),
    .A2(_2244_));
 sg13g2_a21oi_1 _5344_ (.A1(_2242_),
    .A2(_2244_),
    .Y(_0152_),
    .B1(net1754));
 sg13g2_nand2_1 _5345_ (.Y(_2247_),
    .A(_2197_),
    .B(_2205_));
 sg13g2_a21oi_1 _5346_ (.A1(_0692_),
    .A2(net1757),
    .Y(_0153_),
    .B1(_2247_));
 sg13g2_a21oi_1 _5347_ (.A1(_1511_),
    .A2(_2025_),
    .Y(_0154_),
    .B1(net1229));
 sg13g2_nand2_1 _5348_ (.Y(_2248_),
    .A(_0799_),
    .B(_0813_));
 sg13g2_or2_1 _5349_ (.X(_2249_),
    .B(_0785_),
    .A(_0767_));
 sg13g2_o21ai_1 _5350_ (.B1(net1149),
    .Y(_2250_),
    .A1(net1174),
    .A2(net1169));
 sg13g2_o21ai_1 _5351_ (.B1(_2250_),
    .Y(_2251_),
    .A1(net1149),
    .A2(_1910_));
 sg13g2_a21oi_1 _5352_ (.A1(_0764_),
    .A2(_2251_),
    .Y(_2252_),
    .B1(net1140));
 sg13g2_or3_1 _5353_ (.A(_0772_),
    .B(_2249_),
    .C(_2252_),
    .X(_2253_));
 sg13g2_nor2_2 _5354_ (.A(_2248_),
    .B(_2253_),
    .Y(_2254_));
 sg13g2_nor2_1 _5355_ (.A(net1465),
    .B(net958),
    .Y(_2255_));
 sg13g2_nand2_1 _5356_ (.Y(_2256_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[0] ),
    .B(net1170));
 sg13g2_a21oi_1 _5357_ (.A1(net1144),
    .A2(_2256_),
    .Y(_2257_),
    .B1(net1140));
 sg13g2_o21ai_1 _5358_ (.B1(_2257_),
    .Y(_2258_),
    .A1(net1387),
    .A2(net1144));
 sg13g2_a21oi_1 _5359_ (.A1(net958),
    .A2(net1130),
    .Y(_0155_),
    .B1(_2255_));
 sg13g2_nor2_1 _5360_ (.A(net1554),
    .B(net961),
    .Y(_2259_));
 sg13g2_nand2_1 _5361_ (.Y(_2260_),
    .A(net1404),
    .B(net1172));
 sg13g2_a21oi_1 _5362_ (.A1(net1148),
    .A2(_2260_),
    .Y(_2261_),
    .B1(net1141));
 sg13g2_o21ai_1 _5363_ (.B1(_2261_),
    .Y(_2262_),
    .A1(net1347),
    .A2(net1148));
 sg13g2_a21oi_1 _5364_ (.A1(net961),
    .A2(net1126),
    .Y(_0156_),
    .B1(_2259_));
 sg13g2_nor2_1 _5365_ (.A(net1500),
    .B(net961),
    .Y(_2263_));
 sg13g2_nand2_1 _5366_ (.Y(_2264_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[2] ),
    .B(net1172));
 sg13g2_a21oi_1 _5367_ (.A1(net1148),
    .A2(_2264_),
    .Y(_2265_),
    .B1(net1142));
 sg13g2_o21ai_1 _5368_ (.B1(_2265_),
    .Y(_2266_),
    .A1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[2] ),
    .A2(net1148));
 sg13g2_a21oi_1 _5369_ (.A1(net961),
    .A2(net1123),
    .Y(_0157_),
    .B1(_2263_));
 sg13g2_nor2_1 _5370_ (.A(net1473),
    .B(net963),
    .Y(_2267_));
 sg13g2_nand2_1 _5371_ (.Y(_2268_),
    .A(net831),
    .B(net1172));
 sg13g2_a21oi_1 _5372_ (.A1(net1148),
    .A2(_2268_),
    .Y(_2269_),
    .B1(net1141));
 sg13g2_o21ai_1 _5373_ (.B1(_2269_),
    .Y(_2270_),
    .A1(net1379),
    .A2(net1148));
 sg13g2_a21oi_1 _5374_ (.A1(net963),
    .A2(net1120),
    .Y(_0158_),
    .B1(_2267_));
 sg13g2_nor2_1 _5375_ (.A(net1532),
    .B(net962),
    .Y(_2271_));
 sg13g2_nand2_1 _5376_ (.Y(_2272_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[4] ),
    .B(net1170));
 sg13g2_a21oi_1 _5377_ (.A1(net1144),
    .A2(_2272_),
    .Y(_2273_),
    .B1(net1139));
 sg13g2_o21ai_1 _5378_ (.B1(_2273_),
    .Y(_2274_),
    .A1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[4] ),
    .A2(net1144));
 sg13g2_a21oi_1 _5379_ (.A1(net962),
    .A2(net1118),
    .Y(_0159_),
    .B1(_2271_));
 sg13g2_nor2_1 _5380_ (.A(net1458),
    .B(net959),
    .Y(_2275_));
 sg13g2_nand2_1 _5381_ (.Y(_2276_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[5] ),
    .B(net1170));
 sg13g2_a21oi_1 _5382_ (.A1(net1145),
    .A2(_2276_),
    .Y(_2277_),
    .B1(net1139));
 sg13g2_o21ai_1 _5383_ (.B1(_2277_),
    .Y(_2278_),
    .A1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[5] ),
    .A2(net1144));
 sg13g2_a21oi_1 _5384_ (.A1(net959),
    .A2(net1114),
    .Y(_0160_),
    .B1(_2275_));
 sg13g2_nor2_1 _5385_ (.A(net1482),
    .B(net960),
    .Y(_2279_));
 sg13g2_nand2_1 _5386_ (.Y(_2280_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[6] ),
    .B(net1173));
 sg13g2_a21oi_1 _5387_ (.A1(net1149),
    .A2(_2280_),
    .Y(_2281_),
    .B1(net1140));
 sg13g2_o21ai_1 _5388_ (.B1(_2281_),
    .Y(_2282_),
    .A1(net1388),
    .A2(net1149));
 sg13g2_a21oi_1 _5389_ (.A1(net960),
    .A2(net1111),
    .Y(_0161_),
    .B1(_2279_));
 sg13g2_nor2_1 _5390_ (.A(net1421),
    .B(net959),
    .Y(_2283_));
 sg13g2_nand2_1 _5391_ (.Y(_2284_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[7] ),
    .B(net1171));
 sg13g2_a21oi_1 _5392_ (.A1(_0736_),
    .A2(_2284_),
    .Y(_2285_),
    .B1(net1140));
 sg13g2_o21ai_1 _5393_ (.B1(_2285_),
    .Y(_2286_),
    .A1(net1367),
    .A2(_0736_));
 sg13g2_a21oi_1 _5394_ (.A1(net959),
    .A2(net1108),
    .Y(_0162_),
    .B1(_2283_));
 sg13g2_nor2_1 _5395_ (.A(net1548),
    .B(net962),
    .Y(_2287_));
 sg13g2_nand2_1 _5396_ (.Y(_2288_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[8] ),
    .B(net1172));
 sg13g2_a21oi_1 _5397_ (.A1(net1146),
    .A2(_2288_),
    .Y(_2289_),
    .B1(net1141));
 sg13g2_o21ai_1 _5398_ (.B1(_2289_),
    .Y(_2290_),
    .A1(net1506),
    .A2(net1147));
 sg13g2_a21oi_1 _5399_ (.A1(net962),
    .A2(net1107),
    .Y(_0163_),
    .B1(_2287_));
 sg13g2_nor2_1 _5400_ (.A(net1443),
    .B(net963),
    .Y(_2291_));
 sg13g2_nand2_1 _5401_ (.Y(_2292_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[9] ),
    .B(net1171));
 sg13g2_a21oi_1 _5402_ (.A1(net1146),
    .A2(_2292_),
    .Y(_2293_),
    .B1(net1141));
 sg13g2_o21ai_1 _5403_ (.B1(_2293_),
    .Y(_2294_),
    .A1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[9] ),
    .A2(net1146));
 sg13g2_a21oi_1 _5404_ (.A1(net963),
    .A2(net1102),
    .Y(_0164_),
    .B1(_2291_));
 sg13g2_nor2_1 _5405_ (.A(net1542),
    .B(net958),
    .Y(_2295_));
 sg13g2_nand2_1 _5406_ (.Y(_2296_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[10] ),
    .B(net1170));
 sg13g2_a21oi_1 _5407_ (.A1(net1143),
    .A2(_2296_),
    .Y(_2297_),
    .B1(net1139));
 sg13g2_o21ai_1 _5408_ (.B1(_2297_),
    .Y(_2298_),
    .A1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[10] ),
    .A2(net1143));
 sg13g2_a21oi_1 _5409_ (.A1(net958),
    .A2(net1100),
    .Y(_0165_),
    .B1(_2295_));
 sg13g2_nor2_1 _5410_ (.A(net1571),
    .B(net960),
    .Y(_2299_));
 sg13g2_nand2_1 _5411_ (.Y(_2300_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[11] ),
    .B(net1170));
 sg13g2_a21oi_1 _5412_ (.A1(net1143),
    .A2(_2300_),
    .Y(_2301_),
    .B1(net1139));
 sg13g2_o21ai_1 _5413_ (.B1(_2301_),
    .Y(_2302_),
    .A1(net1351),
    .A2(net1143));
 sg13g2_a21oi_1 _5414_ (.A1(net960),
    .A2(net1096),
    .Y(_0166_),
    .B1(_2299_));
 sg13g2_nor2_1 _5415_ (.A(net1601),
    .B(net961),
    .Y(_2303_));
 sg13g2_nand2_1 _5416_ (.Y(_2304_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[12] ),
    .B(net1172));
 sg13g2_a21oi_1 _5417_ (.A1(net1147),
    .A2(_2304_),
    .Y(_2305_),
    .B1(net1141));
 sg13g2_o21ai_1 _5418_ (.B1(_2305_),
    .Y(_2306_),
    .A1(net1370),
    .A2(net1147));
 sg13g2_a21oi_1 _5419_ (.A1(net961),
    .A2(net1092),
    .Y(_0167_),
    .B1(_2303_));
 sg13g2_nor2_1 _5420_ (.A(net1407),
    .B(net963),
    .Y(_2307_));
 sg13g2_nand2_1 _5421_ (.Y(_2308_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[13] ),
    .B(net1172));
 sg13g2_a21oi_1 _5422_ (.A1(net1146),
    .A2(_2308_),
    .Y(_2309_),
    .B1(net1141));
 sg13g2_o21ai_1 _5423_ (.B1(_2309_),
    .Y(_2310_),
    .A1(net1345),
    .A2(net1146));
 sg13g2_a21oi_1 _5424_ (.A1(net963),
    .A2(net1089),
    .Y(_0168_),
    .B1(_2307_));
 sg13g2_nor2_1 _5425_ (.A(net1515),
    .B(net958),
    .Y(_2311_));
 sg13g2_nand2_1 _5426_ (.Y(_2312_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[14] ),
    .B(net1170));
 sg13g2_a21oi_1 _5427_ (.A1(net1143),
    .A2(_2312_),
    .Y(_2313_),
    .B1(net1139));
 sg13g2_o21ai_1 _5428_ (.B1(_2313_),
    .Y(_2314_),
    .A1(net1900),
    .A2(net1143));
 sg13g2_a21oi_1 _5429_ (.A1(net958),
    .A2(net1087),
    .Y(_0169_),
    .B1(_2311_));
 sg13g2_nor2_1 _5430_ (.A(net1527),
    .B(net958),
    .Y(_2315_));
 sg13g2_nand2_1 _5431_ (.Y(_2316_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[15] ),
    .B(net1170));
 sg13g2_a21oi_1 _5432_ (.A1(net1143),
    .A2(_2316_),
    .Y(_2317_),
    .B1(net1139));
 sg13g2_o21ai_1 _5433_ (.B1(_2317_),
    .Y(_2318_),
    .A1(net1902),
    .A2(net1143));
 sg13g2_a21oi_1 _5434_ (.A1(net958),
    .A2(net1083),
    .Y(_0170_),
    .B1(_2315_));
 sg13g2_nor2_1 _5435_ (.A(net1501),
    .B(net959),
    .Y(_2319_));
 sg13g2_nand2_1 _5436_ (.Y(_2320_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[16] ),
    .B(net1171));
 sg13g2_a21oi_1 _5437_ (.A1(net1145),
    .A2(_2320_),
    .Y(_2321_),
    .B1(net1139));
 sg13g2_o21ai_1 _5438_ (.B1(_2321_),
    .Y(_2322_),
    .A1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[16] ),
    .A2(net1145));
 sg13g2_a21oi_1 _5439_ (.A1(net959),
    .A2(net1082),
    .Y(_0171_),
    .B1(_2319_));
 sg13g2_nor2_1 _5440_ (.A(net1428),
    .B(net959),
    .Y(_2323_));
 sg13g2_nand2_1 _5441_ (.Y(_2324_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[17] ),
    .B(net1170));
 sg13g2_a21oi_1 _5442_ (.A1(net1144),
    .A2(_2324_),
    .Y(_2325_),
    .B1(net1139));
 sg13g2_o21ai_1 _5443_ (.B1(_2325_),
    .Y(_2326_),
    .A1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[17] ),
    .A2(net1144));
 sg13g2_a21oi_1 _5444_ (.A1(net959),
    .A2(net1079),
    .Y(_0172_),
    .B1(_2323_));
 sg13g2_nor2_1 _5445_ (.A(net1541),
    .B(net961),
    .Y(_2327_));
 sg13g2_nand2_1 _5446_ (.Y(_2328_),
    .A(net1327),
    .B(net1172));
 sg13g2_a21oi_1 _5447_ (.A1(net1146),
    .A2(_2328_),
    .Y(_2329_),
    .B1(net1141));
 sg13g2_o21ai_1 _5448_ (.B1(_2329_),
    .Y(_2330_),
    .A1(net1377),
    .A2(net1147));
 sg13g2_a21oi_1 _5449_ (.A1(net961),
    .A2(net1074),
    .Y(_0173_),
    .B1(_2327_));
 sg13g2_nor2_1 _5450_ (.A(net1521),
    .B(net960),
    .Y(_2331_));
 sg13g2_nand2_1 _5451_ (.Y(_2332_),
    .A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[19] ),
    .B(net1173));
 sg13g2_a21oi_1 _5452_ (.A1(net1146),
    .A2(_2332_),
    .Y(_2333_),
    .B1(net1141));
 sg13g2_o21ai_1 _5453_ (.B1(_2333_),
    .Y(_2334_),
    .A1(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[19] ),
    .A2(net1146));
 sg13g2_a21oi_1 _5454_ (.A1(net960),
    .A2(net1071),
    .Y(_0174_),
    .B1(_2331_));
 sg13g2_nand2_1 _5455_ (.Y(_2335_),
    .A(net1589),
    .B(net1138));
 sg13g2_a21oi_2 _5456_ (.B1(net3),
    .Y(_2336_),
    .A2(net1138),
    .A1(net1589));
 sg13g2_nand2b_1 _5457_ (.Y(_2337_),
    .B(_2335_),
    .A_N(net3));
 sg13g2_nand2_2 _5458_ (.Y(_2338_),
    .A(net1241),
    .B(_2336_));
 sg13g2_nand4_1 _5459_ (.B(\vga_tetris.msTimer.msTimerQ[3] ),
    .C(\vga_tetris.msTimer.msTimerQ[13] ),
    .A(_0675_),
    .Y(_2339_),
    .D(\vga_tetris.msTimer.msTimerQ[14] ));
 sg13g2_nor4_1 _5460_ (.A(\vga_tetris.msTimer.msTimerQ[1] ),
    .B(\vga_tetris.msTimer.msTimerQ[0] ),
    .C(_1779_),
    .D(_2339_),
    .Y(_2340_));
 sg13g2_nor4_1 _5461_ (.A(\vga_tetris.msTimer.msTimerQ[4] ),
    .B(_0676_),
    .C(\vga_tetris.msTimer.msTimerQ[6] ),
    .D(\vga_tetris.msTimer.msTimerQ[11] ),
    .Y(_2341_));
 sg13g2_nand3_1 _5462_ (.B(_2340_),
    .C(_2341_),
    .A(_1776_),
    .Y(_2342_));
 sg13g2_nor2_1 _5463_ (.A(\vga_tetris._inputs_io_rotateButtonActive ),
    .B(_2342_),
    .Y(_2343_));
 sg13g2_and3_2 _5464_ (.X(_2344_),
    .A(_1776_),
    .B(_2340_),
    .C(_2341_));
 sg13g2_and2_1 _5465_ (.A(_0679_),
    .B(_2344_),
    .X(_2345_));
 sg13g2_nor2_1 _5466_ (.A(net1630),
    .B(_2345_),
    .Y(_2346_));
 sg13g2_and2_1 _5467_ (.A(net1630),
    .B(_2345_),
    .X(_2347_));
 sg13g2_nor3_1 _5468_ (.A(_2338_),
    .B(_2346_),
    .C(_2347_),
    .Y(_0175_));
 sg13g2_nand2_1 _5469_ (.Y(_2348_),
    .A(net1705),
    .B(_2347_));
 sg13g2_xnor2_1 _5470_ (.Y(_2349_),
    .A(net1705),
    .B(_2347_));
 sg13g2_nor2_1 _5471_ (.A(_2338_),
    .B(_2349_),
    .Y(_0176_));
 sg13g2_a21oi_1 _5472_ (.A1(net1705),
    .A2(_2347_),
    .Y(_2350_),
    .B1(net1836));
 sg13g2_and4_1 _5473_ (.A(net1836),
    .B(net1705),
    .C(net1630),
    .D(_2343_),
    .X(_2351_));
 sg13g2_nor3_1 _5474_ (.A(_2337_),
    .B(_2350_),
    .C(_2351_),
    .Y(_2352_));
 sg13g2_and2_1 _5475_ (.A(net1240),
    .B(_2352_),
    .X(_0177_));
 sg13g2_nor2_1 _5476_ (.A(net1842),
    .B(_2351_),
    .Y(_2353_));
 sg13g2_nor3_1 _5477_ (.A(_0680_),
    .B(_0681_),
    .C(_2348_),
    .Y(_2354_));
 sg13g2_nor3_1 _5478_ (.A(_2337_),
    .B(_2353_),
    .C(_2354_),
    .Y(_2355_));
 sg13g2_and2_1 _5479_ (.A(net1241),
    .B(_2355_),
    .X(_0178_));
 sg13g2_and3_2 _5480_ (.X(_2356_),
    .A(\vga_tetris.inputs.buttonTimerQ_0[3] ),
    .B(net1786),
    .C(_2351_));
 sg13g2_o21ai_1 _5481_ (.B1(_2336_),
    .Y(_2357_),
    .A1(net1786),
    .A2(_2354_));
 sg13g2_nor2_1 _5482_ (.A(_2356_),
    .B(_2357_),
    .Y(_2358_));
 sg13g2_nor3_1 _5483_ (.A(net1230),
    .B(_2356_),
    .C(net1787),
    .Y(_0179_));
 sg13g2_o21ai_1 _5484_ (.B1(_2336_),
    .Y(_2359_),
    .A1(net1818),
    .A2(_2356_));
 sg13g2_a21oi_1 _5485_ (.A1(net1818),
    .A2(_2356_),
    .Y(_2360_),
    .B1(_2359_));
 sg13g2_and2_1 _5486_ (.A(net1241),
    .B(net1819),
    .X(_0180_));
 sg13g2_a21oi_1 _5487_ (.A1(\vga_tetris.inputs.buttonTimerQ_0[5] ),
    .A2(_2356_),
    .Y(_2361_),
    .B1(net1394));
 sg13g2_nand3_1 _5488_ (.B(\vga_tetris.inputs.buttonTimerQ_0[5] ),
    .C(_2356_),
    .A(net1394),
    .Y(_2362_));
 sg13g2_nand2b_1 _5489_ (.Y(_2363_),
    .B(_2362_),
    .A_N(_2338_));
 sg13g2_nor2_1 _5490_ (.A(net1395),
    .B(_2363_),
    .Y(_0181_));
 sg13g2_xor2_1 _5491_ (.B(_2362_),
    .A(net1695),
    .X(_2364_));
 sg13g2_nor2_1 _5492_ (.A(_2338_),
    .B(net1696),
    .Y(_0182_));
 sg13g2_nand2_1 _5493_ (.Y(_2365_),
    .A(net1833),
    .B(_1705_));
 sg13g2_a21oi_1 _5494_ (.A1(\vga_tetris._inputs_io_leftButtonActive ),
    .A2(_1705_),
    .Y(_2366_),
    .B1(net1));
 sg13g2_nand2b_1 _5495_ (.Y(_2367_),
    .B(_2365_),
    .A_N(net1));
 sg13g2_nand2_2 _5496_ (.Y(_2368_),
    .A(net1244),
    .B(_2366_));
 sg13g2_nor2_1 _5497_ (.A(\vga_tetris._inputs_io_leftButtonActive ),
    .B(_2342_),
    .Y(_2369_));
 sg13g2_nor2b_1 _5498_ (.A(\vga_tetris._inputs_io_leftButtonActive ),
    .B_N(_2344_),
    .Y(_2370_));
 sg13g2_nor2_1 _5499_ (.A(net1637),
    .B(_2370_),
    .Y(_2371_));
 sg13g2_and2_1 _5500_ (.A(net1637),
    .B(_2370_),
    .X(_2372_));
 sg13g2_nor3_1 _5501_ (.A(_2368_),
    .B(net1638),
    .C(_2372_),
    .Y(_0183_));
 sg13g2_xnor2_1 _5502_ (.Y(_2373_),
    .A(net1715),
    .B(_2372_));
 sg13g2_nor2_1 _5503_ (.A(_2368_),
    .B(net1716),
    .Y(_0184_));
 sg13g2_a21oi_1 _5504_ (.A1(net1715),
    .A2(_2372_),
    .Y(_2374_),
    .B1(net1802));
 sg13g2_and4_1 _5505_ (.A(net1802),
    .B(\vga_tetris.inputs.buttonTimerQ_1[1] ),
    .C(\vga_tetris.inputs.buttonTimerQ_1[0] ),
    .D(_2369_),
    .X(_2375_));
 sg13g2_nor3_1 _5506_ (.A(_2367_),
    .B(_2374_),
    .C(_2375_),
    .Y(_2376_));
 sg13g2_and2_1 _5507_ (.A(net1244),
    .B(net1803),
    .X(_0185_));
 sg13g2_o21ai_1 _5508_ (.B1(_2366_),
    .Y(_2377_),
    .A1(net1814),
    .A2(_2375_));
 sg13g2_a21oi_1 _5509_ (.A1(net1814),
    .A2(_2375_),
    .Y(_2378_),
    .B1(_2377_));
 sg13g2_and2_1 _5510_ (.A(net1241),
    .B(net1815),
    .X(_0186_));
 sg13g2_a21oi_1 _5511_ (.A1(\vga_tetris.inputs.buttonTimerQ_1[3] ),
    .A2(_2375_),
    .Y(_2379_),
    .B1(net1796));
 sg13g2_and3_1 _5512_ (.X(_2380_),
    .A(net1814),
    .B(net1796),
    .C(_2375_));
 sg13g2_nor3_1 _5513_ (.A(_2367_),
    .B(net1797),
    .C(_2380_),
    .Y(_2381_));
 sg13g2_and2_1 _5514_ (.A(net1241),
    .B(net1798),
    .X(_0187_));
 sg13g2_nor2_1 _5515_ (.A(net1837),
    .B(_2380_),
    .Y(_2382_));
 sg13g2_and2_1 _5516_ (.A(net1837),
    .B(_2380_),
    .X(_2383_));
 sg13g2_nor3_1 _5517_ (.A(_2367_),
    .B(_2382_),
    .C(_2383_),
    .Y(_2384_));
 sg13g2_and2_1 _5518_ (.A(net1244),
    .B(_2384_),
    .X(_0188_));
 sg13g2_nor2_1 _5519_ (.A(net1616),
    .B(_2383_),
    .Y(_2385_));
 sg13g2_and2_1 _5520_ (.A(net1616),
    .B(_2383_),
    .X(_2386_));
 sg13g2_nor3_1 _5521_ (.A(_2368_),
    .B(net1617),
    .C(_2386_),
    .Y(_0189_));
 sg13g2_xnor2_1 _5522_ (.Y(_2387_),
    .A(net1631),
    .B(_2386_));
 sg13g2_nor2_1 _5523_ (.A(_2368_),
    .B(net1632),
    .Y(_0190_));
 sg13g2_nand2_1 _5524_ (.Y(_2388_),
    .A(net1843),
    .B(net1138));
 sg13g2_a21oi_1 _5525_ (.A1(net1843),
    .A2(net1138),
    .Y(_2389_),
    .B1(net2));
 sg13g2_nand2b_2 _5526_ (.Y(_2390_),
    .B(_2388_),
    .A_N(net2));
 sg13g2_nand2_2 _5527_ (.Y(_2391_),
    .A(net1240),
    .B(_2389_));
 sg13g2_nor3_1 _5528_ (.A(\vga_tetris._inputs_io_rightButtonActive ),
    .B(_0678_),
    .C(_2342_),
    .Y(_2392_));
 sg13g2_a21oi_1 _5529_ (.A1(_0677_),
    .A2(_2344_),
    .Y(_2393_),
    .B1(net804));
 sg13g2_nor3_1 _5530_ (.A(_2391_),
    .B(_2392_),
    .C(net805),
    .Y(_0191_));
 sg13g2_nor2_1 _5531_ (.A(net1565),
    .B(_2392_),
    .Y(_2394_));
 sg13g2_and2_1 _5532_ (.A(net1565),
    .B(_2392_),
    .X(_2395_));
 sg13g2_nor3_1 _5533_ (.A(_2391_),
    .B(net1566),
    .C(_2395_),
    .Y(_0192_));
 sg13g2_nor2_1 _5534_ (.A(net1831),
    .B(_2395_),
    .Y(_2396_));
 sg13g2_and2_1 _5535_ (.A(net1831),
    .B(_2395_),
    .X(_2397_));
 sg13g2_nor3_1 _5536_ (.A(_2390_),
    .B(_2396_),
    .C(_2397_),
    .Y(_2398_));
 sg13g2_and2_1 _5537_ (.A(net1240),
    .B(net1832),
    .X(_0193_));
 sg13g2_o21ai_1 _5538_ (.B1(_2389_),
    .Y(_2399_),
    .A1(net1823),
    .A2(_2397_));
 sg13g2_a21oi_1 _5539_ (.A1(net1823),
    .A2(_2397_),
    .Y(_2400_),
    .B1(_2399_));
 sg13g2_and2_1 _5540_ (.A(net1240),
    .B(net1824),
    .X(_0194_));
 sg13g2_a21oi_1 _5541_ (.A1(\vga_tetris.inputs.buttonTimerQ_2[3] ),
    .A2(_2397_),
    .Y(_2401_),
    .B1(net1799));
 sg13g2_and3_1 _5542_ (.X(_2402_),
    .A(\vga_tetris.inputs.buttonTimerQ_2[3] ),
    .B(net1799),
    .C(_2397_));
 sg13g2_nor3_1 _5543_ (.A(_2390_),
    .B(net1800),
    .C(_2402_),
    .Y(_2403_));
 sg13g2_and2_1 _5544_ (.A(net1240),
    .B(net1801),
    .X(_0195_));
 sg13g2_nor2_1 _5545_ (.A(net1748),
    .B(_2402_),
    .Y(_2404_));
 sg13g2_and2_1 _5546_ (.A(net1748),
    .B(_2402_),
    .X(_2405_));
 sg13g2_nor4_1 _5547_ (.A(net1228),
    .B(_2390_),
    .C(net1749),
    .D(_2405_),
    .Y(_0196_));
 sg13g2_nand2_1 _5548_ (.Y(_2406_),
    .A(\vga_tetris.inputs.buttonTimerQ_2[6] ),
    .B(_2405_));
 sg13g2_xnor2_1 _5549_ (.Y(_2407_),
    .A(net1689),
    .B(_2405_));
 sg13g2_nor2_1 _5550_ (.A(_2391_),
    .B(net1690),
    .Y(_0197_));
 sg13g2_xor2_1 _5551_ (.B(_2406_),
    .A(net1675),
    .X(_2408_));
 sg13g2_nor2_1 _5552_ (.A(_2391_),
    .B(net1676),
    .Y(_0198_));
 sg13g2_a21o_2 _5553_ (.A2(_1705_),
    .A1(net1684),
    .B1(net4),
    .X(_2409_));
 sg13g2_and2_1 _5554_ (.A(_0683_),
    .B(_2344_),
    .X(_2410_));
 sg13g2_nor3_1 _5555_ (.A(net1684),
    .B(_0685_),
    .C(_2342_),
    .Y(_2411_));
 sg13g2_xnor2_1 _5556_ (.Y(_2412_),
    .A(net1770),
    .B(_2410_));
 sg13g2_nor2_1 _5557_ (.A(net1070),
    .B(_2412_),
    .Y(_2413_));
 sg13g2_nor3_1 _5558_ (.A(net1230),
    .B(net1070),
    .C(_2412_),
    .Y(_0199_));
 sg13g2_nor2_1 _5559_ (.A(net1847),
    .B(_2411_),
    .Y(_2414_));
 sg13g2_and2_1 _5560_ (.A(net1847),
    .B(_2411_),
    .X(_2415_));
 sg13g2_nor3_1 _5561_ (.A(_2409_),
    .B(_2414_),
    .C(_2415_),
    .Y(_2416_));
 sg13g2_and2_1 _5562_ (.A(net1244),
    .B(_2416_),
    .X(_0200_));
 sg13g2_nor2_1 _5563_ (.A(net1844),
    .B(_2415_),
    .Y(_2417_));
 sg13g2_and2_1 _5564_ (.A(net1844),
    .B(_2415_),
    .X(_2418_));
 sg13g2_and4_1 _5565_ (.A(net1770),
    .B(net1895),
    .C(\vga_tetris.inputs.buttonTimerQ_3[2] ),
    .D(_2410_),
    .X(_2419_));
 sg13g2_nor3_1 _5566_ (.A(net1070),
    .B(net1845),
    .C(_2418_),
    .Y(_2420_));
 sg13g2_and2_1 _5567_ (.A(net1244),
    .B(_2420_),
    .X(_0201_));
 sg13g2_xnor2_1 _5568_ (.Y(_2421_),
    .A(net1773),
    .B(_2419_));
 sg13g2_nor2_1 _5569_ (.A(net1070),
    .B(_2421_),
    .Y(_2422_));
 sg13g2_nor3_1 _5570_ (.A(net1229),
    .B(net1070),
    .C(net1774),
    .Y(_0202_));
 sg13g2_a21oi_1 _5571_ (.A1(net1773),
    .A2(net1896),
    .Y(_2423_),
    .B1(net1828));
 sg13g2_and3_1 _5572_ (.X(_2424_),
    .A(net1773),
    .B(net1828),
    .C(_2418_));
 sg13g2_nor3_1 _5573_ (.A(_2409_),
    .B(_2423_),
    .C(_2424_),
    .Y(_2425_));
 sg13g2_and2_1 _5574_ (.A(net1245),
    .B(_2425_),
    .X(_0203_));
 sg13g2_nor2_1 _5575_ (.A(net1841),
    .B(_2424_),
    .Y(_2426_));
 sg13g2_and2_1 _5576_ (.A(net1841),
    .B(_2424_),
    .X(_2427_));
 sg13g2_nand4_1 _5577_ (.B(\vga_tetris.inputs.buttonTimerQ_3[4] ),
    .C(\vga_tetris.inputs.buttonTimerQ_3[5] ),
    .A(\vga_tetris.inputs.buttonTimerQ_3[3] ),
    .Y(_2428_),
    .D(_2419_));
 sg13g2_nor3_1 _5578_ (.A(net1070),
    .B(_2426_),
    .C(_2427_),
    .Y(_2429_));
 sg13g2_and2_1 _5579_ (.A(net1244),
    .B(_2429_),
    .X(_0204_));
 sg13g2_nor2_1 _5580_ (.A(net1829),
    .B(_2427_),
    .Y(_2430_));
 sg13g2_nor2_1 _5581_ (.A(_0686_),
    .B(_2428_),
    .Y(_2431_));
 sg13g2_nor3_1 _5582_ (.A(net1070),
    .B(net1830),
    .C(_2431_),
    .Y(_2432_));
 sg13g2_and2_1 _5583_ (.A(net1244),
    .B(_2432_),
    .X(_0205_));
 sg13g2_a21oi_1 _5584_ (.A1(net1767),
    .A2(_2431_),
    .Y(_2433_),
    .B1(net1070));
 sg13g2_o21ai_1 _5585_ (.B1(net1768),
    .Y(_2434_),
    .A1(net1767),
    .A2(_2431_));
 sg13g2_nor2_1 _5586_ (.A(net1230),
    .B(net1769),
    .Y(_0206_));
 sg13g2_nor3_1 _5587_ (.A(_2352_),
    .B(_2355_),
    .C(_2358_),
    .Y(_2435_));
 sg13g2_nand2_1 _5588_ (.Y(_2436_),
    .A(net1394),
    .B(_2360_));
 sg13g2_o21ai_1 _5589_ (.B1(_0679_),
    .Y(_2437_),
    .A1(_2435_),
    .A2(_2436_));
 sg13g2_nand3_1 _5590_ (.B(_2335_),
    .C(_2437_),
    .A(net1241),
    .Y(_2438_));
 sg13g2_nand2b_1 _5591_ (.Y(_0207_),
    .B(_2438_),
    .A_N(_0182_));
 sg13g2_or3_1 _5592_ (.A(_2376_),
    .B(_2378_),
    .C(_2381_),
    .X(_2439_));
 sg13g2_nand3_1 _5593_ (.B(_2384_),
    .C(_2439_),
    .A(net1616),
    .Y(_2440_));
 sg13g2_nand2b_1 _5594_ (.Y(_2441_),
    .B(_2440_),
    .A_N(net1833));
 sg13g2_nand3_1 _5595_ (.B(_2365_),
    .C(_2441_),
    .A(net1244),
    .Y(_2442_));
 sg13g2_nand2b_1 _5596_ (.Y(_0208_),
    .B(net1834),
    .A_N(_0190_));
 sg13g2_nor3_1 _5597_ (.A(_2398_),
    .B(_2400_),
    .C(_2403_),
    .Y(_2443_));
 sg13g2_nor4_1 _5598_ (.A(_2390_),
    .B(_2404_),
    .C(_2405_),
    .D(_2443_),
    .Y(_2444_));
 sg13g2_a21o_1 _5599_ (.A2(_2444_),
    .A1(net1689),
    .B1(net1843),
    .X(_2445_));
 sg13g2_nand3_1 _5600_ (.B(_2388_),
    .C(_2445_),
    .A(net1240),
    .Y(_2446_));
 sg13g2_nand2b_1 _5601_ (.Y(_0209_),
    .B(_2446_),
    .A_N(_0198_));
 sg13g2_nor4_1 _5602_ (.A(net1684),
    .B(_2413_),
    .C(_2416_),
    .D(_2420_),
    .Y(_2447_));
 sg13g2_nand2b_1 _5603_ (.Y(_2448_),
    .B(_2447_),
    .A_N(_2422_));
 sg13g2_nor4_1 _5604_ (.A(_2425_),
    .B(_2429_),
    .C(_2432_),
    .D(_2448_),
    .Y(_2449_));
 sg13g2_a221oi_1 _5605_ (.B2(_2449_),
    .C1(net1230),
    .B1(_2434_),
    .A1(net1684),
    .Y(_0210_),
    .A2(net1138));
 sg13g2_or2_1 _5606_ (.X(_2450_),
    .B(\vga_tetris._vgaController_io_vSync ),
    .A(net1220));
 sg13g2_nor3_1 _5607_ (.A(net1177),
    .B(net1199),
    .C(_2450_),
    .Y(_0211_));
 sg13g2_nor2_2 _5608_ (.A(_0773_),
    .B(_2252_),
    .Y(_2451_));
 sg13g2_nand3b_1 _5609_ (.B(_2451_),
    .C(_0800_),
    .Y(_2452_),
    .A_N(_0813_));
 sg13g2_nor2_1 _5610_ (.A(_2249_),
    .B(_2452_),
    .Y(_2453_));
 sg13g2_nor2_1 _5611_ (.A(net1539),
    .B(net952),
    .Y(_2454_));
 sg13g2_a21oi_1 _5612_ (.A1(net1131),
    .A2(net952),
    .Y(_0212_),
    .B1(_2454_));
 sg13g2_nor2_1 _5613_ (.A(net1547),
    .B(net954),
    .Y(_2455_));
 sg13g2_a21oi_1 _5614_ (.A1(net1129),
    .A2(net954),
    .Y(_0213_),
    .B1(_2455_));
 sg13g2_nor2_1 _5615_ (.A(net1433),
    .B(net955),
    .Y(_2456_));
 sg13g2_a21oi_1 _5616_ (.A1(_2266_),
    .A2(net955),
    .Y(_0214_),
    .B1(_2456_));
 sg13g2_nor2_1 _5617_ (.A(net1559),
    .B(net954),
    .Y(_2457_));
 sg13g2_a21oi_1 _5618_ (.A1(net1121),
    .A2(net954),
    .Y(_0215_),
    .B1(_2457_));
 sg13g2_nor2_1 _5619_ (.A(net1470),
    .B(net955),
    .Y(_2458_));
 sg13g2_a21oi_1 _5620_ (.A1(_2274_),
    .A2(net955),
    .Y(_0216_),
    .B1(_2458_));
 sg13g2_nor2_1 _5621_ (.A(net1564),
    .B(net951),
    .Y(_2459_));
 sg13g2_a21oi_1 _5622_ (.A1(net1116),
    .A2(net951),
    .Y(_0217_),
    .B1(_2459_));
 sg13g2_nor2_1 _5623_ (.A(net1467),
    .B(net953),
    .Y(_2460_));
 sg13g2_a21oi_1 _5624_ (.A1(_2282_),
    .A2(net953),
    .Y(_0218_),
    .B1(_2460_));
 sg13g2_nor2_1 _5625_ (.A(net1556),
    .B(net953),
    .Y(_2461_));
 sg13g2_a21oi_1 _5626_ (.A1(net1110),
    .A2(net953),
    .Y(_0219_),
    .B1(_2461_));
 sg13g2_nor2_1 _5627_ (.A(net1572),
    .B(net954),
    .Y(_2462_));
 sg13g2_a21oi_1 _5628_ (.A1(net1107),
    .A2(net954),
    .Y(_0220_),
    .B1(_2462_));
 sg13g2_nor2_1 _5629_ (.A(net1466),
    .B(net956),
    .Y(_2463_));
 sg13g2_a21oi_1 _5630_ (.A1(net1104),
    .A2(net956),
    .Y(_0221_),
    .B1(_2463_));
 sg13g2_nor2_1 _5631_ (.A(net1530),
    .B(net951),
    .Y(_2464_));
 sg13g2_a21oi_1 _5632_ (.A1(net1101),
    .A2(net951),
    .Y(_0222_),
    .B1(_2464_));
 sg13g2_nor2_1 _5633_ (.A(net1490),
    .B(net952),
    .Y(_2465_));
 sg13g2_a21oi_1 _5634_ (.A1(net1098),
    .A2(net952),
    .Y(_0223_),
    .B1(_2465_));
 sg13g2_nor2_1 _5635_ (.A(net1474),
    .B(net956),
    .Y(_2466_));
 sg13g2_a21oi_1 _5636_ (.A1(net1095),
    .A2(net956),
    .Y(_0224_),
    .B1(_2466_));
 sg13g2_nor2_1 _5637_ (.A(net1461),
    .B(net956),
    .Y(_2467_));
 sg13g2_a21oi_1 _5638_ (.A1(net1090),
    .A2(net956),
    .Y(_0225_),
    .B1(_2467_));
 sg13g2_nor2_1 _5639_ (.A(net1510),
    .B(net951),
    .Y(_2468_));
 sg13g2_a21oi_1 _5640_ (.A1(net1087),
    .A2(net951),
    .Y(_0226_),
    .B1(_2468_));
 sg13g2_nor2_1 _5641_ (.A(net1398),
    .B(net951),
    .Y(_2469_));
 sg13g2_a21oi_1 _5642_ (.A1(net1085),
    .A2(net951),
    .Y(_0227_),
    .B1(_2469_));
 sg13g2_nor2_1 _5643_ (.A(net1476),
    .B(net957),
    .Y(_2470_));
 sg13g2_a21oi_1 _5644_ (.A1(net1081),
    .A2(net953),
    .Y(_0228_),
    .B1(_2470_));
 sg13g2_nor2_1 _5645_ (.A(net1417),
    .B(net953),
    .Y(_2471_));
 sg13g2_a21oi_1 _5646_ (.A1(net1078),
    .A2(net957),
    .Y(_0229_),
    .B1(_2471_));
 sg13g2_nor2_1 _5647_ (.A(net1568),
    .B(net954),
    .Y(_2472_));
 sg13g2_a21oi_1 _5648_ (.A1(_2330_),
    .A2(net954),
    .Y(_0230_),
    .B1(_2472_));
 sg13g2_nor2_1 _5649_ (.A(net1555),
    .B(net956),
    .Y(_2473_));
 sg13g2_a21oi_1 _5650_ (.A1(net1072),
    .A2(net956),
    .Y(_0231_),
    .B1(_2473_));
 sg13g2_nor2_1 _5651_ (.A(_0800_),
    .B(_0813_),
    .Y(_2474_));
 sg13g2_nand2_2 _5652_ (.Y(_2475_),
    .A(_2451_),
    .B(_2474_));
 sg13g2_nor2_1 _5653_ (.A(_2249_),
    .B(_2475_),
    .Y(_2476_));
 sg13g2_nor2_1 _5654_ (.A(net1430),
    .B(net946),
    .Y(_2477_));
 sg13g2_a21oi_1 _5655_ (.A1(net1131),
    .A2(net946),
    .Y(_0232_),
    .B1(_2477_));
 sg13g2_nor2_1 _5656_ (.A(net1446),
    .B(net948),
    .Y(_2478_));
 sg13g2_a21oi_1 _5657_ (.A1(net1128),
    .A2(net948),
    .Y(_0233_),
    .B1(_2478_));
 sg13g2_nor2_1 _5658_ (.A(net1441),
    .B(net948),
    .Y(_2479_));
 sg13g2_a21oi_1 _5659_ (.A1(net1123),
    .A2(net948),
    .Y(_0234_),
    .B1(_2479_));
 sg13g2_nor2_1 _5660_ (.A(net1391),
    .B(net949),
    .Y(_2480_));
 sg13g2_a21oi_1 _5661_ (.A1(net1120),
    .A2(net949),
    .Y(_0235_),
    .B1(_2480_));
 sg13g2_nor2_1 _5662_ (.A(net1494),
    .B(net947),
    .Y(_2481_));
 sg13g2_a21oi_1 _5663_ (.A1(net1119),
    .A2(net947),
    .Y(_0236_),
    .B1(_2481_));
 sg13g2_nor2_1 _5664_ (.A(net1575),
    .B(net944),
    .Y(_2482_));
 sg13g2_a21oi_1 _5665_ (.A1(net1116),
    .A2(net944),
    .Y(_0237_),
    .B1(_2482_));
 sg13g2_nor2_1 _5666_ (.A(net1511),
    .B(net949),
    .Y(_2483_));
 sg13g2_a21oi_1 _5667_ (.A1(net1111),
    .A2(net949),
    .Y(_0238_),
    .B1(_2483_));
 sg13g2_nor2_1 _5668_ (.A(net1425),
    .B(net945),
    .Y(_2484_));
 sg13g2_a21oi_1 _5669_ (.A1(net1108),
    .A2(net945),
    .Y(_0239_),
    .B1(_2484_));
 sg13g2_nor2_1 _5670_ (.A(net1492),
    .B(net948),
    .Y(_2485_));
 sg13g2_a21oi_1 _5671_ (.A1(net1107),
    .A2(net948),
    .Y(_0240_),
    .B1(_2485_));
 sg13g2_nor2_1 _5672_ (.A(net1397),
    .B(net949),
    .Y(_2486_));
 sg13g2_a21oi_1 _5673_ (.A1(net1102),
    .A2(net949),
    .Y(_0241_),
    .B1(_2486_));
 sg13g2_nor2_1 _5674_ (.A(net1545),
    .B(net944),
    .Y(_2487_));
 sg13g2_a21oi_1 _5675_ (.A1(net1099),
    .A2(net944),
    .Y(_0242_),
    .B1(_2487_));
 sg13g2_nor2_1 _5676_ (.A(net1392),
    .B(net946),
    .Y(_2488_));
 sg13g2_a21oi_1 _5677_ (.A1(net1098),
    .A2(net946),
    .Y(_0243_),
    .B1(_2488_));
 sg13g2_nor2_1 _5678_ (.A(net1546),
    .B(net947),
    .Y(_2489_));
 sg13g2_a21oi_1 _5679_ (.A1(net1094),
    .A2(net947),
    .Y(_0244_),
    .B1(_2489_));
 sg13g2_nor2_1 _5680_ (.A(net1519),
    .B(net947),
    .Y(_2490_));
 sg13g2_a21oi_1 _5681_ (.A1(net1091),
    .A2(net947),
    .Y(_0245_),
    .B1(_2490_));
 sg13g2_nor2_1 _5682_ (.A(net1442),
    .B(net944),
    .Y(_2491_));
 sg13g2_a21oi_1 _5683_ (.A1(net1086),
    .A2(net944),
    .Y(_0246_),
    .B1(_2491_));
 sg13g2_nor2_1 _5684_ (.A(net1485),
    .B(net944),
    .Y(_2492_));
 sg13g2_a21oi_1 _5685_ (.A1(net1083),
    .A2(net944),
    .Y(_0247_),
    .B1(_2492_));
 sg13g2_nor2_1 _5686_ (.A(net1524),
    .B(net945),
    .Y(_2493_));
 sg13g2_a21oi_1 _5687_ (.A1(net1080),
    .A2(net945),
    .Y(_0248_),
    .B1(_2493_));
 sg13g2_nor2_1 _5688_ (.A(net1452),
    .B(net945),
    .Y(_2494_));
 sg13g2_a21oi_1 _5689_ (.A1(net1078),
    .A2(net945),
    .Y(_0249_),
    .B1(_2494_));
 sg13g2_nor2_1 _5690_ (.A(net1427),
    .B(net947),
    .Y(_2495_));
 sg13g2_a21oi_1 _5691_ (.A1(net1075),
    .A2(net947),
    .Y(_0250_),
    .B1(_2495_));
 sg13g2_nor2_1 _5692_ (.A(net1424),
    .B(net949),
    .Y(_2496_));
 sg13g2_a21oi_1 _5693_ (.A1(net1072),
    .A2(net949),
    .Y(_0251_),
    .B1(_2496_));
 sg13g2_nand3_1 _5694_ (.B(_0813_),
    .C(_2451_),
    .A(_0800_),
    .Y(_2497_));
 sg13g2_nor2_2 _5695_ (.A(_2249_),
    .B(_2497_),
    .Y(_2498_));
 sg13g2_nor2_1 _5696_ (.A(net1504),
    .B(net939),
    .Y(_2499_));
 sg13g2_a21oi_1 _5697_ (.A1(net1130),
    .A2(net939),
    .Y(_0252_),
    .B1(_2499_));
 sg13g2_nor2_1 _5698_ (.A(net1513),
    .B(net941),
    .Y(_2500_));
 sg13g2_a21oi_1 _5699_ (.A1(net1128),
    .A2(net942),
    .Y(_0253_),
    .B1(_2500_));
 sg13g2_nor2_1 _5700_ (.A(net1403),
    .B(net942),
    .Y(_2501_));
 sg13g2_a21oi_1 _5701_ (.A1(net1123),
    .A2(net942),
    .Y(_0254_),
    .B1(_2501_));
 sg13g2_nor2_1 _5702_ (.A(net1576),
    .B(net943),
    .Y(_2502_));
 sg13g2_a21oi_1 _5703_ (.A1(net1120),
    .A2(net943),
    .Y(_0255_),
    .B1(_2502_));
 sg13g2_nor2_1 _5704_ (.A(net1551),
    .B(net942),
    .Y(_2503_));
 sg13g2_a21oi_1 _5705_ (.A1(net1117),
    .A2(net942),
    .Y(_0256_),
    .B1(_2503_));
 sg13g2_nor2_1 _5706_ (.A(net1487),
    .B(net938),
    .Y(_2504_));
 sg13g2_a21oi_1 _5707_ (.A1(net1114),
    .A2(net938),
    .Y(_0257_),
    .B1(_2504_));
 sg13g2_nor2_1 _5708_ (.A(net1497),
    .B(net941),
    .Y(_2505_));
 sg13g2_a21oi_1 _5709_ (.A1(net1113),
    .A2(net943),
    .Y(_0258_),
    .B1(_2505_));
 sg13g2_nor2_1 _5710_ (.A(net1422),
    .B(net939),
    .Y(_2506_));
 sg13g2_a21oi_1 _5711_ (.A1(net1110),
    .A2(net939),
    .Y(_0259_),
    .B1(_2506_));
 sg13g2_nor2_1 _5712_ (.A(net1418),
    .B(net943),
    .Y(_2507_));
 sg13g2_a21oi_1 _5713_ (.A1(net1105),
    .A2(net943),
    .Y(_0260_),
    .B1(_2507_));
 sg13g2_nor2_1 _5714_ (.A(net1558),
    .B(net943),
    .Y(_2508_));
 sg13g2_a21oi_1 _5715_ (.A1(net1104),
    .A2(net943),
    .Y(_0261_),
    .B1(_2508_));
 sg13g2_nor2_1 _5716_ (.A(net1451),
    .B(net938),
    .Y(_2509_));
 sg13g2_a21oi_1 _5717_ (.A1(net1099),
    .A2(net938),
    .Y(_0262_),
    .B1(_2509_));
 sg13g2_nor2_1 _5718_ (.A(net1512),
    .B(net940),
    .Y(_2510_));
 sg13g2_a21oi_1 _5719_ (.A1(net1096),
    .A2(net940),
    .Y(_0263_),
    .B1(_2510_));
 sg13g2_nor2_1 _5720_ (.A(net1455),
    .B(net941),
    .Y(_2511_));
 sg13g2_a21oi_1 _5721_ (.A1(net1092),
    .A2(net941),
    .Y(_0264_),
    .B1(_2511_));
 sg13g2_nor2_1 _5722_ (.A(net1528),
    .B(net941),
    .Y(_2512_));
 sg13g2_a21oi_1 _5723_ (.A1(net1091),
    .A2(net941),
    .Y(_0265_),
    .B1(_2512_));
 sg13g2_nor2_1 _5724_ (.A(net1450),
    .B(net938),
    .Y(_2513_));
 sg13g2_a21oi_1 _5725_ (.A1(net1086),
    .A2(net938),
    .Y(_0266_),
    .B1(_2513_));
 sg13g2_nor2_1 _5726_ (.A(net1484),
    .B(net938),
    .Y(_2514_));
 sg13g2_a21oi_1 _5727_ (.A1(net1084),
    .A2(net938),
    .Y(_0267_),
    .B1(_2514_));
 sg13g2_nor2_1 _5728_ (.A(net1437),
    .B(net939),
    .Y(_2515_));
 sg13g2_a21oi_1 _5729_ (.A1(net1082),
    .A2(net939),
    .Y(_0268_),
    .B1(_2515_));
 sg13g2_nor2_1 _5730_ (.A(net1440),
    .B(net939),
    .Y(_2516_));
 sg13g2_a21oi_1 _5731_ (.A1(net1077),
    .A2(net940),
    .Y(_0269_),
    .B1(_2516_));
 sg13g2_nor2_1 _5732_ (.A(net1456),
    .B(net941),
    .Y(_2517_));
 sg13g2_a21oi_1 _5733_ (.A1(net1074),
    .A2(net941),
    .Y(_0270_),
    .B1(_2517_));
 sg13g2_nor2_1 _5734_ (.A(net1574),
    .B(net940),
    .Y(_2518_));
 sg13g2_a21oi_1 _5735_ (.A1(net1071),
    .A2(net940),
    .Y(_0271_),
    .B1(_2518_));
 sg13g2_nand2b_1 _5736_ (.Y(_2519_),
    .B(_2451_),
    .A_N(_2248_));
 sg13g2_or2_1 _5737_ (.X(_2520_),
    .B(_2519_),
    .A(_2249_));
 sg13g2_nand2_1 _5738_ (.Y(_2521_),
    .A(net762),
    .B(net934));
 sg13g2_o21ai_1 _5739_ (.B1(_2521_),
    .Y(_0272_),
    .A1(net1130),
    .A2(net934));
 sg13g2_nand2_1 _5740_ (.Y(_2522_),
    .A(net758),
    .B(net936));
 sg13g2_o21ai_1 _5741_ (.B1(_2522_),
    .Y(_0273_),
    .A1(net1126),
    .A2(net936));
 sg13g2_nand2_1 _5742_ (.Y(_2523_),
    .A(net741),
    .B(net936));
 sg13g2_o21ai_1 _5743_ (.B1(_2523_),
    .Y(_0274_),
    .A1(net1124),
    .A2(net937));
 sg13g2_nand2_1 _5744_ (.Y(_2524_),
    .A(net1316),
    .B(net936));
 sg13g2_o21ai_1 _5745_ (.B1(_2524_),
    .Y(_0275_),
    .A1(net1120),
    .A2(net935));
 sg13g2_nand2_1 _5746_ (.Y(_2525_),
    .A(net1317),
    .B(net935));
 sg13g2_o21ai_1 _5747_ (.B1(_2525_),
    .Y(_0276_),
    .A1(net1118),
    .A2(net935));
 sg13g2_nand2_1 _5748_ (.Y(_2526_),
    .A(net1343),
    .B(net932));
 sg13g2_o21ai_1 _5749_ (.B1(_2526_),
    .Y(_0277_),
    .A1(net1115),
    .A2(net932));
 sg13g2_nand2_1 _5750_ (.Y(_2527_),
    .A(net1355),
    .B(net936));
 sg13g2_o21ai_1 _5751_ (.B1(_2527_),
    .Y(_0278_),
    .A1(net1112),
    .A2(net936));
 sg13g2_nand2_1 _5752_ (.Y(_2528_),
    .A(net1342),
    .B(net933));
 sg13g2_o21ai_1 _5753_ (.B1(_2528_),
    .Y(_0279_),
    .A1(net1108),
    .A2(net933));
 sg13g2_nand2_1 _5754_ (.Y(_2529_),
    .A(net829),
    .B(net935));
 sg13g2_o21ai_1 _5755_ (.B1(_2529_),
    .Y(_0280_),
    .A1(net1106),
    .A2(net935));
 sg13g2_nand2_1 _5756_ (.Y(_2530_),
    .A(net694),
    .B(net937));
 sg13g2_o21ai_1 _5757_ (.B1(_2530_),
    .Y(_0281_),
    .A1(net1104),
    .A2(net937));
 sg13g2_nand2_1 _5758_ (.Y(_2531_),
    .A(net1270),
    .B(net932));
 sg13g2_o21ai_1 _5759_ (.B1(_2531_),
    .Y(_0282_),
    .A1(net1099),
    .A2(net932));
 sg13g2_nand2_1 _5760_ (.Y(_2532_),
    .A(net1323),
    .B(net934));
 sg13g2_o21ai_1 _5761_ (.B1(_2532_),
    .Y(_0283_),
    .A1(net1096),
    .A2(net934));
 sg13g2_nand2_1 _5762_ (.Y(_2533_),
    .A(net1341),
    .B(net935));
 sg13g2_o21ai_1 _5763_ (.B1(_2533_),
    .Y(_0284_),
    .A1(net1093),
    .A2(net936));
 sg13g2_nand2_1 _5764_ (.Y(_2534_),
    .A(net771),
    .B(net937));
 sg13g2_o21ai_1 _5765_ (.B1(_2534_),
    .Y(_0285_),
    .A1(net1089),
    .A2(net937));
 sg13g2_nand2_1 _5766_ (.Y(_2535_),
    .A(net687),
    .B(net932));
 sg13g2_o21ai_1 _5767_ (.B1(_2535_),
    .Y(_0286_),
    .A1(net1086),
    .A2(net932));
 sg13g2_nand2_1 _5768_ (.Y(_2536_),
    .A(net747),
    .B(net932));
 sg13g2_o21ai_1 _5769_ (.B1(_2536_),
    .Y(_0287_),
    .A1(net1083),
    .A2(net932));
 sg13g2_nand2_1 _5770_ (.Y(_2537_),
    .A(net1359),
    .B(net933));
 sg13g2_o21ai_1 _5771_ (.B1(_2537_),
    .Y(_0288_),
    .A1(net1080),
    .A2(net933));
 sg13g2_nand2_1 _5772_ (.Y(_2538_),
    .A(net1252),
    .B(net933));
 sg13g2_o21ai_1 _5773_ (.B1(_2538_),
    .Y(_0289_),
    .A1(net1077),
    .A2(net933));
 sg13g2_nand2_1 _5774_ (.Y(_2539_),
    .A(net1366),
    .B(net935));
 sg13g2_o21ai_1 _5775_ (.B1(_2539_),
    .Y(_0290_),
    .A1(net1074),
    .A2(net935));
 sg13g2_nand2_1 _5776_ (.Y(_2540_),
    .A(net674),
    .B(net937));
 sg13g2_o21ai_1 _5777_ (.B1(_2540_),
    .Y(_0291_),
    .A1(net1072),
    .A2(net937));
 sg13g2_nand2b_2 _5778_ (.Y(_2541_),
    .B(_0767_),
    .A_N(_0785_));
 sg13g2_or2_1 _5779_ (.X(_2542_),
    .B(_2541_),
    .A(_2452_));
 sg13g2_nand2_1 _5780_ (.Y(_2543_),
    .A(net751),
    .B(net926));
 sg13g2_o21ai_1 _5781_ (.B1(_2543_),
    .Y(_0292_),
    .A1(net1131),
    .A2(net926));
 sg13g2_nand2_1 _5782_ (.Y(_2544_),
    .A(net669),
    .B(net930));
 sg13g2_o21ai_1 _5783_ (.B1(_2544_),
    .Y(_0293_),
    .A1(net1126),
    .A2(net930));
 sg13g2_nand2_1 _5784_ (.Y(_2545_),
    .A(net724),
    .B(net930));
 sg13g2_o21ai_1 _5785_ (.B1(_2545_),
    .Y(_0294_),
    .A1(net1123),
    .A2(net930));
 sg13g2_nand2_1 _5786_ (.Y(_2546_),
    .A(net1276),
    .B(net931));
 sg13g2_o21ai_1 _5787_ (.B1(_2546_),
    .Y(_0295_),
    .A1(net1121),
    .A2(net931));
 sg13g2_nand2_1 _5788_ (.Y(_2547_),
    .A(net682),
    .B(net931));
 sg13g2_o21ai_1 _5789_ (.B1(_2547_),
    .Y(_0296_),
    .A1(net1117),
    .A2(net930));
 sg13g2_nand2_1 _5790_ (.Y(_2548_),
    .A(net760),
    .B(net927));
 sg13g2_o21ai_1 _5791_ (.B1(_2548_),
    .Y(_0297_),
    .A1(net1116),
    .A2(net927));
 sg13g2_nand2_1 _5792_ (.Y(_2549_),
    .A(net730),
    .B(net928));
 sg13g2_o21ai_1 _5793_ (.B1(_2549_),
    .Y(_0298_),
    .A1(net1111),
    .A2(net928));
 sg13g2_nand2_1 _5794_ (.Y(_2550_),
    .A(net736),
    .B(net927));
 sg13g2_o21ai_1 _5795_ (.B1(_2550_),
    .Y(_0299_),
    .A1(net1110),
    .A2(net927));
 sg13g2_nand2_1 _5796_ (.Y(_2551_),
    .A(net1318),
    .B(net929));
 sg13g2_o21ai_1 _5797_ (.B1(_2551_),
    .Y(_0300_),
    .A1(net1105),
    .A2(net929));
 sg13g2_nand2_1 _5798_ (.Y(_2552_),
    .A(net1248),
    .B(net929));
 sg13g2_o21ai_1 _5799_ (.B1(_2552_),
    .Y(_0301_),
    .A1(net1102),
    .A2(net929));
 sg13g2_nand2_1 _5800_ (.Y(_2553_),
    .A(net740),
    .B(net925));
 sg13g2_o21ai_1 _5801_ (.B1(_2553_),
    .Y(_0302_),
    .A1(net1100),
    .A2(net925));
 sg13g2_nand2_1 _5802_ (.Y(_2554_),
    .A(net703),
    .B(net925));
 sg13g2_o21ai_1 _5803_ (.B1(_2554_),
    .Y(_0303_),
    .A1(net1097),
    .A2(net925));
 sg13g2_nand2_1 _5804_ (.Y(_2555_),
    .A(net776),
    .B(net929));
 sg13g2_o21ai_1 _5805_ (.B1(_2555_),
    .Y(_0304_),
    .A1(net1093),
    .A2(net930));
 sg13g2_nand2_1 _5806_ (.Y(_2556_),
    .A(net727),
    .B(net929));
 sg13g2_o21ai_1 _5807_ (.B1(_2556_),
    .Y(_0305_),
    .A1(net1089),
    .A2(net929));
 sg13g2_nand2_1 _5808_ (.Y(_2557_),
    .A(net702),
    .B(net925));
 sg13g2_o21ai_1 _5809_ (.B1(_2557_),
    .Y(_0306_),
    .A1(net1087),
    .A2(net925));
 sg13g2_nand2_1 _5810_ (.Y(_2558_),
    .A(net1256),
    .B(net925));
 sg13g2_o21ai_1 _5811_ (.B1(_2558_),
    .Y(_0307_),
    .A1(net1085),
    .A2(net925));
 sg13g2_nand2_1 _5812_ (.Y(_2559_),
    .A(net790),
    .B(net927));
 sg13g2_o21ai_1 _5813_ (.B1(_2559_),
    .Y(_0308_),
    .A1(net1081),
    .A2(net927));
 sg13g2_nand2_1 _5814_ (.Y(_2560_),
    .A(net654),
    .B(net927));
 sg13g2_o21ai_1 _5815_ (.B1(_2560_),
    .Y(_0309_),
    .A1(net1078),
    .A2(net927));
 sg13g2_nand2_1 _5816_ (.Y(_2561_),
    .A(net733),
    .B(net930));
 sg13g2_o21ai_1 _5817_ (.B1(_2561_),
    .Y(_0310_),
    .A1(net1076),
    .A2(net929));
 sg13g2_nand2_1 _5818_ (.Y(_2562_),
    .A(net759),
    .B(net926));
 sg13g2_o21ai_1 _5819_ (.B1(_2562_),
    .Y(_0311_),
    .A1(net1071),
    .A2(net926));
 sg13g2_or2_1 _5820_ (.X(_2563_),
    .B(_2541_),
    .A(_2475_));
 sg13g2_nand2_1 _5821_ (.Y(_2564_),
    .A(net718),
    .B(net919));
 sg13g2_o21ai_1 _5822_ (.B1(_2564_),
    .Y(_0312_),
    .A1(net1130),
    .A2(net919));
 sg13g2_nand2_1 _5823_ (.Y(_2565_),
    .A(net1333),
    .B(net923));
 sg13g2_o21ai_1 _5824_ (.B1(_2565_),
    .Y(_0313_),
    .A1(net1126),
    .A2(net923));
 sg13g2_nand2_1 _5825_ (.Y(_2566_),
    .A(net686),
    .B(net923));
 sg13g2_o21ai_1 _5826_ (.B1(_2566_),
    .Y(_0314_),
    .A1(net1124),
    .A2(net923));
 sg13g2_nand2_1 _5827_ (.Y(_2567_),
    .A(net661),
    .B(net924));
 sg13g2_o21ai_1 _5828_ (.B1(_2567_),
    .Y(_0315_),
    .A1(net1120),
    .A2(net924));
 sg13g2_nand2_1 _5829_ (.Y(_2568_),
    .A(net1281),
    .B(net924));
 sg13g2_o21ai_1 _5830_ (.B1(_2568_),
    .Y(_0316_),
    .A1(net1117),
    .A2(net924));
 sg13g2_nand2_1 _5831_ (.Y(_2569_),
    .A(net715),
    .B(net920));
 sg13g2_o21ai_1 _5832_ (.B1(_2569_),
    .Y(_0317_),
    .A1(net1114),
    .A2(net920));
 sg13g2_nand2_1 _5833_ (.Y(_2570_),
    .A(net1289),
    .B(net921));
 sg13g2_o21ai_1 _5834_ (.B1(_2570_),
    .Y(_0318_),
    .A1(net1111),
    .A2(net921));
 sg13g2_nand2_1 _5835_ (.Y(_2571_),
    .A(net1297),
    .B(net920));
 sg13g2_o21ai_1 _5836_ (.B1(_2571_),
    .Y(_0319_),
    .A1(net1110),
    .A2(net920));
 sg13g2_nand2_1 _5837_ (.Y(_2572_),
    .A(net1268),
    .B(net922));
 sg13g2_o21ai_1 _5838_ (.B1(_2572_),
    .Y(_0320_),
    .A1(net1105),
    .A2(net922));
 sg13g2_nand2_1 _5839_ (.Y(_2573_),
    .A(net1329),
    .B(net922));
 sg13g2_o21ai_1 _5840_ (.B1(_2573_),
    .Y(_0321_),
    .A1(net1103),
    .A2(net922));
 sg13g2_nand2_1 _5841_ (.Y(_2574_),
    .A(net651),
    .B(net919));
 sg13g2_o21ai_1 _5842_ (.B1(_2574_),
    .Y(_0322_),
    .A1(net1101),
    .A2(net919));
 sg13g2_nand2_1 _5843_ (.Y(_2575_),
    .A(net816),
    .B(net921));
 sg13g2_o21ai_1 _5844_ (.B1(_2575_),
    .Y(_0323_),
    .A1(net1096),
    .A2(net921));
 sg13g2_nand2_1 _5845_ (.Y(_2576_),
    .A(net1299),
    .B(net923));
 sg13g2_o21ai_1 _5846_ (.B1(_2576_),
    .Y(_0324_),
    .A1(net1095),
    .A2(net923));
 sg13g2_nand2_1 _5847_ (.Y(_2577_),
    .A(net1309),
    .B(net922));
 sg13g2_o21ai_1 _5848_ (.B1(_2577_),
    .Y(_0325_),
    .A1(net1089),
    .A2(net922));
 sg13g2_nand2_1 _5849_ (.Y(_2578_),
    .A(net815),
    .B(net919));
 sg13g2_o21ai_1 _5850_ (.B1(_2578_),
    .Y(_0326_),
    .A1(net1088),
    .A2(net919));
 sg13g2_nand2_1 _5851_ (.Y(_2579_),
    .A(net1247),
    .B(net919));
 sg13g2_o21ai_1 _5852_ (.B1(_2579_),
    .Y(_0327_),
    .A1(net1085),
    .A2(net919));
 sg13g2_nand2_1 _5853_ (.Y(_2580_),
    .A(net1378),
    .B(net920));
 sg13g2_o21ai_1 _5854_ (.B1(_2580_),
    .Y(_0328_),
    .A1(net1081),
    .A2(net920));
 sg13g2_nand2_1 _5855_ (.Y(_2581_),
    .A(net797),
    .B(net920));
 sg13g2_o21ai_1 _5856_ (.B1(_2581_),
    .Y(_0329_),
    .A1(net1077),
    .A2(net920));
 sg13g2_nand2_1 _5857_ (.Y(_2582_),
    .A(net1312),
    .B(net923));
 sg13g2_o21ai_1 _5858_ (.B1(_2582_),
    .Y(_0330_),
    .A1(net1075),
    .A2(net923));
 sg13g2_nand2_1 _5859_ (.Y(_2583_),
    .A(net783),
    .B(net922));
 sg13g2_o21ai_1 _5860_ (.B1(_2583_),
    .Y(_0331_),
    .A1(net1073),
    .A2(net922));
 sg13g2_or2_1 _5861_ (.X(_2584_),
    .B(_2541_),
    .A(_2497_));
 sg13g2_nand2_1 _5862_ (.Y(_2585_),
    .A(net742),
    .B(net915));
 sg13g2_o21ai_1 _5863_ (.B1(_2585_),
    .Y(_0332_),
    .A1(net1131),
    .A2(net915));
 sg13g2_nand2_1 _5864_ (.Y(_2586_),
    .A(net820),
    .B(net916));
 sg13g2_o21ai_1 _5865_ (.B1(_2586_),
    .Y(_0333_),
    .A1(net1126),
    .A2(net916));
 sg13g2_nand2_1 _5866_ (.Y(_2587_),
    .A(net808),
    .B(net916));
 sg13g2_o21ai_1 _5867_ (.B1(_2587_),
    .Y(_0334_),
    .A1(net1124),
    .A2(net916));
 sg13g2_nand2_1 _5868_ (.Y(_2588_),
    .A(net1348),
    .B(net916));
 sg13g2_o21ai_1 _5869_ (.B1(_2588_),
    .Y(_0335_),
    .A1(net1121),
    .A2(net916));
 sg13g2_nand2_1 _5870_ (.Y(_2589_),
    .A(net752),
    .B(net918));
 sg13g2_o21ai_1 _5871_ (.B1(_2589_),
    .Y(_0336_),
    .A1(net1118),
    .A2(net918));
 sg13g2_nand2_1 _5872_ (.Y(_2590_),
    .A(net745),
    .B(net913));
 sg13g2_o21ai_1 _5873_ (.B1(_2590_),
    .Y(_0337_),
    .A1(net1116),
    .A2(net913));
 sg13g2_nand2_1 _5874_ (.Y(_2591_),
    .A(net1262),
    .B(net916));
 sg13g2_o21ai_1 _5875_ (.B1(_2591_),
    .Y(_0338_),
    .A1(net1112),
    .A2(net916));
 sg13g2_nand2_1 _5876_ (.Y(_2592_),
    .A(net830),
    .B(net914));
 sg13g2_o21ai_1 _5877_ (.B1(_2592_),
    .Y(_0339_),
    .A1(net1108),
    .A2(net914));
 sg13g2_nand2_1 _5878_ (.Y(_2593_),
    .A(net809),
    .B(net917));
 sg13g2_o21ai_1 _5879_ (.B1(_2593_),
    .Y(_0340_),
    .A1(net1105),
    .A2(net918));
 sg13g2_nand2_1 _5880_ (.Y(_2594_),
    .A(net708),
    .B(net918));
 sg13g2_o21ai_1 _5881_ (.B1(_2594_),
    .Y(_0341_),
    .A1(net1102),
    .A2(net918));
 sg13g2_nand2_1 _5882_ (.Y(_2595_),
    .A(net657),
    .B(net913));
 sg13g2_o21ai_1 _5883_ (.B1(_2595_),
    .Y(_0342_),
    .A1(net1099),
    .A2(net913));
 sg13g2_nand2_1 _5884_ (.Y(_2596_),
    .A(net834),
    .B(net915));
 sg13g2_o21ai_1 _5885_ (.B1(_2596_),
    .Y(_0343_),
    .A1(net1098),
    .A2(net915));
 sg13g2_nand2_1 _5886_ (.Y(_2597_),
    .A(net665),
    .B(net917));
 sg13g2_o21ai_1 _5887_ (.B1(_2597_),
    .Y(_0344_),
    .A1(net1093),
    .A2(net917));
 sg13g2_nand2_1 _5888_ (.Y(_2598_),
    .A(net794),
    .B(net917));
 sg13g2_o21ai_1 _5889_ (.B1(_2598_),
    .Y(_0345_),
    .A1(net1091),
    .A2(net917));
 sg13g2_nand2_1 _5890_ (.Y(_2599_),
    .A(net764),
    .B(net913));
 sg13g2_o21ai_1 _5891_ (.B1(_2599_),
    .Y(_0346_),
    .A1(net1087),
    .A2(net913));
 sg13g2_nand2_1 _5892_ (.Y(_2600_),
    .A(net827),
    .B(net913));
 sg13g2_o21ai_1 _5893_ (.B1(_2600_),
    .Y(_0347_),
    .A1(net1083),
    .A2(net913));
 sg13g2_nand2_1 _5894_ (.Y(_2601_),
    .A(net655),
    .B(net914));
 sg13g2_o21ai_1 _5895_ (.B1(_2601_),
    .Y(_0348_),
    .A1(net1082),
    .A2(net914));
 sg13g2_nand2_1 _5896_ (.Y(_2602_),
    .A(net789),
    .B(net914));
 sg13g2_o21ai_1 _5897_ (.B1(_2602_),
    .Y(_0349_),
    .A1(net1078),
    .A2(net914));
 sg13g2_nand2_1 _5898_ (.Y(_2603_),
    .A(net1291),
    .B(net917));
 sg13g2_o21ai_1 _5899_ (.B1(_2603_),
    .Y(_0350_),
    .A1(net1074),
    .A2(net917));
 sg13g2_nand2_1 _5900_ (.Y(_2604_),
    .A(net810),
    .B(net915));
 sg13g2_o21ai_1 _5901_ (.B1(_2604_),
    .Y(_0351_),
    .A1(net1071),
    .A2(net915));
 sg13g2_or2_1 _5902_ (.X(_2605_),
    .B(_2541_),
    .A(_2519_));
 sg13g2_nand2_1 _5903_ (.Y(_2606_),
    .A(net802),
    .B(net909));
 sg13g2_o21ai_1 _5904_ (.B1(_2606_),
    .Y(_0352_),
    .A1(net1131),
    .A2(net909));
 sg13g2_nand2_1 _5905_ (.Y(_2607_),
    .A(net766),
    .B(net911));
 sg13g2_o21ai_1 _5906_ (.B1(_2607_),
    .Y(_0353_),
    .A1(net1127),
    .A2(net911));
 sg13g2_nand2_1 _5907_ (.Y(_2608_),
    .A(net793),
    .B(net912));
 sg13g2_o21ai_1 _5908_ (.B1(_2608_),
    .Y(_0354_),
    .A1(net1124),
    .A2(net912));
 sg13g2_nand2_1 _5909_ (.Y(_2609_),
    .A(net1251),
    .B(net912));
 sg13g2_o21ai_1 _5910_ (.B1(_2609_),
    .Y(_0355_),
    .A1(net1121),
    .A2(net910));
 sg13g2_nand2_1 _5911_ (.Y(_2610_),
    .A(net1319),
    .B(net911));
 sg13g2_o21ai_1 _5912_ (.B1(_2610_),
    .Y(_0356_),
    .A1(net1118),
    .A2(net911));
 sg13g2_nand2_1 _5913_ (.Y(_2611_),
    .A(net668),
    .B(net907));
 sg13g2_o21ai_1 _5914_ (.B1(_2611_),
    .Y(_0357_),
    .A1(net1115),
    .A2(net907));
 sg13g2_nand2_1 _5915_ (.Y(_2612_),
    .A(net788),
    .B(net912));
 sg13g2_o21ai_1 _5916_ (.B1(_2612_),
    .Y(_0358_),
    .A1(net1113),
    .A2(net910));
 sg13g2_nand2_1 _5917_ (.Y(_2613_),
    .A(net821),
    .B(net908));
 sg13g2_o21ai_1 _5918_ (.B1(_2613_),
    .Y(_0359_),
    .A1(net1109),
    .A2(net908));
 sg13g2_nand2_1 _5919_ (.Y(_2614_),
    .A(net1290),
    .B(net910));
 sg13g2_o21ai_1 _5920_ (.B1(_2614_),
    .Y(_0360_),
    .A1(net1106),
    .A2(net910));
 sg13g2_nand2_1 _5921_ (.Y(_2615_),
    .A(net1258),
    .B(net910));
 sg13g2_o21ai_1 _5922_ (.B1(_2615_),
    .Y(_0361_),
    .A1(net1104),
    .A2(net910));
 sg13g2_nand2_1 _5923_ (.Y(_2616_),
    .A(net688),
    .B(net907));
 sg13g2_o21ai_1 _5924_ (.B1(_2616_),
    .Y(_0362_),
    .A1(net1099),
    .A2(net907));
 sg13g2_nand2_1 _5925_ (.Y(_2617_),
    .A(net756),
    .B(net909));
 sg13g2_o21ai_1 _5926_ (.B1(_2617_),
    .Y(_0363_),
    .A1(net1098),
    .A2(net909));
 sg13g2_nand2_1 _5927_ (.Y(_2618_),
    .A(net1344),
    .B(net911));
 sg13g2_o21ai_1 _5928_ (.B1(_2618_),
    .Y(_0364_),
    .A1(net1092),
    .A2(net911));
 sg13g2_nand2_1 _5929_ (.Y(_2619_),
    .A(net667),
    .B(net910));
 sg13g2_o21ai_1 _5930_ (.B1(_2619_),
    .Y(_0365_),
    .A1(net1090),
    .A2(net910));
 sg13g2_nand2_1 _5931_ (.Y(_2620_),
    .A(net695),
    .B(net907));
 sg13g2_o21ai_1 _5932_ (.B1(_2620_),
    .Y(_0366_),
    .A1(net1087),
    .A2(net907));
 sg13g2_nand2_1 _5933_ (.Y(_2621_),
    .A(net707),
    .B(net907));
 sg13g2_o21ai_1 _5934_ (.B1(_2621_),
    .Y(_0367_),
    .A1(net1084),
    .A2(net907));
 sg13g2_nand2_1 _5935_ (.Y(_2622_),
    .A(net1338),
    .B(net908));
 sg13g2_o21ai_1 _5936_ (.B1(_2622_),
    .Y(_0368_),
    .A1(net1080),
    .A2(net908));
 sg13g2_nand2_1 _5937_ (.Y(_2623_),
    .A(net666),
    .B(net908));
 sg13g2_o21ai_1 _5938_ (.B1(_2623_),
    .Y(_0369_),
    .A1(net1078),
    .A2(net908));
 sg13g2_nand2_1 _5939_ (.Y(_2624_),
    .A(net1307),
    .B(net911));
 sg13g2_o21ai_1 _5940_ (.B1(_2624_),
    .Y(_0370_),
    .A1(net1074),
    .A2(net911));
 sg13g2_nand2_1 _5941_ (.Y(_2625_),
    .A(net824),
    .B(net909));
 sg13g2_o21ai_1 _5942_ (.B1(_2625_),
    .Y(_0371_),
    .A1(net1073),
    .A2(net909));
 sg13g2_nand2b_1 _5943_ (.Y(_2626_),
    .B(_0785_),
    .A_N(_0767_));
 sg13g2_or2_1 _5944_ (.X(_2627_),
    .B(_2626_),
    .A(_2452_));
 sg13g2_nand2_1 _5945_ (.Y(_2628_),
    .A(net696),
    .B(net902));
 sg13g2_o21ai_1 _5946_ (.B1(_2628_),
    .Y(_0372_),
    .A1(net1132),
    .A2(net902));
 sg13g2_nand2_1 _5947_ (.Y(_2629_),
    .A(net1340),
    .B(net904));
 sg13g2_o21ai_1 _5948_ (.B1(_2629_),
    .Y(_0373_),
    .A1(net1126),
    .A2(net904));
 sg13g2_nand2_1 _5949_ (.Y(_2630_),
    .A(net1260),
    .B(net904));
 sg13g2_o21ai_1 _5950_ (.B1(_2630_),
    .Y(_0374_),
    .A1(net1125),
    .A2(net904));
 sg13g2_nand2_1 _5951_ (.Y(_2631_),
    .A(net1304),
    .B(net905));
 sg13g2_o21ai_1 _5952_ (.B1(_2631_),
    .Y(_0375_),
    .A1(net1120),
    .A2(net905));
 sg13g2_nand2_1 _5953_ (.Y(_2632_),
    .A(net692),
    .B(net903));
 sg13g2_o21ai_1 _5954_ (.B1(_2632_),
    .Y(_0376_),
    .A1(net1117),
    .A2(net903));
 sg13g2_nand2_1 _5955_ (.Y(_2633_),
    .A(net1255),
    .B(net901));
 sg13g2_o21ai_1 _5956_ (.B1(_2633_),
    .Y(_0377_),
    .A1(net1114),
    .A2(net901));
 sg13g2_nand2_1 _5957_ (.Y(_2634_),
    .A(net782),
    .B(net904));
 sg13g2_o21ai_1 _5958_ (.B1(_2634_),
    .Y(_0378_),
    .A1(net1113),
    .A2(net904));
 sg13g2_nand2_1 _5959_ (.Y(_2635_),
    .A(net662),
    .B(net902));
 sg13g2_o21ai_1 _5960_ (.B1(_2635_),
    .Y(_0379_),
    .A1(net1108),
    .A2(net902));
 sg13g2_nand2_1 _5961_ (.Y(_2636_),
    .A(net709),
    .B(net903));
 sg13g2_o21ai_1 _5962_ (.B1(_2636_),
    .Y(_0380_),
    .A1(net1106),
    .A2(net903));
 sg13g2_nand2_1 _5963_ (.Y(_2637_),
    .A(net693),
    .B(net905));
 sg13g2_o21ai_1 _5964_ (.B1(_2637_),
    .Y(_0381_),
    .A1(net1102),
    .A2(net905));
 sg13g2_nand2_1 _5965_ (.Y(_2638_),
    .A(net1282),
    .B(net902));
 sg13g2_o21ai_1 _5966_ (.B1(_2638_),
    .Y(_0382_),
    .A1(net1101),
    .A2(net906));
 sg13g2_nand2_1 _5967_ (.Y(_2639_),
    .A(net676),
    .B(net902));
 sg13g2_o21ai_1 _5968_ (.B1(_2639_),
    .Y(_0383_),
    .A1(net1096),
    .A2(net902));
 sg13g2_nand2_1 _5969_ (.Y(_2640_),
    .A(net1372),
    .B(net903));
 sg13g2_o21ai_1 _5970_ (.B1(_2640_),
    .Y(_0384_),
    .A1(net1092),
    .A2(net903));
 sg13g2_nand2_1 _5971_ (.Y(_2641_),
    .A(net701),
    .B(net905));
 sg13g2_o21ai_1 _5972_ (.B1(_2641_),
    .Y(_0385_),
    .A1(net1089),
    .A2(net905));
 sg13g2_nand2_1 _5973_ (.Y(_2642_),
    .A(net1356),
    .B(net901));
 sg13g2_o21ai_1 _5974_ (.B1(_2642_),
    .Y(_0386_),
    .A1(net1086),
    .A2(net901));
 sg13g2_nand2_1 _5975_ (.Y(_2643_),
    .A(net1286),
    .B(net901));
 sg13g2_o21ai_1 _5976_ (.B1(_2643_),
    .Y(_0387_),
    .A1(net1083),
    .A2(net901));
 sg13g2_nand2_1 _5977_ (.Y(_2644_),
    .A(net746),
    .B(net901));
 sg13g2_o21ai_1 _5978_ (.B1(_2644_),
    .Y(_0388_),
    .A1(net1080),
    .A2(net901));
 sg13g2_nand2_1 _5979_ (.Y(_2645_),
    .A(net1259),
    .B(net906));
 sg13g2_o21ai_1 _5980_ (.B1(_2645_),
    .Y(_0389_),
    .A1(net1078),
    .A2(net906));
 sg13g2_nand2_1 _5981_ (.Y(_2646_),
    .A(net819),
    .B(net903));
 sg13g2_o21ai_1 _5982_ (.B1(_2646_),
    .Y(_0390_),
    .A1(net1075),
    .A2(net903));
 sg13g2_nand2_1 _5983_ (.Y(_2647_),
    .A(net761),
    .B(net905));
 sg13g2_o21ai_1 _5984_ (.B1(_2647_),
    .Y(_0391_),
    .A1(net1071),
    .A2(net905));
 sg13g2_or2_1 _5985_ (.X(_2648_),
    .B(_2626_),
    .A(_2475_));
 sg13g2_nand2_1 _5986_ (.Y(_2649_),
    .A(net798),
    .B(net897));
 sg13g2_o21ai_1 _5987_ (.B1(_2649_),
    .Y(_0392_),
    .A1(net1132),
    .A2(net897));
 sg13g2_nand2_1 _5988_ (.Y(_2650_),
    .A(net769),
    .B(net898));
 sg13g2_o21ai_1 _5989_ (.B1(_2650_),
    .Y(_0393_),
    .A1(net1129),
    .A2(net898));
 sg13g2_nand2_1 _5990_ (.Y(_2651_),
    .A(net1283),
    .B(net898));
 sg13g2_o21ai_1 _5991_ (.B1(_2651_),
    .Y(_0394_),
    .A1(net1124),
    .A2(net898));
 sg13g2_nand2_1 _5992_ (.Y(_2652_),
    .A(net710),
    .B(net898));
 sg13g2_o21ai_1 _5993_ (.B1(_2652_),
    .Y(_0395_),
    .A1(net1122),
    .A2(net898));
 sg13g2_nand2_1 _5994_ (.Y(_2653_),
    .A(net1325),
    .B(net900));
 sg13g2_o21ai_1 _5995_ (.B1(_2653_),
    .Y(_0396_),
    .A1(net1119),
    .A2(net899));
 sg13g2_nand2_1 _5996_ (.Y(_2654_),
    .A(net1285),
    .B(net896));
 sg13g2_o21ai_1 _5997_ (.B1(_2654_),
    .Y(_0397_),
    .A1(net1114),
    .A2(net896));
 sg13g2_nand2_1 _5998_ (.Y(_2655_),
    .A(net1313),
    .B(net900));
 sg13g2_o21ai_1 _5999_ (.B1(_2655_),
    .Y(_0398_),
    .A1(net1111),
    .A2(net900));
 sg13g2_nand2_1 _6000_ (.Y(_2656_),
    .A(net1263),
    .B(net895));
 sg13g2_o21ai_1 _6001_ (.B1(_2656_),
    .Y(_0399_),
    .A1(net1110),
    .A2(net895));
 sg13g2_nand2_1 _6002_ (.Y(_2657_),
    .A(net735),
    .B(net898));
 sg13g2_o21ai_1 _6003_ (.B1(_2657_),
    .Y(_0400_),
    .A1(net1107),
    .A2(net898));
 sg13g2_nand2_1 _6004_ (.Y(_2658_),
    .A(net750),
    .B(net900));
 sg13g2_o21ai_1 _6005_ (.B1(_2658_),
    .Y(_0401_),
    .A1(net1104),
    .A2(net900));
 sg13g2_nand2_1 _6006_ (.Y(_2659_),
    .A(net713),
    .B(net895));
 sg13g2_o21ai_1 _6007_ (.B1(_2659_),
    .Y(_0402_),
    .A1(net1099),
    .A2(net895));
 sg13g2_nand2_1 _6008_ (.Y(_2660_),
    .A(net670),
    .B(net897));
 sg13g2_o21ai_1 _6009_ (.B1(_2660_),
    .Y(_0403_),
    .A1(net1096),
    .A2(net897));
 sg13g2_nand2_1 _6010_ (.Y(_2661_),
    .A(net753),
    .B(net899));
 sg13g2_o21ai_1 _6011_ (.B1(_2661_),
    .Y(_0404_),
    .A1(net1092),
    .A2(net899));
 sg13g2_nand2_1 _6012_ (.Y(_2662_),
    .A(net823),
    .B(net899));
 sg13g2_o21ai_1 _6013_ (.B1(_2662_),
    .Y(_0405_),
    .A1(net1090),
    .A2(net899));
 sg13g2_nand2_1 _6014_ (.Y(_2663_),
    .A(net1269),
    .B(net895));
 sg13g2_o21ai_1 _6015_ (.B1(_2663_),
    .Y(_0406_),
    .A1(net1086),
    .A2(net895));
 sg13g2_nand2_1 _6016_ (.Y(_2664_),
    .A(net1363),
    .B(net895));
 sg13g2_o21ai_1 _6017_ (.B1(_2664_),
    .Y(_0407_),
    .A1(net1085),
    .A2(net895));
 sg13g2_nand2_1 _6018_ (.Y(_2665_),
    .A(net1277),
    .B(net897));
 sg13g2_o21ai_1 _6019_ (.B1(_2665_),
    .Y(_0408_),
    .A1(net1081),
    .A2(net896));
 sg13g2_nand2_1 _6020_ (.Y(_2666_),
    .A(net763),
    .B(net896));
 sg13g2_o21ai_1 _6021_ (.B1(_2666_),
    .Y(_0409_),
    .A1(net1077),
    .A2(net896));
 sg13g2_nand2_1 _6022_ (.Y(_2667_),
    .A(net739),
    .B(net899));
 sg13g2_o21ai_1 _6023_ (.B1(_2667_),
    .Y(_0410_),
    .A1(net1076),
    .A2(net899));
 sg13g2_nand2_1 _6024_ (.Y(_2668_),
    .A(net786),
    .B(net900));
 sg13g2_o21ai_1 _6025_ (.B1(_2668_),
    .Y(_0411_),
    .A1(net1071),
    .A2(net900));
 sg13g2_or2_1 _6026_ (.X(_2669_),
    .B(_2626_),
    .A(_2497_));
 sg13g2_nand2_1 _6027_ (.Y(_2670_),
    .A(net801),
    .B(net890));
 sg13g2_o21ai_1 _6028_ (.B1(_2670_),
    .Y(_0412_),
    .A1(net1131),
    .A2(net890));
 sg13g2_nand2_1 _6029_ (.Y(_2671_),
    .A(net729),
    .B(net891));
 sg13g2_o21ai_1 _6030_ (.B1(_2671_),
    .Y(_0413_),
    .A1(net1127),
    .A2(net891));
 sg13g2_nand2_1 _6031_ (.Y(_2672_),
    .A(net719),
    .B(net892));
 sg13g2_o21ai_1 _6032_ (.B1(_2672_),
    .Y(_0414_),
    .A1(net1123),
    .A2(net892));
 sg13g2_nand2_1 _6033_ (.Y(_2673_),
    .A(net714),
    .B(net893));
 sg13g2_o21ai_1 _6034_ (.B1(_2673_),
    .Y(_0415_),
    .A1(net1121),
    .A2(net893));
 sg13g2_nand2_1 _6035_ (.Y(_2674_),
    .A(net1330),
    .B(net892));
 sg13g2_o21ai_1 _6036_ (.B1(_2674_),
    .Y(_0416_),
    .A1(net1117),
    .A2(net892));
 sg13g2_nand2_1 _6037_ (.Y(_2675_),
    .A(net1284),
    .B(net889));
 sg13g2_o21ai_1 _6038_ (.B1(_2675_),
    .Y(_0417_),
    .A1(net1115),
    .A2(net889));
 sg13g2_nand2_1 _6039_ (.Y(_2676_),
    .A(net1253),
    .B(net890));
 sg13g2_o21ai_1 _6040_ (.B1(_2676_),
    .Y(_0418_),
    .A1(net1111),
    .A2(net890));
 sg13g2_nand2_1 _6041_ (.Y(_2677_),
    .A(net689),
    .B(net888));
 sg13g2_o21ai_1 _6042_ (.B1(_2677_),
    .Y(_0419_),
    .A1(net1110),
    .A2(net888));
 sg13g2_nand2_1 _6043_ (.Y(_2678_),
    .A(net1320),
    .B(net891));
 sg13g2_o21ai_1 _6044_ (.B1(_2678_),
    .Y(_0420_),
    .A1(net1105),
    .A2(net891));
 sg13g2_nand2_1 _6045_ (.Y(_2679_),
    .A(net706),
    .B(net893));
 sg13g2_o21ai_1 _6046_ (.B1(_2679_),
    .Y(_0421_),
    .A1(net1103),
    .A2(net893));
 sg13g2_nand2_1 _6047_ (.Y(_2680_),
    .A(net1275),
    .B(net890));
 sg13g2_o21ai_1 _6048_ (.B1(_2680_),
    .Y(_0422_),
    .A1(net1101),
    .A2(net894));
 sg13g2_nand2_1 _6049_ (.Y(_2681_),
    .A(net722),
    .B(net890));
 sg13g2_o21ai_1 _6050_ (.B1(_2681_),
    .Y(_0423_),
    .A1(net1098),
    .A2(net894));
 sg13g2_nand2_1 _6051_ (.Y(_2682_),
    .A(net1375),
    .B(net891));
 sg13g2_o21ai_1 _6052_ (.B1(_2682_),
    .Y(_0424_),
    .A1(net1092),
    .A2(net891));
 sg13g2_nand2_1 _6053_ (.Y(_2683_),
    .A(net679),
    .B(net893));
 sg13g2_o21ai_1 _6054_ (.B1(_2683_),
    .Y(_0425_),
    .A1(net1089),
    .A2(net893));
 sg13g2_nand2_1 _6055_ (.Y(_2684_),
    .A(net690),
    .B(net888));
 sg13g2_o21ai_1 _6056_ (.B1(_2684_),
    .Y(_0426_),
    .A1(net1087),
    .A2(net888));
 sg13g2_nand2_1 _6057_ (.Y(_2685_),
    .A(net1267),
    .B(net888));
 sg13g2_o21ai_1 _6058_ (.B1(_2685_),
    .Y(_0427_),
    .A1(net1085),
    .A2(net888));
 sg13g2_nand2_1 _6059_ (.Y(_2686_),
    .A(net1280),
    .B(net888));
 sg13g2_o21ai_1 _6060_ (.B1(_2686_),
    .Y(_0428_),
    .A1(net1081),
    .A2(net888));
 sg13g2_nand2_1 _6061_ (.Y(_2687_),
    .A(net828),
    .B(net889));
 sg13g2_o21ai_1 _6062_ (.B1(_2687_),
    .Y(_0429_),
    .A1(net1077),
    .A2(net889));
 sg13g2_nand2_1 _6063_ (.Y(_2688_),
    .A(net813),
    .B(net891));
 sg13g2_o21ai_1 _6064_ (.B1(_2688_),
    .Y(_0430_),
    .A1(net1074),
    .A2(net891));
 sg13g2_nand2_1 _6065_ (.Y(_2689_),
    .A(net1254),
    .B(net893));
 sg13g2_o21ai_1 _6066_ (.B1(_2689_),
    .Y(_0431_),
    .A1(net1072),
    .A2(net893));
 sg13g2_or2_1 _6067_ (.X(_2690_),
    .B(_2626_),
    .A(_2519_));
 sg13g2_nand2_1 _6068_ (.Y(_2691_),
    .A(net768),
    .B(net884));
 sg13g2_o21ai_1 _6069_ (.B1(_2691_),
    .Y(_0432_),
    .A1(net1130),
    .A2(net882));
 sg13g2_nand2_1 _6070_ (.Y(_2692_),
    .A(net1249),
    .B(net885));
 sg13g2_o21ai_1 _6071_ (.B1(_2692_),
    .Y(_0433_),
    .A1(net1126),
    .A2(net885));
 sg13g2_nand2_1 _6072_ (.Y(_2693_),
    .A(net743),
    .B(net887));
 sg13g2_o21ai_1 _6073_ (.B1(_2693_),
    .Y(_0434_),
    .A1(net1125),
    .A2(net887));
 sg13g2_nand2_1 _6074_ (.Y(_2694_),
    .A(net1310),
    .B(net885));
 sg13g2_o21ai_1 _6075_ (.B1(_2694_),
    .Y(_0435_),
    .A1(net1122),
    .A2(net885));
 sg13g2_nand2_1 _6076_ (.Y(_2695_),
    .A(net781),
    .B(net886));
 sg13g2_o21ai_1 _6077_ (.B1(_2695_),
    .Y(_0436_),
    .A1(net1117),
    .A2(net886));
 sg13g2_nand2_1 _6078_ (.Y(_2696_),
    .A(net814),
    .B(net883));
 sg13g2_o21ai_1 _6079_ (.B1(_2696_),
    .Y(_0437_),
    .A1(net1114),
    .A2(net883));
 sg13g2_nand2_1 _6080_ (.Y(_2697_),
    .A(net772),
    .B(net885));
 sg13g2_o21ai_1 _6081_ (.B1(_2697_),
    .Y(_0438_),
    .A1(net1112),
    .A2(net885));
 sg13g2_nand2_1 _6082_ (.Y(_2698_),
    .A(net1261),
    .B(net883));
 sg13g2_o21ai_1 _6083_ (.B1(_2698_),
    .Y(_0439_),
    .A1(net1109),
    .A2(net882));
 sg13g2_nand2_1 _6084_ (.Y(_2699_),
    .A(net803),
    .B(net885));
 sg13g2_o21ai_1 _6085_ (.B1(_2699_),
    .Y(_0440_),
    .A1(net1107),
    .A2(net885));
 sg13g2_nand2_1 _6086_ (.Y(_2700_),
    .A(net680),
    .B(net887));
 sg13g2_o21ai_1 _6087_ (.B1(_2700_),
    .Y(_0441_),
    .A1(net1102),
    .A2(net887));
 sg13g2_nand2_1 _6088_ (.Y(_2701_),
    .A(net705),
    .B(net882));
 sg13g2_o21ai_1 _6089_ (.B1(_2701_),
    .Y(_0442_),
    .A1(net1099),
    .A2(net882));
 sg13g2_nand2_1 _6090_ (.Y(_2702_),
    .A(net1364),
    .B(net884));
 sg13g2_o21ai_1 _6091_ (.B1(_2702_),
    .Y(_0443_),
    .A1(net1096),
    .A2(net884));
 sg13g2_nand2_1 _6092_ (.Y(_2703_),
    .A(net812),
    .B(net886));
 sg13g2_o21ai_1 _6093_ (.B1(_2703_),
    .Y(_0444_),
    .A1(net1093),
    .A2(net886));
 sg13g2_nand2_1 _6094_ (.Y(_2704_),
    .A(net779),
    .B(net886));
 sg13g2_o21ai_1 _6095_ (.B1(_2704_),
    .Y(_0445_),
    .A1(net1090),
    .A2(net886));
 sg13g2_nand2_1 _6096_ (.Y(_2705_),
    .A(net1257),
    .B(net882));
 sg13g2_o21ai_1 _6097_ (.B1(_2705_),
    .Y(_0446_),
    .A1(net1086),
    .A2(net882));
 sg13g2_nand2_1 _6098_ (.Y(_2706_),
    .A(net1293),
    .B(net882));
 sg13g2_o21ai_1 _6099_ (.B1(_2706_),
    .Y(_0447_),
    .A1(net1084),
    .A2(net882));
 sg13g2_nand2_1 _6100_ (.Y(_2707_),
    .A(net777),
    .B(net883));
 sg13g2_o21ai_1 _6101_ (.B1(_2707_),
    .Y(_0448_),
    .A1(net1081),
    .A2(net883));
 sg13g2_nand2_1 _6102_ (.Y(_2708_),
    .A(net833),
    .B(net883));
 sg13g2_o21ai_1 _6103_ (.B1(_2708_),
    .Y(_0449_),
    .A1(net1078),
    .A2(net883));
 sg13g2_nand2_1 _6104_ (.Y(_2709_),
    .A(net1264),
    .B(net886));
 sg13g2_o21ai_1 _6105_ (.B1(_2709_),
    .Y(_0450_),
    .A1(net1074),
    .A2(net886));
 sg13g2_nand2_1 _6106_ (.Y(_2710_),
    .A(net811),
    .B(net887));
 sg13g2_o21ai_1 _6107_ (.B1(_2710_),
    .Y(_0451_),
    .A1(net1072),
    .A2(net887));
 sg13g2_nand2_1 _6108_ (.Y(_2711_),
    .A(_0767_),
    .B(_0785_));
 sg13g2_or2_1 _6109_ (.X(_2712_),
    .B(_2711_),
    .A(_2452_));
 sg13g2_nand2_1 _6110_ (.Y(_2713_),
    .A(net817),
    .B(net878));
 sg13g2_o21ai_1 _6111_ (.B1(_2713_),
    .Y(_0452_),
    .A1(net1132),
    .A2(net878));
 sg13g2_nand2_1 _6112_ (.Y(_2714_),
    .A(net684),
    .B(net880));
 sg13g2_o21ai_1 _6113_ (.B1(_2714_),
    .Y(_0453_),
    .A1(net1129),
    .A2(net880));
 sg13g2_nand2_1 _6114_ (.Y(_2715_),
    .A(net765),
    .B(net880));
 sg13g2_o21ai_1 _6115_ (.B1(_2715_),
    .Y(_0454_),
    .A1(net1124),
    .A2(_2712_));
 sg13g2_nand2_1 _6116_ (.Y(_2716_),
    .A(net1336),
    .B(net880));
 sg13g2_o21ai_1 _6117_ (.B1(_2716_),
    .Y(_0455_),
    .A1(net1121),
    .A2(net880));
 sg13g2_nand2_1 _6118_ (.Y(_2717_),
    .A(net728),
    .B(net879));
 sg13g2_o21ai_1 _6119_ (.B1(_2717_),
    .Y(_0456_),
    .A1(net1119),
    .A2(net879));
 sg13g2_nand2_1 _6120_ (.Y(_2718_),
    .A(net775),
    .B(net876));
 sg13g2_o21ai_1 _6121_ (.B1(_2718_),
    .Y(_0457_),
    .A1(net1114),
    .A2(net876));
 sg13g2_nand2_1 _6122_ (.Y(_2719_),
    .A(net659),
    .B(net881));
 sg13g2_o21ai_1 _6123_ (.B1(_2719_),
    .Y(_0458_),
    .A1(net1111),
    .A2(net881));
 sg13g2_nand2_1 _6124_ (.Y(_2720_),
    .A(net1335),
    .B(net877));
 sg13g2_o21ai_1 _6125_ (.B1(_2720_),
    .Y(_0459_),
    .A1(net1108),
    .A2(net877));
 sg13g2_nand2_1 _6126_ (.Y(_2721_),
    .A(net807),
    .B(net879));
 sg13g2_o21ai_1 _6127_ (.B1(_2721_),
    .Y(_0460_),
    .A1(net1105),
    .A2(net879));
 sg13g2_nand2_1 _6128_ (.Y(_2722_),
    .A(net677),
    .B(net881));
 sg13g2_o21ai_1 _6129_ (.B1(_2722_),
    .Y(_0461_),
    .A1(net1103),
    .A2(net881));
 sg13g2_nand2_1 _6130_ (.Y(_2723_),
    .A(net1292),
    .B(net876));
 sg13g2_o21ai_1 _6131_ (.B1(_2723_),
    .Y(_0462_),
    .A1(net1099),
    .A2(net876));
 sg13g2_nand2_1 _6132_ (.Y(_2724_),
    .A(net778),
    .B(net881));
 sg13g2_o21ai_1 _6133_ (.B1(_2724_),
    .Y(_0463_),
    .A1(net1097),
    .A2(net878));
 sg13g2_nand2_1 _6134_ (.Y(_2725_),
    .A(net1271),
    .B(net880));
 sg13g2_o21ai_1 _6135_ (.B1(_2725_),
    .Y(_0464_),
    .A1(net1095),
    .A2(net880));
 sg13g2_nand2_1 _6136_ (.Y(_2726_),
    .A(net1266),
    .B(net879));
 sg13g2_o21ai_1 _6137_ (.B1(_2726_),
    .Y(_0465_),
    .A1(net1089),
    .A2(net879));
 sg13g2_nand2_1 _6138_ (.Y(_2727_),
    .A(net836),
    .B(net878));
 sg13g2_o21ai_1 _6139_ (.B1(_2727_),
    .Y(_0466_),
    .A1(net1087),
    .A2(net878));
 sg13g2_nand2_1 _6140_ (.Y(_2728_),
    .A(net1324),
    .B(net876));
 sg13g2_o21ai_1 _6141_ (.B1(_2728_),
    .Y(_0467_),
    .A1(net1083),
    .A2(net876));
 sg13g2_nand2_1 _6142_ (.Y(_2729_),
    .A(net754),
    .B(net876));
 sg13g2_o21ai_1 _6143_ (.B1(_2729_),
    .Y(_0468_),
    .A1(net1080),
    .A2(net876));
 sg13g2_nand2_1 _6144_ (.Y(_2730_),
    .A(net791),
    .B(net877));
 sg13g2_o21ai_1 _6145_ (.B1(_2730_),
    .Y(_0469_),
    .A1(net1077),
    .A2(net877));
 sg13g2_nand2_1 _6146_ (.Y(_2731_),
    .A(net734),
    .B(net879));
 sg13g2_o21ai_1 _6147_ (.B1(_2731_),
    .Y(_0470_),
    .A1(net1076),
    .A2(net879));
 sg13g2_nand2_1 _6148_ (.Y(_2732_),
    .A(net720),
    .B(net881));
 sg13g2_o21ai_1 _6149_ (.B1(_2732_),
    .Y(_0471_),
    .A1(net1073),
    .A2(net881));
 sg13g2_or2_1 _6150_ (.X(_2733_),
    .B(_2711_),
    .A(_2475_));
 sg13g2_nand2_1 _6151_ (.Y(_2734_),
    .A(net822),
    .B(net874));
 sg13g2_o21ai_1 _6152_ (.B1(_2734_),
    .Y(_0472_),
    .A1(net1131),
    .A2(net874));
 sg13g2_nand2_1 _6153_ (.Y(_2735_),
    .A(net1360),
    .B(net872));
 sg13g2_o21ai_1 _6154_ (.B1(_2735_),
    .Y(_0473_),
    .A1(net1128),
    .A2(net872));
 sg13g2_nand2_1 _6155_ (.Y(_2736_),
    .A(net749),
    .B(net872));
 sg13g2_o21ai_1 _6156_ (.B1(_2736_),
    .Y(_0474_),
    .A1(net1125),
    .A2(net872));
 sg13g2_nand2_1 _6157_ (.Y(_2737_),
    .A(net1350),
    .B(net872));
 sg13g2_o21ai_1 _6158_ (.B1(_2737_),
    .Y(_0475_),
    .A1(net1121),
    .A2(net872));
 sg13g2_nand2_1 _6159_ (.Y(_2738_),
    .A(net1315),
    .B(net873));
 sg13g2_o21ai_1 _6160_ (.B1(_2738_),
    .Y(_0476_),
    .A1(net1117),
    .A2(net875));
 sg13g2_nand2_1 _6161_ (.Y(_2739_),
    .A(net1321),
    .B(net870));
 sg13g2_o21ai_1 _6162_ (.B1(_2739_),
    .Y(_0477_),
    .A1(net1116),
    .A2(net870));
 sg13g2_nand2_1 _6163_ (.Y(_2740_),
    .A(net744),
    .B(net872));
 sg13g2_o21ai_1 _6164_ (.B1(_2740_),
    .Y(_0478_),
    .A1(net1112),
    .A2(net872));
 sg13g2_nand2_1 _6165_ (.Y(_2741_),
    .A(net671),
    .B(net871));
 sg13g2_o21ai_1 _6166_ (.B1(_2741_),
    .Y(_0479_),
    .A1(net1108),
    .A2(net871));
 sg13g2_nand2_1 _6167_ (.Y(_2742_),
    .A(net1294),
    .B(net873));
 sg13g2_o21ai_1 _6168_ (.B1(_2742_),
    .Y(_0480_),
    .A1(net1105),
    .A2(net873));
 sg13g2_nand2_1 _6169_ (.Y(_2743_),
    .A(net658),
    .B(net874));
 sg13g2_o21ai_1 _6170_ (.B1(_2743_),
    .Y(_0481_),
    .A1(net1102),
    .A2(net874));
 sg13g2_nand2_1 _6171_ (.Y(_2744_),
    .A(net737),
    .B(net871));
 sg13g2_o21ai_1 _6172_ (.B1(_2744_),
    .Y(_0482_),
    .A1(_2298_),
    .A2(net871));
 sg13g2_nand2_1 _6173_ (.Y(_2745_),
    .A(net683),
    .B(net871));
 sg13g2_o21ai_1 _6174_ (.B1(_2745_),
    .Y(_0483_),
    .A1(net1097),
    .A2(net875));
 sg13g2_nand2_1 _6175_ (.Y(_2746_),
    .A(net767),
    .B(net873));
 sg13g2_o21ai_1 _6176_ (.B1(_2746_),
    .Y(_0484_),
    .A1(net1093),
    .A2(net873));
 sg13g2_nand2_1 _6177_ (.Y(_2747_),
    .A(net673),
    .B(net874));
 sg13g2_o21ai_1 _6178_ (.B1(_2747_),
    .Y(_0485_),
    .A1(net1089),
    .A2(net874));
 sg13g2_nand2_1 _6179_ (.Y(_2748_),
    .A(net1406),
    .B(net870));
 sg13g2_o21ai_1 _6180_ (.B1(_2748_),
    .Y(_0486_),
    .A1(net1088),
    .A2(net870));
 sg13g2_nand2_1 _6181_ (.Y(_2749_),
    .A(net785),
    .B(net870));
 sg13g2_o21ai_1 _6182_ (.B1(_2749_),
    .Y(_0487_),
    .A1(net1083),
    .A2(net870));
 sg13g2_nand2_1 _6183_ (.Y(_2750_),
    .A(net826),
    .B(net870));
 sg13g2_o21ai_1 _6184_ (.B1(_2750_),
    .Y(_0488_),
    .A1(net1080),
    .A2(net870));
 sg13g2_nand2_1 _6185_ (.Y(_2751_),
    .A(net698),
    .B(net871));
 sg13g2_o21ai_1 _6186_ (.B1(_2751_),
    .Y(_0489_),
    .A1(net1079),
    .A2(net871));
 sg13g2_nand2_1 _6187_ (.Y(_2752_),
    .A(net732),
    .B(net873));
 sg13g2_o21ai_1 _6188_ (.B1(_2752_),
    .Y(_0490_),
    .A1(net1075),
    .A2(net873));
 sg13g2_nand2_1 _6189_ (.Y(_2753_),
    .A(net1331),
    .B(net874));
 sg13g2_o21ai_1 _6190_ (.B1(_2753_),
    .Y(_0491_),
    .A1(net1071),
    .A2(net874));
 sg13g2_or2_1 _6191_ (.X(_2754_),
    .B(_2711_),
    .A(_2497_));
 sg13g2_nand2_1 _6192_ (.Y(_2755_),
    .A(net787),
    .B(net866));
 sg13g2_o21ai_1 _6193_ (.B1(_2755_),
    .Y(_0492_),
    .A1(net1130),
    .A2(net866));
 sg13g2_nand2_1 _6194_ (.Y(_2756_),
    .A(net663),
    .B(net867));
 sg13g2_o21ai_1 _6195_ (.B1(_2756_),
    .Y(_0493_),
    .A1(net1128),
    .A2(net867));
 sg13g2_nand2_1 _6196_ (.Y(_2757_),
    .A(net774),
    .B(net867));
 sg13g2_o21ai_1 _6197_ (.B1(_2757_),
    .Y(_0494_),
    .A1(net1124),
    .A2(net867));
 sg13g2_nand2_1 _6198_ (.Y(_2758_),
    .A(net1303),
    .B(net868));
 sg13g2_o21ai_1 _6199_ (.B1(_2758_),
    .Y(_0495_),
    .A1(net1121),
    .A2(net868));
 sg13g2_nand2_1 _6200_ (.Y(_2759_),
    .A(net712),
    .B(net867));
 sg13g2_o21ai_1 _6201_ (.B1(_2759_),
    .Y(_0496_),
    .A1(net1119),
    .A2(net867));
 sg13g2_nand2_1 _6202_ (.Y(_2760_),
    .A(net716),
    .B(net865));
 sg13g2_o21ai_1 _6203_ (.B1(_2760_),
    .Y(_0497_),
    .A1(_2278_),
    .A2(net864));
 sg13g2_nand2_1 _6204_ (.Y(_2761_),
    .A(net755),
    .B(net869));
 sg13g2_o21ai_1 _6205_ (.B1(_2761_),
    .Y(_0498_),
    .A1(net1111),
    .A2(net869));
 sg13g2_nand2_1 _6206_ (.Y(_2762_),
    .A(net660),
    .B(net864));
 sg13g2_o21ai_1 _6207_ (.B1(_2762_),
    .Y(_0499_),
    .A1(net1108),
    .A2(net865));
 sg13g2_nand2_1 _6208_ (.Y(_2763_),
    .A(net792),
    .B(net867));
 sg13g2_o21ai_1 _6209_ (.B1(_2763_),
    .Y(_0500_),
    .A1(net1107),
    .A2(net867));
 sg13g2_nand2_1 _6210_ (.Y(_2764_),
    .A(net1279),
    .B(net869));
 sg13g2_o21ai_1 _6211_ (.B1(_2764_),
    .Y(_0501_),
    .A1(net1102),
    .A2(net869));
 sg13g2_nand2_1 _6212_ (.Y(_2765_),
    .A(net1278),
    .B(net864));
 sg13g2_o21ai_1 _6213_ (.B1(_2765_),
    .Y(_0502_),
    .A1(net1100),
    .A2(net864));
 sg13g2_nand2_1 _6214_ (.Y(_2766_),
    .A(net800),
    .B(net866));
 sg13g2_o21ai_1 _6215_ (.B1(_2766_),
    .Y(_0503_),
    .A1(net1096),
    .A2(net866));
 sg13g2_nand2_1 _6216_ (.Y(_2767_),
    .A(net796),
    .B(net868));
 sg13g2_o21ai_1 _6217_ (.B1(_2767_),
    .Y(_0504_),
    .A1(net1092),
    .A2(net868));
 sg13g2_nand2_1 _6218_ (.Y(_2768_),
    .A(net700),
    .B(net868));
 sg13g2_o21ai_1 _6219_ (.B1(_2768_),
    .Y(_0505_),
    .A1(net1090),
    .A2(net868));
 sg13g2_nand2_1 _6220_ (.Y(_2769_),
    .A(net1298),
    .B(net864));
 sg13g2_o21ai_1 _6221_ (.B1(_2769_),
    .Y(_0506_),
    .A1(net1086),
    .A2(net864));
 sg13g2_nand2_1 _6222_ (.Y(_2770_),
    .A(net1339),
    .B(net864));
 sg13g2_o21ai_1 _6223_ (.B1(_2770_),
    .Y(_0507_),
    .A1(net1083),
    .A2(net864));
 sg13g2_nand2_1 _6224_ (.Y(_2771_),
    .A(net748),
    .B(net865));
 sg13g2_o21ai_1 _6225_ (.B1(_2771_),
    .Y(_0508_),
    .A1(net1081),
    .A2(net865));
 sg13g2_nand2_1 _6226_ (.Y(_2772_),
    .A(net1250),
    .B(net865));
 sg13g2_o21ai_1 _6227_ (.B1(_2772_),
    .Y(_0509_),
    .A1(net1077),
    .A2(net865));
 sg13g2_nand2_1 _6228_ (.Y(_2773_),
    .A(net664),
    .B(net868));
 sg13g2_o21ai_1 _6229_ (.B1(_2773_),
    .Y(_0510_),
    .A1(net1076),
    .A2(net868));
 sg13g2_nand2_1 _6230_ (.Y(_2774_),
    .A(net675),
    .B(net869));
 sg13g2_o21ai_1 _6231_ (.B1(_2774_),
    .Y(_0511_),
    .A1(net1072),
    .A2(net869));
 sg13g2_or2_1 _6232_ (.X(_2775_),
    .B(_2711_),
    .A(_2519_));
 sg13g2_nand2_1 _6233_ (.Y(_2776_),
    .A(net773),
    .B(net858));
 sg13g2_o21ai_1 _6234_ (.B1(_2776_),
    .Y(_0512_),
    .A1(net1130),
    .A2(net858));
 sg13g2_nand2_1 _6235_ (.Y(_2777_),
    .A(net704),
    .B(net861));
 sg13g2_o21ai_1 _6236_ (.B1(_2777_),
    .Y(_0513_),
    .A1(net1127),
    .A2(net861));
 sg13g2_nand2_1 _6237_ (.Y(_2778_),
    .A(net1322),
    .B(net861));
 sg13g2_o21ai_1 _6238_ (.B1(_2778_),
    .Y(_0514_),
    .A1(net1123),
    .A2(net861));
 sg13g2_nand2_1 _6239_ (.Y(_2779_),
    .A(net681),
    .B(net863));
 sg13g2_o21ai_1 _6240_ (.B1(_2779_),
    .Y(_0515_),
    .A1(net1120),
    .A2(net863));
 sg13g2_nand2_1 _6241_ (.Y(_2780_),
    .A(net1314),
    .B(net862));
 sg13g2_o21ai_1 _6242_ (.B1(_2780_),
    .Y(_0516_),
    .A1(net1118),
    .A2(net862));
 sg13g2_nand2_1 _6243_ (.Y(_2781_),
    .A(net1301),
    .B(net859));
 sg13g2_o21ai_1 _6244_ (.B1(_2781_),
    .Y(_0517_),
    .A1(_2278_),
    .A2(net859));
 sg13g2_nand2_1 _6245_ (.Y(_2782_),
    .A(net1334),
    .B(net861));
 sg13g2_o21ai_1 _6246_ (.B1(_2782_),
    .Y(_0518_),
    .A1(net1112),
    .A2(net861));
 sg13g2_nand2_1 _6247_ (.Y(_2783_),
    .A(net1361),
    .B(net859));
 sg13g2_o21ai_1 _6248_ (.B1(_2783_),
    .Y(_0519_),
    .A1(_2286_),
    .A2(net859));
 sg13g2_nand2_1 _6249_ (.Y(_2784_),
    .A(net1265),
    .B(net861));
 sg13g2_o21ai_1 _6250_ (.B1(_2784_),
    .Y(_0520_),
    .A1(net1107),
    .A2(net861));
 sg13g2_nand2_1 _6251_ (.Y(_2785_),
    .A(net672),
    .B(net863));
 sg13g2_o21ai_1 _6252_ (.B1(_2785_),
    .Y(_0521_),
    .A1(net1104),
    .A2(net863));
 sg13g2_nand2_1 _6253_ (.Y(_2786_),
    .A(net1308),
    .B(net858));
 sg13g2_o21ai_1 _6254_ (.B1(_2786_),
    .Y(_0522_),
    .A1(net1101),
    .A2(net858));
 sg13g2_nand2_1 _6255_ (.Y(_2787_),
    .A(net691),
    .B(net860));
 sg13g2_o21ai_1 _6256_ (.B1(_2787_),
    .Y(_0523_),
    .A1(net1097),
    .A2(net860));
 sg13g2_nand2_1 _6257_ (.Y(_2788_),
    .A(net652),
    .B(net862));
 sg13g2_o21ai_1 _6258_ (.B1(_2788_),
    .Y(_0524_),
    .A1(net1095),
    .A2(net862));
 sg13g2_nand2_1 _6259_ (.Y(_2789_),
    .A(net1332),
    .B(net863));
 sg13g2_o21ai_1 _6260_ (.B1(_2789_),
    .Y(_0525_),
    .A1(net1090),
    .A2(net863));
 sg13g2_nand2_1 _6261_ (.Y(_2790_),
    .A(net731),
    .B(net858));
 sg13g2_o21ai_1 _6262_ (.B1(_2790_),
    .Y(_0526_),
    .A1(net1088),
    .A2(net858));
 sg13g2_nand2_1 _6263_ (.Y(_2791_),
    .A(net780),
    .B(net858));
 sg13g2_o21ai_1 _6264_ (.B1(_2791_),
    .Y(_0527_),
    .A1(net1084),
    .A2(net858));
 sg13g2_nand2_1 _6265_ (.Y(_2792_),
    .A(net1371),
    .B(net859));
 sg13g2_o21ai_1 _6266_ (.B1(_2792_),
    .Y(_0528_),
    .A1(net1080),
    .A2(net859));
 sg13g2_nand2_1 _6267_ (.Y(_2793_),
    .A(net725),
    .B(net859));
 sg13g2_o21ai_1 _6268_ (.B1(_2793_),
    .Y(_0529_),
    .A1(net1079),
    .A2(net859));
 sg13g2_nand2_1 _6269_ (.Y(_2794_),
    .A(net1326),
    .B(net862));
 sg13g2_o21ai_1 _6270_ (.B1(_2794_),
    .Y(_0530_),
    .A1(net1075),
    .A2(net862));
 sg13g2_nand2_1 _6271_ (.Y(_2795_),
    .A(net1337),
    .B(net863));
 sg13g2_o21ai_1 _6272_ (.B1(_2795_),
    .Y(_0531_),
    .A1(net1072),
    .A2(net863));
 sg13g2_nor3_2 _6273_ (.A(_0799_),
    .B(_0813_),
    .C(_2253_),
    .Y(_2796_));
 sg13g2_nor2_1 _6274_ (.A(net1444),
    .B(_2796_),
    .Y(_2797_));
 sg13g2_a21oi_1 _6275_ (.A1(net1132),
    .A2(net854),
    .Y(_0532_),
    .B1(_2797_));
 sg13g2_nor2_1 _6276_ (.A(net1462),
    .B(net855),
    .Y(_2798_));
 sg13g2_a21oi_1 _6277_ (.A1(net1126),
    .A2(net855),
    .Y(_0533_),
    .B1(_2798_));
 sg13g2_nor2_1 _6278_ (.A(net1581),
    .B(net856),
    .Y(_2799_));
 sg13g2_a21oi_1 _6279_ (.A1(net1123),
    .A2(net856),
    .Y(_0534_),
    .B1(_2799_));
 sg13g2_nor2_1 _6280_ (.A(net1536),
    .B(net857),
    .Y(_2800_));
 sg13g2_a21oi_1 _6281_ (.A1(net1122),
    .A2(net857),
    .Y(_0535_),
    .B1(_2800_));
 sg13g2_nor2_1 _6282_ (.A(net1472),
    .B(net856),
    .Y(_2801_));
 sg13g2_a21oi_1 _6283_ (.A1(net1117),
    .A2(net856),
    .Y(_0536_),
    .B1(_2801_));
 sg13g2_nor2_1 _6284_ (.A(net1488),
    .B(net853),
    .Y(_2802_));
 sg13g2_a21oi_1 _6285_ (.A1(net1115),
    .A2(net853),
    .Y(_0537_),
    .B1(_2802_));
 sg13g2_nor2_1 _6286_ (.A(net1464),
    .B(net857),
    .Y(_2803_));
 sg13g2_a21oi_1 _6287_ (.A1(net1112),
    .A2(net857),
    .Y(_0538_),
    .B1(_2803_));
 sg13g2_nor2_1 _6288_ (.A(net1509),
    .B(net852),
    .Y(_2804_));
 sg13g2_a21oi_1 _6289_ (.A1(net1109),
    .A2(net852),
    .Y(_0539_),
    .B1(_2804_));
 sg13g2_nor2_1 _6290_ (.A(net1543),
    .B(net856),
    .Y(_2805_));
 sg13g2_a21oi_1 _6291_ (.A1(_2290_),
    .A2(net856),
    .Y(_0540_),
    .B1(_2805_));
 sg13g2_nor2_1 _6292_ (.A(net1480),
    .B(net857),
    .Y(_2806_));
 sg13g2_a21oi_1 _6293_ (.A1(_2294_),
    .A2(net854),
    .Y(_0541_),
    .B1(_2806_));
 sg13g2_nor2_1 _6294_ (.A(net1563),
    .B(net852),
    .Y(_2807_));
 sg13g2_a21oi_1 _6295_ (.A1(net1101),
    .A2(net852),
    .Y(_0542_),
    .B1(_2807_));
 sg13g2_nor2_1 _6296_ (.A(net1414),
    .B(net854),
    .Y(_2808_));
 sg13g2_a21oi_1 _6297_ (.A1(net1097),
    .A2(net854),
    .Y(_0543_),
    .B1(_2808_));
 sg13g2_nor2_1 _6298_ (.A(net1498),
    .B(net855),
    .Y(_2809_));
 sg13g2_a21oi_1 _6299_ (.A1(net1092),
    .A2(net855),
    .Y(_0544_),
    .B1(_2809_));
 sg13g2_nor2_1 _6300_ (.A(net1537),
    .B(net855),
    .Y(_2810_));
 sg13g2_a21oi_1 _6301_ (.A1(net1091),
    .A2(net855),
    .Y(_0545_),
    .B1(_2810_));
 sg13g2_nor2_1 _6302_ (.A(net1439),
    .B(net852),
    .Y(_2811_));
 sg13g2_a21oi_1 _6303_ (.A1(net1088),
    .A2(net852),
    .Y(_0546_),
    .B1(_2811_));
 sg13g2_nor2_1 _6304_ (.A(net1447),
    .B(net852),
    .Y(_2812_));
 sg13g2_a21oi_1 _6305_ (.A1(net1084),
    .A2(net852),
    .Y(_0547_),
    .B1(_2812_));
 sg13g2_nor2_1 _6306_ (.A(net1419),
    .B(net853),
    .Y(_2813_));
 sg13g2_a21oi_1 _6307_ (.A1(net1082),
    .A2(net853),
    .Y(_0548_),
    .B1(_2813_));
 sg13g2_nor2_1 _6308_ (.A(net1569),
    .B(net853),
    .Y(_2814_));
 sg13g2_a21oi_1 _6309_ (.A1(net1079),
    .A2(net853),
    .Y(_0549_),
    .B1(_2814_));
 sg13g2_nor2_1 _6310_ (.A(net1477),
    .B(net855),
    .Y(_2815_));
 sg13g2_a21oi_1 _6311_ (.A1(net1075),
    .A2(net855),
    .Y(_0550_),
    .B1(_2815_));
 sg13g2_nor2_1 _6312_ (.A(net1435),
    .B(net854),
    .Y(_2816_));
 sg13g2_a21oi_1 _6313_ (.A1(net1073),
    .A2(net854),
    .Y(_0551_),
    .B1(_2816_));
 sg13g2_nor2b_2 _6314_ (.A(_2253_),
    .B_N(_2474_),
    .Y(_2817_));
 sg13g2_nor2_1 _6315_ (.A(net1503),
    .B(net846),
    .Y(_2818_));
 sg13g2_a21oi_1 _6316_ (.A1(net1130),
    .A2(net846),
    .Y(_0552_),
    .B1(_2818_));
 sg13g2_nor2_1 _6317_ (.A(net1560),
    .B(net850),
    .Y(_2819_));
 sg13g2_a21oi_1 _6318_ (.A1(net1127),
    .A2(net850),
    .Y(_0553_),
    .B1(_2819_));
 sg13g2_nor2_1 _6319_ (.A(net1426),
    .B(net850),
    .Y(_2820_));
 sg13g2_a21oi_1 _6320_ (.A1(net1123),
    .A2(net850),
    .Y(_0554_),
    .B1(_2820_));
 sg13g2_nor2_1 _6321_ (.A(net1505),
    .B(net851),
    .Y(_2821_));
 sg13g2_a21oi_1 _6322_ (.A1(net1122),
    .A2(net851),
    .Y(_0555_),
    .B1(_2821_));
 sg13g2_nor2_1 _6323_ (.A(net1590),
    .B(net851),
    .Y(_2822_));
 sg13g2_a21oi_1 _6324_ (.A1(net1118),
    .A2(net851),
    .Y(_0556_),
    .B1(_2822_));
 sg13g2_nor2_1 _6325_ (.A(net1432),
    .B(net847),
    .Y(_2823_));
 sg13g2_a21oi_1 _6326_ (.A1(net1116),
    .A2(net847),
    .Y(_0557_),
    .B1(_2823_));
 sg13g2_nor2_1 _6327_ (.A(net1457),
    .B(net849),
    .Y(_2824_));
 sg13g2_a21oi_1 _6328_ (.A1(net1112),
    .A2(net849),
    .Y(_0558_),
    .B1(_2824_));
 sg13g2_nor2_1 _6329_ (.A(net1549),
    .B(net847),
    .Y(_2825_));
 sg13g2_a21oi_1 _6330_ (.A1(_2286_),
    .A2(net847),
    .Y(_0559_),
    .B1(_2825_));
 sg13g2_nor2_1 _6331_ (.A(net1493),
    .B(net849),
    .Y(_2826_));
 sg13g2_a21oi_1 _6332_ (.A1(net1105),
    .A2(net849),
    .Y(_0560_),
    .B1(_2826_));
 sg13g2_nor2_1 _6333_ (.A(net1460),
    .B(net849),
    .Y(_2827_));
 sg13g2_a21oi_1 _6334_ (.A1(net1103),
    .A2(net849),
    .Y(_0561_),
    .B1(_2827_));
 sg13g2_nor2_1 _6335_ (.A(net1495),
    .B(net846),
    .Y(_2828_));
 sg13g2_a21oi_1 _6336_ (.A1(net1101),
    .A2(net846),
    .Y(_0562_),
    .B1(_2828_));
 sg13g2_nor2_1 _6337_ (.A(net1415),
    .B(net848),
    .Y(_2829_));
 sg13g2_a21oi_1 _6338_ (.A1(net1098),
    .A2(net848),
    .Y(_0563_),
    .B1(_2829_));
 sg13g2_nor2_1 _6339_ (.A(net1577),
    .B(net850),
    .Y(_2830_));
 sg13g2_a21oi_1 _6340_ (.A1(net1095),
    .A2(net850),
    .Y(_0564_),
    .B1(_2830_));
 sg13g2_nor2_1 _6341_ (.A(net1522),
    .B(net849),
    .Y(_2831_));
 sg13g2_a21oi_1 _6342_ (.A1(net1090),
    .A2(net849),
    .Y(_0565_),
    .B1(_2831_));
 sg13g2_nor2_1 _6343_ (.A(net1453),
    .B(net846),
    .Y(_2832_));
 sg13g2_a21oi_1 _6344_ (.A1(net1087),
    .A2(net846),
    .Y(_0566_),
    .B1(_2832_));
 sg13g2_nor2_1 _6345_ (.A(net1408),
    .B(net846),
    .Y(_2833_));
 sg13g2_a21oi_1 _6346_ (.A1(net1085),
    .A2(net846),
    .Y(_0567_),
    .B1(_2833_));
 sg13g2_nor2_1 _6347_ (.A(net1531),
    .B(net847),
    .Y(_2834_));
 sg13g2_a21oi_1 _6348_ (.A1(net1081),
    .A2(net847),
    .Y(_0568_),
    .B1(_2834_));
 sg13g2_nor2_1 _6349_ (.A(net1514),
    .B(net847),
    .Y(_2835_));
 sg13g2_a21oi_1 _6350_ (.A1(net1078),
    .A2(net847),
    .Y(_0569_),
    .B1(_2835_));
 sg13g2_nor2_1 _6351_ (.A(net1423),
    .B(net850),
    .Y(_2836_));
 sg13g2_a21oi_1 _6352_ (.A1(net1074),
    .A2(net850),
    .Y(_0570_),
    .B1(_2836_));
 sg13g2_nor2_1 _6353_ (.A(net1431),
    .B(net848),
    .Y(_2837_));
 sg13g2_a21oi_1 _6354_ (.A1(net1071),
    .A2(net848),
    .Y(_0571_),
    .B1(_2837_));
 sg13g2_nor4_1 _6355_ (.A(_0799_),
    .B(_0811_),
    .C(_0812_),
    .D(_2253_),
    .Y(_2838_));
 sg13g2_nor2_1 _6356_ (.A(net1410),
    .B(net844),
    .Y(_2839_));
 sg13g2_a21oi_1 _6357_ (.A1(net1131),
    .A2(net844),
    .Y(_0572_),
    .B1(_2839_));
 sg13g2_nor2_1 _6358_ (.A(net1525),
    .B(net842),
    .Y(_2840_));
 sg13g2_a21oi_1 _6359_ (.A1(net1128),
    .A2(net842),
    .Y(_0573_),
    .B1(_2840_));
 sg13g2_nor2_1 _6360_ (.A(net1463),
    .B(net842),
    .Y(_2841_));
 sg13g2_a21oi_1 _6361_ (.A1(net1124),
    .A2(net842),
    .Y(_0574_),
    .B1(_2841_));
 sg13g2_nor2_1 _6362_ (.A(net1526),
    .B(net842),
    .Y(_2842_));
 sg13g2_a21oi_1 _6363_ (.A1(net1120),
    .A2(net842),
    .Y(_0575_),
    .B1(_2842_));
 sg13g2_nor2_1 _6364_ (.A(net1588),
    .B(net844),
    .Y(_2843_));
 sg13g2_a21oi_1 _6365_ (.A1(net1119),
    .A2(net845),
    .Y(_0576_),
    .B1(_2843_));
 sg13g2_nor2_1 _6366_ (.A(net1516),
    .B(net839),
    .Y(_2844_));
 sg13g2_a21oi_1 _6367_ (.A1(net1114),
    .A2(net839),
    .Y(_0577_),
    .B1(_2844_));
 sg13g2_nor2_1 _6368_ (.A(net1573),
    .B(net842),
    .Y(_2845_));
 sg13g2_a21oi_1 _6369_ (.A1(net1112),
    .A2(net842),
    .Y(_0578_),
    .B1(_2845_));
 sg13g2_nor2_1 _6370_ (.A(net1499),
    .B(net840),
    .Y(_2846_));
 sg13g2_a21oi_1 _6371_ (.A1(net1109),
    .A2(net840),
    .Y(_0579_),
    .B1(_2846_));
 sg13g2_nor2_1 _6372_ (.A(net1517),
    .B(net843),
    .Y(_2847_));
 sg13g2_a21oi_1 _6373_ (.A1(net1106),
    .A2(net843),
    .Y(_0580_),
    .B1(_2847_));
 sg13g2_nor2_1 _6374_ (.A(net1448),
    .B(net844),
    .Y(_2848_));
 sg13g2_a21oi_1 _6375_ (.A1(_2294_),
    .A2(net844),
    .Y(_0581_),
    .B1(_2848_));
 sg13g2_nor2_1 _6376_ (.A(net1540),
    .B(net839),
    .Y(_2849_));
 sg13g2_a21oi_1 _6377_ (.A1(net1100),
    .A2(net839),
    .Y(_0582_),
    .B1(_2849_));
 sg13g2_nor2_1 _6378_ (.A(net1508),
    .B(net841),
    .Y(_2850_));
 sg13g2_a21oi_1 _6379_ (.A1(net1097),
    .A2(net841),
    .Y(_0583_),
    .B1(_2850_));
 sg13g2_nor2_1 _6380_ (.A(net1486),
    .B(net843),
    .Y(_2851_));
 sg13g2_a21oi_1 _6381_ (.A1(net1094),
    .A2(net843),
    .Y(_0584_),
    .B1(_2851_));
 sg13g2_nor2_1 _6382_ (.A(net1557),
    .B(net843),
    .Y(_2852_));
 sg13g2_a21oi_1 _6383_ (.A1(net1090),
    .A2(net843),
    .Y(_0585_),
    .B1(_2852_));
 sg13g2_nor2_1 _6384_ (.A(net1459),
    .B(net839),
    .Y(_2853_));
 sg13g2_a21oi_1 _6385_ (.A1(net1086),
    .A2(net839),
    .Y(_0586_),
    .B1(_2853_));
 sg13g2_nor2_1 _6386_ (.A(net1469),
    .B(net839),
    .Y(_2854_));
 sg13g2_a21oi_1 _6387_ (.A1(net1084),
    .A2(net839),
    .Y(_0587_),
    .B1(_2854_));
 sg13g2_nor2_1 _6388_ (.A(net1496),
    .B(net840),
    .Y(_2855_));
 sg13g2_a21oi_1 _6389_ (.A1(net1080),
    .A2(net840),
    .Y(_0588_),
    .B1(_2855_));
 sg13g2_nor2_1 _6390_ (.A(net1402),
    .B(net840),
    .Y(_2856_));
 sg13g2_a21oi_1 _6391_ (.A1(net1077),
    .A2(net840),
    .Y(_0589_),
    .B1(_2856_));
 sg13g2_nor2_1 _6392_ (.A(net1454),
    .B(net843),
    .Y(_2857_));
 sg13g2_a21oi_1 _6393_ (.A1(net1076),
    .A2(net843),
    .Y(_0590_),
    .B1(_2857_));
 sg13g2_nor2_1 _6394_ (.A(net1489),
    .B(net844),
    .Y(_2858_));
 sg13g2_a21oi_1 _6395_ (.A1(net1072),
    .A2(net844),
    .Y(_0591_),
    .B1(_2858_));
 sg13g2_nor3_1 _6396_ (.A(net1176),
    .B(net1220),
    .C(net1612),
    .Y(_0592_));
 sg13g2_nor4_1 _6397_ (.A(\vga_tetris.vgaController.verticalCounterQ[5] ),
    .B(\vga_tetris.vgaController.verticalCounterQ[4] ),
    .C(\vga_tetris.vgaController.verticalCounterQ[1] ),
    .D(\vga_tetris.vgaController.verticalCounterQ[0] ),
    .Y(_2859_));
 sg13g2_nor4_1 _6398_ (.A(_0629_),
    .B(\vga_tetris.vgaController.verticalCounterQ[8] ),
    .C(\vga_tetris.vgaController.verticalCounterQ[7] ),
    .D(\vga_tetris.vgaController.verticalCounterQ[6] ),
    .Y(_2860_));
 sg13g2_nand4_1 _6399_ (.B(\vga_tetris.vgaController.verticalCounterQ[2] ),
    .C(_2859_),
    .A(\vga_tetris.vgaController.verticalCounterQ[3] ),
    .Y(_2861_),
    .D(_2860_));
 sg13g2_inv_1 _6400_ (.Y(_2862_),
    .A(_2861_));
 sg13g2_nor3_2 _6401_ (.A(_1752_),
    .B(net1067),
    .C(_2862_),
    .Y(_2863_));
 sg13g2_o21ai_1 _6402_ (.B1(net1234),
    .Y(_2864_),
    .A1(net1478),
    .A2(_2863_));
 sg13g2_a21oi_1 _6403_ (.A1(net1478),
    .A2(_1760_),
    .Y(_0593_),
    .B1(_2864_));
 sg13g2_a21oi_1 _6404_ (.A1(net1478),
    .A2(_1760_),
    .Y(_2865_),
    .B1(net1582));
 sg13g2_nand2_1 _6405_ (.Y(_2866_),
    .A(net1582),
    .B(net1478));
 sg13g2_nand2_1 _6406_ (.Y(_2867_),
    .A(net1234),
    .B(_2866_));
 sg13g2_a21oi_1 _6407_ (.A1(net1063),
    .A2(_2867_),
    .Y(_0594_),
    .B1(_2865_));
 sg13g2_nand2_1 _6408_ (.Y(_2868_),
    .A(net1606),
    .B(_1761_));
 sg13g2_nand3_1 _6409_ (.B(net1582),
    .C(net1478),
    .A(\vga_tetris.vgaController.verticalCounterQ[2] ),
    .Y(_2869_));
 sg13g2_xor2_1 _6410_ (.B(_2866_),
    .A(net1606),
    .X(_2870_));
 sg13g2_nand2_2 _6411_ (.Y(_2871_),
    .A(net1234),
    .B(_2863_));
 sg13g2_o21ai_1 _6412_ (.B1(_2868_),
    .Y(_0595_),
    .A1(_2870_),
    .A2(_2871_));
 sg13g2_nand2_1 _6413_ (.Y(_2872_),
    .A(net1593),
    .B(_1761_));
 sg13g2_nor2_1 _6414_ (.A(_0631_),
    .B(_2869_),
    .Y(_2873_));
 sg13g2_xnor2_1 _6415_ (.Y(_2874_),
    .A(_0631_),
    .B(_2869_));
 sg13g2_o21ai_1 _6416_ (.B1(_2872_),
    .Y(_0596_),
    .A1(_2871_),
    .A2(_2874_));
 sg13g2_a21oi_1 _6417_ (.A1(_1760_),
    .A2(_2873_),
    .Y(_2875_),
    .B1(net1591));
 sg13g2_and3_1 _6418_ (.X(_2876_),
    .A(net1591),
    .B(_1760_),
    .C(_2873_));
 sg13g2_nor3_1 _6419_ (.A(net1219),
    .B(net1592),
    .C(_2876_),
    .Y(_0597_));
 sg13g2_and2_1 _6420_ (.A(net1775),
    .B(_2876_),
    .X(_2877_));
 sg13g2_o21ai_1 _6421_ (.B1(net1235),
    .Y(_2878_),
    .A1(net1775),
    .A2(_2876_));
 sg13g2_nor2_1 _6422_ (.A(_2877_),
    .B(_2878_),
    .Y(_0598_));
 sg13g2_xnor2_1 _6423_ (.Y(_2879_),
    .A(net1728),
    .B(_2877_));
 sg13g2_nor2_1 _6424_ (.A(net1223),
    .B(net1729),
    .Y(_0599_));
 sg13g2_a21o_1 _6425_ (.A2(_2877_),
    .A1(net1728),
    .B1(net1809),
    .X(_2880_));
 sg13g2_nand3_1 _6426_ (.B(net1728),
    .C(_2877_),
    .A(net1809),
    .Y(_2881_));
 sg13g2_and3_1 _6427_ (.X(_0600_),
    .A(net1235),
    .B(_2880_),
    .C(_2881_));
 sg13g2_nand3_1 _6428_ (.B(_1099_),
    .C(_2873_),
    .A(net1591),
    .Y(_2882_));
 sg13g2_nand2_1 _6429_ (.Y(_2883_),
    .A(net1235),
    .B(_2882_));
 sg13g2_a22oi_1 _6430_ (.Y(_0601_),
    .B1(_2883_),
    .B2(net1063),
    .A2(_2881_),
    .A1(_0630_));
 sg13g2_o21ai_1 _6431_ (.B1(_0629_),
    .Y(_2884_),
    .A1(_2871_),
    .A2(_2882_));
 sg13g2_nor2_1 _6432_ (.A(_0629_),
    .B(_2882_),
    .Y(_2885_));
 sg13g2_o21ai_1 _6433_ (.B1(net1063),
    .Y(_2886_),
    .A1(_2871_),
    .A2(_2885_));
 sg13g2_and2_1 _6434_ (.A(net1827),
    .B(_2886_),
    .X(_0602_));
 sg13g2_xnor2_1 _6435_ (.Y(_2887_),
    .A(net1723),
    .B(net1067));
 sg13g2_nor2_1 _6436_ (.A(net1063),
    .B(_2887_),
    .Y(_0603_));
 sg13g2_nor2b_2 _6437_ (.A(net1067),
    .B_N(_1752_),
    .Y(_2888_));
 sg13g2_nand2_1 _6438_ (.Y(_2889_),
    .A(net1599),
    .B(_2888_));
 sg13g2_nand3_1 _6439_ (.B(_1207_),
    .C(net1067),
    .A(_0872_),
    .Y(_2890_));
 sg13g2_a21oi_1 _6440_ (.A1(_2889_),
    .A2(_2890_),
    .Y(_0604_),
    .B1(net1219));
 sg13g2_xnor2_1 _6441_ (.Y(_2891_),
    .A(net1198),
    .B(_0872_));
 sg13g2_a22oi_1 _6442_ (.Y(_2892_),
    .B1(_2891_),
    .B2(net1067),
    .A2(_2888_),
    .A1(net1198));
 sg13g2_nor2_1 _6443_ (.A(net1219),
    .B(_2892_),
    .Y(_0605_));
 sg13g2_a22oi_1 _6444_ (.Y(_2893_),
    .B1(_2888_),
    .B2(net1782),
    .A2(net1067),
    .A1(_0876_));
 sg13g2_o21ai_1 _6445_ (.B1(net1234),
    .Y(_2894_),
    .A1(net1782),
    .A2(_0874_));
 sg13g2_nor2_1 _6446_ (.A(_2893_),
    .B(_2894_),
    .Y(_0606_));
 sg13g2_a22oi_1 _6447_ (.Y(_2895_),
    .B1(_2888_),
    .B2(net1196),
    .A2(_1759_),
    .A1(_1753_));
 sg13g2_o21ai_1 _6448_ (.B1(net1237),
    .Y(_2896_),
    .A1(net1195),
    .A2(_0875_));
 sg13g2_nor2_1 _6449_ (.A(net1882),
    .B(_2896_),
    .Y(_0607_));
 sg13g2_a22oi_1 _6450_ (.Y(_2897_),
    .B1(_2888_),
    .B2(net1194),
    .A2(_1759_),
    .A1(_1755_));
 sg13g2_a21oi_1 _6451_ (.A1(net1196),
    .A2(_0875_),
    .Y(_2898_),
    .B1(net1194));
 sg13g2_nor3_1 _6452_ (.A(net1220),
    .B(_2897_),
    .C(net1859),
    .Y(_0608_));
 sg13g2_a22oi_1 _6453_ (.Y(_2899_),
    .B1(_2888_),
    .B2(net1191),
    .A2(_1759_),
    .A1(_1756_));
 sg13g2_o21ai_1 _6454_ (.B1(net1237),
    .Y(_2900_),
    .A1(net1191),
    .A2(_1754_));
 sg13g2_nor2_1 _6455_ (.A(net1891),
    .B(_2900_),
    .Y(_0609_));
 sg13g2_nand3_1 _6456_ (.B(net1192),
    .C(_1754_),
    .A(net1190),
    .Y(_2901_));
 sg13g2_and2_1 _6457_ (.A(_1757_),
    .B(_2901_),
    .X(_2902_));
 sg13g2_a22oi_1 _6458_ (.Y(_2903_),
    .B1(_2902_),
    .B2(_0626_),
    .A2(_2888_),
    .A1(net1724));
 sg13g2_nor2_1 _6459_ (.A(net1218),
    .B(net1725),
    .Y(_0610_));
 sg13g2_nor2_2 _6460_ (.A(net1887),
    .B(_2901_),
    .Y(_2904_));
 sg13g2_nor2b_1 _6461_ (.A(_1760_),
    .B_N(net1579),
    .Y(_2905_));
 sg13g2_o21ai_1 _6462_ (.B1(net1234),
    .Y(_2906_),
    .A1(_2904_),
    .A2(_2905_));
 sg13g2_a21oi_1 _6463_ (.A1(net1579),
    .A2(_2904_),
    .Y(_0611_),
    .B1(_2906_));
 sg13g2_nor2_1 _6464_ (.A(_1758_),
    .B(_2904_),
    .Y(_2907_));
 sg13g2_nor2_1 _6465_ (.A(_1199_),
    .B(_2907_),
    .Y(_2908_));
 sg13g2_nor2_1 _6466_ (.A(_2888_),
    .B(_2908_),
    .Y(_2909_));
 sg13g2_nor2_1 _6467_ (.A(net1219),
    .B(_2909_),
    .Y(_0612_));
 sg13g2_nand2b_1 _6468_ (.Y(_2910_),
    .B(_1214_),
    .A_N(net1181));
 sg13g2_a21oi_1 _6469_ (.A1(_1203_),
    .A2(_2910_),
    .Y(_2911_),
    .B1(\vga_tetris._vgaController_io_pixelPosY[9] ));
 sg13g2_and2_1 _6470_ (.A(_2863_),
    .B(_2911_),
    .X(_2912_));
 sg13g2_o21ai_1 _6471_ (.B1(_1760_),
    .Y(_2913_),
    .A1(_2862_),
    .A2(_2911_));
 sg13g2_inv_1 _6472_ (.Y(_2914_),
    .A(_2913_));
 sg13g2_o21ai_1 _6473_ (.B1(net1234),
    .Y(_2915_),
    .A1(net1610),
    .A2(net1061));
 sg13g2_a21oi_1 _6474_ (.A1(net1610),
    .A2(_2914_),
    .Y(_0613_),
    .B1(_2915_));
 sg13g2_xor2_1 _6475_ (.B(net1610),
    .A(net1779),
    .X(_2916_));
 sg13g2_a22oi_1 _6476_ (.Y(_2917_),
    .B1(_2916_),
    .B2(net1061),
    .A2(_2913_),
    .A1(net1779));
 sg13g2_nor2_1 _6477_ (.A(net1219),
    .B(_2917_),
    .Y(_0614_));
 sg13g2_a21o_1 _6478_ (.A2(\vga_tetris._vgaController_io_pixelPosY[0] ),
    .A1(\vga_tetris._vgaController_io_pixelPosY[1] ),
    .B1(net1188),
    .X(_2918_));
 sg13g2_and2_1 _6479_ (.A(_0877_),
    .B(_2918_),
    .X(_2919_));
 sg13g2_a22oi_1 _6480_ (.Y(_2920_),
    .B1(_2919_),
    .B2(net1061),
    .A2(_2913_),
    .A1(net1188));
 sg13g2_nor2_1 _6481_ (.A(net1219),
    .B(net1862),
    .Y(_0615_));
 sg13g2_xnor2_1 _6482_ (.Y(_2921_),
    .A(net1187),
    .B(_0877_));
 sg13g2_a22oi_1 _6483_ (.Y(_2922_),
    .B1(_2921_),
    .B2(net1061),
    .A2(_2913_),
    .A1(net1187));
 sg13g2_nor2_1 _6484_ (.A(net1219),
    .B(_2922_),
    .Y(_0616_));
 sg13g2_xnor2_1 _6485_ (.Y(_2923_),
    .A(net1182),
    .B(_0878_));
 sg13g2_a22oi_1 _6486_ (.Y(_2924_),
    .B1(_2923_),
    .B2(net1061),
    .A2(_2913_),
    .A1(net1182));
 sg13g2_nor2_1 _6487_ (.A(net1218),
    .B(net1893),
    .Y(_0617_));
 sg13g2_nor2_1 _6488_ (.A(_0878_),
    .B(_1230_),
    .Y(_2925_));
 sg13g2_inv_1 _6489_ (.Y(_2926_),
    .A(_2925_));
 sg13g2_a21oi_1 _6490_ (.A1(_2912_),
    .A2(_2926_),
    .Y(_2927_),
    .B1(_2913_));
 sg13g2_nand2b_1 _6491_ (.Y(_2928_),
    .B(net1233),
    .A_N(_2927_));
 sg13g2_o21ai_1 _6492_ (.B1(_2910_),
    .Y(_2929_),
    .A1(net1180),
    .A2(net1061));
 sg13g2_nor2_1 _6493_ (.A(_2928_),
    .B(_2929_),
    .Y(_0618_));
 sg13g2_and2_1 _6494_ (.A(net1061),
    .B(_2925_),
    .X(_2930_));
 sg13g2_o21ai_1 _6495_ (.B1(net1233),
    .Y(_2931_),
    .A1(net1179),
    .A2(_2930_));
 sg13g2_a21oi_1 _6496_ (.A1(net1179),
    .A2(_2927_),
    .Y(_0619_),
    .B1(_2931_));
 sg13g2_nand2_1 _6497_ (.Y(_2932_),
    .A(net1179),
    .B(_2930_));
 sg13g2_nand3_1 _6498_ (.B(_0781_),
    .C(net1061),
    .A(net1233),
    .Y(_2933_));
 sg13g2_and2_1 _6499_ (.A(_2928_),
    .B(_2933_),
    .X(_2934_));
 sg13g2_a21oi_1 _6500_ (.A1(_0625_),
    .A2(_2932_),
    .Y(_0620_),
    .B1(_2934_));
 sg13g2_nand2b_1 _6501_ (.Y(_2935_),
    .B(net1640),
    .A_N(_2934_));
 sg13g2_nand2_1 _6502_ (.Y(_2936_),
    .A(net1233),
    .B(_1210_));
 sg13g2_o21ai_1 _6503_ (.B1(_2935_),
    .Y(_0621_),
    .A1(_2932_),
    .A2(_2936_));
 sg13g2_nor3_1 _6504_ (.A(_0624_),
    .B(net1218),
    .C(_2914_),
    .Y(_0622_));
 sg13g2_a21oi_1 _6505_ (.A1(net1175),
    .A2(net1199),
    .Y(_0623_),
    .B1(_2450_));
 sg13g2_dfrbpq_2 _6506_ (.RESET_B(net328),
    .D(_0000_),
    .Q(\vga_tetris.tetrisLogic.stateQ[0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6507_ (.RESET_B(net548),
    .D(_0001_),
    .Q(\vga_tetris.tetrisLogic.stateQ[1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6508_ (.RESET_B(net546),
    .D(net1682),
    .Q(\vga_tetris.tetrisLogic.stateQ[3] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6509_ (.RESET_B(net544),
    .D(net1869),
    .Q(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[2] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _6510_ (.RESET_B(net543),
    .D(_0004_),
    .Q(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[3] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _6511_ (.RESET_B(net542),
    .D(_0005_),
    .Q(\vga_tetris.vgaController.horizontalCounterQ[0] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6512_ (.RESET_B(net541),
    .D(_0006_),
    .Q(\vga_tetris.vgaController.horizontalCounterQ[1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6513_ (.RESET_B(net540),
    .D(_0007_),
    .Q(\vga_tetris.vgaController.horizontalCounterQ[2] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6514_ (.RESET_B(net539),
    .D(_0008_),
    .Q(\vga_tetris.vgaController.horizontalCounterQ[3] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6515_ (.RESET_B(net538),
    .D(_0009_),
    .Q(\vga_tetris.vgaController.horizontalCounterQ[4] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _6516_ (.RESET_B(net537),
    .D(net1649),
    .Q(\vga_tetris.vgaController.horizontalCounterQ[5] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _6517_ (.RESET_B(net536),
    .D(net1679),
    .Q(\vga_tetris.vgaController.horizontalCounterQ[6] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6518_ (.RESET_B(net535),
    .D(_0012_),
    .Q(\vga_tetris.vgaController.horizontalCounterQ[7] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _6519_ (.RESET_B(net534),
    .D(_0013_),
    .Q(\vga_tetris.vgaController.horizontalCounterQ[8] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6520_ (.RESET_B(net533),
    .D(_0014_),
    .Q(\vga_tetris.vgaController.horizontalCounterQ[9] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _6521_ (.RESET_B(net532),
    .D(net647),
    .Q(\vga_tetris.msTimer.msTimerQ[0] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _6522_ (.RESET_B(net531),
    .D(_0016_),
    .Q(\vga_tetris.msTimer.msTimerQ[1] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6523_ (.RESET_B(net530),
    .D(net1386),
    .Q(\vga_tetris.msTimer.msTimerQ[2] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _6524_ (.RESET_B(net529),
    .D(net1636),
    .Q(\vga_tetris.msTimer.msTimerQ[3] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _6525_ (.RESET_B(net528),
    .D(net1646),
    .Q(\vga_tetris.msTimer.msTimerQ[4] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6526_ (.RESET_B(net527),
    .D(net1659),
    .Q(\vga_tetris.msTimer.msTimerQ[5] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6527_ (.RESET_B(net526),
    .D(_0021_),
    .Q(\vga_tetris.msTimer.msTimerQ[6] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6528_ (.RESET_B(net525),
    .D(net1655),
    .Q(\vga_tetris.msTimer.msTimerQ[7] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6529_ (.RESET_B(net524),
    .D(_0023_),
    .Q(\vga_tetris.msTimer.msTimerQ[8] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6530_ (.RESET_B(net523),
    .D(_0024_),
    .Q(\vga_tetris.msTimer.msTimerQ[9] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6531_ (.RESET_B(net522),
    .D(net1735),
    .Q(\vga_tetris.msTimer.msTimerQ[10] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6532_ (.RESET_B(net521),
    .D(_0026_),
    .Q(\vga_tetris.msTimer.msTimerQ[11] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6533_ (.RESET_B(net520),
    .D(net1732),
    .Q(\vga_tetris.msTimer.msTimerQ[12] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6534_ (.RESET_B(net519),
    .D(net1354),
    .Q(\vga_tetris.msTimer.msTimerQ[13] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6535_ (.RESET_B(net518),
    .D(_0029_),
    .Q(\vga_tetris.msTimer.msTimerQ[14] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6536_ (.RESET_B(net517),
    .D(_0030_),
    .Q(\vga_tetris.tetrisLogic.adderSubtracter.io_a[0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6537_ (.RESET_B(net515),
    .D(_0031_),
    .Q(\vga_tetris.tetrisLogic.adderSubtracter.io_a[1] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6538_ (.RESET_B(net513),
    .D(_0032_),
    .Q(\vga_tetris.tetrisLogic.adderSubtracter.io_a[2] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6539_ (.RESET_B(net511),
    .D(_0033_),
    .Q(\vga_tetris.tetrisLogic.adderSubtracter.io_a[3] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6540_ (.RESET_B(net509),
    .D(_0034_),
    .Q(\vga_tetris.tetrisLogic.adderSubtracter.io_a[4] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6541_ (.RESET_B(net507),
    .D(_0035_),
    .Q(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6542_ (.RESET_B(net505),
    .D(_0036_),
    .Q(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[1] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _6543_ (.RESET_B(net503),
    .D(_0037_),
    .Q(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[2] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6544_ (.RESET_B(net501),
    .D(_0038_),
    .Q(\vga_tetris.tetrisLogic.rotationQ[0] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6545_ (.RESET_B(net499),
    .D(_0039_),
    .Q(\vga_tetris.tetrisLogic.rotationQ[1] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _6546_ (.RESET_B(net497),
    .D(_0040_),
    .Q(\vga_tetris.tetrisLogic.stateQ[2] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6547_ (.RESET_B(net495),
    .D(net1855),
    .Q(\vga_tetris.tetrisLogic.stateQ[4] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6548_ (.RESET_B(net493),
    .D(_0042_),
    .Q(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6549_ (.RESET_B(net492),
    .D(_0043_),
    .Q(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _6550_ (.RESET_B(net491),
    .D(_0044_),
    .Q(\vga_tetris.tetrisLogic.shapeDropTimerQ[0] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6551_ (.RESET_B(net490),
    .D(net1535),
    .Q(\vga_tetris.tetrisLogic.shapeDropTimerQ[1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6552_ (.RESET_B(net489),
    .D(_0046_),
    .Q(\vga_tetris.tetrisLogic.shapeDropTimerQ[2] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6553_ (.RESET_B(net488),
    .D(net1694),
    .Q(\vga_tetris.tetrisLogic.shapeDropTimerQ[3] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6554_ (.RESET_B(net487),
    .D(_0048_),
    .Q(\vga_tetris.tetrisLogic.shapeDropTimerQ[4] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6555_ (.RESET_B(net486),
    .D(_0049_),
    .Q(\vga_tetris.tetrisLogic.shapeDropTimerQ[5] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6556_ (.RESET_B(net485),
    .D(_0050_),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _6557_ (.RESET_B(net483),
    .D(net1584),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[1] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6558_ (.RESET_B(net481),
    .D(_0052_),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[2] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6559_ (.RESET_B(net479),
    .D(net1296),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[3] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6560_ (.RESET_B(net477),
    .D(_0054_),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[4] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6561_ (.RESET_B(net475),
    .D(_0055_),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[5] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6562_ (.RESET_B(net473),
    .D(_0056_),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[6] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6563_ (.RESET_B(net471),
    .D(net1383),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[7] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6564_ (.RESET_B(net469),
    .D(net1306),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[8] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6565_ (.RESET_B(net467),
    .D(_0059_),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[9] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _6566_ (.RESET_B(net465),
    .D(_0060_),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[10] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6567_ (.RESET_B(net463),
    .D(_0061_),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[11] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6568_ (.RESET_B(net461),
    .D(net1627),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[12] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6569_ (.RESET_B(net459),
    .D(_0063_),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[13] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6570_ (.RESET_B(net457),
    .D(net1358),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[14] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6571_ (.RESET_B(net455),
    .D(_0065_),
    .Q(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[15] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _6572_ (.RESET_B(net453),
    .D(_0066_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_done ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6573_ (.RESET_B(net452),
    .D(net1727),
    .Q(\vga_tetris.tetrisLogic.addOrRemoveShape.stateQ[0] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6574_ (.RESET_B(net451),
    .D(net649),
    .Q(\vga_tetris.tetrisLogic.addOrRemoveShape.stateQ[1] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6575_ (.RESET_B(net450),
    .D(_0069_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_rowIndex[0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _6576_ (.RESET_B(net448),
    .D(net1712),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_rowIndex[1] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6577_ (.RESET_B(net446),
    .D(_0071_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[0] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6578_ (.RESET_B(net444),
    .D(_0072_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[1] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6579_ (.RESET_B(net442),
    .D(_0073_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[2] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6580_ (.RESET_B(net440),
    .D(_0074_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[3] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6581_ (.RESET_B(net438),
    .D(_0075_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[4] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6582_ (.RESET_B(net436),
    .D(_0076_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[5] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6583_ (.RESET_B(net434),
    .D(net1390),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[6] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6584_ (.RESET_B(net432),
    .D(net1369),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[7] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6585_ (.RESET_B(net430),
    .D(net1507),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[8] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6586_ (.RESET_B(net428),
    .D(_0080_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[9] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6587_ (.RESET_B(net426),
    .D(_0081_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[10] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6588_ (.RESET_B(net424),
    .D(net1352),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[11] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6589_ (.RESET_B(net422),
    .D(_0083_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[12] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6590_ (.RESET_B(net420),
    .D(net1346),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[13] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6591_ (.RESET_B(net418),
    .D(_0085_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[14] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6592_ (.RESET_B(net416),
    .D(_0086_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[15] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6593_ (.RESET_B(net414),
    .D(_0087_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[16] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6594_ (.RESET_B(net412),
    .D(_0088_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[17] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6595_ (.RESET_B(net410),
    .D(_0089_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[18] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6596_ (.RESET_B(net408),
    .D(_0090_),
    .Q(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[19] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _6597_ (.RESET_B(net406),
    .D(net1721),
    .Q(\vga_tetris.tetrisLogic.gameOverResetHappenedQ ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6598_ (.RESET_B(net405),
    .D(_0092_),
    .Q(\vga_tetris.tetrisLogic.checkMoveAllowed.checkIsRunningQ ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _6599_ (.RESET_B(net404),
    .D(_0093_),
    .Q(\vga_tetris.tetrisLogic.addOrRemoveShape.clearingQ ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _6600_ (.RESET_B(net403),
    .D(net1288),
    .Q(\vga_tetris.tetrisLogic._checkMoveAllowed_io_rowIndex[0] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6601_ (.RESET_B(net401),
    .D(net1381),
    .Q(\vga_tetris.tetrisLogic._checkMoveAllowed_io_rowIndex[1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6602_ (.RESET_B(net399),
    .D(net1865),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.operationIsRunningQ ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _6603_ (.RESET_B(net398),
    .D(net1812),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[0] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6604_ (.RESET_B(net397),
    .D(_0098_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6605_ (.RESET_B(net396),
    .D(_0099_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _6606_ (.RESET_B(net395),
    .D(_0100_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _6607_ (.RESET_B(net394),
    .D(net1840),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[4] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6608_ (.RESET_B(net393),
    .D(net1878),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[0] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6609_ (.RESET_B(net392),
    .D(_0103_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6610_ (.RESET_B(net391),
    .D(net1765),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[2] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6611_ (.RESET_B(net390),
    .D(net1747),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[3] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6612_ (.RESET_B(net389),
    .D(net1808),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[4] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _6613_ (.RESET_B(net388),
    .D(_0107_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[0] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6614_ (.RESET_B(net386),
    .D(net1652),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[1] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6615_ (.RESET_B(net384),
    .D(net1553),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[2] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6616_ (.RESET_B(net382),
    .D(net1605),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[3] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6617_ (.RESET_B(net380),
    .D(_0111_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[4] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6618_ (.RESET_B(net378),
    .D(_0112_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6619_ (.RESET_B(net377),
    .D(_0113_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[1] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _6620_ (.RESET_B(net376),
    .D(_0114_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6621_ (.RESET_B(net375),
    .D(_0115_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[0] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6622_ (.RESET_B(net373),
    .D(net1405),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6623_ (.RESET_B(net371),
    .D(net1672),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[2] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6624_ (.RESET_B(net369),
    .D(net832),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[3] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6625_ (.RESET_B(net367),
    .D(_0119_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[4] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6626_ (.RESET_B(net365),
    .D(net1274),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[5] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6627_ (.RESET_B(net363),
    .D(_0121_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[6] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6628_ (.RESET_B(net361),
    .D(_0122_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[7] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6629_ (.RESET_B(net359),
    .D(_0123_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[8] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6630_ (.RESET_B(net357),
    .D(_0124_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[9] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _6631_ (.RESET_B(net355),
    .D(_0125_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[10] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6632_ (.RESET_B(net353),
    .D(_0126_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[11] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6633_ (.RESET_B(net351),
    .D(_0127_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[12] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6634_ (.RESET_B(net349),
    .D(_0128_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[13] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6635_ (.RESET_B(net347),
    .D(_0129_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[14] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6636_ (.RESET_B(net345),
    .D(_0130_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[15] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6637_ (.RESET_B(net343),
    .D(_0131_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[16] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6638_ (.RESET_B(net341),
    .D(_0132_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[17] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6639_ (.RESET_B(net339),
    .D(net1328),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[18] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6640_ (.RESET_B(net337),
    .D(_0134_),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[19] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _6641_ (.RESET_B(net335),
    .D(net1662),
    .Q(\vga_tetris._tetrisLogic_io_score_3[0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _6642_ (.RESET_B(net334),
    .D(net1688),
    .Q(\vga_tetris._tetrisLogic_io_score_3[1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _6643_ (.RESET_B(net333),
    .D(net1742),
    .Q(\vga_tetris._tetrisLogic_io_score_3[2] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _6644_ (.RESET_B(net332),
    .D(_0138_),
    .Q(\vga_tetris._tetrisLogic_io_score_3[3] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6645_ (.RESET_B(net331),
    .D(net1413),
    .Q(\vga_tetris.tetrisLogic.gameOverLogic.buttonPressesCounterQ[0] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6646_ (.RESET_B(net329),
    .D(_0140_),
    .Q(\vga_tetris.tetrisLogic.gameOverLogic.buttonPressesCounterQ[1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6647_ (.RESET_B(net327),
    .D(_0141_),
    .Q(\vga_tetris.tetrisLogic._checkMoveAllowed_io_checkDone ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6648_ (.RESET_B(net326),
    .D(_0142_),
    .Q(\vga_tetris._tetrisLogic_io_score_2[0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _6649_ (.RESET_B(net325),
    .D(_0143_),
    .Q(\vga_tetris._tetrisLogic_io_score_2[1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _6650_ (.RESET_B(net324),
    .D(net1587),
    .Q(\vga_tetris._tetrisLogic_io_score_2[2] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6651_ (.RESET_B(net323),
    .D(_0145_),
    .Q(\vga_tetris._tetrisLogic_io_score_2[3] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6652_ (.RESET_B(net322),
    .D(net1817),
    .Q(\vga_tetris._tetrisLogic_io_score_1[0] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _6653_ (.RESET_B(net321),
    .D(_0147_),
    .Q(\vga_tetris._tetrisLogic_io_score_1[1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6654_ (.RESET_B(net320),
    .D(net1598),
    .Q(\vga_tetris._tetrisLogic_io_score_1[2] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _6655_ (.RESET_B(net319),
    .D(net1760),
    .Q(\vga_tetris._tetrisLogic_io_score_1[3] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6656_ (.RESET_B(net318),
    .D(net1822),
    .Q(\vga_tetris._tetrisLogic_io_score_0[0] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _6657_ (.RESET_B(net317),
    .D(_0151_),
    .Q(\vga_tetris._tetrisLogic_io_score_0[1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _6658_ (.RESET_B(net316),
    .D(net1755),
    .Q(\vga_tetris._tetrisLogic_io_score_0[2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _6659_ (.RESET_B(net315),
    .D(net1758),
    .Q(\vga_tetris._tetrisLogic_io_score_0[3] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _6660_ (.RESET_B(net314),
    .D(net1850),
    .Q(\vga_tetris._tetrisLogic_io_gameOver ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6661_ (.RESET_B(net313),
    .D(_0155_),
    .Q(\vga_tetris.boardMem.board_19[0] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _6662_ (.RESET_B(net312),
    .D(_0156_),
    .Q(\vga_tetris.boardMem.board_19[1] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6663_ (.RESET_B(net311),
    .D(_0157_),
    .Q(\vga_tetris.boardMem.board_19[2] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6664_ (.RESET_B(net310),
    .D(_0158_),
    .Q(\vga_tetris.boardMem.board_19[3] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6665_ (.RESET_B(net309),
    .D(_0159_),
    .Q(\vga_tetris.boardMem.board_19[4] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _6666_ (.RESET_B(net308),
    .D(_0160_),
    .Q(\vga_tetris.boardMem.board_19[5] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6667_ (.RESET_B(net307),
    .D(_0161_),
    .Q(\vga_tetris.boardMem.board_19[6] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _6668_ (.RESET_B(net306),
    .D(_0162_),
    .Q(\vga_tetris.boardMem.board_19[7] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6669_ (.RESET_B(net305),
    .D(_0163_),
    .Q(\vga_tetris.boardMem.board_19[8] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6670_ (.RESET_B(net304),
    .D(_0164_),
    .Q(\vga_tetris.boardMem.board_19[9] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6671_ (.RESET_B(net303),
    .D(_0165_),
    .Q(\vga_tetris.boardMem.board_19[10] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _6672_ (.RESET_B(net302),
    .D(_0166_),
    .Q(\vga_tetris.boardMem.board_19[11] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _6673_ (.RESET_B(net301),
    .D(_0167_),
    .Q(\vga_tetris.boardMem.board_19[12] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6674_ (.RESET_B(net300),
    .D(_0168_),
    .Q(\vga_tetris.boardMem.board_19[13] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6675_ (.RESET_B(net299),
    .D(_0169_),
    .Q(\vga_tetris.boardMem.board_19[14] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _6676_ (.RESET_B(net298),
    .D(_0170_),
    .Q(\vga_tetris.boardMem.board_19[15] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6677_ (.RESET_B(net297),
    .D(net1502),
    .Q(\vga_tetris.boardMem.board_19[16] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6678_ (.RESET_B(net296),
    .D(net1429),
    .Q(\vga_tetris.boardMem.board_19[17] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6679_ (.RESET_B(net295),
    .D(_0173_),
    .Q(\vga_tetris.boardMem.board_19[18] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6680_ (.RESET_B(net294),
    .D(_0174_),
    .Q(\vga_tetris.boardMem.board_19[19] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _6681_ (.RESET_B(net293),
    .D(_0175_),
    .Q(\vga_tetris.inputs.buttonTimerQ_0[0] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _6682_ (.RESET_B(net292),
    .D(_0176_),
    .Q(\vga_tetris.inputs.buttonTimerQ_0[1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6683_ (.RESET_B(net291),
    .D(_0177_),
    .Q(\vga_tetris.inputs.buttonTimerQ_0[2] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6684_ (.RESET_B(net290),
    .D(_0178_),
    .Q(\vga_tetris.inputs.buttonTimerQ_0[3] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6685_ (.RESET_B(net289),
    .D(net1788),
    .Q(\vga_tetris.inputs.buttonTimerQ_0[4] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6686_ (.RESET_B(net288),
    .D(_0180_),
    .Q(\vga_tetris.inputs.buttonTimerQ_0[5] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6687_ (.RESET_B(net287),
    .D(net1396),
    .Q(\vga_tetris.inputs.buttonTimerQ_0[6] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6688_ (.RESET_B(net286),
    .D(_0182_),
    .Q(\vga_tetris.inputs.buttonTimerQ_0[7] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6689_ (.RESET_B(net285),
    .D(net1639),
    .Q(\vga_tetris.inputs.buttonTimerQ_1[0] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6690_ (.RESET_B(net284),
    .D(net1717),
    .Q(\vga_tetris.inputs.buttonTimerQ_1[1] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6691_ (.RESET_B(net283),
    .D(_0185_),
    .Q(\vga_tetris.inputs.buttonTimerQ_1[2] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6692_ (.RESET_B(net282),
    .D(_0186_),
    .Q(\vga_tetris.inputs.buttonTimerQ_1[3] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6693_ (.RESET_B(net281),
    .D(_0187_),
    .Q(\vga_tetris.inputs.buttonTimerQ_1[4] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6694_ (.RESET_B(net280),
    .D(_0188_),
    .Q(\vga_tetris.inputs.buttonTimerQ_1[5] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6695_ (.RESET_B(net279),
    .D(net1618),
    .Q(\vga_tetris.inputs.buttonTimerQ_1[6] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6696_ (.RESET_B(net278),
    .D(net1633),
    .Q(\vga_tetris.inputs.buttonTimerQ_1[7] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6697_ (.RESET_B(net277),
    .D(net806),
    .Q(\vga_tetris.inputs.buttonTimerQ_2[0] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6698_ (.RESET_B(net276),
    .D(net1567),
    .Q(\vga_tetris.inputs.buttonTimerQ_2[1] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6699_ (.RESET_B(net275),
    .D(_0193_),
    .Q(\vga_tetris.inputs.buttonTimerQ_2[2] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6700_ (.RESET_B(net274),
    .D(_0194_),
    .Q(\vga_tetris.inputs.buttonTimerQ_2[3] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6701_ (.RESET_B(net273),
    .D(_0195_),
    .Q(\vga_tetris.inputs.buttonTimerQ_2[4] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6702_ (.RESET_B(net272),
    .D(net1750),
    .Q(\vga_tetris.inputs.buttonTimerQ_2[5] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6703_ (.RESET_B(net271),
    .D(net1691),
    .Q(\vga_tetris.inputs.buttonTimerQ_2[6] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6704_ (.RESET_B(net270),
    .D(net1677),
    .Q(\vga_tetris.inputs.buttonTimerQ_2[7] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6705_ (.RESET_B(net269),
    .D(_0199_),
    .Q(\vga_tetris.inputs.buttonTimerQ_3[0] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6706_ (.RESET_B(net268),
    .D(_0200_),
    .Q(\vga_tetris.inputs.buttonTimerQ_3[1] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6707_ (.RESET_B(net267),
    .D(_0201_),
    .Q(\vga_tetris.inputs.buttonTimerQ_3[2] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6708_ (.RESET_B(net266),
    .D(_0202_),
    .Q(\vga_tetris.inputs.buttonTimerQ_3[3] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6709_ (.RESET_B(net265),
    .D(_0203_),
    .Q(\vga_tetris.inputs.buttonTimerQ_3[4] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6710_ (.RESET_B(net264),
    .D(_0204_),
    .Q(\vga_tetris.inputs.buttonTimerQ_3[5] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6711_ (.RESET_B(net263),
    .D(_0205_),
    .Q(\vga_tetris.inputs.buttonTimerQ_3[6] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6712_ (.RESET_B(net262),
    .D(_0206_),
    .Q(\vga_tetris.inputs.buttonTimerQ_3[7] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6713_ (.RESET_B(net261),
    .D(_0207_),
    .Q(\vga_tetris._inputs_io_rotateButtonActive ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6714_ (.RESET_B(net260),
    .D(net1835),
    .Q(\vga_tetris._inputs_io_leftButtonActive ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _6715_ (.RESET_B(net259),
    .D(_0209_),
    .Q(\vga_tetris._inputs_io_rightButtonActive ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _6716_ (.RESET_B(net258),
    .D(net1685),
    .Q(\vga_tetris._inputs_io_downButtonActive ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6717_ (.RESET_B(net257),
    .D(net1772),
    .Q(\vga_tetris.startTetrisLogicQ ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6718_ (.RESET_B(net256),
    .D(_0212_),
    .Q(\vga_tetris.boardMem.board_0[0] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _6719_ (.RESET_B(net255),
    .D(_0213_),
    .Q(\vga_tetris.boardMem.board_0[1] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6720_ (.RESET_B(net254),
    .D(net1434),
    .Q(\vga_tetris.boardMem.board_0[2] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6721_ (.RESET_B(net253),
    .D(_0215_),
    .Q(\vga_tetris.boardMem.board_0[3] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6722_ (.RESET_B(net252),
    .D(net1471),
    .Q(\vga_tetris.boardMem.board_0[4] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6723_ (.RESET_B(net251),
    .D(_0217_),
    .Q(\vga_tetris.boardMem.board_0[5] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6724_ (.RESET_B(net250),
    .D(net1468),
    .Q(\vga_tetris.boardMem.board_0[6] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6725_ (.RESET_B(net249),
    .D(_0219_),
    .Q(\vga_tetris.boardMem.board_0[7] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6726_ (.RESET_B(net248),
    .D(_0220_),
    .Q(\vga_tetris.boardMem.board_0[8] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6727_ (.RESET_B(net247),
    .D(_0221_),
    .Q(\vga_tetris.boardMem.board_0[9] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6728_ (.RESET_B(net246),
    .D(_0222_),
    .Q(\vga_tetris.boardMem.board_0[10] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _6729_ (.RESET_B(net245),
    .D(net1491),
    .Q(\vga_tetris.boardMem.board_0[11] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _6730_ (.RESET_B(net244),
    .D(net1475),
    .Q(\vga_tetris.boardMem.board_0[12] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6731_ (.RESET_B(net243),
    .D(_0225_),
    .Q(\vga_tetris.boardMem.board_0[13] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6732_ (.RESET_B(net242),
    .D(_0226_),
    .Q(\vga_tetris.boardMem.board_0[14] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6733_ (.RESET_B(net241),
    .D(net1399),
    .Q(\vga_tetris.boardMem.board_0[15] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6734_ (.RESET_B(net240),
    .D(_0228_),
    .Q(\vga_tetris.boardMem.board_0[16] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6735_ (.RESET_B(net239),
    .D(_0229_),
    .Q(\vga_tetris.boardMem.board_0[17] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6736_ (.RESET_B(net238),
    .D(_0230_),
    .Q(\vga_tetris.boardMem.board_0[18] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6737_ (.RESET_B(net237),
    .D(_0231_),
    .Q(\vga_tetris.boardMem.board_0[19] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _6738_ (.RESET_B(net236),
    .D(_0232_),
    .Q(\vga_tetris.boardMem.board_1[0] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _6739_ (.RESET_B(net235),
    .D(_0233_),
    .Q(\vga_tetris.boardMem.board_1[1] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6740_ (.RESET_B(net234),
    .D(_0234_),
    .Q(\vga_tetris.boardMem.board_1[2] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6741_ (.RESET_B(net233),
    .D(_0235_),
    .Q(\vga_tetris.boardMem.board_1[3] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6742_ (.RESET_B(net232),
    .D(_0236_),
    .Q(\vga_tetris.boardMem.board_1[4] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6743_ (.RESET_B(net231),
    .D(_0237_),
    .Q(\vga_tetris.boardMem.board_1[5] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6744_ (.RESET_B(net230),
    .D(_0238_),
    .Q(\vga_tetris.boardMem.board_1[6] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6745_ (.RESET_B(net229),
    .D(_0239_),
    .Q(\vga_tetris.boardMem.board_1[7] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6746_ (.RESET_B(net228),
    .D(_0240_),
    .Q(\vga_tetris.boardMem.board_1[8] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6747_ (.RESET_B(net227),
    .D(_0241_),
    .Q(\vga_tetris.boardMem.board_1[9] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6748_ (.RESET_B(net226),
    .D(_0242_),
    .Q(\vga_tetris.boardMem.board_1[10] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _6749_ (.RESET_B(net225),
    .D(net1393),
    .Q(\vga_tetris.boardMem.board_1[11] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _6750_ (.RESET_B(net224),
    .D(_0244_),
    .Q(\vga_tetris.boardMem.board_1[12] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6751_ (.RESET_B(net223),
    .D(net1520),
    .Q(\vga_tetris.boardMem.board_1[13] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6752_ (.RESET_B(net222),
    .D(_0246_),
    .Q(\vga_tetris.boardMem.board_1[14] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _6753_ (.RESET_B(net221),
    .D(_0247_),
    .Q(\vga_tetris.boardMem.board_1[15] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6754_ (.RESET_B(net220),
    .D(_0248_),
    .Q(\vga_tetris.boardMem.board_1[16] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6755_ (.RESET_B(net219),
    .D(_0249_),
    .Q(\vga_tetris.boardMem.board_1[17] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6756_ (.RESET_B(net218),
    .D(_0250_),
    .Q(\vga_tetris.boardMem.board_1[18] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6757_ (.RESET_B(net217),
    .D(_0251_),
    .Q(\vga_tetris.boardMem.board_1[19] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _6758_ (.RESET_B(net216),
    .D(_0252_),
    .Q(\vga_tetris.boardMem.board_2[0] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _6759_ (.RESET_B(net215),
    .D(_0253_),
    .Q(\vga_tetris.boardMem.board_2[1] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6760_ (.RESET_B(net214),
    .D(_0254_),
    .Q(\vga_tetris.boardMem.board_2[2] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6761_ (.RESET_B(net213),
    .D(_0255_),
    .Q(\vga_tetris.boardMem.board_2[3] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6762_ (.RESET_B(net212),
    .D(_0256_),
    .Q(\vga_tetris.boardMem.board_2[4] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _6763_ (.RESET_B(net211),
    .D(_0257_),
    .Q(\vga_tetris.boardMem.board_2[5] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6764_ (.RESET_B(net210),
    .D(_0258_),
    .Q(\vga_tetris.boardMem.board_2[6] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6765_ (.RESET_B(net209),
    .D(_0259_),
    .Q(\vga_tetris.boardMem.board_2[7] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6766_ (.RESET_B(net208),
    .D(_0260_),
    .Q(\vga_tetris.boardMem.board_2[8] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6767_ (.RESET_B(net207),
    .D(_0261_),
    .Q(\vga_tetris.boardMem.board_2[9] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6768_ (.RESET_B(net206),
    .D(_0262_),
    .Q(\vga_tetris.boardMem.board_2[10] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _6769_ (.RESET_B(net205),
    .D(_0263_),
    .Q(\vga_tetris.boardMem.board_2[11] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _6770_ (.RESET_B(net204),
    .D(_0264_),
    .Q(\vga_tetris.boardMem.board_2[12] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6771_ (.RESET_B(net203),
    .D(net1529),
    .Q(\vga_tetris.boardMem.board_2[13] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6772_ (.RESET_B(net202),
    .D(_0266_),
    .Q(\vga_tetris.boardMem.board_2[14] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _6773_ (.RESET_B(net201),
    .D(_0267_),
    .Q(\vga_tetris.boardMem.board_2[15] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6774_ (.RESET_B(net200),
    .D(net1438),
    .Q(\vga_tetris.boardMem.board_2[16] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6775_ (.RESET_B(net199),
    .D(_0269_),
    .Q(\vga_tetris.boardMem.board_2[17] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6776_ (.RESET_B(net198),
    .D(_0270_),
    .Q(\vga_tetris.boardMem.board_2[18] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6777_ (.RESET_B(net197),
    .D(_0271_),
    .Q(\vga_tetris.boardMem.board_2[19] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _6778_ (.RESET_B(net196),
    .D(_0272_),
    .Q(\vga_tetris.boardMem.board_3[0] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _6779_ (.RESET_B(net195),
    .D(_0273_),
    .Q(\vga_tetris.boardMem.board_3[1] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _6780_ (.RESET_B(net194),
    .D(_0274_),
    .Q(\vga_tetris.boardMem.board_3[2] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6781_ (.RESET_B(net193),
    .D(_0275_),
    .Q(\vga_tetris.boardMem.board_3[3] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6782_ (.RESET_B(net192),
    .D(_0276_),
    .Q(\vga_tetris.boardMem.board_3[4] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6783_ (.RESET_B(net191),
    .D(_0277_),
    .Q(\vga_tetris.boardMem.board_3[5] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6784_ (.RESET_B(net190),
    .D(_0278_),
    .Q(\vga_tetris.boardMem.board_3[6] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6785_ (.RESET_B(net189),
    .D(_0279_),
    .Q(\vga_tetris.boardMem.board_3[7] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6786_ (.RESET_B(net188),
    .D(_0280_),
    .Q(\vga_tetris.boardMem.board_3[8] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6787_ (.RESET_B(net187),
    .D(_0281_),
    .Q(\vga_tetris.boardMem.board_3[9] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6788_ (.RESET_B(net186),
    .D(_0282_),
    .Q(\vga_tetris.boardMem.board_3[10] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _6789_ (.RESET_B(net185),
    .D(_0283_),
    .Q(\vga_tetris.boardMem.board_3[11] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _6790_ (.RESET_B(net184),
    .D(_0284_),
    .Q(\vga_tetris.boardMem.board_3[12] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6791_ (.RESET_B(net183),
    .D(_0285_),
    .Q(\vga_tetris.boardMem.board_3[13] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6792_ (.RESET_B(net182),
    .D(_0286_),
    .Q(\vga_tetris.boardMem.board_3[14] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6793_ (.RESET_B(net181),
    .D(_0287_),
    .Q(\vga_tetris.boardMem.board_3[15] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6794_ (.RESET_B(net180),
    .D(_0288_),
    .Q(\vga_tetris.boardMem.board_3[16] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6795_ (.RESET_B(net179),
    .D(_0289_),
    .Q(\vga_tetris.boardMem.board_3[17] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6796_ (.RESET_B(net178),
    .D(_0290_),
    .Q(\vga_tetris.boardMem.board_3[18] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6797_ (.RESET_B(net177),
    .D(_0291_),
    .Q(\vga_tetris.boardMem.board_3[19] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6798_ (.RESET_B(net176),
    .D(_0292_),
    .Q(\vga_tetris.boardMem.board_4[0] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _6799_ (.RESET_B(net175),
    .D(_0293_),
    .Q(\vga_tetris.boardMem.board_4[1] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6800_ (.RESET_B(net174),
    .D(_0294_),
    .Q(\vga_tetris.boardMem.board_4[2] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6801_ (.RESET_B(net173),
    .D(_0295_),
    .Q(\vga_tetris.boardMem.board_4[3] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6802_ (.RESET_B(net172),
    .D(_0296_),
    .Q(\vga_tetris.boardMem.board_4[4] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6803_ (.RESET_B(net171),
    .D(_0297_),
    .Q(\vga_tetris.boardMem.board_4[5] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6804_ (.RESET_B(net170),
    .D(_0298_),
    .Q(\vga_tetris.boardMem.board_4[6] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _6805_ (.RESET_B(net169),
    .D(_0299_),
    .Q(\vga_tetris.boardMem.board_4[7] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6806_ (.RESET_B(net168),
    .D(_0300_),
    .Q(\vga_tetris.boardMem.board_4[8] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6807_ (.RESET_B(net167),
    .D(_0301_),
    .Q(\vga_tetris.boardMem.board_4[9] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6808_ (.RESET_B(net166),
    .D(_0302_),
    .Q(\vga_tetris.boardMem.board_4[10] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _6809_ (.RESET_B(net165),
    .D(_0303_),
    .Q(\vga_tetris.boardMem.board_4[11] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _6810_ (.RESET_B(net164),
    .D(_0304_),
    .Q(\vga_tetris.boardMem.board_4[12] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6811_ (.RESET_B(net163),
    .D(_0305_),
    .Q(\vga_tetris.boardMem.board_4[13] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6812_ (.RESET_B(net162),
    .D(_0306_),
    .Q(\vga_tetris.boardMem.board_4[14] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _6813_ (.RESET_B(net161),
    .D(_0307_),
    .Q(\vga_tetris.boardMem.board_4[15] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6814_ (.RESET_B(net160),
    .D(_0308_),
    .Q(\vga_tetris.boardMem.board_4[16] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6815_ (.RESET_B(net159),
    .D(_0309_),
    .Q(\vga_tetris.boardMem.board_4[17] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6816_ (.RESET_B(net158),
    .D(_0310_),
    .Q(\vga_tetris.boardMem.board_4[18] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6817_ (.RESET_B(net157),
    .D(_0311_),
    .Q(\vga_tetris.boardMem.board_4[19] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _6818_ (.RESET_B(net156),
    .D(_0312_),
    .Q(\vga_tetris.boardMem.board_5[0] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _6819_ (.RESET_B(net155),
    .D(_0313_),
    .Q(\vga_tetris.boardMem.board_5[1] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _6820_ (.RESET_B(net154),
    .D(_0314_),
    .Q(\vga_tetris.boardMem.board_5[2] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6821_ (.RESET_B(net153),
    .D(_0315_),
    .Q(\vga_tetris.boardMem.board_5[3] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6822_ (.RESET_B(net152),
    .D(_0316_),
    .Q(\vga_tetris.boardMem.board_5[4] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6823_ (.RESET_B(net151),
    .D(_0317_),
    .Q(\vga_tetris.boardMem.board_5[5] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6824_ (.RESET_B(net150),
    .D(_0318_),
    .Q(\vga_tetris.boardMem.board_5[6] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _6825_ (.RESET_B(net149),
    .D(_0319_),
    .Q(\vga_tetris.boardMem.board_5[7] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6826_ (.RESET_B(net148),
    .D(_0320_),
    .Q(\vga_tetris.boardMem.board_5[8] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6827_ (.RESET_B(net147),
    .D(_0321_),
    .Q(\vga_tetris.boardMem.board_5[9] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6828_ (.RESET_B(net146),
    .D(_0322_),
    .Q(\vga_tetris.boardMem.board_5[10] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _6829_ (.RESET_B(net145),
    .D(_0323_),
    .Q(\vga_tetris.boardMem.board_5[11] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _6830_ (.RESET_B(net144),
    .D(net1300),
    .Q(\vga_tetris.boardMem.board_5[12] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6831_ (.RESET_B(net143),
    .D(_0325_),
    .Q(\vga_tetris.boardMem.board_5[13] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6832_ (.RESET_B(net142),
    .D(_0326_),
    .Q(\vga_tetris.boardMem.board_5[14] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _6833_ (.RESET_B(net141),
    .D(_0327_),
    .Q(\vga_tetris.boardMem.board_5[15] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6834_ (.RESET_B(net140),
    .D(_0328_),
    .Q(\vga_tetris.boardMem.board_5[16] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6835_ (.RESET_B(net139),
    .D(_0329_),
    .Q(\vga_tetris.boardMem.board_5[17] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6836_ (.RESET_B(net138),
    .D(_0330_),
    .Q(\vga_tetris.boardMem.board_5[18] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6837_ (.RESET_B(net137),
    .D(net784),
    .Q(\vga_tetris.boardMem.board_5[19] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6838_ (.RESET_B(net136),
    .D(_0332_),
    .Q(\vga_tetris.boardMem.board_6[0] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _6839_ (.RESET_B(net135),
    .D(_0333_),
    .Q(\vga_tetris.boardMem.board_6[1] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6840_ (.RESET_B(net134),
    .D(_0334_),
    .Q(\vga_tetris.boardMem.board_6[2] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6841_ (.RESET_B(net133),
    .D(_0335_),
    .Q(\vga_tetris.boardMem.board_6[3] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6842_ (.RESET_B(net132),
    .D(_0336_),
    .Q(\vga_tetris.boardMem.board_6[4] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6843_ (.RESET_B(net131),
    .D(_0337_),
    .Q(\vga_tetris.boardMem.board_6[5] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6844_ (.RESET_B(net130),
    .D(_0338_),
    .Q(\vga_tetris.boardMem.board_6[6] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6845_ (.RESET_B(net129),
    .D(_0339_),
    .Q(\vga_tetris.boardMem.board_6[7] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6846_ (.RESET_B(net128),
    .D(_0340_),
    .Q(\vga_tetris.boardMem.board_6[8] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6847_ (.RESET_B(net127),
    .D(_0341_),
    .Q(\vga_tetris.boardMem.board_6[9] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6848_ (.RESET_B(net126),
    .D(_0342_),
    .Q(\vga_tetris.boardMem.board_6[10] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _6849_ (.RESET_B(net125),
    .D(net835),
    .Q(\vga_tetris.boardMem.board_6[11] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _6850_ (.RESET_B(net124),
    .D(_0344_),
    .Q(\vga_tetris.boardMem.board_6[12] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6851_ (.RESET_B(net123),
    .D(net795),
    .Q(\vga_tetris.boardMem.board_6[13] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6852_ (.RESET_B(net122),
    .D(_0346_),
    .Q(\vga_tetris.boardMem.board_6[14] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _6853_ (.RESET_B(net121),
    .D(_0347_),
    .Q(\vga_tetris.boardMem.board_6[15] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6854_ (.RESET_B(net120),
    .D(net656),
    .Q(\vga_tetris.boardMem.board_6[16] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6855_ (.RESET_B(net119),
    .D(_0349_),
    .Q(\vga_tetris.boardMem.board_6[17] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6856_ (.RESET_B(net118),
    .D(_0350_),
    .Q(\vga_tetris.boardMem.board_6[18] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6857_ (.RESET_B(net117),
    .D(_0351_),
    .Q(\vga_tetris.boardMem.board_6[19] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _6858_ (.RESET_B(net116),
    .D(_0352_),
    .Q(\vga_tetris.boardMem.board_7[0] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _6859_ (.RESET_B(net115),
    .D(_0353_),
    .Q(\vga_tetris.boardMem.board_7[1] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6860_ (.RESET_B(net114),
    .D(_0354_),
    .Q(\vga_tetris.boardMem.board_7[2] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6861_ (.RESET_B(net113),
    .D(_0355_),
    .Q(\vga_tetris.boardMem.board_7[3] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6862_ (.RESET_B(net112),
    .D(_0356_),
    .Q(\vga_tetris.boardMem.board_7[4] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6863_ (.RESET_B(net111),
    .D(_0357_),
    .Q(\vga_tetris.boardMem.board_7[5] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6864_ (.RESET_B(net110),
    .D(_0358_),
    .Q(\vga_tetris.boardMem.board_7[6] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6865_ (.RESET_B(net109),
    .D(_0359_),
    .Q(\vga_tetris.boardMem.board_7[7] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6866_ (.RESET_B(net108),
    .D(_0360_),
    .Q(\vga_tetris.boardMem.board_7[8] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6867_ (.RESET_B(net107),
    .D(_0361_),
    .Q(\vga_tetris.boardMem.board_7[9] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6868_ (.RESET_B(net106),
    .D(_0362_),
    .Q(\vga_tetris.boardMem.board_7[10] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _6869_ (.RESET_B(net105),
    .D(net757),
    .Q(\vga_tetris.boardMem.board_7[11] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _6870_ (.RESET_B(net104),
    .D(_0364_),
    .Q(\vga_tetris.boardMem.board_7[12] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6871_ (.RESET_B(net103),
    .D(_0365_),
    .Q(\vga_tetris.boardMem.board_7[13] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6872_ (.RESET_B(net102),
    .D(_0366_),
    .Q(\vga_tetris.boardMem.board_7[14] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _6873_ (.RESET_B(net101),
    .D(_0367_),
    .Q(\vga_tetris.boardMem.board_7[15] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _6874_ (.RESET_B(net100),
    .D(_0368_),
    .Q(\vga_tetris.boardMem.board_7[16] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6875_ (.RESET_B(net99),
    .D(_0369_),
    .Q(\vga_tetris.boardMem.board_7[17] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6876_ (.RESET_B(net98),
    .D(_0370_),
    .Q(\vga_tetris.boardMem.board_7[18] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6877_ (.RESET_B(net97),
    .D(net825),
    .Q(\vga_tetris.boardMem.board_7[19] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _6878_ (.RESET_B(net96),
    .D(net697),
    .Q(\vga_tetris.boardMem.board_8[0] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _6879_ (.RESET_B(net95),
    .D(_0373_),
    .Q(\vga_tetris.boardMem.board_8[1] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6880_ (.RESET_B(net94),
    .D(_0374_),
    .Q(\vga_tetris.boardMem.board_8[2] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6881_ (.RESET_B(net93),
    .D(_0375_),
    .Q(\vga_tetris.boardMem.board_8[3] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6882_ (.RESET_B(net92),
    .D(_0376_),
    .Q(\vga_tetris.boardMem.board_8[4] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6883_ (.RESET_B(net91),
    .D(_0377_),
    .Q(\vga_tetris.boardMem.board_8[5] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6884_ (.RESET_B(net90),
    .D(_0378_),
    .Q(\vga_tetris.boardMem.board_8[6] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6885_ (.RESET_B(net89),
    .D(_0379_),
    .Q(\vga_tetris.boardMem.board_8[7] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6886_ (.RESET_B(net88),
    .D(_0380_),
    .Q(\vga_tetris.boardMem.board_8[8] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6887_ (.RESET_B(net87),
    .D(_0381_),
    .Q(\vga_tetris.boardMem.board_8[9] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6888_ (.RESET_B(net86),
    .D(_0382_),
    .Q(\vga_tetris.boardMem.board_8[10] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _6889_ (.RESET_B(net85),
    .D(_0383_),
    .Q(\vga_tetris.boardMem.board_8[11] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _6890_ (.RESET_B(net84),
    .D(_0384_),
    .Q(\vga_tetris.boardMem.board_8[12] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6891_ (.RESET_B(net83),
    .D(_0385_),
    .Q(\vga_tetris.boardMem.board_8[13] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6892_ (.RESET_B(net82),
    .D(_0386_),
    .Q(\vga_tetris.boardMem.board_8[14] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _6893_ (.RESET_B(net81),
    .D(_0387_),
    .Q(\vga_tetris.boardMem.board_8[15] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6894_ (.RESET_B(net80),
    .D(_0388_),
    .Q(\vga_tetris.boardMem.board_8[16] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6895_ (.RESET_B(net79),
    .D(_0389_),
    .Q(\vga_tetris.boardMem.board_8[17] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6896_ (.RESET_B(net78),
    .D(_0390_),
    .Q(\vga_tetris.boardMem.board_8[18] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6897_ (.RESET_B(net77),
    .D(_0391_),
    .Q(\vga_tetris.boardMem.board_8[19] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6898_ (.RESET_B(net76),
    .D(net799),
    .Q(\vga_tetris.boardMem.board_9[0] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _6899_ (.RESET_B(net75),
    .D(net770),
    .Q(\vga_tetris.boardMem.board_9[1] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6900_ (.RESET_B(net74),
    .D(_0394_),
    .Q(\vga_tetris.boardMem.board_9[2] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6901_ (.RESET_B(net73),
    .D(net711),
    .Q(\vga_tetris.boardMem.board_9[3] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6902_ (.RESET_B(net72),
    .D(_0396_),
    .Q(\vga_tetris.boardMem.board_9[4] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6903_ (.RESET_B(net71),
    .D(_0397_),
    .Q(\vga_tetris.boardMem.board_9[5] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6904_ (.RESET_B(net70),
    .D(_0398_),
    .Q(\vga_tetris.boardMem.board_9[6] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _6905_ (.RESET_B(net69),
    .D(_0399_),
    .Q(\vga_tetris.boardMem.board_9[7] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6906_ (.RESET_B(net68),
    .D(_0400_),
    .Q(\vga_tetris.boardMem.board_9[8] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6907_ (.RESET_B(net67),
    .D(_0401_),
    .Q(\vga_tetris.boardMem.board_9[9] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6908_ (.RESET_B(net66),
    .D(_0402_),
    .Q(\vga_tetris.boardMem.board_9[10] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _6909_ (.RESET_B(net65),
    .D(_0403_),
    .Q(\vga_tetris.boardMem.board_9[11] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _6910_ (.RESET_B(net64),
    .D(_0404_),
    .Q(\vga_tetris.boardMem.board_9[12] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6911_ (.RESET_B(net63),
    .D(_0405_),
    .Q(\vga_tetris.boardMem.board_9[13] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6912_ (.RESET_B(net62),
    .D(_0406_),
    .Q(\vga_tetris.boardMem.board_9[14] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6913_ (.RESET_B(net61),
    .D(_0407_),
    .Q(\vga_tetris.boardMem.board_9[15] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6914_ (.RESET_B(net60),
    .D(_0408_),
    .Q(\vga_tetris.boardMem.board_9[16] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6915_ (.RESET_B(net59),
    .D(_0409_),
    .Q(\vga_tetris.boardMem.board_9[17] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6916_ (.RESET_B(net58),
    .D(_0410_),
    .Q(\vga_tetris.boardMem.board_9[18] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6917_ (.RESET_B(net57),
    .D(_0411_),
    .Q(\vga_tetris.boardMem.board_9[19] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6918_ (.RESET_B(net56),
    .D(_0412_),
    .Q(\vga_tetris.boardMem.board_10[0] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6919_ (.RESET_B(net55),
    .D(_0413_),
    .Q(\vga_tetris.boardMem.board_10[1] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6920_ (.RESET_B(net54),
    .D(_0414_),
    .Q(\vga_tetris.boardMem.board_10[2] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6921_ (.RESET_B(net53),
    .D(_0415_),
    .Q(\vga_tetris.boardMem.board_10[3] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6922_ (.RESET_B(net52),
    .D(_0416_),
    .Q(\vga_tetris.boardMem.board_10[4] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _6923_ (.RESET_B(net51),
    .D(_0417_),
    .Q(\vga_tetris.boardMem.board_10[5] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6924_ (.RESET_B(net50),
    .D(_0418_),
    .Q(\vga_tetris.boardMem.board_10[6] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _6925_ (.RESET_B(net49),
    .D(_0419_),
    .Q(\vga_tetris.boardMem.board_10[7] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6926_ (.RESET_B(net48),
    .D(_0420_),
    .Q(\vga_tetris.boardMem.board_10[8] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6927_ (.RESET_B(net47),
    .D(_0421_),
    .Q(\vga_tetris.boardMem.board_10[9] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6928_ (.RESET_B(net46),
    .D(_0422_),
    .Q(\vga_tetris.boardMem.board_10[10] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _6929_ (.RESET_B(net45),
    .D(net723),
    .Q(\vga_tetris.boardMem.board_10[11] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _6930_ (.RESET_B(net44),
    .D(_0424_),
    .Q(\vga_tetris.boardMem.board_10[12] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6931_ (.RESET_B(net43),
    .D(_0425_),
    .Q(\vga_tetris.boardMem.board_10[13] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6932_ (.RESET_B(net42),
    .D(_0426_),
    .Q(\vga_tetris.boardMem.board_10[14] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _6933_ (.RESET_B(net41),
    .D(_0427_),
    .Q(\vga_tetris.boardMem.board_10[15] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6934_ (.RESET_B(net40),
    .D(_0428_),
    .Q(\vga_tetris.boardMem.board_10[16] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6935_ (.RESET_B(net39),
    .D(_0429_),
    .Q(\vga_tetris.boardMem.board_10[17] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6936_ (.RESET_B(net38),
    .D(_0430_),
    .Q(\vga_tetris.boardMem.board_10[18] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6937_ (.RESET_B(net37),
    .D(_0431_),
    .Q(\vga_tetris.boardMem.board_10[19] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6938_ (.RESET_B(net36),
    .D(_0432_),
    .Q(\vga_tetris.boardMem.board_11[0] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _6939_ (.RESET_B(net35),
    .D(_0433_),
    .Q(\vga_tetris.boardMem.board_11[1] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6940_ (.RESET_B(net34),
    .D(_0434_),
    .Q(\vga_tetris.boardMem.board_11[2] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6941_ (.RESET_B(net33),
    .D(net1311),
    .Q(\vga_tetris.boardMem.board_11[3] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6942_ (.RESET_B(net32),
    .D(_0436_),
    .Q(\vga_tetris.boardMem.board_11[4] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6943_ (.RESET_B(net31),
    .D(_0437_),
    .Q(\vga_tetris.boardMem.board_11[5] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6944_ (.RESET_B(net30),
    .D(_0438_),
    .Q(\vga_tetris.boardMem.board_11[6] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6945_ (.RESET_B(net29),
    .D(_0439_),
    .Q(\vga_tetris.boardMem.board_11[7] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6946_ (.RESET_B(net28),
    .D(_0440_),
    .Q(\vga_tetris.boardMem.board_11[8] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6947_ (.RESET_B(net27),
    .D(_0441_),
    .Q(\vga_tetris.boardMem.board_11[9] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6948_ (.RESET_B(net26),
    .D(_0442_),
    .Q(\vga_tetris.boardMem.board_11[10] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _6949_ (.RESET_B(net25),
    .D(_0443_),
    .Q(\vga_tetris.boardMem.board_11[11] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _6950_ (.RESET_B(net24),
    .D(_0444_),
    .Q(\vga_tetris.boardMem.board_11[12] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6951_ (.RESET_B(net23),
    .D(_0445_),
    .Q(\vga_tetris.boardMem.board_11[13] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6952_ (.RESET_B(net22),
    .D(_0446_),
    .Q(\vga_tetris.boardMem.board_11[14] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6953_ (.RESET_B(net21),
    .D(_0447_),
    .Q(\vga_tetris.boardMem.board_11[15] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6954_ (.RESET_B(net644),
    .D(_0448_),
    .Q(\vga_tetris.boardMem.board_11[16] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6955_ (.RESET_B(net643),
    .D(_0449_),
    .Q(\vga_tetris.boardMem.board_11[17] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6956_ (.RESET_B(net642),
    .D(_0450_),
    .Q(\vga_tetris.boardMem.board_11[18] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6957_ (.RESET_B(net641),
    .D(_0451_),
    .Q(\vga_tetris.boardMem.board_11[19] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6958_ (.RESET_B(net640),
    .D(net818),
    .Q(\vga_tetris.boardMem.board_12[0] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _6959_ (.RESET_B(net639),
    .D(net685),
    .Q(\vga_tetris.boardMem.board_12[1] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6960_ (.RESET_B(net638),
    .D(_0454_),
    .Q(\vga_tetris.boardMem.board_12[2] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6961_ (.RESET_B(net637),
    .D(_0455_),
    .Q(\vga_tetris.boardMem.board_12[3] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6962_ (.RESET_B(net636),
    .D(_0456_),
    .Q(\vga_tetris.boardMem.board_12[4] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6963_ (.RESET_B(net635),
    .D(_0457_),
    .Q(\vga_tetris.boardMem.board_12[5] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6964_ (.RESET_B(net634),
    .D(_0458_),
    .Q(\vga_tetris.boardMem.board_12[6] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6965_ (.RESET_B(net633),
    .D(_0459_),
    .Q(\vga_tetris.boardMem.board_12[7] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6966_ (.RESET_B(net632),
    .D(_0460_),
    .Q(\vga_tetris.boardMem.board_12[8] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6967_ (.RESET_B(net631),
    .D(_0461_),
    .Q(\vga_tetris.boardMem.board_12[9] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6968_ (.RESET_B(net630),
    .D(_0462_),
    .Q(\vga_tetris.boardMem.board_12[10] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _6969_ (.RESET_B(net629),
    .D(_0463_),
    .Q(\vga_tetris.boardMem.board_12[11] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _6970_ (.RESET_B(net628),
    .D(net1272),
    .Q(\vga_tetris.boardMem.board_12[12] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6971_ (.RESET_B(net627),
    .D(_0465_),
    .Q(\vga_tetris.boardMem.board_12[13] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6972_ (.RESET_B(net626),
    .D(_0466_),
    .Q(\vga_tetris.boardMem.board_12[14] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _6973_ (.RESET_B(net625),
    .D(_0467_),
    .Q(\vga_tetris.boardMem.board_12[15] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6974_ (.RESET_B(net624),
    .D(_0468_),
    .Q(\vga_tetris.boardMem.board_12[16] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6975_ (.RESET_B(net623),
    .D(_0469_),
    .Q(\vga_tetris.boardMem.board_12[17] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6976_ (.RESET_B(net622),
    .D(_0470_),
    .Q(\vga_tetris.boardMem.board_12[18] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6977_ (.RESET_B(net621),
    .D(net721),
    .Q(\vga_tetris.boardMem.board_12[19] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6978_ (.RESET_B(net620),
    .D(_0472_),
    .Q(\vga_tetris.boardMem.board_13[0] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6979_ (.RESET_B(net619),
    .D(_0473_),
    .Q(\vga_tetris.boardMem.board_13[1] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6980_ (.RESET_B(net618),
    .D(_0474_),
    .Q(\vga_tetris.boardMem.board_13[2] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6981_ (.RESET_B(net617),
    .D(_0475_),
    .Q(\vga_tetris.boardMem.board_13[3] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6982_ (.RESET_B(net616),
    .D(_0476_),
    .Q(\vga_tetris.boardMem.board_13[4] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6983_ (.RESET_B(net615),
    .D(_0477_),
    .Q(\vga_tetris.boardMem.board_13[5] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6984_ (.RESET_B(net614),
    .D(_0478_),
    .Q(\vga_tetris.boardMem.board_13[6] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6985_ (.RESET_B(net613),
    .D(_0479_),
    .Q(\vga_tetris.boardMem.board_13[7] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6986_ (.RESET_B(net612),
    .D(_0480_),
    .Q(\vga_tetris.boardMem.board_13[8] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6987_ (.RESET_B(net611),
    .D(_0481_),
    .Q(\vga_tetris.boardMem.board_13[9] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6988_ (.RESET_B(net610),
    .D(net738),
    .Q(\vga_tetris.boardMem.board_13[10] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _6989_ (.RESET_B(net609),
    .D(_0483_),
    .Q(\vga_tetris.boardMem.board_13[11] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _6990_ (.RESET_B(net608),
    .D(_0484_),
    .Q(\vga_tetris.boardMem.board_13[12] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6991_ (.RESET_B(net607),
    .D(_0485_),
    .Q(\vga_tetris.boardMem.board_13[13] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6992_ (.RESET_B(net606),
    .D(_0486_),
    .Q(\vga_tetris.boardMem.board_13[14] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6993_ (.RESET_B(net605),
    .D(_0487_),
    .Q(\vga_tetris.boardMem.board_13[15] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6994_ (.RESET_B(net604),
    .D(_0488_),
    .Q(\vga_tetris.boardMem.board_13[16] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6995_ (.RESET_B(net603),
    .D(net699),
    .Q(\vga_tetris.boardMem.board_13[17] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6996_ (.RESET_B(net602),
    .D(_0490_),
    .Q(\vga_tetris.boardMem.board_13[18] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6997_ (.RESET_B(net601),
    .D(_0491_),
    .Q(\vga_tetris.boardMem.board_13[19] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _6998_ (.RESET_B(net600),
    .D(_0492_),
    .Q(\vga_tetris.boardMem.board_14[0] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _6999_ (.RESET_B(net599),
    .D(_0493_),
    .Q(\vga_tetris.boardMem.board_14[1] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _7000_ (.RESET_B(net598),
    .D(_0494_),
    .Q(\vga_tetris.boardMem.board_14[2] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _7001_ (.RESET_B(net597),
    .D(_0495_),
    .Q(\vga_tetris.boardMem.board_14[3] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _7002_ (.RESET_B(net596),
    .D(_0496_),
    .Q(\vga_tetris.boardMem.board_14[4] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _7003_ (.RESET_B(net595),
    .D(net717),
    .Q(\vga_tetris.boardMem.board_14[5] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _7004_ (.RESET_B(net594),
    .D(_0498_),
    .Q(\vga_tetris.boardMem.board_14[6] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _7005_ (.RESET_B(net593),
    .D(_0499_),
    .Q(\vga_tetris.boardMem.board_14[7] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _7006_ (.RESET_B(net592),
    .D(_0500_),
    .Q(\vga_tetris.boardMem.board_14[8] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _7007_ (.RESET_B(net591),
    .D(_0501_),
    .Q(\vga_tetris.boardMem.board_14[9] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _7008_ (.RESET_B(net590),
    .D(_0502_),
    .Q(\vga_tetris.boardMem.board_14[10] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _7009_ (.RESET_B(net589),
    .D(_0503_),
    .Q(\vga_tetris.boardMem.board_14[11] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _7010_ (.RESET_B(net588),
    .D(_0504_),
    .Q(\vga_tetris.boardMem.board_14[12] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _7011_ (.RESET_B(net587),
    .D(_0505_),
    .Q(\vga_tetris.boardMem.board_14[13] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _7012_ (.RESET_B(net586),
    .D(_0506_),
    .Q(\vga_tetris.boardMem.board_14[14] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _7013_ (.RESET_B(net585),
    .D(_0507_),
    .Q(\vga_tetris.boardMem.board_14[15] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _7014_ (.RESET_B(net584),
    .D(_0508_),
    .Q(\vga_tetris.boardMem.board_14[16] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _7015_ (.RESET_B(net583),
    .D(_0509_),
    .Q(\vga_tetris.boardMem.board_14[17] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _7016_ (.RESET_B(net582),
    .D(_0510_),
    .Q(\vga_tetris.boardMem.board_14[18] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _7017_ (.RESET_B(net581),
    .D(_0511_),
    .Q(\vga_tetris.boardMem.board_14[19] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _7018_ (.RESET_B(net580),
    .D(_0512_),
    .Q(\vga_tetris.boardMem.board_15[0] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _7019_ (.RESET_B(net579),
    .D(_0513_),
    .Q(\vga_tetris.boardMem.board_15[1] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _7020_ (.RESET_B(net578),
    .D(_0514_),
    .Q(\vga_tetris.boardMem.board_15[2] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _7021_ (.RESET_B(net577),
    .D(_0515_),
    .Q(\vga_tetris.boardMem.board_15[3] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _7022_ (.RESET_B(net576),
    .D(_0516_),
    .Q(\vga_tetris.boardMem.board_15[4] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _7023_ (.RESET_B(net575),
    .D(net1302),
    .Q(\vga_tetris.boardMem.board_15[5] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _7024_ (.RESET_B(net574),
    .D(_0518_),
    .Q(\vga_tetris.boardMem.board_15[6] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _7025_ (.RESET_B(net573),
    .D(net1362),
    .Q(\vga_tetris.boardMem.board_15[7] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _7026_ (.RESET_B(net572),
    .D(_0520_),
    .Q(\vga_tetris.boardMem.board_15[8] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _7027_ (.RESET_B(net571),
    .D(_0521_),
    .Q(\vga_tetris.boardMem.board_15[9] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _7028_ (.RESET_B(net570),
    .D(_0522_),
    .Q(\vga_tetris.boardMem.board_15[10] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _7029_ (.RESET_B(net569),
    .D(_0523_),
    .Q(\vga_tetris.boardMem.board_15[11] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _7030_ (.RESET_B(net568),
    .D(net653),
    .Q(\vga_tetris.boardMem.board_15[12] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _7031_ (.RESET_B(net567),
    .D(_0525_),
    .Q(\vga_tetris.boardMem.board_15[13] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _7032_ (.RESET_B(net566),
    .D(_0526_),
    .Q(\vga_tetris.boardMem.board_15[14] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _7033_ (.RESET_B(net565),
    .D(_0527_),
    .Q(\vga_tetris.boardMem.board_15[15] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _7034_ (.RESET_B(net564),
    .D(_0528_),
    .Q(\vga_tetris.boardMem.board_15[16] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _7035_ (.RESET_B(net563),
    .D(net726),
    .Q(\vga_tetris.boardMem.board_15[17] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _7036_ (.RESET_B(net562),
    .D(_0530_),
    .Q(\vga_tetris.boardMem.board_15[18] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _7037_ (.RESET_B(net561),
    .D(_0531_),
    .Q(\vga_tetris.boardMem.board_15[19] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _7038_ (.RESET_B(net560),
    .D(net1445),
    .Q(\vga_tetris.boardMem.board_16[0] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _7039_ (.RESET_B(net559),
    .D(_0533_),
    .Q(\vga_tetris.boardMem.board_16[1] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _7040_ (.RESET_B(net558),
    .D(_0534_),
    .Q(\vga_tetris.boardMem.board_16[2] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _7041_ (.RESET_B(net557),
    .D(_0535_),
    .Q(\vga_tetris.boardMem.board_16[3] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _7042_ (.RESET_B(net556),
    .D(_0536_),
    .Q(\vga_tetris.boardMem.board_16[4] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _7043_ (.RESET_B(net555),
    .D(_0537_),
    .Q(\vga_tetris.boardMem.board_16[5] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _7044_ (.RESET_B(net554),
    .D(_0538_),
    .Q(\vga_tetris.boardMem.board_16[6] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _7045_ (.RESET_B(net553),
    .D(_0539_),
    .Q(\vga_tetris.boardMem.board_16[7] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _7046_ (.RESET_B(net552),
    .D(net1544),
    .Q(\vga_tetris.boardMem.board_16[8] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _7047_ (.RESET_B(net551),
    .D(net1481),
    .Q(\vga_tetris.boardMem.board_16[9] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _7048_ (.RESET_B(net550),
    .D(_0542_),
    .Q(\vga_tetris.boardMem.board_16[10] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _7049_ (.RESET_B(net549),
    .D(_0543_),
    .Q(\vga_tetris.boardMem.board_16[11] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _7050_ (.RESET_B(net547),
    .D(_0544_),
    .Q(\vga_tetris.boardMem.board_16[12] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _7051_ (.RESET_B(net545),
    .D(net1538),
    .Q(\vga_tetris.boardMem.board_16[13] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _7052_ (.RESET_B(net516),
    .D(_0546_),
    .Q(\vga_tetris.boardMem.board_16[14] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _7053_ (.RESET_B(net514),
    .D(_0547_),
    .Q(\vga_tetris.boardMem.board_16[15] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _7054_ (.RESET_B(net512),
    .D(net1420),
    .Q(\vga_tetris.boardMem.board_16[16] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _7055_ (.RESET_B(net510),
    .D(net1570),
    .Q(\vga_tetris.boardMem.board_16[17] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _7056_ (.RESET_B(net508),
    .D(_0550_),
    .Q(\vga_tetris.boardMem.board_16[18] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _7057_ (.RESET_B(net506),
    .D(net1436),
    .Q(\vga_tetris.boardMem.board_16[19] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _7058_ (.RESET_B(net504),
    .D(_0552_),
    .Q(\vga_tetris.boardMem.board_17[0] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _7059_ (.RESET_B(net502),
    .D(_0553_),
    .Q(\vga_tetris.boardMem.board_17[1] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _7060_ (.RESET_B(net500),
    .D(_0554_),
    .Q(\vga_tetris.boardMem.board_17[2] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _7061_ (.RESET_B(net498),
    .D(_0555_),
    .Q(\vga_tetris.boardMem.board_17[3] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _7062_ (.RESET_B(net496),
    .D(_0556_),
    .Q(\vga_tetris.boardMem.board_17[4] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _7063_ (.RESET_B(net494),
    .D(_0557_),
    .Q(\vga_tetris.boardMem.board_17[5] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _7064_ (.RESET_B(net484),
    .D(_0558_),
    .Q(\vga_tetris.boardMem.board_17[6] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _7065_ (.RESET_B(net482),
    .D(net1550),
    .Q(\vga_tetris.boardMem.board_17[7] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _7066_ (.RESET_B(net480),
    .D(_0560_),
    .Q(\vga_tetris.boardMem.board_17[8] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _7067_ (.RESET_B(net478),
    .D(_0561_),
    .Q(\vga_tetris.boardMem.board_17[9] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _7068_ (.RESET_B(net476),
    .D(_0562_),
    .Q(\vga_tetris.boardMem.board_17[10] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _7069_ (.RESET_B(net474),
    .D(net1416),
    .Q(\vga_tetris.boardMem.board_17[11] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _7070_ (.RESET_B(net472),
    .D(net1578),
    .Q(\vga_tetris.boardMem.board_17[12] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _7071_ (.RESET_B(net470),
    .D(_0565_),
    .Q(\vga_tetris.boardMem.board_17[13] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _7072_ (.RESET_B(net468),
    .D(_0566_),
    .Q(\vga_tetris.boardMem.board_17[14] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _7073_ (.RESET_B(net466),
    .D(net1409),
    .Q(\vga_tetris.boardMem.board_17[15] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _7074_ (.RESET_B(net464),
    .D(_0568_),
    .Q(\vga_tetris.boardMem.board_17[16] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _7075_ (.RESET_B(net462),
    .D(_0569_),
    .Q(\vga_tetris.boardMem.board_17[17] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _7076_ (.RESET_B(net460),
    .D(_0570_),
    .Q(\vga_tetris.boardMem.board_17[18] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _7077_ (.RESET_B(net458),
    .D(_0571_),
    .Q(\vga_tetris.boardMem.board_17[19] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _7078_ (.RESET_B(net456),
    .D(_0572_),
    .Q(\vga_tetris.boardMem.board_18[0] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _7079_ (.RESET_B(net454),
    .D(_0573_),
    .Q(\vga_tetris.boardMem.board_18[1] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _7080_ (.RESET_B(net449),
    .D(_0574_),
    .Q(\vga_tetris.boardMem.board_18[2] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _7081_ (.RESET_B(net447),
    .D(_0575_),
    .Q(\vga_tetris.boardMem.board_18[3] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _7082_ (.RESET_B(net445),
    .D(_0576_),
    .Q(\vga_tetris.boardMem.board_18[4] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _7083_ (.RESET_B(net443),
    .D(_0577_),
    .Q(\vga_tetris.boardMem.board_18[5] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _7084_ (.RESET_B(net441),
    .D(_0578_),
    .Q(\vga_tetris.boardMem.board_18[6] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _7085_ (.RESET_B(net439),
    .D(_0579_),
    .Q(\vga_tetris.boardMem.board_18[7] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _7086_ (.RESET_B(net437),
    .D(_0580_),
    .Q(\vga_tetris.boardMem.board_18[8] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _7087_ (.RESET_B(net435),
    .D(net1449),
    .Q(\vga_tetris.boardMem.board_18[9] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _7088_ (.RESET_B(net433),
    .D(_0582_),
    .Q(\vga_tetris.boardMem.board_18[10] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _7089_ (.RESET_B(net431),
    .D(_0583_),
    .Q(\vga_tetris.boardMem.board_18[11] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _7090_ (.RESET_B(net429),
    .D(_0584_),
    .Q(\vga_tetris.boardMem.board_18[12] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _7091_ (.RESET_B(net427),
    .D(_0585_),
    .Q(\vga_tetris.boardMem.board_18[13] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _7092_ (.RESET_B(net425),
    .D(_0586_),
    .Q(\vga_tetris.boardMem.board_18[14] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _7093_ (.RESET_B(net423),
    .D(_0587_),
    .Q(\vga_tetris.boardMem.board_18[15] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _7094_ (.RESET_B(net421),
    .D(_0588_),
    .Q(\vga_tetris.boardMem.board_18[16] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _7095_ (.RESET_B(net419),
    .D(_0589_),
    .Q(\vga_tetris.boardMem.board_18[17] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _7096_ (.RESET_B(net417),
    .D(_0590_),
    .Q(\vga_tetris.boardMem.board_18[18] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _7097_ (.RESET_B(net415),
    .D(_0591_),
    .Q(\vga_tetris.boardMem.board_18[19] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _7098_ (.RESET_B(net413),
    .D(net1613),
    .Q(\vga_tetris.tetrisLogic.shiftTheBoard.internalStartTriggerQ ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _7099_ (.RESET_B(net411),
    .D(net1479),
    .Q(\vga_tetris.vgaController.verticalCounterQ[0] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _7100_ (.RESET_B(net407),
    .D(_0594_),
    .Q(\vga_tetris.vgaController.verticalCounterQ[1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _7101_ (.RESET_B(net400),
    .D(net1607),
    .Q(\vga_tetris.vgaController.verticalCounterQ[2] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _7102_ (.RESET_B(net385),
    .D(net1594),
    .Q(\vga_tetris.vgaController.verticalCounterQ[3] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _7103_ (.RESET_B(net381),
    .D(_0597_),
    .Q(\vga_tetris.vgaController.verticalCounterQ[4] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _7104_ (.RESET_B(net374),
    .D(_0598_),
    .Q(\vga_tetris.vgaController.verticalCounterQ[5] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _7105_ (.RESET_B(net370),
    .D(_0599_),
    .Q(\vga_tetris.vgaController.verticalCounterQ[6] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _7106_ (.RESET_B(net366),
    .D(_0600_),
    .Q(\vga_tetris.vgaController.verticalCounterQ[7] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _7107_ (.RESET_B(net362),
    .D(net1603),
    .Q(\vga_tetris.vgaController.verticalCounterQ[8] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _7108_ (.RESET_B(net358),
    .D(_0602_),
    .Q(\vga_tetris.vgaController.verticalCounterQ[9] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _7109_ (.RESET_B(net354),
    .D(_0603_),
    .Q(\vga_tetris._vgaController_io_pixelPosX[0] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _7110_ (.RESET_B(net350),
    .D(net1600),
    .Q(\vga_tetris._vgaController_io_pixelPosX[1] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _7111_ (.RESET_B(net346),
    .D(_0605_),
    .Q(\vga_tetris._vgaController_io_pixelPosX[2] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _7112_ (.RESET_B(net342),
    .D(net1783),
    .Q(\vga_tetris._vgaController_io_pixelPosX[3] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _7113_ (.RESET_B(net338),
    .D(_0607_),
    .Q(\vga_tetris._vgaController_io_pixelPosX[4] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _7114_ (.RESET_B(net330),
    .D(net1860),
    .Q(\vga_tetris._vgaController_io_pixelPosX[5] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _7115_ (.RESET_B(net409),
    .D(_0609_),
    .Q(\vga_tetris._vgaController_io_pixelPosX[6] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _7116_ (.RESET_B(net387),
    .D(_0610_),
    .Q(\vga_tetris._vgaController_io_pixelPosX[7] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _7117_ (.RESET_B(net379),
    .D(net1580),
    .Q(\vga_tetris._vgaController_io_pixelPosX[8] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _7118_ (.RESET_B(net368),
    .D(_0612_),
    .Q(\vga_tetris._vgaController_io_pixelPosX[9] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _7119_ (.RESET_B(net360),
    .D(_0613_),
    .Q(\vga_tetris._vgaController_io_pixelPosY[0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _7120_ (.RESET_B(net352),
    .D(_0614_),
    .Q(\vga_tetris._vgaController_io_pixelPosY[1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _7121_ (.RESET_B(net344),
    .D(_0615_),
    .Q(\vga_tetris._vgaController_io_pixelPosY[2] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _7122_ (.RESET_B(net336),
    .D(_0616_),
    .Q(\vga_tetris._vgaController_io_pixelPosY[3] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _7123_ (.RESET_B(net402),
    .D(_0617_),
    .Q(\vga_tetris._tetrisDisplay_io_boardYCoord[0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _7124_ (.RESET_B(net372),
    .D(_0618_),
    .Q(\vga_tetris._tetrisDisplay_io_boardYCoord[1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _7125_ (.RESET_B(net356),
    .D(_0619_),
    .Q(\vga_tetris._vgaController_io_pixelPosY[6] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _7126_ (.RESET_B(net340),
    .D(net1704),
    .Q(\vga_tetris._vgaController_io_pixelPosY[7] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _7127_ (.RESET_B(net383),
    .D(net1641),
    .Q(\vga_tetris._vgaController_io_pixelPosY[8] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _7128_ (.RESET_B(net348),
    .D(_0622_),
    .Q(\vga_tetris._vgaController_io_pixelPosY[9] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _7129_ (.RESET_B(net364),
    .D(_0623_),
    .Q(\vga_tetris.runningTetrisLogicQ ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_tiehi _6952__22 (.L_HI(net22));
 sg13g2_tiehi _6951__23 (.L_HI(net23));
 sg13g2_tiehi _6950__24 (.L_HI(net24));
 sg13g2_tiehi _6949__25 (.L_HI(net25));
 sg13g2_tiehi _6948__26 (.L_HI(net26));
 sg13g2_tiehi _6947__27 (.L_HI(net27));
 sg13g2_tiehi _6946__28 (.L_HI(net28));
 sg13g2_tiehi _6945__29 (.L_HI(net29));
 sg13g2_tiehi _6944__30 (.L_HI(net30));
 sg13g2_tiehi _6943__31 (.L_HI(net31));
 sg13g2_tiehi _6942__32 (.L_HI(net32));
 sg13g2_tiehi _6941__33 (.L_HI(net33));
 sg13g2_tiehi _6940__34 (.L_HI(net34));
 sg13g2_tiehi _6939__35 (.L_HI(net35));
 sg13g2_tiehi _6938__36 (.L_HI(net36));
 sg13g2_tiehi _6937__37 (.L_HI(net37));
 sg13g2_tiehi _6936__38 (.L_HI(net38));
 sg13g2_tiehi _6935__39 (.L_HI(net39));
 sg13g2_tiehi _6934__40 (.L_HI(net40));
 sg13g2_tiehi _6933__41 (.L_HI(net41));
 sg13g2_tiehi _6932__42 (.L_HI(net42));
 sg13g2_tiehi _6931__43 (.L_HI(net43));
 sg13g2_tiehi _6930__44 (.L_HI(net44));
 sg13g2_tiehi _6929__45 (.L_HI(net45));
 sg13g2_tiehi _6928__46 (.L_HI(net46));
 sg13g2_tiehi _6927__47 (.L_HI(net47));
 sg13g2_tiehi _6926__48 (.L_HI(net48));
 sg13g2_tiehi _6925__49 (.L_HI(net49));
 sg13g2_tiehi _6924__50 (.L_HI(net50));
 sg13g2_tiehi _6923__51 (.L_HI(net51));
 sg13g2_tiehi _6922__52 (.L_HI(net52));
 sg13g2_tiehi _6921__53 (.L_HI(net53));
 sg13g2_tiehi _6920__54 (.L_HI(net54));
 sg13g2_tiehi _6919__55 (.L_HI(net55));
 sg13g2_tiehi _6918__56 (.L_HI(net56));
 sg13g2_tiehi _6917__57 (.L_HI(net57));
 sg13g2_tiehi _6916__58 (.L_HI(net58));
 sg13g2_tiehi _6915__59 (.L_HI(net59));
 sg13g2_tiehi _6914__60 (.L_HI(net60));
 sg13g2_tiehi _6913__61 (.L_HI(net61));
 sg13g2_tiehi _6912__62 (.L_HI(net62));
 sg13g2_tiehi _6911__63 (.L_HI(net63));
 sg13g2_tiehi _6910__64 (.L_HI(net64));
 sg13g2_tiehi _6909__65 (.L_HI(net65));
 sg13g2_tiehi _6908__66 (.L_HI(net66));
 sg13g2_tiehi _6907__67 (.L_HI(net67));
 sg13g2_tiehi _6906__68 (.L_HI(net68));
 sg13g2_tiehi _6905__69 (.L_HI(net69));
 sg13g2_tiehi _6904__70 (.L_HI(net70));
 sg13g2_tiehi _6903__71 (.L_HI(net71));
 sg13g2_tiehi _6902__72 (.L_HI(net72));
 sg13g2_tiehi _6901__73 (.L_HI(net73));
 sg13g2_tiehi _6900__74 (.L_HI(net74));
 sg13g2_tiehi _6899__75 (.L_HI(net75));
 sg13g2_tiehi _6898__76 (.L_HI(net76));
 sg13g2_tiehi _6897__77 (.L_HI(net77));
 sg13g2_tiehi _6896__78 (.L_HI(net78));
 sg13g2_tiehi _6895__79 (.L_HI(net79));
 sg13g2_tiehi _6894__80 (.L_HI(net80));
 sg13g2_tiehi _6893__81 (.L_HI(net81));
 sg13g2_tiehi _6892__82 (.L_HI(net82));
 sg13g2_tiehi _6891__83 (.L_HI(net83));
 sg13g2_tiehi _6890__84 (.L_HI(net84));
 sg13g2_tiehi _6889__85 (.L_HI(net85));
 sg13g2_tiehi _6888__86 (.L_HI(net86));
 sg13g2_tiehi _6887__87 (.L_HI(net87));
 sg13g2_tiehi _6886__88 (.L_HI(net88));
 sg13g2_tiehi _6885__89 (.L_HI(net89));
 sg13g2_tiehi _6884__90 (.L_HI(net90));
 sg13g2_tiehi _6883__91 (.L_HI(net91));
 sg13g2_tiehi _6882__92 (.L_HI(net92));
 sg13g2_tiehi _6881__93 (.L_HI(net93));
 sg13g2_tiehi _6880__94 (.L_HI(net94));
 sg13g2_tiehi _6879__95 (.L_HI(net95));
 sg13g2_tiehi _6878__96 (.L_HI(net96));
 sg13g2_tiehi _6877__97 (.L_HI(net97));
 sg13g2_tiehi _6876__98 (.L_HI(net98));
 sg13g2_tiehi _6875__99 (.L_HI(net99));
 sg13g2_tiehi _6874__100 (.L_HI(net100));
 sg13g2_tiehi _6873__101 (.L_HI(net101));
 sg13g2_tiehi _6872__102 (.L_HI(net102));
 sg13g2_tiehi _6871__103 (.L_HI(net103));
 sg13g2_tiehi _6870__104 (.L_HI(net104));
 sg13g2_tiehi _6869__105 (.L_HI(net105));
 sg13g2_tiehi _6868__106 (.L_HI(net106));
 sg13g2_tiehi _6867__107 (.L_HI(net107));
 sg13g2_tiehi _6866__108 (.L_HI(net108));
 sg13g2_tiehi _6865__109 (.L_HI(net109));
 sg13g2_tiehi _6864__110 (.L_HI(net110));
 sg13g2_tiehi _6863__111 (.L_HI(net111));
 sg13g2_tiehi _6862__112 (.L_HI(net112));
 sg13g2_tiehi _6861__113 (.L_HI(net113));
 sg13g2_tiehi _6860__114 (.L_HI(net114));
 sg13g2_tiehi _6859__115 (.L_HI(net115));
 sg13g2_tiehi _6858__116 (.L_HI(net116));
 sg13g2_tiehi _6857__117 (.L_HI(net117));
 sg13g2_tiehi _6856__118 (.L_HI(net118));
 sg13g2_tiehi _6855__119 (.L_HI(net119));
 sg13g2_tiehi _6854__120 (.L_HI(net120));
 sg13g2_tiehi _6853__121 (.L_HI(net121));
 sg13g2_tiehi _6852__122 (.L_HI(net122));
 sg13g2_tiehi _6851__123 (.L_HI(net123));
 sg13g2_tiehi _6850__124 (.L_HI(net124));
 sg13g2_tiehi _6849__125 (.L_HI(net125));
 sg13g2_tiehi _6848__126 (.L_HI(net126));
 sg13g2_tiehi _6847__127 (.L_HI(net127));
 sg13g2_tiehi _6846__128 (.L_HI(net128));
 sg13g2_tiehi _6845__129 (.L_HI(net129));
 sg13g2_tiehi _6844__130 (.L_HI(net130));
 sg13g2_tiehi _6843__131 (.L_HI(net131));
 sg13g2_tiehi _6842__132 (.L_HI(net132));
 sg13g2_tiehi _6841__133 (.L_HI(net133));
 sg13g2_tiehi _6840__134 (.L_HI(net134));
 sg13g2_tiehi _6839__135 (.L_HI(net135));
 sg13g2_tiehi _6838__136 (.L_HI(net136));
 sg13g2_tiehi _6837__137 (.L_HI(net137));
 sg13g2_tiehi _6836__138 (.L_HI(net138));
 sg13g2_tiehi _6835__139 (.L_HI(net139));
 sg13g2_tiehi _6834__140 (.L_HI(net140));
 sg13g2_tiehi _6833__141 (.L_HI(net141));
 sg13g2_tiehi _6832__142 (.L_HI(net142));
 sg13g2_tiehi _6831__143 (.L_HI(net143));
 sg13g2_tiehi _6830__144 (.L_HI(net144));
 sg13g2_tiehi _6829__145 (.L_HI(net145));
 sg13g2_tiehi _6828__146 (.L_HI(net146));
 sg13g2_tiehi _6827__147 (.L_HI(net147));
 sg13g2_tiehi _6826__148 (.L_HI(net148));
 sg13g2_tiehi _6825__149 (.L_HI(net149));
 sg13g2_tiehi _6824__150 (.L_HI(net150));
 sg13g2_tiehi _6823__151 (.L_HI(net151));
 sg13g2_tiehi _6822__152 (.L_HI(net152));
 sg13g2_tiehi _6821__153 (.L_HI(net153));
 sg13g2_tiehi _6820__154 (.L_HI(net154));
 sg13g2_tiehi _6819__155 (.L_HI(net155));
 sg13g2_tiehi _6818__156 (.L_HI(net156));
 sg13g2_tiehi _6817__157 (.L_HI(net157));
 sg13g2_tiehi _6816__158 (.L_HI(net158));
 sg13g2_tiehi _6815__159 (.L_HI(net159));
 sg13g2_tiehi _6814__160 (.L_HI(net160));
 sg13g2_tiehi _6813__161 (.L_HI(net161));
 sg13g2_tiehi _6812__162 (.L_HI(net162));
 sg13g2_tiehi _6811__163 (.L_HI(net163));
 sg13g2_tiehi _6810__164 (.L_HI(net164));
 sg13g2_tiehi _6809__165 (.L_HI(net165));
 sg13g2_tiehi _6808__166 (.L_HI(net166));
 sg13g2_tiehi _6807__167 (.L_HI(net167));
 sg13g2_tiehi _6806__168 (.L_HI(net168));
 sg13g2_tiehi _6805__169 (.L_HI(net169));
 sg13g2_tiehi _6804__170 (.L_HI(net170));
 sg13g2_tiehi _6803__171 (.L_HI(net171));
 sg13g2_tiehi _6802__172 (.L_HI(net172));
 sg13g2_tiehi _6801__173 (.L_HI(net173));
 sg13g2_tiehi _6800__174 (.L_HI(net174));
 sg13g2_tiehi _6799__175 (.L_HI(net175));
 sg13g2_tiehi _6798__176 (.L_HI(net176));
 sg13g2_tiehi _6797__177 (.L_HI(net177));
 sg13g2_tiehi _6796__178 (.L_HI(net178));
 sg13g2_tiehi _6795__179 (.L_HI(net179));
 sg13g2_tiehi _6794__180 (.L_HI(net180));
 sg13g2_tiehi _6793__181 (.L_HI(net181));
 sg13g2_tiehi _6792__182 (.L_HI(net182));
 sg13g2_tiehi _6791__183 (.L_HI(net183));
 sg13g2_tiehi _6790__184 (.L_HI(net184));
 sg13g2_tiehi _6789__185 (.L_HI(net185));
 sg13g2_tiehi _6788__186 (.L_HI(net186));
 sg13g2_tiehi _6787__187 (.L_HI(net187));
 sg13g2_tiehi _6786__188 (.L_HI(net188));
 sg13g2_tiehi _6785__189 (.L_HI(net189));
 sg13g2_tiehi _6784__190 (.L_HI(net190));
 sg13g2_tiehi _6783__191 (.L_HI(net191));
 sg13g2_tiehi _6782__192 (.L_HI(net192));
 sg13g2_tiehi _6781__193 (.L_HI(net193));
 sg13g2_tiehi _6780__194 (.L_HI(net194));
 sg13g2_tiehi _6779__195 (.L_HI(net195));
 sg13g2_tiehi _6778__196 (.L_HI(net196));
 sg13g2_tiehi _6777__197 (.L_HI(net197));
 sg13g2_tiehi _6776__198 (.L_HI(net198));
 sg13g2_tiehi _6775__199 (.L_HI(net199));
 sg13g2_tiehi _6774__200 (.L_HI(net200));
 sg13g2_tiehi _6773__201 (.L_HI(net201));
 sg13g2_tiehi _6772__202 (.L_HI(net202));
 sg13g2_tiehi _6771__203 (.L_HI(net203));
 sg13g2_tiehi _6770__204 (.L_HI(net204));
 sg13g2_tiehi _6769__205 (.L_HI(net205));
 sg13g2_tiehi _6768__206 (.L_HI(net206));
 sg13g2_tiehi _6767__207 (.L_HI(net207));
 sg13g2_tiehi _6766__208 (.L_HI(net208));
 sg13g2_tiehi _6765__209 (.L_HI(net209));
 sg13g2_tiehi _6764__210 (.L_HI(net210));
 sg13g2_tiehi _6763__211 (.L_HI(net211));
 sg13g2_tiehi _6762__212 (.L_HI(net212));
 sg13g2_tiehi _6761__213 (.L_HI(net213));
 sg13g2_tiehi _6760__214 (.L_HI(net214));
 sg13g2_tiehi _6759__215 (.L_HI(net215));
 sg13g2_tiehi _6758__216 (.L_HI(net216));
 sg13g2_tiehi _6757__217 (.L_HI(net217));
 sg13g2_tiehi _6756__218 (.L_HI(net218));
 sg13g2_tiehi _6755__219 (.L_HI(net219));
 sg13g2_tiehi _6754__220 (.L_HI(net220));
 sg13g2_tiehi _6753__221 (.L_HI(net221));
 sg13g2_tiehi _6752__222 (.L_HI(net222));
 sg13g2_tiehi _6751__223 (.L_HI(net223));
 sg13g2_tiehi _6750__224 (.L_HI(net224));
 sg13g2_tiehi _6749__225 (.L_HI(net225));
 sg13g2_tiehi _6748__226 (.L_HI(net226));
 sg13g2_tiehi _6747__227 (.L_HI(net227));
 sg13g2_tiehi _6746__228 (.L_HI(net228));
 sg13g2_tiehi _6745__229 (.L_HI(net229));
 sg13g2_tiehi _6744__230 (.L_HI(net230));
 sg13g2_tiehi _6743__231 (.L_HI(net231));
 sg13g2_tiehi _6742__232 (.L_HI(net232));
 sg13g2_tiehi _6741__233 (.L_HI(net233));
 sg13g2_tiehi _6740__234 (.L_HI(net234));
 sg13g2_tiehi _6739__235 (.L_HI(net235));
 sg13g2_tiehi _6738__236 (.L_HI(net236));
 sg13g2_tiehi _6737__237 (.L_HI(net237));
 sg13g2_tiehi _6736__238 (.L_HI(net238));
 sg13g2_tiehi _6735__239 (.L_HI(net239));
 sg13g2_tiehi _6734__240 (.L_HI(net240));
 sg13g2_tiehi _6733__241 (.L_HI(net241));
 sg13g2_tiehi _6732__242 (.L_HI(net242));
 sg13g2_tiehi _6731__243 (.L_HI(net243));
 sg13g2_tiehi _6730__244 (.L_HI(net244));
 sg13g2_tiehi _6729__245 (.L_HI(net245));
 sg13g2_tiehi _6728__246 (.L_HI(net246));
 sg13g2_tiehi _6727__247 (.L_HI(net247));
 sg13g2_tiehi _6726__248 (.L_HI(net248));
 sg13g2_tiehi _6725__249 (.L_HI(net249));
 sg13g2_tiehi _6724__250 (.L_HI(net250));
 sg13g2_tiehi _6723__251 (.L_HI(net251));
 sg13g2_tiehi _6722__252 (.L_HI(net252));
 sg13g2_tiehi _6721__253 (.L_HI(net253));
 sg13g2_tiehi _6720__254 (.L_HI(net254));
 sg13g2_tiehi _6719__255 (.L_HI(net255));
 sg13g2_tiehi _6718__256 (.L_HI(net256));
 sg13g2_tiehi _6717__257 (.L_HI(net257));
 sg13g2_tiehi _6716__258 (.L_HI(net258));
 sg13g2_tiehi _6715__259 (.L_HI(net259));
 sg13g2_tiehi _6714__260 (.L_HI(net260));
 sg13g2_tiehi _6713__261 (.L_HI(net261));
 sg13g2_tiehi _6712__262 (.L_HI(net262));
 sg13g2_tiehi _6711__263 (.L_HI(net263));
 sg13g2_tiehi _6710__264 (.L_HI(net264));
 sg13g2_tiehi _6709__265 (.L_HI(net265));
 sg13g2_tiehi _6708__266 (.L_HI(net266));
 sg13g2_tiehi _6707__267 (.L_HI(net267));
 sg13g2_tiehi _6706__268 (.L_HI(net268));
 sg13g2_tiehi _6705__269 (.L_HI(net269));
 sg13g2_tiehi _6704__270 (.L_HI(net270));
 sg13g2_tiehi _6703__271 (.L_HI(net271));
 sg13g2_tiehi _6702__272 (.L_HI(net272));
 sg13g2_tiehi _6701__273 (.L_HI(net273));
 sg13g2_tiehi _6700__274 (.L_HI(net274));
 sg13g2_tiehi _6699__275 (.L_HI(net275));
 sg13g2_tiehi _6698__276 (.L_HI(net276));
 sg13g2_tiehi _6697__277 (.L_HI(net277));
 sg13g2_tiehi _6696__278 (.L_HI(net278));
 sg13g2_tiehi _6695__279 (.L_HI(net279));
 sg13g2_tiehi _6694__280 (.L_HI(net280));
 sg13g2_tiehi _6693__281 (.L_HI(net281));
 sg13g2_tiehi _6692__282 (.L_HI(net282));
 sg13g2_tiehi _6691__283 (.L_HI(net283));
 sg13g2_tiehi _6690__284 (.L_HI(net284));
 sg13g2_tiehi _6689__285 (.L_HI(net285));
 sg13g2_tiehi _6688__286 (.L_HI(net286));
 sg13g2_tiehi _6687__287 (.L_HI(net287));
 sg13g2_tiehi _6686__288 (.L_HI(net288));
 sg13g2_tiehi _6685__289 (.L_HI(net289));
 sg13g2_tiehi _6684__290 (.L_HI(net290));
 sg13g2_tiehi _6683__291 (.L_HI(net291));
 sg13g2_tiehi _6682__292 (.L_HI(net292));
 sg13g2_tiehi _6681__293 (.L_HI(net293));
 sg13g2_tiehi _6680__294 (.L_HI(net294));
 sg13g2_tiehi _6679__295 (.L_HI(net295));
 sg13g2_tiehi _6678__296 (.L_HI(net296));
 sg13g2_tiehi _6677__297 (.L_HI(net297));
 sg13g2_tiehi _6676__298 (.L_HI(net298));
 sg13g2_tiehi _6675__299 (.L_HI(net299));
 sg13g2_tiehi _6674__300 (.L_HI(net300));
 sg13g2_tiehi _6673__301 (.L_HI(net301));
 sg13g2_tiehi _6672__302 (.L_HI(net302));
 sg13g2_tiehi _6671__303 (.L_HI(net303));
 sg13g2_tiehi _6670__304 (.L_HI(net304));
 sg13g2_tiehi _6669__305 (.L_HI(net305));
 sg13g2_tiehi _6668__306 (.L_HI(net306));
 sg13g2_tiehi _6667__307 (.L_HI(net307));
 sg13g2_tiehi _6666__308 (.L_HI(net308));
 sg13g2_tiehi _6665__309 (.L_HI(net309));
 sg13g2_tiehi _6664__310 (.L_HI(net310));
 sg13g2_tiehi _6663__311 (.L_HI(net311));
 sg13g2_tiehi _6662__312 (.L_HI(net312));
 sg13g2_tiehi _6661__313 (.L_HI(net313));
 sg13g2_tiehi _6660__314 (.L_HI(net314));
 sg13g2_tiehi _6659__315 (.L_HI(net315));
 sg13g2_tiehi _6658__316 (.L_HI(net316));
 sg13g2_tiehi _6657__317 (.L_HI(net317));
 sg13g2_tiehi _6656__318 (.L_HI(net318));
 sg13g2_tiehi _6655__319 (.L_HI(net319));
 sg13g2_tiehi _6654__320 (.L_HI(net320));
 sg13g2_tiehi _6653__321 (.L_HI(net321));
 sg13g2_tiehi _6652__322 (.L_HI(net322));
 sg13g2_tiehi _6651__323 (.L_HI(net323));
 sg13g2_tiehi _6650__324 (.L_HI(net324));
 sg13g2_tiehi _6649__325 (.L_HI(net325));
 sg13g2_tiehi _6648__326 (.L_HI(net326));
 sg13g2_tiehi _6647__327 (.L_HI(net327));
 sg13g2_tiehi _6506__328 (.L_HI(net328));
 sg13g2_tiehi _6646__329 (.L_HI(net329));
 sg13g2_tiehi _7114__330 (.L_HI(net330));
 sg13g2_tiehi _6645__331 (.L_HI(net331));
 sg13g2_tiehi _6644__332 (.L_HI(net332));
 sg13g2_tiehi _6643__333 (.L_HI(net333));
 sg13g2_tiehi _6642__334 (.L_HI(net334));
 sg13g2_tiehi _6641__335 (.L_HI(net335));
 sg13g2_tiehi _7122__336 (.L_HI(net336));
 sg13g2_tiehi _6640__337 (.L_HI(net337));
 sg13g2_tiehi _7113__338 (.L_HI(net338));
 sg13g2_tiehi _6639__339 (.L_HI(net339));
 sg13g2_tiehi _7126__340 (.L_HI(net340));
 sg13g2_tiehi _6638__341 (.L_HI(net341));
 sg13g2_tiehi _7112__342 (.L_HI(net342));
 sg13g2_tiehi _6637__343 (.L_HI(net343));
 sg13g2_tiehi _7121__344 (.L_HI(net344));
 sg13g2_tiehi _6636__345 (.L_HI(net345));
 sg13g2_tiehi _7111__346 (.L_HI(net346));
 sg13g2_tiehi _6635__347 (.L_HI(net347));
 sg13g2_tiehi _7128__348 (.L_HI(net348));
 sg13g2_tiehi _6634__349 (.L_HI(net349));
 sg13g2_tiehi _7110__350 (.L_HI(net350));
 sg13g2_tiehi _6633__351 (.L_HI(net351));
 sg13g2_tiehi _7120__352 (.L_HI(net352));
 sg13g2_tiehi _6632__353 (.L_HI(net353));
 sg13g2_tiehi _7109__354 (.L_HI(net354));
 sg13g2_tiehi _6631__355 (.L_HI(net355));
 sg13g2_tiehi _7125__356 (.L_HI(net356));
 sg13g2_tiehi _6630__357 (.L_HI(net357));
 sg13g2_tiehi _7108__358 (.L_HI(net358));
 sg13g2_tiehi _6629__359 (.L_HI(net359));
 sg13g2_tiehi _7119__360 (.L_HI(net360));
 sg13g2_tiehi _6628__361 (.L_HI(net361));
 sg13g2_tiehi _7107__362 (.L_HI(net362));
 sg13g2_tiehi _6627__363 (.L_HI(net363));
 sg13g2_tiehi _7129__364 (.L_HI(net364));
 sg13g2_tiehi _6626__365 (.L_HI(net365));
 sg13g2_tiehi _7106__366 (.L_HI(net366));
 sg13g2_tiehi _6625__367 (.L_HI(net367));
 sg13g2_tiehi _7118__368 (.L_HI(net368));
 sg13g2_tiehi _6624__369 (.L_HI(net369));
 sg13g2_tiehi _7105__370 (.L_HI(net370));
 sg13g2_tiehi _6623__371 (.L_HI(net371));
 sg13g2_tiehi _7124__372 (.L_HI(net372));
 sg13g2_tiehi _6622__373 (.L_HI(net373));
 sg13g2_tiehi _7104__374 (.L_HI(net374));
 sg13g2_tiehi _6621__375 (.L_HI(net375));
 sg13g2_tiehi _6620__376 (.L_HI(net376));
 sg13g2_tiehi _6619__377 (.L_HI(net377));
 sg13g2_tiehi _6618__378 (.L_HI(net378));
 sg13g2_tiehi _7117__379 (.L_HI(net379));
 sg13g2_tiehi _6617__380 (.L_HI(net380));
 sg13g2_tiehi _7103__381 (.L_HI(net381));
 sg13g2_tiehi _6616__382 (.L_HI(net382));
 sg13g2_tiehi _7127__383 (.L_HI(net383));
 sg13g2_tiehi _6615__384 (.L_HI(net384));
 sg13g2_tiehi _7102__385 (.L_HI(net385));
 sg13g2_tiehi _6614__386 (.L_HI(net386));
 sg13g2_tiehi _7116__387 (.L_HI(net387));
 sg13g2_tiehi _6613__388 (.L_HI(net388));
 sg13g2_tiehi _6612__389 (.L_HI(net389));
 sg13g2_tiehi _6611__390 (.L_HI(net390));
 sg13g2_tiehi _6610__391 (.L_HI(net391));
 sg13g2_tiehi _6609__392 (.L_HI(net392));
 sg13g2_tiehi _6608__393 (.L_HI(net393));
 sg13g2_tiehi _6607__394 (.L_HI(net394));
 sg13g2_tiehi _6606__395 (.L_HI(net395));
 sg13g2_tiehi _6605__396 (.L_HI(net396));
 sg13g2_tiehi _6604__397 (.L_HI(net397));
 sg13g2_tiehi _6603__398 (.L_HI(net398));
 sg13g2_tiehi _6602__399 (.L_HI(net399));
 sg13g2_tiehi _7101__400 (.L_HI(net400));
 sg13g2_tiehi _6601__401 (.L_HI(net401));
 sg13g2_tiehi _7123__402 (.L_HI(net402));
 sg13g2_tiehi _6600__403 (.L_HI(net403));
 sg13g2_tiehi _6599__404 (.L_HI(net404));
 sg13g2_tiehi _6598__405 (.L_HI(net405));
 sg13g2_tiehi _6597__406 (.L_HI(net406));
 sg13g2_tiehi _7100__407 (.L_HI(net407));
 sg13g2_tiehi _6596__408 (.L_HI(net408));
 sg13g2_tiehi _7115__409 (.L_HI(net409));
 sg13g2_tiehi _6595__410 (.L_HI(net410));
 sg13g2_tiehi _7099__411 (.L_HI(net411));
 sg13g2_tiehi _6594__412 (.L_HI(net412));
 sg13g2_tiehi _7098__413 (.L_HI(net413));
 sg13g2_tiehi _6593__414 (.L_HI(net414));
 sg13g2_tiehi _7097__415 (.L_HI(net415));
 sg13g2_tiehi _6592__416 (.L_HI(net416));
 sg13g2_tiehi _7096__417 (.L_HI(net417));
 sg13g2_tiehi _6591__418 (.L_HI(net418));
 sg13g2_tiehi _7095__419 (.L_HI(net419));
 sg13g2_tiehi _6590__420 (.L_HI(net420));
 sg13g2_tiehi _7094__421 (.L_HI(net421));
 sg13g2_tiehi _6589__422 (.L_HI(net422));
 sg13g2_tiehi _7093__423 (.L_HI(net423));
 sg13g2_tiehi _6588__424 (.L_HI(net424));
 sg13g2_tiehi _7092__425 (.L_HI(net425));
 sg13g2_tiehi _6587__426 (.L_HI(net426));
 sg13g2_tiehi _7091__427 (.L_HI(net427));
 sg13g2_tiehi _6586__428 (.L_HI(net428));
 sg13g2_tiehi _7090__429 (.L_HI(net429));
 sg13g2_tiehi _6585__430 (.L_HI(net430));
 sg13g2_tiehi _7089__431 (.L_HI(net431));
 sg13g2_tiehi _6584__432 (.L_HI(net432));
 sg13g2_tiehi _7088__433 (.L_HI(net433));
 sg13g2_tiehi _6583__434 (.L_HI(net434));
 sg13g2_tiehi _7087__435 (.L_HI(net435));
 sg13g2_tiehi _6582__436 (.L_HI(net436));
 sg13g2_tiehi _7086__437 (.L_HI(net437));
 sg13g2_tiehi _6581__438 (.L_HI(net438));
 sg13g2_tiehi _7085__439 (.L_HI(net439));
 sg13g2_tiehi _6580__440 (.L_HI(net440));
 sg13g2_tiehi _7084__441 (.L_HI(net441));
 sg13g2_tiehi _6579__442 (.L_HI(net442));
 sg13g2_tiehi _7083__443 (.L_HI(net443));
 sg13g2_tiehi _6578__444 (.L_HI(net444));
 sg13g2_tiehi _7082__445 (.L_HI(net445));
 sg13g2_tiehi _6577__446 (.L_HI(net446));
 sg13g2_tiehi _7081__447 (.L_HI(net447));
 sg13g2_tiehi _6576__448 (.L_HI(net448));
 sg13g2_tiehi _7080__449 (.L_HI(net449));
 sg13g2_tiehi _6575__450 (.L_HI(net450));
 sg13g2_tiehi _6574__451 (.L_HI(net451));
 sg13g2_tiehi _6573__452 (.L_HI(net452));
 sg13g2_tiehi _6572__453 (.L_HI(net453));
 sg13g2_tiehi _7079__454 (.L_HI(net454));
 sg13g2_tiehi _6571__455 (.L_HI(net455));
 sg13g2_tiehi _7078__456 (.L_HI(net456));
 sg13g2_tiehi _6570__457 (.L_HI(net457));
 sg13g2_tiehi _7077__458 (.L_HI(net458));
 sg13g2_tiehi _6569__459 (.L_HI(net459));
 sg13g2_tiehi _7076__460 (.L_HI(net460));
 sg13g2_tiehi _6568__461 (.L_HI(net461));
 sg13g2_tiehi _7075__462 (.L_HI(net462));
 sg13g2_tiehi _6567__463 (.L_HI(net463));
 sg13g2_tiehi _7074__464 (.L_HI(net464));
 sg13g2_tiehi _6566__465 (.L_HI(net465));
 sg13g2_tiehi _7073__466 (.L_HI(net466));
 sg13g2_tiehi _6565__467 (.L_HI(net467));
 sg13g2_tiehi _7072__468 (.L_HI(net468));
 sg13g2_tiehi _6564__469 (.L_HI(net469));
 sg13g2_tiehi _7071__470 (.L_HI(net470));
 sg13g2_tiehi _6563__471 (.L_HI(net471));
 sg13g2_tiehi _7070__472 (.L_HI(net472));
 sg13g2_tiehi _6562__473 (.L_HI(net473));
 sg13g2_tiehi _7069__474 (.L_HI(net474));
 sg13g2_tiehi _6561__475 (.L_HI(net475));
 sg13g2_tiehi _7068__476 (.L_HI(net476));
 sg13g2_tiehi _6560__477 (.L_HI(net477));
 sg13g2_tiehi _7067__478 (.L_HI(net478));
 sg13g2_tiehi _6559__479 (.L_HI(net479));
 sg13g2_tiehi _7066__480 (.L_HI(net480));
 sg13g2_tiehi _6558__481 (.L_HI(net481));
 sg13g2_tiehi _7065__482 (.L_HI(net482));
 sg13g2_tiehi _6557__483 (.L_HI(net483));
 sg13g2_tiehi _7064__484 (.L_HI(net484));
 sg13g2_tiehi _6556__485 (.L_HI(net485));
 sg13g2_tiehi _6555__486 (.L_HI(net486));
 sg13g2_tiehi _6554__487 (.L_HI(net487));
 sg13g2_tiehi _6553__488 (.L_HI(net488));
 sg13g2_tiehi _6552__489 (.L_HI(net489));
 sg13g2_tiehi _6551__490 (.L_HI(net490));
 sg13g2_tiehi _6550__491 (.L_HI(net491));
 sg13g2_tiehi _6549__492 (.L_HI(net492));
 sg13g2_tiehi _6548__493 (.L_HI(net493));
 sg13g2_tiehi _7063__494 (.L_HI(net494));
 sg13g2_tiehi _6547__495 (.L_HI(net495));
 sg13g2_tiehi _7062__496 (.L_HI(net496));
 sg13g2_tiehi _6546__497 (.L_HI(net497));
 sg13g2_tiehi _7061__498 (.L_HI(net498));
 sg13g2_tiehi _6545__499 (.L_HI(net499));
 sg13g2_tiehi _7060__500 (.L_HI(net500));
 sg13g2_tiehi _6544__501 (.L_HI(net501));
 sg13g2_tiehi _7059__502 (.L_HI(net502));
 sg13g2_tiehi _6543__503 (.L_HI(net503));
 sg13g2_tiehi _7058__504 (.L_HI(net504));
 sg13g2_tiehi _6542__505 (.L_HI(net505));
 sg13g2_tiehi _7057__506 (.L_HI(net506));
 sg13g2_tiehi _6541__507 (.L_HI(net507));
 sg13g2_tiehi _7056__508 (.L_HI(net508));
 sg13g2_tiehi _6540__509 (.L_HI(net509));
 sg13g2_tiehi _7055__510 (.L_HI(net510));
 sg13g2_tiehi _6539__511 (.L_HI(net511));
 sg13g2_tiehi _7054__512 (.L_HI(net512));
 sg13g2_tiehi _6538__513 (.L_HI(net513));
 sg13g2_tiehi _7053__514 (.L_HI(net514));
 sg13g2_tiehi _6537__515 (.L_HI(net515));
 sg13g2_tiehi _7052__516 (.L_HI(net516));
 sg13g2_tiehi _6536__517 (.L_HI(net517));
 sg13g2_tiehi _6535__518 (.L_HI(net518));
 sg13g2_tiehi _6534__519 (.L_HI(net519));
 sg13g2_tiehi _6533__520 (.L_HI(net520));
 sg13g2_tiehi _6532__521 (.L_HI(net521));
 sg13g2_tiehi _6531__522 (.L_HI(net522));
 sg13g2_tiehi _6530__523 (.L_HI(net523));
 sg13g2_tiehi _6529__524 (.L_HI(net524));
 sg13g2_tiehi _6528__525 (.L_HI(net525));
 sg13g2_tiehi _6527__526 (.L_HI(net526));
 sg13g2_tiehi _6526__527 (.L_HI(net527));
 sg13g2_tiehi _6525__528 (.L_HI(net528));
 sg13g2_tiehi _6524__529 (.L_HI(net529));
 sg13g2_tiehi _6523__530 (.L_HI(net530));
 sg13g2_tiehi _6522__531 (.L_HI(net531));
 sg13g2_tiehi _6521__532 (.L_HI(net532));
 sg13g2_tiehi _6520__533 (.L_HI(net533));
 sg13g2_tiehi _6519__534 (.L_HI(net534));
 sg13g2_tiehi _6518__535 (.L_HI(net535));
 sg13g2_tiehi _6517__536 (.L_HI(net536));
 sg13g2_tiehi _6516__537 (.L_HI(net537));
 sg13g2_tiehi _6515__538 (.L_HI(net538));
 sg13g2_tiehi _6514__539 (.L_HI(net539));
 sg13g2_tiehi _6513__540 (.L_HI(net540));
 sg13g2_tiehi _6512__541 (.L_HI(net541));
 sg13g2_tiehi _6511__542 (.L_HI(net542));
 sg13g2_tiehi _6510__543 (.L_HI(net543));
 sg13g2_tiehi _6509__544 (.L_HI(net544));
 sg13g2_tiehi _7051__545 (.L_HI(net545));
 sg13g2_tiehi _6508__546 (.L_HI(net546));
 sg13g2_tiehi _7050__547 (.L_HI(net547));
 sg13g2_tiehi _6507__548 (.L_HI(net548));
 sg13g2_tiehi _7049__549 (.L_HI(net549));
 sg13g2_tiehi _7048__550 (.L_HI(net550));
 sg13g2_tiehi _7047__551 (.L_HI(net551));
 sg13g2_tiehi _7046__552 (.L_HI(net552));
 sg13g2_tiehi _7045__553 (.L_HI(net553));
 sg13g2_tiehi _7044__554 (.L_HI(net554));
 sg13g2_tiehi _7043__555 (.L_HI(net555));
 sg13g2_tiehi _7042__556 (.L_HI(net556));
 sg13g2_tiehi _7041__557 (.L_HI(net557));
 sg13g2_tiehi _7040__558 (.L_HI(net558));
 sg13g2_tiehi _7039__559 (.L_HI(net559));
 sg13g2_tiehi _7038__560 (.L_HI(net560));
 sg13g2_tiehi _7037__561 (.L_HI(net561));
 sg13g2_tiehi _7036__562 (.L_HI(net562));
 sg13g2_tiehi _7035__563 (.L_HI(net563));
 sg13g2_tiehi _7034__564 (.L_HI(net564));
 sg13g2_tiehi _7033__565 (.L_HI(net565));
 sg13g2_tiehi _7032__566 (.L_HI(net566));
 sg13g2_tiehi _7031__567 (.L_HI(net567));
 sg13g2_tiehi _7030__568 (.L_HI(net568));
 sg13g2_tiehi _7029__569 (.L_HI(net569));
 sg13g2_tiehi _7028__570 (.L_HI(net570));
 sg13g2_tiehi _7027__571 (.L_HI(net571));
 sg13g2_tiehi _7026__572 (.L_HI(net572));
 sg13g2_tiehi _7025__573 (.L_HI(net573));
 sg13g2_tiehi _7024__574 (.L_HI(net574));
 sg13g2_tiehi _7023__575 (.L_HI(net575));
 sg13g2_tiehi _7022__576 (.L_HI(net576));
 sg13g2_tiehi _7021__577 (.L_HI(net577));
 sg13g2_tiehi _7020__578 (.L_HI(net578));
 sg13g2_tiehi _7019__579 (.L_HI(net579));
 sg13g2_tiehi _7018__580 (.L_HI(net580));
 sg13g2_tiehi _7017__581 (.L_HI(net581));
 sg13g2_tiehi _7016__582 (.L_HI(net582));
 sg13g2_tiehi _7015__583 (.L_HI(net583));
 sg13g2_tiehi _7014__584 (.L_HI(net584));
 sg13g2_tiehi _7013__585 (.L_HI(net585));
 sg13g2_tiehi _7012__586 (.L_HI(net586));
 sg13g2_tiehi _7011__587 (.L_HI(net587));
 sg13g2_tiehi _7010__588 (.L_HI(net588));
 sg13g2_tiehi _7009__589 (.L_HI(net589));
 sg13g2_tiehi _7008__590 (.L_HI(net590));
 sg13g2_tiehi _7007__591 (.L_HI(net591));
 sg13g2_tiehi _7006__592 (.L_HI(net592));
 sg13g2_tiehi _7005__593 (.L_HI(net593));
 sg13g2_tiehi _7004__594 (.L_HI(net594));
 sg13g2_tiehi _7003__595 (.L_HI(net595));
 sg13g2_tiehi _7002__596 (.L_HI(net596));
 sg13g2_tiehi _7001__597 (.L_HI(net597));
 sg13g2_tiehi _7000__598 (.L_HI(net598));
 sg13g2_tiehi _6999__599 (.L_HI(net599));
 sg13g2_tiehi _6998__600 (.L_HI(net600));
 sg13g2_tiehi _6997__601 (.L_HI(net601));
 sg13g2_tiehi _6996__602 (.L_HI(net602));
 sg13g2_tiehi _6995__603 (.L_HI(net603));
 sg13g2_tiehi _6994__604 (.L_HI(net604));
 sg13g2_tiehi _6993__605 (.L_HI(net605));
 sg13g2_tiehi _6992__606 (.L_HI(net606));
 sg13g2_tiehi _6991__607 (.L_HI(net607));
 sg13g2_tiehi _6990__608 (.L_HI(net608));
 sg13g2_tiehi _6989__609 (.L_HI(net609));
 sg13g2_tiehi _6988__610 (.L_HI(net610));
 sg13g2_tiehi _6987__611 (.L_HI(net611));
 sg13g2_tiehi _6986__612 (.L_HI(net612));
 sg13g2_tiehi _6985__613 (.L_HI(net613));
 sg13g2_tiehi _6984__614 (.L_HI(net614));
 sg13g2_tiehi _6983__615 (.L_HI(net615));
 sg13g2_tiehi _6982__616 (.L_HI(net616));
 sg13g2_tiehi _6981__617 (.L_HI(net617));
 sg13g2_tiehi _6980__618 (.L_HI(net618));
 sg13g2_tiehi _6979__619 (.L_HI(net619));
 sg13g2_tiehi _6978__620 (.L_HI(net620));
 sg13g2_tiehi _6977__621 (.L_HI(net621));
 sg13g2_tiehi _6976__622 (.L_HI(net622));
 sg13g2_tiehi _6975__623 (.L_HI(net623));
 sg13g2_tiehi _6974__624 (.L_HI(net624));
 sg13g2_tiehi _6973__625 (.L_HI(net625));
 sg13g2_tiehi _6972__626 (.L_HI(net626));
 sg13g2_tiehi _6971__627 (.L_HI(net627));
 sg13g2_tiehi _6970__628 (.L_HI(net628));
 sg13g2_tiehi _6969__629 (.L_HI(net629));
 sg13g2_tiehi _6968__630 (.L_HI(net630));
 sg13g2_tiehi _6967__631 (.L_HI(net631));
 sg13g2_tiehi _6966__632 (.L_HI(net632));
 sg13g2_tiehi _6965__633 (.L_HI(net633));
 sg13g2_tiehi _6964__634 (.L_HI(net634));
 sg13g2_tiehi _6963__635 (.L_HI(net635));
 sg13g2_tiehi _6962__636 (.L_HI(net636));
 sg13g2_tiehi _6961__637 (.L_HI(net637));
 sg13g2_tiehi _6960__638 (.L_HI(net638));
 sg13g2_tiehi _6959__639 (.L_HI(net639));
 sg13g2_tiehi _6958__640 (.L_HI(net640));
 sg13g2_tiehi _6957__641 (.L_HI(net641));
 sg13g2_tiehi _6956__642 (.L_HI(net642));
 sg13g2_tiehi _6955__643 (.L_HI(net643));
 sg13g2_tiehi _6954__644 (.L_HI(net644));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_vga_tetris_6 (.L_LO(net6));
 sg13g2_tielo tt_um_vga_tetris_7 (.L_LO(net7));
 sg13g2_tielo tt_um_vga_tetris_8 (.L_LO(net8));
 sg13g2_tielo tt_um_vga_tetris_9 (.L_LO(net9));
 sg13g2_tielo tt_um_vga_tetris_10 (.L_LO(net10));
 sg13g2_tielo tt_um_vga_tetris_11 (.L_LO(net11));
 sg13g2_tielo tt_um_vga_tetris_12 (.L_LO(net12));
 sg13g2_tielo tt_um_vga_tetris_13 (.L_LO(net13));
 sg13g2_tielo tt_um_vga_tetris_14 (.L_LO(net14));
 sg13g2_tielo tt_um_vga_tetris_15 (.L_LO(net15));
 sg13g2_tielo tt_um_vga_tetris_16 (.L_LO(net16));
 sg13g2_tielo tt_um_vga_tetris_17 (.L_LO(net17));
 sg13g2_tielo tt_um_vga_tetris_18 (.L_LO(net18));
 sg13g2_tielo tt_um_vga_tetris_19 (.L_LO(net19));
 sg13g2_tielo tt_um_vga_tetris_20 (.L_LO(net20));
 sg13g2_tiehi _6953__21 (.L_HI(net21));
 sg13g2_buf_1 _7770_ (.A(\vga_tetris._vgaController_io_vSync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _7771_ (.A(vga_hs),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout837 (.A(_1658_),
    .X(net837));
 sg13g2_buf_8 fanout838 (.A(_2134_),
    .X(net838));
 sg13g2_buf_8 fanout839 (.A(net841),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(net841),
    .X(net840));
 sg13g2_buf_8 fanout841 (.A(net845),
    .X(net841));
 sg13g2_buf_8 fanout842 (.A(net845),
    .X(net842));
 sg13g2_buf_8 fanout843 (.A(net844),
    .X(net843));
 sg13g2_buf_8 fanout844 (.A(net845),
    .X(net844));
 sg13g2_buf_8 fanout845 (.A(_2838_),
    .X(net845));
 sg13g2_buf_8 fanout846 (.A(net848),
    .X(net846));
 sg13g2_buf_8 fanout847 (.A(net848),
    .X(net847));
 sg13g2_buf_8 fanout848 (.A(_2817_),
    .X(net848));
 sg13g2_buf_8 fanout849 (.A(net851),
    .X(net849));
 sg13g2_buf_8 fanout850 (.A(net851),
    .X(net850));
 sg13g2_buf_8 fanout851 (.A(_2817_),
    .X(net851));
 sg13g2_buf_8 fanout852 (.A(net854),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(net854),
    .X(net853));
 sg13g2_buf_8 fanout854 (.A(_2796_),
    .X(net854));
 sg13g2_buf_8 fanout855 (.A(net857),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(net857),
    .X(net856));
 sg13g2_buf_8 fanout857 (.A(_2796_),
    .X(net857));
 sg13g2_buf_8 fanout858 (.A(net860),
    .X(net858));
 sg13g2_buf_8 fanout859 (.A(net860),
    .X(net859));
 sg13g2_buf_8 fanout860 (.A(_2775_),
    .X(net860));
 sg13g2_buf_8 fanout861 (.A(net862),
    .X(net861));
 sg13g2_buf_8 fanout862 (.A(_2775_),
    .X(net862));
 sg13g2_buf_8 fanout863 (.A(_2775_),
    .X(net863));
 sg13g2_buf_8 fanout864 (.A(net866),
    .X(net864));
 sg13g2_buf_8 fanout865 (.A(net866),
    .X(net865));
 sg13g2_buf_8 fanout866 (.A(_2754_),
    .X(net866));
 sg13g2_buf_8 fanout867 (.A(net869),
    .X(net867));
 sg13g2_buf_8 fanout868 (.A(net869),
    .X(net868));
 sg13g2_buf_8 fanout869 (.A(_2754_),
    .X(net869));
 sg13g2_buf_8 fanout870 (.A(net871),
    .X(net870));
 sg13g2_buf_8 fanout871 (.A(net875),
    .X(net871));
 sg13g2_buf_8 fanout872 (.A(net873),
    .X(net872));
 sg13g2_buf_8 fanout873 (.A(net875),
    .X(net873));
 sg13g2_buf_8 fanout874 (.A(net875),
    .X(net874));
 sg13g2_buf_8 fanout875 (.A(_2733_),
    .X(net875));
 sg13g2_buf_8 fanout876 (.A(net878),
    .X(net876));
 sg13g2_buf_1 fanout877 (.A(net878),
    .X(net877));
 sg13g2_buf_8 fanout878 (.A(_2712_),
    .X(net878));
 sg13g2_buf_8 fanout879 (.A(net880),
    .X(net879));
 sg13g2_buf_8 fanout880 (.A(net881),
    .X(net880));
 sg13g2_buf_8 fanout881 (.A(_2712_),
    .X(net881));
 sg13g2_buf_8 fanout882 (.A(net884),
    .X(net882));
 sg13g2_buf_8 fanout883 (.A(net884),
    .X(net883));
 sg13g2_buf_8 fanout884 (.A(_2690_),
    .X(net884));
 sg13g2_buf_8 fanout885 (.A(net887),
    .X(net885));
 sg13g2_buf_8 fanout886 (.A(net887),
    .X(net886));
 sg13g2_buf_8 fanout887 (.A(_2690_),
    .X(net887));
 sg13g2_buf_8 fanout888 (.A(net890),
    .X(net888));
 sg13g2_buf_1 fanout889 (.A(net890),
    .X(net889));
 sg13g2_buf_8 fanout890 (.A(net894),
    .X(net890));
 sg13g2_buf_8 fanout891 (.A(net894),
    .X(net891));
 sg13g2_buf_1 fanout892 (.A(net894),
    .X(net892));
 sg13g2_buf_8 fanout893 (.A(net894),
    .X(net893));
 sg13g2_buf_8 fanout894 (.A(_2669_),
    .X(net894));
 sg13g2_buf_8 fanout895 (.A(net897),
    .X(net895));
 sg13g2_buf_8 fanout896 (.A(net897),
    .X(net896));
 sg13g2_buf_8 fanout897 (.A(_2648_),
    .X(net897));
 sg13g2_buf_8 fanout898 (.A(net899),
    .X(net898));
 sg13g2_buf_8 fanout899 (.A(net900),
    .X(net899));
 sg13g2_buf_8 fanout900 (.A(_2648_),
    .X(net900));
 sg13g2_buf_8 fanout901 (.A(net902),
    .X(net901));
 sg13g2_buf_8 fanout902 (.A(net906),
    .X(net902));
 sg13g2_buf_8 fanout903 (.A(net906),
    .X(net903));
 sg13g2_buf_8 fanout904 (.A(net906),
    .X(net904));
 sg13g2_buf_8 fanout905 (.A(net906),
    .X(net905));
 sg13g2_buf_8 fanout906 (.A(_2627_),
    .X(net906));
 sg13g2_buf_8 fanout907 (.A(net909),
    .X(net907));
 sg13g2_buf_8 fanout908 (.A(net909),
    .X(net908));
 sg13g2_buf_8 fanout909 (.A(_2605_),
    .X(net909));
 sg13g2_buf_8 fanout910 (.A(net912),
    .X(net910));
 sg13g2_buf_8 fanout911 (.A(net912),
    .X(net911));
 sg13g2_buf_8 fanout912 (.A(_2605_),
    .X(net912));
 sg13g2_buf_8 fanout913 (.A(net915),
    .X(net913));
 sg13g2_buf_8 fanout914 (.A(net915),
    .X(net914));
 sg13g2_buf_8 fanout915 (.A(_2584_),
    .X(net915));
 sg13g2_buf_8 fanout916 (.A(net917),
    .X(net916));
 sg13g2_buf_8 fanout917 (.A(net918),
    .X(net917));
 sg13g2_buf_8 fanout918 (.A(_2584_),
    .X(net918));
 sg13g2_buf_8 fanout919 (.A(net921),
    .X(net919));
 sg13g2_buf_8 fanout920 (.A(net921),
    .X(net920));
 sg13g2_buf_8 fanout921 (.A(_2563_),
    .X(net921));
 sg13g2_buf_8 fanout922 (.A(net924),
    .X(net922));
 sg13g2_buf_8 fanout923 (.A(net924),
    .X(net923));
 sg13g2_buf_8 fanout924 (.A(_2563_),
    .X(net924));
 sg13g2_buf_8 fanout925 (.A(net928),
    .X(net925));
 sg13g2_buf_1 fanout926 (.A(net928),
    .X(net926));
 sg13g2_buf_8 fanout927 (.A(net928),
    .X(net927));
 sg13g2_buf_8 fanout928 (.A(net931),
    .X(net928));
 sg13g2_buf_8 fanout929 (.A(net930),
    .X(net929));
 sg13g2_buf_8 fanout930 (.A(net931),
    .X(net930));
 sg13g2_buf_8 fanout931 (.A(_2542_),
    .X(net931));
 sg13g2_buf_8 fanout932 (.A(net934),
    .X(net932));
 sg13g2_buf_2 fanout933 (.A(net934),
    .X(net933));
 sg13g2_buf_8 fanout934 (.A(_2520_),
    .X(net934));
 sg13g2_buf_8 fanout935 (.A(net936),
    .X(net935));
 sg13g2_buf_8 fanout936 (.A(net937),
    .X(net936));
 sg13g2_buf_8 fanout937 (.A(_2520_),
    .X(net937));
 sg13g2_buf_8 fanout938 (.A(net939),
    .X(net938));
 sg13g2_buf_8 fanout939 (.A(net940),
    .X(net939));
 sg13g2_buf_8 fanout940 (.A(_2498_),
    .X(net940));
 sg13g2_buf_8 fanout941 (.A(_2498_),
    .X(net941));
 sg13g2_buf_2 fanout942 (.A(net943),
    .X(net942));
 sg13g2_buf_8 fanout943 (.A(_2498_),
    .X(net943));
 sg13g2_buf_8 fanout944 (.A(net946),
    .X(net944));
 sg13g2_buf_8 fanout945 (.A(net946),
    .X(net945));
 sg13g2_buf_8 fanout946 (.A(net950),
    .X(net946));
 sg13g2_buf_8 fanout947 (.A(net950),
    .X(net947));
 sg13g2_buf_2 fanout948 (.A(net950),
    .X(net948));
 sg13g2_buf_8 fanout949 (.A(net950),
    .X(net949));
 sg13g2_buf_8 fanout950 (.A(_2476_),
    .X(net950));
 sg13g2_buf_8 fanout951 (.A(net953),
    .X(net951));
 sg13g2_buf_1 fanout952 (.A(net953),
    .X(net952));
 sg13g2_buf_8 fanout953 (.A(net957),
    .X(net953));
 sg13g2_buf_8 fanout954 (.A(net955),
    .X(net954));
 sg13g2_buf_8 fanout955 (.A(net957),
    .X(net955));
 sg13g2_buf_8 fanout956 (.A(net957),
    .X(net956));
 sg13g2_buf_8 fanout957 (.A(_2453_),
    .X(net957));
 sg13g2_buf_8 fanout958 (.A(net960),
    .X(net958));
 sg13g2_buf_8 fanout959 (.A(net960),
    .X(net959));
 sg13g2_buf_8 fanout960 (.A(_2254_),
    .X(net960));
 sg13g2_buf_8 fanout961 (.A(net963),
    .X(net961));
 sg13g2_buf_1 fanout962 (.A(net963),
    .X(net962));
 sg13g2_buf_8 fanout963 (.A(_2254_),
    .X(net963));
 sg13g2_buf_8 fanout964 (.A(net966),
    .X(net964));
 sg13g2_buf_8 fanout965 (.A(net966),
    .X(net965));
 sg13g2_buf_8 fanout966 (.A(_0833_),
    .X(net966));
 sg13g2_buf_8 fanout967 (.A(_0832_),
    .X(net967));
 sg13g2_buf_8 fanout968 (.A(_0832_),
    .X(net968));
 sg13g2_buf_8 fanout969 (.A(_0857_),
    .X(net969));
 sg13g2_buf_8 fanout970 (.A(_0857_),
    .X(net970));
 sg13g2_buf_8 fanout971 (.A(_0856_),
    .X(net971));
 sg13g2_buf_8 fanout972 (.A(_0854_),
    .X(net972));
 sg13g2_buf_8 fanout973 (.A(_0854_),
    .X(net973));
 sg13g2_buf_8 fanout974 (.A(_0853_),
    .X(net974));
 sg13g2_buf_8 fanout975 (.A(_0853_),
    .X(net975));
 sg13g2_buf_8 fanout976 (.A(net977),
    .X(net976));
 sg13g2_buf_8 fanout977 (.A(_0851_),
    .X(net977));
 sg13g2_buf_8 fanout978 (.A(_0850_),
    .X(net978));
 sg13g2_buf_8 fanout979 (.A(net980),
    .X(net979));
 sg13g2_buf_8 fanout980 (.A(_0846_),
    .X(net980));
 sg13g2_buf_8 fanout981 (.A(_0845_),
    .X(net981));
 sg13g2_buf_8 fanout982 (.A(_0845_),
    .X(net982));
 sg13g2_buf_8 fanout983 (.A(_0843_),
    .X(net983));
 sg13g2_buf_8 fanout984 (.A(_0843_),
    .X(net984));
 sg13g2_buf_8 fanout985 (.A(_0842_),
    .X(net985));
 sg13g2_buf_8 fanout986 (.A(_0842_),
    .X(net986));
 sg13g2_buf_8 fanout987 (.A(_0841_),
    .X(net987));
 sg13g2_buf_8 fanout988 (.A(_0841_),
    .X(net988));
 sg13g2_buf_8 fanout989 (.A(net990),
    .X(net989));
 sg13g2_buf_8 fanout990 (.A(_0839_),
    .X(net990));
 sg13g2_buf_8 fanout991 (.A(_0837_),
    .X(net991));
 sg13g2_buf_8 fanout992 (.A(_0834_),
    .X(net992));
 sg13g2_buf_8 fanout993 (.A(net994),
    .X(net993));
 sg13g2_buf_8 fanout994 (.A(_0831_),
    .X(net994));
 sg13g2_buf_8 fanout995 (.A(net996),
    .X(net995));
 sg13g2_buf_8 fanout996 (.A(_0829_),
    .X(net996));
 sg13g2_buf_8 fanout997 (.A(_0827_),
    .X(net997));
 sg13g2_buf_8 fanout998 (.A(_0827_),
    .X(net998));
 sg13g2_buf_8 fanout999 (.A(_0825_),
    .X(net999));
 sg13g2_buf_8 fanout1000 (.A(_0825_),
    .X(net1000));
 sg13g2_buf_8 fanout1001 (.A(_0821_),
    .X(net1001));
 sg13g2_buf_8 fanout1002 (.A(net1003),
    .X(net1002));
 sg13g2_buf_8 fanout1003 (.A(_0818_),
    .X(net1003));
 sg13g2_buf_8 fanout1004 (.A(net1005),
    .X(net1004));
 sg13g2_buf_8 fanout1005 (.A(_0844_),
    .X(net1005));
 sg13g2_buf_8 fanout1006 (.A(net1007),
    .X(net1006));
 sg13g2_buf_8 fanout1007 (.A(_0844_),
    .X(net1007));
 sg13g2_buf_8 fanout1008 (.A(net1012),
    .X(net1008));
 sg13g2_buf_1 fanout1009 (.A(net1012),
    .X(net1009));
 sg13g2_buf_8 fanout1010 (.A(net1011),
    .X(net1010));
 sg13g2_buf_2 fanout1011 (.A(net1012),
    .X(net1011));
 sg13g2_buf_8 fanout1012 (.A(net1016),
    .X(net1012));
 sg13g2_buf_8 fanout1013 (.A(net1014),
    .X(net1013));
 sg13g2_buf_8 fanout1014 (.A(net1016),
    .X(net1014));
 sg13g2_buf_8 fanout1015 (.A(net1016),
    .X(net1015));
 sg13g2_buf_8 fanout1016 (.A(_0836_),
    .X(net1016));
 sg13g2_buf_8 fanout1017 (.A(net1022),
    .X(net1017));
 sg13g2_buf_8 fanout1018 (.A(net1019),
    .X(net1018));
 sg13g2_buf_8 fanout1019 (.A(net1022),
    .X(net1019));
 sg13g2_buf_8 fanout1020 (.A(net1021),
    .X(net1020));
 sg13g2_buf_8 fanout1021 (.A(net1022),
    .X(net1021));
 sg13g2_buf_8 fanout1022 (.A(_0830_),
    .X(net1022));
 sg13g2_buf_8 fanout1023 (.A(net1025),
    .X(net1023));
 sg13g2_buf_8 fanout1024 (.A(net1025),
    .X(net1024));
 sg13g2_buf_8 fanout1025 (.A(_0828_),
    .X(net1025));
 sg13g2_buf_8 fanout1026 (.A(_0828_),
    .X(net1026));
 sg13g2_buf_2 fanout1027 (.A(_0828_),
    .X(net1027));
 sg13g2_buf_8 fanout1028 (.A(net1031),
    .X(net1028));
 sg13g2_buf_8 fanout1029 (.A(net1030),
    .X(net1029));
 sg13g2_buf_8 fanout1030 (.A(net1031),
    .X(net1030));
 sg13g2_buf_8 fanout1031 (.A(_0824_),
    .X(net1031));
 sg13g2_buf_8 fanout1032 (.A(net1034),
    .X(net1032));
 sg13g2_buf_1 fanout1033 (.A(net1034),
    .X(net1033));
 sg13g2_buf_8 fanout1034 (.A(_0824_),
    .X(net1034));
 sg13g2_buf_8 fanout1035 (.A(net1036),
    .X(net1035));
 sg13g2_buf_8 fanout1036 (.A(_0823_),
    .X(net1036));
 sg13g2_buf_8 fanout1037 (.A(_0823_),
    .X(net1037));
 sg13g2_buf_8 fanout1038 (.A(net1039),
    .X(net1038));
 sg13g2_buf_8 fanout1039 (.A(net1040),
    .X(net1039));
 sg13g2_buf_8 fanout1040 (.A(_0823_),
    .X(net1040));
 sg13g2_buf_8 fanout1041 (.A(net1043),
    .X(net1041));
 sg13g2_buf_8 fanout1042 (.A(net1043),
    .X(net1042));
 sg13g2_buf_8 fanout1043 (.A(_0820_),
    .X(net1043));
 sg13g2_buf_8 fanout1044 (.A(net1045),
    .X(net1044));
 sg13g2_buf_8 fanout1045 (.A(_0820_),
    .X(net1045));
 sg13g2_buf_8 fanout1046 (.A(net1051),
    .X(net1046));
 sg13g2_buf_2 fanout1047 (.A(net1051),
    .X(net1047));
 sg13g2_buf_8 fanout1048 (.A(net1049),
    .X(net1048));
 sg13g2_buf_8 fanout1049 (.A(net1051),
    .X(net1049));
 sg13g2_buf_8 fanout1050 (.A(net1051),
    .X(net1050));
 sg13g2_buf_8 fanout1051 (.A(_0817_),
    .X(net1051));
 sg13g2_buf_8 fanout1052 (.A(net1055),
    .X(net1052));
 sg13g2_buf_1 fanout1053 (.A(net1055),
    .X(net1053));
 sg13g2_buf_8 fanout1054 (.A(net1055),
    .X(net1054));
 sg13g2_buf_8 fanout1055 (.A(_0789_),
    .X(net1055));
 sg13g2_buf_8 fanout1056 (.A(net1058),
    .X(net1056));
 sg13g2_buf_1 fanout1057 (.A(net1058),
    .X(net1057));
 sg13g2_buf_8 fanout1058 (.A(_0789_),
    .X(net1058));
 sg13g2_buf_8 fanout1059 (.A(net1060),
    .X(net1059));
 sg13g2_buf_2 fanout1060 (.A(_1610_),
    .X(net1060));
 sg13g2_buf_8 fanout1061 (.A(_2912_),
    .X(net1061));
 sg13g2_buf_8 fanout1062 (.A(_1623_),
    .X(net1062));
 sg13g2_buf_8 fanout1063 (.A(_1762_),
    .X(net1063));
 sg13g2_buf_8 fanout1064 (.A(_1539_),
    .X(net1064));
 sg13g2_buf_8 fanout1065 (.A(_0892_),
    .X(net1065));
 sg13g2_buf_8 fanout1066 (.A(_0892_),
    .X(net1066));
 sg13g2_buf_8 fanout1067 (.A(_1759_),
    .X(net1067));
 sg13g2_buf_8 fanout1068 (.A(_0891_),
    .X(net1068));
 sg13g2_buf_8 fanout1069 (.A(_1576_),
    .X(net1069));
 sg13g2_buf_8 fanout1070 (.A(_2409_),
    .X(net1070));
 sg13g2_buf_8 fanout1071 (.A(net1073),
    .X(net1071));
 sg13g2_buf_8 fanout1072 (.A(net1073),
    .X(net1072));
 sg13g2_buf_8 fanout1073 (.A(_2334_),
    .X(net1073));
 sg13g2_buf_8 fanout1074 (.A(net1075),
    .X(net1074));
 sg13g2_buf_8 fanout1075 (.A(net1076),
    .X(net1075));
 sg13g2_buf_8 fanout1076 (.A(_2330_),
    .X(net1076));
 sg13g2_buf_8 fanout1077 (.A(net1079),
    .X(net1077));
 sg13g2_buf_8 fanout1078 (.A(net1079),
    .X(net1078));
 sg13g2_buf_8 fanout1079 (.A(_2326_),
    .X(net1079));
 sg13g2_buf_8 fanout1080 (.A(net1082),
    .X(net1080));
 sg13g2_buf_8 fanout1081 (.A(net1082),
    .X(net1081));
 sg13g2_buf_8 fanout1082 (.A(_2322_),
    .X(net1082));
 sg13g2_buf_8 fanout1083 (.A(net1085),
    .X(net1083));
 sg13g2_buf_2 fanout1084 (.A(net1085),
    .X(net1084));
 sg13g2_buf_8 fanout1085 (.A(net1903),
    .X(net1085));
 sg13g2_buf_8 fanout1086 (.A(net1088),
    .X(net1086));
 sg13g2_buf_8 fanout1087 (.A(net1088),
    .X(net1087));
 sg13g2_buf_8 fanout1088 (.A(_2314_),
    .X(net1088));
 sg13g2_buf_8 fanout1089 (.A(net1091),
    .X(net1089));
 sg13g2_buf_8 fanout1090 (.A(net1091),
    .X(net1090));
 sg13g2_buf_8 fanout1091 (.A(_2310_),
    .X(net1091));
 sg13g2_buf_8 fanout1092 (.A(net1094),
    .X(net1092));
 sg13g2_buf_1 fanout1093 (.A(net1094),
    .X(net1093));
 sg13g2_buf_1 fanout1094 (.A(net1095),
    .X(net1094));
 sg13g2_buf_8 fanout1095 (.A(_2306_),
    .X(net1095));
 sg13g2_buf_8 fanout1096 (.A(net1098),
    .X(net1096));
 sg13g2_buf_2 fanout1097 (.A(net1098),
    .X(net1097));
 sg13g2_buf_8 fanout1098 (.A(_2302_),
    .X(net1098));
 sg13g2_buf_8 fanout1099 (.A(net1100),
    .X(net1099));
 sg13g2_buf_8 fanout1100 (.A(net1101),
    .X(net1100));
 sg13g2_buf_8 fanout1101 (.A(_2298_),
    .X(net1101));
 sg13g2_buf_8 fanout1102 (.A(net1104),
    .X(net1102));
 sg13g2_buf_1 fanout1103 (.A(net1104),
    .X(net1103));
 sg13g2_buf_8 fanout1104 (.A(_2294_),
    .X(net1104));
 sg13g2_buf_8 fanout1105 (.A(net1106),
    .X(net1105));
 sg13g2_buf_8 fanout1106 (.A(net1107),
    .X(net1106));
 sg13g2_buf_8 fanout1107 (.A(_2290_),
    .X(net1107));
 sg13g2_buf_8 fanout1108 (.A(net1110),
    .X(net1108));
 sg13g2_buf_1 fanout1109 (.A(net1110),
    .X(net1109));
 sg13g2_buf_8 fanout1110 (.A(_2286_),
    .X(net1110));
 sg13g2_buf_8 fanout1111 (.A(_2282_),
    .X(net1111));
 sg13g2_buf_8 fanout1112 (.A(net1113),
    .X(net1112));
 sg13g2_buf_1 fanout1113 (.A(_2282_),
    .X(net1113));
 sg13g2_buf_8 fanout1114 (.A(net1116),
    .X(net1114));
 sg13g2_buf_1 fanout1115 (.A(net1116),
    .X(net1115));
 sg13g2_buf_8 fanout1116 (.A(_2278_),
    .X(net1116));
 sg13g2_buf_8 fanout1117 (.A(net1119),
    .X(net1117));
 sg13g2_buf_2 fanout1118 (.A(net1119),
    .X(net1118));
 sg13g2_buf_8 fanout1119 (.A(_2274_),
    .X(net1119));
 sg13g2_buf_8 fanout1120 (.A(net1122),
    .X(net1120));
 sg13g2_buf_8 fanout1121 (.A(net1122),
    .X(net1121));
 sg13g2_buf_8 fanout1122 (.A(_2270_),
    .X(net1122));
 sg13g2_buf_8 fanout1123 (.A(net1125),
    .X(net1123));
 sg13g2_buf_8 fanout1124 (.A(_2266_),
    .X(net1124));
 sg13g2_buf_2 fanout1125 (.A(_2266_),
    .X(net1125));
 sg13g2_buf_8 fanout1126 (.A(net1128),
    .X(net1126));
 sg13g2_buf_1 fanout1127 (.A(net1128),
    .X(net1127));
 sg13g2_buf_8 fanout1128 (.A(net1129),
    .X(net1128));
 sg13g2_buf_8 fanout1129 (.A(_2262_),
    .X(net1129));
 sg13g2_buf_8 fanout1130 (.A(net1132),
    .X(net1130));
 sg13g2_buf_8 fanout1131 (.A(net1132),
    .X(net1131));
 sg13g2_buf_8 fanout1132 (.A(_2258_),
    .X(net1132));
 sg13g2_buf_8 fanout1133 (.A(_2206_),
    .X(net1133));
 sg13g2_buf_1 fanout1134 (.A(_2206_),
    .X(net1134));
 sg13g2_buf_8 fanout1135 (.A(_1782_),
    .X(net1135));
 sg13g2_buf_8 fanout1136 (.A(_2056_),
    .X(net1136));
 sg13g2_buf_8 fanout1137 (.A(_2053_),
    .X(net1137));
 sg13g2_buf_8 fanout1138 (.A(_1705_),
    .X(net1138));
 sg13g2_buf_8 fanout1139 (.A(net1140),
    .X(net1139));
 sg13g2_buf_8 fanout1140 (.A(net1142),
    .X(net1140));
 sg13g2_buf_8 fanout1141 (.A(net1142),
    .X(net1141));
 sg13g2_buf_8 fanout1142 (.A(_1507_),
    .X(net1142));
 sg13g2_buf_8 fanout1143 (.A(net1144),
    .X(net1143));
 sg13g2_buf_8 fanout1144 (.A(net1145),
    .X(net1144));
 sg13g2_buf_1 fanout1145 (.A(net1149),
    .X(net1145));
 sg13g2_buf_8 fanout1146 (.A(net1148),
    .X(net1146));
 sg13g2_buf_1 fanout1147 (.A(net1148),
    .X(net1147));
 sg13g2_buf_8 fanout1148 (.A(net1149),
    .X(net1148));
 sg13g2_buf_8 fanout1149 (.A(_0736_),
    .X(net1149));
 sg13g2_buf_8 fanout1150 (.A(_0710_),
    .X(net1150));
 sg13g2_buf_8 fanout1151 (.A(net1152),
    .X(net1151));
 sg13g2_buf_8 fanout1152 (.A(net1153),
    .X(net1152));
 sg13g2_buf_8 fanout1153 (.A(net1155),
    .X(net1153));
 sg13g2_buf_8 fanout1154 (.A(net1155),
    .X(net1154));
 sg13g2_buf_8 fanout1155 (.A(_2170_),
    .X(net1155));
 sg13g2_buf_8 fanout1156 (.A(net1157),
    .X(net1156));
 sg13g2_buf_8 fanout1157 (.A(net1160),
    .X(net1157));
 sg13g2_buf_8 fanout1158 (.A(net1159),
    .X(net1158));
 sg13g2_buf_8 fanout1159 (.A(net1160),
    .X(net1159));
 sg13g2_buf_8 fanout1160 (.A(_1669_),
    .X(net1160));
 sg13g2_buf_2 fanout1161 (.A(net1163),
    .X(net1161));
 sg13g2_buf_1 fanout1162 (.A(net1163),
    .X(net1162));
 sg13g2_buf_8 fanout1163 (.A(net1164),
    .X(net1163));
 sg13g2_buf_8 fanout1164 (.A(_0887_),
    .X(net1164));
 sg13g2_buf_8 fanout1165 (.A(net1166),
    .X(net1165));
 sg13g2_buf_8 fanout1166 (.A(net1167),
    .X(net1166));
 sg13g2_buf_2 fanout1167 (.A(_0887_),
    .X(net1167));
 sg13g2_buf_8 fanout1168 (.A(net1169),
    .X(net1168));
 sg13g2_buf_8 fanout1169 (.A(_0702_),
    .X(net1169));
 sg13g2_buf_8 fanout1170 (.A(net1171),
    .X(net1170));
 sg13g2_buf_2 fanout1171 (.A(net1172),
    .X(net1171));
 sg13g2_buf_8 fanout1172 (.A(net1173),
    .X(net1172));
 sg13g2_buf_8 fanout1173 (.A(_0699_),
    .X(net1173));
 sg13g2_buf_8 fanout1174 (.A(_0698_),
    .X(net1174));
 sg13g2_buf_8 fanout1175 (.A(_0662_),
    .X(net1175));
 sg13g2_buf_8 fanout1176 (.A(_0659_),
    .X(net1176));
 sg13g2_buf_8 fanout1177 (.A(net1771),
    .X(net1177));
 sg13g2_buf_1 fanout1178 (.A(\vga_tetris.runningTetrisLogicQ ),
    .X(net1178));
 sg13g2_buf_8 fanout1179 (.A(net1793),
    .X(net1179));
 sg13g2_buf_8 fanout1180 (.A(net1181),
    .X(net1180));
 sg13g2_buf_8 fanout1181 (.A(net1889),
    .X(net1181));
 sg13g2_buf_8 fanout1182 (.A(net1184),
    .X(net1182));
 sg13g2_buf_1 fanout1183 (.A(net1184),
    .X(net1183));
 sg13g2_buf_8 fanout1184 (.A(\vga_tetris._tetrisDisplay_io_boardYCoord[0] ),
    .X(net1184));
 sg13g2_buf_8 fanout1185 (.A(net1186),
    .X(net1185));
 sg13g2_buf_1 fanout1186 (.A(net1187),
    .X(net1186));
 sg13g2_buf_2 fanout1187 (.A(net1856),
    .X(net1187));
 sg13g2_buf_8 fanout1188 (.A(net1861),
    .X(net1188));
 sg13g2_buf_1 fanout1189 (.A(\vga_tetris._vgaController_io_pixelPosY[2] ),
    .X(net1189));
 sg13g2_buf_8 fanout1190 (.A(\vga_tetris._vgaController_io_pixelPosX[7] ),
    .X(net1190));
 sg13g2_buf_8 fanout1191 (.A(net1192),
    .X(net1191));
 sg13g2_buf_8 fanout1192 (.A(net1890),
    .X(net1192));
 sg13g2_buf_8 fanout1193 (.A(net1858),
    .X(net1193));
 sg13g2_buf_1 fanout1194 (.A(net1858),
    .X(net1194));
 sg13g2_buf_8 fanout1195 (.A(net1196),
    .X(net1195));
 sg13g2_buf_8 fanout1196 (.A(net1197),
    .X(net1196));
 sg13g2_buf_8 fanout1197 (.A(net1881),
    .X(net1197));
 sg13g2_buf_8 fanout1198 (.A(net1857),
    .X(net1198));
 sg13g2_buf_8 fanout1199 (.A(net1726),
    .X(net1199));
 sg13g2_buf_8 fanout1200 (.A(net1849),
    .X(net1200));
 sg13g2_buf_8 fanout1201 (.A(net1877),
    .X(net1201));
 sg13g2_buf_8 fanout1202 (.A(net1863),
    .X(net1202));
 sg13g2_buf_8 fanout1203 (.A(net1863),
    .X(net1203));
 sg13g2_buf_8 fanout1204 (.A(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[1] ),
    .X(net1204));
 sg13g2_buf_8 fanout1205 (.A(net1854),
    .X(net1205));
 sg13g2_buf_1 fanout1206 (.A(\vga_tetris.tetrisLogic.stateQ[4] ),
    .X(net1206));
 sg13g2_buf_8 fanout1207 (.A(net1208),
    .X(net1207));
 sg13g2_buf_2 fanout1208 (.A(net1851),
    .X(net1208));
 sg13g2_buf_8 fanout1209 (.A(net1210),
    .X(net1209));
 sg13g2_buf_8 fanout1210 (.A(net1875),
    .X(net1210));
 sg13g2_buf_8 fanout1211 (.A(net1736),
    .X(net1211));
 sg13g2_buf_8 fanout1212 (.A(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[1] ),
    .X(net1212));
 sg13g2_buf_8 fanout1213 (.A(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[3] ),
    .X(net1213));
 sg13g2_buf_8 fanout1214 (.A(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[2] ),
    .X(net1214));
 sg13g2_buf_8 fanout1215 (.A(\vga_tetris.tetrisLogic.stateQ[1] ),
    .X(net1215));
 sg13g2_buf_1 fanout1216 (.A(net1739),
    .X(net1216));
 sg13g2_buf_8 fanout1217 (.A(net1879),
    .X(net1217));
 sg13g2_buf_8 fanout1218 (.A(net1224),
    .X(net1218));
 sg13g2_buf_8 fanout1219 (.A(net1223),
    .X(net1219));
 sg13g2_buf_8 fanout1220 (.A(net1222),
    .X(net1220));
 sg13g2_buf_8 fanout1221 (.A(net1222),
    .X(net1221));
 sg13g2_buf_8 fanout1222 (.A(net1223),
    .X(net1222));
 sg13g2_buf_8 fanout1223 (.A(net1224),
    .X(net1223));
 sg13g2_buf_8 fanout1224 (.A(_0684_),
    .X(net1224));
 sg13g2_buf_8 fanout1225 (.A(net1226),
    .X(net1225));
 sg13g2_buf_8 fanout1226 (.A(net1227),
    .X(net1226));
 sg13g2_buf_8 fanout1227 (.A(_0684_),
    .X(net1227));
 sg13g2_buf_8 fanout1228 (.A(net1230),
    .X(net1228));
 sg13g2_buf_8 fanout1229 (.A(net1230),
    .X(net1229));
 sg13g2_buf_8 fanout1230 (.A(_0684_),
    .X(net1230));
 sg13g2_buf_8 fanout1231 (.A(net1232),
    .X(net1231));
 sg13g2_buf_8 fanout1232 (.A(net1233),
    .X(net1232));
 sg13g2_buf_2 fanout1233 (.A(net1237),
    .X(net1233));
 sg13g2_buf_8 fanout1234 (.A(net1236),
    .X(net1234));
 sg13g2_buf_2 fanout1235 (.A(net1236),
    .X(net1235));
 sg13g2_buf_8 fanout1236 (.A(net1237),
    .X(net1236));
 sg13g2_buf_8 fanout1237 (.A(net1246),
    .X(net1237));
 sg13g2_buf_8 fanout1238 (.A(net1239),
    .X(net1238));
 sg13g2_buf_8 fanout1239 (.A(net1246),
    .X(net1239));
 sg13g2_buf_8 fanout1240 (.A(net1242),
    .X(net1240));
 sg13g2_buf_2 fanout1241 (.A(net1242),
    .X(net1241));
 sg13g2_buf_8 fanout1242 (.A(net1246),
    .X(net1242));
 sg13g2_buf_8 fanout1243 (.A(net1245),
    .X(net1243));
 sg13g2_buf_8 fanout1244 (.A(net1245),
    .X(net1244));
 sg13g2_buf_8 fanout1245 (.A(net1246),
    .X(net1245));
 sg13g2_buf_8 fanout1246 (.A(rst_n),
    .X(net1246));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_tielo tt_um_vga_tetris_5 (.L_LO(net5));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_4_7_0_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\vga_tetris.vgaController.horizontalCounterQ[0] ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold2 (.A(\vga_tetris.msTimer.msTimerQ[0] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0015_),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold4 (.A(\vga_tetris.tetrisLogic.addOrRemoveShape.stateQ[1] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0068_),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold6 (.A(\vga_tetris.vgaController.horizontalCounterQ[1] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold7 (.A(\vga_tetris.boardMem.board_5[10] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold8 (.A(\vga_tetris.boardMem.board_15[12] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0524_),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold10 (.A(\vga_tetris.boardMem.board_4[17] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold11 (.A(\vga_tetris.boardMem.board_6[16] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0348_),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold13 (.A(\vga_tetris.boardMem.board_6[10] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold14 (.A(\vga_tetris.boardMem.board_13[9] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold15 (.A(\vga_tetris.boardMem.board_12[6] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold16 (.A(\vga_tetris.boardMem.board_14[7] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold17 (.A(\vga_tetris.boardMem.board_5[3] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold18 (.A(\vga_tetris.boardMem.board_8[7] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold19 (.A(\vga_tetris.boardMem.board_14[1] ),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold20 (.A(\vga_tetris.boardMem.board_14[18] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold21 (.A(\vga_tetris.boardMem.board_6[12] ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold22 (.A(\vga_tetris.boardMem.board_7[17] ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold23 (.A(\vga_tetris.boardMem.board_7[13] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold24 (.A(\vga_tetris.boardMem.board_7[5] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold25 (.A(\vga_tetris.boardMem.board_4[1] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold26 (.A(\vga_tetris.boardMem.board_9[11] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold27 (.A(\vga_tetris.boardMem.board_13[7] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold28 (.A(\vga_tetris.boardMem.board_15[9] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold29 (.A(\vga_tetris.boardMem.board_13[13] ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold30 (.A(\vga_tetris.boardMem.board_3[19] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold31 (.A(\vga_tetris.boardMem.board_14[19] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold32 (.A(\vga_tetris.boardMem.board_8[11] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold33 (.A(\vga_tetris.boardMem.board_12[9] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold34 (.A(\vga_tetris.vgaController.horizontalCounterQ[2] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold35 (.A(\vga_tetris.boardMem.board_10[13] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold36 (.A(\vga_tetris.boardMem.board_11[9] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold37 (.A(\vga_tetris.boardMem.board_15[3] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold38 (.A(\vga_tetris.boardMem.board_4[4] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold39 (.A(\vga_tetris.boardMem.board_13[11] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold40 (.A(\vga_tetris.boardMem.board_12[1] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0453_),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold42 (.A(\vga_tetris.boardMem.board_5[2] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold43 (.A(\vga_tetris.boardMem.board_3[14] ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold44 (.A(\vga_tetris.boardMem.board_7[10] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold45 (.A(\vga_tetris.boardMem.board_10[7] ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold46 (.A(\vga_tetris.boardMem.board_10[14] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold47 (.A(\vga_tetris.boardMem.board_15[11] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold48 (.A(\vga_tetris.boardMem.board_8[4] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold49 (.A(\vga_tetris.boardMem.board_8[9] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold50 (.A(\vga_tetris.boardMem.board_3[9] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold51 (.A(\vga_tetris.boardMem.board_7[14] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold52 (.A(\vga_tetris.boardMem.board_8[0] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0372_),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold54 (.A(\vga_tetris.boardMem.board_13[17] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0489_),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold56 (.A(\vga_tetris.boardMem.board_14[13] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold57 (.A(\vga_tetris.boardMem.board_8[13] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold58 (.A(\vga_tetris.boardMem.board_4[14] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold59 (.A(\vga_tetris.boardMem.board_4[11] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold60 (.A(\vga_tetris.boardMem.board_15[1] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold61 (.A(\vga_tetris.boardMem.board_11[10] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold62 (.A(\vga_tetris.boardMem.board_10[9] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold63 (.A(\vga_tetris.boardMem.board_7[15] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold64 (.A(\vga_tetris.boardMem.board_6[9] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold65 (.A(\vga_tetris.boardMem.board_8[8] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold66 (.A(\vga_tetris.boardMem.board_9[3] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0395_),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold68 (.A(\vga_tetris.boardMem.board_14[4] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold69 (.A(\vga_tetris.boardMem.board_9[10] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold70 (.A(\vga_tetris.boardMem.board_10[3] ),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold71 (.A(\vga_tetris.boardMem.board_5[5] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold72 (.A(\vga_tetris.boardMem.board_14[5] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0497_),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold74 (.A(\vga_tetris.boardMem.board_5[0] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold75 (.A(\vga_tetris.boardMem.board_10[2] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold76 (.A(\vga_tetris.boardMem.board_12[19] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0471_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold78 (.A(\vga_tetris.boardMem.board_10[11] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0423_),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold80 (.A(\vga_tetris.boardMem.board_4[2] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold81 (.A(\vga_tetris.boardMem.board_15[17] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0529_),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold83 (.A(\vga_tetris.boardMem.board_4[13] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold84 (.A(\vga_tetris.boardMem.board_12[4] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold85 (.A(\vga_tetris.boardMem.board_10[1] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold86 (.A(\vga_tetris.boardMem.board_4[6] ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold87 (.A(\vga_tetris.boardMem.board_15[14] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold88 (.A(\vga_tetris.boardMem.board_13[18] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold89 (.A(\vga_tetris.boardMem.board_4[18] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold90 (.A(\vga_tetris.boardMem.board_12[18] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold91 (.A(\vga_tetris.boardMem.board_9[8] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold92 (.A(\vga_tetris.boardMem.board_4[7] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold93 (.A(\vga_tetris.boardMem.board_13[10] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0482_),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold95 (.A(\vga_tetris.boardMem.board_9[18] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold96 (.A(\vga_tetris.boardMem.board_4[10] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold97 (.A(\vga_tetris.boardMem.board_3[2] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold98 (.A(\vga_tetris.boardMem.board_6[0] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold99 (.A(\vga_tetris.boardMem.board_11[2] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold100 (.A(\vga_tetris.boardMem.board_13[6] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold101 (.A(\vga_tetris.boardMem.board_6[5] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold102 (.A(\vga_tetris.boardMem.board_8[16] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold103 (.A(\vga_tetris.boardMem.board_3[15] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold104 (.A(\vga_tetris.boardMem.board_14[16] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold105 (.A(\vga_tetris.boardMem.board_13[2] ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold106 (.A(\vga_tetris.boardMem.board_9[9] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold107 (.A(\vga_tetris.boardMem.board_4[0] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold108 (.A(\vga_tetris.boardMem.board_6[4] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold109 (.A(\vga_tetris.boardMem.board_9[12] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold110 (.A(\vga_tetris.boardMem.board_12[16] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold111 (.A(\vga_tetris.boardMem.board_14[6] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold112 (.A(\vga_tetris.boardMem.board_7[11] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0363_),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold114 (.A(\vga_tetris.boardMem.board_3[1] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold115 (.A(\vga_tetris.boardMem.board_4[19] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold116 (.A(\vga_tetris.boardMem.board_4[5] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold117 (.A(\vga_tetris.boardMem.board_8[19] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold118 (.A(\vga_tetris.boardMem.board_3[0] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold119 (.A(\vga_tetris.boardMem.board_9[17] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold120 (.A(\vga_tetris.boardMem.board_6[14] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold121 (.A(\vga_tetris.boardMem.board_12[2] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold122 (.A(\vga_tetris.boardMem.board_7[1] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold123 (.A(\vga_tetris.boardMem.board_13[12] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold124 (.A(\vga_tetris.boardMem.board_11[0] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold125 (.A(\vga_tetris.boardMem.board_9[1] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0393_),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold127 (.A(\vga_tetris.boardMem.board_3[13] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold128 (.A(\vga_tetris.boardMem.board_11[6] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold129 (.A(\vga_tetris.boardMem.board_15[0] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold130 (.A(\vga_tetris.boardMem.board_14[2] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold131 (.A(\vga_tetris.boardMem.board_12[5] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold132 (.A(\vga_tetris.boardMem.board_4[12] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold133 (.A(\vga_tetris.boardMem.board_11[16] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold134 (.A(\vga_tetris.boardMem.board_12[11] ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold135 (.A(\vga_tetris.boardMem.board_11[13] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold136 (.A(\vga_tetris.boardMem.board_15[15] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold137 (.A(\vga_tetris.boardMem.board_11[4] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold138 (.A(\vga_tetris.boardMem.board_8[6] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold139 (.A(\vga_tetris.boardMem.board_5[19] ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0331_),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold141 (.A(\vga_tetris.boardMem.board_13[15] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold142 (.A(\vga_tetris.boardMem.board_9[19] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold143 (.A(\vga_tetris.boardMem.board_14[0] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold144 (.A(\vga_tetris.boardMem.board_7[6] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold145 (.A(\vga_tetris.boardMem.board_6[17] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold146 (.A(\vga_tetris.boardMem.board_4[16] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold147 (.A(\vga_tetris.boardMem.board_12[17] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold148 (.A(\vga_tetris.boardMem.board_14[8] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold149 (.A(\vga_tetris.boardMem.board_7[2] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold150 (.A(\vga_tetris.boardMem.board_6[13] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0345_),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold152 (.A(\vga_tetris.boardMem.board_14[12] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold153 (.A(\vga_tetris.boardMem.board_5[17] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold154 (.A(\vga_tetris.boardMem.board_9[0] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0392_),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold156 (.A(\vga_tetris.boardMem.board_14[11] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold157 (.A(\vga_tetris.boardMem.board_10[0] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold158 (.A(\vga_tetris.boardMem.board_7[0] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold159 (.A(\vga_tetris.boardMem.board_11[8] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold160 (.A(\vga_tetris.inputs.buttonTimerQ_2[0] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold161 (.A(_2393_),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0191_),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold163 (.A(\vga_tetris.boardMem.board_12[8] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold164 (.A(\vga_tetris.boardMem.board_6[2] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold165 (.A(\vga_tetris.boardMem.board_6[8] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold166 (.A(\vga_tetris.boardMem.board_6[19] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold167 (.A(\vga_tetris.boardMem.board_11[19] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold168 (.A(\vga_tetris.boardMem.board_11[12] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold169 (.A(\vga_tetris.boardMem.board_10[18] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold170 (.A(\vga_tetris.boardMem.board_11[5] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold171 (.A(\vga_tetris.boardMem.board_5[14] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold172 (.A(\vga_tetris.boardMem.board_5[11] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold173 (.A(\vga_tetris.boardMem.board_12[0] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0452_),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold175 (.A(\vga_tetris.boardMem.board_8[18] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold176 (.A(\vga_tetris.boardMem.board_6[1] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold177 (.A(\vga_tetris.boardMem.board_7[7] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold178 (.A(\vga_tetris.boardMem.board_13[0] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold179 (.A(\vga_tetris.boardMem.board_9[13] ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold180 (.A(\vga_tetris.boardMem.board_7[19] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0371_),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold182 (.A(\vga_tetris.boardMem.board_13[16] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold183 (.A(\vga_tetris.boardMem.board_6[15] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold184 (.A(\vga_tetris.boardMem.board_10[17] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold185 (.A(\vga_tetris.boardMem.board_3[8] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold186 (.A(\vga_tetris.boardMem.board_6[7] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold187 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[3] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0118_),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold189 (.A(\vga_tetris.boardMem.board_11[17] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold190 (.A(\vga_tetris.boardMem.board_6[11] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0343_),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold192 (.A(\vga_tetris.boardMem.board_12[14] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold193 (.A(\vga_tetris.boardMem.board_5[15] ),
    .X(net1247));
 sg13g2_dlygate4sd3_1 hold194 (.A(\vga_tetris.boardMem.board_4[9] ),
    .X(net1248));
 sg13g2_dlygate4sd3_1 hold195 (.A(\vga_tetris.boardMem.board_11[1] ),
    .X(net1249));
 sg13g2_dlygate4sd3_1 hold196 (.A(\vga_tetris.boardMem.board_14[17] ),
    .X(net1250));
 sg13g2_dlygate4sd3_1 hold197 (.A(\vga_tetris.boardMem.board_7[3] ),
    .X(net1251));
 sg13g2_dlygate4sd3_1 hold198 (.A(\vga_tetris.boardMem.board_3[17] ),
    .X(net1252));
 sg13g2_dlygate4sd3_1 hold199 (.A(\vga_tetris.boardMem.board_10[6] ),
    .X(net1253));
 sg13g2_dlygate4sd3_1 hold200 (.A(\vga_tetris.boardMem.board_10[19] ),
    .X(net1254));
 sg13g2_dlygate4sd3_1 hold201 (.A(\vga_tetris.boardMem.board_8[5] ),
    .X(net1255));
 sg13g2_dlygate4sd3_1 hold202 (.A(\vga_tetris.boardMem.board_4[15] ),
    .X(net1256));
 sg13g2_dlygate4sd3_1 hold203 (.A(\vga_tetris.boardMem.board_11[14] ),
    .X(net1257));
 sg13g2_dlygate4sd3_1 hold204 (.A(\vga_tetris.boardMem.board_7[9] ),
    .X(net1258));
 sg13g2_dlygate4sd3_1 hold205 (.A(\vga_tetris.boardMem.board_8[17] ),
    .X(net1259));
 sg13g2_dlygate4sd3_1 hold206 (.A(\vga_tetris.boardMem.board_8[2] ),
    .X(net1260));
 sg13g2_dlygate4sd3_1 hold207 (.A(\vga_tetris.boardMem.board_11[7] ),
    .X(net1261));
 sg13g2_dlygate4sd3_1 hold208 (.A(\vga_tetris.boardMem.board_6[6] ),
    .X(net1262));
 sg13g2_dlygate4sd3_1 hold209 (.A(\vga_tetris.boardMem.board_9[7] ),
    .X(net1263));
 sg13g2_dlygate4sd3_1 hold210 (.A(\vga_tetris.boardMem.board_11[18] ),
    .X(net1264));
 sg13g2_dlygate4sd3_1 hold211 (.A(\vga_tetris.boardMem.board_15[8] ),
    .X(net1265));
 sg13g2_dlygate4sd3_1 hold212 (.A(\vga_tetris.boardMem.board_12[13] ),
    .X(net1266));
 sg13g2_dlygate4sd3_1 hold213 (.A(\vga_tetris.boardMem.board_10[15] ),
    .X(net1267));
 sg13g2_dlygate4sd3_1 hold214 (.A(\vga_tetris.boardMem.board_5[8] ),
    .X(net1268));
 sg13g2_dlygate4sd3_1 hold215 (.A(\vga_tetris.boardMem.board_9[14] ),
    .X(net1269));
 sg13g2_dlygate4sd3_1 hold216 (.A(\vga_tetris.boardMem.board_3[10] ),
    .X(net1270));
 sg13g2_dlygate4sd3_1 hold217 (.A(\vga_tetris.boardMem.board_12[12] ),
    .X(net1271));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0464_),
    .X(net1272));
 sg13g2_dlygate4sd3_1 hold219 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[5] ),
    .X(net1273));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0120_),
    .X(net1274));
 sg13g2_dlygate4sd3_1 hold221 (.A(\vga_tetris.boardMem.board_10[10] ),
    .X(net1275));
 sg13g2_dlygate4sd3_1 hold222 (.A(\vga_tetris.boardMem.board_4[3] ),
    .X(net1276));
 sg13g2_dlygate4sd3_1 hold223 (.A(\vga_tetris.boardMem.board_9[16] ),
    .X(net1277));
 sg13g2_dlygate4sd3_1 hold224 (.A(\vga_tetris.boardMem.board_14[10] ),
    .X(net1278));
 sg13g2_dlygate4sd3_1 hold225 (.A(\vga_tetris.boardMem.board_14[9] ),
    .X(net1279));
 sg13g2_dlygate4sd3_1 hold226 (.A(\vga_tetris.boardMem.board_10[16] ),
    .X(net1280));
 sg13g2_dlygate4sd3_1 hold227 (.A(\vga_tetris.boardMem.board_5[4] ),
    .X(net1281));
 sg13g2_dlygate4sd3_1 hold228 (.A(\vga_tetris.boardMem.board_8[10] ),
    .X(net1282));
 sg13g2_dlygate4sd3_1 hold229 (.A(\vga_tetris.boardMem.board_9[2] ),
    .X(net1283));
 sg13g2_dlygate4sd3_1 hold230 (.A(\vga_tetris.boardMem.board_10[5] ),
    .X(net1284));
 sg13g2_dlygate4sd3_1 hold231 (.A(\vga_tetris.boardMem.board_9[5] ),
    .X(net1285));
 sg13g2_dlygate4sd3_1 hold232 (.A(\vga_tetris.boardMem.board_8[15] ),
    .X(net1286));
 sg13g2_dlygate4sd3_1 hold233 (.A(\vga_tetris.tetrisLogic._checkMoveAllowed_io_rowIndex[0] ),
    .X(net1287));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0094_),
    .X(net1288));
 sg13g2_dlygate4sd3_1 hold235 (.A(\vga_tetris.boardMem.board_5[6] ),
    .X(net1289));
 sg13g2_dlygate4sd3_1 hold236 (.A(\vga_tetris.boardMem.board_7[8] ),
    .X(net1290));
 sg13g2_dlygate4sd3_1 hold237 (.A(\vga_tetris.boardMem.board_6[18] ),
    .X(net1291));
 sg13g2_dlygate4sd3_1 hold238 (.A(\vga_tetris.boardMem.board_12[10] ),
    .X(net1292));
 sg13g2_dlygate4sd3_1 hold239 (.A(\vga_tetris.boardMem.board_11[15] ),
    .X(net1293));
 sg13g2_dlygate4sd3_1 hold240 (.A(\vga_tetris.boardMem.board_13[8] ),
    .X(net1294));
 sg13g2_dlygate4sd3_1 hold241 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[3] ),
    .X(net1295));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0053_),
    .X(net1296));
 sg13g2_dlygate4sd3_1 hold243 (.A(\vga_tetris.boardMem.board_5[7] ),
    .X(net1297));
 sg13g2_dlygate4sd3_1 hold244 (.A(\vga_tetris.boardMem.board_14[14] ),
    .X(net1298));
 sg13g2_dlygate4sd3_1 hold245 (.A(\vga_tetris.boardMem.board_5[12] ),
    .X(net1299));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0324_),
    .X(net1300));
 sg13g2_dlygate4sd3_1 hold247 (.A(\vga_tetris.boardMem.board_15[5] ),
    .X(net1301));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0517_),
    .X(net1302));
 sg13g2_dlygate4sd3_1 hold249 (.A(\vga_tetris.boardMem.board_14[3] ),
    .X(net1303));
 sg13g2_dlygate4sd3_1 hold250 (.A(\vga_tetris.boardMem.board_8[3] ),
    .X(net1304));
 sg13g2_dlygate4sd3_1 hold251 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[8] ),
    .X(net1305));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0058_),
    .X(net1306));
 sg13g2_dlygate4sd3_1 hold253 (.A(\vga_tetris.boardMem.board_7[18] ),
    .X(net1307));
 sg13g2_dlygate4sd3_1 hold254 (.A(\vga_tetris.boardMem.board_15[10] ),
    .X(net1308));
 sg13g2_dlygate4sd3_1 hold255 (.A(\vga_tetris.boardMem.board_5[13] ),
    .X(net1309));
 sg13g2_dlygate4sd3_1 hold256 (.A(\vga_tetris.boardMem.board_11[3] ),
    .X(net1310));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0435_),
    .X(net1311));
 sg13g2_dlygate4sd3_1 hold258 (.A(\vga_tetris.boardMem.board_5[18] ),
    .X(net1312));
 sg13g2_dlygate4sd3_1 hold259 (.A(\vga_tetris.boardMem.board_9[6] ),
    .X(net1313));
 sg13g2_dlygate4sd3_1 hold260 (.A(\vga_tetris.boardMem.board_15[4] ),
    .X(net1314));
 sg13g2_dlygate4sd3_1 hold261 (.A(\vga_tetris.boardMem.board_13[4] ),
    .X(net1315));
 sg13g2_dlygate4sd3_1 hold262 (.A(\vga_tetris.boardMem.board_3[3] ),
    .X(net1316));
 sg13g2_dlygate4sd3_1 hold263 (.A(\vga_tetris.boardMem.board_3[4] ),
    .X(net1317));
 sg13g2_dlygate4sd3_1 hold264 (.A(\vga_tetris.boardMem.board_4[8] ),
    .X(net1318));
 sg13g2_dlygate4sd3_1 hold265 (.A(\vga_tetris.boardMem.board_7[4] ),
    .X(net1319));
 sg13g2_dlygate4sd3_1 hold266 (.A(\vga_tetris.boardMem.board_10[8] ),
    .X(net1320));
 sg13g2_dlygate4sd3_1 hold267 (.A(\vga_tetris.boardMem.board_13[5] ),
    .X(net1321));
 sg13g2_dlygate4sd3_1 hold268 (.A(\vga_tetris.boardMem.board_15[2] ),
    .X(net1322));
 sg13g2_dlygate4sd3_1 hold269 (.A(\vga_tetris.boardMem.board_3[11] ),
    .X(net1323));
 sg13g2_dlygate4sd3_1 hold270 (.A(\vga_tetris.boardMem.board_12[15] ),
    .X(net1324));
 sg13g2_dlygate4sd3_1 hold271 (.A(\vga_tetris.boardMem.board_9[4] ),
    .X(net1325));
 sg13g2_dlygate4sd3_1 hold272 (.A(\vga_tetris.boardMem.board_15[18] ),
    .X(net1326));
 sg13g2_dlygate4sd3_1 hold273 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[18] ),
    .X(net1327));
 sg13g2_dlygate4sd3_1 hold274 (.A(_0133_),
    .X(net1328));
 sg13g2_dlygate4sd3_1 hold275 (.A(\vga_tetris.boardMem.board_5[9] ),
    .X(net1329));
 sg13g2_dlygate4sd3_1 hold276 (.A(\vga_tetris.boardMem.board_10[4] ),
    .X(net1330));
 sg13g2_dlygate4sd3_1 hold277 (.A(\vga_tetris.boardMem.board_13[19] ),
    .X(net1331));
 sg13g2_dlygate4sd3_1 hold278 (.A(\vga_tetris.boardMem.board_15[13] ),
    .X(net1332));
 sg13g2_dlygate4sd3_1 hold279 (.A(\vga_tetris.boardMem.board_5[1] ),
    .X(net1333));
 sg13g2_dlygate4sd3_1 hold280 (.A(\vga_tetris.boardMem.board_15[6] ),
    .X(net1334));
 sg13g2_dlygate4sd3_1 hold281 (.A(\vga_tetris.boardMem.board_12[7] ),
    .X(net1335));
 sg13g2_dlygate4sd3_1 hold282 (.A(\vga_tetris.boardMem.board_12[3] ),
    .X(net1336));
 sg13g2_dlygate4sd3_1 hold283 (.A(\vga_tetris.boardMem.board_15[19] ),
    .X(net1337));
 sg13g2_dlygate4sd3_1 hold284 (.A(\vga_tetris.boardMem.board_7[16] ),
    .X(net1338));
 sg13g2_dlygate4sd3_1 hold285 (.A(\vga_tetris.boardMem.board_14[15] ),
    .X(net1339));
 sg13g2_dlygate4sd3_1 hold286 (.A(\vga_tetris.boardMem.board_8[1] ),
    .X(net1340));
 sg13g2_dlygate4sd3_1 hold287 (.A(\vga_tetris.boardMem.board_3[12] ),
    .X(net1341));
 sg13g2_dlygate4sd3_1 hold288 (.A(\vga_tetris.boardMem.board_3[7] ),
    .X(net1342));
 sg13g2_dlygate4sd3_1 hold289 (.A(\vga_tetris.boardMem.board_3[5] ),
    .X(net1343));
 sg13g2_dlygate4sd3_1 hold290 (.A(\vga_tetris.boardMem.board_7[12] ),
    .X(net1344));
 sg13g2_dlygate4sd3_1 hold291 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[13] ),
    .X(net1345));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0084_),
    .X(net1346));
 sg13g2_dlygate4sd3_1 hold293 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[1] ),
    .X(net1347));
 sg13g2_dlygate4sd3_1 hold294 (.A(\vga_tetris.boardMem.board_6[3] ),
    .X(net1348));
 sg13g2_dlygate4sd3_1 hold295 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[9] ),
    .X(net1349));
 sg13g2_dlygate4sd3_1 hold296 (.A(\vga_tetris.boardMem.board_13[3] ),
    .X(net1350));
 sg13g2_dlygate4sd3_1 hold297 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[11] ),
    .X(net1351));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0082_),
    .X(net1352));
 sg13g2_dlygate4sd3_1 hold299 (.A(\vga_tetris.msTimer.msTimerQ[13] ),
    .X(net1353));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0028_),
    .X(net1354));
 sg13g2_dlygate4sd3_1 hold301 (.A(\vga_tetris.boardMem.board_3[6] ),
    .X(net1355));
 sg13g2_dlygate4sd3_1 hold302 (.A(\vga_tetris.boardMem.board_8[14] ),
    .X(net1356));
 sg13g2_dlygate4sd3_1 hold303 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[14] ),
    .X(net1357));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0064_),
    .X(net1358));
 sg13g2_dlygate4sd3_1 hold305 (.A(\vga_tetris.boardMem.board_3[16] ),
    .X(net1359));
 sg13g2_dlygate4sd3_1 hold306 (.A(\vga_tetris.boardMem.board_13[1] ),
    .X(net1360));
 sg13g2_dlygate4sd3_1 hold307 (.A(\vga_tetris.boardMem.board_15[7] ),
    .X(net1361));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0519_),
    .X(net1362));
 sg13g2_dlygate4sd3_1 hold309 (.A(\vga_tetris.boardMem.board_9[15] ),
    .X(net1363));
 sg13g2_dlygate4sd3_1 hold310 (.A(\vga_tetris.boardMem.board_11[11] ),
    .X(net1364));
 sg13g2_dlygate4sd3_1 hold311 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[4] ),
    .X(net1365));
 sg13g2_dlygate4sd3_1 hold312 (.A(\vga_tetris.boardMem.board_3[18] ),
    .X(net1366));
 sg13g2_dlygate4sd3_1 hold313 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[7] ),
    .X(net1367));
 sg13g2_dlygate4sd3_1 hold314 (.A(_1958_),
    .X(net1368));
 sg13g2_dlygate4sd3_1 hold315 (.A(_0078_),
    .X(net1369));
 sg13g2_dlygate4sd3_1 hold316 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[12] ),
    .X(net1370));
 sg13g2_dlygate4sd3_1 hold317 (.A(\vga_tetris.boardMem.board_15[16] ),
    .X(net1371));
 sg13g2_dlygate4sd3_1 hold318 (.A(\vga_tetris.boardMem.board_8[12] ),
    .X(net1372));
 sg13g2_dlygate4sd3_1 hold319 (.A(\vga_tetris.msTimer.msTimerQ[14] ),
    .X(net1373));
 sg13g2_dlygate4sd3_1 hold320 (.A(_1808_),
    .X(net1374));
 sg13g2_dlygate4sd3_1 hold321 (.A(\vga_tetris.boardMem.board_10[12] ),
    .X(net1375));
 sg13g2_dlygate4sd3_1 hold322 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[5] ),
    .X(net1376));
 sg13g2_dlygate4sd3_1 hold323 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[18] ),
    .X(net1377));
 sg13g2_dlygate4sd3_1 hold324 (.A(\vga_tetris.boardMem.board_5[16] ),
    .X(net1378));
 sg13g2_dlygate4sd3_1 hold325 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[3] ),
    .X(net1379));
 sg13g2_dlygate4sd3_1 hold326 (.A(\vga_tetris.tetrisLogic._checkMoveAllowed_io_rowIndex[1] ),
    .X(net1380));
 sg13g2_dlygate4sd3_1 hold327 (.A(_0095_),
    .X(net1381));
 sg13g2_dlygate4sd3_1 hold328 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[6] ),
    .X(net1382));
 sg13g2_dlygate4sd3_1 hold329 (.A(_0057_),
    .X(net1383));
 sg13g2_dlygate4sd3_1 hold330 (.A(\vga_tetris.msTimer.msTimerQ[2] ),
    .X(net1384));
 sg13g2_dlygate4sd3_1 hold331 (.A(_1786_),
    .X(net1385));
 sg13g2_dlygate4sd3_1 hold332 (.A(_0017_),
    .X(net1386));
 sg13g2_dlygate4sd3_1 hold333 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[0] ),
    .X(net1387));
 sg13g2_dlygate4sd3_1 hold334 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[6] ),
    .X(net1388));
 sg13g2_dlygate4sd3_1 hold335 (.A(_1951_),
    .X(net1389));
 sg13g2_dlygate4sd3_1 hold336 (.A(_0077_),
    .X(net1390));
 sg13g2_dlygate4sd3_1 hold337 (.A(\vga_tetris.boardMem.board_1[3] ),
    .X(net1391));
 sg13g2_dlygate4sd3_1 hold338 (.A(\vga_tetris.boardMem.board_1[11] ),
    .X(net1392));
 sg13g2_dlygate4sd3_1 hold339 (.A(_0243_),
    .X(net1393));
 sg13g2_dlygate4sd3_1 hold340 (.A(\vga_tetris.inputs.buttonTimerQ_0[6] ),
    .X(net1394));
 sg13g2_dlygate4sd3_1 hold341 (.A(_2361_),
    .X(net1395));
 sg13g2_dlygate4sd3_1 hold342 (.A(_0181_),
    .X(net1396));
 sg13g2_dlygate4sd3_1 hold343 (.A(\vga_tetris.boardMem.board_1[9] ),
    .X(net1397));
 sg13g2_dlygate4sd3_1 hold344 (.A(\vga_tetris.boardMem.board_0[15] ),
    .X(net1398));
 sg13g2_dlygate4sd3_1 hold345 (.A(_0227_),
    .X(net1399));
 sg13g2_dlygate4sd3_1 hold346 (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[0] ),
    .X(net1400));
 sg13g2_dlygate4sd3_1 hold347 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[10] ),
    .X(net1401));
 sg13g2_dlygate4sd3_1 hold348 (.A(\vga_tetris.boardMem.board_18[17] ),
    .X(net1402));
 sg13g2_dlygate4sd3_1 hold349 (.A(\vga_tetris.boardMem.board_2[2] ),
    .X(net1403));
 sg13g2_dlygate4sd3_1 hold350 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[1] ),
    .X(net1404));
 sg13g2_dlygate4sd3_1 hold351 (.A(_0116_),
    .X(net1405));
 sg13g2_dlygate4sd3_1 hold352 (.A(\vga_tetris.boardMem.board_13[14] ),
    .X(net1406));
 sg13g2_dlygate4sd3_1 hold353 (.A(\vga_tetris.boardMem.board_19[13] ),
    .X(net1407));
 sg13g2_dlygate4sd3_1 hold354 (.A(\vga_tetris.boardMem.board_17[15] ),
    .X(net1408));
 sg13g2_dlygate4sd3_1 hold355 (.A(_0567_),
    .X(net1409));
 sg13g2_dlygate4sd3_1 hold356 (.A(\vga_tetris.boardMem.board_18[0] ),
    .X(net1410));
 sg13g2_dlygate4sd3_1 hold357 (.A(\vga_tetris.tetrisLogic.gameOverLogic.buttonPressesCounterQ[0] ),
    .X(net1411));
 sg13g2_dlygate4sd3_1 hold358 (.A(_2218_),
    .X(net1412));
 sg13g2_dlygate4sd3_1 hold359 (.A(_0139_),
    .X(net1413));
 sg13g2_dlygate4sd3_1 hold360 (.A(\vga_tetris.boardMem.board_16[11] ),
    .X(net1414));
 sg13g2_dlygate4sd3_1 hold361 (.A(\vga_tetris.boardMem.board_17[11] ),
    .X(net1415));
 sg13g2_dlygate4sd3_1 hold362 (.A(_0563_),
    .X(net1416));
 sg13g2_dlygate4sd3_1 hold363 (.A(\vga_tetris.boardMem.board_0[17] ),
    .X(net1417));
 sg13g2_dlygate4sd3_1 hold364 (.A(\vga_tetris.boardMem.board_2[8] ),
    .X(net1418));
 sg13g2_dlygate4sd3_1 hold365 (.A(\vga_tetris.boardMem.board_16[16] ),
    .X(net1419));
 sg13g2_dlygate4sd3_1 hold366 (.A(_0548_),
    .X(net1420));
 sg13g2_dlygate4sd3_1 hold367 (.A(\vga_tetris.boardMem.board_19[7] ),
    .X(net1421));
 sg13g2_dlygate4sd3_1 hold368 (.A(\vga_tetris.boardMem.board_2[7] ),
    .X(net1422));
 sg13g2_dlygate4sd3_1 hold369 (.A(\vga_tetris.boardMem.board_17[18] ),
    .X(net1423));
 sg13g2_dlygate4sd3_1 hold370 (.A(\vga_tetris.boardMem.board_1[19] ),
    .X(net1424));
 sg13g2_dlygate4sd3_1 hold371 (.A(\vga_tetris.boardMem.board_1[7] ),
    .X(net1425));
 sg13g2_dlygate4sd3_1 hold372 (.A(\vga_tetris.boardMem.board_17[2] ),
    .X(net1426));
 sg13g2_dlygate4sd3_1 hold373 (.A(\vga_tetris.boardMem.board_1[18] ),
    .X(net1427));
 sg13g2_dlygate4sd3_1 hold374 (.A(\vga_tetris.boardMem.board_19[17] ),
    .X(net1428));
 sg13g2_dlygate4sd3_1 hold375 (.A(_0172_),
    .X(net1429));
 sg13g2_dlygate4sd3_1 hold376 (.A(\vga_tetris.boardMem.board_1[0] ),
    .X(net1430));
 sg13g2_dlygate4sd3_1 hold377 (.A(\vga_tetris.boardMem.board_17[19] ),
    .X(net1431));
 sg13g2_dlygate4sd3_1 hold378 (.A(\vga_tetris.boardMem.board_17[5] ),
    .X(net1432));
 sg13g2_dlygate4sd3_1 hold379 (.A(\vga_tetris.boardMem.board_0[2] ),
    .X(net1433));
 sg13g2_dlygate4sd3_1 hold380 (.A(_0214_),
    .X(net1434));
 sg13g2_dlygate4sd3_1 hold381 (.A(\vga_tetris.boardMem.board_16[19] ),
    .X(net1435));
 sg13g2_dlygate4sd3_1 hold382 (.A(_0551_),
    .X(net1436));
 sg13g2_dlygate4sd3_1 hold383 (.A(\vga_tetris.boardMem.board_2[16] ),
    .X(net1437));
 sg13g2_dlygate4sd3_1 hold384 (.A(_0268_),
    .X(net1438));
 sg13g2_dlygate4sd3_1 hold385 (.A(\vga_tetris.boardMem.board_16[14] ),
    .X(net1439));
 sg13g2_dlygate4sd3_1 hold386 (.A(\vga_tetris.boardMem.board_2[17] ),
    .X(net1440));
 sg13g2_dlygate4sd3_1 hold387 (.A(\vga_tetris.boardMem.board_1[2] ),
    .X(net1441));
 sg13g2_dlygate4sd3_1 hold388 (.A(\vga_tetris.boardMem.board_1[14] ),
    .X(net1442));
 sg13g2_dlygate4sd3_1 hold389 (.A(\vga_tetris.boardMem.board_19[9] ),
    .X(net1443));
 sg13g2_dlygate4sd3_1 hold390 (.A(\vga_tetris.boardMem.board_16[0] ),
    .X(net1444));
 sg13g2_dlygate4sd3_1 hold391 (.A(_0532_),
    .X(net1445));
 sg13g2_dlygate4sd3_1 hold392 (.A(\vga_tetris.boardMem.board_1[1] ),
    .X(net1446));
 sg13g2_dlygate4sd3_1 hold393 (.A(\vga_tetris.boardMem.board_16[15] ),
    .X(net1447));
 sg13g2_dlygate4sd3_1 hold394 (.A(\vga_tetris.boardMem.board_18[9] ),
    .X(net1448));
 sg13g2_dlygate4sd3_1 hold395 (.A(_0581_),
    .X(net1449));
 sg13g2_dlygate4sd3_1 hold396 (.A(\vga_tetris.boardMem.board_2[14] ),
    .X(net1450));
 sg13g2_dlygate4sd3_1 hold397 (.A(\vga_tetris.boardMem.board_2[10] ),
    .X(net1451));
 sg13g2_dlygate4sd3_1 hold398 (.A(\vga_tetris.boardMem.board_1[17] ),
    .X(net1452));
 sg13g2_dlygate4sd3_1 hold399 (.A(\vga_tetris.boardMem.board_17[14] ),
    .X(net1453));
 sg13g2_dlygate4sd3_1 hold400 (.A(\vga_tetris.boardMem.board_18[18] ),
    .X(net1454));
 sg13g2_dlygate4sd3_1 hold401 (.A(\vga_tetris.boardMem.board_2[12] ),
    .X(net1455));
 sg13g2_dlygate4sd3_1 hold402 (.A(\vga_tetris.boardMem.board_2[18] ),
    .X(net1456));
 sg13g2_dlygate4sd3_1 hold403 (.A(\vga_tetris.boardMem.board_17[6] ),
    .X(net1457));
 sg13g2_dlygate4sd3_1 hold404 (.A(\vga_tetris.boardMem.board_19[5] ),
    .X(net1458));
 sg13g2_dlygate4sd3_1 hold405 (.A(\vga_tetris.boardMem.board_18[14] ),
    .X(net1459));
 sg13g2_dlygate4sd3_1 hold406 (.A(\vga_tetris.boardMem.board_17[9] ),
    .X(net1460));
 sg13g2_dlygate4sd3_1 hold407 (.A(\vga_tetris.boardMem.board_0[13] ),
    .X(net1461));
 sg13g2_dlygate4sd3_1 hold408 (.A(\vga_tetris.boardMem.board_16[1] ),
    .X(net1462));
 sg13g2_dlygate4sd3_1 hold409 (.A(\vga_tetris.boardMem.board_18[2] ),
    .X(net1463));
 sg13g2_dlygate4sd3_1 hold410 (.A(\vga_tetris.boardMem.board_16[6] ),
    .X(net1464));
 sg13g2_dlygate4sd3_1 hold411 (.A(\vga_tetris.boardMem.board_19[0] ),
    .X(net1465));
 sg13g2_dlygate4sd3_1 hold412 (.A(\vga_tetris.boardMem.board_0[9] ),
    .X(net1466));
 sg13g2_dlygate4sd3_1 hold413 (.A(\vga_tetris.boardMem.board_0[6] ),
    .X(net1467));
 sg13g2_dlygate4sd3_1 hold414 (.A(_0218_),
    .X(net1468));
 sg13g2_dlygate4sd3_1 hold415 (.A(\vga_tetris.boardMem.board_18[15] ),
    .X(net1469));
 sg13g2_dlygate4sd3_1 hold416 (.A(\vga_tetris.boardMem.board_0[4] ),
    .X(net1470));
 sg13g2_dlygate4sd3_1 hold417 (.A(_0216_),
    .X(net1471));
 sg13g2_dlygate4sd3_1 hold418 (.A(\vga_tetris.boardMem.board_16[4] ),
    .X(net1472));
 sg13g2_dlygate4sd3_1 hold419 (.A(\vga_tetris.boardMem.board_19[3] ),
    .X(net1473));
 sg13g2_dlygate4sd3_1 hold420 (.A(\vga_tetris.boardMem.board_0[12] ),
    .X(net1474));
 sg13g2_dlygate4sd3_1 hold421 (.A(_0224_),
    .X(net1475));
 sg13g2_dlygate4sd3_1 hold422 (.A(\vga_tetris.boardMem.board_0[16] ),
    .X(net1476));
 sg13g2_dlygate4sd3_1 hold423 (.A(\vga_tetris.boardMem.board_16[18] ),
    .X(net1477));
 sg13g2_dlygate4sd3_1 hold424 (.A(\vga_tetris.vgaController.verticalCounterQ[0] ),
    .X(net1478));
 sg13g2_dlygate4sd3_1 hold425 (.A(_0593_),
    .X(net1479));
 sg13g2_dlygate4sd3_1 hold426 (.A(\vga_tetris.boardMem.board_16[9] ),
    .X(net1480));
 sg13g2_dlygate4sd3_1 hold427 (.A(_0541_),
    .X(net1481));
 sg13g2_dlygate4sd3_1 hold428 (.A(\vga_tetris.boardMem.board_19[6] ),
    .X(net1482));
 sg13g2_dlygate4sd3_1 hold429 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[5] ),
    .X(net1483));
 sg13g2_dlygate4sd3_1 hold430 (.A(\vga_tetris.boardMem.board_2[15] ),
    .X(net1484));
 sg13g2_dlygate4sd3_1 hold431 (.A(\vga_tetris.boardMem.board_1[15] ),
    .X(net1485));
 sg13g2_dlygate4sd3_1 hold432 (.A(\vga_tetris.boardMem.board_18[12] ),
    .X(net1486));
 sg13g2_dlygate4sd3_1 hold433 (.A(\vga_tetris.boardMem.board_2[5] ),
    .X(net1487));
 sg13g2_dlygate4sd3_1 hold434 (.A(\vga_tetris.boardMem.board_16[5] ),
    .X(net1488));
 sg13g2_dlygate4sd3_1 hold435 (.A(\vga_tetris.boardMem.board_18[19] ),
    .X(net1489));
 sg13g2_dlygate4sd3_1 hold436 (.A(\vga_tetris.boardMem.board_0[11] ),
    .X(net1490));
 sg13g2_dlygate4sd3_1 hold437 (.A(_0223_),
    .X(net1491));
 sg13g2_dlygate4sd3_1 hold438 (.A(\vga_tetris.boardMem.board_1[8] ),
    .X(net1492));
 sg13g2_dlygate4sd3_1 hold439 (.A(\vga_tetris.boardMem.board_17[8] ),
    .X(net1493));
 sg13g2_dlygate4sd3_1 hold440 (.A(\vga_tetris.boardMem.board_1[4] ),
    .X(net1494));
 sg13g2_dlygate4sd3_1 hold441 (.A(\vga_tetris.boardMem.board_17[10] ),
    .X(net1495));
 sg13g2_dlygate4sd3_1 hold442 (.A(\vga_tetris.boardMem.board_18[16] ),
    .X(net1496));
 sg13g2_dlygate4sd3_1 hold443 (.A(\vga_tetris.boardMem.board_2[6] ),
    .X(net1497));
 sg13g2_dlygate4sd3_1 hold444 (.A(\vga_tetris.boardMem.board_16[12] ),
    .X(net1498));
 sg13g2_dlygate4sd3_1 hold445 (.A(\vga_tetris.boardMem.board_18[7] ),
    .X(net1499));
 sg13g2_dlygate4sd3_1 hold446 (.A(\vga_tetris.boardMem.board_19[2] ),
    .X(net1500));
 sg13g2_dlygate4sd3_1 hold447 (.A(\vga_tetris.boardMem.board_19[16] ),
    .X(net1501));
 sg13g2_dlygate4sd3_1 hold448 (.A(_0171_),
    .X(net1502));
 sg13g2_dlygate4sd3_1 hold449 (.A(\vga_tetris.boardMem.board_17[0] ),
    .X(net1503));
 sg13g2_dlygate4sd3_1 hold450 (.A(\vga_tetris.boardMem.board_2[0] ),
    .X(net1504));
 sg13g2_dlygate4sd3_1 hold451 (.A(\vga_tetris.boardMem.board_17[3] ),
    .X(net1505));
 sg13g2_dlygate4sd3_1 hold452 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[8] ),
    .X(net1506));
 sg13g2_dlygate4sd3_1 hold453 (.A(_0079_),
    .X(net1507));
 sg13g2_dlygate4sd3_1 hold454 (.A(\vga_tetris.boardMem.board_18[11] ),
    .X(net1508));
 sg13g2_dlygate4sd3_1 hold455 (.A(\vga_tetris.boardMem.board_16[7] ),
    .X(net1509));
 sg13g2_dlygate4sd3_1 hold456 (.A(\vga_tetris.boardMem.board_0[14] ),
    .X(net1510));
 sg13g2_dlygate4sd3_1 hold457 (.A(\vga_tetris.boardMem.board_1[6] ),
    .X(net1511));
 sg13g2_dlygate4sd3_1 hold458 (.A(\vga_tetris.boardMem.board_2[11] ),
    .X(net1512));
 sg13g2_dlygate4sd3_1 hold459 (.A(\vga_tetris.boardMem.board_2[1] ),
    .X(net1513));
 sg13g2_dlygate4sd3_1 hold460 (.A(\vga_tetris.boardMem.board_17[17] ),
    .X(net1514));
 sg13g2_dlygate4sd3_1 hold461 (.A(\vga_tetris.boardMem.board_19[14] ),
    .X(net1515));
 sg13g2_dlygate4sd3_1 hold462 (.A(\vga_tetris.boardMem.board_18[5] ),
    .X(net1516));
 sg13g2_dlygate4sd3_1 hold463 (.A(\vga_tetris.boardMem.board_18[8] ),
    .X(net1517));
 sg13g2_dlygate4sd3_1 hold464 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[10] ),
    .X(net1518));
 sg13g2_dlygate4sd3_1 hold465 (.A(\vga_tetris.boardMem.board_1[13] ),
    .X(net1519));
 sg13g2_dlygate4sd3_1 hold466 (.A(_0245_),
    .X(net1520));
 sg13g2_dlygate4sd3_1 hold467 (.A(\vga_tetris.boardMem.board_19[19] ),
    .X(net1521));
 sg13g2_dlygate4sd3_1 hold468 (.A(\vga_tetris.boardMem.board_17[13] ),
    .X(net1522));
 sg13g2_dlygate4sd3_1 hold469 (.A(\vga_tetris.vgaController.horizontalCounterQ[3] ),
    .X(net1523));
 sg13g2_dlygate4sd3_1 hold470 (.A(\vga_tetris.boardMem.board_1[16] ),
    .X(net1524));
 sg13g2_dlygate4sd3_1 hold471 (.A(\vga_tetris.boardMem.board_18[1] ),
    .X(net1525));
 sg13g2_dlygate4sd3_1 hold472 (.A(\vga_tetris.boardMem.board_18[3] ),
    .X(net1526));
 sg13g2_dlygate4sd3_1 hold473 (.A(\vga_tetris.boardMem.board_19[15] ),
    .X(net1527));
 sg13g2_dlygate4sd3_1 hold474 (.A(\vga_tetris.boardMem.board_2[13] ),
    .X(net1528));
 sg13g2_dlygate4sd3_1 hold475 (.A(_0265_),
    .X(net1529));
 sg13g2_dlygate4sd3_1 hold476 (.A(\vga_tetris.boardMem.board_0[10] ),
    .X(net1530));
 sg13g2_dlygate4sd3_1 hold477 (.A(\vga_tetris.boardMem.board_17[16] ),
    .X(net1531));
 sg13g2_dlygate4sd3_1 hold478 (.A(\vga_tetris.boardMem.board_19[4] ),
    .X(net1532));
 sg13g2_dlygate4sd3_1 hold479 (.A(\vga_tetris.tetrisLogic.shapeDropTimerQ[1] ),
    .X(net1533));
 sg13g2_dlygate4sd3_1 hold480 (.A(_1881_),
    .X(net1534));
 sg13g2_dlygate4sd3_1 hold481 (.A(_0045_),
    .X(net1535));
 sg13g2_dlygate4sd3_1 hold482 (.A(\vga_tetris.boardMem.board_16[3] ),
    .X(net1536));
 sg13g2_dlygate4sd3_1 hold483 (.A(\vga_tetris.boardMem.board_16[13] ),
    .X(net1537));
 sg13g2_dlygate4sd3_1 hold484 (.A(_0545_),
    .X(net1538));
 sg13g2_dlygate4sd3_1 hold485 (.A(\vga_tetris.boardMem.board_0[0] ),
    .X(net1539));
 sg13g2_dlygate4sd3_1 hold486 (.A(\vga_tetris.boardMem.board_18[10] ),
    .X(net1540));
 sg13g2_dlygate4sd3_1 hold487 (.A(\vga_tetris.boardMem.board_19[18] ),
    .X(net1541));
 sg13g2_dlygate4sd3_1 hold488 (.A(\vga_tetris.boardMem.board_19[10] ),
    .X(net1542));
 sg13g2_dlygate4sd3_1 hold489 (.A(\vga_tetris.boardMem.board_16[8] ),
    .X(net1543));
 sg13g2_dlygate4sd3_1 hold490 (.A(_0540_),
    .X(net1544));
 sg13g2_dlygate4sd3_1 hold491 (.A(\vga_tetris.boardMem.board_1[10] ),
    .X(net1545));
 sg13g2_dlygate4sd3_1 hold492 (.A(\vga_tetris.boardMem.board_1[12] ),
    .X(net1546));
 sg13g2_dlygate4sd3_1 hold493 (.A(\vga_tetris.boardMem.board_0[1] ),
    .X(net1547));
 sg13g2_dlygate4sd3_1 hold494 (.A(\vga_tetris.boardMem.board_19[8] ),
    .X(net1548));
 sg13g2_dlygate4sd3_1 hold495 (.A(\vga_tetris.boardMem.board_17[7] ),
    .X(net1549));
 sg13g2_dlygate4sd3_1 hold496 (.A(_0559_),
    .X(net1550));
 sg13g2_dlygate4sd3_1 hold497 (.A(\vga_tetris.boardMem.board_2[4] ),
    .X(net1551));
 sg13g2_dlygate4sd3_1 hold498 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[2] ),
    .X(net1552));
 sg13g2_dlygate4sd3_1 hold499 (.A(_0109_),
    .X(net1553));
 sg13g2_dlygate4sd3_1 hold500 (.A(\vga_tetris.boardMem.board_19[1] ),
    .X(net1554));
 sg13g2_dlygate4sd3_1 hold501 (.A(\vga_tetris.boardMem.board_0[19] ),
    .X(net1555));
 sg13g2_dlygate4sd3_1 hold502 (.A(\vga_tetris.boardMem.board_0[7] ),
    .X(net1556));
 sg13g2_dlygate4sd3_1 hold503 (.A(\vga_tetris.boardMem.board_18[13] ),
    .X(net1557));
 sg13g2_dlygate4sd3_1 hold504 (.A(\vga_tetris.boardMem.board_2[9] ),
    .X(net1558));
 sg13g2_dlygate4sd3_1 hold505 (.A(\vga_tetris.boardMem.board_0[3] ),
    .X(net1559));
 sg13g2_dlygate4sd3_1 hold506 (.A(\vga_tetris.boardMem.board_17[1] ),
    .X(net1560));
 sg13g2_dlygate4sd3_1 hold507 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[15] ),
    .X(net1561));
 sg13g2_dlygate4sd3_1 hold508 (.A(\vga_tetris.tetrisLogic.checkMoveAllowed.checkIsRunningQ ),
    .X(net1562));
 sg13g2_dlygate4sd3_1 hold509 (.A(\vga_tetris.boardMem.board_16[10] ),
    .X(net1563));
 sg13g2_dlygate4sd3_1 hold510 (.A(\vga_tetris.boardMem.board_0[5] ),
    .X(net1564));
 sg13g2_dlygate4sd3_1 hold511 (.A(\vga_tetris.inputs.buttonTimerQ_2[1] ),
    .X(net1565));
 sg13g2_dlygate4sd3_1 hold512 (.A(_2394_),
    .X(net1566));
 sg13g2_dlygate4sd3_1 hold513 (.A(_0192_),
    .X(net1567));
 sg13g2_dlygate4sd3_1 hold514 (.A(\vga_tetris.boardMem.board_0[18] ),
    .X(net1568));
 sg13g2_dlygate4sd3_1 hold515 (.A(\vga_tetris.boardMem.board_16[17] ),
    .X(net1569));
 sg13g2_dlygate4sd3_1 hold516 (.A(_0549_),
    .X(net1570));
 sg13g2_dlygate4sd3_1 hold517 (.A(\vga_tetris.boardMem.board_19[11] ),
    .X(net1571));
 sg13g2_dlygate4sd3_1 hold518 (.A(\vga_tetris.boardMem.board_0[8] ),
    .X(net1572));
 sg13g2_dlygate4sd3_1 hold519 (.A(\vga_tetris.boardMem.board_18[6] ),
    .X(net1573));
 sg13g2_dlygate4sd3_1 hold520 (.A(\vga_tetris.boardMem.board_2[19] ),
    .X(net1574));
 sg13g2_dlygate4sd3_1 hold521 (.A(\vga_tetris.boardMem.board_1[5] ),
    .X(net1575));
 sg13g2_dlygate4sd3_1 hold522 (.A(\vga_tetris.boardMem.board_2[3] ),
    .X(net1576));
 sg13g2_dlygate4sd3_1 hold523 (.A(\vga_tetris.boardMem.board_17[12] ),
    .X(net1577));
 sg13g2_dlygate4sd3_1 hold524 (.A(_0564_),
    .X(net1578));
 sg13g2_dlygate4sd3_1 hold525 (.A(\vga_tetris._vgaController_io_pixelPosX[8] ),
    .X(net1579));
 sg13g2_dlygate4sd3_1 hold526 (.A(_0611_),
    .X(net1580));
 sg13g2_dlygate4sd3_1 hold527 (.A(\vga_tetris.boardMem.board_16[2] ),
    .X(net1581));
 sg13g2_dlygate4sd3_1 hold528 (.A(\vga_tetris.vgaController.verticalCounterQ[1] ),
    .X(net1582));
 sg13g2_dlygate4sd3_1 hold529 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[1] ),
    .X(net1583));
 sg13g2_dlygate4sd3_1 hold530 (.A(_0051_),
    .X(net1584));
 sg13g2_dlygate4sd3_1 hold531 (.A(\vga_tetris._tetrisLogic_io_score_2[2] ),
    .X(net1585));
 sg13g2_dlygate4sd3_1 hold532 (.A(_2228_),
    .X(net1586));
 sg13g2_dlygate4sd3_1 hold533 (.A(_0144_),
    .X(net1587));
 sg13g2_dlygate4sd3_1 hold534 (.A(\vga_tetris.boardMem.board_18[4] ),
    .X(net1588));
 sg13g2_dlygate4sd3_1 hold535 (.A(\vga_tetris._inputs_io_rotateButtonActive ),
    .X(net1589));
 sg13g2_dlygate4sd3_1 hold536 (.A(\vga_tetris.boardMem.board_17[4] ),
    .X(net1590));
 sg13g2_dlygate4sd3_1 hold537 (.A(\vga_tetris.vgaController.verticalCounterQ[4] ),
    .X(net1591));
 sg13g2_dlygate4sd3_1 hold538 (.A(_2875_),
    .X(net1592));
 sg13g2_dlygate4sd3_1 hold539 (.A(\vga_tetris.vgaController.verticalCounterQ[3] ),
    .X(net1593));
 sg13g2_dlygate4sd3_1 hold540 (.A(_0596_),
    .X(net1594));
 sg13g2_dlygate4sd3_1 hold541 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[2] ),
    .X(net1595));
 sg13g2_dlygate4sd3_1 hold542 (.A(\vga_tetris._tetrisLogic_io_score_1[2] ),
    .X(net1596));
 sg13g2_dlygate4sd3_1 hold543 (.A(_2236_),
    .X(net1597));
 sg13g2_dlygate4sd3_1 hold544 (.A(_0148_),
    .X(net1598));
 sg13g2_dlygate4sd3_1 hold545 (.A(\vga_tetris._vgaController_io_pixelPosX[1] ),
    .X(net1599));
 sg13g2_dlygate4sd3_1 hold546 (.A(_0604_),
    .X(net1600));
 sg13g2_dlygate4sd3_1 hold547 (.A(\vga_tetris.boardMem.board_19[12] ),
    .X(net1601));
 sg13g2_dlygate4sd3_1 hold548 (.A(\vga_tetris.vgaController.verticalCounterQ[8] ),
    .X(net1602));
 sg13g2_dlygate4sd3_1 hold549 (.A(_0601_),
    .X(net1603));
 sg13g2_dlygate4sd3_1 hold550 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[3] ),
    .X(net1604));
 sg13g2_dlygate4sd3_1 hold551 (.A(_0110_),
    .X(net1605));
 sg13g2_dlygate4sd3_1 hold552 (.A(\vga_tetris.vgaController.verticalCounterQ[2] ),
    .X(net1606));
 sg13g2_dlygate4sd3_1 hold553 (.A(_0595_),
    .X(net1607));
 sg13g2_dlygate4sd3_1 hold554 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[15] ),
    .X(net1608));
 sg13g2_dlygate4sd3_1 hold555 (.A(_2004_),
    .X(net1609));
 sg13g2_dlygate4sd3_1 hold556 (.A(\vga_tetris._vgaController_io_pixelPosY[0] ),
    .X(net1610));
 sg13g2_dlygate4sd3_1 hold557 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[2] ),
    .X(net1611));
 sg13g2_dlygate4sd3_1 hold558 (.A(_2090_),
    .X(net1612));
 sg13g2_dlygate4sd3_1 hold559 (.A(_0592_),
    .X(net1613));
 sg13g2_dlygate4sd3_1 hold560 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[0] ),
    .X(net1614));
 sg13g2_dlygate4sd3_1 hold561 (.A(_1839_),
    .X(net1615));
 sg13g2_dlygate4sd3_1 hold562 (.A(\vga_tetris.inputs.buttonTimerQ_1[6] ),
    .X(net1616));
 sg13g2_dlygate4sd3_1 hold563 (.A(_2385_),
    .X(net1617));
 sg13g2_dlygate4sd3_1 hold564 (.A(_0189_),
    .X(net1618));
 sg13g2_dlygate4sd3_1 hold565 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[4] ),
    .X(net1619));
 sg13g2_dlygate4sd3_1 hold566 (.A(_1947_),
    .X(net1620));
 sg13g2_dlygate4sd3_1 hold567 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[19] ),
    .X(net1621));
 sg13g2_dlygate4sd3_1 hold568 (.A(_2024_),
    .X(net1622));
 sg13g2_dlygate4sd3_1 hold569 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_rowIndex[1] ),
    .X(net1623));
 sg13g2_dlygate4sd3_1 hold570 (.A(_1911_),
    .X(net1624));
 sg13g2_dlygate4sd3_1 hold571 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[14] ),
    .X(net1625));
 sg13g2_dlygate4sd3_1 hold572 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[12] ),
    .X(net1626));
 sg13g2_dlygate4sd3_1 hold573 (.A(_0062_),
    .X(net1627));
 sg13g2_dlygate4sd3_1 hold574 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[11] ),
    .X(net1628));
 sg13g2_dlygate4sd3_1 hold575 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[9] ),
    .X(net1629));
 sg13g2_dlygate4sd3_1 hold576 (.A(\vga_tetris.inputs.buttonTimerQ_0[0] ),
    .X(net1630));
 sg13g2_dlygate4sd3_1 hold577 (.A(\vga_tetris.inputs.buttonTimerQ_1[7] ),
    .X(net1631));
 sg13g2_dlygate4sd3_1 hold578 (.A(_2387_),
    .X(net1632));
 sg13g2_dlygate4sd3_1 hold579 (.A(_0190_),
    .X(net1633));
 sg13g2_dlygate4sd3_1 hold580 (.A(\vga_tetris.msTimer.msTimerQ[3] ),
    .X(net1634));
 sg13g2_dlygate4sd3_1 hold581 (.A(_1788_),
    .X(net1635));
 sg13g2_dlygate4sd3_1 hold582 (.A(_0018_),
    .X(net1636));
 sg13g2_dlygate4sd3_1 hold583 (.A(\vga_tetris.inputs.buttonTimerQ_1[0] ),
    .X(net1637));
 sg13g2_dlygate4sd3_1 hold584 (.A(_2371_),
    .X(net1638));
 sg13g2_dlygate4sd3_1 hold585 (.A(_0183_),
    .X(net1639));
 sg13g2_dlygate4sd3_1 hold586 (.A(\vga_tetris._vgaController_io_pixelPosY[8] ),
    .X(net1640));
 sg13g2_dlygate4sd3_1 hold587 (.A(_0621_),
    .X(net1641));
 sg13g2_dlygate4sd3_1 hold588 (.A(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[1] ),
    .X(net1642));
 sg13g2_dlygate4sd3_1 hold589 (.A(_1840_),
    .X(net1643));
 sg13g2_dlygate4sd3_1 hold590 (.A(\vga_tetris.msTimer.msTimerQ[4] ),
    .X(net1644));
 sg13g2_dlygate4sd3_1 hold591 (.A(_1790_),
    .X(net1645));
 sg13g2_dlygate4sd3_1 hold592 (.A(_0019_),
    .X(net1646));
 sg13g2_dlygate4sd3_1 hold593 (.A(\vga_tetris.vgaController.horizontalCounterQ[5] ),
    .X(net1647));
 sg13g2_dlygate4sd3_1 hold594 (.A(_1768_),
    .X(net1648));
 sg13g2_dlygate4sd3_1 hold595 (.A(_0010_),
    .X(net1649));
 sg13g2_dlygate4sd3_1 hold596 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[10] ),
    .X(net1650));
 sg13g2_dlygate4sd3_1 hold597 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[1] ),
    .X(net1651));
 sg13g2_dlygate4sd3_1 hold598 (.A(_0108_),
    .X(net1652));
 sg13g2_dlygate4sd3_1 hold599 (.A(\vga_tetris.msTimer.msTimerQ[7] ),
    .X(net1653));
 sg13g2_dlygate4sd3_1 hold600 (.A(_1795_),
    .X(net1654));
 sg13g2_dlygate4sd3_1 hold601 (.A(_0022_),
    .X(net1655));
 sg13g2_dlygate4sd3_1 hold602 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[14] ),
    .X(net1656));
 sg13g2_dlygate4sd3_1 hold603 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[13] ),
    .X(net1657));
 sg13g2_dlygate4sd3_1 hold604 (.A(\vga_tetris.msTimer.msTimerQ[5] ),
    .X(net1658));
 sg13g2_dlygate4sd3_1 hold605 (.A(_0020_),
    .X(net1659));
 sg13g2_dlygate4sd3_1 hold606 (.A(\vga_tetris._tetrisLogic_io_score_3[0] ),
    .X(net1660));
 sg13g2_dlygate4sd3_1 hold607 (.A(_2204_),
    .X(net1661));
 sg13g2_dlygate4sd3_1 hold608 (.A(_0135_),
    .X(net1662));
 sg13g2_dlygate4sd3_1 hold609 (.A(\vga_tetris.tetrisLogic.tetrisLFSRPseudoRandomNumGen.lfsrQ[13] ),
    .X(net1663));
 sg13g2_dlygate4sd3_1 hold610 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[8] ),
    .X(net1664));
 sg13g2_dlygate4sd3_1 hold611 (.A(\vga_tetris.vgaController.horizontalCounterQ[7] ),
    .X(net1665));
 sg13g2_dlygate4sd3_1 hold612 (.A(_1772_),
    .X(net1666));
 sg13g2_dlygate4sd3_1 hold613 (.A(\vga_tetris._vgaController_io_pixelPosY[9] ),
    .X(net1667));
 sg13g2_dlygate4sd3_1 hold614 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[11] ),
    .X(net1668));
 sg13g2_dlygate4sd3_1 hold615 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[6] ),
    .X(net1669));
 sg13g2_dlygate4sd3_1 hold616 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[2] ),
    .X(net1670));
 sg13g2_dlygate4sd3_1 hold617 (.A(_2174_),
    .X(net1671));
 sg13g2_dlygate4sd3_1 hold618 (.A(_0117_),
    .X(net1672));
 sg13g2_dlygate4sd3_1 hold619 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[15] ),
    .X(net1673));
 sg13g2_dlygate4sd3_1 hold620 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[4] ),
    .X(net1674));
 sg13g2_dlygate4sd3_1 hold621 (.A(\vga_tetris.inputs.buttonTimerQ_2[7] ),
    .X(net1675));
 sg13g2_dlygate4sd3_1 hold622 (.A(_2408_),
    .X(net1676));
 sg13g2_dlygate4sd3_1 hold623 (.A(_0198_),
    .X(net1677));
 sg13g2_dlygate4sd3_1 hold624 (.A(\vga_tetris.vgaController.horizontalCounterQ[6] ),
    .X(net1678));
 sg13g2_dlygate4sd3_1 hold625 (.A(_0011_),
    .X(net1679));
 sg13g2_dlygate4sd3_1 hold626 (.A(\vga_tetris.tetrisLogic.stateQ[3] ),
    .X(net1680));
 sg13g2_dlygate4sd3_1 hold627 (.A(_1720_),
    .X(net1681));
 sg13g2_dlygate4sd3_1 hold628 (.A(_0002_),
    .X(net1682));
 sg13g2_dlygate4sd3_1 hold629 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[12] ),
    .X(net1683));
 sg13g2_dlygate4sd3_1 hold630 (.A(\vga_tetris._inputs_io_downButtonActive ),
    .X(net1684));
 sg13g2_dlygate4sd3_1 hold631 (.A(_0210_),
    .X(net1685));
 sg13g2_dlygate4sd3_1 hold632 (.A(\vga_tetris._tetrisLogic_io_score_3[3] ),
    .X(net1686));
 sg13g2_dlygate4sd3_1 hold633 (.A(_2211_),
    .X(net1687));
 sg13g2_dlygate4sd3_1 hold634 (.A(_0136_),
    .X(net1688));
 sg13g2_dlygate4sd3_1 hold635 (.A(\vga_tetris.inputs.buttonTimerQ_2[6] ),
    .X(net1689));
 sg13g2_dlygate4sd3_1 hold636 (.A(_2407_),
    .X(net1690));
 sg13g2_dlygate4sd3_1 hold637 (.A(_0197_),
    .X(net1691));
 sg13g2_dlygate4sd3_1 hold638 (.A(\vga_tetris.tetrisLogic.shapeDropTimerQ[3] ),
    .X(net1692));
 sg13g2_dlygate4sd3_1 hold639 (.A(_1885_),
    .X(net1693));
 sg13g2_dlygate4sd3_1 hold640 (.A(_0047_),
    .X(net1694));
 sg13g2_dlygate4sd3_1 hold641 (.A(\vga_tetris.inputs.buttonTimerQ_0[7] ),
    .X(net1695));
 sg13g2_dlygate4sd3_1 hold642 (.A(_2364_),
    .X(net1696));
 sg13g2_dlygate4sd3_1 hold643 (.A(\vga_tetris.msTimer.msTimerQ[6] ),
    .X(net1697));
 sg13g2_dlygate4sd3_1 hold644 (.A(\vga_tetris.msTimer.msTimerQ[8] ),
    .X(net1698));
 sg13g2_dlygate4sd3_1 hold645 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[0] ),
    .X(net1699));
 sg13g2_dlygate4sd3_1 hold646 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[9] ),
    .X(net1700));
 sg13g2_dlygate4sd3_1 hold647 (.A(\vga_tetris.tetrisLogic.shapeDropTimerQ[2] ),
    .X(net1701));
 sg13g2_dlygate4sd3_1 hold648 (.A(_1883_),
    .X(net1702));
 sg13g2_dlygate4sd3_1 hold649 (.A(\vga_tetris._vgaController_io_pixelPosY[7] ),
    .X(net1703));
 sg13g2_dlygate4sd3_1 hold650 (.A(_0620_),
    .X(net1704));
 sg13g2_dlygate4sd3_1 hold651 (.A(\vga_tetris.inputs.buttonTimerQ_0[1] ),
    .X(net1705));
 sg13g2_dlygate4sd3_1 hold652 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[4] ),
    .X(net1706));
 sg13g2_dlygate4sd3_1 hold653 (.A(\vga_tetris.msTimer.msTimerQ[1] ),
    .X(net1707));
 sg13g2_dlygate4sd3_1 hold654 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[16] ),
    .X(net1708));
 sg13g2_dlygate4sd3_1 hold655 (.A(\vga_tetris.tetrisLogic.shapeDropTimerQ[0] ),
    .X(net1709));
 sg13g2_dlygate4sd3_1 hold656 (.A(_1880_),
    .X(net1710));
 sg13g2_dlygate4sd3_1 hold657 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_rowIndex[0] ),
    .X(net1711));
 sg13g2_dlygate4sd3_1 hold658 (.A(_0070_),
    .X(net1712));
 sg13g2_dlygate4sd3_1 hold659 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[17] ),
    .X(net1713));
 sg13g2_dlygate4sd3_1 hold660 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[19] ),
    .X(net1714));
 sg13g2_dlygate4sd3_1 hold661 (.A(\vga_tetris.inputs.buttonTimerQ_1[1] ),
    .X(net1715));
 sg13g2_dlygate4sd3_1 hold662 (.A(_2373_),
    .X(net1716));
 sg13g2_dlygate4sd3_1 hold663 (.A(_0184_),
    .X(net1717));
 sg13g2_dlygate4sd3_1 hold664 (.A(\vga_tetris.tetrisLogic.shapeDropTimerQ[4] ),
    .X(net1718));
 sg13g2_dlygate4sd3_1 hold665 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[2] ),
    .X(net1719));
 sg13g2_dlygate4sd3_1 hold666 (.A(\vga_tetris.tetrisLogic.gameOverResetHappenedQ ),
    .X(net1720));
 sg13g2_dlygate4sd3_1 hold667 (.A(_0091_),
    .X(net1721));
 sg13g2_dlygate4sd3_1 hold668 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.boardRowDataQ[7] ),
    .X(net1722));
 sg13g2_dlygate4sd3_1 hold669 (.A(\vga_tetris._vgaController_io_pixelPosX[0] ),
    .X(net1723));
 sg13g2_dlygate4sd3_1 hold670 (.A(\vga_tetris._vgaController_io_pixelPosX[7] ),
    .X(net1724));
 sg13g2_dlygate4sd3_1 hold671 (.A(_2903_),
    .X(net1725));
 sg13g2_dlygate4sd3_1 hold672 (.A(\vga_tetris.startTetrisLogicQ ),
    .X(net1726));
 sg13g2_dlygate4sd3_1 hold673 (.A(_0067_),
    .X(net1727));
 sg13g2_dlygate4sd3_1 hold674 (.A(\vga_tetris.vgaController.verticalCounterQ[6] ),
    .X(net1728));
 sg13g2_dlygate4sd3_1 hold675 (.A(_2879_),
    .X(net1729));
 sg13g2_dlygate4sd3_1 hold676 (.A(\vga_tetris.msTimer.msTimerQ[12] ),
    .X(net1730));
 sg13g2_dlygate4sd3_1 hold677 (.A(_1806_),
    .X(net1731));
 sg13g2_dlygate4sd3_1 hold678 (.A(_0027_),
    .X(net1732));
 sg13g2_dlygate4sd3_1 hold679 (.A(\vga_tetris.msTimer.msTimerQ[10] ),
    .X(net1733));
 sg13g2_dlygate4sd3_1 hold680 (.A(_1802_),
    .X(net1734));
 sg13g2_dlygate4sd3_1 hold681 (.A(_0025_),
    .X(net1735));
 sg13g2_dlygate4sd3_1 hold682 (.A(\vga_tetris.tetrisLogic.shapeDataProvider.io_shapeSelector[2] ),
    .X(net1736));
 sg13g2_dlygate4sd3_1 hold683 (.A(_1841_),
    .X(net1737));
 sg13g2_dlygate4sd3_1 hold684 (.A(\vga_tetris.tetrisLogic.shapeDropTimerQ[5] ),
    .X(net1738));
 sg13g2_dlygate4sd3_1 hold685 (.A(\vga_tetris.tetrisLogic.stateQ[1] ),
    .X(net1739));
 sg13g2_dlygate4sd3_1 hold686 (.A(\vga_tetris._tetrisLogic_io_score_3[2] ),
    .X(net1740));
 sg13g2_dlygate4sd3_1 hold687 (.A(_2214_),
    .X(net1741));
 sg13g2_dlygate4sd3_1 hold688 (.A(_0137_),
    .X(net1742));
 sg13g2_dlygate4sd3_1 hold689 (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[3] ),
    .X(net1743));
 sg13g2_dlygate4sd3_1 hold690 (.A(\vga_tetris.msTimer.msTimerQ[9] ),
    .X(net1744));
 sg13g2_dlygate4sd3_1 hold691 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[3] ),
    .X(net1745));
 sg13g2_dlygate4sd3_1 hold692 (.A(_2127_),
    .X(net1746));
 sg13g2_dlygate4sd3_1 hold693 (.A(_0105_),
    .X(net1747));
 sg13g2_dlygate4sd3_1 hold694 (.A(\vga_tetris.inputs.buttonTimerQ_2[5] ),
    .X(net1748));
 sg13g2_dlygate4sd3_1 hold695 (.A(_2404_),
    .X(net1749));
 sg13g2_dlygate4sd3_1 hold696 (.A(_0196_),
    .X(net1750));
 sg13g2_dlygate4sd3_1 hold697 (.A(\vga_tetris.vgaController.horizontalCounterQ[9] ),
    .X(net1751));
 sg13g2_dlygate4sd3_1 hold698 (.A(_1775_),
    .X(net1752));
 sg13g2_dlygate4sd3_1 hold699 (.A(\vga_tetris._tetrisLogic_io_score_0[3] ),
    .X(net1753));
 sg13g2_dlygate4sd3_1 hold700 (.A(_2246_),
    .X(net1754));
 sg13g2_dlygate4sd3_1 hold701 (.A(_0152_),
    .X(net1755));
 sg13g2_dlygate4sd3_1 hold702 (.A(\vga_tetris._tetrisLogic_io_score_0[2] ),
    .X(net1756));
 sg13g2_dlygate4sd3_1 hold703 (.A(_2244_),
    .X(net1757));
 sg13g2_dlygate4sd3_1 hold704 (.A(_0153_),
    .X(net1758));
 sg13g2_dlygate4sd3_1 hold705 (.A(\vga_tetris._tetrisLogic_io_score_1[3] ),
    .X(net1759));
 sg13g2_dlygate4sd3_1 hold706 (.A(_0149_),
    .X(net1760));
 sg13g2_dlygate4sd3_1 hold707 (.A(\vga_tetris.tetrisLogic.stateQ[2] ),
    .X(net1761));
 sg13g2_dlygate4sd3_1 hold708 (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[4] ),
    .X(net1762));
 sg13g2_dlygate4sd3_1 hold709 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[2] ),
    .X(net1763));
 sg13g2_dlygate4sd3_1 hold710 (.A(_2124_),
    .X(net1764));
 sg13g2_dlygate4sd3_1 hold711 (.A(_0104_),
    .X(net1765));
 sg13g2_dlygate4sd3_1 hold712 (.A(\vga_tetris.vgaController.horizontalCounterQ[8] ),
    .X(net1766));
 sg13g2_dlygate4sd3_1 hold713 (.A(\vga_tetris.inputs.buttonTimerQ_3[7] ),
    .X(net1767));
 sg13g2_dlygate4sd3_1 hold714 (.A(_2433_),
    .X(net1768));
 sg13g2_dlygate4sd3_1 hold715 (.A(_2434_),
    .X(net1769));
 sg13g2_dlygate4sd3_1 hold716 (.A(\vga_tetris.inputs.buttonTimerQ_3[0] ),
    .X(net1770));
 sg13g2_dlygate4sd3_1 hold717 (.A(\vga_tetris.runningTetrisLogicQ ),
    .X(net1771));
 sg13g2_dlygate4sd3_1 hold718 (.A(_0211_),
    .X(net1772));
 sg13g2_dlygate4sd3_1 hold719 (.A(\vga_tetris.inputs.buttonTimerQ_3[3] ),
    .X(net1773));
 sg13g2_dlygate4sd3_1 hold720 (.A(_2421_),
    .X(net1774));
 sg13g2_dlygate4sd3_1 hold721 (.A(\vga_tetris.vgaController.verticalCounterQ[5] ),
    .X(net1775));
 sg13g2_dlygate4sd3_1 hold722 (.A(\vga_tetris.tetrisLogic.addOrRemoveShape.stateQ[0] ),
    .X(net1776));
 sg13g2_dlygate4sd3_1 hold723 (.A(_1918_),
    .X(net1777));
 sg13g2_dlygate4sd3_1 hold724 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[16] ),
    .X(net1778));
 sg13g2_dlygate4sd3_1 hold725 (.A(\vga_tetris._vgaController_io_pixelPosY[1] ),
    .X(net1779));
 sg13g2_dlygate4sd3_1 hold726 (.A(\vga_tetris.msTimer.msTimerQ[11] ),
    .X(net1780));
 sg13g2_dlygate4sd3_1 hold727 (.A(\vga_tetris.vgaController.horizontalCounterQ[4] ),
    .X(net1781));
 sg13g2_dlygate4sd3_1 hold728 (.A(\vga_tetris._vgaController_io_pixelPosX[3] ),
    .X(net1782));
 sg13g2_dlygate4sd3_1 hold729 (.A(_0606_),
    .X(net1783));
 sg13g2_dlygate4sd3_1 hold730 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[17] ),
    .X(net1784));
 sg13g2_dlygate4sd3_1 hold731 (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[2] ),
    .X(net1785));
 sg13g2_dlygate4sd3_1 hold732 (.A(\vga_tetris.inputs.buttonTimerQ_0[4] ),
    .X(net1786));
 sg13g2_dlygate4sd3_1 hold733 (.A(_2357_),
    .X(net1787));
 sg13g2_dlygate4sd3_1 hold734 (.A(_0179_),
    .X(net1788));
 sg13g2_dlygate4sd3_1 hold735 (.A(\vga_tetris._tetrisLogic_io_score_1[1] ),
    .X(net1789));
 sg13g2_dlygate4sd3_1 hold736 (.A(\vga_tetris.tetrisLogic.gameOverLogic.buttonPressesCounterQ[1] ),
    .X(net1790));
 sg13g2_dlygate4sd3_1 hold737 (.A(_2221_),
    .X(net1791));
 sg13g2_dlygate4sd3_1 hold738 (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[1] ),
    .X(net1792));
 sg13g2_dlygate4sd3_1 hold739 (.A(\vga_tetris._vgaController_io_pixelPosY[6] ),
    .X(net1793));
 sg13g2_dlygate4sd3_1 hold740 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_done ),
    .X(net1794));
 sg13g2_dlygate4sd3_1 hold741 (.A(_2033_),
    .X(net1795));
 sg13g2_dlygate4sd3_1 hold742 (.A(\vga_tetris.inputs.buttonTimerQ_1[4] ),
    .X(net1796));
 sg13g2_dlygate4sd3_1 hold743 (.A(_2379_),
    .X(net1797));
 sg13g2_dlygate4sd3_1 hold744 (.A(_2381_),
    .X(net1798));
 sg13g2_dlygate4sd3_1 hold745 (.A(\vga_tetris.inputs.buttonTimerQ_2[4] ),
    .X(net1799));
 sg13g2_dlygate4sd3_1 hold746 (.A(_2401_),
    .X(net1800));
 sg13g2_dlygate4sd3_1 hold747 (.A(_2403_),
    .X(net1801));
 sg13g2_dlygate4sd3_1 hold748 (.A(\vga_tetris.inputs.buttonTimerQ_1[2] ),
    .X(net1802));
 sg13g2_dlygate4sd3_1 hold749 (.A(_2376_),
    .X(net1803));
 sg13g2_dlygate4sd3_1 hold750 (.A(\vga_tetris._tetrisLogic_io_score_2[3] ),
    .X(net1804));
 sg13g2_dlygate4sd3_1 hold751 (.A(_2225_),
    .X(net1805));
 sg13g2_dlygate4sd3_1 hold752 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[4] ),
    .X(net1806));
 sg13g2_dlygate4sd3_1 hold753 (.A(_2130_),
    .X(net1807));
 sg13g2_dlygate4sd3_1 hold754 (.A(_0106_),
    .X(net1808));
 sg13g2_dlygate4sd3_1 hold755 (.A(\vga_tetris.vgaController.verticalCounterQ[7] ),
    .X(net1809));
 sg13g2_dlygate4sd3_1 hold756 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[0] ),
    .X(net1810));
 sg13g2_dlygate4sd3_1 hold757 (.A(_2059_),
    .X(net1811));
 sg13g2_dlygate4sd3_1 hold758 (.A(_0097_),
    .X(net1812));
 sg13g2_dlygate4sd3_1 hold759 (.A(\vga_tetris._tetrisLogic_io_score_2[0] ),
    .X(net1813));
 sg13g2_dlygate4sd3_1 hold760 (.A(\vga_tetris.inputs.buttonTimerQ_1[3] ),
    .X(net1814));
 sg13g2_dlygate4sd3_1 hold761 (.A(_2378_),
    .X(net1815));
 sg13g2_dlygate4sd3_1 hold762 (.A(\vga_tetris._tetrisLogic_io_score_1[0] ),
    .X(net1816));
 sg13g2_dlygate4sd3_1 hold763 (.A(_0146_),
    .X(net1817));
 sg13g2_dlygate4sd3_1 hold764 (.A(\vga_tetris.inputs.buttonTimerQ_0[5] ),
    .X(net1818));
 sg13g2_dlygate4sd3_1 hold765 (.A(_2360_),
    .X(net1819));
 sg13g2_dlygate4sd3_1 hold766 (.A(\vga_tetris._tetrisLogic_io_score_0[0] ),
    .X(net1820));
 sg13g2_dlygate4sd3_1 hold767 (.A(_2239_),
    .X(net1821));
 sg13g2_dlygate4sd3_1 hold768 (.A(_0150_),
    .X(net1822));
 sg13g2_dlygate4sd3_1 hold769 (.A(\vga_tetris.inputs.buttonTimerQ_2[3] ),
    .X(net1823));
 sg13g2_dlygate4sd3_1 hold770 (.A(_2400_),
    .X(net1824));
 sg13g2_dlygate4sd3_1 hold771 (.A(\vga_tetris._tetrisLogic_io_score_0[1] ),
    .X(net1825));
 sg13g2_dlygate4sd3_1 hold772 (.A(\vga_tetris.vgaController.verticalCounterQ[9] ),
    .X(net1826));
 sg13g2_dlygate4sd3_1 hold773 (.A(_2884_),
    .X(net1827));
 sg13g2_dlygate4sd3_1 hold774 (.A(\vga_tetris.inputs.buttonTimerQ_3[4] ),
    .X(net1828));
 sg13g2_dlygate4sd3_1 hold775 (.A(\vga_tetris.inputs.buttonTimerQ_3[6] ),
    .X(net1829));
 sg13g2_dlygate4sd3_1 hold776 (.A(_2430_),
    .X(net1830));
 sg13g2_dlygate4sd3_1 hold777 (.A(\vga_tetris.inputs.buttonTimerQ_2[2] ),
    .X(net1831));
 sg13g2_dlygate4sd3_1 hold778 (.A(_2398_),
    .X(net1832));
 sg13g2_dlygate4sd3_1 hold779 (.A(\vga_tetris._inputs_io_leftButtonActive ),
    .X(net1833));
 sg13g2_dlygate4sd3_1 hold780 (.A(_2442_),
    .X(net1834));
 sg13g2_dlygate4sd3_1 hold781 (.A(_0208_),
    .X(net1835));
 sg13g2_dlygate4sd3_1 hold782 (.A(\vga_tetris.inputs.buttonTimerQ_0[2] ),
    .X(net1836));
 sg13g2_dlygate4sd3_1 hold783 (.A(\vga_tetris.inputs.buttonTimerQ_1[5] ),
    .X(net1837));
 sg13g2_dlygate4sd3_1 hold784 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[4] ),
    .X(net1838));
 sg13g2_dlygate4sd3_1 hold785 (.A(_2088_),
    .X(net1839));
 sg13g2_dlygate4sd3_1 hold786 (.A(_0101_),
    .X(net1840));
 sg13g2_dlygate4sd3_1 hold787 (.A(\vga_tetris.inputs.buttonTimerQ_3[5] ),
    .X(net1841));
 sg13g2_dlygate4sd3_1 hold788 (.A(\vga_tetris.inputs.buttonTimerQ_0[3] ),
    .X(net1842));
 sg13g2_dlygate4sd3_1 hold789 (.A(\vga_tetris._inputs_io_rightButtonActive ),
    .X(net1843));
 sg13g2_dlygate4sd3_1 hold790 (.A(\vga_tetris.inputs.buttonTimerQ_3[2] ),
    .X(net1844));
 sg13g2_dlygate4sd3_1 hold791 (.A(_2417_),
    .X(net1845));
 sg13g2_dlygate4sd3_1 hold792 (.A(\vga_tetris._tetrisLogic_io_score_3[1] ),
    .X(net1846));
 sg13g2_dlygate4sd3_1 hold793 (.A(\vga_tetris.inputs.buttonTimerQ_3[1] ),
    .X(net1847));
 sg13g2_dlygate4sd3_1 hold794 (.A(\vga_tetris._inputs_io_rotateButtonActive ),
    .X(net1848));
 sg13g2_dlygate4sd3_1 hold795 (.A(\vga_tetris._tetrisLogic_io_gameOver ),
    .X(net1849));
 sg13g2_dlygate4sd3_1 hold796 (.A(_0154_),
    .X(net1850));
 sg13g2_dlygate4sd3_1 hold797 (.A(\vga_tetris.tetrisLogic.rotationQ[1] ),
    .X(net1851));
 sg13g2_dlygate4sd3_1 hold798 (.A(_1853_),
    .X(net1852));
 sg13g2_dlygate4sd3_1 hold799 (.A(\vga_tetris.vgaController.verticalCounterQ[6] ),
    .X(net1853));
 sg13g2_dlygate4sd3_1 hold800 (.A(\vga_tetris.tetrisLogic.stateQ[4] ),
    .X(net1854));
 sg13g2_dlygate4sd3_1 hold801 (.A(_0041_),
    .X(net1855));
 sg13g2_dlygate4sd3_1 hold802 (.A(\vga_tetris._vgaController_io_pixelPosY[3] ),
    .X(net1856));
 sg13g2_dlygate4sd3_1 hold803 (.A(\vga_tetris._vgaController_io_pixelPosX[2] ),
    .X(net1857));
 sg13g2_dlygate4sd3_1 hold804 (.A(\vga_tetris._vgaController_io_pixelPosX[5] ),
    .X(net1858));
 sg13g2_dlygate4sd3_1 hold805 (.A(_2898_),
    .X(net1859));
 sg13g2_dlygate4sd3_1 hold806 (.A(_0608_),
    .X(net1860));
 sg13g2_dlygate4sd3_1 hold807 (.A(\vga_tetris._vgaController_io_pixelPosY[2] ),
    .X(net1861));
 sg13g2_dlygate4sd3_1 hold808 (.A(_2920_),
    .X(net1862));
 sg13g2_dlygate4sd3_1 hold809 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.operationIsRunningQ ),
    .X(net1863));
 sg13g2_dlygate4sd3_1 hold810 (.A(_2037_),
    .X(net1864));
 sg13g2_dlygate4sd3_1 hold811 (.A(_0096_),
    .X(net1865));
 sg13g2_dlygate4sd3_1 hold812 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.linesToShiftQ[0] ),
    .X(net1866));
 sg13g2_dlygate4sd3_1 hold813 (.A(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[2] ),
    .X(net1867));
 sg13g2_dlygate4sd3_1 hold814 (.A(_1729_),
    .X(net1868));
 sg13g2_dlygate4sd3_1 hold815 (.A(_0003_),
    .X(net1869));
 sg13g2_dlygate4sd3_1 hold816 (.A(\vga_tetris._tetrisLogic_io_score_2[1] ),
    .X(net1870));
 sg13g2_dlygate4sd3_1 hold817 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[1] ),
    .X(net1871));
 sg13g2_dlygate4sd3_1 hold818 (.A(_2067_),
    .X(net1872));
 sg13g2_dlygate4sd3_1 hold819 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[1] ),
    .X(net1873));
 sg13g2_dlygate4sd3_1 hold820 (.A(_2107_),
    .X(net1874));
 sg13g2_dlygate4sd3_1 hold821 (.A(\vga_tetris.tetrisLogic.rotationQ[0] ),
    .X(net1875));
 sg13g2_dlygate4sd3_1 hold822 (.A(_1849_),
    .X(net1876));
 sg13g2_dlygate4sd3_1 hold823 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[0] ),
    .X(net1877));
 sg13g2_dlygate4sd3_1 hold824 (.A(_0102_),
    .X(net1878));
 sg13g2_dlygate4sd3_1 hold825 (.A(\vga_tetris.tetrisLogic.stateQ[0] ),
    .X(net1879));
 sg13g2_dlygate4sd3_1 hold826 (.A(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[0] ),
    .X(net1880));
 sg13g2_dlygate4sd3_1 hold827 (.A(\vga_tetris._vgaController_io_pixelPosX[4] ),
    .X(net1881));
 sg13g2_dlygate4sd3_1 hold828 (.A(_2895_),
    .X(net1882));
 sg13g2_dlygate4sd3_1 hold829 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[3] ),
    .X(net1883));
 sg13g2_dlygate4sd3_1 hold830 (.A(\vga_tetris.tetrisLogic.addOrRemoveShape.io_shapeXCoord[3] ),
    .X(net1884));
 sg13g2_dlygate4sd3_1 hold831 (.A(_1747_),
    .X(net1885));
 sg13g2_dlygate4sd3_1 hold832 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.rowIndexQ[1] ),
    .X(net1886));
 sg13g2_dlygate4sd3_1 hold833 (.A(\vga_tetris._vgaController_io_pixelPosX[9] ),
    .X(net1887));
 sg13g2_dlygate4sd3_1 hold834 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.shiftStartPosQ[2] ),
    .X(net1888));
 sg13g2_dlygate4sd3_1 hold835 (.A(\vga_tetris._tetrisDisplay_io_boardYCoord[1] ),
    .X(net1889));
 sg13g2_dlygate4sd3_1 hold836 (.A(\vga_tetris._vgaController_io_pixelPosX[6] ),
    .X(net1890));
 sg13g2_dlygate4sd3_1 hold837 (.A(_2899_),
    .X(net1891));
 sg13g2_dlygate4sd3_1 hold838 (.A(\vga_tetris._vgaController_io_pixelPosY[0] ),
    .X(net1892));
 sg13g2_dlygate4sd3_1 hold839 (.A(_2924_),
    .X(net1893));
 sg13g2_dlygate4sd3_1 hold840 (.A(\vga_tetris.tetrisLogic.shiftTheBoard.stateQ[0] ),
    .X(net1894));
 sg13g2_dlygate4sd3_1 hold841 (.A(\vga_tetris.inputs.buttonTimerQ_3[1] ),
    .X(net1895));
 sg13g2_dlygate4sd3_1 hold842 (.A(_2419_),
    .X(net1896));
 sg13g2_dlygate4sd3_1 hold843 (.A(\vga_tetris.vgaController.horizontalCounterQ[5] ),
    .X(net1897));
 sg13g2_dlygate4sd3_1 hold844 (.A(_1751_),
    .X(net1898));
 sg13g2_dlygate4sd3_1 hold845 (.A(\vga_tetris.tetrisLogic.shapeDropTimerQ[0] ),
    .X(net1899));
 sg13g2_dlygate4sd3_1 hold846 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[14] ),
    .X(net1900));
 sg13g2_dlygate4sd3_1 hold847 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_done ),
    .X(net1901));
 sg13g2_dlygate4sd3_1 hold848 (.A(\vga_tetris.tetrisLogic._addOrRemoveShape_io_boardRowDataOut[15] ),
    .X(net1902));
 sg13g2_dlygate4sd3_1 hold849 (.A(_2318_),
    .X(net1903));
 sg13g2_dlygate4sd3_1 hold850 (.A(\vga_tetris.tetrisLogic.adderSubtracter.io_a[2] ),
    .X(net1904));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_4 FILLER_4_546 ();
 sg13g2_fill_2 FILLER_4_550 ();
 sg13g2_decap_8 FILLER_4_556 ();
 sg13g2_decap_8 FILLER_4_563 ();
 sg13g2_decap_8 FILLER_4_570 ();
 sg13g2_decap_8 FILLER_4_577 ();
 sg13g2_decap_8 FILLER_4_584 ();
 sg13g2_decap_8 FILLER_4_591 ();
 sg13g2_decap_8 FILLER_4_598 ();
 sg13g2_decap_8 FILLER_4_605 ();
 sg13g2_decap_8 FILLER_4_612 ();
 sg13g2_decap_8 FILLER_4_619 ();
 sg13g2_decap_8 FILLER_4_626 ();
 sg13g2_decap_8 FILLER_4_633 ();
 sg13g2_decap_8 FILLER_4_640 ();
 sg13g2_decap_8 FILLER_4_647 ();
 sg13g2_decap_8 FILLER_4_654 ();
 sg13g2_decap_8 FILLER_4_661 ();
 sg13g2_decap_8 FILLER_4_668 ();
 sg13g2_decap_8 FILLER_4_675 ();
 sg13g2_decap_8 FILLER_4_682 ();
 sg13g2_decap_8 FILLER_4_689 ();
 sg13g2_decap_8 FILLER_4_696 ();
 sg13g2_decap_8 FILLER_4_703 ();
 sg13g2_decap_8 FILLER_4_710 ();
 sg13g2_decap_8 FILLER_4_717 ();
 sg13g2_decap_8 FILLER_4_724 ();
 sg13g2_decap_8 FILLER_4_731 ();
 sg13g2_decap_8 FILLER_4_738 ();
 sg13g2_decap_8 FILLER_4_745 ();
 sg13g2_decap_8 FILLER_4_752 ();
 sg13g2_decap_8 FILLER_4_759 ();
 sg13g2_decap_8 FILLER_4_766 ();
 sg13g2_decap_8 FILLER_4_773 ();
 sg13g2_decap_8 FILLER_4_780 ();
 sg13g2_decap_8 FILLER_4_787 ();
 sg13g2_decap_8 FILLER_4_794 ();
 sg13g2_decap_8 FILLER_4_801 ();
 sg13g2_decap_8 FILLER_4_808 ();
 sg13g2_decap_8 FILLER_4_815 ();
 sg13g2_decap_8 FILLER_4_822 ();
 sg13g2_decap_8 FILLER_4_829 ();
 sg13g2_decap_8 FILLER_4_836 ();
 sg13g2_decap_8 FILLER_4_843 ();
 sg13g2_decap_8 FILLER_4_850 ();
 sg13g2_decap_4 FILLER_4_857 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_fill_2 FILLER_5_490 ();
 sg13g2_fill_2 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_503 ();
 sg13g2_decap_8 FILLER_5_510 ();
 sg13g2_decap_8 FILLER_5_517 ();
 sg13g2_decap_8 FILLER_5_524 ();
 sg13g2_decap_8 FILLER_5_531 ();
 sg13g2_decap_4 FILLER_5_538 ();
 sg13g2_decap_8 FILLER_5_569 ();
 sg13g2_decap_8 FILLER_5_576 ();
 sg13g2_decap_8 FILLER_5_583 ();
 sg13g2_decap_8 FILLER_5_590 ();
 sg13g2_decap_8 FILLER_5_597 ();
 sg13g2_decap_8 FILLER_5_604 ();
 sg13g2_decap_8 FILLER_5_611 ();
 sg13g2_decap_8 FILLER_5_618 ();
 sg13g2_decap_8 FILLER_5_625 ();
 sg13g2_decap_8 FILLER_5_632 ();
 sg13g2_decap_8 FILLER_5_639 ();
 sg13g2_decap_8 FILLER_5_646 ();
 sg13g2_decap_8 FILLER_5_653 ();
 sg13g2_decap_8 FILLER_5_660 ();
 sg13g2_decap_8 FILLER_5_667 ();
 sg13g2_decap_8 FILLER_5_674 ();
 sg13g2_decap_8 FILLER_5_681 ();
 sg13g2_decap_8 FILLER_5_688 ();
 sg13g2_decap_8 FILLER_5_695 ();
 sg13g2_decap_8 FILLER_5_702 ();
 sg13g2_decap_8 FILLER_5_709 ();
 sg13g2_decap_8 FILLER_5_716 ();
 sg13g2_decap_8 FILLER_5_723 ();
 sg13g2_decap_8 FILLER_5_730 ();
 sg13g2_decap_8 FILLER_5_737 ();
 sg13g2_decap_8 FILLER_5_744 ();
 sg13g2_decap_8 FILLER_5_751 ();
 sg13g2_decap_8 FILLER_5_758 ();
 sg13g2_decap_8 FILLER_5_765 ();
 sg13g2_decap_8 FILLER_5_772 ();
 sg13g2_decap_8 FILLER_5_779 ();
 sg13g2_decap_8 FILLER_5_786 ();
 sg13g2_decap_8 FILLER_5_793 ();
 sg13g2_decap_8 FILLER_5_800 ();
 sg13g2_decap_8 FILLER_5_807 ();
 sg13g2_decap_8 FILLER_5_814 ();
 sg13g2_decap_8 FILLER_5_821 ();
 sg13g2_decap_8 FILLER_5_828 ();
 sg13g2_decap_8 FILLER_5_835 ();
 sg13g2_decap_8 FILLER_5_842 ();
 sg13g2_decap_8 FILLER_5_849 ();
 sg13g2_decap_4 FILLER_5_856 ();
 sg13g2_fill_2 FILLER_5_860 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_fill_1 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_278 ();
 sg13g2_decap_8 FILLER_6_285 ();
 sg13g2_decap_8 FILLER_6_292 ();
 sg13g2_decap_8 FILLER_6_299 ();
 sg13g2_decap_8 FILLER_6_306 ();
 sg13g2_fill_2 FILLER_6_313 ();
 sg13g2_decap_8 FILLER_6_319 ();
 sg13g2_decap_8 FILLER_6_326 ();
 sg13g2_decap_4 FILLER_6_333 ();
 sg13g2_decap_8 FILLER_6_342 ();
 sg13g2_decap_8 FILLER_6_349 ();
 sg13g2_decap_8 FILLER_6_356 ();
 sg13g2_decap_8 FILLER_6_363 ();
 sg13g2_decap_8 FILLER_6_370 ();
 sg13g2_fill_2 FILLER_6_377 ();
 sg13g2_decap_8 FILLER_6_388 ();
 sg13g2_fill_1 FILLER_6_404 ();
 sg13g2_decap_8 FILLER_6_414 ();
 sg13g2_decap_4 FILLER_6_421 ();
 sg13g2_fill_1 FILLER_6_452 ();
 sg13g2_decap_8 FILLER_6_457 ();
 sg13g2_fill_2 FILLER_6_464 ();
 sg13g2_decap_8 FILLER_6_475 ();
 sg13g2_decap_4 FILLER_6_482 ();
 sg13g2_fill_1 FILLER_6_486 ();
 sg13g2_decap_8 FILLER_6_523 ();
 sg13g2_decap_8 FILLER_6_530 ();
 sg13g2_fill_2 FILLER_6_537 ();
 sg13g2_fill_2 FILLER_6_552 ();
 sg13g2_fill_1 FILLER_6_554 ();
 sg13g2_fill_2 FILLER_6_559 ();
 sg13g2_fill_1 FILLER_6_561 ();
 sg13g2_fill_2 FILLER_6_571 ();
 sg13g2_fill_1 FILLER_6_577 ();
 sg13g2_fill_2 FILLER_6_587 ();
 sg13g2_fill_1 FILLER_6_589 ();
 sg13g2_fill_2 FILLER_6_608 ();
 sg13g2_fill_1 FILLER_6_610 ();
 sg13g2_decap_4 FILLER_6_615 ();
 sg13g2_fill_2 FILLER_6_619 ();
 sg13g2_fill_1 FILLER_6_648 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_683 ();
 sg13g2_decap_8 FILLER_6_690 ();
 sg13g2_decap_8 FILLER_6_697 ();
 sg13g2_decap_8 FILLER_6_704 ();
 sg13g2_decap_8 FILLER_6_711 ();
 sg13g2_decap_8 FILLER_6_718 ();
 sg13g2_decap_8 FILLER_6_725 ();
 sg13g2_decap_8 FILLER_6_732 ();
 sg13g2_decap_8 FILLER_6_739 ();
 sg13g2_decap_8 FILLER_6_746 ();
 sg13g2_decap_8 FILLER_6_753 ();
 sg13g2_decap_8 FILLER_6_760 ();
 sg13g2_decap_8 FILLER_6_767 ();
 sg13g2_decap_8 FILLER_6_774 ();
 sg13g2_decap_8 FILLER_6_781 ();
 sg13g2_decap_8 FILLER_6_788 ();
 sg13g2_decap_8 FILLER_6_795 ();
 sg13g2_decap_8 FILLER_6_802 ();
 sg13g2_decap_8 FILLER_6_809 ();
 sg13g2_decap_8 FILLER_6_816 ();
 sg13g2_decap_8 FILLER_6_823 ();
 sg13g2_decap_8 FILLER_6_830 ();
 sg13g2_decap_8 FILLER_6_837 ();
 sg13g2_decap_8 FILLER_6_844 ();
 sg13g2_decap_8 FILLER_6_851 ();
 sg13g2_decap_4 FILLER_6_858 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_fill_2 FILLER_7_98 ();
 sg13g2_fill_1 FILLER_7_100 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_fill_2 FILLER_7_161 ();
 sg13g2_fill_2 FILLER_7_167 ();
 sg13g2_fill_1 FILLER_7_169 ();
 sg13g2_decap_8 FILLER_7_174 ();
 sg13g2_decap_8 FILLER_7_181 ();
 sg13g2_decap_8 FILLER_7_188 ();
 sg13g2_fill_2 FILLER_7_195 ();
 sg13g2_fill_1 FILLER_7_197 ();
 sg13g2_decap_8 FILLER_7_206 ();
 sg13g2_decap_8 FILLER_7_213 ();
 sg13g2_decap_8 FILLER_7_220 ();
 sg13g2_decap_8 FILLER_7_227 ();
 sg13g2_decap_8 FILLER_7_234 ();
 sg13g2_decap_8 FILLER_7_241 ();
 sg13g2_decap_8 FILLER_7_248 ();
 sg13g2_decap_8 FILLER_7_255 ();
 sg13g2_decap_8 FILLER_7_262 ();
 sg13g2_decap_4 FILLER_7_300 ();
 sg13g2_fill_1 FILLER_7_304 ();
 sg13g2_fill_1 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_fill_1 FILLER_7_371 ();
 sg13g2_fill_2 FILLER_7_403 ();
 sg13g2_fill_2 FILLER_7_477 ();
 sg13g2_fill_1 FILLER_7_479 ();
 sg13g2_decap_4 FILLER_7_485 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_fill_2 FILLER_7_504 ();
 sg13g2_fill_1 FILLER_7_533 ();
 sg13g2_fill_2 FILLER_7_566 ();
 sg13g2_fill_1 FILLER_7_671 ();
 sg13g2_decap_8 FILLER_7_699 ();
 sg13g2_decap_8 FILLER_7_706 ();
 sg13g2_decap_8 FILLER_7_713 ();
 sg13g2_decap_8 FILLER_7_720 ();
 sg13g2_decap_8 FILLER_7_727 ();
 sg13g2_decap_8 FILLER_7_734 ();
 sg13g2_decap_8 FILLER_7_741 ();
 sg13g2_decap_8 FILLER_7_748 ();
 sg13g2_decap_8 FILLER_7_755 ();
 sg13g2_decap_8 FILLER_7_762 ();
 sg13g2_decap_8 FILLER_7_769 ();
 sg13g2_decap_8 FILLER_7_776 ();
 sg13g2_decap_8 FILLER_7_783 ();
 sg13g2_decap_8 FILLER_7_790 ();
 sg13g2_decap_8 FILLER_7_797 ();
 sg13g2_decap_8 FILLER_7_804 ();
 sg13g2_decap_8 FILLER_7_811 ();
 sg13g2_decap_8 FILLER_7_818 ();
 sg13g2_decap_8 FILLER_7_825 ();
 sg13g2_decap_8 FILLER_7_832 ();
 sg13g2_decap_8 FILLER_7_839 ();
 sg13g2_decap_8 FILLER_7_846 ();
 sg13g2_decap_8 FILLER_7_853 ();
 sg13g2_fill_2 FILLER_7_860 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_4 FILLER_8_63 ();
 sg13g2_decap_4 FILLER_8_71 ();
 sg13g2_decap_8 FILLER_8_80 ();
 sg13g2_decap_8 FILLER_8_87 ();
 sg13g2_fill_2 FILLER_8_94 ();
 sg13g2_fill_2 FILLER_8_123 ();
 sg13g2_decap_8 FILLER_8_129 ();
 sg13g2_fill_1 FILLER_8_136 ();
 sg13g2_decap_8 FILLER_8_146 ();
 sg13g2_decap_4 FILLER_8_153 ();
 sg13g2_fill_1 FILLER_8_157 ();
 sg13g2_fill_2 FILLER_8_185 ();
 sg13g2_fill_2 FILLER_8_268 ();
 sg13g2_fill_1 FILLER_8_270 ();
 sg13g2_fill_2 FILLER_8_289 ();
 sg13g2_fill_1 FILLER_8_291 ();
 sg13g2_fill_2 FILLER_8_305 ();
 sg13g2_fill_2 FILLER_8_317 ();
 sg13g2_fill_1 FILLER_8_323 ();
 sg13g2_fill_2 FILLER_8_342 ();
 sg13g2_fill_1 FILLER_8_344 ();
 sg13g2_fill_1 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_360 ();
 sg13g2_decap_4 FILLER_8_367 ();
 sg13g2_decap_8 FILLER_8_389 ();
 sg13g2_decap_4 FILLER_8_396 ();
 sg13g2_fill_1 FILLER_8_400 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_decap_4 FILLER_8_416 ();
 sg13g2_fill_2 FILLER_8_420 ();
 sg13g2_decap_4 FILLER_8_435 ();
 sg13g2_fill_1 FILLER_8_439 ();
 sg13g2_decap_4 FILLER_8_450 ();
 sg13g2_fill_1 FILLER_8_454 ();
 sg13g2_decap_8 FILLER_8_459 ();
 sg13g2_decap_8 FILLER_8_466 ();
 sg13g2_fill_2 FILLER_8_473 ();
 sg13g2_fill_2 FILLER_8_520 ();
 sg13g2_decap_4 FILLER_8_535 ();
 sg13g2_fill_2 FILLER_8_539 ();
 sg13g2_fill_1 FILLER_8_545 ();
 sg13g2_fill_1 FILLER_8_564 ();
 sg13g2_decap_8 FILLER_8_579 ();
 sg13g2_decap_8 FILLER_8_586 ();
 sg13g2_fill_2 FILLER_8_593 ();
 sg13g2_fill_2 FILLER_8_604 ();
 sg13g2_fill_2 FILLER_8_642 ();
 sg13g2_fill_1 FILLER_8_644 ();
 sg13g2_fill_2 FILLER_8_653 ();
 sg13g2_decap_4 FILLER_8_659 ();
 sg13g2_decap_8 FILLER_8_704 ();
 sg13g2_fill_1 FILLER_8_711 ();
 sg13g2_fill_2 FILLER_8_717 ();
 sg13g2_decap_8 FILLER_8_723 ();
 sg13g2_decap_8 FILLER_8_730 ();
 sg13g2_decap_8 FILLER_8_737 ();
 sg13g2_decap_8 FILLER_8_744 ();
 sg13g2_decap_8 FILLER_8_751 ();
 sg13g2_decap_8 FILLER_8_758 ();
 sg13g2_decap_8 FILLER_8_765 ();
 sg13g2_decap_8 FILLER_8_772 ();
 sg13g2_decap_8 FILLER_8_779 ();
 sg13g2_decap_8 FILLER_8_786 ();
 sg13g2_decap_8 FILLER_8_793 ();
 sg13g2_decap_8 FILLER_8_800 ();
 sg13g2_decap_8 FILLER_8_807 ();
 sg13g2_decap_8 FILLER_8_814 ();
 sg13g2_decap_8 FILLER_8_821 ();
 sg13g2_decap_8 FILLER_8_828 ();
 sg13g2_decap_8 FILLER_8_835 ();
 sg13g2_decap_8 FILLER_8_842 ();
 sg13g2_decap_8 FILLER_8_849 ();
 sg13g2_decap_4 FILLER_8_856 ();
 sg13g2_fill_2 FILLER_8_860 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_4 FILLER_9_35 ();
 sg13g2_fill_1 FILLER_9_70 ();
 sg13g2_decap_4 FILLER_9_98 ();
 sg13g2_fill_1 FILLER_9_102 ();
 sg13g2_fill_2 FILLER_9_108 ();
 sg13g2_fill_2 FILLER_9_214 ();
 sg13g2_fill_2 FILLER_9_229 ();
 sg13g2_fill_1 FILLER_9_231 ();
 sg13g2_fill_2 FILLER_9_241 ();
 sg13g2_fill_1 FILLER_9_243 ();
 sg13g2_fill_2 FILLER_9_270 ();
 sg13g2_fill_1 FILLER_9_272 ();
 sg13g2_fill_2 FILLER_9_314 ();
 sg13g2_fill_1 FILLER_9_316 ();
 sg13g2_fill_1 FILLER_9_371 ();
 sg13g2_decap_4 FILLER_9_458 ();
 sg13g2_fill_2 FILLER_9_462 ();
 sg13g2_fill_2 FILLER_9_469 ();
 sg13g2_fill_1 FILLER_9_475 ();
 sg13g2_decap_4 FILLER_9_485 ();
 sg13g2_fill_1 FILLER_9_489 ();
 sg13g2_decap_4 FILLER_9_495 ();
 sg13g2_fill_1 FILLER_9_514 ();
 sg13g2_fill_2 FILLER_9_520 ();
 sg13g2_decap_4 FILLER_9_581 ();
 sg13g2_fill_2 FILLER_9_671 ();
 sg13g2_fill_1 FILLER_9_673 ();
 sg13g2_fill_2 FILLER_9_731 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_772 ();
 sg13g2_decap_8 FILLER_9_779 ();
 sg13g2_decap_8 FILLER_9_786 ();
 sg13g2_decap_8 FILLER_9_793 ();
 sg13g2_decap_8 FILLER_9_800 ();
 sg13g2_decap_8 FILLER_9_807 ();
 sg13g2_decap_8 FILLER_9_814 ();
 sg13g2_decap_8 FILLER_9_821 ();
 sg13g2_decap_8 FILLER_9_828 ();
 sg13g2_decap_8 FILLER_9_835 ();
 sg13g2_decap_8 FILLER_9_842 ();
 sg13g2_decap_8 FILLER_9_849 ();
 sg13g2_decap_4 FILLER_9_856 ();
 sg13g2_fill_2 FILLER_9_860 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_fill_1 FILLER_10_42 ();
 sg13g2_fill_2 FILLER_10_75 ();
 sg13g2_decap_4 FILLER_10_81 ();
 sg13g2_fill_2 FILLER_10_98 ();
 sg13g2_fill_2 FILLER_10_105 ();
 sg13g2_fill_1 FILLER_10_107 ();
 sg13g2_decap_8 FILLER_10_136 ();
 sg13g2_fill_1 FILLER_10_143 ();
 sg13g2_fill_2 FILLER_10_176 ();
 sg13g2_fill_1 FILLER_10_178 ();
 sg13g2_decap_8 FILLER_10_215 ();
 sg13g2_decap_8 FILLER_10_222 ();
 sg13g2_fill_2 FILLER_10_229 ();
 sg13g2_fill_1 FILLER_10_236 ();
 sg13g2_fill_2 FILLER_10_259 ();
 sg13g2_fill_2 FILLER_10_266 ();
 sg13g2_fill_1 FILLER_10_300 ();
 sg13g2_decap_4 FILLER_10_332 ();
 sg13g2_fill_1 FILLER_10_340 ();
 sg13g2_decap_4 FILLER_10_353 ();
 sg13g2_fill_2 FILLER_10_357 ();
 sg13g2_fill_2 FILLER_10_368 ();
 sg13g2_fill_2 FILLER_10_374 ();
 sg13g2_fill_1 FILLER_10_376 ();
 sg13g2_fill_2 FILLER_10_385 ();
 sg13g2_fill_2 FILLER_10_400 ();
 sg13g2_decap_4 FILLER_10_412 ();
 sg13g2_fill_2 FILLER_10_435 ();
 sg13g2_decap_8 FILLER_10_445 ();
 sg13g2_fill_1 FILLER_10_452 ();
 sg13g2_decap_8 FILLER_10_557 ();
 sg13g2_fill_2 FILLER_10_564 ();
 sg13g2_fill_1 FILLER_10_566 ();
 sg13g2_fill_1 FILLER_10_597 ();
 sg13g2_fill_1 FILLER_10_634 ();
 sg13g2_fill_2 FILLER_10_653 ();
 sg13g2_fill_1 FILLER_10_660 ();
 sg13g2_fill_2 FILLER_10_683 ();
 sg13g2_fill_1 FILLER_10_685 ();
 sg13g2_fill_1 FILLER_10_716 ();
 sg13g2_fill_2 FILLER_10_744 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_fill_2 FILLER_11_21 ();
 sg13g2_decap_4 FILLER_11_28 ();
 sg13g2_fill_2 FILLER_11_36 ();
 sg13g2_fill_1 FILLER_11_38 ();
 sg13g2_fill_1 FILLER_11_80 ();
 sg13g2_decap_8 FILLER_11_134 ();
 sg13g2_decap_4 FILLER_11_141 ();
 sg13g2_fill_1 FILLER_11_199 ();
 sg13g2_decap_8 FILLER_11_213 ();
 sg13g2_fill_2 FILLER_11_251 ();
 sg13g2_fill_2 FILLER_11_307 ();
 sg13g2_fill_1 FILLER_11_309 ();
 sg13g2_decap_4 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_4 FILLER_11_357 ();
 sg13g2_fill_2 FILLER_11_361 ();
 sg13g2_fill_2 FILLER_11_417 ();
 sg13g2_fill_1 FILLER_11_419 ();
 sg13g2_fill_1 FILLER_11_455 ();
 sg13g2_fill_2 FILLER_11_513 ();
 sg13g2_fill_2 FILLER_11_537 ();
 sg13g2_fill_1 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_fill_1 FILLER_11_595 ();
 sg13g2_decap_4 FILLER_11_601 ();
 sg13g2_fill_2 FILLER_11_605 ();
 sg13g2_decap_4 FILLER_11_633 ();
 sg13g2_fill_1 FILLER_11_637 ();
 sg13g2_fill_2 FILLER_11_642 ();
 sg13g2_fill_2 FILLER_11_679 ();
 sg13g2_fill_1 FILLER_11_681 ();
 sg13g2_decap_4 FILLER_11_740 ();
 sg13g2_fill_2 FILLER_11_744 ();
 sg13g2_decap_4 FILLER_11_751 ();
 sg13g2_fill_2 FILLER_11_759 ();
 sg13g2_fill_1 FILLER_11_761 ();
 sg13g2_fill_1 FILLER_11_766 ();
 sg13g2_decap_8 FILLER_11_776 ();
 sg13g2_decap_8 FILLER_11_783 ();
 sg13g2_decap_8 FILLER_11_790 ();
 sg13g2_decap_8 FILLER_11_797 ();
 sg13g2_decap_8 FILLER_11_804 ();
 sg13g2_decap_8 FILLER_11_811 ();
 sg13g2_decap_8 FILLER_11_818 ();
 sg13g2_decap_8 FILLER_11_825 ();
 sg13g2_decap_8 FILLER_11_832 ();
 sg13g2_decap_8 FILLER_11_839 ();
 sg13g2_decap_8 FILLER_11_846 ();
 sg13g2_decap_8 FILLER_11_853 ();
 sg13g2_fill_2 FILLER_11_860 ();
 sg13g2_decap_4 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_4 ();
 sg13g2_fill_2 FILLER_12_41 ();
 sg13g2_fill_1 FILLER_12_43 ();
 sg13g2_decap_8 FILLER_12_48 ();
 sg13g2_decap_8 FILLER_12_55 ();
 sg13g2_fill_1 FILLER_12_75 ();
 sg13g2_fill_1 FILLER_12_93 ();
 sg13g2_fill_2 FILLER_12_115 ();
 sg13g2_decap_4 FILLER_12_175 ();
 sg13g2_fill_1 FILLER_12_228 ();
 sg13g2_decap_8 FILLER_12_233 ();
 sg13g2_fill_1 FILLER_12_240 ();
 sg13g2_decap_4 FILLER_12_255 ();
 sg13g2_decap_4 FILLER_12_280 ();
 sg13g2_decap_4 FILLER_12_297 ();
 sg13g2_fill_1 FILLER_12_310 ();
 sg13g2_fill_1 FILLER_12_319 ();
 sg13g2_fill_2 FILLER_12_338 ();
 sg13g2_fill_1 FILLER_12_340 ();
 sg13g2_fill_2 FILLER_12_368 ();
 sg13g2_fill_1 FILLER_12_370 ();
 sg13g2_fill_2 FILLER_12_389 ();
 sg13g2_fill_1 FILLER_12_428 ();
 sg13g2_decap_4 FILLER_12_485 ();
 sg13g2_fill_1 FILLER_12_489 ();
 sg13g2_decap_8 FILLER_12_503 ();
 sg13g2_fill_2 FILLER_12_510 ();
 sg13g2_decap_4 FILLER_12_516 ();
 sg13g2_fill_2 FILLER_12_520 ();
 sg13g2_decap_8 FILLER_12_535 ();
 sg13g2_decap_8 FILLER_12_542 ();
 sg13g2_decap_4 FILLER_12_549 ();
 sg13g2_fill_1 FILLER_12_553 ();
 sg13g2_fill_2 FILLER_12_558 ();
 sg13g2_fill_1 FILLER_12_560 ();
 sg13g2_fill_1 FILLER_12_575 ();
 sg13g2_fill_2 FILLER_12_580 ();
 sg13g2_fill_1 FILLER_12_582 ();
 sg13g2_fill_2 FILLER_12_610 ();
 sg13g2_decap_4 FILLER_12_656 ();
 sg13g2_fill_1 FILLER_12_660 ();
 sg13g2_decap_4 FILLER_12_674 ();
 sg13g2_fill_1 FILLER_12_682 ();
 sg13g2_fill_2 FILLER_12_710 ();
 sg13g2_fill_1 FILLER_12_712 ();
 sg13g2_fill_2 FILLER_12_745 ();
 sg13g2_fill_1 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_7 ();
 sg13g2_fill_1 FILLER_13_9 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_fill_1 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_27 ();
 sg13g2_decap_4 FILLER_13_43 ();
 sg13g2_fill_2 FILLER_13_47 ();
 sg13g2_fill_2 FILLER_13_62 ();
 sg13g2_fill_2 FILLER_13_69 ();
 sg13g2_fill_1 FILLER_13_71 ();
 sg13g2_fill_1 FILLER_13_117 ();
 sg13g2_fill_2 FILLER_13_132 ();
 sg13g2_fill_1 FILLER_13_134 ();
 sg13g2_decap_8 FILLER_13_157 ();
 sg13g2_decap_4 FILLER_13_164 ();
 sg13g2_decap_8 FILLER_13_187 ();
 sg13g2_decap_4 FILLER_13_194 ();
 sg13g2_fill_1 FILLER_13_198 ();
 sg13g2_fill_2 FILLER_13_204 ();
 sg13g2_fill_1 FILLER_13_206 ();
 sg13g2_decap_4 FILLER_13_220 ();
 sg13g2_fill_2 FILLER_13_264 ();
 sg13g2_fill_1 FILLER_13_266 ();
 sg13g2_fill_2 FILLER_13_294 ();
 sg13g2_fill_2 FILLER_13_332 ();
 sg13g2_fill_1 FILLER_13_347 ();
 sg13g2_fill_2 FILLER_13_393 ();
 sg13g2_fill_2 FILLER_13_439 ();
 sg13g2_fill_1 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_fill_1 FILLER_13_462 ();
 sg13g2_fill_2 FILLER_13_467 ();
 sg13g2_fill_1 FILLER_13_469 ();
 sg13g2_fill_2 FILLER_13_475 ();
 sg13g2_fill_2 FILLER_13_522 ();
 sg13g2_decap_4 FILLER_13_551 ();
 sg13g2_fill_1 FILLER_13_555 ();
 sg13g2_decap_8 FILLER_13_565 ();
 sg13g2_fill_2 FILLER_13_572 ();
 sg13g2_decap_4 FILLER_13_595 ();
 sg13g2_fill_2 FILLER_13_599 ();
 sg13g2_fill_2 FILLER_13_605 ();
 sg13g2_decap_4 FILLER_13_616 ();
 sg13g2_fill_1 FILLER_13_620 ();
 sg13g2_fill_2 FILLER_13_675 ();
 sg13g2_fill_1 FILLER_13_677 ();
 sg13g2_fill_1 FILLER_13_687 ();
 sg13g2_decap_4 FILLER_13_715 ();
 sg13g2_fill_1 FILLER_13_719 ();
 sg13g2_decap_8 FILLER_13_724 ();
 sg13g2_fill_1 FILLER_13_731 ();
 sg13g2_decap_4 FILLER_13_741 ();
 sg13g2_fill_2 FILLER_13_745 ();
 sg13g2_decap_8 FILLER_13_778 ();
 sg13g2_decap_8 FILLER_13_790 ();
 sg13g2_decap_8 FILLER_13_797 ();
 sg13g2_decap_8 FILLER_13_804 ();
 sg13g2_decap_8 FILLER_13_811 ();
 sg13g2_decap_8 FILLER_13_818 ();
 sg13g2_decap_8 FILLER_13_825 ();
 sg13g2_decap_8 FILLER_13_832 ();
 sg13g2_decap_8 FILLER_13_839 ();
 sg13g2_decap_8 FILLER_13_846 ();
 sg13g2_decap_8 FILLER_13_853 ();
 sg13g2_fill_2 FILLER_13_860 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_2 ();
 sg13g2_decap_8 FILLER_14_75 ();
 sg13g2_fill_2 FILLER_14_82 ();
 sg13g2_decap_4 FILLER_14_89 ();
 sg13g2_fill_1 FILLER_14_98 ();
 sg13g2_fill_1 FILLER_14_148 ();
 sg13g2_fill_1 FILLER_14_154 ();
 sg13g2_decap_4 FILLER_14_159 ();
 sg13g2_fill_1 FILLER_14_163 ();
 sg13g2_decap_4 FILLER_14_177 ();
 sg13g2_fill_2 FILLER_14_181 ();
 sg13g2_fill_2 FILLER_14_196 ();
 sg13g2_fill_1 FILLER_14_225 ();
 sg13g2_decap_4 FILLER_14_235 ();
 sg13g2_fill_2 FILLER_14_239 ();
 sg13g2_fill_1 FILLER_14_245 ();
 sg13g2_fill_2 FILLER_14_251 ();
 sg13g2_fill_1 FILLER_14_253 ();
 sg13g2_decap_4 FILLER_14_258 ();
 sg13g2_fill_2 FILLER_14_262 ();
 sg13g2_fill_2 FILLER_14_269 ();
 sg13g2_fill_1 FILLER_14_271 ();
 sg13g2_decap_4 FILLER_14_276 ();
 sg13g2_decap_8 FILLER_14_289 ();
 sg13g2_decap_4 FILLER_14_296 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_4 FILLER_14_315 ();
 sg13g2_fill_1 FILLER_14_319 ();
 sg13g2_fill_1 FILLER_14_338 ();
 sg13g2_fill_2 FILLER_14_382 ();
 sg13g2_decap_4 FILLER_14_437 ();
 sg13g2_decap_8 FILLER_14_486 ();
 sg13g2_fill_2 FILLER_14_493 ();
 sg13g2_fill_1 FILLER_14_495 ();
 sg13g2_fill_1 FILLER_14_512 ();
 sg13g2_fill_1 FILLER_14_527 ();
 sg13g2_fill_2 FILLER_14_591 ();
 sg13g2_fill_1 FILLER_14_593 ();
 sg13g2_fill_2 FILLER_14_603 ();
 sg13g2_fill_1 FILLER_14_605 ();
 sg13g2_fill_2 FILLER_14_663 ();
 sg13g2_fill_1 FILLER_14_665 ();
 sg13g2_fill_1 FILLER_14_693 ();
 sg13g2_decap_8 FILLER_14_698 ();
 sg13g2_decap_4 FILLER_14_705 ();
 sg13g2_fill_1 FILLER_14_709 ();
 sg13g2_fill_2 FILLER_14_742 ();
 sg13g2_fill_1 FILLER_14_744 ();
 sg13g2_fill_1 FILLER_14_762 ();
 sg13g2_fill_1 FILLER_14_785 ();
 sg13g2_decap_8 FILLER_14_813 ();
 sg13g2_decap_8 FILLER_14_824 ();
 sg13g2_decap_8 FILLER_14_831 ();
 sg13g2_decap_8 FILLER_14_838 ();
 sg13g2_decap_8 FILLER_14_845 ();
 sg13g2_decap_8 FILLER_14_852 ();
 sg13g2_fill_2 FILLER_14_859 ();
 sg13g2_fill_1 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_13 ();
 sg13g2_decap_4 FILLER_15_20 ();
 sg13g2_fill_1 FILLER_15_24 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_fill_2 FILLER_15_49 ();
 sg13g2_decap_4 FILLER_15_83 ();
 sg13g2_fill_2 FILLER_15_87 ();
 sg13g2_fill_2 FILLER_15_102 ();
 sg13g2_fill_1 FILLER_15_104 ();
 sg13g2_fill_1 FILLER_15_131 ();
 sg13g2_fill_2 FILLER_15_136 ();
 sg13g2_fill_2 FILLER_15_203 ();
 sg13g2_decap_4 FILLER_15_231 ();
 sg13g2_fill_1 FILLER_15_240 ();
 sg13g2_decap_8 FILLER_15_269 ();
 sg13g2_fill_2 FILLER_15_276 ();
 sg13g2_fill_1 FILLER_15_278 ();
 sg13g2_fill_1 FILLER_15_336 ();
 sg13g2_fill_1 FILLER_15_355 ();
 sg13g2_fill_2 FILLER_15_396 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_4 FILLER_15_417 ();
 sg13g2_fill_2 FILLER_15_421 ();
 sg13g2_fill_1 FILLER_15_432 ();
 sg13g2_decap_4 FILLER_15_451 ();
 sg13g2_fill_2 FILLER_15_455 ();
 sg13g2_fill_1 FILLER_15_475 ();
 sg13g2_fill_1 FILLER_15_490 ();
 sg13g2_decap_4 FILLER_15_496 ();
 sg13g2_fill_1 FILLER_15_500 ();
 sg13g2_fill_2 FILLER_15_505 ();
 sg13g2_fill_1 FILLER_15_507 ();
 sg13g2_fill_2 FILLER_15_522 ();
 sg13g2_fill_1 FILLER_15_524 ();
 sg13g2_fill_2 FILLER_15_552 ();
 sg13g2_fill_1 FILLER_15_554 ();
 sg13g2_fill_2 FILLER_15_559 ();
 sg13g2_fill_2 FILLER_15_602 ();
 sg13g2_fill_1 FILLER_15_604 ();
 sg13g2_decap_4 FILLER_15_632 ();
 sg13g2_fill_1 FILLER_15_636 ();
 sg13g2_fill_1 FILLER_15_650 ();
 sg13g2_fill_1 FILLER_15_678 ();
 sg13g2_decap_8 FILLER_15_683 ();
 sg13g2_fill_2 FILLER_15_690 ();
 sg13g2_fill_1 FILLER_15_692 ();
 sg13g2_fill_1 FILLER_15_724 ();
 sg13g2_fill_2 FILLER_15_736 ();
 sg13g2_decap_4 FILLER_15_742 ();
 sg13g2_fill_2 FILLER_15_746 ();
 sg13g2_decap_4 FILLER_15_753 ();
 sg13g2_decap_4 FILLER_15_770 ();
 sg13g2_decap_8 FILLER_15_842 ();
 sg13g2_decap_8 FILLER_15_849 ();
 sg13g2_decap_4 FILLER_15_856 ();
 sg13g2_fill_2 FILLER_15_860 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_2 ();
 sg13g2_fill_1 FILLER_16_34 ();
 sg13g2_fill_2 FILLER_16_62 ();
 sg13g2_fill_1 FILLER_16_64 ();
 sg13g2_fill_2 FILLER_16_75 ();
 sg13g2_fill_1 FILLER_16_77 ();
 sg13g2_fill_1 FILLER_16_105 ();
 sg13g2_fill_2 FILLER_16_142 ();
 sg13g2_fill_1 FILLER_16_144 ();
 sg13g2_fill_2 FILLER_16_157 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_fill_1 FILLER_16_290 ();
 sg13g2_fill_1 FILLER_16_300 ();
 sg13g2_fill_2 FILLER_16_324 ();
 sg13g2_fill_2 FILLER_16_339 ();
 sg13g2_decap_8 FILLER_16_376 ();
 sg13g2_fill_1 FILLER_16_383 ();
 sg13g2_fill_2 FILLER_16_397 ();
 sg13g2_fill_2 FILLER_16_448 ();
 sg13g2_fill_2 FILLER_16_486 ();
 sg13g2_fill_2 FILLER_16_524 ();
 sg13g2_fill_1 FILLER_16_526 ();
 sg13g2_decap_4 FILLER_16_541 ();
 sg13g2_decap_4 FILLER_16_558 ();
 sg13g2_fill_1 FILLER_16_567 ();
 sg13g2_fill_2 FILLER_16_581 ();
 sg13g2_fill_1 FILLER_16_583 ();
 sg13g2_decap_8 FILLER_16_590 ();
 sg13g2_decap_8 FILLER_16_597 ();
 sg13g2_fill_2 FILLER_16_604 ();
 sg13g2_fill_1 FILLER_16_606 ();
 sg13g2_decap_4 FILLER_16_612 ();
 sg13g2_decap_8 FILLER_16_620 ();
 sg13g2_fill_1 FILLER_16_627 ();
 sg13g2_fill_2 FILLER_16_637 ();
 sg13g2_fill_1 FILLER_16_639 ();
 sg13g2_fill_2 FILLER_16_664 ();
 sg13g2_fill_1 FILLER_16_666 ();
 sg13g2_fill_1 FILLER_16_676 ();
 sg13g2_fill_2 FILLER_16_708 ();
 sg13g2_fill_1 FILLER_16_728 ();
 sg13g2_fill_2 FILLER_16_787 ();
 sg13g2_fill_1 FILLER_16_789 ();
 sg13g2_fill_2 FILLER_16_821 ();
 sg13g2_fill_1 FILLER_16_823 ();
 sg13g2_decap_8 FILLER_16_846 ();
 sg13g2_decap_8 FILLER_16_853 ();
 sg13g2_fill_2 FILLER_16_860 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_7 ();
 sg13g2_decap_4 FILLER_17_12 ();
 sg13g2_fill_2 FILLER_17_26 ();
 sg13g2_fill_1 FILLER_17_28 ();
 sg13g2_fill_1 FILLER_17_38 ();
 sg13g2_fill_2 FILLER_17_52 ();
 sg13g2_decap_4 FILLER_17_90 ();
 sg13g2_fill_2 FILLER_17_99 ();
 sg13g2_fill_2 FILLER_17_114 ();
 sg13g2_fill_1 FILLER_17_116 ();
 sg13g2_fill_2 FILLER_17_126 ();
 sg13g2_fill_1 FILLER_17_128 ();
 sg13g2_fill_1 FILLER_17_138 ();
 sg13g2_decap_4 FILLER_17_171 ();
 sg13g2_decap_4 FILLER_17_179 ();
 sg13g2_fill_1 FILLER_17_183 ();
 sg13g2_fill_1 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_223 ();
 sg13g2_fill_1 FILLER_17_230 ();
 sg13g2_decap_4 FILLER_17_239 ();
 sg13g2_fill_2 FILLER_17_261 ();
 sg13g2_fill_1 FILLER_17_263 ();
 sg13g2_fill_1 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_355 ();
 sg13g2_decap_8 FILLER_17_362 ();
 sg13g2_fill_2 FILLER_17_369 ();
 sg13g2_fill_1 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_412 ();
 sg13g2_fill_2 FILLER_17_419 ();
 sg13g2_fill_2 FILLER_17_434 ();
 sg13g2_fill_1 FILLER_17_463 ();
 sg13g2_decap_4 FILLER_17_468 ();
 sg13g2_fill_1 FILLER_17_472 ();
 sg13g2_decap_8 FILLER_17_477 ();
 sg13g2_fill_1 FILLER_17_489 ();
 sg13g2_fill_2 FILLER_17_498 ();
 sg13g2_fill_1 FILLER_17_500 ();
 sg13g2_fill_1 FILLER_17_516 ();
 sg13g2_decap_8 FILLER_17_521 ();
 sg13g2_fill_2 FILLER_17_533 ();
 sg13g2_decap_4 FILLER_17_639 ();
 sg13g2_fill_2 FILLER_17_643 ();
 sg13g2_fill_2 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_4 FILLER_17_707 ();
 sg13g2_fill_1 FILLER_17_711 ();
 sg13g2_fill_2 FILLER_17_728 ();
 sg13g2_fill_1 FILLER_17_734 ();
 sg13g2_decap_4 FILLER_17_808 ();
 sg13g2_fill_2 FILLER_17_821 ();
 sg13g2_fill_1 FILLER_17_823 ();
 sg13g2_decap_8 FILLER_17_851 ();
 sg13g2_decap_4 FILLER_17_858 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_2 ();
 sg13g2_decap_8 FILLER_18_43 ();
 sg13g2_fill_1 FILLER_18_55 ();
 sg13g2_fill_1 FILLER_18_104 ();
 sg13g2_fill_1 FILLER_18_114 ();
 sg13g2_fill_2 FILLER_18_128 ();
 sg13g2_fill_1 FILLER_18_130 ();
 sg13g2_fill_2 FILLER_18_136 ();
 sg13g2_fill_1 FILLER_18_138 ();
 sg13g2_decap_8 FILLER_18_157 ();
 sg13g2_decap_4 FILLER_18_164 ();
 sg13g2_fill_2 FILLER_18_168 ();
 sg13g2_fill_1 FILLER_18_197 ();
 sg13g2_fill_2 FILLER_18_215 ();
 sg13g2_decap_4 FILLER_18_249 ();
 sg13g2_fill_2 FILLER_18_294 ();
 sg13g2_fill_1 FILLER_18_296 ();
 sg13g2_decap_8 FILLER_18_311 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_fill_2 FILLER_18_382 ();
 sg13g2_fill_1 FILLER_18_384 ();
 sg13g2_fill_2 FILLER_18_412 ();
 sg13g2_decap_4 FILLER_18_422 ();
 sg13g2_fill_1 FILLER_18_439 ();
 sg13g2_fill_2 FILLER_18_455 ();
 sg13g2_fill_1 FILLER_18_457 ();
 sg13g2_fill_2 FILLER_18_467 ();
 sg13g2_fill_1 FILLER_18_469 ();
 sg13g2_fill_2 FILLER_18_510 ();
 sg13g2_fill_2 FILLER_18_556 ();
 sg13g2_fill_1 FILLER_18_590 ();
 sg13g2_fill_2 FILLER_18_600 ();
 sg13g2_fill_2 FILLER_18_625 ();
 sg13g2_fill_2 FILLER_18_631 ();
 sg13g2_fill_1 FILLER_18_654 ();
 sg13g2_decap_4 FILLER_18_659 ();
 sg13g2_fill_2 FILLER_18_663 ();
 sg13g2_fill_1 FILLER_18_686 ();
 sg13g2_decap_4 FILLER_18_700 ();
 sg13g2_fill_1 FILLER_18_708 ();
 sg13g2_fill_2 FILLER_18_717 ();
 sg13g2_fill_1 FILLER_18_719 ();
 sg13g2_fill_2 FILLER_18_761 ();
 sg13g2_fill_1 FILLER_18_834 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_4 ();
 sg13g2_decap_8 FILLER_19_13 ();
 sg13g2_fill_2 FILLER_19_20 ();
 sg13g2_fill_2 FILLER_19_27 ();
 sg13g2_fill_2 FILLER_19_69 ();
 sg13g2_fill_1 FILLER_19_71 ();
 sg13g2_fill_2 FILLER_19_81 ();
 sg13g2_fill_1 FILLER_19_97 ();
 sg13g2_fill_2 FILLER_19_109 ();
 sg13g2_fill_1 FILLER_19_111 ();
 sg13g2_fill_1 FILLER_19_160 ();
 sg13g2_decap_8 FILLER_19_179 ();
 sg13g2_decap_8 FILLER_19_250 ();
 sg13g2_fill_2 FILLER_19_257 ();
 sg13g2_fill_1 FILLER_19_267 ();
 sg13g2_decap_4 FILLER_19_272 ();
 sg13g2_fill_1 FILLER_19_276 ();
 sg13g2_fill_1 FILLER_19_290 ();
 sg13g2_fill_2 FILLER_19_318 ();
 sg13g2_fill_1 FILLER_19_320 ();
 sg13g2_decap_8 FILLER_19_330 ();
 sg13g2_decap_8 FILLER_19_337 ();
 sg13g2_fill_2 FILLER_19_344 ();
 sg13g2_fill_1 FILLER_19_346 ();
 sg13g2_fill_2 FILLER_19_356 ();
 sg13g2_fill_2 FILLER_19_373 ();
 sg13g2_fill_1 FILLER_19_380 ();
 sg13g2_decap_8 FILLER_19_426 ();
 sg13g2_fill_1 FILLER_19_433 ();
 sg13g2_decap_4 FILLER_19_496 ();
 sg13g2_decap_8 FILLER_19_504 ();
 sg13g2_decap_8 FILLER_19_511 ();
 sg13g2_decap_4 FILLER_19_549 ();
 sg13g2_fill_2 FILLER_19_553 ();
 sg13g2_fill_1 FILLER_19_591 ();
 sg13g2_fill_2 FILLER_19_655 ();
 sg13g2_fill_1 FILLER_19_657 ();
 sg13g2_fill_2 FILLER_19_685 ();
 sg13g2_fill_2 FILLER_19_736 ();
 sg13g2_decap_8 FILLER_19_751 ();
 sg13g2_decap_8 FILLER_19_789 ();
 sg13g2_fill_2 FILLER_19_835 ();
 sg13g2_fill_2 FILLER_19_846 ();
 sg13g2_fill_1 FILLER_19_861 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_44 ();
 sg13g2_fill_1 FILLER_20_46 ();
 sg13g2_decap_4 FILLER_20_87 ();
 sg13g2_decap_4 FILLER_20_128 ();
 sg13g2_fill_2 FILLER_20_132 ();
 sg13g2_fill_2 FILLER_20_161 ();
 sg13g2_fill_1 FILLER_20_163 ();
 sg13g2_decap_8 FILLER_20_191 ();
 sg13g2_fill_1 FILLER_20_198 ();
 sg13g2_fill_2 FILLER_20_211 ();
 sg13g2_decap_4 FILLER_20_222 ();
 sg13g2_fill_1 FILLER_20_226 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_fill_2 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_244 ();
 sg13g2_decap_8 FILLER_20_251 ();
 sg13g2_fill_2 FILLER_20_258 ();
 sg13g2_fill_2 FILLER_20_300 ();
 sg13g2_fill_1 FILLER_20_302 ();
 sg13g2_fill_2 FILLER_20_344 ();
 sg13g2_decap_4 FILLER_20_373 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_fill_2 FILLER_20_405 ();
 sg13g2_decap_4 FILLER_20_440 ();
 sg13g2_fill_1 FILLER_20_444 ();
 sg13g2_decap_8 FILLER_20_449 ();
 sg13g2_decap_8 FILLER_20_456 ();
 sg13g2_fill_1 FILLER_20_463 ();
 sg13g2_fill_1 FILLER_20_522 ();
 sg13g2_fill_2 FILLER_20_558 ();
 sg13g2_decap_8 FILLER_20_564 ();
 sg13g2_decap_8 FILLER_20_571 ();
 sg13g2_decap_4 FILLER_20_578 ();
 sg13g2_fill_2 FILLER_20_582 ();
 sg13g2_fill_2 FILLER_20_594 ();
 sg13g2_decap_4 FILLER_20_605 ();
 sg13g2_fill_1 FILLER_20_609 ();
 sg13g2_fill_1 FILLER_20_628 ();
 sg13g2_fill_2 FILLER_20_669 ();
 sg13g2_fill_1 FILLER_20_671 ();
 sg13g2_fill_2 FILLER_20_681 ();
 sg13g2_fill_1 FILLER_20_683 ();
 sg13g2_fill_1 FILLER_20_697 ();
 sg13g2_fill_1 FILLER_20_707 ();
 sg13g2_fill_1 FILLER_20_721 ();
 sg13g2_decap_8 FILLER_20_766 ();
 sg13g2_decap_4 FILLER_20_805 ();
 sg13g2_decap_4 FILLER_20_858 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_fill_2 FILLER_21_28 ();
 sg13g2_fill_2 FILLER_21_35 ();
 sg13g2_decap_4 FILLER_21_41 ();
 sg13g2_decap_8 FILLER_21_58 ();
 sg13g2_decap_8 FILLER_21_65 ();
 sg13g2_decap_8 FILLER_21_85 ();
 sg13g2_decap_8 FILLER_21_92 ();
 sg13g2_decap_4 FILLER_21_99 ();
 sg13g2_fill_1 FILLER_21_103 ();
 sg13g2_decap_8 FILLER_21_117 ();
 sg13g2_fill_1 FILLER_21_124 ();
 sg13g2_decap_4 FILLER_21_134 ();
 sg13g2_fill_1 FILLER_21_147 ();
 sg13g2_decap_4 FILLER_21_152 ();
 sg13g2_fill_2 FILLER_21_165 ();
 sg13g2_fill_1 FILLER_21_225 ();
 sg13g2_decap_8 FILLER_21_262 ();
 sg13g2_fill_1 FILLER_21_269 ();
 sg13g2_decap_4 FILLER_21_274 ();
 sg13g2_fill_2 FILLER_21_278 ();
 sg13g2_fill_2 FILLER_21_291 ();
 sg13g2_fill_1 FILLER_21_293 ();
 sg13g2_fill_1 FILLER_21_307 ();
 sg13g2_fill_2 FILLER_21_317 ();
 sg13g2_decap_8 FILLER_21_356 ();
 sg13g2_decap_4 FILLER_21_363 ();
 sg13g2_decap_8 FILLER_21_404 ();
 sg13g2_fill_2 FILLER_21_411 ();
 sg13g2_fill_1 FILLER_21_413 ();
 sg13g2_fill_1 FILLER_21_418 ();
 sg13g2_decap_4 FILLER_21_423 ();
 sg13g2_fill_1 FILLER_21_427 ();
 sg13g2_fill_2 FILLER_21_446 ();
 sg13g2_fill_1 FILLER_21_448 ();
 sg13g2_decap_8 FILLER_21_455 ();
 sg13g2_fill_1 FILLER_21_462 ();
 sg13g2_fill_1 FILLER_21_499 ();
 sg13g2_fill_2 FILLER_21_510 ();
 sg13g2_decap_4 FILLER_21_521 ();
 sg13g2_fill_2 FILLER_21_525 ();
 sg13g2_fill_1 FILLER_21_553 ();
 sg13g2_decap_8 FILLER_21_563 ();
 sg13g2_decap_4 FILLER_21_570 ();
 sg13g2_fill_1 FILLER_21_574 ();
 sg13g2_decap_4 FILLER_21_580 ();
 sg13g2_fill_2 FILLER_21_584 ();
 sg13g2_decap_4 FILLER_21_591 ();
 sg13g2_fill_1 FILLER_21_595 ();
 sg13g2_fill_2 FILLER_21_602 ();
 sg13g2_fill_1 FILLER_21_604 ();
 sg13g2_decap_8 FILLER_21_669 ();
 sg13g2_decap_8 FILLER_21_676 ();
 sg13g2_fill_2 FILLER_21_719 ();
 sg13g2_fill_1 FILLER_21_721 ();
 sg13g2_fill_1 FILLER_21_731 ();
 sg13g2_fill_2 FILLER_21_746 ();
 sg13g2_fill_1 FILLER_21_748 ();
 sg13g2_decap_4 FILLER_21_776 ();
 sg13g2_fill_1 FILLER_21_780 ();
 sg13g2_fill_1 FILLER_21_789 ();
 sg13g2_fill_2 FILLER_21_803 ();
 sg13g2_fill_1 FILLER_21_805 ();
 sg13g2_fill_2 FILLER_21_833 ();
 sg13g2_fill_1 FILLER_21_835 ();
 sg13g2_fill_1 FILLER_21_844 ();
 sg13g2_decap_8 FILLER_21_854 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_fill_2 FILLER_22_21 ();
 sg13g2_fill_1 FILLER_22_50 ();
 sg13g2_fill_2 FILLER_22_88 ();
 sg13g2_fill_1 FILLER_22_90 ();
 sg13g2_fill_2 FILLER_22_104 ();
 sg13g2_fill_1 FILLER_22_106 ();
 sg13g2_fill_2 FILLER_22_134 ();
 sg13g2_fill_1 FILLER_22_136 ();
 sg13g2_decap_4 FILLER_22_142 ();
 sg13g2_fill_1 FILLER_22_146 ();
 sg13g2_decap_8 FILLER_22_205 ();
 sg13g2_fill_1 FILLER_22_212 ();
 sg13g2_decap_8 FILLER_22_272 ();
 sg13g2_decap_4 FILLER_22_279 ();
 sg13g2_fill_2 FILLER_22_289 ();
 sg13g2_fill_2 FILLER_22_318 ();
 sg13g2_fill_1 FILLER_22_347 ();
 sg13g2_fill_1 FILLER_22_366 ();
 sg13g2_fill_2 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_424 ();
 sg13g2_fill_1 FILLER_22_466 ();
 sg13g2_fill_1 FILLER_22_496 ();
 sg13g2_fill_2 FILLER_22_541 ();
 sg13g2_fill_1 FILLER_22_573 ();
 sg13g2_decap_4 FILLER_22_607 ();
 sg13g2_decap_4 FILLER_22_628 ();
 sg13g2_fill_1 FILLER_22_632 ();
 sg13g2_decap_8 FILLER_22_653 ();
 sg13g2_decap_8 FILLER_22_664 ();
 sg13g2_fill_2 FILLER_22_671 ();
 sg13g2_decap_4 FILLER_22_684 ();
 sg13g2_fill_1 FILLER_22_688 ();
 sg13g2_fill_2 FILLER_22_701 ();
 sg13g2_fill_1 FILLER_22_748 ();
 sg13g2_decap_4 FILLER_22_759 ();
 sg13g2_fill_1 FILLER_22_763 ();
 sg13g2_fill_2 FILLER_22_773 ();
 sg13g2_fill_1 FILLER_22_787 ();
 sg13g2_fill_2 FILLER_22_798 ();
 sg13g2_fill_1 FILLER_22_800 ();
 sg13g2_fill_1 FILLER_22_828 ();
 sg13g2_fill_1 FILLER_22_834 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_4 FILLER_23_45 ();
 sg13g2_fill_2 FILLER_23_49 ();
 sg13g2_fill_2 FILLER_23_90 ();
 sg13g2_fill_2 FILLER_23_109 ();
 sg13g2_fill_1 FILLER_23_111 ();
 sg13g2_decap_8 FILLER_23_116 ();
 sg13g2_decap_8 FILLER_23_123 ();
 sg13g2_decap_4 FILLER_23_130 ();
 sg13g2_decap_4 FILLER_23_177 ();
 sg13g2_fill_2 FILLER_23_212 ();
 sg13g2_decap_8 FILLER_23_223 ();
 sg13g2_fill_1 FILLER_23_230 ();
 sg13g2_fill_2 FILLER_23_287 ();
 sg13g2_fill_2 FILLER_23_295 ();
 sg13g2_fill_1 FILLER_23_314 ();
 sg13g2_fill_1 FILLER_23_324 ();
 sg13g2_fill_2 FILLER_23_329 ();
 sg13g2_fill_1 FILLER_23_331 ();
 sg13g2_decap_4 FILLER_23_341 ();
 sg13g2_fill_1 FILLER_23_345 ();
 sg13g2_decap_4 FILLER_23_351 ();
 sg13g2_fill_1 FILLER_23_355 ();
 sg13g2_fill_2 FILLER_23_392 ();
 sg13g2_decap_4 FILLER_23_421 ();
 sg13g2_decap_8 FILLER_23_438 ();
 sg13g2_decap_8 FILLER_23_445 ();
 sg13g2_decap_4 FILLER_23_452 ();
 sg13g2_fill_1 FILLER_23_534 ();
 sg13g2_fill_1 FILLER_23_562 ();
 sg13g2_fill_2 FILLER_23_566 ();
 sg13g2_fill_2 FILLER_23_583 ();
 sg13g2_decap_4 FILLER_23_589 ();
 sg13g2_fill_2 FILLER_23_632 ();
 sg13g2_fill_1 FILLER_23_634 ();
 sg13g2_fill_2 FILLER_23_653 ();
 sg13g2_fill_1 FILLER_23_688 ();
 sg13g2_fill_1 FILLER_23_695 ();
 sg13g2_decap_8 FILLER_23_711 ();
 sg13g2_fill_2 FILLER_23_718 ();
 sg13g2_fill_1 FILLER_23_720 ();
 sg13g2_fill_2 FILLER_23_738 ();
 sg13g2_fill_1 FILLER_23_776 ();
 sg13g2_fill_2 FILLER_23_786 ();
 sg13g2_fill_2 FILLER_23_821 ();
 sg13g2_fill_1 FILLER_23_823 ();
 sg13g2_fill_1 FILLER_23_837 ();
 sg13g2_fill_1 FILLER_23_842 ();
 sg13g2_decap_8 FILLER_23_852 ();
 sg13g2_fill_2 FILLER_23_859 ();
 sg13g2_fill_1 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_7 ();
 sg13g2_fill_1 FILLER_24_40 ();
 sg13g2_fill_2 FILLER_24_62 ();
 sg13g2_fill_1 FILLER_24_64 ();
 sg13g2_fill_2 FILLER_24_70 ();
 sg13g2_fill_1 FILLER_24_72 ();
 sg13g2_fill_1 FILLER_24_109 ();
 sg13g2_decap_4 FILLER_24_166 ();
 sg13g2_fill_1 FILLER_24_170 ();
 sg13g2_decap_4 FILLER_24_180 ();
 sg13g2_fill_2 FILLER_24_184 ();
 sg13g2_fill_1 FILLER_24_190 ();
 sg13g2_fill_2 FILLER_24_197 ();
 sg13g2_fill_2 FILLER_24_205 ();
 sg13g2_fill_1 FILLER_24_207 ();
 sg13g2_decap_4 FILLER_24_217 ();
 sg13g2_fill_2 FILLER_24_221 ();
 sg13g2_decap_8 FILLER_24_228 ();
 sg13g2_fill_1 FILLER_24_235 ();
 sg13g2_fill_2 FILLER_24_251 ();
 sg13g2_fill_2 FILLER_24_258 ();
 sg13g2_fill_1 FILLER_24_260 ();
 sg13g2_fill_2 FILLER_24_276 ();
 sg13g2_fill_1 FILLER_24_288 ();
 sg13g2_fill_1 FILLER_24_295 ();
 sg13g2_fill_2 FILLER_24_328 ();
 sg13g2_fill_2 FILLER_24_334 ();
 sg13g2_fill_1 FILLER_24_336 ();
 sg13g2_fill_2 FILLER_24_373 ();
 sg13g2_fill_1 FILLER_24_375 ();
 sg13g2_decap_8 FILLER_24_403 ();
 sg13g2_fill_2 FILLER_24_410 ();
 sg13g2_fill_2 FILLER_24_462 ();
 sg13g2_decap_8 FILLER_24_501 ();
 sg13g2_fill_2 FILLER_24_508 ();
 sg13g2_fill_2 FILLER_24_523 ();
 sg13g2_decap_4 FILLER_24_562 ();
 sg13g2_fill_2 FILLER_24_566 ();
 sg13g2_fill_1 FILLER_24_573 ();
 sg13g2_decap_8 FILLER_24_578 ();
 sg13g2_decap_8 FILLER_24_585 ();
 sg13g2_decap_8 FILLER_24_592 ();
 sg13g2_fill_1 FILLER_24_599 ();
 sg13g2_decap_8 FILLER_24_658 ();
 sg13g2_fill_1 FILLER_24_665 ();
 sg13g2_fill_1 FILLER_24_679 ();
 sg13g2_fill_1 FILLER_24_729 ();
 sg13g2_fill_2 FILLER_24_756 ();
 sg13g2_fill_1 FILLER_24_758 ();
 sg13g2_fill_1 FILLER_24_772 ();
 sg13g2_decap_4 FILLER_24_778 ();
 sg13g2_fill_2 FILLER_24_782 ();
 sg13g2_fill_1 FILLER_24_788 ();
 sg13g2_fill_2 FILLER_24_794 ();
 sg13g2_decap_4 FILLER_24_810 ();
 sg13g2_fill_1 FILLER_24_814 ();
 sg13g2_fill_2 FILLER_24_819 ();
 sg13g2_fill_1 FILLER_24_821 ();
 sg13g2_fill_2 FILLER_24_831 ();
 sg13g2_fill_2 FILLER_24_860 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_7 ();
 sg13g2_fill_2 FILLER_25_11 ();
 sg13g2_decap_8 FILLER_25_17 ();
 sg13g2_fill_1 FILLER_25_24 ();
 sg13g2_decap_4 FILLER_25_74 ();
 sg13g2_decap_8 FILLER_25_82 ();
 sg13g2_decap_4 FILLER_25_89 ();
 sg13g2_fill_1 FILLER_25_93 ();
 sg13g2_fill_2 FILLER_25_152 ();
 sg13g2_decap_8 FILLER_25_190 ();
 sg13g2_fill_1 FILLER_25_197 ();
 sg13g2_fill_2 FILLER_25_204 ();
 sg13g2_fill_1 FILLER_25_280 ();
 sg13g2_fill_2 FILLER_25_316 ();
 sg13g2_fill_1 FILLER_25_318 ();
 sg13g2_fill_1 FILLER_25_366 ();
 sg13g2_decap_4 FILLER_25_411 ();
 sg13g2_fill_2 FILLER_25_415 ();
 sg13g2_decap_4 FILLER_25_421 ();
 sg13g2_fill_2 FILLER_25_425 ();
 sg13g2_fill_2 FILLER_25_436 ();
 sg13g2_fill_1 FILLER_25_438 ();
 sg13g2_fill_1 FILLER_25_448 ();
 sg13g2_fill_2 FILLER_25_454 ();
 sg13g2_fill_2 FILLER_25_505 ();
 sg13g2_decap_4 FILLER_25_516 ();
 sg13g2_fill_1 FILLER_25_520 ();
 sg13g2_fill_2 FILLER_25_558 ();
 sg13g2_fill_1 FILLER_25_560 ();
 sg13g2_fill_2 FILLER_25_566 ();
 sg13g2_fill_1 FILLER_25_568 ();
 sg13g2_decap_4 FILLER_25_596 ();
 sg13g2_fill_2 FILLER_25_600 ();
 sg13g2_decap_8 FILLER_25_628 ();
 sg13g2_fill_2 FILLER_25_665 ();
 sg13g2_fill_1 FILLER_25_699 ();
 sg13g2_fill_1 FILLER_25_713 ();
 sg13g2_decap_4 FILLER_25_723 ();
 sg13g2_fill_1 FILLER_25_727 ();
 sg13g2_decap_8 FILLER_25_733 ();
 sg13g2_fill_2 FILLER_25_740 ();
 sg13g2_fill_1 FILLER_25_742 ();
 sg13g2_decap_8 FILLER_25_837 ();
 sg13g2_decap_8 FILLER_25_844 ();
 sg13g2_decap_8 FILLER_25_851 ();
 sg13g2_decap_4 FILLER_25_858 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_14 ();
 sg13g2_decap_4 FILLER_26_19 ();
 sg13g2_fill_2 FILLER_26_23 ();
 sg13g2_decap_8 FILLER_26_30 ();
 sg13g2_decap_8 FILLER_26_41 ();
 sg13g2_fill_2 FILLER_26_48 ();
 sg13g2_decap_8 FILLER_26_54 ();
 sg13g2_fill_2 FILLER_26_61 ();
 sg13g2_fill_1 FILLER_26_63 ();
 sg13g2_fill_2 FILLER_26_79 ();
 sg13g2_decap_4 FILLER_26_89 ();
 sg13g2_fill_1 FILLER_26_93 ();
 sg13g2_fill_1 FILLER_26_103 ();
 sg13g2_fill_1 FILLER_26_149 ();
 sg13g2_fill_1 FILLER_26_167 ();
 sg13g2_fill_2 FILLER_26_181 ();
 sg13g2_fill_2 FILLER_26_188 ();
 sg13g2_decap_8 FILLER_26_194 ();
 sg13g2_decap_4 FILLER_26_201 ();
 sg13g2_fill_2 FILLER_26_222 ();
 sg13g2_fill_1 FILLER_26_224 ();
 sg13g2_fill_1 FILLER_26_314 ();
 sg13g2_fill_2 FILLER_26_324 ();
 sg13g2_fill_1 FILLER_26_326 ();
 sg13g2_fill_1 FILLER_26_358 ();
 sg13g2_fill_2 FILLER_26_373 ();
 sg13g2_fill_1 FILLER_26_375 ();
 sg13g2_fill_1 FILLER_26_389 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_fill_1 FILLER_26_409 ();
 sg13g2_fill_2 FILLER_26_415 ();
 sg13g2_decap_4 FILLER_26_421 ();
 sg13g2_fill_1 FILLER_26_435 ();
 sg13g2_fill_1 FILLER_26_445 ();
 sg13g2_fill_1 FILLER_26_473 ();
 sg13g2_fill_1 FILLER_26_478 ();
 sg13g2_decap_4 FILLER_26_492 ();
 sg13g2_fill_1 FILLER_26_536 ();
 sg13g2_fill_2 FILLER_26_550 ();
 sg13g2_fill_1 FILLER_26_606 ();
 sg13g2_fill_2 FILLER_26_634 ();
 sg13g2_fill_1 FILLER_26_671 ();
 sg13g2_decap_8 FILLER_26_676 ();
 sg13g2_decap_8 FILLER_26_683 ();
 sg13g2_fill_1 FILLER_26_690 ();
 sg13g2_decap_8 FILLER_26_767 ();
 sg13g2_decap_8 FILLER_26_778 ();
 sg13g2_decap_8 FILLER_26_785 ();
 sg13g2_fill_1 FILLER_26_792 ();
 sg13g2_decap_8 FILLER_26_819 ();
 sg13g2_fill_2 FILLER_26_826 ();
 sg13g2_decap_8 FILLER_26_833 ();
 sg13g2_decap_8 FILLER_26_844 ();
 sg13g2_decap_8 FILLER_26_851 ();
 sg13g2_decap_4 FILLER_26_858 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_7 ();
 sg13g2_fill_1 FILLER_27_9 ();
 sg13g2_fill_2 FILLER_27_42 ();
 sg13g2_fill_1 FILLER_27_44 ();
 sg13g2_fill_2 FILLER_27_90 ();
 sg13g2_fill_2 FILLER_27_109 ();
 sg13g2_fill_2 FILLER_27_138 ();
 sg13g2_fill_1 FILLER_27_140 ();
 sg13g2_fill_2 FILLER_27_149 ();
 sg13g2_decap_8 FILLER_27_173 ();
 sg13g2_fill_2 FILLER_27_220 ();
 sg13g2_fill_1 FILLER_27_222 ();
 sg13g2_fill_1 FILLER_27_228 ();
 sg13g2_fill_1 FILLER_27_269 ();
 sg13g2_fill_1 FILLER_27_284 ();
 sg13g2_fill_2 FILLER_27_370 ();
 sg13g2_fill_2 FILLER_27_390 ();
 sg13g2_fill_1 FILLER_27_392 ();
 sg13g2_fill_2 FILLER_27_443 ();
 sg13g2_fill_1 FILLER_27_445 ();
 sg13g2_fill_1 FILLER_27_466 ();
 sg13g2_fill_2 FILLER_27_476 ();
 sg13g2_fill_1 FILLER_27_491 ();
 sg13g2_decap_4 FILLER_27_518 ();
 sg13g2_fill_1 FILLER_27_522 ();
 sg13g2_fill_2 FILLER_27_573 ();
 sg13g2_fill_1 FILLER_27_575 ();
 sg13g2_fill_2 FILLER_27_607 ();
 sg13g2_decap_4 FILLER_27_636 ();
 sg13g2_decap_4 FILLER_27_649 ();
 sg13g2_fill_1 FILLER_27_653 ();
 sg13g2_fill_2 FILLER_27_698 ();
 sg13g2_fill_1 FILLER_27_700 ();
 sg13g2_decap_4 FILLER_27_726 ();
 sg13g2_fill_2 FILLER_27_730 ();
 sg13g2_fill_2 FILLER_27_736 ();
 sg13g2_fill_1 FILLER_27_738 ();
 sg13g2_decap_8 FILLER_27_748 ();
 sg13g2_fill_2 FILLER_27_755 ();
 sg13g2_fill_1 FILLER_27_757 ();
 sg13g2_fill_1 FILLER_27_763 ();
 sg13g2_fill_2 FILLER_27_802 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_2 ();
 sg13g2_decap_4 FILLER_28_48 ();
 sg13g2_fill_2 FILLER_28_79 ();
 sg13g2_fill_1 FILLER_28_81 ();
 sg13g2_fill_1 FILLER_28_95 ();
 sg13g2_fill_1 FILLER_28_141 ();
 sg13g2_fill_1 FILLER_28_156 ();
 sg13g2_fill_2 FILLER_28_182 ();
 sg13g2_fill_1 FILLER_28_184 ();
 sg13g2_fill_2 FILLER_28_193 ();
 sg13g2_fill_1 FILLER_28_195 ();
 sg13g2_decap_4 FILLER_28_202 ();
 sg13g2_fill_1 FILLER_28_247 ();
 sg13g2_decap_4 FILLER_28_261 ();
 sg13g2_fill_1 FILLER_28_265 ();
 sg13g2_fill_2 FILLER_28_308 ();
 sg13g2_fill_2 FILLER_28_378 ();
 sg13g2_decap_4 FILLER_28_420 ();
 sg13g2_fill_1 FILLER_28_424 ();
 sg13g2_decap_4 FILLER_28_460 ();
 sg13g2_fill_2 FILLER_28_464 ();
 sg13g2_decap_4 FILLER_28_541 ();
 sg13g2_fill_1 FILLER_28_545 ();
 sg13g2_fill_2 FILLER_28_550 ();
 sg13g2_fill_1 FILLER_28_552 ();
 sg13g2_decap_8 FILLER_28_565 ();
 sg13g2_decap_4 FILLER_28_594 ();
 sg13g2_fill_1 FILLER_28_598 ();
 sg13g2_fill_1 FILLER_28_604 ();
 sg13g2_fill_1 FILLER_28_626 ();
 sg13g2_fill_2 FILLER_28_654 ();
 sg13g2_fill_1 FILLER_28_656 ();
 sg13g2_fill_1 FILLER_28_670 ();
 sg13g2_fill_2 FILLER_28_712 ();
 sg13g2_fill_1 FILLER_28_714 ();
 sg13g2_fill_2 FILLER_28_726 ();
 sg13g2_fill_1 FILLER_28_728 ();
 sg13g2_decap_4 FILLER_28_733 ();
 sg13g2_fill_2 FILLER_28_737 ();
 sg13g2_decap_4 FILLER_28_782 ();
 sg13g2_fill_2 FILLER_28_786 ();
 sg13g2_fill_2 FILLER_28_797 ();
 sg13g2_fill_1 FILLER_28_799 ();
 sg13g2_decap_8 FILLER_28_822 ();
 sg13g2_fill_1 FILLER_28_833 ();
 sg13g2_decap_4 FILLER_28_856 ();
 sg13g2_fill_2 FILLER_28_860 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_35 ();
 sg13g2_fill_1 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_61 ();
 sg13g2_fill_1 FILLER_29_68 ();
 sg13g2_fill_2 FILLER_29_94 ();
 sg13g2_fill_1 FILLER_29_96 ();
 sg13g2_decap_4 FILLER_29_129 ();
 sg13g2_fill_1 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_169 ();
 sg13g2_fill_1 FILLER_29_203 ();
 sg13g2_decap_4 FILLER_29_212 ();
 sg13g2_fill_2 FILLER_29_216 ();
 sg13g2_fill_2 FILLER_29_248 ();
 sg13g2_fill_1 FILLER_29_250 ();
 sg13g2_fill_2 FILLER_29_264 ();
 sg13g2_fill_1 FILLER_29_266 ();
 sg13g2_fill_2 FILLER_29_280 ();
 sg13g2_fill_2 FILLER_29_296 ();
 sg13g2_fill_1 FILLER_29_329 ();
 sg13g2_fill_2 FILLER_29_343 ();
 sg13g2_decap_8 FILLER_29_358 ();
 sg13g2_decap_4 FILLER_29_365 ();
 sg13g2_fill_2 FILLER_29_421 ();
 sg13g2_fill_1 FILLER_29_423 ();
 sg13g2_fill_2 FILLER_29_429 ();
 sg13g2_fill_2 FILLER_29_440 ();
 sg13g2_fill_1 FILLER_29_442 ();
 sg13g2_fill_2 FILLER_29_482 ();
 sg13g2_decap_8 FILLER_29_493 ();
 sg13g2_fill_2 FILLER_29_554 ();
 sg13g2_fill_1 FILLER_29_556 ();
 sg13g2_decap_4 FILLER_29_571 ();
 sg13g2_fill_1 FILLER_29_575 ();
 sg13g2_fill_1 FILLER_29_603 ();
 sg13g2_fill_1 FILLER_29_631 ();
 sg13g2_decap_4 FILLER_29_636 ();
 sg13g2_fill_1 FILLER_29_653 ();
 sg13g2_fill_1 FILLER_29_699 ();
 sg13g2_fill_2 FILLER_29_709 ();
 sg13g2_fill_2 FILLER_29_800 ();
 sg13g2_fill_1 FILLER_29_834 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_44 ();
 sg13g2_fill_1 FILLER_30_87 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_4 FILLER_30_112 ();
 sg13g2_decap_4 FILLER_30_125 ();
 sg13g2_fill_1 FILLER_30_160 ();
 sg13g2_decap_4 FILLER_30_218 ();
 sg13g2_decap_8 FILLER_30_240 ();
 sg13g2_fill_1 FILLER_30_247 ();
 sg13g2_fill_2 FILLER_30_325 ();
 sg13g2_fill_1 FILLER_30_327 ();
 sg13g2_fill_1 FILLER_30_332 ();
 sg13g2_decap_8 FILLER_30_337 ();
 sg13g2_fill_1 FILLER_30_354 ();
 sg13g2_decap_4 FILLER_30_364 ();
 sg13g2_fill_1 FILLER_30_368 ();
 sg13g2_fill_2 FILLER_30_382 ();
 sg13g2_fill_1 FILLER_30_384 ();
 sg13g2_fill_2 FILLER_30_390 ();
 sg13g2_fill_1 FILLER_30_392 ();
 sg13g2_fill_2 FILLER_30_415 ();
 sg13g2_fill_1 FILLER_30_417 ();
 sg13g2_fill_2 FILLER_30_467 ();
 sg13g2_fill_1 FILLER_30_477 ();
 sg13g2_fill_2 FILLER_30_513 ();
 sg13g2_decap_4 FILLER_30_532 ();
 sg13g2_fill_2 FILLER_30_536 ();
 sg13g2_fill_1 FILLER_30_583 ();
 sg13g2_decap_8 FILLER_30_629 ();
 sg13g2_decap_8 FILLER_30_636 ();
 sg13g2_fill_1 FILLER_30_643 ();
 sg13g2_fill_2 FILLER_30_649 ();
 sg13g2_fill_1 FILLER_30_651 ();
 sg13g2_fill_1 FILLER_30_656 ();
 sg13g2_fill_2 FILLER_30_665 ();
 sg13g2_fill_1 FILLER_30_667 ();
 sg13g2_decap_8 FILLER_30_690 ();
 sg13g2_fill_1 FILLER_30_719 ();
 sg13g2_fill_2 FILLER_30_724 ();
 sg13g2_fill_1 FILLER_30_726 ();
 sg13g2_fill_1 FILLER_30_736 ();
 sg13g2_fill_1 FILLER_30_746 ();
 sg13g2_fill_1 FILLER_30_762 ();
 sg13g2_fill_2 FILLER_30_781 ();
 sg13g2_decap_4 FILLER_30_789 ();
 sg13g2_fill_1 FILLER_30_793 ();
 sg13g2_fill_1 FILLER_30_798 ();
 sg13g2_fill_2 FILLER_30_803 ();
 sg13g2_fill_2 FILLER_30_827 ();
 sg13g2_fill_1 FILLER_30_829 ();
 sg13g2_decap_4 FILLER_30_857 ();
 sg13g2_fill_1 FILLER_30_861 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_7 ();
 sg13g2_fill_1 FILLER_31_9 ();
 sg13g2_fill_1 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_19 ();
 sg13g2_fill_2 FILLER_31_26 ();
 sg13g2_fill_2 FILLER_31_33 ();
 sg13g2_fill_1 FILLER_31_35 ();
 sg13g2_decap_4 FILLER_31_54 ();
 sg13g2_fill_2 FILLER_31_58 ();
 sg13g2_fill_2 FILLER_31_86 ();
 sg13g2_fill_1 FILLER_31_88 ();
 sg13g2_fill_2 FILLER_31_116 ();
 sg13g2_fill_1 FILLER_31_162 ();
 sg13g2_decap_4 FILLER_31_167 ();
 sg13g2_fill_1 FILLER_31_171 ();
 sg13g2_decap_8 FILLER_31_219 ();
 sg13g2_fill_2 FILLER_31_226 ();
 sg13g2_fill_1 FILLER_31_271 ();
 sg13g2_decap_4 FILLER_31_285 ();
 sg13g2_fill_1 FILLER_31_289 ();
 sg13g2_fill_2 FILLER_31_298 ();
 sg13g2_fill_1 FILLER_31_300 ();
 sg13g2_fill_2 FILLER_31_306 ();
 sg13g2_fill_1 FILLER_31_308 ();
 sg13g2_fill_1 FILLER_31_322 ();
 sg13g2_decap_4 FILLER_31_435 ();
 sg13g2_fill_2 FILLER_31_439 ();
 sg13g2_fill_2 FILLER_31_446 ();
 sg13g2_fill_1 FILLER_31_448 ();
 sg13g2_decap_4 FILLER_31_510 ();
 sg13g2_fill_1 FILLER_31_514 ();
 sg13g2_fill_2 FILLER_31_541 ();
 sg13g2_decap_4 FILLER_31_551 ();
 sg13g2_fill_1 FILLER_31_555 ();
 sg13g2_decap_8 FILLER_31_565 ();
 sg13g2_fill_2 FILLER_31_572 ();
 sg13g2_fill_1 FILLER_31_574 ();
 sg13g2_fill_2 FILLER_31_588 ();
 sg13g2_fill_1 FILLER_31_680 ();
 sg13g2_fill_2 FILLER_31_690 ();
 sg13g2_decap_4 FILLER_31_724 ();
 sg13g2_fill_2 FILLER_31_768 ();
 sg13g2_fill_1 FILLER_31_770 ();
 sg13g2_fill_1 FILLER_31_798 ();
 sg13g2_fill_2 FILLER_31_831 ();
 sg13g2_fill_1 FILLER_31_833 ();
 sg13g2_decap_8 FILLER_31_847 ();
 sg13g2_decap_8 FILLER_31_854 ();
 sg13g2_fill_1 FILLER_31_861 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_9 ();
 sg13g2_fill_2 FILLER_32_51 ();
 sg13g2_fill_1 FILLER_32_53 ();
 sg13g2_fill_2 FILLER_32_95 ();
 sg13g2_fill_1 FILLER_32_97 ();
 sg13g2_decap_8 FILLER_32_111 ();
 sg13g2_decap_4 FILLER_32_118 ();
 sg13g2_fill_2 FILLER_32_122 ();
 sg13g2_fill_1 FILLER_32_128 ();
 sg13g2_fill_2 FILLER_32_142 ();
 sg13g2_decap_4 FILLER_32_180 ();
 sg13g2_fill_2 FILLER_32_184 ();
 sg13g2_fill_1 FILLER_32_194 ();
 sg13g2_fill_1 FILLER_32_200 ();
 sg13g2_fill_1 FILLER_32_249 ();
 sg13g2_decap_4 FILLER_32_254 ();
 sg13g2_fill_2 FILLER_32_289 ();
 sg13g2_fill_1 FILLER_32_330 ();
 sg13g2_decap_4 FILLER_32_344 ();
 sg13g2_fill_2 FILLER_32_362 ();
 sg13g2_decap_8 FILLER_32_400 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_4 FILLER_32_422 ();
 sg13g2_fill_1 FILLER_32_430 ();
 sg13g2_fill_2 FILLER_32_436 ();
 sg13g2_decap_4 FILLER_32_486 ();
 sg13g2_fill_1 FILLER_32_490 ();
 sg13g2_decap_4 FILLER_32_495 ();
 sg13g2_fill_2 FILLER_32_499 ();
 sg13g2_fill_2 FILLER_32_507 ();
 sg13g2_fill_1 FILLER_32_509 ();
 sg13g2_fill_1 FILLER_32_523 ();
 sg13g2_fill_1 FILLER_32_537 ();
 sg13g2_fill_2 FILLER_32_565 ();
 sg13g2_fill_2 FILLER_32_643 ();
 sg13g2_decap_8 FILLER_32_649 ();
 sg13g2_fill_2 FILLER_32_656 ();
 sg13g2_fill_2 FILLER_32_664 ();
 sg13g2_fill_1 FILLER_32_666 ();
 sg13g2_decap_8 FILLER_32_721 ();
 sg13g2_decap_4 FILLER_32_728 ();
 sg13g2_fill_1 FILLER_32_732 ();
 sg13g2_decap_8 FILLER_32_737 ();
 sg13g2_decap_8 FILLER_32_744 ();
 sg13g2_fill_2 FILLER_32_751 ();
 sg13g2_fill_1 FILLER_32_753 ();
 sg13g2_fill_2 FILLER_32_758 ();
 sg13g2_fill_1 FILLER_32_764 ();
 sg13g2_fill_1 FILLER_32_782 ();
 sg13g2_decap_4 FILLER_32_792 ();
 sg13g2_fill_2 FILLER_32_801 ();
 sg13g2_fill_1 FILLER_32_803 ();
 sg13g2_decap_4 FILLER_32_830 ();
 sg13g2_fill_1 FILLER_32_834 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_51 ();
 sg13g2_fill_1 FILLER_33_58 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_4 FILLER_33_70 ();
 sg13g2_fill_1 FILLER_33_74 ();
 sg13g2_fill_2 FILLER_33_134 ();
 sg13g2_decap_4 FILLER_33_181 ();
 sg13g2_fill_1 FILLER_33_185 ();
 sg13g2_decap_4 FILLER_33_218 ();
 sg13g2_fill_1 FILLER_33_222 ();
 sg13g2_fill_1 FILLER_33_269 ();
 sg13g2_fill_2 FILLER_33_310 ();
 sg13g2_fill_1 FILLER_33_312 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_fill_1 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_33_460 ();
 sg13g2_decap_4 FILLER_33_516 ();
 sg13g2_fill_1 FILLER_33_520 ();
 sg13g2_decap_4 FILLER_33_547 ();
 sg13g2_fill_1 FILLER_33_564 ();
 sg13g2_decap_4 FILLER_33_583 ();
 sg13g2_fill_2 FILLER_33_587 ();
 sg13g2_fill_1 FILLER_33_593 ();
 sg13g2_fill_1 FILLER_33_620 ();
 sg13g2_decap_8 FILLER_33_648 ();
 sg13g2_fill_2 FILLER_33_661 ();
 sg13g2_fill_1 FILLER_33_663 ();
 sg13g2_fill_2 FILLER_33_669 ();
 sg13g2_fill_1 FILLER_33_671 ();
 sg13g2_fill_2 FILLER_33_676 ();
 sg13g2_fill_2 FILLER_33_710 ();
 sg13g2_fill_1 FILLER_33_712 ();
 sg13g2_decap_8 FILLER_33_740 ();
 sg13g2_decap_4 FILLER_33_747 ();
 sg13g2_fill_1 FILLER_33_751 ();
 sg13g2_fill_2 FILLER_33_790 ();
 sg13g2_fill_1 FILLER_33_824 ();
 sg13g2_fill_1 FILLER_33_834 ();
 sg13g2_decap_4 FILLER_33_857 ();
 sg13g2_fill_1 FILLER_33_861 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_4 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_4 FILLER_34_28 ();
 sg13g2_fill_1 FILLER_34_32 ();
 sg13g2_decap_8 FILLER_34_47 ();
 sg13g2_decap_4 FILLER_34_76 ();
 sg13g2_fill_2 FILLER_34_98 ();
 sg13g2_fill_1 FILLER_34_100 ();
 sg13g2_fill_2 FILLER_34_105 ();
 sg13g2_fill_1 FILLER_34_156 ();
 sg13g2_fill_2 FILLER_34_193 ();
 sg13g2_fill_2 FILLER_34_205 ();
 sg13g2_fill_1 FILLER_34_207 ();
 sg13g2_fill_2 FILLER_34_213 ();
 sg13g2_decap_4 FILLER_34_219 ();
 sg13g2_fill_1 FILLER_34_223 ();
 sg13g2_decap_8 FILLER_34_228 ();
 sg13g2_decap_4 FILLER_34_248 ();
 sg13g2_decap_4 FILLER_34_258 ();
 sg13g2_fill_2 FILLER_34_275 ();
 sg13g2_fill_1 FILLER_34_277 ();
 sg13g2_decap_4 FILLER_34_371 ();
 sg13g2_decap_8 FILLER_34_419 ();
 sg13g2_fill_1 FILLER_34_426 ();
 sg13g2_decap_4 FILLER_34_469 ();
 sg13g2_fill_2 FILLER_34_473 ();
 sg13g2_decap_8 FILLER_34_493 ();
 sg13g2_decap_4 FILLER_34_500 ();
 sg13g2_fill_2 FILLER_34_504 ();
 sg13g2_fill_1 FILLER_34_511 ();
 sg13g2_fill_2 FILLER_34_516 ();
 sg13g2_decap_4 FILLER_34_549 ();
 sg13g2_fill_1 FILLER_34_584 ();
 sg13g2_decap_4 FILLER_34_621 ();
 sg13g2_decap_8 FILLER_34_666 ();
 sg13g2_fill_1 FILLER_34_673 ();
 sg13g2_fill_2 FILLER_34_679 ();
 sg13g2_fill_2 FILLER_34_685 ();
 sg13g2_fill_2 FILLER_34_700 ();
 sg13g2_fill_2 FILLER_34_733 ();
 sg13g2_fill_1 FILLER_34_761 ();
 sg13g2_fill_2 FILLER_34_774 ();
 sg13g2_fill_1 FILLER_34_785 ();
 sg13g2_fill_2 FILLER_34_792 ();
 sg13g2_fill_1 FILLER_34_794 ();
 sg13g2_decap_4 FILLER_34_799 ();
 sg13g2_fill_2 FILLER_34_820 ();
 sg13g2_fill_1 FILLER_34_822 ();
 sg13g2_fill_1 FILLER_34_828 ();
 sg13g2_decap_4 FILLER_34_856 ();
 sg13g2_fill_2 FILLER_34_860 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_4 ();
 sg13g2_fill_2 FILLER_35_41 ();
 sg13g2_fill_1 FILLER_35_43 ();
 sg13g2_fill_1 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_54 ();
 sg13g2_fill_2 FILLER_35_61 ();
 sg13g2_fill_1 FILLER_35_90 ();
 sg13g2_fill_1 FILLER_35_100 ();
 sg13g2_decap_4 FILLER_35_106 ();
 sg13g2_fill_2 FILLER_35_110 ();
 sg13g2_fill_2 FILLER_35_135 ();
 sg13g2_fill_2 FILLER_35_181 ();
 sg13g2_fill_1 FILLER_35_183 ();
 sg13g2_fill_2 FILLER_35_207 ();
 sg13g2_decap_8 FILLER_35_236 ();
 sg13g2_fill_1 FILLER_35_243 ();
 sg13g2_decap_4 FILLER_35_324 ();
 sg13g2_fill_2 FILLER_35_328 ();
 sg13g2_fill_2 FILLER_35_343 ();
 sg13g2_fill_1 FILLER_35_350 ();
 sg13g2_decap_4 FILLER_35_364 ();
 sg13g2_fill_1 FILLER_35_390 ();
 sg13g2_fill_2 FILLER_35_404 ();
 sg13g2_fill_2 FILLER_35_486 ();
 sg13g2_fill_1 FILLER_35_488 ();
 sg13g2_decap_4 FILLER_35_499 ();
 sg13g2_fill_2 FILLER_35_530 ();
 sg13g2_fill_2 FILLER_35_537 ();
 sg13g2_fill_1 FILLER_35_539 ();
 sg13g2_fill_1 FILLER_35_574 ();
 sg13g2_fill_1 FILLER_35_579 ();
 sg13g2_fill_2 FILLER_35_593 ();
 sg13g2_decap_4 FILLER_35_599 ();
 sg13g2_decap_4 FILLER_35_612 ();
 sg13g2_fill_2 FILLER_35_624 ();
 sg13g2_fill_1 FILLER_35_649 ();
 sg13g2_decap_4 FILLER_35_664 ();
 sg13g2_fill_1 FILLER_35_715 ();
 sg13g2_decap_4 FILLER_35_720 ();
 sg13g2_decap_8 FILLER_35_742 ();
 sg13g2_fill_2 FILLER_35_749 ();
 sg13g2_fill_1 FILLER_35_751 ();
 sg13g2_decap_8 FILLER_35_826 ();
 sg13g2_decap_8 FILLER_35_850 ();
 sg13g2_decap_4 FILLER_35_857 ();
 sg13g2_fill_1 FILLER_35_861 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_12 ();
 sg13g2_fill_2 FILLER_36_19 ();
 sg13g2_fill_1 FILLER_36_21 ();
 sg13g2_fill_2 FILLER_36_76 ();
 sg13g2_fill_2 FILLER_36_83 ();
 sg13g2_fill_1 FILLER_36_90 ();
 sg13g2_fill_2 FILLER_36_96 ();
 sg13g2_fill_1 FILLER_36_98 ();
 sg13g2_decap_4 FILLER_36_103 ();
 sg13g2_fill_2 FILLER_36_107 ();
 sg13g2_fill_2 FILLER_36_150 ();
 sg13g2_fill_2 FILLER_36_184 ();
 sg13g2_fill_2 FILLER_36_200 ();
 sg13g2_fill_1 FILLER_36_202 ();
 sg13g2_fill_1 FILLER_36_211 ();
 sg13g2_fill_2 FILLER_36_253 ();
 sg13g2_fill_1 FILLER_36_255 ();
 sg13g2_decap_4 FILLER_36_261 ();
 sg13g2_fill_2 FILLER_36_265 ();
 sg13g2_fill_2 FILLER_36_278 ();
 sg13g2_fill_1 FILLER_36_280 ();
 sg13g2_fill_2 FILLER_36_304 ();
 sg13g2_fill_1 FILLER_36_306 ();
 sg13g2_fill_2 FILLER_36_355 ();
 sg13g2_fill_1 FILLER_36_357 ();
 sg13g2_decap_8 FILLER_36_376 ();
 sg13g2_fill_2 FILLER_36_383 ();
 sg13g2_fill_1 FILLER_36_385 ();
 sg13g2_fill_1 FILLER_36_391 ();
 sg13g2_fill_1 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_36_446 ();
 sg13g2_decap_4 FILLER_36_453 ();
 sg13g2_fill_2 FILLER_36_457 ();
 sg13g2_decap_4 FILLER_36_512 ();
 sg13g2_fill_2 FILLER_36_539 ();
 sg13g2_fill_1 FILLER_36_587 ();
 sg13g2_fill_1 FILLER_36_615 ();
 sg13g2_fill_1 FILLER_36_652 ();
 sg13g2_fill_2 FILLER_36_685 ();
 sg13g2_fill_1 FILLER_36_691 ();
 sg13g2_decap_4 FILLER_36_707 ();
 sg13g2_fill_1 FILLER_36_765 ();
 sg13g2_decap_4 FILLER_36_770 ();
 sg13g2_fill_1 FILLER_36_774 ();
 sg13g2_fill_2 FILLER_36_796 ();
 sg13g2_fill_1 FILLER_36_798 ();
 sg13g2_decap_4 FILLER_36_817 ();
 sg13g2_fill_2 FILLER_36_821 ();
 sg13g2_fill_2 FILLER_36_859 ();
 sg13g2_fill_1 FILLER_36_861 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_2 ();
 sg13g2_fill_1 FILLER_37_44 ();
 sg13g2_fill_2 FILLER_37_87 ();
 sg13g2_fill_2 FILLER_37_125 ();
 sg13g2_fill_2 FILLER_37_141 ();
 sg13g2_fill_2 FILLER_37_174 ();
 sg13g2_fill_2 FILLER_37_216 ();
 sg13g2_decap_8 FILLER_37_237 ();
 sg13g2_fill_2 FILLER_37_271 ();
 sg13g2_fill_1 FILLER_37_273 ();
 sg13g2_fill_1 FILLER_37_290 ();
 sg13g2_fill_2 FILLER_37_344 ();
 sg13g2_fill_2 FILLER_37_372 ();
 sg13g2_decap_8 FILLER_37_397 ();
 sg13g2_decap_4 FILLER_37_404 ();
 sg13g2_decap_4 FILLER_37_452 ();
 sg13g2_fill_2 FILLER_37_456 ();
 sg13g2_fill_2 FILLER_37_485 ();
 sg13g2_decap_4 FILLER_37_496 ();
 sg13g2_fill_2 FILLER_37_500 ();
 sg13g2_decap_8 FILLER_37_512 ();
 sg13g2_decap_4 FILLER_37_519 ();
 sg13g2_fill_1 FILLER_37_523 ();
 sg13g2_decap_8 FILLER_37_551 ();
 sg13g2_decap_8 FILLER_37_558 ();
 sg13g2_decap_4 FILLER_37_593 ();
 sg13g2_fill_1 FILLER_37_597 ();
 sg13g2_decap_8 FILLER_37_630 ();
 sg13g2_decap_8 FILLER_37_637 ();
 sg13g2_decap_8 FILLER_37_644 ();
 sg13g2_fill_1 FILLER_37_651 ();
 sg13g2_fill_2 FILLER_37_669 ();
 sg13g2_fill_1 FILLER_37_706 ();
 sg13g2_decap_8 FILLER_37_712 ();
 sg13g2_decap_8 FILLER_37_719 ();
 sg13g2_fill_1 FILLER_37_726 ();
 sg13g2_decap_4 FILLER_37_731 ();
 sg13g2_fill_2 FILLER_37_743 ();
 sg13g2_fill_1 FILLER_37_745 ();
 sg13g2_decap_4 FILLER_37_755 ();
 sg13g2_fill_2 FILLER_37_759 ();
 sg13g2_fill_2 FILLER_37_799 ();
 sg13g2_decap_4 FILLER_37_828 ();
 sg13g2_decap_8 FILLER_37_845 ();
 sg13g2_decap_8 FILLER_37_852 ();
 sg13g2_fill_2 FILLER_37_859 ();
 sg13g2_fill_1 FILLER_37_861 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_34 ();
 sg13g2_fill_2 FILLER_38_44 ();
 sg13g2_fill_1 FILLER_38_46 ();
 sg13g2_decap_4 FILLER_38_64 ();
 sg13g2_fill_2 FILLER_38_73 ();
 sg13g2_fill_1 FILLER_38_75 ();
 sg13g2_fill_1 FILLER_38_89 ();
 sg13g2_fill_2 FILLER_38_98 ();
 sg13g2_fill_1 FILLER_38_118 ();
 sg13g2_fill_2 FILLER_38_150 ();
 sg13g2_fill_1 FILLER_38_199 ();
 sg13g2_decap_8 FILLER_38_227 ();
 sg13g2_fill_1 FILLER_38_234 ();
 sg13g2_fill_1 FILLER_38_267 ();
 sg13g2_fill_2 FILLER_38_272 ();
 sg13g2_fill_2 FILLER_38_287 ();
 sg13g2_fill_1 FILLER_38_289 ();
 sg13g2_decap_8 FILLER_38_307 ();
 sg13g2_decap_8 FILLER_38_314 ();
 sg13g2_decap_4 FILLER_38_321 ();
 sg13g2_decap_8 FILLER_38_343 ();
 sg13g2_fill_2 FILLER_38_368 ();
 sg13g2_fill_1 FILLER_38_399 ();
 sg13g2_decap_8 FILLER_38_413 ();
 sg13g2_fill_2 FILLER_38_420 ();
 sg13g2_fill_2 FILLER_38_448 ();
 sg13g2_decap_4 FILLER_38_481 ();
 sg13g2_fill_2 FILLER_38_503 ();
 sg13g2_fill_2 FILLER_38_514 ();
 sg13g2_fill_1 FILLER_38_516 ();
 sg13g2_decap_4 FILLER_38_522 ();
 sg13g2_fill_1 FILLER_38_526 ();
 sg13g2_fill_2 FILLER_38_561 ();
 sg13g2_fill_2 FILLER_38_577 ();
 sg13g2_fill_1 FILLER_38_579 ();
 sg13g2_decap_4 FILLER_38_596 ();
 sg13g2_fill_1 FILLER_38_600 ();
 sg13g2_decap_4 FILLER_38_633 ();
 sg13g2_fill_1 FILLER_38_673 ();
 sg13g2_decap_4 FILLER_38_706 ();
 sg13g2_fill_1 FILLER_38_715 ();
 sg13g2_decap_4 FILLER_38_724 ();
 sg13g2_decap_8 FILLER_38_781 ();
 sg13g2_decap_8 FILLER_38_788 ();
 sg13g2_fill_2 FILLER_38_795 ();
 sg13g2_fill_2 FILLER_38_801 ();
 sg13g2_fill_1 FILLER_38_803 ();
 sg13g2_decap_4 FILLER_38_857 ();
 sg13g2_fill_1 FILLER_38_861 ();
 sg13g2_decap_4 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_4 ();
 sg13g2_fill_2 FILLER_39_10 ();
 sg13g2_decap_4 FILLER_39_16 ();
 sg13g2_fill_1 FILLER_39_49 ();
 sg13g2_fill_2 FILLER_39_82 ();
 sg13g2_fill_1 FILLER_39_137 ();
 sg13g2_fill_2 FILLER_39_155 ();
 sg13g2_fill_1 FILLER_39_157 ();
 sg13g2_fill_2 FILLER_39_197 ();
 sg13g2_fill_1 FILLER_39_199 ();
 sg13g2_fill_1 FILLER_39_213 ();
 sg13g2_decap_8 FILLER_39_233 ();
 sg13g2_fill_2 FILLER_39_240 ();
 sg13g2_decap_8 FILLER_39_260 ();
 sg13g2_fill_1 FILLER_39_267 ();
 sg13g2_decap_8 FILLER_39_277 ();
 sg13g2_decap_4 FILLER_39_284 ();
 sg13g2_decap_4 FILLER_39_315 ();
 sg13g2_fill_1 FILLER_39_319 ();
 sg13g2_decap_8 FILLER_39_350 ();
 sg13g2_fill_2 FILLER_39_357 ();
 sg13g2_decap_8 FILLER_39_364 ();
 sg13g2_decap_8 FILLER_39_371 ();
 sg13g2_fill_2 FILLER_39_378 ();
 sg13g2_fill_1 FILLER_39_380 ();
 sg13g2_decap_8 FILLER_39_394 ();
 sg13g2_fill_2 FILLER_39_401 ();
 sg13g2_decap_4 FILLER_39_455 ();
 sg13g2_fill_1 FILLER_39_463 ();
 sg13g2_decap_8 FILLER_39_477 ();
 sg13g2_decap_4 FILLER_39_484 ();
 sg13g2_fill_2 FILLER_39_488 ();
 sg13g2_fill_1 FILLER_39_517 ();
 sg13g2_decap_4 FILLER_39_539 ();
 sg13g2_fill_2 FILLER_39_543 ();
 sg13g2_fill_1 FILLER_39_581 ();
 sg13g2_fill_1 FILLER_39_614 ();
 sg13g2_decap_4 FILLER_39_646 ();
 sg13g2_fill_1 FILLER_39_650 ();
 sg13g2_decap_4 FILLER_39_655 ();
 sg13g2_fill_2 FILLER_39_659 ();
 sg13g2_fill_2 FILLER_39_665 ();
 sg13g2_decap_8 FILLER_39_672 ();
 sg13g2_fill_2 FILLER_39_684 ();
 sg13g2_decap_8 FILLER_39_694 ();
 sg13g2_decap_4 FILLER_39_701 ();
 sg13g2_fill_2 FILLER_39_741 ();
 sg13g2_fill_1 FILLER_39_743 ();
 sg13g2_fill_1 FILLER_39_766 ();
 sg13g2_fill_2 FILLER_39_803 ();
 sg13g2_fill_1 FILLER_39_818 ();
 sg13g2_decap_8 FILLER_39_837 ();
 sg13g2_decap_8 FILLER_39_844 ();
 sg13g2_decap_8 FILLER_39_851 ();
 sg13g2_decap_4 FILLER_39_858 ();
 sg13g2_fill_1 FILLER_40_0 ();
 sg13g2_decap_4 FILLER_40_45 ();
 sg13g2_decap_4 FILLER_40_66 ();
 sg13g2_fill_1 FILLER_40_70 ();
 sg13g2_decap_4 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_101 ();
 sg13g2_decap_4 FILLER_40_108 ();
 sg13g2_fill_1 FILLER_40_126 ();
 sg13g2_fill_2 FILLER_40_136 ();
 sg13g2_fill_1 FILLER_40_183 ();
 sg13g2_fill_2 FILLER_40_252 ();
 sg13g2_fill_1 FILLER_40_286 ();
 sg13g2_fill_1 FILLER_40_297 ();
 sg13g2_fill_2 FILLER_40_324 ();
 sg13g2_decap_8 FILLER_40_363 ();
 sg13g2_fill_2 FILLER_40_374 ();
 sg13g2_fill_1 FILLER_40_376 ();
 sg13g2_decap_4 FILLER_40_382 ();
 sg13g2_fill_2 FILLER_40_386 ();
 sg13g2_decap_8 FILLER_40_401 ();
 sg13g2_fill_1 FILLER_40_413 ();
 sg13g2_fill_2 FILLER_40_427 ();
 sg13g2_decap_8 FILLER_40_469 ();
 sg13g2_fill_2 FILLER_40_476 ();
 sg13g2_fill_1 FILLER_40_478 ();
 sg13g2_fill_1 FILLER_40_506 ();
 sg13g2_fill_2 FILLER_40_512 ();
 sg13g2_fill_2 FILLER_40_523 ();
 sg13g2_fill_1 FILLER_40_525 ();
 sg13g2_fill_2 FILLER_40_539 ();
 sg13g2_decap_8 FILLER_40_553 ();
 sg13g2_decap_8 FILLER_40_560 ();
 sg13g2_fill_2 FILLER_40_567 ();
 sg13g2_fill_1 FILLER_40_569 ();
 sg13g2_decap_8 FILLER_40_575 ();
 sg13g2_fill_2 FILLER_40_582 ();
 sg13g2_fill_1 FILLER_40_584 ();
 sg13g2_fill_2 FILLER_40_589 ();
 sg13g2_fill_1 FILLER_40_617 ();
 sg13g2_decap_8 FILLER_40_631 ();
 sg13g2_fill_2 FILLER_40_638 ();
 sg13g2_decap_8 FILLER_40_716 ();
 sg13g2_decap_8 FILLER_40_723 ();
 sg13g2_fill_1 FILLER_40_730 ();
 sg13g2_fill_1 FILLER_40_736 ();
 sg13g2_fill_1 FILLER_40_741 ();
 sg13g2_fill_2 FILLER_40_748 ();
 sg13g2_fill_1 FILLER_40_750 ();
 sg13g2_decap_4 FILLER_40_785 ();
 sg13g2_decap_8 FILLER_40_804 ();
 sg13g2_decap_4 FILLER_40_811 ();
 sg13g2_decap_8 FILLER_40_842 ();
 sg13g2_decap_8 FILLER_40_849 ();
 sg13g2_decap_4 FILLER_40_856 ();
 sg13g2_fill_2 FILLER_40_860 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_7 ();
 sg13g2_decap_4 FILLER_41_13 ();
 sg13g2_fill_2 FILLER_41_39 ();
 sg13g2_fill_1 FILLER_41_41 ();
 sg13g2_fill_2 FILLER_41_47 ();
 sg13g2_decap_8 FILLER_41_53 ();
 sg13g2_decap_8 FILLER_41_60 ();
 sg13g2_fill_1 FILLER_41_67 ();
 sg13g2_decap_8 FILLER_41_73 ();
 sg13g2_fill_1 FILLER_41_80 ();
 sg13g2_decap_4 FILLER_41_104 ();
 sg13g2_fill_2 FILLER_41_135 ();
 sg13g2_fill_1 FILLER_41_137 ();
 sg13g2_fill_2 FILLER_41_156 ();
 sg13g2_fill_1 FILLER_41_158 ();
 sg13g2_decap_8 FILLER_41_163 ();
 sg13g2_fill_1 FILLER_41_170 ();
 sg13g2_decap_4 FILLER_41_176 ();
 sg13g2_fill_1 FILLER_41_180 ();
 sg13g2_decap_4 FILLER_41_202 ();
 sg13g2_fill_2 FILLER_41_206 ();
 sg13g2_decap_4 FILLER_41_217 ();
 sg13g2_decap_8 FILLER_41_227 ();
 sg13g2_decap_4 FILLER_41_234 ();
 sg13g2_fill_1 FILLER_41_247 ();
 sg13g2_fill_1 FILLER_41_281 ();
 sg13g2_fill_2 FILLER_41_287 ();
 sg13g2_decap_4 FILLER_41_302 ();
 sg13g2_fill_1 FILLER_41_306 ();
 sg13g2_decap_4 FILLER_41_312 ();
 sg13g2_fill_1 FILLER_41_316 ();
 sg13g2_decap_8 FILLER_41_321 ();
 sg13g2_fill_1 FILLER_41_328 ();
 sg13g2_fill_1 FILLER_41_353 ();
 sg13g2_fill_1 FILLER_41_358 ();
 sg13g2_fill_2 FILLER_41_372 ();
 sg13g2_fill_2 FILLER_41_401 ();
 sg13g2_fill_1 FILLER_41_403 ();
 sg13g2_decap_8 FILLER_41_436 ();
 sg13g2_decap_4 FILLER_41_443 ();
 sg13g2_decap_4 FILLER_41_451 ();
 sg13g2_decap_4 FILLER_41_465 ();
 sg13g2_fill_1 FILLER_41_478 ();
 sg13g2_fill_2 FILLER_41_493 ();
 sg13g2_fill_2 FILLER_41_525 ();
 sg13g2_fill_2 FILLER_41_558 ();
 sg13g2_fill_1 FILLER_41_560 ();
 sg13g2_decap_8 FILLER_41_638 ();
 sg13g2_fill_1 FILLER_41_645 ();
 sg13g2_decap_8 FILLER_41_650 ();
 sg13g2_decap_4 FILLER_41_657 ();
 sg13g2_fill_2 FILLER_41_667 ();
 sg13g2_fill_1 FILLER_41_669 ();
 sg13g2_fill_2 FILLER_41_679 ();
 sg13g2_decap_8 FILLER_41_685 ();
 sg13g2_decap_8 FILLER_41_692 ();
 sg13g2_fill_2 FILLER_41_717 ();
 sg13g2_fill_1 FILLER_41_719 ();
 sg13g2_fill_2 FILLER_41_760 ();
 sg13g2_decap_8 FILLER_41_789 ();
 sg13g2_decap_4 FILLER_41_796 ();
 sg13g2_decap_8 FILLER_41_836 ();
 sg13g2_decap_8 FILLER_41_843 ();
 sg13g2_decap_8 FILLER_41_850 ();
 sg13g2_decap_4 FILLER_41_857 ();
 sg13g2_fill_1 FILLER_41_861 ();
 sg13g2_decap_4 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_31 ();
 sg13g2_fill_1 FILLER_42_33 ();
 sg13g2_fill_1 FILLER_42_83 ();
 sg13g2_decap_4 FILLER_42_89 ();
 sg13g2_fill_1 FILLER_42_93 ();
 sg13g2_decap_8 FILLER_42_99 ();
 sg13g2_decap_8 FILLER_42_123 ();
 sg13g2_fill_1 FILLER_42_130 ();
 sg13g2_decap_8 FILLER_42_135 ();
 sg13g2_decap_8 FILLER_42_142 ();
 sg13g2_decap_4 FILLER_42_149 ();
 sg13g2_fill_1 FILLER_42_153 ();
 sg13g2_fill_1 FILLER_42_232 ();
 sg13g2_fill_1 FILLER_42_246 ();
 sg13g2_fill_1 FILLER_42_260 ();
 sg13g2_fill_2 FILLER_42_288 ();
 sg13g2_fill_2 FILLER_42_294 ();
 sg13g2_decap_4 FILLER_42_305 ();
 sg13g2_decap_4 FILLER_42_345 ();
 sg13g2_fill_1 FILLER_42_376 ();
 sg13g2_fill_2 FILLER_42_411 ();
 sg13g2_fill_1 FILLER_42_413 ();
 sg13g2_fill_2 FILLER_42_418 ();
 sg13g2_fill_1 FILLER_42_420 ();
 sg13g2_decap_4 FILLER_42_470 ();
 sg13g2_fill_1 FILLER_42_494 ();
 sg13g2_fill_2 FILLER_42_505 ();
 sg13g2_fill_2 FILLER_42_548 ();
 sg13g2_decap_4 FILLER_42_577 ();
 sg13g2_fill_2 FILLER_42_600 ();
 sg13g2_fill_1 FILLER_42_602 ();
 sg13g2_decap_4 FILLER_42_612 ();
 sg13g2_fill_2 FILLER_42_620 ();
 sg13g2_fill_1 FILLER_42_622 ();
 sg13g2_decap_8 FILLER_42_632 ();
 sg13g2_fill_1 FILLER_42_683 ();
 sg13g2_fill_2 FILLER_42_688 ();
 sg13g2_fill_1 FILLER_42_690 ();
 sg13g2_decap_8 FILLER_42_709 ();
 sg13g2_decap_4 FILLER_42_716 ();
 sg13g2_fill_2 FILLER_42_720 ();
 sg13g2_decap_8 FILLER_42_731 ();
 sg13g2_decap_8 FILLER_42_747 ();
 sg13g2_fill_2 FILLER_42_754 ();
 sg13g2_fill_1 FILLER_42_756 ();
 sg13g2_fill_1 FILLER_42_763 ();
 sg13g2_decap_4 FILLER_42_768 ();
 sg13g2_fill_1 FILLER_42_772 ();
 sg13g2_fill_2 FILLER_42_783 ();
 sg13g2_fill_1 FILLER_42_785 ();
 sg13g2_fill_2 FILLER_42_790 ();
 sg13g2_fill_1 FILLER_42_792 ();
 sg13g2_fill_2 FILLER_42_802 ();
 sg13g2_fill_1 FILLER_42_817 ();
 sg13g2_decap_8 FILLER_42_831 ();
 sg13g2_decap_8 FILLER_42_838 ();
 sg13g2_decap_8 FILLER_42_845 ();
 sg13g2_decap_8 FILLER_42_852 ();
 sg13g2_fill_2 FILLER_42_859 ();
 sg13g2_fill_1 FILLER_42_861 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_7 ();
 sg13g2_fill_2 FILLER_43_36 ();
 sg13g2_fill_1 FILLER_43_38 ();
 sg13g2_fill_1 FILLER_43_57 ();
 sg13g2_fill_2 FILLER_43_72 ();
 sg13g2_fill_1 FILLER_43_74 ();
 sg13g2_fill_2 FILLER_43_89 ();
 sg13g2_fill_1 FILLER_43_91 ();
 sg13g2_fill_1 FILLER_43_101 ();
 sg13g2_decap_4 FILLER_43_106 ();
 sg13g2_fill_2 FILLER_43_110 ();
 sg13g2_fill_2 FILLER_43_130 ();
 sg13g2_fill_1 FILLER_43_132 ();
 sg13g2_decap_4 FILLER_43_162 ();
 sg13g2_fill_1 FILLER_43_166 ();
 sg13g2_decap_8 FILLER_43_173 ();
 sg13g2_fill_2 FILLER_43_180 ();
 sg13g2_fill_1 FILLER_43_182 ();
 sg13g2_fill_2 FILLER_43_188 ();
 sg13g2_fill_1 FILLER_43_190 ();
 sg13g2_decap_4 FILLER_43_199 ();
 sg13g2_fill_2 FILLER_43_203 ();
 sg13g2_fill_2 FILLER_43_321 ();
 sg13g2_fill_1 FILLER_43_323 ();
 sg13g2_decap_8 FILLER_43_346 ();
 sg13g2_fill_1 FILLER_43_353 ();
 sg13g2_fill_2 FILLER_43_385 ();
 sg13g2_fill_1 FILLER_43_387 ();
 sg13g2_fill_1 FILLER_43_430 ();
 sg13g2_decap_8 FILLER_43_440 ();
 sg13g2_fill_2 FILLER_43_462 ();
 sg13g2_fill_1 FILLER_43_464 ();
 sg13g2_fill_2 FILLER_43_503 ();
 sg13g2_decap_4 FILLER_43_518 ();
 sg13g2_fill_1 FILLER_43_522 ();
 sg13g2_fill_1 FILLER_43_532 ();
 sg13g2_fill_2 FILLER_43_556 ();
 sg13g2_fill_1 FILLER_43_558 ();
 sg13g2_decap_4 FILLER_43_568 ();
 sg13g2_fill_1 FILLER_43_572 ();
 sg13g2_decap_4 FILLER_43_581 ();
 sg13g2_decap_8 FILLER_43_588 ();
 sg13g2_fill_1 FILLER_43_595 ();
 sg13g2_fill_2 FILLER_43_649 ();
 sg13g2_fill_2 FILLER_43_660 ();
 sg13g2_fill_1 FILLER_43_668 ();
 sg13g2_fill_2 FILLER_43_773 ();
 sg13g2_fill_2 FILLER_43_807 ();
 sg13g2_decap_8 FILLER_43_841 ();
 sg13g2_decap_8 FILLER_43_848 ();
 sg13g2_decap_8 FILLER_43_855 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_18 ();
 sg13g2_fill_2 FILLER_44_25 ();
 sg13g2_fill_1 FILLER_44_27 ();
 sg13g2_fill_1 FILLER_44_86 ();
 sg13g2_decap_4 FILLER_44_114 ();
 sg13g2_fill_2 FILLER_44_145 ();
 sg13g2_fill_1 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_166 ();
 sg13g2_fill_1 FILLER_44_173 ();
 sg13g2_fill_2 FILLER_44_219 ();
 sg13g2_fill_1 FILLER_44_221 ();
 sg13g2_fill_2 FILLER_44_249 ();
 sg13g2_fill_2 FILLER_44_260 ();
 sg13g2_fill_1 FILLER_44_262 ();
 sg13g2_fill_2 FILLER_44_284 ();
 sg13g2_fill_1 FILLER_44_301 ();
 sg13g2_fill_1 FILLER_44_311 ();
 sg13g2_fill_2 FILLER_44_317 ();
 sg13g2_decap_4 FILLER_44_328 ();
 sg13g2_fill_1 FILLER_44_332 ();
 sg13g2_fill_2 FILLER_44_351 ();
 sg13g2_fill_2 FILLER_44_393 ();
 sg13g2_fill_1 FILLER_44_395 ();
 sg13g2_fill_1 FILLER_44_402 ();
 sg13g2_fill_1 FILLER_44_407 ();
 sg13g2_fill_1 FILLER_44_412 ();
 sg13g2_fill_2 FILLER_44_426 ();
 sg13g2_fill_1 FILLER_44_428 ();
 sg13g2_decap_8 FILLER_44_442 ();
 sg13g2_decap_8 FILLER_44_449 ();
 sg13g2_decap_8 FILLER_44_456 ();
 sg13g2_fill_2 FILLER_44_463 ();
 sg13g2_decap_4 FILLER_44_482 ();
 sg13g2_fill_2 FILLER_44_513 ();
 sg13g2_fill_1 FILLER_44_515 ();
 sg13g2_fill_1 FILLER_44_521 ();
 sg13g2_fill_2 FILLER_44_540 ();
 sg13g2_fill_1 FILLER_44_559 ();
 sg13g2_fill_1 FILLER_44_590 ();
 sg13g2_fill_2 FILLER_44_627 ();
 sg13g2_fill_1 FILLER_44_629 ();
 sg13g2_decap_8 FILLER_44_662 ();
 sg13g2_decap_4 FILLER_44_669 ();
 sg13g2_fill_1 FILLER_44_673 ();
 sg13g2_fill_1 FILLER_44_688 ();
 sg13g2_fill_1 FILLER_44_708 ();
 sg13g2_fill_2 FILLER_44_715 ();
 sg13g2_decap_4 FILLER_44_734 ();
 sg13g2_fill_1 FILLER_44_738 ();
 sg13g2_decap_4 FILLER_44_744 ();
 sg13g2_fill_2 FILLER_44_748 ();
 sg13g2_fill_1 FILLER_44_763 ();
 sg13g2_fill_2 FILLER_44_792 ();
 sg13g2_fill_1 FILLER_44_794 ();
 sg13g2_fill_2 FILLER_44_804 ();
 sg13g2_fill_1 FILLER_44_806 ();
 sg13g2_fill_2 FILLER_44_811 ();
 sg13g2_fill_2 FILLER_44_822 ();
 sg13g2_decap_8 FILLER_44_837 ();
 sg13g2_decap_8 FILLER_44_844 ();
 sg13g2_decap_8 FILLER_44_851 ();
 sg13g2_decap_4 FILLER_44_858 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_4 FILLER_45_28 ();
 sg13g2_fill_2 FILLER_45_32 ();
 sg13g2_decap_4 FILLER_45_38 ();
 sg13g2_fill_2 FILLER_45_51 ();
 sg13g2_fill_1 FILLER_45_53 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_4 FILLER_45_70 ();
 sg13g2_fill_1 FILLER_45_74 ();
 sg13g2_fill_2 FILLER_45_107 ();
 sg13g2_fill_1 FILLER_45_122 ();
 sg13g2_decap_8 FILLER_45_127 ();
 sg13g2_decap_8 FILLER_45_134 ();
 sg13g2_fill_2 FILLER_45_141 ();
 sg13g2_fill_2 FILLER_45_183 ();
 sg13g2_fill_1 FILLER_45_190 ();
 sg13g2_decap_4 FILLER_45_213 ();
 sg13g2_fill_2 FILLER_45_217 ();
 sg13g2_decap_8 FILLER_45_227 ();
 sg13g2_decap_4 FILLER_45_234 ();
 sg13g2_fill_2 FILLER_45_238 ();
 sg13g2_fill_2 FILLER_45_267 ();
 sg13g2_decap_4 FILLER_45_315 ();
 sg13g2_fill_1 FILLER_45_319 ();
 sg13g2_decap_4 FILLER_45_388 ();
 sg13g2_decap_4 FILLER_45_400 ();
 sg13g2_fill_2 FILLER_45_404 ();
 sg13g2_fill_2 FILLER_45_446 ();
 sg13g2_fill_1 FILLER_45_448 ();
 sg13g2_fill_1 FILLER_45_476 ();
 sg13g2_fill_2 FILLER_45_524 ();
 sg13g2_fill_1 FILLER_45_526 ();
 sg13g2_fill_1 FILLER_45_575 ();
 sg13g2_fill_1 FILLER_45_634 ();
 sg13g2_fill_1 FILLER_45_657 ();
 sg13g2_fill_2 FILLER_45_680 ();
 sg13g2_decap_4 FILLER_45_795 ();
 sg13g2_fill_2 FILLER_45_799 ();
 sg13g2_decap_8 FILLER_45_828 ();
 sg13g2_decap_8 FILLER_45_835 ();
 sg13g2_decap_8 FILLER_45_842 ();
 sg13g2_decap_8 FILLER_45_849 ();
 sg13g2_decap_4 FILLER_45_856 ();
 sg13g2_fill_2 FILLER_45_860 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_fill_1 FILLER_46_42 ();
 sg13g2_decap_4 FILLER_46_70 ();
 sg13g2_fill_2 FILLER_46_74 ();
 sg13g2_fill_1 FILLER_46_115 ();
 sg13g2_decap_4 FILLER_46_121 ();
 sg13g2_decap_8 FILLER_46_129 ();
 sg13g2_decap_8 FILLER_46_136 ();
 sg13g2_fill_2 FILLER_46_180 ();
 sg13g2_fill_1 FILLER_46_209 ();
 sg13g2_decap_8 FILLER_46_235 ();
 sg13g2_fill_2 FILLER_46_242 ();
 sg13g2_fill_1 FILLER_46_244 ();
 sg13g2_fill_1 FILLER_46_249 ();
 sg13g2_fill_2 FILLER_46_264 ();
 sg13g2_fill_1 FILLER_46_266 ();
 sg13g2_decap_4 FILLER_46_307 ();
 sg13g2_fill_2 FILLER_46_311 ();
 sg13g2_decap_8 FILLER_46_326 ();
 sg13g2_fill_2 FILLER_46_344 ();
 sg13g2_fill_1 FILLER_46_346 ();
 sg13g2_fill_1 FILLER_46_369 ();
 sg13g2_decap_8 FILLER_46_379 ();
 sg13g2_fill_1 FILLER_46_386 ();
 sg13g2_fill_2 FILLER_46_396 ();
 sg13g2_fill_1 FILLER_46_398 ();
 sg13g2_fill_2 FILLER_46_417 ();
 sg13g2_fill_1 FILLER_46_419 ();
 sg13g2_fill_1 FILLER_46_451 ();
 sg13g2_fill_2 FILLER_46_460 ();
 sg13g2_fill_2 FILLER_46_476 ();
 sg13g2_decap_8 FILLER_46_487 ();
 sg13g2_decap_8 FILLER_46_494 ();
 sg13g2_fill_2 FILLER_46_501 ();
 sg13g2_decap_4 FILLER_46_536 ();
 sg13g2_fill_2 FILLER_46_557 ();
 sg13g2_fill_1 FILLER_46_559 ();
 sg13g2_fill_1 FILLER_46_601 ();
 sg13g2_fill_1 FILLER_46_610 ();
 sg13g2_fill_2 FILLER_46_679 ();
 sg13g2_fill_1 FILLER_46_681 ();
 sg13g2_fill_1 FILLER_46_686 ();
 sg13g2_decap_4 FILLER_46_691 ();
 sg13g2_fill_2 FILLER_46_695 ();
 sg13g2_fill_2 FILLER_46_706 ();
 sg13g2_fill_1 FILLER_46_708 ();
 sg13g2_decap_4 FILLER_46_718 ();
 sg13g2_decap_8 FILLER_46_731 ();
 sg13g2_fill_2 FILLER_46_738 ();
 sg13g2_fill_1 FILLER_46_740 ();
 sg13g2_fill_2 FILLER_46_745 ();
 sg13g2_fill_1 FILLER_46_747 ();
 sg13g2_decap_4 FILLER_46_752 ();
 sg13g2_fill_1 FILLER_46_756 ();
 sg13g2_fill_2 FILLER_46_766 ();
 sg13g2_fill_1 FILLER_46_768 ();
 sg13g2_decap_4 FILLER_46_777 ();
 sg13g2_fill_2 FILLER_46_781 ();
 sg13g2_decap_8 FILLER_46_792 ();
 sg13g2_decap_8 FILLER_46_799 ();
 sg13g2_decap_8 FILLER_46_810 ();
 sg13g2_decap_8 FILLER_46_817 ();
 sg13g2_decap_8 FILLER_46_824 ();
 sg13g2_decap_8 FILLER_46_831 ();
 sg13g2_decap_8 FILLER_46_838 ();
 sg13g2_decap_8 FILLER_46_845 ();
 sg13g2_decap_8 FILLER_46_852 ();
 sg13g2_fill_2 FILLER_46_859 ();
 sg13g2_fill_1 FILLER_46_861 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_4 FILLER_47_42 ();
 sg13g2_fill_1 FILLER_47_46 ();
 sg13g2_decap_8 FILLER_47_55 ();
 sg13g2_fill_1 FILLER_47_62 ();
 sg13g2_fill_2 FILLER_47_99 ();
 sg13g2_fill_1 FILLER_47_101 ();
 sg13g2_decap_4 FILLER_47_159 ();
 sg13g2_fill_2 FILLER_47_163 ();
 sg13g2_decap_4 FILLER_47_212 ();
 sg13g2_fill_2 FILLER_47_216 ();
 sg13g2_decap_4 FILLER_47_228 ();
 sg13g2_fill_2 FILLER_47_232 ();
 sg13g2_decap_8 FILLER_47_238 ();
 sg13g2_fill_2 FILLER_47_245 ();
 sg13g2_fill_1 FILLER_47_247 ();
 sg13g2_fill_1 FILLER_47_257 ();
 sg13g2_fill_2 FILLER_47_267 ();
 sg13g2_fill_2 FILLER_47_305 ();
 sg13g2_fill_1 FILLER_47_307 ();
 sg13g2_decap_8 FILLER_47_330 ();
 sg13g2_fill_2 FILLER_47_337 ();
 sg13g2_fill_1 FILLER_47_339 ();
 sg13g2_fill_2 FILLER_47_363 ();
 sg13g2_decap_8 FILLER_47_374 ();
 sg13g2_fill_2 FILLER_47_381 ();
 sg13g2_fill_2 FILLER_47_401 ();
 sg13g2_decap_8 FILLER_47_436 ();
 sg13g2_decap_4 FILLER_47_443 ();
 sg13g2_fill_1 FILLER_47_474 ();
 sg13g2_fill_2 FILLER_47_510 ();
 sg13g2_fill_1 FILLER_47_512 ();
 sg13g2_fill_2 FILLER_47_517 ();
 sg13g2_decap_4 FILLER_47_532 ();
 sg13g2_fill_2 FILLER_47_536 ();
 sg13g2_fill_1 FILLER_47_543 ();
 sg13g2_fill_2 FILLER_47_548 ();
 sg13g2_fill_2 FILLER_47_572 ();
 sg13g2_fill_1 FILLER_47_601 ();
 sg13g2_decap_4 FILLER_47_615 ();
 sg13g2_fill_2 FILLER_47_619 ();
 sg13g2_decap_8 FILLER_47_625 ();
 sg13g2_decap_8 FILLER_47_632 ();
 sg13g2_decap_4 FILLER_47_639 ();
 sg13g2_fill_1 FILLER_47_643 ();
 sg13g2_decap_8 FILLER_47_648 ();
 sg13g2_decap_8 FILLER_47_655 ();
 sg13g2_decap_8 FILLER_47_689 ();
 sg13g2_decap_8 FILLER_47_696 ();
 sg13g2_decap_8 FILLER_47_703 ();
 sg13g2_decap_8 FILLER_47_710 ();
 sg13g2_decap_8 FILLER_47_717 ();
 sg13g2_decap_8 FILLER_47_724 ();
 sg13g2_decap_8 FILLER_47_731 ();
 sg13g2_decap_8 FILLER_47_738 ();
 sg13g2_decap_8 FILLER_47_745 ();
 sg13g2_decap_8 FILLER_47_752 ();
 sg13g2_decap_8 FILLER_47_759 ();
 sg13g2_decap_8 FILLER_47_766 ();
 sg13g2_decap_8 FILLER_47_773 ();
 sg13g2_decap_8 FILLER_47_780 ();
 sg13g2_decap_8 FILLER_47_787 ();
 sg13g2_decap_8 FILLER_47_794 ();
 sg13g2_decap_8 FILLER_47_801 ();
 sg13g2_decap_8 FILLER_47_808 ();
 sg13g2_decap_8 FILLER_47_815 ();
 sg13g2_decap_8 FILLER_47_822 ();
 sg13g2_decap_8 FILLER_47_829 ();
 sg13g2_decap_8 FILLER_47_836 ();
 sg13g2_decap_8 FILLER_47_843 ();
 sg13g2_decap_8 FILLER_47_850 ();
 sg13g2_decap_4 FILLER_47_857 ();
 sg13g2_fill_1 FILLER_47_861 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_4 FILLER_48_56 ();
 sg13g2_fill_2 FILLER_48_60 ();
 sg13g2_decap_8 FILLER_48_75 ();
 sg13g2_fill_1 FILLER_48_82 ();
 sg13g2_fill_1 FILLER_48_131 ();
 sg13g2_fill_1 FILLER_48_199 ();
 sg13g2_fill_2 FILLER_48_227 ();
 sg13g2_fill_2 FILLER_48_256 ();
 sg13g2_fill_1 FILLER_48_258 ();
 sg13g2_fill_2 FILLER_48_268 ();
 sg13g2_fill_2 FILLER_48_280 ();
 sg13g2_fill_1 FILLER_48_282 ();
 sg13g2_decap_8 FILLER_48_291 ();
 sg13g2_fill_1 FILLER_48_298 ();
 sg13g2_fill_1 FILLER_48_312 ();
 sg13g2_decap_4 FILLER_48_327 ();
 sg13g2_fill_2 FILLER_48_362 ();
 sg13g2_fill_1 FILLER_48_364 ();
 sg13g2_fill_1 FILLER_48_406 ();
 sg13g2_fill_2 FILLER_48_412 ();
 sg13g2_fill_1 FILLER_48_414 ();
 sg13g2_fill_2 FILLER_48_429 ();
 sg13g2_fill_1 FILLER_48_431 ();
 sg13g2_decap_4 FILLER_48_445 ();
 sg13g2_fill_2 FILLER_48_449 ();
 sg13g2_fill_2 FILLER_48_459 ();
 sg13g2_fill_1 FILLER_48_461 ();
 sg13g2_fill_2 FILLER_48_481 ();
 sg13g2_fill_2 FILLER_48_496 ();
 sg13g2_fill_1 FILLER_48_498 ();
 sg13g2_decap_8 FILLER_48_512 ();
 sg13g2_fill_2 FILLER_48_529 ();
 sg13g2_fill_2 FILLER_48_536 ();
 sg13g2_fill_1 FILLER_48_538 ();
 sg13g2_decap_8 FILLER_48_570 ();
 sg13g2_decap_8 FILLER_48_577 ();
 sg13g2_fill_2 FILLER_48_607 ();
 sg13g2_fill_1 FILLER_48_609 ();
 sg13g2_decap_8 FILLER_48_650 ();
 sg13g2_decap_8 FILLER_48_657 ();
 sg13g2_decap_4 FILLER_48_664 ();
 sg13g2_fill_2 FILLER_48_672 ();
 sg13g2_fill_1 FILLER_48_674 ();
 sg13g2_decap_8 FILLER_48_684 ();
 sg13g2_decap_8 FILLER_48_691 ();
 sg13g2_decap_8 FILLER_48_698 ();
 sg13g2_decap_8 FILLER_48_705 ();
 sg13g2_decap_8 FILLER_48_712 ();
 sg13g2_decap_8 FILLER_48_719 ();
 sg13g2_decap_8 FILLER_48_726 ();
 sg13g2_decap_8 FILLER_48_733 ();
 sg13g2_decap_8 FILLER_48_740 ();
 sg13g2_decap_8 FILLER_48_747 ();
 sg13g2_decap_8 FILLER_48_754 ();
 sg13g2_decap_8 FILLER_48_761 ();
 sg13g2_decap_8 FILLER_48_768 ();
 sg13g2_decap_8 FILLER_48_775 ();
 sg13g2_decap_8 FILLER_48_782 ();
 sg13g2_decap_8 FILLER_48_789 ();
 sg13g2_decap_8 FILLER_48_796 ();
 sg13g2_decap_8 FILLER_48_803 ();
 sg13g2_decap_8 FILLER_48_810 ();
 sg13g2_decap_8 FILLER_48_817 ();
 sg13g2_decap_8 FILLER_48_824 ();
 sg13g2_decap_8 FILLER_48_831 ();
 sg13g2_decap_8 FILLER_48_838 ();
 sg13g2_decap_8 FILLER_48_845 ();
 sg13g2_decap_8 FILLER_48_852 ();
 sg13g2_fill_2 FILLER_48_859 ();
 sg13g2_fill_1 FILLER_48_861 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_4 FILLER_49_84 ();
 sg13g2_decap_4 FILLER_49_92 ();
 sg13g2_fill_2 FILLER_49_96 ();
 sg13g2_fill_2 FILLER_49_175 ();
 sg13g2_fill_1 FILLER_49_177 ();
 sg13g2_decap_8 FILLER_49_182 ();
 sg13g2_fill_1 FILLER_49_189 ();
 sg13g2_decap_4 FILLER_49_199 ();
 sg13g2_fill_2 FILLER_49_203 ();
 sg13g2_decap_8 FILLER_49_209 ();
 sg13g2_decap_4 FILLER_49_216 ();
 sg13g2_fill_1 FILLER_49_220 ();
 sg13g2_decap_8 FILLER_49_234 ();
 sg13g2_decap_4 FILLER_49_241 ();
 sg13g2_fill_1 FILLER_49_245 ();
 sg13g2_fill_2 FILLER_49_261 ();
 sg13g2_fill_1 FILLER_49_263 ();
 sg13g2_fill_2 FILLER_49_273 ();
 sg13g2_fill_1 FILLER_49_275 ();
 sg13g2_decap_8 FILLER_49_298 ();
 sg13g2_fill_1 FILLER_49_305 ();
 sg13g2_fill_1 FILLER_49_355 ();
 sg13g2_decap_8 FILLER_49_365 ();
 sg13g2_fill_2 FILLER_49_372 ();
 sg13g2_fill_1 FILLER_49_374 ();
 sg13g2_fill_2 FILLER_49_403 ();
 sg13g2_fill_2 FILLER_49_423 ();
 sg13g2_decap_8 FILLER_49_457 ();
 sg13g2_decap_8 FILLER_49_464 ();
 sg13g2_fill_1 FILLER_49_471 ();
 sg13g2_fill_2 FILLER_49_527 ();
 sg13g2_fill_1 FILLER_49_529 ();
 sg13g2_fill_2 FILLER_49_557 ();
 sg13g2_decap_4 FILLER_49_578 ();
 sg13g2_decap_8 FILLER_49_635 ();
 sg13g2_decap_8 FILLER_49_642 ();
 sg13g2_decap_8 FILLER_49_649 ();
 sg13g2_decap_8 FILLER_49_656 ();
 sg13g2_decap_8 FILLER_49_663 ();
 sg13g2_decap_8 FILLER_49_670 ();
 sg13g2_decap_8 FILLER_49_677 ();
 sg13g2_decap_8 FILLER_49_684 ();
 sg13g2_decap_8 FILLER_49_691 ();
 sg13g2_decap_8 FILLER_49_698 ();
 sg13g2_decap_8 FILLER_49_705 ();
 sg13g2_decap_8 FILLER_49_712 ();
 sg13g2_fill_1 FILLER_49_719 ();
 sg13g2_decap_8 FILLER_49_733 ();
 sg13g2_decap_8 FILLER_49_740 ();
 sg13g2_decap_8 FILLER_49_747 ();
 sg13g2_decap_8 FILLER_49_754 ();
 sg13g2_decap_8 FILLER_49_761 ();
 sg13g2_decap_8 FILLER_49_768 ();
 sg13g2_decap_8 FILLER_49_775 ();
 sg13g2_decap_8 FILLER_49_782 ();
 sg13g2_decap_8 FILLER_49_789 ();
 sg13g2_decap_8 FILLER_49_796 ();
 sg13g2_decap_8 FILLER_49_803 ();
 sg13g2_decap_8 FILLER_49_810 ();
 sg13g2_decap_8 FILLER_49_817 ();
 sg13g2_decap_8 FILLER_49_824 ();
 sg13g2_decap_8 FILLER_49_831 ();
 sg13g2_decap_8 FILLER_49_838 ();
 sg13g2_decap_8 FILLER_49_845 ();
 sg13g2_decap_8 FILLER_49_852 ();
 sg13g2_fill_2 FILLER_49_859 ();
 sg13g2_fill_1 FILLER_49_861 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_98 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_decap_8 FILLER_50_112 ();
 sg13g2_decap_4 FILLER_50_132 ();
 sg13g2_fill_2 FILLER_50_136 ();
 sg13g2_decap_8 FILLER_50_151 ();
 sg13g2_fill_1 FILLER_50_158 ();
 sg13g2_decap_8 FILLER_50_172 ();
 sg13g2_decap_4 FILLER_50_179 ();
 sg13g2_fill_1 FILLER_50_183 ();
 sg13g2_decap_4 FILLER_50_238 ();
 sg13g2_fill_1 FILLER_50_242 ();
 sg13g2_fill_2 FILLER_50_267 ();
 sg13g2_fill_1 FILLER_50_274 ();
 sg13g2_fill_1 FILLER_50_288 ();
 sg13g2_decap_4 FILLER_50_309 ();
 sg13g2_fill_1 FILLER_50_313 ();
 sg13g2_fill_2 FILLER_50_319 ();
 sg13g2_fill_1 FILLER_50_321 ();
 sg13g2_fill_1 FILLER_50_346 ();
 sg13g2_fill_1 FILLER_50_383 ();
 sg13g2_decap_4 FILLER_50_402 ();
 sg13g2_decap_4 FILLER_50_423 ();
 sg13g2_fill_1 FILLER_50_427 ();
 sg13g2_fill_2 FILLER_50_442 ();
 sg13g2_fill_2 FILLER_50_460 ();
 sg13g2_decap_8 FILLER_50_472 ();
 sg13g2_decap_8 FILLER_50_479 ();
 sg13g2_decap_4 FILLER_50_486 ();
 sg13g2_fill_1 FILLER_50_490 ();
 sg13g2_decap_4 FILLER_50_500 ();
 sg13g2_fill_1 FILLER_50_562 ();
 sg13g2_fill_2 FILLER_50_590 ();
 sg13g2_decap_4 FILLER_50_610 ();
 sg13g2_decap_8 FILLER_50_640 ();
 sg13g2_decap_8 FILLER_50_647 ();
 sg13g2_decap_8 FILLER_50_654 ();
 sg13g2_decap_4 FILLER_50_661 ();
 sg13g2_fill_2 FILLER_50_665 ();
 sg13g2_decap_8 FILLER_50_680 ();
 sg13g2_decap_8 FILLER_50_687 ();
 sg13g2_decap_8 FILLER_50_694 ();
 sg13g2_decap_8 FILLER_50_701 ();
 sg13g2_decap_8 FILLER_50_708 ();
 sg13g2_decap_8 FILLER_50_715 ();
 sg13g2_decap_8 FILLER_50_722 ();
 sg13g2_decap_8 FILLER_50_729 ();
 sg13g2_decap_8 FILLER_50_736 ();
 sg13g2_decap_8 FILLER_50_743 ();
 sg13g2_decap_8 FILLER_50_750 ();
 sg13g2_decap_8 FILLER_50_757 ();
 sg13g2_decap_8 FILLER_50_764 ();
 sg13g2_decap_8 FILLER_50_771 ();
 sg13g2_decap_8 FILLER_50_778 ();
 sg13g2_decap_8 FILLER_50_785 ();
 sg13g2_decap_8 FILLER_50_792 ();
 sg13g2_decap_8 FILLER_50_799 ();
 sg13g2_decap_8 FILLER_50_806 ();
 sg13g2_decap_8 FILLER_50_813 ();
 sg13g2_decap_8 FILLER_50_820 ();
 sg13g2_decap_8 FILLER_50_827 ();
 sg13g2_decap_8 FILLER_50_834 ();
 sg13g2_decap_8 FILLER_50_841 ();
 sg13g2_decap_8 FILLER_50_848 ();
 sg13g2_decap_8 FILLER_50_855 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_fill_2 FILLER_51_49 ();
 sg13g2_fill_1 FILLER_51_51 ();
 sg13g2_decap_8 FILLER_51_65 ();
 sg13g2_decap_8 FILLER_51_72 ();
 sg13g2_decap_8 FILLER_51_79 ();
 sg13g2_decap_4 FILLER_51_86 ();
 sg13g2_fill_2 FILLER_51_90 ();
 sg13g2_decap_8 FILLER_51_96 ();
 sg13g2_decap_8 FILLER_51_103 ();
 sg13g2_decap_8 FILLER_51_110 ();
 sg13g2_decap_8 FILLER_51_117 ();
 sg13g2_decap_8 FILLER_51_124 ();
 sg13g2_fill_1 FILLER_51_131 ();
 sg13g2_fill_1 FILLER_51_213 ();
 sg13g2_fill_2 FILLER_51_230 ();
 sg13g2_decap_8 FILLER_51_241 ();
 sg13g2_fill_2 FILLER_51_248 ();
 sg13g2_fill_1 FILLER_51_250 ();
 sg13g2_fill_2 FILLER_51_273 ();
 sg13g2_fill_1 FILLER_51_275 ();
 sg13g2_fill_1 FILLER_51_294 ();
 sg13g2_decap_8 FILLER_51_305 ();
 sg13g2_decap_4 FILLER_51_324 ();
 sg13g2_fill_1 FILLER_51_360 ();
 sg13g2_fill_1 FILLER_51_369 ();
 sg13g2_fill_2 FILLER_51_379 ();
 sg13g2_fill_2 FILLER_51_400 ();
 sg13g2_fill_2 FILLER_51_411 ();
 sg13g2_fill_1 FILLER_51_413 ();
 sg13g2_fill_2 FILLER_51_418 ();
 sg13g2_fill_2 FILLER_51_432 ();
 sg13g2_fill_2 FILLER_51_451 ();
 sg13g2_decap_4 FILLER_51_474 ();
 sg13g2_fill_1 FILLER_51_478 ();
 sg13g2_fill_2 FILLER_51_495 ();
 sg13g2_fill_1 FILLER_51_497 ();
 sg13g2_fill_1 FILLER_51_526 ();
 sg13g2_fill_2 FILLER_51_531 ();
 sg13g2_decap_8 FILLER_51_537 ();
 sg13g2_fill_1 FILLER_51_544 ();
 sg13g2_decap_4 FILLER_51_551 ();
 sg13g2_fill_2 FILLER_51_592 ();
 sg13g2_fill_1 FILLER_51_594 ();
 sg13g2_decap_8 FILLER_51_609 ();
 sg13g2_fill_1 FILLER_51_616 ();
 sg13g2_fill_1 FILLER_51_645 ();
 sg13g2_fill_2 FILLER_51_657 ();
 sg13g2_fill_1 FILLER_51_672 ();
 sg13g2_decap_8 FILLER_51_682 ();
 sg13g2_decap_8 FILLER_51_689 ();
 sg13g2_decap_8 FILLER_51_696 ();
 sg13g2_decap_8 FILLER_51_703 ();
 sg13g2_decap_8 FILLER_51_710 ();
 sg13g2_decap_8 FILLER_51_717 ();
 sg13g2_decap_8 FILLER_51_724 ();
 sg13g2_decap_8 FILLER_51_731 ();
 sg13g2_decap_8 FILLER_51_738 ();
 sg13g2_decap_8 FILLER_51_745 ();
 sg13g2_decap_8 FILLER_51_752 ();
 sg13g2_decap_8 FILLER_51_759 ();
 sg13g2_decap_8 FILLER_51_766 ();
 sg13g2_decap_8 FILLER_51_773 ();
 sg13g2_decap_8 FILLER_51_780 ();
 sg13g2_decap_8 FILLER_51_787 ();
 sg13g2_decap_8 FILLER_51_794 ();
 sg13g2_decap_8 FILLER_51_801 ();
 sg13g2_decap_8 FILLER_51_808 ();
 sg13g2_decap_8 FILLER_51_815 ();
 sg13g2_decap_8 FILLER_51_822 ();
 sg13g2_decap_8 FILLER_51_829 ();
 sg13g2_decap_8 FILLER_51_836 ();
 sg13g2_decap_8 FILLER_51_843 ();
 sg13g2_decap_8 FILLER_51_850 ();
 sg13g2_decap_4 FILLER_51_857 ();
 sg13g2_fill_1 FILLER_51_861 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_fill_1 FILLER_52_84 ();
 sg13g2_fill_1 FILLER_52_141 ();
 sg13g2_fill_1 FILLER_52_151 ();
 sg13g2_decap_8 FILLER_52_156 ();
 sg13g2_decap_4 FILLER_52_163 ();
 sg13g2_fill_2 FILLER_52_167 ();
 sg13g2_fill_2 FILLER_52_173 ();
 sg13g2_fill_2 FILLER_52_179 ();
 sg13g2_fill_1 FILLER_52_199 ();
 sg13g2_decap_4 FILLER_52_246 ();
 sg13g2_fill_2 FILLER_52_267 ();
 sg13g2_fill_1 FILLER_52_269 ();
 sg13g2_fill_2 FILLER_52_282 ();
 sg13g2_fill_1 FILLER_52_303 ();
 sg13g2_decap_8 FILLER_52_327 ();
 sg13g2_decap_4 FILLER_52_334 ();
 sg13g2_fill_2 FILLER_52_342 ();
 sg13g2_fill_1 FILLER_52_344 ();
 sg13g2_fill_1 FILLER_52_376 ();
 sg13g2_fill_1 FILLER_52_387 ();
 sg13g2_fill_2 FILLER_52_424 ();
 sg13g2_fill_1 FILLER_52_438 ();
 sg13g2_fill_2 FILLER_52_463 ();
 sg13g2_fill_1 FILLER_52_465 ();
 sg13g2_fill_2 FILLER_52_472 ();
 sg13g2_fill_1 FILLER_52_474 ();
 sg13g2_decap_8 FILLER_52_497 ();
 sg13g2_fill_2 FILLER_52_504 ();
 sg13g2_fill_1 FILLER_52_506 ();
 sg13g2_fill_2 FILLER_52_526 ();
 sg13g2_fill_1 FILLER_52_528 ();
 sg13g2_decap_4 FILLER_52_591 ();
 sg13g2_fill_1 FILLER_52_595 ();
 sg13g2_fill_1 FILLER_52_601 ();
 sg13g2_decap_4 FILLER_52_607 ();
 sg13g2_fill_2 FILLER_52_611 ();
 sg13g2_fill_1 FILLER_52_643 ();
 sg13g2_fill_1 FILLER_52_649 ();
 sg13g2_fill_2 FILLER_52_655 ();
 sg13g2_fill_1 FILLER_52_657 ();
 sg13g2_decap_8 FILLER_52_686 ();
 sg13g2_decap_8 FILLER_52_693 ();
 sg13g2_decap_8 FILLER_52_700 ();
 sg13g2_decap_8 FILLER_52_707 ();
 sg13g2_decap_8 FILLER_52_714 ();
 sg13g2_decap_8 FILLER_52_721 ();
 sg13g2_decap_8 FILLER_52_728 ();
 sg13g2_decap_8 FILLER_52_735 ();
 sg13g2_decap_8 FILLER_52_742 ();
 sg13g2_decap_8 FILLER_52_749 ();
 sg13g2_decap_8 FILLER_52_756 ();
 sg13g2_decap_8 FILLER_52_763 ();
 sg13g2_decap_8 FILLER_52_770 ();
 sg13g2_decap_8 FILLER_52_777 ();
 sg13g2_decap_8 FILLER_52_784 ();
 sg13g2_decap_8 FILLER_52_791 ();
 sg13g2_decap_8 FILLER_52_798 ();
 sg13g2_decap_8 FILLER_52_805 ();
 sg13g2_decap_8 FILLER_52_812 ();
 sg13g2_decap_8 FILLER_52_819 ();
 sg13g2_decap_8 FILLER_52_826 ();
 sg13g2_decap_8 FILLER_52_833 ();
 sg13g2_decap_8 FILLER_52_840 ();
 sg13g2_decap_8 FILLER_52_847 ();
 sg13g2_decap_8 FILLER_52_854 ();
 sg13g2_fill_1 FILLER_52_861 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_4 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_64 ();
 sg13g2_decap_8 FILLER_53_71 ();
 sg13g2_decap_8 FILLER_53_110 ();
 sg13g2_fill_1 FILLER_53_117 ();
 sg13g2_fill_2 FILLER_53_127 ();
 sg13g2_fill_2 FILLER_53_175 ();
 sg13g2_fill_1 FILLER_53_225 ();
 sg13g2_decap_8 FILLER_53_239 ();
 sg13g2_decap_4 FILLER_53_246 ();
 sg13g2_decap_8 FILLER_53_255 ();
 sg13g2_decap_4 FILLER_53_262 ();
 sg13g2_decap_4 FILLER_53_270 ();
 sg13g2_fill_1 FILLER_53_274 ();
 sg13g2_decap_4 FILLER_53_326 ();
 sg13g2_fill_2 FILLER_53_330 ();
 sg13g2_decap_8 FILLER_53_340 ();
 sg13g2_decap_8 FILLER_53_347 ();
 sg13g2_decap_8 FILLER_53_354 ();
 sg13g2_fill_1 FILLER_53_361 ();
 sg13g2_fill_1 FILLER_53_391 ();
 sg13g2_fill_1 FILLER_53_405 ();
 sg13g2_decap_4 FILLER_53_415 ();
 sg13g2_fill_1 FILLER_53_419 ();
 sg13g2_decap_8 FILLER_53_434 ();
 sg13g2_decap_8 FILLER_53_441 ();
 sg13g2_decap_4 FILLER_53_468 ();
 sg13g2_decap_8 FILLER_53_491 ();
 sg13g2_decap_8 FILLER_53_498 ();
 sg13g2_decap_4 FILLER_53_505 ();
 sg13g2_fill_1 FILLER_53_509 ();
 sg13g2_decap_4 FILLER_53_524 ();
 sg13g2_fill_2 FILLER_53_528 ();
 sg13g2_decap_8 FILLER_53_534 ();
 sg13g2_fill_2 FILLER_53_541 ();
 sg13g2_decap_8 FILLER_53_549 ();
 sg13g2_fill_2 FILLER_53_575 ();
 sg13g2_fill_1 FILLER_53_577 ();
 sg13g2_fill_2 FILLER_53_583 ();
 sg13g2_decap_8 FILLER_53_588 ();
 sg13g2_fill_2 FILLER_53_617 ();
 sg13g2_fill_1 FILLER_53_619 ();
 sg13g2_fill_2 FILLER_53_631 ();
 sg13g2_fill_1 FILLER_53_633 ();
 sg13g2_fill_1 FILLER_53_638 ();
 sg13g2_fill_2 FILLER_53_657 ();
 sg13g2_decap_4 FILLER_53_667 ();
 sg13g2_decap_8 FILLER_53_688 ();
 sg13g2_decap_8 FILLER_53_695 ();
 sg13g2_decap_8 FILLER_53_702 ();
 sg13g2_decap_8 FILLER_53_709 ();
 sg13g2_decap_8 FILLER_53_716 ();
 sg13g2_decap_8 FILLER_53_723 ();
 sg13g2_decap_8 FILLER_53_730 ();
 sg13g2_decap_8 FILLER_53_737 ();
 sg13g2_decap_8 FILLER_53_744 ();
 sg13g2_decap_8 FILLER_53_751 ();
 sg13g2_decap_8 FILLER_53_758 ();
 sg13g2_decap_8 FILLER_53_765 ();
 sg13g2_decap_8 FILLER_53_772 ();
 sg13g2_decap_8 FILLER_53_779 ();
 sg13g2_decap_8 FILLER_53_786 ();
 sg13g2_decap_8 FILLER_53_793 ();
 sg13g2_decap_8 FILLER_53_800 ();
 sg13g2_decap_8 FILLER_53_807 ();
 sg13g2_decap_8 FILLER_53_814 ();
 sg13g2_decap_8 FILLER_53_821 ();
 sg13g2_decap_8 FILLER_53_828 ();
 sg13g2_decap_8 FILLER_53_835 ();
 sg13g2_decap_8 FILLER_53_842 ();
 sg13g2_decap_8 FILLER_53_849 ();
 sg13g2_decap_4 FILLER_53_856 ();
 sg13g2_fill_2 FILLER_53_860 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_fill_1 FILLER_54_28 ();
 sg13g2_fill_2 FILLER_54_33 ();
 sg13g2_fill_1 FILLER_54_35 ();
 sg13g2_fill_1 FILLER_54_50 ();
 sg13g2_fill_1 FILLER_54_111 ();
 sg13g2_decap_8 FILLER_54_142 ();
 sg13g2_decap_4 FILLER_54_149 ();
 sg13g2_fill_2 FILLER_54_158 ();
 sg13g2_fill_2 FILLER_54_163 ();
 sg13g2_fill_1 FILLER_54_165 ();
 sg13g2_fill_2 FILLER_54_174 ();
 sg13g2_fill_2 FILLER_54_189 ();
 sg13g2_fill_2 FILLER_54_195 ();
 sg13g2_fill_1 FILLER_54_197 ();
 sg13g2_fill_2 FILLER_54_207 ();
 sg13g2_fill_2 FILLER_54_220 ();
 sg13g2_fill_1 FILLER_54_222 ();
 sg13g2_decap_8 FILLER_54_239 ();
 sg13g2_decap_8 FILLER_54_246 ();
 sg13g2_fill_1 FILLER_54_253 ();
 sg13g2_fill_1 FILLER_54_259 ();
 sg13g2_decap_8 FILLER_54_276 ();
 sg13g2_decap_8 FILLER_54_283 ();
 sg13g2_fill_2 FILLER_54_290 ();
 sg13g2_fill_1 FILLER_54_292 ();
 sg13g2_decap_4 FILLER_54_297 ();
 sg13g2_decap_4 FILLER_54_306 ();
 sg13g2_fill_2 FILLER_54_315 ();
 sg13g2_fill_1 FILLER_54_317 ();
 sg13g2_decap_8 FILLER_54_348 ();
 sg13g2_fill_2 FILLER_54_355 ();
 sg13g2_fill_1 FILLER_54_357 ();
 sg13g2_fill_2 FILLER_54_376 ();
 sg13g2_fill_1 FILLER_54_378 ();
 sg13g2_decap_4 FILLER_54_407 ();
 sg13g2_fill_2 FILLER_54_443 ();
 sg13g2_fill_1 FILLER_54_445 ();
 sg13g2_fill_2 FILLER_54_452 ();
 sg13g2_fill_1 FILLER_54_464 ();
 sg13g2_fill_2 FILLER_54_470 ();
 sg13g2_decap_4 FILLER_54_478 ();
 sg13g2_decap_4 FILLER_54_487 ();
 sg13g2_fill_2 FILLER_54_491 ();
 sg13g2_fill_1 FILLER_54_505 ();
 sg13g2_decap_4 FILLER_54_531 ();
 sg13g2_fill_2 FILLER_54_569 ();
 sg13g2_fill_1 FILLER_54_571 ();
 sg13g2_fill_1 FILLER_54_585 ();
 sg13g2_decap_4 FILLER_54_600 ();
 sg13g2_fill_1 FILLER_54_604 ();
 sg13g2_decap_8 FILLER_54_610 ();
 sg13g2_fill_2 FILLER_54_617 ();
 sg13g2_decap_4 FILLER_54_624 ();
 sg13g2_fill_1 FILLER_54_628 ();
 sg13g2_decap_8 FILLER_54_635 ();
 sg13g2_fill_2 FILLER_54_642 ();
 sg13g2_fill_1 FILLER_54_644 ();
 sg13g2_fill_1 FILLER_54_654 ();
 sg13g2_decap_8 FILLER_54_671 ();
 sg13g2_fill_2 FILLER_54_684 ();
 sg13g2_decap_8 FILLER_54_693 ();
 sg13g2_decap_8 FILLER_54_700 ();
 sg13g2_decap_8 FILLER_54_707 ();
 sg13g2_decap_8 FILLER_54_714 ();
 sg13g2_decap_8 FILLER_54_721 ();
 sg13g2_decap_8 FILLER_54_728 ();
 sg13g2_decap_8 FILLER_54_735 ();
 sg13g2_decap_8 FILLER_54_742 ();
 sg13g2_decap_8 FILLER_54_749 ();
 sg13g2_decap_8 FILLER_54_756 ();
 sg13g2_decap_8 FILLER_54_763 ();
 sg13g2_decap_8 FILLER_54_770 ();
 sg13g2_decap_8 FILLER_54_777 ();
 sg13g2_decap_8 FILLER_54_784 ();
 sg13g2_decap_8 FILLER_54_791 ();
 sg13g2_decap_8 FILLER_54_798 ();
 sg13g2_decap_8 FILLER_54_805 ();
 sg13g2_decap_8 FILLER_54_812 ();
 sg13g2_decap_8 FILLER_54_819 ();
 sg13g2_decap_8 FILLER_54_826 ();
 sg13g2_decap_8 FILLER_54_833 ();
 sg13g2_decap_8 FILLER_54_840 ();
 sg13g2_decap_8 FILLER_54_847 ();
 sg13g2_decap_8 FILLER_54_854 ();
 sg13g2_fill_1 FILLER_54_861 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_7 ();
 sg13g2_fill_1 FILLER_55_9 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_fill_2 FILLER_55_21 ();
 sg13g2_fill_1 FILLER_55_23 ();
 sg13g2_decap_8 FILLER_55_65 ();
 sg13g2_decap_4 FILLER_55_72 ();
 sg13g2_fill_1 FILLER_55_76 ();
 sg13g2_fill_2 FILLER_55_103 ();
 sg13g2_fill_1 FILLER_55_105 ();
 sg13g2_fill_2 FILLER_55_154 ();
 sg13g2_fill_1 FILLER_55_173 ();
 sg13g2_decap_4 FILLER_55_193 ();
 sg13g2_decap_8 FILLER_55_219 ();
 sg13g2_decap_4 FILLER_55_226 ();
 sg13g2_decap_4 FILLER_55_242 ();
 sg13g2_decap_8 FILLER_55_273 ();
 sg13g2_decap_8 FILLER_55_280 ();
 sg13g2_decap_8 FILLER_55_287 ();
 sg13g2_fill_2 FILLER_55_294 ();
 sg13g2_fill_1 FILLER_55_296 ();
 sg13g2_decap_4 FILLER_55_304 ();
 sg13g2_decap_8 FILLER_55_314 ();
 sg13g2_fill_2 FILLER_55_321 ();
 sg13g2_decap_8 FILLER_55_339 ();
 sg13g2_fill_1 FILLER_55_346 ();
 sg13g2_decap_4 FILLER_55_384 ();
 sg13g2_decap_8 FILLER_55_400 ();
 sg13g2_fill_1 FILLER_55_407 ();
 sg13g2_fill_1 FILLER_55_421 ();
 sg13g2_decap_8 FILLER_55_436 ();
 sg13g2_decap_8 FILLER_55_443 ();
 sg13g2_fill_1 FILLER_55_450 ();
 sg13g2_fill_1 FILLER_55_457 ();
 sg13g2_fill_2 FILLER_55_461 ();
 sg13g2_fill_1 FILLER_55_463 ();
 sg13g2_fill_2 FILLER_55_482 ();
 sg13g2_fill_2 FILLER_55_500 ();
 sg13g2_fill_1 FILLER_55_502 ();
 sg13g2_decap_8 FILLER_55_519 ();
 sg13g2_decap_8 FILLER_55_526 ();
 sg13g2_fill_1 FILLER_55_533 ();
 sg13g2_decap_8 FILLER_55_546 ();
 sg13g2_fill_2 FILLER_55_553 ();
 sg13g2_fill_2 FILLER_55_578 ();
 sg13g2_fill_1 FILLER_55_580 ();
 sg13g2_decap_8 FILLER_55_599 ();
 sg13g2_fill_2 FILLER_55_606 ();
 sg13g2_fill_1 FILLER_55_608 ();
 sg13g2_fill_2 FILLER_55_614 ();
 sg13g2_fill_1 FILLER_55_620 ();
 sg13g2_decap_8 FILLER_55_634 ();
 sg13g2_fill_2 FILLER_55_654 ();
 sg13g2_fill_2 FILLER_55_669 ();
 sg13g2_fill_1 FILLER_55_671 ();
 sg13g2_decap_4 FILLER_55_682 ();
 sg13g2_decap_8 FILLER_55_699 ();
 sg13g2_decap_8 FILLER_55_706 ();
 sg13g2_decap_8 FILLER_55_713 ();
 sg13g2_decap_8 FILLER_55_720 ();
 sg13g2_decap_8 FILLER_55_727 ();
 sg13g2_decap_8 FILLER_55_734 ();
 sg13g2_decap_8 FILLER_55_741 ();
 sg13g2_decap_8 FILLER_55_748 ();
 sg13g2_decap_8 FILLER_55_755 ();
 sg13g2_decap_8 FILLER_55_762 ();
 sg13g2_decap_8 FILLER_55_769 ();
 sg13g2_decap_8 FILLER_55_776 ();
 sg13g2_decap_8 FILLER_55_783 ();
 sg13g2_decap_8 FILLER_55_790 ();
 sg13g2_decap_8 FILLER_55_797 ();
 sg13g2_decap_8 FILLER_55_804 ();
 sg13g2_decap_8 FILLER_55_811 ();
 sg13g2_decap_8 FILLER_55_818 ();
 sg13g2_decap_8 FILLER_55_825 ();
 sg13g2_decap_8 FILLER_55_832 ();
 sg13g2_decap_8 FILLER_55_839 ();
 sg13g2_decap_8 FILLER_55_846 ();
 sg13g2_decap_8 FILLER_55_853 ();
 sg13g2_fill_2 FILLER_55_860 ();
 sg13g2_decap_4 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_50 ();
 sg13g2_fill_1 FILLER_56_57 ();
 sg13g2_fill_1 FILLER_56_98 ();
 sg13g2_fill_2 FILLER_56_113 ();
 sg13g2_fill_1 FILLER_56_115 ();
 sg13g2_fill_2 FILLER_56_125 ();
 sg13g2_decap_8 FILLER_56_132 ();
 sg13g2_fill_1 FILLER_56_139 ();
 sg13g2_decap_8 FILLER_56_144 ();
 sg13g2_fill_2 FILLER_56_164 ();
 sg13g2_fill_1 FILLER_56_166 ();
 sg13g2_fill_2 FILLER_56_173 ();
 sg13g2_decap_8 FILLER_56_217 ();
 sg13g2_decap_8 FILLER_56_224 ();
 sg13g2_fill_1 FILLER_56_231 ();
 sg13g2_decap_8 FILLER_56_237 ();
 sg13g2_decap_4 FILLER_56_244 ();
 sg13g2_fill_1 FILLER_56_258 ();
 sg13g2_decap_8 FILLER_56_268 ();
 sg13g2_fill_2 FILLER_56_275 ();
 sg13g2_fill_1 FILLER_56_277 ();
 sg13g2_fill_1 FILLER_56_285 ();
 sg13g2_decap_8 FILLER_56_291 ();
 sg13g2_decap_4 FILLER_56_298 ();
 sg13g2_decap_8 FILLER_56_306 ();
 sg13g2_decap_8 FILLER_56_313 ();
 sg13g2_fill_1 FILLER_56_320 ();
 sg13g2_fill_2 FILLER_56_332 ();
 sg13g2_fill_1 FILLER_56_344 ();
 sg13g2_fill_2 FILLER_56_362 ();
 sg13g2_fill_2 FILLER_56_372 ();
 sg13g2_fill_2 FILLER_56_390 ();
 sg13g2_fill_1 FILLER_56_392 ();
 sg13g2_decap_4 FILLER_56_406 ();
 sg13g2_fill_1 FILLER_56_410 ();
 sg13g2_decap_8 FILLER_56_424 ();
 sg13g2_decap_8 FILLER_56_431 ();
 sg13g2_fill_2 FILLER_56_438 ();
 sg13g2_decap_8 FILLER_56_461 ();
 sg13g2_decap_4 FILLER_56_468 ();
 sg13g2_fill_2 FILLER_56_477 ();
 sg13g2_fill_1 FILLER_56_479 ();
 sg13g2_decap_4 FILLER_56_494 ();
 sg13g2_fill_1 FILLER_56_498 ();
 sg13g2_fill_2 FILLER_56_504 ();
 sg13g2_fill_1 FILLER_56_506 ();
 sg13g2_fill_1 FILLER_56_519 ();
 sg13g2_fill_2 FILLER_56_528 ();
 sg13g2_fill_2 FILLER_56_544 ();
 sg13g2_fill_2 FILLER_56_554 ();
 sg13g2_fill_2 FILLER_56_561 ();
 sg13g2_fill_1 FILLER_56_563 ();
 sg13g2_decap_4 FILLER_56_608 ();
 sg13g2_decap_8 FILLER_56_634 ();
 sg13g2_decap_4 FILLER_56_641 ();
 sg13g2_decap_8 FILLER_56_650 ();
 sg13g2_decap_8 FILLER_56_707 ();
 sg13g2_decap_8 FILLER_56_714 ();
 sg13g2_decap_8 FILLER_56_721 ();
 sg13g2_decap_8 FILLER_56_728 ();
 sg13g2_decap_8 FILLER_56_735 ();
 sg13g2_decap_8 FILLER_56_742 ();
 sg13g2_decap_8 FILLER_56_749 ();
 sg13g2_decap_8 FILLER_56_756 ();
 sg13g2_decap_8 FILLER_56_763 ();
 sg13g2_decap_8 FILLER_56_770 ();
 sg13g2_decap_8 FILLER_56_777 ();
 sg13g2_decap_8 FILLER_56_784 ();
 sg13g2_decap_8 FILLER_56_791 ();
 sg13g2_decap_8 FILLER_56_798 ();
 sg13g2_decap_8 FILLER_56_805 ();
 sg13g2_decap_8 FILLER_56_812 ();
 sg13g2_decap_8 FILLER_56_819 ();
 sg13g2_decap_8 FILLER_56_826 ();
 sg13g2_decap_8 FILLER_56_833 ();
 sg13g2_decap_8 FILLER_56_840 ();
 sg13g2_decap_8 FILLER_56_847 ();
 sg13g2_decap_8 FILLER_56_854 ();
 sg13g2_fill_1 FILLER_56_861 ();
 sg13g2_decap_4 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_32 ();
 sg13g2_fill_1 FILLER_57_34 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_fill_1 FILLER_57_63 ();
 sg13g2_decap_4 FILLER_57_68 ();
 sg13g2_fill_2 FILLER_57_72 ();
 sg13g2_decap_8 FILLER_57_160 ();
 sg13g2_decap_4 FILLER_57_167 ();
 sg13g2_decap_8 FILLER_57_191 ();
 sg13g2_decap_4 FILLER_57_198 ();
 sg13g2_fill_2 FILLER_57_214 ();
 sg13g2_fill_2 FILLER_57_240 ();
 sg13g2_fill_1 FILLER_57_242 ();
 sg13g2_fill_1 FILLER_57_253 ();
 sg13g2_fill_2 FILLER_57_273 ();
 sg13g2_fill_1 FILLER_57_275 ();
 sg13g2_fill_2 FILLER_57_351 ();
 sg13g2_fill_1 FILLER_57_353 ();
 sg13g2_decap_8 FILLER_57_360 ();
 sg13g2_decap_8 FILLER_57_372 ();
 sg13g2_decap_4 FILLER_57_379 ();
 sg13g2_fill_2 FILLER_57_383 ();
 sg13g2_fill_2 FILLER_57_390 ();
 sg13g2_decap_8 FILLER_57_401 ();
 sg13g2_decap_8 FILLER_57_408 ();
 sg13g2_fill_1 FILLER_57_415 ();
 sg13g2_fill_2 FILLER_57_465 ();
 sg13g2_decap_8 FILLER_57_471 ();
 sg13g2_decap_4 FILLER_57_478 ();
 sg13g2_fill_2 FILLER_57_482 ();
 sg13g2_decap_8 FILLER_57_497 ();
 sg13g2_fill_1 FILLER_57_504 ();
 sg13g2_fill_1 FILLER_57_526 ();
 sg13g2_fill_1 FILLER_57_545 ();
 sg13g2_decap_4 FILLER_57_553 ();
 sg13g2_fill_1 FILLER_57_574 ();
 sg13g2_decap_8 FILLER_57_593 ();
 sg13g2_decap_8 FILLER_57_600 ();
 sg13g2_fill_2 FILLER_57_607 ();
 sg13g2_fill_1 FILLER_57_609 ();
 sg13g2_decap_8 FILLER_57_634 ();
 sg13g2_decap_8 FILLER_57_685 ();
 sg13g2_decap_8 FILLER_57_692 ();
 sg13g2_decap_8 FILLER_57_699 ();
 sg13g2_decap_8 FILLER_57_706 ();
 sg13g2_decap_8 FILLER_57_713 ();
 sg13g2_decap_8 FILLER_57_720 ();
 sg13g2_decap_8 FILLER_57_727 ();
 sg13g2_fill_2 FILLER_57_734 ();
 sg13g2_fill_1 FILLER_57_736 ();
 sg13g2_decap_8 FILLER_57_741 ();
 sg13g2_fill_2 FILLER_57_748 ();
 sg13g2_decap_4 FILLER_57_755 ();
 sg13g2_fill_2 FILLER_57_759 ();
 sg13g2_decap_8 FILLER_57_779 ();
 sg13g2_decap_8 FILLER_57_786 ();
 sg13g2_decap_8 FILLER_57_796 ();
 sg13g2_decap_8 FILLER_57_803 ();
 sg13g2_decap_8 FILLER_57_810 ();
 sg13g2_decap_8 FILLER_57_817 ();
 sg13g2_decap_8 FILLER_57_824 ();
 sg13g2_decap_8 FILLER_57_831 ();
 sg13g2_decap_8 FILLER_57_838 ();
 sg13g2_decap_8 FILLER_57_845 ();
 sg13g2_decap_8 FILLER_57_852 ();
 sg13g2_fill_2 FILLER_57_859 ();
 sg13g2_fill_1 FILLER_57_861 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_7 ();
 sg13g2_fill_2 FILLER_58_13 ();
 sg13g2_fill_2 FILLER_58_47 ();
 sg13g2_fill_1 FILLER_58_49 ();
 sg13g2_fill_1 FILLER_58_56 ();
 sg13g2_fill_1 FILLER_58_112 ();
 sg13g2_decap_4 FILLER_58_128 ();
 sg13g2_fill_1 FILLER_58_136 ();
 sg13g2_decap_8 FILLER_58_141 ();
 sg13g2_decap_8 FILLER_58_148 ();
 sg13g2_decap_8 FILLER_58_155 ();
 sg13g2_fill_2 FILLER_58_162 ();
 sg13g2_fill_1 FILLER_58_164 ();
 sg13g2_fill_1 FILLER_58_175 ();
 sg13g2_fill_1 FILLER_58_200 ();
 sg13g2_fill_2 FILLER_58_219 ();
 sg13g2_fill_2 FILLER_58_230 ();
 sg13g2_fill_1 FILLER_58_232 ();
 sg13g2_fill_2 FILLER_58_238 ();
 sg13g2_fill_1 FILLER_58_240 ();
 sg13g2_fill_1 FILLER_58_247 ();
 sg13g2_fill_1 FILLER_58_257 ();
 sg13g2_decap_4 FILLER_58_298 ();
 sg13g2_decap_8 FILLER_58_315 ();
 sg13g2_fill_2 FILLER_58_322 ();
 sg13g2_fill_1 FILLER_58_324 ();
 sg13g2_decap_8 FILLER_58_334 ();
 sg13g2_fill_1 FILLER_58_341 ();
 sg13g2_decap_4 FILLER_58_365 ();
 sg13g2_fill_1 FILLER_58_369 ();
 sg13g2_fill_2 FILLER_58_392 ();
 sg13g2_decap_4 FILLER_58_399 ();
 sg13g2_fill_2 FILLER_58_403 ();
 sg13g2_fill_2 FILLER_58_418 ();
 sg13g2_fill_1 FILLER_58_420 ();
 sg13g2_decap_4 FILLER_58_425 ();
 sg13g2_fill_2 FILLER_58_429 ();
 sg13g2_fill_2 FILLER_58_490 ();
 sg13g2_fill_1 FILLER_58_492 ();
 sg13g2_fill_2 FILLER_58_506 ();
 sg13g2_fill_1 FILLER_58_508 ();
 sg13g2_decap_8 FILLER_58_513 ();
 sg13g2_decap_8 FILLER_58_520 ();
 sg13g2_decap_8 FILLER_58_527 ();
 sg13g2_decap_8 FILLER_58_534 ();
 sg13g2_fill_2 FILLER_58_541 ();
 sg13g2_fill_2 FILLER_58_551 ();
 sg13g2_fill_1 FILLER_58_558 ();
 sg13g2_fill_1 FILLER_58_565 ();
 sg13g2_decap_4 FILLER_58_638 ();
 sg13g2_decap_4 FILLER_58_656 ();
 sg13g2_decap_8 FILLER_58_701 ();
 sg13g2_decap_8 FILLER_58_712 ();
 sg13g2_decap_4 FILLER_58_719 ();
 sg13g2_decap_4 FILLER_58_728 ();
 sg13g2_fill_2 FILLER_58_764 ();
 sg13g2_decap_8 FILLER_58_802 ();
 sg13g2_decap_8 FILLER_58_809 ();
 sg13g2_decap_8 FILLER_58_816 ();
 sg13g2_decap_8 FILLER_58_823 ();
 sg13g2_decap_8 FILLER_58_830 ();
 sg13g2_decap_8 FILLER_58_837 ();
 sg13g2_decap_8 FILLER_58_844 ();
 sg13g2_decap_8 FILLER_58_851 ();
 sg13g2_decap_4 FILLER_58_858 ();
 sg13g2_fill_1 FILLER_59_0 ();
 sg13g2_fill_2 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_55 ();
 sg13g2_fill_1 FILLER_59_62 ();
 sg13g2_decap_8 FILLER_59_83 ();
 sg13g2_fill_1 FILLER_59_90 ();
 sg13g2_fill_2 FILLER_59_132 ();
 sg13g2_fill_1 FILLER_59_134 ();
 sg13g2_decap_4 FILLER_59_148 ();
 sg13g2_fill_1 FILLER_59_177 ();
 sg13g2_decap_8 FILLER_59_193 ();
 sg13g2_decap_8 FILLER_59_200 ();
 sg13g2_fill_1 FILLER_59_207 ();
 sg13g2_fill_2 FILLER_59_217 ();
 sg13g2_decap_4 FILLER_59_224 ();
 sg13g2_fill_2 FILLER_59_244 ();
 sg13g2_fill_1 FILLER_59_250 ();
 sg13g2_decap_8 FILLER_59_255 ();
 sg13g2_fill_2 FILLER_59_262 ();
 sg13g2_decap_4 FILLER_59_268 ();
 sg13g2_fill_2 FILLER_59_272 ();
 sg13g2_decap_4 FILLER_59_287 ();
 sg13g2_fill_2 FILLER_59_291 ();
 sg13g2_fill_2 FILLER_59_303 ();
 sg13g2_fill_1 FILLER_59_305 ();
 sg13g2_fill_2 FILLER_59_347 ();
 sg13g2_fill_1 FILLER_59_349 ();
 sg13g2_fill_2 FILLER_59_370 ();
 sg13g2_decap_8 FILLER_59_391 ();
 sg13g2_decap_8 FILLER_59_398 ();
 sg13g2_decap_8 FILLER_59_465 ();
 sg13g2_fill_2 FILLER_59_472 ();
 sg13g2_decap_8 FILLER_59_487 ();
 sg13g2_decap_4 FILLER_59_494 ();
 sg13g2_fill_1 FILLER_59_498 ();
 sg13g2_fill_2 FILLER_59_579 ();
 sg13g2_fill_1 FILLER_59_581 ();
 sg13g2_fill_1 FILLER_59_587 ();
 sg13g2_decap_8 FILLER_59_591 ();
 sg13g2_decap_8 FILLER_59_598 ();
 sg13g2_decap_4 FILLER_59_605 ();
 sg13g2_fill_1 FILLER_59_609 ();
 sg13g2_fill_1 FILLER_59_647 ();
 sg13g2_fill_2 FILLER_59_652 ();
 sg13g2_fill_1 FILLER_59_654 ();
 sg13g2_fill_2 FILLER_59_701 ();
 sg13g2_fill_2 FILLER_59_730 ();
 sg13g2_fill_1 FILLER_59_732 ();
 sg13g2_fill_2 FILLER_59_746 ();
 sg13g2_decap_8 FILLER_59_796 ();
 sg13g2_decap_8 FILLER_59_803 ();
 sg13g2_decap_8 FILLER_59_810 ();
 sg13g2_decap_8 FILLER_59_817 ();
 sg13g2_decap_8 FILLER_59_824 ();
 sg13g2_decap_8 FILLER_59_831 ();
 sg13g2_decap_8 FILLER_59_838 ();
 sg13g2_decap_8 FILLER_59_845 ();
 sg13g2_decap_8 FILLER_59_852 ();
 sg13g2_fill_2 FILLER_59_859 ();
 sg13g2_fill_1 FILLER_59_861 ();
 sg13g2_decap_4 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_4 ();
 sg13g2_decap_8 FILLER_60_10 ();
 sg13g2_fill_2 FILLER_60_54 ();
 sg13g2_fill_1 FILLER_60_56 ();
 sg13g2_decap_4 FILLER_60_78 ();
 sg13g2_fill_2 FILLER_60_101 ();
 sg13g2_fill_1 FILLER_60_103 ();
 sg13g2_fill_1 FILLER_60_113 ();
 sg13g2_fill_1 FILLER_60_119 ();
 sg13g2_decap_8 FILLER_60_124 ();
 sg13g2_fill_1 FILLER_60_131 ();
 sg13g2_fill_2 FILLER_60_153 ();
 sg13g2_fill_1 FILLER_60_164 ();
 sg13g2_decap_8 FILLER_60_170 ();
 sg13g2_fill_2 FILLER_60_177 ();
 sg13g2_fill_2 FILLER_60_189 ();
 sg13g2_decap_8 FILLER_60_196 ();
 sg13g2_decap_8 FILLER_60_203 ();
 sg13g2_decap_4 FILLER_60_210 ();
 sg13g2_fill_1 FILLER_60_214 ();
 sg13g2_fill_2 FILLER_60_305 ();
 sg13g2_decap_4 FILLER_60_315 ();
 sg13g2_fill_2 FILLER_60_319 ();
 sg13g2_fill_1 FILLER_60_339 ();
 sg13g2_fill_2 FILLER_60_353 ();
 sg13g2_fill_1 FILLER_60_355 ();
 sg13g2_decap_8 FILLER_60_364 ();
 sg13g2_decap_8 FILLER_60_371 ();
 sg13g2_decap_8 FILLER_60_394 ();
 sg13g2_decap_4 FILLER_60_401 ();
 sg13g2_fill_1 FILLER_60_405 ();
 sg13g2_fill_2 FILLER_60_419 ();
 sg13g2_fill_1 FILLER_60_425 ();
 sg13g2_fill_1 FILLER_60_435 ();
 sg13g2_fill_1 FILLER_60_446 ();
 sg13g2_fill_1 FILLER_60_452 ();
 sg13g2_fill_2 FILLER_60_459 ();
 sg13g2_fill_1 FILLER_60_461 ();
 sg13g2_decap_4 FILLER_60_503 ();
 sg13g2_fill_1 FILLER_60_507 ();
 sg13g2_decap_8 FILLER_60_516 ();
 sg13g2_decap_4 FILLER_60_523 ();
 sg13g2_fill_2 FILLER_60_527 ();
 sg13g2_decap_4 FILLER_60_551 ();
 sg13g2_fill_1 FILLER_60_573 ();
 sg13g2_fill_1 FILLER_60_582 ();
 sg13g2_fill_1 FILLER_60_624 ();
 sg13g2_decap_8 FILLER_60_633 ();
 sg13g2_fill_2 FILLER_60_640 ();
 sg13g2_fill_1 FILLER_60_642 ();
 sg13g2_fill_2 FILLER_60_696 ();
 sg13g2_decap_8 FILLER_60_707 ();
 sg13g2_decap_8 FILLER_60_714 ();
 sg13g2_fill_1 FILLER_60_721 ();
 sg13g2_fill_1 FILLER_60_725 ();
 sg13g2_fill_2 FILLER_60_731 ();
 sg13g2_fill_1 FILLER_60_747 ();
 sg13g2_decap_4 FILLER_60_761 ();
 sg13g2_fill_2 FILLER_60_773 ();
 sg13g2_decap_8 FILLER_60_802 ();
 sg13g2_decap_8 FILLER_60_809 ();
 sg13g2_decap_8 FILLER_60_816 ();
 sg13g2_decap_8 FILLER_60_823 ();
 sg13g2_decap_8 FILLER_60_830 ();
 sg13g2_decap_8 FILLER_60_837 ();
 sg13g2_decap_8 FILLER_60_844 ();
 sg13g2_decap_8 FILLER_60_851 ();
 sg13g2_decap_4 FILLER_60_858 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_29 ();
 sg13g2_fill_1 FILLER_61_31 ();
 sg13g2_fill_1 FILLER_61_41 ();
 sg13g2_fill_1 FILLER_61_86 ();
 sg13g2_fill_2 FILLER_61_100 ();
 sg13g2_decap_8 FILLER_61_129 ();
 sg13g2_decap_8 FILLER_61_136 ();
 sg13g2_decap_4 FILLER_61_171 ();
 sg13g2_decap_4 FILLER_61_179 ();
 sg13g2_fill_1 FILLER_61_183 ();
 sg13g2_fill_2 FILLER_61_200 ();
 sg13g2_fill_1 FILLER_61_202 ();
 sg13g2_decap_4 FILLER_61_214 ();
 sg13g2_fill_2 FILLER_61_223 ();
 sg13g2_fill_1 FILLER_61_234 ();
 sg13g2_decap_8 FILLER_61_268 ();
 sg13g2_fill_1 FILLER_61_275 ();
 sg13g2_fill_1 FILLER_61_333 ();
 sg13g2_decap_4 FILLER_61_368 ();
 sg13g2_fill_2 FILLER_61_372 ();
 sg13g2_fill_1 FILLER_61_379 ();
 sg13g2_decap_8 FILLER_61_408 ();
 sg13g2_fill_1 FILLER_61_415 ();
 sg13g2_fill_2 FILLER_61_467 ();
 sg13g2_decap_8 FILLER_61_493 ();
 sg13g2_decap_4 FILLER_61_500 ();
 sg13g2_fill_1 FILLER_61_509 ();
 sg13g2_fill_1 FILLER_61_523 ();
 sg13g2_decap_8 FILLER_61_537 ();
 sg13g2_fill_2 FILLER_61_544 ();
 sg13g2_fill_1 FILLER_61_546 ();
 sg13g2_fill_1 FILLER_61_557 ();
 sg13g2_decap_8 FILLER_61_566 ();
 sg13g2_decap_8 FILLER_61_573 ();
 sg13g2_fill_1 FILLER_61_580 ();
 sg13g2_fill_1 FILLER_61_589 ();
 sg13g2_fill_2 FILLER_61_598 ();
 sg13g2_decap_8 FILLER_61_617 ();
 sg13g2_decap_8 FILLER_61_624 ();
 sg13g2_fill_2 FILLER_61_631 ();
 sg13g2_fill_1 FILLER_61_633 ();
 sg13g2_fill_2 FILLER_61_779 ();
 sg13g2_decap_8 FILLER_61_809 ();
 sg13g2_decap_8 FILLER_61_816 ();
 sg13g2_decap_8 FILLER_61_823 ();
 sg13g2_decap_8 FILLER_61_830 ();
 sg13g2_decap_8 FILLER_61_837 ();
 sg13g2_decap_8 FILLER_61_844 ();
 sg13g2_decap_8 FILLER_61_851 ();
 sg13g2_decap_4 FILLER_61_858 ();
 sg13g2_decap_4 FILLER_62_0 ();
 sg13g2_fill_2 FILLER_62_4 ();
 sg13g2_decap_8 FILLER_62_61 ();
 sg13g2_decap_4 FILLER_62_68 ();
 sg13g2_decap_4 FILLER_62_75 ();
 sg13g2_fill_2 FILLER_62_79 ();
 sg13g2_fill_1 FILLER_62_118 ();
 sg13g2_decap_8 FILLER_62_129 ();
 sg13g2_fill_1 FILLER_62_136 ();
 sg13g2_decap_8 FILLER_62_143 ();
 sg13g2_decap_4 FILLER_62_150 ();
 sg13g2_decap_8 FILLER_62_168 ();
 sg13g2_decap_4 FILLER_62_175 ();
 sg13g2_fill_1 FILLER_62_213 ();
 sg13g2_fill_2 FILLER_62_227 ();
 sg13g2_fill_2 FILLER_62_257 ();
 sg13g2_decap_8 FILLER_62_272 ();
 sg13g2_decap_4 FILLER_62_279 ();
 sg13g2_decap_8 FILLER_62_304 ();
 sg13g2_fill_1 FILLER_62_311 ();
 sg13g2_fill_2 FILLER_62_365 ();
 sg13g2_fill_1 FILLER_62_367 ();
 sg13g2_fill_1 FILLER_62_390 ();
 sg13g2_decap_8 FILLER_62_413 ();
 sg13g2_decap_8 FILLER_62_424 ();
 sg13g2_fill_1 FILLER_62_431 ();
 sg13g2_fill_2 FILLER_62_441 ();
 sg13g2_fill_1 FILLER_62_443 ();
 sg13g2_fill_2 FILLER_62_449 ();
 sg13g2_fill_1 FILLER_62_451 ();
 sg13g2_fill_1 FILLER_62_457 ();
 sg13g2_fill_2 FILLER_62_471 ();
 sg13g2_fill_1 FILLER_62_473 ();
 sg13g2_fill_2 FILLER_62_478 ();
 sg13g2_fill_1 FILLER_62_480 ();
 sg13g2_decap_8 FILLER_62_513 ();
 sg13g2_decap_8 FILLER_62_520 ();
 sg13g2_fill_1 FILLER_62_546 ();
 sg13g2_fill_2 FILLER_62_552 ();
 sg13g2_fill_1 FILLER_62_554 ();
 sg13g2_fill_1 FILLER_62_582 ();
 sg13g2_fill_2 FILLER_62_600 ();
 sg13g2_fill_1 FILLER_62_602 ();
 sg13g2_decap_8 FILLER_62_631 ();
 sg13g2_fill_1 FILLER_62_642 ();
 sg13g2_fill_1 FILLER_62_647 ();
 sg13g2_fill_2 FILLER_62_708 ();
 sg13g2_fill_1 FILLER_62_710 ();
 sg13g2_fill_2 FILLER_62_715 ();
 sg13g2_fill_1 FILLER_62_727 ();
 sg13g2_decap_4 FILLER_62_737 ();
 sg13g2_fill_2 FILLER_62_741 ();
 sg13g2_fill_2 FILLER_62_747 ();
 sg13g2_fill_1 FILLER_62_786 ();
 sg13g2_fill_2 FILLER_62_791 ();
 sg13g2_decap_8 FILLER_62_806 ();
 sg13g2_decap_8 FILLER_62_813 ();
 sg13g2_decap_8 FILLER_62_820 ();
 sg13g2_decap_8 FILLER_62_827 ();
 sg13g2_decap_8 FILLER_62_834 ();
 sg13g2_decap_8 FILLER_62_841 ();
 sg13g2_decap_8 FILLER_62_848 ();
 sg13g2_decap_8 FILLER_62_855 ();
 sg13g2_fill_2 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_45 ();
 sg13g2_fill_2 FILLER_63_91 ();
 sg13g2_fill_2 FILLER_63_153 ();
 sg13g2_fill_1 FILLER_63_155 ();
 sg13g2_fill_2 FILLER_63_201 ();
 sg13g2_decap_8 FILLER_63_207 ();
 sg13g2_fill_2 FILLER_63_214 ();
 sg13g2_fill_1 FILLER_63_216 ();
 sg13g2_decap_4 FILLER_63_226 ();
 sg13g2_fill_2 FILLER_63_230 ();
 sg13g2_fill_1 FILLER_63_248 ();
 sg13g2_fill_2 FILLER_63_258 ();
 sg13g2_decap_8 FILLER_63_304 ();
 sg13g2_decap_8 FILLER_63_311 ();
 sg13g2_fill_1 FILLER_63_322 ();
 sg13g2_fill_1 FILLER_63_337 ();
 sg13g2_fill_2 FILLER_63_370 ();
 sg13g2_fill_1 FILLER_63_372 ();
 sg13g2_fill_2 FILLER_63_378 ();
 sg13g2_fill_1 FILLER_63_388 ();
 sg13g2_decap_4 FILLER_63_409 ();
 sg13g2_fill_1 FILLER_63_484 ();
 sg13g2_fill_2 FILLER_63_498 ();
 sg13g2_fill_1 FILLER_63_500 ();
 sg13g2_decap_8 FILLER_63_514 ();
 sg13g2_decap_8 FILLER_63_521 ();
 sg13g2_decap_4 FILLER_63_532 ();
 sg13g2_fill_2 FILLER_63_546 ();
 sg13g2_fill_1 FILLER_63_548 ();
 sg13g2_decap_4 FILLER_63_554 ();
 sg13g2_fill_1 FILLER_63_558 ();
 sg13g2_decap_8 FILLER_63_569 ();
 sg13g2_decap_4 FILLER_63_576 ();
 sg13g2_fill_1 FILLER_63_580 ();
 sg13g2_fill_1 FILLER_63_593 ();
 sg13g2_fill_2 FILLER_63_603 ();
 sg13g2_fill_1 FILLER_63_605 ();
 sg13g2_fill_2 FILLER_63_637 ();
 sg13g2_fill_2 FILLER_63_673 ();
 sg13g2_fill_1 FILLER_63_757 ();
 sg13g2_fill_2 FILLER_63_774 ();
 sg13g2_fill_2 FILLER_63_786 ();
 sg13g2_decap_8 FILLER_63_818 ();
 sg13g2_decap_8 FILLER_63_825 ();
 sg13g2_decap_8 FILLER_63_832 ();
 sg13g2_decap_8 FILLER_63_839 ();
 sg13g2_decap_8 FILLER_63_846 ();
 sg13g2_decap_8 FILLER_63_853 ();
 sg13g2_fill_2 FILLER_63_860 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_4 FILLER_64_15 ();
 sg13g2_fill_1 FILLER_64_60 ();
 sg13g2_decap_4 FILLER_64_65 ();
 sg13g2_fill_1 FILLER_64_69 ();
 sg13g2_fill_2 FILLER_64_87 ();
 sg13g2_fill_1 FILLER_64_89 ();
 sg13g2_fill_2 FILLER_64_102 ();
 sg13g2_fill_2 FILLER_64_145 ();
 sg13g2_fill_2 FILLER_64_156 ();
 sg13g2_fill_1 FILLER_64_158 ();
 sg13g2_fill_1 FILLER_64_169 ();
 sg13g2_fill_2 FILLER_64_187 ();
 sg13g2_decap_8 FILLER_64_194 ();
 sg13g2_fill_1 FILLER_64_201 ();
 sg13g2_fill_2 FILLER_64_210 ();
 sg13g2_fill_1 FILLER_64_212 ();
 sg13g2_decap_4 FILLER_64_221 ();
 sg13g2_decap_8 FILLER_64_270 ();
 sg13g2_decap_4 FILLER_64_277 ();
 sg13g2_fill_2 FILLER_64_281 ();
 sg13g2_fill_2 FILLER_64_366 ();
 sg13g2_fill_1 FILLER_64_368 ();
 sg13g2_fill_2 FILLER_64_384 ();
 sg13g2_decap_8 FILLER_64_406 ();
 sg13g2_decap_4 FILLER_64_413 ();
 sg13g2_fill_2 FILLER_64_417 ();
 sg13g2_decap_8 FILLER_64_423 ();
 sg13g2_decap_4 FILLER_64_430 ();
 sg13g2_fill_1 FILLER_64_471 ();
 sg13g2_decap_4 FILLER_64_500 ();
 sg13g2_decap_8 FILLER_64_530 ();
 sg13g2_fill_2 FILLER_64_537 ();
 sg13g2_fill_1 FILLER_64_544 ();
 sg13g2_decap_4 FILLER_64_550 ();
 sg13g2_fill_2 FILLER_64_554 ();
 sg13g2_decap_8 FILLER_64_570 ();
 sg13g2_decap_4 FILLER_64_577 ();
 sg13g2_fill_2 FILLER_64_581 ();
 sg13g2_fill_2 FILLER_64_604 ();
 sg13g2_fill_2 FILLER_64_615 ();
 sg13g2_fill_1 FILLER_64_641 ();
 sg13g2_decap_4 FILLER_64_670 ();
 sg13g2_fill_1 FILLER_64_674 ();
 sg13g2_fill_1 FILLER_64_684 ();
 sg13g2_fill_1 FILLER_64_720 ();
 sg13g2_decap_4 FILLER_64_763 ();
 sg13g2_fill_1 FILLER_64_767 ();
 sg13g2_fill_2 FILLER_64_812 ();
 sg13g2_fill_1 FILLER_64_814 ();
 sg13g2_decap_8 FILLER_64_824 ();
 sg13g2_decap_8 FILLER_64_831 ();
 sg13g2_decap_8 FILLER_64_838 ();
 sg13g2_decap_8 FILLER_64_845 ();
 sg13g2_decap_8 FILLER_64_852 ();
 sg13g2_fill_2 FILLER_64_859 ();
 sg13g2_fill_1 FILLER_64_861 ();
 sg13g2_decap_4 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_4 ();
 sg13g2_fill_2 FILLER_65_50 ();
 sg13g2_decap_4 FILLER_65_56 ();
 sg13g2_fill_2 FILLER_65_88 ();
 sg13g2_fill_1 FILLER_65_104 ();
 sg13g2_fill_2 FILLER_65_109 ();
 sg13g2_decap_8 FILLER_65_120 ();
 sg13g2_decap_8 FILLER_65_127 ();
 sg13g2_decap_8 FILLER_65_134 ();
 sg13g2_decap_4 FILLER_65_141 ();
 sg13g2_fill_2 FILLER_65_145 ();
 sg13g2_decap_8 FILLER_65_164 ();
 sg13g2_fill_1 FILLER_65_171 ();
 sg13g2_decap_8 FILLER_65_176 ();
 sg13g2_decap_8 FILLER_65_183 ();
 sg13g2_decap_4 FILLER_65_190 ();
 sg13g2_decap_8 FILLER_65_212 ();
 sg13g2_decap_4 FILLER_65_219 ();
 sg13g2_fill_2 FILLER_65_223 ();
 sg13g2_decap_8 FILLER_65_252 ();
 sg13g2_decap_4 FILLER_65_320 ();
 sg13g2_fill_1 FILLER_65_324 ();
 sg13g2_decap_8 FILLER_65_329 ();
 sg13g2_decap_4 FILLER_65_336 ();
 sg13g2_fill_1 FILLER_65_340 ();
 sg13g2_decap_4 FILLER_65_362 ();
 sg13g2_decap_4 FILLER_65_403 ();
 sg13g2_fill_1 FILLER_65_407 ();
 sg13g2_fill_2 FILLER_65_427 ();
 sg13g2_fill_2 FILLER_65_452 ();
 sg13g2_fill_1 FILLER_65_474 ();
 sg13g2_decap_4 FILLER_65_503 ();
 sg13g2_fill_2 FILLER_65_519 ();
 sg13g2_fill_1 FILLER_65_521 ();
 sg13g2_decap_4 FILLER_65_540 ();
 sg13g2_fill_1 FILLER_65_544 ();
 sg13g2_decap_8 FILLER_65_551 ();
 sg13g2_fill_2 FILLER_65_558 ();
 sg13g2_fill_1 FILLER_65_560 ();
 sg13g2_decap_8 FILLER_65_585 ();
 sg13g2_fill_2 FILLER_65_638 ();
 sg13g2_fill_2 FILLER_65_662 ();
 sg13g2_fill_1 FILLER_65_664 ();
 sg13g2_fill_2 FILLER_65_674 ();
 sg13g2_fill_2 FILLER_65_703 ();
 sg13g2_fill_2 FILLER_65_755 ();
 sg13g2_fill_1 FILLER_65_757 ();
 sg13g2_decap_8 FILLER_65_782 ();
 sg13g2_fill_1 FILLER_65_789 ();
 sg13g2_decap_8 FILLER_65_803 ();
 sg13g2_decap_8 FILLER_65_810 ();
 sg13g2_decap_8 FILLER_65_817 ();
 sg13g2_decap_8 FILLER_65_824 ();
 sg13g2_decap_8 FILLER_65_831 ();
 sg13g2_decap_8 FILLER_65_838 ();
 sg13g2_decap_8 FILLER_65_845 ();
 sg13g2_decap_8 FILLER_65_852 ();
 sg13g2_fill_2 FILLER_65_859 ();
 sg13g2_fill_1 FILLER_65_861 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_35 ();
 sg13g2_fill_1 FILLER_66_37 ();
 sg13g2_fill_2 FILLER_66_83 ();
 sg13g2_fill_1 FILLER_66_85 ();
 sg13g2_decap_4 FILLER_66_126 ();
 sg13g2_fill_2 FILLER_66_130 ();
 sg13g2_fill_2 FILLER_66_143 ();
 sg13g2_decap_8 FILLER_66_161 ();
 sg13g2_fill_2 FILLER_66_182 ();
 sg13g2_fill_1 FILLER_66_213 ();
 sg13g2_decap_8 FILLER_66_222 ();
 sg13g2_fill_1 FILLER_66_229 ();
 sg13g2_decap_4 FILLER_66_234 ();
 sg13g2_fill_1 FILLER_66_238 ();
 sg13g2_decap_8 FILLER_66_252 ();
 sg13g2_fill_1 FILLER_66_259 ();
 sg13g2_fill_1 FILLER_66_268 ();
 sg13g2_fill_2 FILLER_66_300 ();
 sg13g2_fill_2 FILLER_66_332 ();
 sg13g2_fill_2 FILLER_66_350 ();
 sg13g2_decap_8 FILLER_66_366 ();
 sg13g2_decap_4 FILLER_66_373 ();
 sg13g2_fill_1 FILLER_66_377 ();
 sg13g2_fill_2 FILLER_66_391 ();
 sg13g2_decap_4 FILLER_66_397 ();
 sg13g2_fill_1 FILLER_66_401 ();
 sg13g2_decap_8 FILLER_66_425 ();
 sg13g2_fill_1 FILLER_66_438 ();
 sg13g2_fill_2 FILLER_66_445 ();
 sg13g2_fill_1 FILLER_66_447 ();
 sg13g2_decap_4 FILLER_66_473 ();
 sg13g2_fill_1 FILLER_66_477 ();
 sg13g2_fill_2 FILLER_66_488 ();
 sg13g2_fill_1 FILLER_66_490 ();
 sg13g2_fill_2 FILLER_66_497 ();
 sg13g2_fill_1 FILLER_66_499 ();
 sg13g2_decap_8 FILLER_66_507 ();
 sg13g2_decap_4 FILLER_66_514 ();
 sg13g2_fill_2 FILLER_66_533 ();
 sg13g2_fill_2 FILLER_66_548 ();
 sg13g2_fill_1 FILLER_66_550 ();
 sg13g2_fill_2 FILLER_66_556 ();
 sg13g2_fill_1 FILLER_66_558 ();
 sg13g2_decap_8 FILLER_66_577 ();
 sg13g2_fill_2 FILLER_66_584 ();
 sg13g2_fill_1 FILLER_66_586 ();
 sg13g2_fill_2 FILLER_66_614 ();
 sg13g2_fill_2 FILLER_66_673 ();
 sg13g2_fill_2 FILLER_66_684 ();
 sg13g2_fill_1 FILLER_66_686 ();
 sg13g2_fill_2 FILLER_66_710 ();
 sg13g2_fill_2 FILLER_66_729 ();
 sg13g2_decap_8 FILLER_66_788 ();
 sg13g2_decap_8 FILLER_66_795 ();
 sg13g2_decap_8 FILLER_66_802 ();
 sg13g2_decap_8 FILLER_66_809 ();
 sg13g2_decap_8 FILLER_66_816 ();
 sg13g2_decap_8 FILLER_66_823 ();
 sg13g2_decap_8 FILLER_66_830 ();
 sg13g2_decap_8 FILLER_66_837 ();
 sg13g2_decap_8 FILLER_66_844 ();
 sg13g2_decap_8 FILLER_66_851 ();
 sg13g2_decap_4 FILLER_66_858 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_4 FILLER_67_7 ();
 sg13g2_fill_1 FILLER_67_11 ();
 sg13g2_decap_8 FILLER_67_16 ();
 sg13g2_decap_4 FILLER_67_23 ();
 sg13g2_fill_1 FILLER_67_27 ();
 sg13g2_fill_1 FILLER_67_63 ();
 sg13g2_fill_2 FILLER_67_132 ();
 sg13g2_fill_1 FILLER_67_147 ();
 sg13g2_decap_8 FILLER_67_184 ();
 sg13g2_fill_2 FILLER_67_191 ();
 sg13g2_fill_1 FILLER_67_193 ();
 sg13g2_decap_8 FILLER_67_212 ();
 sg13g2_decap_8 FILLER_67_219 ();
 sg13g2_decap_8 FILLER_67_226 ();
 sg13g2_decap_8 FILLER_67_233 ();
 sg13g2_fill_1 FILLER_67_240 ();
 sg13g2_fill_1 FILLER_67_282 ();
 sg13g2_fill_2 FILLER_67_337 ();
 sg13g2_fill_2 FILLER_67_352 ();
 sg13g2_fill_1 FILLER_67_381 ();
 sg13g2_fill_2 FILLER_67_396 ();
 sg13g2_decap_4 FILLER_67_407 ();
 sg13g2_fill_1 FILLER_67_411 ();
 sg13g2_fill_1 FILLER_67_453 ();
 sg13g2_decap_4 FILLER_67_469 ();
 sg13g2_fill_2 FILLER_67_473 ();
 sg13g2_fill_2 FILLER_67_498 ();
 sg13g2_decap_8 FILLER_67_504 ();
 sg13g2_decap_4 FILLER_67_511 ();
 sg13g2_fill_1 FILLER_67_515 ();
 sg13g2_decap_4 FILLER_67_542 ();
 sg13g2_fill_2 FILLER_67_546 ();
 sg13g2_decap_8 FILLER_67_576 ();
 sg13g2_fill_2 FILLER_67_583 ();
 sg13g2_fill_2 FILLER_67_616 ();
 sg13g2_fill_1 FILLER_67_627 ();
 sg13g2_fill_1 FILLER_67_654 ();
 sg13g2_fill_2 FILLER_67_668 ();
 sg13g2_decap_4 FILLER_67_730 ();
 sg13g2_fill_2 FILLER_67_734 ();
 sg13g2_fill_2 FILLER_67_740 ();
 sg13g2_fill_1 FILLER_67_742 ();
 sg13g2_decap_4 FILLER_67_747 ();
 sg13g2_fill_2 FILLER_67_751 ();
 sg13g2_fill_2 FILLER_67_761 ();
 sg13g2_decap_8 FILLER_67_798 ();
 sg13g2_decap_8 FILLER_67_805 ();
 sg13g2_decap_8 FILLER_67_812 ();
 sg13g2_decap_8 FILLER_67_819 ();
 sg13g2_decap_8 FILLER_67_826 ();
 sg13g2_decap_8 FILLER_67_833 ();
 sg13g2_decap_8 FILLER_67_840 ();
 sg13g2_decap_8 FILLER_67_847 ();
 sg13g2_decap_8 FILLER_67_854 ();
 sg13g2_fill_1 FILLER_67_861 ();
 sg13g2_decap_4 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_72 ();
 sg13g2_fill_1 FILLER_68_74 ();
 sg13g2_fill_2 FILLER_68_89 ();
 sg13g2_fill_2 FILLER_68_99 ();
 sg13g2_fill_1 FILLER_68_101 ();
 sg13g2_fill_1 FILLER_68_115 ();
 sg13g2_decap_4 FILLER_68_121 ();
 sg13g2_fill_1 FILLER_68_125 ();
 sg13g2_decap_8 FILLER_68_130 ();
 sg13g2_decap_8 FILLER_68_137 ();
 sg13g2_decap_8 FILLER_68_144 ();
 sg13g2_fill_2 FILLER_68_151 ();
 sg13g2_fill_1 FILLER_68_153 ();
 sg13g2_decap_8 FILLER_68_158 ();
 sg13g2_fill_1 FILLER_68_175 ();
 sg13g2_decap_8 FILLER_68_181 ();
 sg13g2_fill_1 FILLER_68_188 ();
 sg13g2_decap_8 FILLER_68_199 ();
 sg13g2_decap_8 FILLER_68_206 ();
 sg13g2_decap_4 FILLER_68_241 ();
 sg13g2_fill_1 FILLER_68_245 ();
 sg13g2_fill_1 FILLER_68_259 ();
 sg13g2_fill_1 FILLER_68_278 ();
 sg13g2_fill_2 FILLER_68_332 ();
 sg13g2_fill_1 FILLER_68_334 ();
 sg13g2_decap_4 FILLER_68_355 ();
 sg13g2_fill_1 FILLER_68_359 ();
 sg13g2_fill_2 FILLER_68_368 ();
 sg13g2_fill_1 FILLER_68_370 ();
 sg13g2_fill_1 FILLER_68_416 ();
 sg13g2_decap_8 FILLER_68_421 ();
 sg13g2_decap_8 FILLER_68_428 ();
 sg13g2_decap_8 FILLER_68_470 ();
 sg13g2_fill_2 FILLER_68_477 ();
 sg13g2_fill_2 FILLER_68_497 ();
 sg13g2_fill_2 FILLER_68_526 ();
 sg13g2_decap_8 FILLER_68_532 ();
 sg13g2_decap_4 FILLER_68_539 ();
 sg13g2_fill_1 FILLER_68_543 ();
 sg13g2_fill_1 FILLER_68_547 ();
 sg13g2_fill_2 FILLER_68_590 ();
 sg13g2_fill_1 FILLER_68_592 ();
 sg13g2_fill_2 FILLER_68_606 ();
 sg13g2_fill_2 FILLER_68_613 ();
 sg13g2_fill_2 FILLER_68_686 ();
 sg13g2_decap_8 FILLER_68_721 ();
 sg13g2_fill_2 FILLER_68_728 ();
 sg13g2_decap_8 FILLER_68_808 ();
 sg13g2_decap_8 FILLER_68_815 ();
 sg13g2_decap_8 FILLER_68_822 ();
 sg13g2_decap_8 FILLER_68_829 ();
 sg13g2_decap_8 FILLER_68_836 ();
 sg13g2_decap_8 FILLER_68_843 ();
 sg13g2_decap_8 FILLER_68_850 ();
 sg13g2_decap_4 FILLER_68_857 ();
 sg13g2_fill_1 FILLER_68_861 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_7 ();
 sg13g2_fill_2 FILLER_69_17 ();
 sg13g2_fill_1 FILLER_69_19 ();
 sg13g2_fill_2 FILLER_69_41 ();
 sg13g2_fill_1 FILLER_69_43 ();
 sg13g2_fill_1 FILLER_69_76 ();
 sg13g2_decap_8 FILLER_69_149 ();
 sg13g2_fill_1 FILLER_69_156 ();
 sg13g2_decap_4 FILLER_69_189 ();
 sg13g2_fill_1 FILLER_69_193 ();
 sg13g2_decap_8 FILLER_69_199 ();
 sg13g2_decap_4 FILLER_69_210 ();
 sg13g2_fill_1 FILLER_69_214 ();
 sg13g2_fill_2 FILLER_69_269 ();
 sg13g2_fill_1 FILLER_69_307 ();
 sg13g2_fill_1 FILLER_69_323 ();
 sg13g2_decap_4 FILLER_69_342 ();
 sg13g2_decap_8 FILLER_69_369 ();
 sg13g2_fill_2 FILLER_69_381 ();
 sg13g2_fill_1 FILLER_69_400 ();
 sg13g2_decap_8 FILLER_69_414 ();
 sg13g2_decap_8 FILLER_69_421 ();
 sg13g2_decap_4 FILLER_69_428 ();
 sg13g2_decap_4 FILLER_69_436 ();
 sg13g2_decap_4 FILLER_69_481 ();
 sg13g2_fill_2 FILLER_69_504 ();
 sg13g2_decap_4 FILLER_69_534 ();
 sg13g2_decap_4 FILLER_69_556 ();
 sg13g2_fill_2 FILLER_69_586 ();
 sg13g2_fill_2 FILLER_69_638 ();
 sg13g2_fill_1 FILLER_69_640 ();
 sg13g2_fill_1 FILLER_69_650 ();
 sg13g2_decap_4 FILLER_69_659 ();
 sg13g2_fill_1 FILLER_69_663 ();
 sg13g2_decap_8 FILLER_69_668 ();
 sg13g2_fill_2 FILLER_69_675 ();
 sg13g2_decap_4 FILLER_69_681 ();
 sg13g2_fill_1 FILLER_69_685 ();
 sg13g2_fill_1 FILLER_69_694 ();
 sg13g2_decap_8 FILLER_69_722 ();
 sg13g2_decap_4 FILLER_69_729 ();
 sg13g2_fill_2 FILLER_69_733 ();
 sg13g2_fill_1 FILLER_69_739 ();
 sg13g2_decap_4 FILLER_69_744 ();
 sg13g2_fill_1 FILLER_69_748 ();
 sg13g2_fill_1 FILLER_69_784 ();
 sg13g2_decap_8 FILLER_69_816 ();
 sg13g2_decap_8 FILLER_69_823 ();
 sg13g2_decap_8 FILLER_69_830 ();
 sg13g2_decap_8 FILLER_69_837 ();
 sg13g2_decap_8 FILLER_69_844 ();
 sg13g2_decap_8 FILLER_69_851 ();
 sg13g2_decap_4 FILLER_69_858 ();
 sg13g2_fill_2 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_2 ();
 sg13g2_fill_2 FILLER_70_52 ();
 sg13g2_fill_1 FILLER_70_54 ();
 sg13g2_fill_1 FILLER_70_96 ();
 sg13g2_fill_2 FILLER_70_110 ();
 sg13g2_fill_2 FILLER_70_129 ();
 sg13g2_fill_1 FILLER_70_159 ();
 sg13g2_decap_4 FILLER_70_193 ();
 sg13g2_fill_1 FILLER_70_197 ();
 sg13g2_decap_4 FILLER_70_216 ();
 sg13g2_fill_2 FILLER_70_220 ();
 sg13g2_fill_1 FILLER_70_231 ();
 sg13g2_decap_8 FILLER_70_245 ();
 sg13g2_fill_2 FILLER_70_252 ();
 sg13g2_fill_2 FILLER_70_268 ();
 sg13g2_fill_1 FILLER_70_296 ();
 sg13g2_decap_8 FILLER_70_313 ();
 sg13g2_decap_8 FILLER_70_320 ();
 sg13g2_decap_4 FILLER_70_327 ();
 sg13g2_decap_8 FILLER_70_365 ();
 sg13g2_decap_8 FILLER_70_372 ();
 sg13g2_fill_1 FILLER_70_379 ();
 sg13g2_fill_2 FILLER_70_390 ();
 sg13g2_fill_2 FILLER_70_441 ();
 sg13g2_fill_1 FILLER_70_443 ();
 sg13g2_decap_4 FILLER_70_458 ();
 sg13g2_fill_2 FILLER_70_462 ();
 sg13g2_fill_1 FILLER_70_505 ();
 sg13g2_fill_2 FILLER_70_542 ();
 sg13g2_fill_1 FILLER_70_544 ();
 sg13g2_decap_4 FILLER_70_576 ();
 sg13g2_fill_2 FILLER_70_580 ();
 sg13g2_fill_1 FILLER_70_595 ();
 sg13g2_fill_1 FILLER_70_609 ();
 sg13g2_fill_2 FILLER_70_624 ();
 sg13g2_fill_2 FILLER_70_654 ();
 sg13g2_fill_2 FILLER_70_688 ();
 sg13g2_decap_4 FILLER_70_695 ();
 sg13g2_fill_2 FILLER_70_707 ();
 sg13g2_fill_2 FILLER_70_737 ();
 sg13g2_fill_1 FILLER_70_795 ();
 sg13g2_decap_8 FILLER_70_824 ();
 sg13g2_decap_8 FILLER_70_831 ();
 sg13g2_decap_8 FILLER_70_838 ();
 sg13g2_decap_8 FILLER_70_845 ();
 sg13g2_decap_8 FILLER_70_852 ();
 sg13g2_fill_2 FILLER_70_859 ();
 sg13g2_fill_1 FILLER_70_861 ();
 sg13g2_decap_4 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_4 ();
 sg13g2_fill_1 FILLER_71_32 ();
 sg13g2_fill_2 FILLER_71_65 ();
 sg13g2_fill_1 FILLER_71_81 ();
 sg13g2_fill_2 FILLER_71_91 ();
 sg13g2_fill_2 FILLER_71_102 ();
 sg13g2_fill_1 FILLER_71_131 ();
 sg13g2_decap_8 FILLER_71_154 ();
 sg13g2_fill_2 FILLER_71_161 ();
 sg13g2_decap_8 FILLER_71_187 ();
 sg13g2_fill_1 FILLER_71_194 ();
 sg13g2_fill_2 FILLER_71_218 ();
 sg13g2_fill_1 FILLER_71_220 ();
 sg13g2_fill_2 FILLER_71_239 ();
 sg13g2_fill_1 FILLER_71_241 ();
 sg13g2_decap_4 FILLER_71_246 ();
 sg13g2_fill_2 FILLER_71_264 ();
 sg13g2_fill_1 FILLER_71_266 ();
 sg13g2_fill_2 FILLER_71_286 ();
 sg13g2_fill_1 FILLER_71_288 ();
 sg13g2_decap_8 FILLER_71_304 ();
 sg13g2_decap_8 FILLER_71_324 ();
 sg13g2_decap_4 FILLER_71_331 ();
 sg13g2_decap_4 FILLER_71_347 ();
 sg13g2_decap_4 FILLER_71_366 ();
 sg13g2_fill_2 FILLER_71_370 ();
 sg13g2_decap_8 FILLER_71_392 ();
 sg13g2_fill_2 FILLER_71_399 ();
 sg13g2_fill_1 FILLER_71_401 ();
 sg13g2_decap_8 FILLER_71_427 ();
 sg13g2_fill_2 FILLER_71_434 ();
 sg13g2_fill_1 FILLER_71_436 ();
 sg13g2_fill_1 FILLER_71_468 ();
 sg13g2_fill_2 FILLER_71_477 ();
 sg13g2_fill_1 FILLER_71_532 ();
 sg13g2_decap_4 FILLER_71_537 ();
 sg13g2_decap_8 FILLER_71_567 ();
 sg13g2_decap_4 FILLER_71_574 ();
 sg13g2_fill_2 FILLER_71_578 ();
 sg13g2_fill_2 FILLER_71_616 ();
 sg13g2_fill_1 FILLER_71_618 ();
 sg13g2_fill_2 FILLER_71_636 ();
 sg13g2_fill_1 FILLER_71_638 ();
 sg13g2_fill_2 FILLER_71_652 ();
 sg13g2_fill_2 FILLER_71_667 ();
 sg13g2_fill_1 FILLER_71_677 ();
 sg13g2_fill_1 FILLER_71_714 ();
 sg13g2_decap_4 FILLER_71_719 ();
 sg13g2_decap_4 FILLER_71_732 ();
 sg13g2_fill_1 FILLER_71_778 ();
 sg13g2_decap_8 FILLER_71_829 ();
 sg13g2_decap_8 FILLER_71_836 ();
 sg13g2_decap_8 FILLER_71_843 ();
 sg13g2_decap_8 FILLER_71_850 ();
 sg13g2_decap_4 FILLER_71_857 ();
 sg13g2_fill_1 FILLER_71_861 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_7 ();
 sg13g2_fill_1 FILLER_72_9 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_fill_2 FILLER_72_21 ();
 sg13g2_fill_1 FILLER_72_42 ();
 sg13g2_fill_2 FILLER_72_47 ();
 sg13g2_fill_1 FILLER_72_58 ();
 sg13g2_fill_1 FILLER_72_105 ();
 sg13g2_fill_2 FILLER_72_114 ();
 sg13g2_fill_1 FILLER_72_116 ();
 sg13g2_fill_2 FILLER_72_147 ();
 sg13g2_fill_1 FILLER_72_149 ();
 sg13g2_decap_8 FILLER_72_154 ();
 sg13g2_decap_8 FILLER_72_177 ();
 sg13g2_decap_8 FILLER_72_184 ();
 sg13g2_fill_2 FILLER_72_191 ();
 sg13g2_decap_4 FILLER_72_233 ();
 sg13g2_fill_1 FILLER_72_277 ();
 sg13g2_fill_2 FILLER_72_290 ();
 sg13g2_fill_1 FILLER_72_292 ();
 sg13g2_decap_8 FILLER_72_316 ();
 sg13g2_fill_2 FILLER_72_323 ();
 sg13g2_fill_2 FILLER_72_355 ();
 sg13g2_fill_1 FILLER_72_357 ();
 sg13g2_decap_8 FILLER_72_367 ();
 sg13g2_fill_2 FILLER_72_374 ();
 sg13g2_fill_1 FILLER_72_394 ();
 sg13g2_fill_2 FILLER_72_433 ();
 sg13g2_decap_8 FILLER_72_452 ();
 sg13g2_fill_2 FILLER_72_459 ();
 sg13g2_fill_2 FILLER_72_506 ();
 sg13g2_fill_1 FILLER_72_517 ();
 sg13g2_fill_1 FILLER_72_523 ();
 sg13g2_fill_2 FILLER_72_537 ();
 sg13g2_fill_2 FILLER_72_575 ();
 sg13g2_fill_1 FILLER_72_590 ();
 sg13g2_fill_1 FILLER_72_613 ();
 sg13g2_fill_2 FILLER_72_663 ();
 sg13g2_fill_1 FILLER_72_665 ();
 sg13g2_decap_4 FILLER_72_696 ();
 sg13g2_fill_2 FILLER_72_709 ();
 sg13g2_fill_1 FILLER_72_711 ();
 sg13g2_fill_2 FILLER_72_759 ();
 sg13g2_fill_2 FILLER_72_777 ();
 sg13g2_fill_2 FILLER_72_792 ();
 sg13g2_fill_1 FILLER_72_794 ();
 sg13g2_decap_8 FILLER_72_836 ();
 sg13g2_decap_8 FILLER_72_843 ();
 sg13g2_decap_8 FILLER_72_850 ();
 sg13g2_decap_4 FILLER_72_857 ();
 sg13g2_fill_1 FILLER_72_861 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_fill_2 FILLER_73_56 ();
 sg13g2_fill_1 FILLER_73_99 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_4 FILLER_73_133 ();
 sg13g2_fill_1 FILLER_73_137 ();
 sg13g2_decap_4 FILLER_73_141 ();
 sg13g2_decap_4 FILLER_73_153 ();
 sg13g2_fill_2 FILLER_73_165 ();
 sg13g2_decap_8 FILLER_73_186 ();
 sg13g2_decap_8 FILLER_73_206 ();
 sg13g2_decap_4 FILLER_73_213 ();
 sg13g2_fill_2 FILLER_73_217 ();
 sg13g2_fill_2 FILLER_73_263 ();
 sg13g2_fill_2 FILLER_73_294 ();
 sg13g2_fill_1 FILLER_73_296 ();
 sg13g2_decap_8 FILLER_73_310 ();
 sg13g2_fill_2 FILLER_73_317 ();
 sg13g2_fill_1 FILLER_73_319 ();
 sg13g2_decap_4 FILLER_73_333 ();
 sg13g2_fill_2 FILLER_73_337 ();
 sg13g2_fill_2 FILLER_73_349 ();
 sg13g2_fill_2 FILLER_73_359 ();
 sg13g2_fill_1 FILLER_73_361 ();
 sg13g2_decap_4 FILLER_73_375 ();
 sg13g2_fill_2 FILLER_73_379 ();
 sg13g2_fill_2 FILLER_73_390 ();
 sg13g2_fill_2 FILLER_73_397 ();
 sg13g2_decap_4 FILLER_73_416 ();
 sg13g2_fill_2 FILLER_73_420 ();
 sg13g2_fill_2 FILLER_73_435 ();
 sg13g2_fill_1 FILLER_73_437 ();
 sg13g2_fill_2 FILLER_73_465 ();
 sg13g2_fill_1 FILLER_73_467 ();
 sg13g2_fill_1 FILLER_73_499 ();
 sg13g2_fill_2 FILLER_73_535 ();
 sg13g2_fill_1 FILLER_73_542 ();
 sg13g2_fill_2 FILLER_73_557 ();
 sg13g2_decap_8 FILLER_73_568 ();
 sg13g2_fill_2 FILLER_73_575 ();
 sg13g2_fill_1 FILLER_73_577 ();
 sg13g2_fill_1 FILLER_73_680 ();
 sg13g2_fill_2 FILLER_73_695 ();
 sg13g2_fill_1 FILLER_73_697 ();
 sg13g2_fill_2 FILLER_73_764 ();
 sg13g2_fill_2 FILLER_73_782 ();
 sg13g2_decap_8 FILLER_73_831 ();
 sg13g2_decap_8 FILLER_73_838 ();
 sg13g2_decap_8 FILLER_73_845 ();
 sg13g2_decap_8 FILLER_73_852 ();
 sg13g2_fill_2 FILLER_73_859 ();
 sg13g2_fill_1 FILLER_73_861 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_4 FILLER_74_49 ();
 sg13g2_fill_2 FILLER_74_53 ();
 sg13g2_fill_1 FILLER_74_151 ();
 sg13g2_fill_2 FILLER_74_175 ();
 sg13g2_fill_1 FILLER_74_177 ();
 sg13g2_fill_1 FILLER_74_218 ();
 sg13g2_fill_2 FILLER_74_269 ();
 sg13g2_decap_4 FILLER_74_289 ();
 sg13g2_fill_1 FILLER_74_293 ();
 sg13g2_decap_4 FILLER_74_308 ();
 sg13g2_decap_4 FILLER_74_330 ();
 sg13g2_fill_1 FILLER_74_334 ();
 sg13g2_fill_1 FILLER_74_344 ();
 sg13g2_decap_4 FILLER_74_365 ();
 sg13g2_fill_2 FILLER_74_369 ();
 sg13g2_fill_2 FILLER_74_393 ();
 sg13g2_fill_1 FILLER_74_395 ();
 sg13g2_fill_1 FILLER_74_428 ();
 sg13g2_fill_2 FILLER_74_488 ();
 sg13g2_fill_1 FILLER_74_490 ();
 sg13g2_fill_2 FILLER_74_546 ();
 sg13g2_fill_1 FILLER_74_548 ();
 sg13g2_fill_1 FILLER_74_576 ();
 sg13g2_fill_2 FILLER_74_582 ();
 sg13g2_fill_1 FILLER_74_584 ();
 sg13g2_fill_1 FILLER_74_603 ();
 sg13g2_fill_2 FILLER_74_644 ();
 sg13g2_fill_1 FILLER_74_646 ();
 sg13g2_fill_1 FILLER_74_651 ();
 sg13g2_fill_1 FILLER_74_666 ();
 sg13g2_fill_2 FILLER_74_685 ();
 sg13g2_fill_1 FILLER_74_687 ();
 sg13g2_fill_2 FILLER_74_701 ();
 sg13g2_decap_8 FILLER_74_707 ();
 sg13g2_fill_2 FILLER_74_714 ();
 sg13g2_fill_1 FILLER_74_716 ();
 sg13g2_fill_2 FILLER_74_787 ();
 sg13g2_fill_1 FILLER_74_789 ();
 sg13g2_decap_8 FILLER_74_826 ();
 sg13g2_decap_8 FILLER_74_833 ();
 sg13g2_decap_8 FILLER_74_840 ();
 sg13g2_decap_8 FILLER_74_847 ();
 sg13g2_decap_8 FILLER_74_854 ();
 sg13g2_fill_1 FILLER_74_861 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_fill_2 FILLER_75_49 ();
 sg13g2_fill_2 FILLER_75_78 ();
 sg13g2_fill_1 FILLER_75_112 ();
 sg13g2_fill_2 FILLER_75_122 ();
 sg13g2_fill_2 FILLER_75_133 ();
 sg13g2_fill_1 FILLER_75_135 ();
 sg13g2_decap_4 FILLER_75_142 ();
 sg13g2_fill_2 FILLER_75_168 ();
 sg13g2_fill_1 FILLER_75_170 ();
 sg13g2_fill_2 FILLER_75_202 ();
 sg13g2_decap_4 FILLER_75_213 ();
 sg13g2_fill_2 FILLER_75_217 ();
 sg13g2_fill_2 FILLER_75_288 ();
 sg13g2_fill_1 FILLER_75_290 ();
 sg13g2_decap_4 FILLER_75_318 ();
 sg13g2_fill_2 FILLER_75_331 ();
 sg13g2_decap_4 FILLER_75_346 ();
 sg13g2_fill_1 FILLER_75_350 ();
 sg13g2_fill_2 FILLER_75_377 ();
 sg13g2_decap_8 FILLER_75_383 ();
 sg13g2_decap_8 FILLER_75_390 ();
 sg13g2_fill_1 FILLER_75_419 ();
 sg13g2_fill_2 FILLER_75_437 ();
 sg13g2_decap_8 FILLER_75_447 ();
 sg13g2_fill_2 FILLER_75_481 ();
 sg13g2_decap_4 FILLER_75_550 ();
 sg13g2_fill_2 FILLER_75_622 ();
 sg13g2_fill_2 FILLER_75_665 ();
 sg13g2_fill_1 FILLER_75_690 ();
 sg13g2_fill_2 FILLER_75_727 ();
 sg13g2_fill_1 FILLER_75_729 ();
 sg13g2_fill_1 FILLER_75_799 ();
 sg13g2_decap_8 FILLER_75_818 ();
 sg13g2_decap_8 FILLER_75_825 ();
 sg13g2_decap_8 FILLER_75_832 ();
 sg13g2_decap_8 FILLER_75_839 ();
 sg13g2_decap_8 FILLER_75_846 ();
 sg13g2_decap_8 FILLER_75_853 ();
 sg13g2_fill_2 FILLER_75_860 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_fill_2 FILLER_76_56 ();
 sg13g2_fill_2 FILLER_76_86 ();
 sg13g2_decap_4 FILLER_76_115 ();
 sg13g2_fill_2 FILLER_76_119 ();
 sg13g2_fill_2 FILLER_76_147 ();
 sg13g2_fill_1 FILLER_76_149 ();
 sg13g2_fill_1 FILLER_76_155 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_fill_1 FILLER_76_168 ();
 sg13g2_fill_1 FILLER_76_174 ();
 sg13g2_fill_2 FILLER_76_213 ();
 sg13g2_decap_4 FILLER_76_222 ();
 sg13g2_fill_2 FILLER_76_277 ();
 sg13g2_decap_4 FILLER_76_347 ();
 sg13g2_decap_8 FILLER_76_372 ();
 sg13g2_decap_8 FILLER_76_379 ();
 sg13g2_fill_1 FILLER_76_386 ();
 sg13g2_fill_1 FILLER_76_391 ();
 sg13g2_decap_8 FILLER_76_451 ();
 sg13g2_fill_1 FILLER_76_458 ();
 sg13g2_fill_1 FILLER_76_463 ();
 sg13g2_fill_2 FILLER_76_514 ();
 sg13g2_fill_1 FILLER_76_532 ();
 sg13g2_decap_8 FILLER_76_537 ();
 sg13g2_decap_4 FILLER_76_544 ();
 sg13g2_fill_2 FILLER_76_548 ();
 sg13g2_fill_2 FILLER_76_567 ();
 sg13g2_fill_2 FILLER_76_595 ();
 sg13g2_fill_1 FILLER_76_597 ();
 sg13g2_fill_1 FILLER_76_615 ();
 sg13g2_fill_2 FILLER_76_626 ();
 sg13g2_fill_1 FILLER_76_628 ();
 sg13g2_decap_4 FILLER_76_642 ();
 sg13g2_fill_2 FILLER_76_646 ();
 sg13g2_decap_4 FILLER_76_652 ();
 sg13g2_fill_1 FILLER_76_661 ();
 sg13g2_fill_2 FILLER_76_667 ();
 sg13g2_decap_4 FILLER_76_700 ();
 sg13g2_fill_2 FILLER_76_704 ();
 sg13g2_fill_1 FILLER_76_710 ();
 sg13g2_fill_1 FILLER_76_756 ();
 sg13g2_fill_1 FILLER_76_761 ();
 sg13g2_fill_2 FILLER_76_771 ();
 sg13g2_decap_8 FILLER_76_813 ();
 sg13g2_decap_8 FILLER_76_820 ();
 sg13g2_decap_8 FILLER_76_827 ();
 sg13g2_decap_8 FILLER_76_834 ();
 sg13g2_decap_8 FILLER_76_841 ();
 sg13g2_decap_8 FILLER_76_848 ();
 sg13g2_decap_8 FILLER_76_855 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_67 ();
 sg13g2_fill_2 FILLER_77_129 ();
 sg13g2_fill_2 FILLER_77_152 ();
 sg13g2_fill_1 FILLER_77_154 ();
 sg13g2_decap_4 FILLER_77_168 ();
 sg13g2_fill_2 FILLER_77_172 ();
 sg13g2_fill_1 FILLER_77_195 ();
 sg13g2_fill_2 FILLER_77_204 ();
 sg13g2_fill_1 FILLER_77_206 ();
 sg13g2_fill_1 FILLER_77_221 ();
 sg13g2_decap_8 FILLER_77_231 ();
 sg13g2_fill_2 FILLER_77_238 ();
 sg13g2_fill_2 FILLER_77_272 ();
 sg13g2_fill_2 FILLER_77_290 ();
 sg13g2_fill_1 FILLER_77_292 ();
 sg13g2_fill_2 FILLER_77_311 ();
 sg13g2_fill_1 FILLER_77_313 ();
 sg13g2_fill_2 FILLER_77_337 ();
 sg13g2_decap_8 FILLER_77_352 ();
 sg13g2_decap_4 FILLER_77_364 ();
 sg13g2_fill_1 FILLER_77_368 ();
 sg13g2_decap_8 FILLER_77_373 ();
 sg13g2_fill_2 FILLER_77_380 ();
 sg13g2_fill_1 FILLER_77_409 ();
 sg13g2_fill_2 FILLER_77_440 ();
 sg13g2_fill_2 FILLER_77_450 ();
 sg13g2_fill_1 FILLER_77_452 ();
 sg13g2_fill_1 FILLER_77_527 ();
 sg13g2_fill_2 FILLER_77_555 ();
 sg13g2_fill_1 FILLER_77_627 ();
 sg13g2_fill_1 FILLER_77_655 ();
 sg13g2_decap_8 FILLER_77_692 ();
 sg13g2_decap_8 FILLER_77_699 ();
 sg13g2_decap_4 FILLER_77_706 ();
 sg13g2_fill_1 FILLER_77_710 ();
 sg13g2_decap_8 FILLER_77_724 ();
 sg13g2_decap_8 FILLER_77_731 ();
 sg13g2_decap_4 FILLER_77_742 ();
 sg13g2_fill_1 FILLER_77_746 ();
 sg13g2_decap_4 FILLER_77_774 ();
 sg13g2_fill_2 FILLER_77_782 ();
 sg13g2_fill_1 FILLER_77_784 ();
 sg13g2_fill_2 FILLER_77_789 ();
 sg13g2_fill_1 FILLER_77_791 ();
 sg13g2_fill_2 FILLER_77_797 ();
 sg13g2_decap_8 FILLER_77_803 ();
 sg13g2_decap_8 FILLER_77_810 ();
 sg13g2_decap_8 FILLER_77_817 ();
 sg13g2_decap_8 FILLER_77_824 ();
 sg13g2_decap_8 FILLER_77_831 ();
 sg13g2_decap_8 FILLER_77_838 ();
 sg13g2_decap_8 FILLER_77_845 ();
 sg13g2_decap_8 FILLER_77_852 ();
 sg13g2_fill_2 FILLER_77_859 ();
 sg13g2_fill_1 FILLER_77_861 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_fill_2 FILLER_78_104 ();
 sg13g2_fill_1 FILLER_78_106 ();
 sg13g2_fill_1 FILLER_78_135 ();
 sg13g2_fill_2 FILLER_78_165 ();
 sg13g2_fill_1 FILLER_78_176 ();
 sg13g2_fill_2 FILLER_78_191 ();
 sg13g2_fill_2 FILLER_78_239 ();
 sg13g2_fill_2 FILLER_78_277 ();
 sg13g2_decap_4 FILLER_78_311 ();
 sg13g2_fill_2 FILLER_78_361 ();
 sg13g2_fill_1 FILLER_78_363 ();
 sg13g2_fill_1 FILLER_78_391 ();
 sg13g2_fill_2 FILLER_78_439 ();
 sg13g2_fill_2 FILLER_78_467 ();
 sg13g2_fill_1 FILLER_78_469 ();
 sg13g2_fill_2 FILLER_78_521 ();
 sg13g2_fill_2 FILLER_78_532 ();
 sg13g2_fill_1 FILLER_78_627 ();
 sg13g2_fill_1 FILLER_78_641 ();
 sg13g2_fill_2 FILLER_78_659 ();
 sg13g2_decap_8 FILLER_78_665 ();
 sg13g2_decap_4 FILLER_78_672 ();
 sg13g2_decap_8 FILLER_78_689 ();
 sg13g2_decap_8 FILLER_78_696 ();
 sg13g2_decap_8 FILLER_78_703 ();
 sg13g2_decap_8 FILLER_78_710 ();
 sg13g2_decap_8 FILLER_78_717 ();
 sg13g2_decap_8 FILLER_78_724 ();
 sg13g2_decap_8 FILLER_78_731 ();
 sg13g2_decap_8 FILLER_78_738 ();
 sg13g2_decap_4 FILLER_78_745 ();
 sg13g2_decap_8 FILLER_78_757 ();
 sg13g2_fill_2 FILLER_78_764 ();
 sg13g2_decap_8 FILLER_78_775 ();
 sg13g2_decap_8 FILLER_78_782 ();
 sg13g2_decap_8 FILLER_78_793 ();
 sg13g2_decap_8 FILLER_78_800 ();
 sg13g2_decap_8 FILLER_78_807 ();
 sg13g2_decap_8 FILLER_78_814 ();
 sg13g2_decap_8 FILLER_78_821 ();
 sg13g2_decap_8 FILLER_78_828 ();
 sg13g2_decap_8 FILLER_78_835 ();
 sg13g2_decap_8 FILLER_78_842 ();
 sg13g2_decap_8 FILLER_78_849 ();
 sg13g2_decap_4 FILLER_78_856 ();
 sg13g2_fill_2 FILLER_78_860 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_94 ();
 sg13g2_decap_8 FILLER_79_101 ();
 sg13g2_decap_4 FILLER_79_108 ();
 sg13g2_fill_1 FILLER_79_112 ();
 sg13g2_decap_4 FILLER_79_117 ();
 sg13g2_fill_2 FILLER_79_121 ();
 sg13g2_decap_8 FILLER_79_230 ();
 sg13g2_decap_8 FILLER_79_237 ();
 sg13g2_fill_1 FILLER_79_293 ();
 sg13g2_fill_2 FILLER_79_334 ();
 sg13g2_fill_2 FILLER_79_349 ();
 sg13g2_fill_1 FILLER_79_351 ();
 sg13g2_fill_2 FILLER_79_356 ();
 sg13g2_fill_2 FILLER_79_470 ();
 sg13g2_fill_2 FILLER_79_519 ();
 sg13g2_fill_1 FILLER_79_521 ();
 sg13g2_fill_1 FILLER_79_549 ();
 sg13g2_fill_2 FILLER_79_565 ();
 sg13g2_fill_1 FILLER_79_567 ();
 sg13g2_fill_1 FILLER_79_621 ();
 sg13g2_decap_8 FILLER_79_649 ();
 sg13g2_decap_8 FILLER_79_656 ();
 sg13g2_decap_8 FILLER_79_663 ();
 sg13g2_decap_8 FILLER_79_670 ();
 sg13g2_decap_8 FILLER_79_677 ();
 sg13g2_decap_8 FILLER_79_684 ();
 sg13g2_decap_8 FILLER_79_691 ();
 sg13g2_decap_8 FILLER_79_698 ();
 sg13g2_decap_8 FILLER_79_705 ();
 sg13g2_decap_8 FILLER_79_712 ();
 sg13g2_decap_8 FILLER_79_719 ();
 sg13g2_decap_8 FILLER_79_726 ();
 sg13g2_decap_8 FILLER_79_733 ();
 sg13g2_decap_8 FILLER_79_740 ();
 sg13g2_decap_8 FILLER_79_747 ();
 sg13g2_decap_8 FILLER_79_754 ();
 sg13g2_decap_8 FILLER_79_761 ();
 sg13g2_decap_8 FILLER_79_768 ();
 sg13g2_decap_8 FILLER_79_775 ();
 sg13g2_decap_8 FILLER_79_782 ();
 sg13g2_decap_8 FILLER_79_789 ();
 sg13g2_decap_8 FILLER_79_796 ();
 sg13g2_decap_8 FILLER_79_803 ();
 sg13g2_decap_8 FILLER_79_810 ();
 sg13g2_decap_8 FILLER_79_817 ();
 sg13g2_decap_8 FILLER_79_824 ();
 sg13g2_decap_8 FILLER_79_831 ();
 sg13g2_decap_8 FILLER_79_838 ();
 sg13g2_decap_8 FILLER_79_845 ();
 sg13g2_decap_8 FILLER_79_852 ();
 sg13g2_fill_2 FILLER_79_859 ();
 sg13g2_fill_1 FILLER_79_861 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_fill_2 FILLER_80_108 ();
 sg13g2_fill_1 FILLER_80_110 ();
 sg13g2_fill_1 FILLER_80_180 ();
 sg13g2_fill_2 FILLER_80_189 ();
 sg13g2_decap_4 FILLER_80_233 ();
 sg13g2_fill_1 FILLER_80_237 ();
 sg13g2_fill_1 FILLER_80_270 ();
 sg13g2_fill_2 FILLER_80_275 ();
 sg13g2_fill_1 FILLER_80_277 ();
 sg13g2_fill_2 FILLER_80_314 ();
 sg13g2_fill_2 FILLER_80_429 ();
 sg13g2_fill_1 FILLER_80_431 ();
 sg13g2_fill_2 FILLER_80_437 ();
 sg13g2_fill_1 FILLER_80_467 ();
 sg13g2_fill_2 FILLER_80_477 ();
 sg13g2_fill_1 FILLER_80_479 ();
 sg13g2_fill_2 FILLER_80_516 ();
 sg13g2_fill_1 FILLER_80_594 ();
 sg13g2_fill_1 FILLER_80_604 ();
 sg13g2_fill_1 FILLER_80_614 ();
 sg13g2_fill_2 FILLER_80_633 ();
 sg13g2_decap_8 FILLER_80_656 ();
 sg13g2_decap_8 FILLER_80_663 ();
 sg13g2_decap_8 FILLER_80_670 ();
 sg13g2_decap_8 FILLER_80_677 ();
 sg13g2_decap_8 FILLER_80_684 ();
 sg13g2_decap_8 FILLER_80_691 ();
 sg13g2_decap_8 FILLER_80_698 ();
 sg13g2_decap_8 FILLER_80_705 ();
 sg13g2_decap_8 FILLER_80_712 ();
 sg13g2_decap_8 FILLER_80_719 ();
 sg13g2_decap_8 FILLER_80_726 ();
 sg13g2_decap_8 FILLER_80_733 ();
 sg13g2_decap_8 FILLER_80_740 ();
 sg13g2_decap_8 FILLER_80_747 ();
 sg13g2_decap_8 FILLER_80_754 ();
 sg13g2_decap_8 FILLER_80_761 ();
 sg13g2_decap_8 FILLER_80_768 ();
 sg13g2_decap_8 FILLER_80_775 ();
 sg13g2_decap_8 FILLER_80_782 ();
 sg13g2_decap_8 FILLER_80_789 ();
 sg13g2_decap_8 FILLER_80_796 ();
 sg13g2_decap_8 FILLER_80_803 ();
 sg13g2_decap_8 FILLER_80_810 ();
 sg13g2_decap_8 FILLER_80_817 ();
 sg13g2_decap_8 FILLER_80_824 ();
 sg13g2_decap_8 FILLER_80_831 ();
 sg13g2_decap_8 FILLER_80_838 ();
 sg13g2_decap_8 FILLER_80_845 ();
 sg13g2_decap_8 FILLER_80_852 ();
 sg13g2_fill_2 FILLER_80_859 ();
 sg13g2_fill_1 FILLER_80_861 ();
 assign uio_oe[0] = net5;
 assign uio_oe[1] = net6;
 assign uio_oe[2] = net7;
 assign uio_oe[3] = net8;
 assign uio_oe[4] = net9;
 assign uio_oe[5] = net10;
 assign uio_oe[6] = net11;
 assign uio_oe[7] = net12;
 assign uio_out[0] = net13;
 assign uio_out[1] = net14;
 assign uio_out[2] = net15;
 assign uio_out[3] = net16;
 assign uio_out[4] = net17;
 assign uio_out[5] = net18;
 assign uio_out[6] = net19;
 assign uio_out[7] = net20;
endmodule
