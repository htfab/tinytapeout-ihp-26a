module tt_um_ezrawolf_tinydcim_ihp26a (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire clknet_0_clk;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net4;
 wire net5;
 wire net6;
 wire net1;
 wire net2;
 wire net3;
 wire net7;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;

 sg13g2_inv_2 _053_ (.Y(_008_),
    .A(net4));
 sg13g2_o21ai_1 _054_ (.B1(net1),
    .Y(_009_),
    .A1(net2),
    .A2(net31));
 sg13g2_a21oi_1 _055_ (.A1(net6),
    .A2(net31),
    .Y(_000_),
    .B1(_009_));
 sg13g2_nor2b_1 _056_ (.A(net3),
    .B_N(net39),
    .Y(_010_));
 sg13g2_xnor2_1 _057_ (.Y(_011_),
    .A(net39),
    .B(net3));
 sg13g2_xnor2_1 _058_ (.Y(_012_),
    .A(net31),
    .B(_011_));
 sg13g2_o21ai_1 _059_ (.B1(net1),
    .Y(_013_),
    .A1(net6),
    .A2(net39));
 sg13g2_a21oi_1 _060_ (.A1(net6),
    .A2(_012_),
    .Y(_001_),
    .B1(_013_));
 sg13g2_a21oi_2 _061_ (.B1(_010_),
    .Y(_014_),
    .A2(_011_),
    .A1(net31));
 sg13g2_xnor2_1 _062_ (.Y(_015_),
    .A(net42),
    .B(net4));
 sg13g2_nor2b_1 _063_ (.A(_014_),
    .B_N(_015_),
    .Y(_016_));
 sg13g2_xor2_1 _064_ (.B(_015_),
    .A(_014_),
    .X(_017_));
 sg13g2_o21ai_1 _065_ (.B1(net1),
    .Y(_018_),
    .A1(net6),
    .A2(net42));
 sg13g2_a21oi_1 _066_ (.A1(net6),
    .A2(_017_),
    .Y(_002_),
    .B1(_018_));
 sg13g2_xnor2_1 _067_ (.Y(_019_),
    .A(net34),
    .B(net4));
 sg13g2_a21o_1 _068_ (.A2(_008_),
    .A1(uo_out[2]),
    .B1(_016_),
    .X(_020_));
 sg13g2_xnor2_1 _069_ (.Y(_021_),
    .A(_019_),
    .B(_020_));
 sg13g2_o21ai_1 _070_ (.B1(net1),
    .Y(_022_),
    .A1(net6),
    .A2(net34));
 sg13g2_a21oi_1 _071_ (.A1(net6),
    .A2(_021_),
    .Y(_003_),
    .B1(_022_));
 sg13g2_nand2_1 _072_ (.Y(_023_),
    .A(_015_),
    .B(_019_));
 sg13g2_o21ai_1 _073_ (.B1(_008_),
    .Y(_024_),
    .A1(uo_out[3]),
    .A2(uo_out[2]));
 sg13g2_o21ai_1 _074_ (.B1(_024_),
    .Y(_025_),
    .A1(_014_),
    .A2(_023_));
 sg13g2_nor2b_1 _075_ (.A(net4),
    .B_N(uo_out[4]),
    .Y(_026_));
 sg13g2_xnor2_1 _076_ (.Y(_027_),
    .A(net40),
    .B(net4));
 sg13g2_inv_1 _077_ (.Y(_028_),
    .A(_027_));
 sg13g2_xnor2_1 _078_ (.Y(_029_),
    .A(_025_),
    .B(_027_));
 sg13g2_o21ai_1 _079_ (.B1(net1),
    .Y(_030_),
    .A1(net5),
    .A2(net40));
 sg13g2_a21oi_1 _080_ (.A1(net5),
    .A2(_029_),
    .Y(_004_),
    .B1(_030_));
 sg13g2_xor2_1 _081_ (.B(net4),
    .A(net37),
    .X(_031_));
 sg13g2_a21oi_1 _082_ (.A1(_025_),
    .A2(_027_),
    .Y(_032_),
    .B1(_026_));
 sg13g2_xnor2_1 _083_ (.Y(_033_),
    .A(_031_),
    .B(_032_));
 sg13g2_o21ai_1 _084_ (.B1(net1),
    .Y(_034_),
    .A1(net5),
    .A2(net37));
 sg13g2_a21oi_1 _085_ (.A1(net5),
    .A2(_033_),
    .Y(_005_),
    .B1(_034_));
 sg13g2_nand2_1 _086_ (.Y(_035_),
    .A(net32),
    .B(_008_));
 sg13g2_xor2_1 _087_ (.B(net4),
    .A(net32),
    .X(_036_));
 sg13g2_nor2_1 _088_ (.A(_028_),
    .B(_031_),
    .Y(_037_));
 sg13g2_a221oi_1 _089_ (.B2(_037_),
    .C1(_026_),
    .B1(_025_),
    .A1(uo_out[5]),
    .Y(_038_),
    .A2(_008_));
 sg13g2_xnor2_1 _090_ (.Y(_039_),
    .A(_036_),
    .B(_038_));
 sg13g2_o21ai_1 _091_ (.B1(net1),
    .Y(_040_),
    .A1(net5),
    .A2(net32));
 sg13g2_a21oi_1 _092_ (.A1(net5),
    .A2(_039_),
    .Y(_006_),
    .B1(_040_));
 sg13g2_o21ai_1 _093_ (.B1(_035_),
    .Y(_041_),
    .A1(_036_),
    .A2(_038_));
 sg13g2_xnor2_1 _094_ (.Y(_042_),
    .A(net36),
    .B(net4));
 sg13g2_xnor2_1 _095_ (.Y(_043_),
    .A(_041_),
    .B(_042_));
 sg13g2_o21ai_1 _096_ (.B1(net1),
    .Y(_044_),
    .A1(net36),
    .A2(net5));
 sg13g2_a21oi_1 _097_ (.A1(net5),
    .A2(_043_),
    .Y(_007_),
    .B1(_044_));
 sg13g2_dfrbpq_2 _098_ (.RESET_B(net23),
    .D(_000_),
    .Q(uo_out[0]),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_2 _099_ (.RESET_B(net30),
    .D(_001_),
    .Q(uo_out[1]),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_2 _100_ (.RESET_B(net28),
    .D(_002_),
    .Q(uo_out[2]),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_2 _101_ (.RESET_B(net26),
    .D(net35),
    .Q(uo_out[3]),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_2 _102_ (.RESET_B(net24),
    .D(net41),
    .Q(uo_out[4]),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_2 _103_ (.RESET_B(net29),
    .D(net38),
    .Q(uo_out[5]),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_2 _104_ (.RESET_B(net25),
    .D(net33),
    .Q(uo_out[6]),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_2 _105_ (.RESET_B(net27),
    .D(_007_),
    .Q(uo_out[7]),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_tiehi _102__21 (.L_HI(net24));
 sg13g2_tiehi _104__22 (.L_HI(net25));
 sg13g2_tiehi _101__23 (.L_HI(net26));
 sg13g2_tiehi _105__24 (.L_HI(net27));
 sg13g2_tiehi _100__25 (.L_HI(net28));
 sg13g2_tiehi _103__26 (.L_HI(net29));
 sg13g2_tiehi _099__27 (.L_HI(net30));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_ezrawolf_tinydcim_ihp26a_5 (.L_LO(net8));
 sg13g2_tielo tt_um_ezrawolf_tinydcim_ihp26a_6 (.L_LO(net9));
 sg13g2_tielo tt_um_ezrawolf_tinydcim_ihp26a_7 (.L_LO(net10));
 sg13g2_tielo tt_um_ezrawolf_tinydcim_ihp26a_8 (.L_LO(net11));
 sg13g2_tielo tt_um_ezrawolf_tinydcim_ihp26a_9 (.L_LO(net12));
 sg13g2_tielo tt_um_ezrawolf_tinydcim_ihp26a_10 (.L_LO(net13));
 sg13g2_tielo tt_um_ezrawolf_tinydcim_ihp26a_11 (.L_LO(net14));
 sg13g2_tielo tt_um_ezrawolf_tinydcim_ihp26a_12 (.L_LO(net15));
 sg13g2_tielo tt_um_ezrawolf_tinydcim_ihp26a_13 (.L_LO(net16));
 sg13g2_tielo tt_um_ezrawolf_tinydcim_ihp26a_14 (.L_LO(net17));
 sg13g2_tielo tt_um_ezrawolf_tinydcim_ihp26a_15 (.L_LO(net18));
 sg13g2_tielo tt_um_ezrawolf_tinydcim_ihp26a_16 (.L_LO(net19));
 sg13g2_tielo tt_um_ezrawolf_tinydcim_ihp26a_17 (.L_LO(net20));
 sg13g2_tielo tt_um_ezrawolf_tinydcim_ihp26a_18 (.L_LO(net21));
 sg13g2_tielo tt_um_ezrawolf_tinydcim_ihp26a_19 (.L_LO(net22));
 sg13g2_tiehi _098__20 (.L_HI(net23));
 sg13g2_buf_8 fanout4 (.A(net3),
    .X(net4));
 sg13g2_buf_8 fanout5 (.A(net6),
    .X(net5));
 sg13g2_buf_8 fanout6 (.A(net2),
    .X(net6));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_tielo tt_um_ezrawolf_tinydcim_ihp26a_4 (.L_LO(net7));
 sg13g2_buf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(uo_out[0]),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold2 (.A(uo_out[6]),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold3 (.A(_006_),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold4 (.A(uo_out[3]),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold5 (.A(_003_),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold6 (.A(uo_out[7]),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold7 (.A(uo_out[5]),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold8 (.A(_005_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold9 (.A(uo_out[1]),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold10 (.A(uo_out[4]),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold11 (.A(_004_),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold12 (.A(uo_out[2]),
    .X(net42));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_decap_8 FILLER_0_875 ();
 sg13g2_decap_8 FILLER_0_882 ();
 sg13g2_decap_8 FILLER_0_889 ();
 sg13g2_decap_8 FILLER_0_896 ();
 sg13g2_decap_8 FILLER_0_903 ();
 sg13g2_decap_8 FILLER_0_910 ();
 sg13g2_decap_8 FILLER_0_917 ();
 sg13g2_decap_8 FILLER_0_924 ();
 sg13g2_decap_8 FILLER_0_931 ();
 sg13g2_decap_8 FILLER_0_938 ();
 sg13g2_decap_8 FILLER_0_945 ();
 sg13g2_decap_8 FILLER_0_952 ();
 sg13g2_decap_8 FILLER_0_959 ();
 sg13g2_decap_8 FILLER_0_966 ();
 sg13g2_decap_8 FILLER_0_973 ();
 sg13g2_decap_8 FILLER_0_980 ();
 sg13g2_decap_8 FILLER_0_987 ();
 sg13g2_decap_8 FILLER_0_994 ();
 sg13g2_decap_8 FILLER_0_1001 ();
 sg13g2_decap_8 FILLER_0_1008 ();
 sg13g2_decap_8 FILLER_0_1015 ();
 sg13g2_decap_8 FILLER_0_1022 ();
 sg13g2_decap_8 FILLER_0_1029 ();
 sg13g2_decap_8 FILLER_0_1036 ();
 sg13g2_decap_8 FILLER_0_1043 ();
 sg13g2_decap_8 FILLER_0_1050 ();
 sg13g2_decap_8 FILLER_0_1057 ();
 sg13g2_decap_8 FILLER_0_1064 ();
 sg13g2_decap_8 FILLER_0_1071 ();
 sg13g2_decap_8 FILLER_0_1078 ();
 sg13g2_decap_8 FILLER_0_1085 ();
 sg13g2_decap_8 FILLER_0_1092 ();
 sg13g2_decap_8 FILLER_0_1099 ();
 sg13g2_decap_8 FILLER_0_1106 ();
 sg13g2_decap_8 FILLER_0_1113 ();
 sg13g2_decap_8 FILLER_0_1120 ();
 sg13g2_decap_8 FILLER_0_1127 ();
 sg13g2_decap_8 FILLER_0_1134 ();
 sg13g2_decap_8 FILLER_0_1141 ();
 sg13g2_decap_8 FILLER_0_1148 ();
 sg13g2_decap_8 FILLER_0_1155 ();
 sg13g2_decap_8 FILLER_0_1162 ();
 sg13g2_decap_8 FILLER_0_1169 ();
 sg13g2_decap_8 FILLER_0_1176 ();
 sg13g2_decap_8 FILLER_0_1183 ();
 sg13g2_decap_8 FILLER_0_1190 ();
 sg13g2_decap_8 FILLER_0_1197 ();
 sg13g2_decap_8 FILLER_0_1204 ();
 sg13g2_decap_8 FILLER_0_1211 ();
 sg13g2_decap_8 FILLER_0_1218 ();
 sg13g2_decap_8 FILLER_0_1225 ();
 sg13g2_decap_8 FILLER_0_1232 ();
 sg13g2_decap_8 FILLER_0_1239 ();
 sg13g2_decap_8 FILLER_0_1246 ();
 sg13g2_decap_8 FILLER_0_1253 ();
 sg13g2_decap_8 FILLER_0_1260 ();
 sg13g2_decap_8 FILLER_0_1267 ();
 sg13g2_decap_8 FILLER_0_1274 ();
 sg13g2_decap_8 FILLER_0_1281 ();
 sg13g2_decap_8 FILLER_0_1288 ();
 sg13g2_decap_8 FILLER_0_1295 ();
 sg13g2_decap_8 FILLER_0_1302 ();
 sg13g2_decap_8 FILLER_0_1309 ();
 sg13g2_decap_8 FILLER_0_1316 ();
 sg13g2_decap_8 FILLER_0_1323 ();
 sg13g2_decap_8 FILLER_0_1330 ();
 sg13g2_decap_8 FILLER_0_1337 ();
 sg13g2_decap_8 FILLER_0_1344 ();
 sg13g2_decap_8 FILLER_0_1351 ();
 sg13g2_decap_8 FILLER_0_1358 ();
 sg13g2_decap_8 FILLER_0_1365 ();
 sg13g2_decap_8 FILLER_0_1372 ();
 sg13g2_decap_8 FILLER_0_1379 ();
 sg13g2_decap_8 FILLER_0_1386 ();
 sg13g2_decap_8 FILLER_0_1393 ();
 sg13g2_decap_8 FILLER_0_1400 ();
 sg13g2_decap_8 FILLER_0_1407 ();
 sg13g2_decap_8 FILLER_0_1414 ();
 sg13g2_decap_8 FILLER_0_1421 ();
 sg13g2_decap_8 FILLER_0_1428 ();
 sg13g2_decap_8 FILLER_0_1435 ();
 sg13g2_decap_8 FILLER_0_1442 ();
 sg13g2_decap_8 FILLER_0_1449 ();
 sg13g2_decap_8 FILLER_0_1456 ();
 sg13g2_decap_8 FILLER_0_1463 ();
 sg13g2_decap_8 FILLER_0_1470 ();
 sg13g2_decap_8 FILLER_0_1477 ();
 sg13g2_decap_8 FILLER_0_1484 ();
 sg13g2_decap_8 FILLER_0_1491 ();
 sg13g2_decap_8 FILLER_0_1498 ();
 sg13g2_decap_8 FILLER_0_1505 ();
 sg13g2_decap_8 FILLER_0_1512 ();
 sg13g2_decap_8 FILLER_0_1519 ();
 sg13g2_decap_8 FILLER_0_1526 ();
 sg13g2_decap_8 FILLER_0_1533 ();
 sg13g2_decap_8 FILLER_0_1540 ();
 sg13g2_decap_8 FILLER_0_1547 ();
 sg13g2_decap_8 FILLER_0_1554 ();
 sg13g2_decap_8 FILLER_0_1561 ();
 sg13g2_decap_8 FILLER_0_1568 ();
 sg13g2_decap_8 FILLER_0_1575 ();
 sg13g2_decap_8 FILLER_0_1582 ();
 sg13g2_decap_8 FILLER_0_1589 ();
 sg13g2_decap_8 FILLER_0_1596 ();
 sg13g2_decap_8 FILLER_0_1603 ();
 sg13g2_decap_8 FILLER_0_1610 ();
 sg13g2_decap_8 FILLER_0_1617 ();
 sg13g2_decap_8 FILLER_0_1624 ();
 sg13g2_decap_8 FILLER_0_1631 ();
 sg13g2_decap_8 FILLER_0_1638 ();
 sg13g2_decap_8 FILLER_0_1645 ();
 sg13g2_decap_8 FILLER_0_1652 ();
 sg13g2_decap_8 FILLER_0_1659 ();
 sg13g2_decap_8 FILLER_0_1666 ();
 sg13g2_decap_8 FILLER_0_1673 ();
 sg13g2_decap_8 FILLER_0_1680 ();
 sg13g2_decap_8 FILLER_0_1687 ();
 sg13g2_decap_8 FILLER_0_1694 ();
 sg13g2_decap_8 FILLER_0_1701 ();
 sg13g2_decap_8 FILLER_0_1708 ();
 sg13g2_decap_8 FILLER_0_1715 ();
 sg13g2_decap_8 FILLER_0_1722 ();
 sg13g2_decap_8 FILLER_0_1729 ();
 sg13g2_decap_8 FILLER_0_1736 ();
 sg13g2_decap_8 FILLER_0_1743 ();
 sg13g2_decap_8 FILLER_0_1750 ();
 sg13g2_decap_8 FILLER_0_1757 ();
 sg13g2_decap_8 FILLER_0_1764 ();
 sg13g2_decap_8 FILLER_0_1771 ();
 sg13g2_decap_8 FILLER_0_1778 ();
 sg13g2_decap_8 FILLER_0_1785 ();
 sg13g2_decap_8 FILLER_0_1792 ();
 sg13g2_decap_8 FILLER_0_1799 ();
 sg13g2_decap_8 FILLER_0_1806 ();
 sg13g2_decap_8 FILLER_0_1813 ();
 sg13g2_decap_8 FILLER_0_1820 ();
 sg13g2_decap_8 FILLER_0_1827 ();
 sg13g2_decap_8 FILLER_0_1834 ();
 sg13g2_decap_8 FILLER_0_1841 ();
 sg13g2_decap_8 FILLER_0_1848 ();
 sg13g2_decap_8 FILLER_0_1855 ();
 sg13g2_decap_8 FILLER_0_1862 ();
 sg13g2_decap_8 FILLER_0_1869 ();
 sg13g2_decap_8 FILLER_0_1876 ();
 sg13g2_decap_8 FILLER_0_1883 ();
 sg13g2_decap_8 FILLER_0_1890 ();
 sg13g2_decap_8 FILLER_0_1897 ();
 sg13g2_decap_8 FILLER_0_1904 ();
 sg13g2_decap_8 FILLER_0_1911 ();
 sg13g2_decap_8 FILLER_0_1918 ();
 sg13g2_decap_8 FILLER_0_1925 ();
 sg13g2_decap_8 FILLER_0_1932 ();
 sg13g2_decap_8 FILLER_0_1939 ();
 sg13g2_decap_8 FILLER_0_1946 ();
 sg13g2_decap_8 FILLER_0_1953 ();
 sg13g2_decap_8 FILLER_0_1960 ();
 sg13g2_decap_8 FILLER_0_1967 ();
 sg13g2_decap_8 FILLER_0_1974 ();
 sg13g2_decap_8 FILLER_0_1981 ();
 sg13g2_decap_8 FILLER_0_1988 ();
 sg13g2_decap_8 FILLER_0_1995 ();
 sg13g2_decap_8 FILLER_0_2002 ();
 sg13g2_decap_8 FILLER_0_2009 ();
 sg13g2_decap_8 FILLER_0_2016 ();
 sg13g2_decap_8 FILLER_0_2023 ();
 sg13g2_decap_8 FILLER_0_2030 ();
 sg13g2_decap_8 FILLER_0_2037 ();
 sg13g2_decap_8 FILLER_0_2044 ();
 sg13g2_decap_8 FILLER_0_2051 ();
 sg13g2_decap_8 FILLER_0_2058 ();
 sg13g2_decap_8 FILLER_0_2065 ();
 sg13g2_decap_8 FILLER_0_2072 ();
 sg13g2_decap_8 FILLER_0_2079 ();
 sg13g2_decap_8 FILLER_0_2086 ();
 sg13g2_decap_8 FILLER_0_2093 ();
 sg13g2_decap_8 FILLER_0_2100 ();
 sg13g2_decap_8 FILLER_0_2107 ();
 sg13g2_decap_8 FILLER_0_2114 ();
 sg13g2_decap_8 FILLER_0_2121 ();
 sg13g2_decap_8 FILLER_0_2128 ();
 sg13g2_decap_8 FILLER_0_2135 ();
 sg13g2_decap_8 FILLER_0_2142 ();
 sg13g2_decap_8 FILLER_0_2149 ();
 sg13g2_decap_8 FILLER_0_2156 ();
 sg13g2_decap_8 FILLER_0_2163 ();
 sg13g2_decap_8 FILLER_0_2170 ();
 sg13g2_decap_8 FILLER_0_2177 ();
 sg13g2_decap_8 FILLER_0_2184 ();
 sg13g2_decap_8 FILLER_0_2191 ();
 sg13g2_decap_8 FILLER_0_2198 ();
 sg13g2_decap_8 FILLER_0_2205 ();
 sg13g2_decap_8 FILLER_0_2212 ();
 sg13g2_decap_8 FILLER_0_2219 ();
 sg13g2_decap_8 FILLER_0_2226 ();
 sg13g2_decap_8 FILLER_0_2233 ();
 sg13g2_decap_8 FILLER_0_2240 ();
 sg13g2_decap_8 FILLER_0_2247 ();
 sg13g2_decap_8 FILLER_0_2254 ();
 sg13g2_decap_8 FILLER_0_2261 ();
 sg13g2_decap_8 FILLER_0_2268 ();
 sg13g2_decap_8 FILLER_0_2275 ();
 sg13g2_decap_8 FILLER_0_2282 ();
 sg13g2_decap_8 FILLER_0_2289 ();
 sg13g2_decap_8 FILLER_0_2296 ();
 sg13g2_decap_8 FILLER_0_2303 ();
 sg13g2_decap_8 FILLER_0_2310 ();
 sg13g2_decap_8 FILLER_0_2317 ();
 sg13g2_decap_8 FILLER_0_2324 ();
 sg13g2_decap_8 FILLER_0_2331 ();
 sg13g2_decap_8 FILLER_0_2338 ();
 sg13g2_decap_8 FILLER_0_2345 ();
 sg13g2_decap_8 FILLER_0_2352 ();
 sg13g2_decap_8 FILLER_0_2359 ();
 sg13g2_decap_8 FILLER_0_2366 ();
 sg13g2_decap_8 FILLER_0_2373 ();
 sg13g2_decap_8 FILLER_0_2380 ();
 sg13g2_decap_8 FILLER_0_2387 ();
 sg13g2_decap_8 FILLER_0_2394 ();
 sg13g2_decap_8 FILLER_0_2401 ();
 sg13g2_decap_8 FILLER_0_2408 ();
 sg13g2_decap_8 FILLER_0_2415 ();
 sg13g2_decap_8 FILLER_0_2422 ();
 sg13g2_decap_8 FILLER_0_2429 ();
 sg13g2_decap_8 FILLER_0_2436 ();
 sg13g2_decap_8 FILLER_0_2443 ();
 sg13g2_decap_8 FILLER_0_2450 ();
 sg13g2_decap_8 FILLER_0_2457 ();
 sg13g2_decap_8 FILLER_0_2464 ();
 sg13g2_decap_8 FILLER_0_2471 ();
 sg13g2_decap_8 FILLER_0_2478 ();
 sg13g2_decap_8 FILLER_0_2485 ();
 sg13g2_decap_8 FILLER_0_2492 ();
 sg13g2_decap_8 FILLER_0_2499 ();
 sg13g2_decap_8 FILLER_0_2506 ();
 sg13g2_decap_8 FILLER_0_2513 ();
 sg13g2_decap_8 FILLER_0_2520 ();
 sg13g2_decap_8 FILLER_0_2527 ();
 sg13g2_decap_8 FILLER_0_2534 ();
 sg13g2_decap_8 FILLER_0_2541 ();
 sg13g2_decap_8 FILLER_0_2548 ();
 sg13g2_decap_8 FILLER_0_2555 ();
 sg13g2_decap_8 FILLER_0_2562 ();
 sg13g2_decap_8 FILLER_0_2569 ();
 sg13g2_decap_8 FILLER_0_2576 ();
 sg13g2_decap_8 FILLER_0_2583 ();
 sg13g2_decap_8 FILLER_0_2590 ();
 sg13g2_decap_8 FILLER_0_2597 ();
 sg13g2_decap_8 FILLER_0_2604 ();
 sg13g2_decap_8 FILLER_0_2611 ();
 sg13g2_decap_8 FILLER_0_2618 ();
 sg13g2_decap_8 FILLER_0_2625 ();
 sg13g2_decap_8 FILLER_0_2632 ();
 sg13g2_decap_8 FILLER_0_2639 ();
 sg13g2_decap_8 FILLER_0_2646 ();
 sg13g2_decap_8 FILLER_0_2653 ();
 sg13g2_decap_8 FILLER_0_2660 ();
 sg13g2_decap_8 FILLER_0_2667 ();
 sg13g2_decap_8 FILLER_0_2674 ();
 sg13g2_decap_8 FILLER_0_2681 ();
 sg13g2_decap_8 FILLER_0_2688 ();
 sg13g2_decap_8 FILLER_0_2695 ();
 sg13g2_decap_8 FILLER_0_2702 ();
 sg13g2_decap_8 FILLER_0_2709 ();
 sg13g2_decap_8 FILLER_0_2716 ();
 sg13g2_decap_8 FILLER_0_2723 ();
 sg13g2_decap_8 FILLER_0_2730 ();
 sg13g2_decap_8 FILLER_0_2737 ();
 sg13g2_decap_8 FILLER_0_2744 ();
 sg13g2_decap_8 FILLER_0_2751 ();
 sg13g2_decap_8 FILLER_0_2758 ();
 sg13g2_decap_8 FILLER_0_2765 ();
 sg13g2_decap_8 FILLER_0_2772 ();
 sg13g2_decap_8 FILLER_0_2779 ();
 sg13g2_decap_8 FILLER_0_2786 ();
 sg13g2_decap_8 FILLER_0_2793 ();
 sg13g2_decap_8 FILLER_0_2800 ();
 sg13g2_decap_8 FILLER_0_2807 ();
 sg13g2_decap_8 FILLER_0_2814 ();
 sg13g2_decap_8 FILLER_0_2821 ();
 sg13g2_decap_8 FILLER_0_2828 ();
 sg13g2_decap_8 FILLER_0_2835 ();
 sg13g2_decap_8 FILLER_0_2842 ();
 sg13g2_decap_8 FILLER_0_2849 ();
 sg13g2_decap_8 FILLER_0_2856 ();
 sg13g2_decap_8 FILLER_0_2863 ();
 sg13g2_decap_8 FILLER_0_2870 ();
 sg13g2_decap_8 FILLER_0_2877 ();
 sg13g2_decap_8 FILLER_0_2884 ();
 sg13g2_decap_8 FILLER_0_2891 ();
 sg13g2_decap_8 FILLER_0_2898 ();
 sg13g2_decap_8 FILLER_0_2905 ();
 sg13g2_decap_8 FILLER_0_2912 ();
 sg13g2_decap_8 FILLER_0_2919 ();
 sg13g2_decap_8 FILLER_0_2926 ();
 sg13g2_decap_8 FILLER_0_2933 ();
 sg13g2_decap_8 FILLER_0_2940 ();
 sg13g2_decap_8 FILLER_0_2947 ();
 sg13g2_decap_8 FILLER_0_2954 ();
 sg13g2_decap_8 FILLER_0_2961 ();
 sg13g2_decap_8 FILLER_0_2968 ();
 sg13g2_decap_8 FILLER_0_2975 ();
 sg13g2_decap_8 FILLER_0_2982 ();
 sg13g2_decap_8 FILLER_0_2989 ();
 sg13g2_decap_8 FILLER_0_2996 ();
 sg13g2_decap_8 FILLER_0_3003 ();
 sg13g2_decap_8 FILLER_0_3010 ();
 sg13g2_decap_8 FILLER_0_3017 ();
 sg13g2_decap_8 FILLER_0_3024 ();
 sg13g2_decap_8 FILLER_0_3031 ();
 sg13g2_decap_8 FILLER_0_3038 ();
 sg13g2_decap_8 FILLER_0_3045 ();
 sg13g2_decap_8 FILLER_0_3052 ();
 sg13g2_decap_8 FILLER_0_3059 ();
 sg13g2_decap_8 FILLER_0_3066 ();
 sg13g2_decap_8 FILLER_0_3073 ();
 sg13g2_decap_8 FILLER_0_3080 ();
 sg13g2_decap_8 FILLER_0_3087 ();
 sg13g2_decap_8 FILLER_0_3094 ();
 sg13g2_decap_8 FILLER_0_3101 ();
 sg13g2_decap_8 FILLER_0_3108 ();
 sg13g2_decap_8 FILLER_0_3115 ();
 sg13g2_decap_8 FILLER_0_3122 ();
 sg13g2_decap_8 FILLER_0_3129 ();
 sg13g2_decap_8 FILLER_0_3136 ();
 sg13g2_decap_8 FILLER_0_3143 ();
 sg13g2_decap_8 FILLER_0_3150 ();
 sg13g2_decap_8 FILLER_0_3157 ();
 sg13g2_decap_8 FILLER_0_3164 ();
 sg13g2_decap_8 FILLER_0_3171 ();
 sg13g2_decap_8 FILLER_0_3178 ();
 sg13g2_decap_8 FILLER_0_3185 ();
 sg13g2_decap_8 FILLER_0_3192 ();
 sg13g2_decap_8 FILLER_0_3199 ();
 sg13g2_decap_8 FILLER_0_3206 ();
 sg13g2_decap_8 FILLER_0_3213 ();
 sg13g2_decap_8 FILLER_0_3220 ();
 sg13g2_decap_8 FILLER_0_3227 ();
 sg13g2_decap_8 FILLER_0_3234 ();
 sg13g2_decap_8 FILLER_0_3241 ();
 sg13g2_decap_8 FILLER_0_3248 ();
 sg13g2_decap_8 FILLER_0_3255 ();
 sg13g2_decap_8 FILLER_0_3262 ();
 sg13g2_decap_8 FILLER_0_3269 ();
 sg13g2_decap_8 FILLER_0_3276 ();
 sg13g2_decap_8 FILLER_0_3283 ();
 sg13g2_decap_8 FILLER_0_3290 ();
 sg13g2_decap_8 FILLER_0_3297 ();
 sg13g2_decap_8 FILLER_0_3304 ();
 sg13g2_decap_8 FILLER_0_3311 ();
 sg13g2_decap_8 FILLER_0_3318 ();
 sg13g2_decap_8 FILLER_0_3325 ();
 sg13g2_decap_8 FILLER_0_3332 ();
 sg13g2_decap_8 FILLER_0_3339 ();
 sg13g2_decap_8 FILLER_0_3346 ();
 sg13g2_decap_8 FILLER_0_3353 ();
 sg13g2_decap_8 FILLER_0_3360 ();
 sg13g2_decap_8 FILLER_0_3367 ();
 sg13g2_decap_8 FILLER_0_3374 ();
 sg13g2_decap_8 FILLER_0_3381 ();
 sg13g2_decap_8 FILLER_0_3388 ();
 sg13g2_decap_8 FILLER_0_3395 ();
 sg13g2_decap_8 FILLER_0_3402 ();
 sg13g2_decap_8 FILLER_0_3409 ();
 sg13g2_decap_8 FILLER_0_3416 ();
 sg13g2_decap_8 FILLER_0_3423 ();
 sg13g2_decap_8 FILLER_0_3430 ();
 sg13g2_decap_8 FILLER_0_3437 ();
 sg13g2_decap_8 FILLER_0_3444 ();
 sg13g2_decap_8 FILLER_0_3451 ();
 sg13g2_decap_8 FILLER_0_3458 ();
 sg13g2_decap_8 FILLER_0_3465 ();
 sg13g2_decap_8 FILLER_0_3472 ();
 sg13g2_decap_8 FILLER_0_3479 ();
 sg13g2_decap_8 FILLER_0_3486 ();
 sg13g2_decap_8 FILLER_0_3493 ();
 sg13g2_decap_8 FILLER_0_3500 ();
 sg13g2_decap_8 FILLER_0_3507 ();
 sg13g2_decap_8 FILLER_0_3514 ();
 sg13g2_decap_8 FILLER_0_3521 ();
 sg13g2_decap_8 FILLER_0_3528 ();
 sg13g2_decap_8 FILLER_0_3535 ();
 sg13g2_decap_8 FILLER_0_3542 ();
 sg13g2_decap_8 FILLER_0_3549 ();
 sg13g2_decap_8 FILLER_0_3556 ();
 sg13g2_decap_8 FILLER_0_3563 ();
 sg13g2_decap_8 FILLER_0_3570 ();
 sg13g2_fill_2 FILLER_0_3577 ();
 sg13g2_fill_1 FILLER_0_3579 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_decap_8 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_1_868 ();
 sg13g2_decap_8 FILLER_1_875 ();
 sg13g2_decap_8 FILLER_1_882 ();
 sg13g2_decap_8 FILLER_1_889 ();
 sg13g2_decap_8 FILLER_1_896 ();
 sg13g2_decap_8 FILLER_1_903 ();
 sg13g2_decap_8 FILLER_1_910 ();
 sg13g2_decap_8 FILLER_1_917 ();
 sg13g2_decap_8 FILLER_1_924 ();
 sg13g2_decap_8 FILLER_1_931 ();
 sg13g2_decap_8 FILLER_1_938 ();
 sg13g2_decap_8 FILLER_1_945 ();
 sg13g2_decap_8 FILLER_1_952 ();
 sg13g2_decap_8 FILLER_1_959 ();
 sg13g2_decap_8 FILLER_1_966 ();
 sg13g2_decap_8 FILLER_1_973 ();
 sg13g2_decap_8 FILLER_1_980 ();
 sg13g2_decap_8 FILLER_1_987 ();
 sg13g2_decap_8 FILLER_1_994 ();
 sg13g2_decap_8 FILLER_1_1001 ();
 sg13g2_decap_8 FILLER_1_1008 ();
 sg13g2_decap_8 FILLER_1_1015 ();
 sg13g2_decap_8 FILLER_1_1022 ();
 sg13g2_decap_8 FILLER_1_1029 ();
 sg13g2_decap_8 FILLER_1_1036 ();
 sg13g2_decap_8 FILLER_1_1043 ();
 sg13g2_decap_8 FILLER_1_1050 ();
 sg13g2_decap_8 FILLER_1_1057 ();
 sg13g2_decap_8 FILLER_1_1064 ();
 sg13g2_decap_8 FILLER_1_1071 ();
 sg13g2_decap_8 FILLER_1_1078 ();
 sg13g2_decap_8 FILLER_1_1085 ();
 sg13g2_decap_8 FILLER_1_1092 ();
 sg13g2_decap_8 FILLER_1_1099 ();
 sg13g2_decap_8 FILLER_1_1106 ();
 sg13g2_decap_8 FILLER_1_1113 ();
 sg13g2_decap_8 FILLER_1_1120 ();
 sg13g2_decap_8 FILLER_1_1127 ();
 sg13g2_decap_8 FILLER_1_1134 ();
 sg13g2_decap_8 FILLER_1_1141 ();
 sg13g2_decap_8 FILLER_1_1148 ();
 sg13g2_decap_8 FILLER_1_1155 ();
 sg13g2_decap_8 FILLER_1_1162 ();
 sg13g2_decap_8 FILLER_1_1169 ();
 sg13g2_decap_8 FILLER_1_1176 ();
 sg13g2_decap_8 FILLER_1_1183 ();
 sg13g2_decap_8 FILLER_1_1190 ();
 sg13g2_decap_8 FILLER_1_1197 ();
 sg13g2_decap_8 FILLER_1_1204 ();
 sg13g2_decap_8 FILLER_1_1211 ();
 sg13g2_decap_8 FILLER_1_1218 ();
 sg13g2_decap_8 FILLER_1_1225 ();
 sg13g2_decap_8 FILLER_1_1232 ();
 sg13g2_decap_8 FILLER_1_1239 ();
 sg13g2_decap_8 FILLER_1_1246 ();
 sg13g2_decap_8 FILLER_1_1253 ();
 sg13g2_decap_8 FILLER_1_1260 ();
 sg13g2_decap_8 FILLER_1_1267 ();
 sg13g2_decap_8 FILLER_1_1274 ();
 sg13g2_decap_8 FILLER_1_1281 ();
 sg13g2_decap_8 FILLER_1_1288 ();
 sg13g2_decap_8 FILLER_1_1295 ();
 sg13g2_decap_8 FILLER_1_1302 ();
 sg13g2_decap_8 FILLER_1_1309 ();
 sg13g2_decap_8 FILLER_1_1316 ();
 sg13g2_decap_8 FILLER_1_1323 ();
 sg13g2_decap_8 FILLER_1_1330 ();
 sg13g2_decap_8 FILLER_1_1337 ();
 sg13g2_decap_8 FILLER_1_1344 ();
 sg13g2_decap_8 FILLER_1_1351 ();
 sg13g2_decap_8 FILLER_1_1358 ();
 sg13g2_decap_8 FILLER_1_1365 ();
 sg13g2_decap_8 FILLER_1_1372 ();
 sg13g2_decap_8 FILLER_1_1379 ();
 sg13g2_decap_8 FILLER_1_1386 ();
 sg13g2_decap_8 FILLER_1_1393 ();
 sg13g2_decap_8 FILLER_1_1400 ();
 sg13g2_decap_8 FILLER_1_1407 ();
 sg13g2_decap_8 FILLER_1_1414 ();
 sg13g2_decap_8 FILLER_1_1421 ();
 sg13g2_decap_8 FILLER_1_1428 ();
 sg13g2_decap_8 FILLER_1_1435 ();
 sg13g2_decap_8 FILLER_1_1442 ();
 sg13g2_decap_8 FILLER_1_1449 ();
 sg13g2_decap_8 FILLER_1_1456 ();
 sg13g2_decap_8 FILLER_1_1463 ();
 sg13g2_decap_8 FILLER_1_1470 ();
 sg13g2_decap_8 FILLER_1_1477 ();
 sg13g2_decap_8 FILLER_1_1484 ();
 sg13g2_decap_8 FILLER_1_1491 ();
 sg13g2_decap_8 FILLER_1_1498 ();
 sg13g2_decap_8 FILLER_1_1505 ();
 sg13g2_decap_8 FILLER_1_1512 ();
 sg13g2_decap_8 FILLER_1_1519 ();
 sg13g2_decap_8 FILLER_1_1526 ();
 sg13g2_decap_8 FILLER_1_1533 ();
 sg13g2_decap_8 FILLER_1_1540 ();
 sg13g2_decap_8 FILLER_1_1547 ();
 sg13g2_decap_8 FILLER_1_1554 ();
 sg13g2_decap_8 FILLER_1_1561 ();
 sg13g2_decap_8 FILLER_1_1568 ();
 sg13g2_decap_8 FILLER_1_1575 ();
 sg13g2_decap_8 FILLER_1_1582 ();
 sg13g2_decap_8 FILLER_1_1589 ();
 sg13g2_decap_8 FILLER_1_1596 ();
 sg13g2_decap_8 FILLER_1_1603 ();
 sg13g2_decap_8 FILLER_1_1610 ();
 sg13g2_decap_8 FILLER_1_1617 ();
 sg13g2_decap_8 FILLER_1_1624 ();
 sg13g2_decap_8 FILLER_1_1631 ();
 sg13g2_decap_8 FILLER_1_1638 ();
 sg13g2_decap_8 FILLER_1_1645 ();
 sg13g2_decap_8 FILLER_1_1652 ();
 sg13g2_decap_8 FILLER_1_1659 ();
 sg13g2_decap_8 FILLER_1_1666 ();
 sg13g2_decap_8 FILLER_1_1673 ();
 sg13g2_decap_8 FILLER_1_1680 ();
 sg13g2_decap_8 FILLER_1_1687 ();
 sg13g2_decap_8 FILLER_1_1694 ();
 sg13g2_decap_8 FILLER_1_1701 ();
 sg13g2_decap_8 FILLER_1_1708 ();
 sg13g2_decap_8 FILLER_1_1715 ();
 sg13g2_decap_8 FILLER_1_1722 ();
 sg13g2_decap_8 FILLER_1_1729 ();
 sg13g2_decap_8 FILLER_1_1736 ();
 sg13g2_decap_8 FILLER_1_1743 ();
 sg13g2_decap_8 FILLER_1_1750 ();
 sg13g2_decap_8 FILLER_1_1757 ();
 sg13g2_decap_8 FILLER_1_1764 ();
 sg13g2_decap_8 FILLER_1_1771 ();
 sg13g2_decap_8 FILLER_1_1778 ();
 sg13g2_decap_8 FILLER_1_1785 ();
 sg13g2_decap_8 FILLER_1_1792 ();
 sg13g2_decap_8 FILLER_1_1799 ();
 sg13g2_decap_8 FILLER_1_1806 ();
 sg13g2_decap_8 FILLER_1_1813 ();
 sg13g2_decap_8 FILLER_1_1820 ();
 sg13g2_decap_8 FILLER_1_1827 ();
 sg13g2_decap_8 FILLER_1_1834 ();
 sg13g2_decap_8 FILLER_1_1841 ();
 sg13g2_decap_8 FILLER_1_1848 ();
 sg13g2_decap_8 FILLER_1_1855 ();
 sg13g2_decap_8 FILLER_1_1862 ();
 sg13g2_decap_8 FILLER_1_1869 ();
 sg13g2_decap_8 FILLER_1_1876 ();
 sg13g2_decap_8 FILLER_1_1883 ();
 sg13g2_decap_8 FILLER_1_1890 ();
 sg13g2_decap_8 FILLER_1_1897 ();
 sg13g2_decap_8 FILLER_1_1904 ();
 sg13g2_decap_8 FILLER_1_1911 ();
 sg13g2_decap_8 FILLER_1_1918 ();
 sg13g2_decap_8 FILLER_1_1925 ();
 sg13g2_decap_8 FILLER_1_1932 ();
 sg13g2_decap_8 FILLER_1_1939 ();
 sg13g2_decap_8 FILLER_1_1946 ();
 sg13g2_decap_8 FILLER_1_1953 ();
 sg13g2_decap_8 FILLER_1_1960 ();
 sg13g2_decap_8 FILLER_1_1967 ();
 sg13g2_decap_8 FILLER_1_1974 ();
 sg13g2_decap_8 FILLER_1_1981 ();
 sg13g2_decap_8 FILLER_1_1988 ();
 sg13g2_decap_8 FILLER_1_1995 ();
 sg13g2_decap_8 FILLER_1_2002 ();
 sg13g2_decap_8 FILLER_1_2009 ();
 sg13g2_decap_8 FILLER_1_2016 ();
 sg13g2_decap_8 FILLER_1_2023 ();
 sg13g2_decap_8 FILLER_1_2030 ();
 sg13g2_decap_8 FILLER_1_2037 ();
 sg13g2_decap_8 FILLER_1_2044 ();
 sg13g2_decap_8 FILLER_1_2051 ();
 sg13g2_decap_8 FILLER_1_2058 ();
 sg13g2_decap_8 FILLER_1_2065 ();
 sg13g2_decap_8 FILLER_1_2072 ();
 sg13g2_decap_8 FILLER_1_2079 ();
 sg13g2_decap_8 FILLER_1_2086 ();
 sg13g2_decap_8 FILLER_1_2093 ();
 sg13g2_decap_8 FILLER_1_2100 ();
 sg13g2_decap_8 FILLER_1_2107 ();
 sg13g2_decap_8 FILLER_1_2114 ();
 sg13g2_decap_8 FILLER_1_2121 ();
 sg13g2_decap_8 FILLER_1_2128 ();
 sg13g2_decap_8 FILLER_1_2135 ();
 sg13g2_decap_8 FILLER_1_2142 ();
 sg13g2_decap_8 FILLER_1_2149 ();
 sg13g2_decap_8 FILLER_1_2156 ();
 sg13g2_decap_8 FILLER_1_2163 ();
 sg13g2_decap_8 FILLER_1_2170 ();
 sg13g2_decap_8 FILLER_1_2177 ();
 sg13g2_decap_8 FILLER_1_2184 ();
 sg13g2_decap_8 FILLER_1_2191 ();
 sg13g2_decap_8 FILLER_1_2198 ();
 sg13g2_decap_8 FILLER_1_2205 ();
 sg13g2_decap_8 FILLER_1_2212 ();
 sg13g2_decap_8 FILLER_1_2219 ();
 sg13g2_decap_8 FILLER_1_2226 ();
 sg13g2_decap_8 FILLER_1_2233 ();
 sg13g2_decap_8 FILLER_1_2240 ();
 sg13g2_decap_8 FILLER_1_2247 ();
 sg13g2_decap_8 FILLER_1_2254 ();
 sg13g2_decap_8 FILLER_1_2261 ();
 sg13g2_decap_8 FILLER_1_2268 ();
 sg13g2_decap_8 FILLER_1_2275 ();
 sg13g2_decap_8 FILLER_1_2282 ();
 sg13g2_decap_8 FILLER_1_2289 ();
 sg13g2_decap_8 FILLER_1_2296 ();
 sg13g2_decap_8 FILLER_1_2303 ();
 sg13g2_decap_8 FILLER_1_2310 ();
 sg13g2_decap_8 FILLER_1_2317 ();
 sg13g2_decap_8 FILLER_1_2324 ();
 sg13g2_decap_8 FILLER_1_2331 ();
 sg13g2_decap_8 FILLER_1_2338 ();
 sg13g2_decap_8 FILLER_1_2345 ();
 sg13g2_decap_8 FILLER_1_2352 ();
 sg13g2_decap_8 FILLER_1_2359 ();
 sg13g2_decap_8 FILLER_1_2366 ();
 sg13g2_decap_8 FILLER_1_2373 ();
 sg13g2_decap_8 FILLER_1_2380 ();
 sg13g2_decap_8 FILLER_1_2387 ();
 sg13g2_decap_8 FILLER_1_2394 ();
 sg13g2_decap_8 FILLER_1_2401 ();
 sg13g2_decap_8 FILLER_1_2408 ();
 sg13g2_decap_8 FILLER_1_2415 ();
 sg13g2_decap_8 FILLER_1_2422 ();
 sg13g2_decap_8 FILLER_1_2429 ();
 sg13g2_decap_8 FILLER_1_2436 ();
 sg13g2_decap_8 FILLER_1_2443 ();
 sg13g2_decap_8 FILLER_1_2450 ();
 sg13g2_decap_8 FILLER_1_2457 ();
 sg13g2_decap_8 FILLER_1_2464 ();
 sg13g2_decap_8 FILLER_1_2471 ();
 sg13g2_decap_8 FILLER_1_2478 ();
 sg13g2_decap_8 FILLER_1_2485 ();
 sg13g2_decap_8 FILLER_1_2492 ();
 sg13g2_decap_8 FILLER_1_2499 ();
 sg13g2_decap_8 FILLER_1_2506 ();
 sg13g2_decap_8 FILLER_1_2513 ();
 sg13g2_decap_8 FILLER_1_2520 ();
 sg13g2_decap_8 FILLER_1_2527 ();
 sg13g2_decap_8 FILLER_1_2534 ();
 sg13g2_decap_8 FILLER_1_2541 ();
 sg13g2_decap_8 FILLER_1_2548 ();
 sg13g2_decap_8 FILLER_1_2555 ();
 sg13g2_decap_8 FILLER_1_2562 ();
 sg13g2_decap_8 FILLER_1_2569 ();
 sg13g2_decap_8 FILLER_1_2576 ();
 sg13g2_decap_8 FILLER_1_2583 ();
 sg13g2_decap_8 FILLER_1_2590 ();
 sg13g2_decap_8 FILLER_1_2597 ();
 sg13g2_decap_8 FILLER_1_2604 ();
 sg13g2_decap_8 FILLER_1_2611 ();
 sg13g2_decap_8 FILLER_1_2618 ();
 sg13g2_decap_8 FILLER_1_2625 ();
 sg13g2_decap_8 FILLER_1_2632 ();
 sg13g2_decap_8 FILLER_1_2639 ();
 sg13g2_decap_8 FILLER_1_2646 ();
 sg13g2_decap_8 FILLER_1_2653 ();
 sg13g2_decap_8 FILLER_1_2660 ();
 sg13g2_decap_8 FILLER_1_2667 ();
 sg13g2_decap_8 FILLER_1_2674 ();
 sg13g2_decap_8 FILLER_1_2681 ();
 sg13g2_decap_8 FILLER_1_2688 ();
 sg13g2_decap_8 FILLER_1_2695 ();
 sg13g2_decap_8 FILLER_1_2702 ();
 sg13g2_decap_8 FILLER_1_2709 ();
 sg13g2_decap_8 FILLER_1_2716 ();
 sg13g2_decap_8 FILLER_1_2723 ();
 sg13g2_decap_8 FILLER_1_2730 ();
 sg13g2_decap_8 FILLER_1_2737 ();
 sg13g2_decap_8 FILLER_1_2744 ();
 sg13g2_decap_8 FILLER_1_2751 ();
 sg13g2_decap_8 FILLER_1_2758 ();
 sg13g2_decap_8 FILLER_1_2765 ();
 sg13g2_decap_8 FILLER_1_2772 ();
 sg13g2_decap_8 FILLER_1_2779 ();
 sg13g2_decap_8 FILLER_1_2786 ();
 sg13g2_decap_8 FILLER_1_2793 ();
 sg13g2_decap_8 FILLER_1_2800 ();
 sg13g2_decap_8 FILLER_1_2807 ();
 sg13g2_decap_8 FILLER_1_2814 ();
 sg13g2_decap_8 FILLER_1_2821 ();
 sg13g2_decap_8 FILLER_1_2828 ();
 sg13g2_decap_8 FILLER_1_2835 ();
 sg13g2_decap_8 FILLER_1_2842 ();
 sg13g2_decap_8 FILLER_1_2849 ();
 sg13g2_decap_8 FILLER_1_2856 ();
 sg13g2_decap_8 FILLER_1_2863 ();
 sg13g2_decap_8 FILLER_1_2870 ();
 sg13g2_decap_8 FILLER_1_2877 ();
 sg13g2_decap_8 FILLER_1_2884 ();
 sg13g2_decap_8 FILLER_1_2891 ();
 sg13g2_decap_8 FILLER_1_2898 ();
 sg13g2_decap_8 FILLER_1_2905 ();
 sg13g2_decap_8 FILLER_1_2912 ();
 sg13g2_decap_8 FILLER_1_2919 ();
 sg13g2_decap_8 FILLER_1_2926 ();
 sg13g2_decap_8 FILLER_1_2933 ();
 sg13g2_decap_8 FILLER_1_2940 ();
 sg13g2_decap_8 FILLER_1_2947 ();
 sg13g2_decap_8 FILLER_1_2954 ();
 sg13g2_decap_8 FILLER_1_2961 ();
 sg13g2_decap_8 FILLER_1_2968 ();
 sg13g2_decap_8 FILLER_1_2975 ();
 sg13g2_decap_8 FILLER_1_2982 ();
 sg13g2_decap_8 FILLER_1_2989 ();
 sg13g2_decap_8 FILLER_1_2996 ();
 sg13g2_decap_8 FILLER_1_3003 ();
 sg13g2_decap_8 FILLER_1_3010 ();
 sg13g2_decap_8 FILLER_1_3017 ();
 sg13g2_decap_8 FILLER_1_3024 ();
 sg13g2_decap_8 FILLER_1_3031 ();
 sg13g2_decap_8 FILLER_1_3038 ();
 sg13g2_decap_8 FILLER_1_3045 ();
 sg13g2_decap_8 FILLER_1_3052 ();
 sg13g2_decap_8 FILLER_1_3059 ();
 sg13g2_decap_8 FILLER_1_3066 ();
 sg13g2_decap_8 FILLER_1_3073 ();
 sg13g2_decap_8 FILLER_1_3080 ();
 sg13g2_decap_8 FILLER_1_3087 ();
 sg13g2_decap_8 FILLER_1_3094 ();
 sg13g2_decap_8 FILLER_1_3101 ();
 sg13g2_decap_8 FILLER_1_3108 ();
 sg13g2_decap_8 FILLER_1_3115 ();
 sg13g2_decap_8 FILLER_1_3122 ();
 sg13g2_decap_8 FILLER_1_3129 ();
 sg13g2_decap_8 FILLER_1_3136 ();
 sg13g2_decap_8 FILLER_1_3143 ();
 sg13g2_decap_8 FILLER_1_3150 ();
 sg13g2_decap_8 FILLER_1_3157 ();
 sg13g2_decap_8 FILLER_1_3164 ();
 sg13g2_decap_8 FILLER_1_3171 ();
 sg13g2_decap_8 FILLER_1_3178 ();
 sg13g2_decap_8 FILLER_1_3185 ();
 sg13g2_decap_8 FILLER_1_3192 ();
 sg13g2_decap_8 FILLER_1_3199 ();
 sg13g2_decap_8 FILLER_1_3206 ();
 sg13g2_decap_8 FILLER_1_3213 ();
 sg13g2_decap_8 FILLER_1_3220 ();
 sg13g2_decap_8 FILLER_1_3227 ();
 sg13g2_decap_8 FILLER_1_3234 ();
 sg13g2_decap_8 FILLER_1_3241 ();
 sg13g2_decap_8 FILLER_1_3248 ();
 sg13g2_decap_8 FILLER_1_3255 ();
 sg13g2_decap_8 FILLER_1_3262 ();
 sg13g2_decap_8 FILLER_1_3269 ();
 sg13g2_decap_8 FILLER_1_3276 ();
 sg13g2_decap_8 FILLER_1_3283 ();
 sg13g2_decap_8 FILLER_1_3290 ();
 sg13g2_decap_8 FILLER_1_3297 ();
 sg13g2_decap_8 FILLER_1_3304 ();
 sg13g2_decap_8 FILLER_1_3311 ();
 sg13g2_decap_8 FILLER_1_3318 ();
 sg13g2_decap_8 FILLER_1_3325 ();
 sg13g2_decap_8 FILLER_1_3332 ();
 sg13g2_decap_8 FILLER_1_3339 ();
 sg13g2_decap_8 FILLER_1_3346 ();
 sg13g2_decap_8 FILLER_1_3353 ();
 sg13g2_decap_8 FILLER_1_3360 ();
 sg13g2_decap_8 FILLER_1_3367 ();
 sg13g2_decap_8 FILLER_1_3374 ();
 sg13g2_decap_8 FILLER_1_3381 ();
 sg13g2_decap_8 FILLER_1_3388 ();
 sg13g2_decap_8 FILLER_1_3395 ();
 sg13g2_decap_8 FILLER_1_3402 ();
 sg13g2_decap_8 FILLER_1_3409 ();
 sg13g2_decap_8 FILLER_1_3416 ();
 sg13g2_decap_8 FILLER_1_3423 ();
 sg13g2_decap_8 FILLER_1_3430 ();
 sg13g2_decap_8 FILLER_1_3437 ();
 sg13g2_decap_8 FILLER_1_3444 ();
 sg13g2_decap_8 FILLER_1_3451 ();
 sg13g2_decap_8 FILLER_1_3458 ();
 sg13g2_decap_8 FILLER_1_3465 ();
 sg13g2_decap_8 FILLER_1_3472 ();
 sg13g2_decap_8 FILLER_1_3479 ();
 sg13g2_decap_8 FILLER_1_3486 ();
 sg13g2_decap_8 FILLER_1_3493 ();
 sg13g2_decap_8 FILLER_1_3500 ();
 sg13g2_decap_8 FILLER_1_3507 ();
 sg13g2_decap_8 FILLER_1_3514 ();
 sg13g2_decap_8 FILLER_1_3521 ();
 sg13g2_decap_8 FILLER_1_3528 ();
 sg13g2_decap_8 FILLER_1_3535 ();
 sg13g2_decap_8 FILLER_1_3542 ();
 sg13g2_decap_8 FILLER_1_3549 ();
 sg13g2_decap_8 FILLER_1_3556 ();
 sg13g2_decap_8 FILLER_1_3563 ();
 sg13g2_decap_8 FILLER_1_3570 ();
 sg13g2_fill_2 FILLER_1_3577 ();
 sg13g2_fill_1 FILLER_1_3579 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_decap_8 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_2_868 ();
 sg13g2_decap_8 FILLER_2_875 ();
 sg13g2_decap_8 FILLER_2_882 ();
 sg13g2_decap_8 FILLER_2_889 ();
 sg13g2_decap_8 FILLER_2_896 ();
 sg13g2_decap_8 FILLER_2_903 ();
 sg13g2_decap_8 FILLER_2_910 ();
 sg13g2_decap_8 FILLER_2_917 ();
 sg13g2_decap_8 FILLER_2_924 ();
 sg13g2_decap_8 FILLER_2_931 ();
 sg13g2_decap_8 FILLER_2_938 ();
 sg13g2_decap_8 FILLER_2_945 ();
 sg13g2_decap_8 FILLER_2_952 ();
 sg13g2_decap_8 FILLER_2_959 ();
 sg13g2_decap_8 FILLER_2_966 ();
 sg13g2_decap_8 FILLER_2_973 ();
 sg13g2_decap_8 FILLER_2_980 ();
 sg13g2_decap_8 FILLER_2_987 ();
 sg13g2_decap_8 FILLER_2_994 ();
 sg13g2_decap_8 FILLER_2_1001 ();
 sg13g2_decap_8 FILLER_2_1008 ();
 sg13g2_decap_8 FILLER_2_1015 ();
 sg13g2_decap_8 FILLER_2_1022 ();
 sg13g2_decap_8 FILLER_2_1029 ();
 sg13g2_decap_8 FILLER_2_1036 ();
 sg13g2_decap_8 FILLER_2_1043 ();
 sg13g2_decap_8 FILLER_2_1050 ();
 sg13g2_decap_8 FILLER_2_1057 ();
 sg13g2_decap_8 FILLER_2_1064 ();
 sg13g2_decap_8 FILLER_2_1071 ();
 sg13g2_decap_8 FILLER_2_1078 ();
 sg13g2_decap_8 FILLER_2_1085 ();
 sg13g2_decap_8 FILLER_2_1092 ();
 sg13g2_decap_8 FILLER_2_1099 ();
 sg13g2_decap_8 FILLER_2_1106 ();
 sg13g2_decap_8 FILLER_2_1113 ();
 sg13g2_decap_8 FILLER_2_1120 ();
 sg13g2_decap_8 FILLER_2_1127 ();
 sg13g2_decap_8 FILLER_2_1134 ();
 sg13g2_decap_8 FILLER_2_1141 ();
 sg13g2_decap_8 FILLER_2_1148 ();
 sg13g2_decap_8 FILLER_2_1155 ();
 sg13g2_decap_8 FILLER_2_1162 ();
 sg13g2_decap_8 FILLER_2_1169 ();
 sg13g2_decap_8 FILLER_2_1176 ();
 sg13g2_decap_8 FILLER_2_1183 ();
 sg13g2_decap_8 FILLER_2_1190 ();
 sg13g2_decap_8 FILLER_2_1197 ();
 sg13g2_decap_8 FILLER_2_1204 ();
 sg13g2_decap_8 FILLER_2_1211 ();
 sg13g2_decap_8 FILLER_2_1218 ();
 sg13g2_decap_8 FILLER_2_1225 ();
 sg13g2_decap_8 FILLER_2_1232 ();
 sg13g2_decap_8 FILLER_2_1239 ();
 sg13g2_decap_8 FILLER_2_1246 ();
 sg13g2_decap_8 FILLER_2_1253 ();
 sg13g2_decap_8 FILLER_2_1260 ();
 sg13g2_decap_8 FILLER_2_1267 ();
 sg13g2_decap_8 FILLER_2_1274 ();
 sg13g2_decap_8 FILLER_2_1281 ();
 sg13g2_decap_8 FILLER_2_1288 ();
 sg13g2_decap_8 FILLER_2_1295 ();
 sg13g2_decap_8 FILLER_2_1302 ();
 sg13g2_decap_8 FILLER_2_1309 ();
 sg13g2_decap_8 FILLER_2_1316 ();
 sg13g2_decap_8 FILLER_2_1323 ();
 sg13g2_decap_8 FILLER_2_1330 ();
 sg13g2_decap_8 FILLER_2_1337 ();
 sg13g2_decap_8 FILLER_2_1344 ();
 sg13g2_decap_8 FILLER_2_1351 ();
 sg13g2_decap_8 FILLER_2_1358 ();
 sg13g2_decap_8 FILLER_2_1365 ();
 sg13g2_decap_8 FILLER_2_1372 ();
 sg13g2_decap_8 FILLER_2_1379 ();
 sg13g2_decap_8 FILLER_2_1386 ();
 sg13g2_decap_8 FILLER_2_1393 ();
 sg13g2_decap_8 FILLER_2_1400 ();
 sg13g2_decap_8 FILLER_2_1407 ();
 sg13g2_decap_8 FILLER_2_1414 ();
 sg13g2_decap_8 FILLER_2_1421 ();
 sg13g2_decap_8 FILLER_2_1428 ();
 sg13g2_decap_8 FILLER_2_1435 ();
 sg13g2_decap_8 FILLER_2_1442 ();
 sg13g2_decap_8 FILLER_2_1449 ();
 sg13g2_decap_8 FILLER_2_1456 ();
 sg13g2_decap_8 FILLER_2_1463 ();
 sg13g2_decap_8 FILLER_2_1470 ();
 sg13g2_decap_8 FILLER_2_1477 ();
 sg13g2_decap_8 FILLER_2_1484 ();
 sg13g2_decap_8 FILLER_2_1491 ();
 sg13g2_decap_8 FILLER_2_1498 ();
 sg13g2_decap_8 FILLER_2_1505 ();
 sg13g2_decap_8 FILLER_2_1512 ();
 sg13g2_decap_8 FILLER_2_1519 ();
 sg13g2_decap_8 FILLER_2_1526 ();
 sg13g2_decap_8 FILLER_2_1533 ();
 sg13g2_decap_8 FILLER_2_1540 ();
 sg13g2_decap_8 FILLER_2_1547 ();
 sg13g2_decap_8 FILLER_2_1554 ();
 sg13g2_decap_8 FILLER_2_1561 ();
 sg13g2_decap_8 FILLER_2_1568 ();
 sg13g2_decap_8 FILLER_2_1575 ();
 sg13g2_decap_8 FILLER_2_1582 ();
 sg13g2_decap_8 FILLER_2_1589 ();
 sg13g2_decap_8 FILLER_2_1596 ();
 sg13g2_decap_8 FILLER_2_1603 ();
 sg13g2_decap_8 FILLER_2_1610 ();
 sg13g2_decap_8 FILLER_2_1617 ();
 sg13g2_decap_8 FILLER_2_1624 ();
 sg13g2_decap_8 FILLER_2_1631 ();
 sg13g2_decap_8 FILLER_2_1638 ();
 sg13g2_decap_8 FILLER_2_1645 ();
 sg13g2_decap_8 FILLER_2_1652 ();
 sg13g2_decap_8 FILLER_2_1659 ();
 sg13g2_decap_8 FILLER_2_1666 ();
 sg13g2_decap_8 FILLER_2_1673 ();
 sg13g2_decap_8 FILLER_2_1680 ();
 sg13g2_decap_8 FILLER_2_1687 ();
 sg13g2_decap_8 FILLER_2_1694 ();
 sg13g2_decap_8 FILLER_2_1701 ();
 sg13g2_decap_8 FILLER_2_1708 ();
 sg13g2_decap_8 FILLER_2_1715 ();
 sg13g2_decap_8 FILLER_2_1722 ();
 sg13g2_decap_8 FILLER_2_1729 ();
 sg13g2_decap_8 FILLER_2_1736 ();
 sg13g2_decap_8 FILLER_2_1743 ();
 sg13g2_decap_8 FILLER_2_1750 ();
 sg13g2_decap_8 FILLER_2_1757 ();
 sg13g2_decap_8 FILLER_2_1764 ();
 sg13g2_decap_8 FILLER_2_1771 ();
 sg13g2_decap_8 FILLER_2_1778 ();
 sg13g2_decap_8 FILLER_2_1785 ();
 sg13g2_decap_8 FILLER_2_1792 ();
 sg13g2_decap_8 FILLER_2_1799 ();
 sg13g2_decap_8 FILLER_2_1806 ();
 sg13g2_decap_8 FILLER_2_1813 ();
 sg13g2_decap_8 FILLER_2_1820 ();
 sg13g2_decap_8 FILLER_2_1827 ();
 sg13g2_decap_8 FILLER_2_1834 ();
 sg13g2_decap_8 FILLER_2_1841 ();
 sg13g2_decap_8 FILLER_2_1848 ();
 sg13g2_decap_8 FILLER_2_1855 ();
 sg13g2_decap_8 FILLER_2_1862 ();
 sg13g2_decap_8 FILLER_2_1869 ();
 sg13g2_decap_8 FILLER_2_1876 ();
 sg13g2_decap_8 FILLER_2_1883 ();
 sg13g2_decap_8 FILLER_2_1890 ();
 sg13g2_decap_8 FILLER_2_1897 ();
 sg13g2_decap_8 FILLER_2_1904 ();
 sg13g2_decap_8 FILLER_2_1911 ();
 sg13g2_decap_8 FILLER_2_1918 ();
 sg13g2_decap_8 FILLER_2_1925 ();
 sg13g2_decap_8 FILLER_2_1932 ();
 sg13g2_decap_8 FILLER_2_1939 ();
 sg13g2_decap_8 FILLER_2_1946 ();
 sg13g2_decap_8 FILLER_2_1953 ();
 sg13g2_decap_8 FILLER_2_1960 ();
 sg13g2_decap_8 FILLER_2_1967 ();
 sg13g2_decap_8 FILLER_2_1974 ();
 sg13g2_decap_8 FILLER_2_1981 ();
 sg13g2_decap_8 FILLER_2_1988 ();
 sg13g2_decap_8 FILLER_2_1995 ();
 sg13g2_decap_8 FILLER_2_2002 ();
 sg13g2_decap_8 FILLER_2_2009 ();
 sg13g2_decap_8 FILLER_2_2016 ();
 sg13g2_decap_8 FILLER_2_2023 ();
 sg13g2_decap_8 FILLER_2_2030 ();
 sg13g2_decap_8 FILLER_2_2037 ();
 sg13g2_decap_8 FILLER_2_2044 ();
 sg13g2_decap_8 FILLER_2_2051 ();
 sg13g2_decap_8 FILLER_2_2058 ();
 sg13g2_decap_8 FILLER_2_2065 ();
 sg13g2_decap_8 FILLER_2_2072 ();
 sg13g2_decap_8 FILLER_2_2079 ();
 sg13g2_decap_8 FILLER_2_2086 ();
 sg13g2_decap_8 FILLER_2_2093 ();
 sg13g2_decap_8 FILLER_2_2100 ();
 sg13g2_decap_8 FILLER_2_2107 ();
 sg13g2_decap_8 FILLER_2_2114 ();
 sg13g2_decap_8 FILLER_2_2121 ();
 sg13g2_decap_8 FILLER_2_2128 ();
 sg13g2_decap_8 FILLER_2_2135 ();
 sg13g2_decap_8 FILLER_2_2142 ();
 sg13g2_decap_8 FILLER_2_2149 ();
 sg13g2_decap_8 FILLER_2_2156 ();
 sg13g2_decap_8 FILLER_2_2163 ();
 sg13g2_decap_8 FILLER_2_2170 ();
 sg13g2_decap_8 FILLER_2_2177 ();
 sg13g2_decap_8 FILLER_2_2184 ();
 sg13g2_decap_8 FILLER_2_2191 ();
 sg13g2_decap_8 FILLER_2_2198 ();
 sg13g2_decap_8 FILLER_2_2205 ();
 sg13g2_decap_8 FILLER_2_2212 ();
 sg13g2_decap_8 FILLER_2_2219 ();
 sg13g2_decap_8 FILLER_2_2226 ();
 sg13g2_decap_8 FILLER_2_2233 ();
 sg13g2_decap_8 FILLER_2_2240 ();
 sg13g2_decap_8 FILLER_2_2247 ();
 sg13g2_decap_8 FILLER_2_2254 ();
 sg13g2_decap_8 FILLER_2_2261 ();
 sg13g2_decap_8 FILLER_2_2268 ();
 sg13g2_decap_8 FILLER_2_2275 ();
 sg13g2_decap_8 FILLER_2_2282 ();
 sg13g2_decap_8 FILLER_2_2289 ();
 sg13g2_decap_8 FILLER_2_2296 ();
 sg13g2_decap_8 FILLER_2_2303 ();
 sg13g2_decap_8 FILLER_2_2310 ();
 sg13g2_decap_8 FILLER_2_2317 ();
 sg13g2_decap_8 FILLER_2_2324 ();
 sg13g2_decap_8 FILLER_2_2331 ();
 sg13g2_decap_8 FILLER_2_2338 ();
 sg13g2_decap_8 FILLER_2_2345 ();
 sg13g2_decap_8 FILLER_2_2352 ();
 sg13g2_decap_8 FILLER_2_2359 ();
 sg13g2_decap_8 FILLER_2_2366 ();
 sg13g2_decap_8 FILLER_2_2373 ();
 sg13g2_decap_8 FILLER_2_2380 ();
 sg13g2_decap_8 FILLER_2_2387 ();
 sg13g2_decap_8 FILLER_2_2394 ();
 sg13g2_decap_8 FILLER_2_2401 ();
 sg13g2_decap_8 FILLER_2_2408 ();
 sg13g2_decap_8 FILLER_2_2415 ();
 sg13g2_decap_8 FILLER_2_2422 ();
 sg13g2_decap_8 FILLER_2_2429 ();
 sg13g2_decap_8 FILLER_2_2436 ();
 sg13g2_decap_8 FILLER_2_2443 ();
 sg13g2_decap_8 FILLER_2_2450 ();
 sg13g2_decap_8 FILLER_2_2457 ();
 sg13g2_decap_8 FILLER_2_2464 ();
 sg13g2_decap_8 FILLER_2_2471 ();
 sg13g2_decap_8 FILLER_2_2478 ();
 sg13g2_decap_8 FILLER_2_2485 ();
 sg13g2_decap_8 FILLER_2_2492 ();
 sg13g2_decap_8 FILLER_2_2499 ();
 sg13g2_decap_8 FILLER_2_2506 ();
 sg13g2_decap_8 FILLER_2_2513 ();
 sg13g2_decap_8 FILLER_2_2520 ();
 sg13g2_decap_8 FILLER_2_2527 ();
 sg13g2_decap_8 FILLER_2_2534 ();
 sg13g2_decap_8 FILLER_2_2541 ();
 sg13g2_decap_8 FILLER_2_2548 ();
 sg13g2_decap_8 FILLER_2_2555 ();
 sg13g2_decap_8 FILLER_2_2562 ();
 sg13g2_decap_8 FILLER_2_2569 ();
 sg13g2_decap_8 FILLER_2_2576 ();
 sg13g2_decap_8 FILLER_2_2583 ();
 sg13g2_decap_8 FILLER_2_2590 ();
 sg13g2_decap_8 FILLER_2_2597 ();
 sg13g2_decap_8 FILLER_2_2604 ();
 sg13g2_decap_8 FILLER_2_2611 ();
 sg13g2_decap_8 FILLER_2_2618 ();
 sg13g2_decap_8 FILLER_2_2625 ();
 sg13g2_decap_8 FILLER_2_2632 ();
 sg13g2_decap_8 FILLER_2_2639 ();
 sg13g2_decap_8 FILLER_2_2646 ();
 sg13g2_decap_8 FILLER_2_2653 ();
 sg13g2_decap_8 FILLER_2_2660 ();
 sg13g2_decap_8 FILLER_2_2667 ();
 sg13g2_decap_8 FILLER_2_2674 ();
 sg13g2_decap_8 FILLER_2_2681 ();
 sg13g2_decap_8 FILLER_2_2688 ();
 sg13g2_decap_8 FILLER_2_2695 ();
 sg13g2_decap_8 FILLER_2_2702 ();
 sg13g2_decap_8 FILLER_2_2709 ();
 sg13g2_decap_8 FILLER_2_2716 ();
 sg13g2_decap_8 FILLER_2_2723 ();
 sg13g2_decap_8 FILLER_2_2730 ();
 sg13g2_decap_8 FILLER_2_2737 ();
 sg13g2_decap_8 FILLER_2_2744 ();
 sg13g2_decap_8 FILLER_2_2751 ();
 sg13g2_decap_8 FILLER_2_2758 ();
 sg13g2_decap_8 FILLER_2_2765 ();
 sg13g2_decap_8 FILLER_2_2772 ();
 sg13g2_decap_8 FILLER_2_2779 ();
 sg13g2_decap_8 FILLER_2_2786 ();
 sg13g2_decap_8 FILLER_2_2793 ();
 sg13g2_decap_8 FILLER_2_2800 ();
 sg13g2_decap_8 FILLER_2_2807 ();
 sg13g2_decap_8 FILLER_2_2814 ();
 sg13g2_decap_8 FILLER_2_2821 ();
 sg13g2_decap_8 FILLER_2_2828 ();
 sg13g2_decap_8 FILLER_2_2835 ();
 sg13g2_decap_8 FILLER_2_2842 ();
 sg13g2_decap_8 FILLER_2_2849 ();
 sg13g2_decap_8 FILLER_2_2856 ();
 sg13g2_decap_8 FILLER_2_2863 ();
 sg13g2_decap_8 FILLER_2_2870 ();
 sg13g2_decap_8 FILLER_2_2877 ();
 sg13g2_decap_8 FILLER_2_2884 ();
 sg13g2_decap_8 FILLER_2_2891 ();
 sg13g2_decap_8 FILLER_2_2898 ();
 sg13g2_decap_8 FILLER_2_2905 ();
 sg13g2_decap_8 FILLER_2_2912 ();
 sg13g2_decap_8 FILLER_2_2919 ();
 sg13g2_decap_8 FILLER_2_2926 ();
 sg13g2_decap_8 FILLER_2_2933 ();
 sg13g2_decap_8 FILLER_2_2940 ();
 sg13g2_decap_8 FILLER_2_2947 ();
 sg13g2_decap_8 FILLER_2_2954 ();
 sg13g2_decap_8 FILLER_2_2961 ();
 sg13g2_decap_8 FILLER_2_2968 ();
 sg13g2_decap_8 FILLER_2_2975 ();
 sg13g2_decap_8 FILLER_2_2982 ();
 sg13g2_decap_8 FILLER_2_2989 ();
 sg13g2_decap_8 FILLER_2_2996 ();
 sg13g2_decap_8 FILLER_2_3003 ();
 sg13g2_decap_8 FILLER_2_3010 ();
 sg13g2_decap_8 FILLER_2_3017 ();
 sg13g2_decap_8 FILLER_2_3024 ();
 sg13g2_decap_8 FILLER_2_3031 ();
 sg13g2_decap_8 FILLER_2_3038 ();
 sg13g2_decap_8 FILLER_2_3045 ();
 sg13g2_decap_8 FILLER_2_3052 ();
 sg13g2_decap_8 FILLER_2_3059 ();
 sg13g2_decap_8 FILLER_2_3066 ();
 sg13g2_decap_8 FILLER_2_3073 ();
 sg13g2_decap_8 FILLER_2_3080 ();
 sg13g2_decap_8 FILLER_2_3087 ();
 sg13g2_decap_8 FILLER_2_3094 ();
 sg13g2_decap_8 FILLER_2_3101 ();
 sg13g2_decap_8 FILLER_2_3108 ();
 sg13g2_decap_8 FILLER_2_3115 ();
 sg13g2_decap_8 FILLER_2_3122 ();
 sg13g2_decap_8 FILLER_2_3129 ();
 sg13g2_decap_8 FILLER_2_3136 ();
 sg13g2_decap_8 FILLER_2_3143 ();
 sg13g2_decap_8 FILLER_2_3150 ();
 sg13g2_decap_8 FILLER_2_3157 ();
 sg13g2_decap_8 FILLER_2_3164 ();
 sg13g2_decap_8 FILLER_2_3171 ();
 sg13g2_decap_8 FILLER_2_3178 ();
 sg13g2_decap_8 FILLER_2_3185 ();
 sg13g2_decap_8 FILLER_2_3192 ();
 sg13g2_decap_8 FILLER_2_3199 ();
 sg13g2_decap_8 FILLER_2_3206 ();
 sg13g2_decap_8 FILLER_2_3213 ();
 sg13g2_decap_8 FILLER_2_3220 ();
 sg13g2_decap_8 FILLER_2_3227 ();
 sg13g2_decap_8 FILLER_2_3234 ();
 sg13g2_decap_8 FILLER_2_3241 ();
 sg13g2_decap_8 FILLER_2_3248 ();
 sg13g2_decap_8 FILLER_2_3255 ();
 sg13g2_decap_8 FILLER_2_3262 ();
 sg13g2_decap_8 FILLER_2_3269 ();
 sg13g2_decap_8 FILLER_2_3276 ();
 sg13g2_decap_8 FILLER_2_3283 ();
 sg13g2_decap_8 FILLER_2_3290 ();
 sg13g2_decap_8 FILLER_2_3297 ();
 sg13g2_decap_8 FILLER_2_3304 ();
 sg13g2_decap_8 FILLER_2_3311 ();
 sg13g2_decap_8 FILLER_2_3318 ();
 sg13g2_decap_8 FILLER_2_3325 ();
 sg13g2_decap_8 FILLER_2_3332 ();
 sg13g2_decap_8 FILLER_2_3339 ();
 sg13g2_decap_8 FILLER_2_3346 ();
 sg13g2_decap_8 FILLER_2_3353 ();
 sg13g2_decap_8 FILLER_2_3360 ();
 sg13g2_decap_8 FILLER_2_3367 ();
 sg13g2_decap_8 FILLER_2_3374 ();
 sg13g2_decap_8 FILLER_2_3381 ();
 sg13g2_decap_8 FILLER_2_3388 ();
 sg13g2_decap_8 FILLER_2_3395 ();
 sg13g2_decap_8 FILLER_2_3402 ();
 sg13g2_decap_8 FILLER_2_3409 ();
 sg13g2_decap_8 FILLER_2_3416 ();
 sg13g2_decap_8 FILLER_2_3423 ();
 sg13g2_decap_8 FILLER_2_3430 ();
 sg13g2_decap_8 FILLER_2_3437 ();
 sg13g2_decap_8 FILLER_2_3444 ();
 sg13g2_decap_8 FILLER_2_3451 ();
 sg13g2_decap_8 FILLER_2_3458 ();
 sg13g2_decap_8 FILLER_2_3465 ();
 sg13g2_decap_8 FILLER_2_3472 ();
 sg13g2_decap_8 FILLER_2_3479 ();
 sg13g2_decap_8 FILLER_2_3486 ();
 sg13g2_decap_8 FILLER_2_3493 ();
 sg13g2_decap_8 FILLER_2_3500 ();
 sg13g2_decap_8 FILLER_2_3507 ();
 sg13g2_decap_8 FILLER_2_3514 ();
 sg13g2_decap_8 FILLER_2_3521 ();
 sg13g2_decap_8 FILLER_2_3528 ();
 sg13g2_decap_8 FILLER_2_3535 ();
 sg13g2_decap_8 FILLER_2_3542 ();
 sg13g2_decap_8 FILLER_2_3549 ();
 sg13g2_decap_8 FILLER_2_3556 ();
 sg13g2_decap_8 FILLER_2_3563 ();
 sg13g2_decap_8 FILLER_2_3570 ();
 sg13g2_fill_2 FILLER_2_3577 ();
 sg13g2_fill_1 FILLER_2_3579 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_decap_8 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_3_868 ();
 sg13g2_decap_8 FILLER_3_875 ();
 sg13g2_decap_8 FILLER_3_882 ();
 sg13g2_decap_8 FILLER_3_889 ();
 sg13g2_decap_8 FILLER_3_896 ();
 sg13g2_decap_8 FILLER_3_903 ();
 sg13g2_decap_8 FILLER_3_910 ();
 sg13g2_decap_8 FILLER_3_917 ();
 sg13g2_decap_8 FILLER_3_924 ();
 sg13g2_decap_8 FILLER_3_931 ();
 sg13g2_decap_8 FILLER_3_938 ();
 sg13g2_decap_8 FILLER_3_945 ();
 sg13g2_decap_8 FILLER_3_952 ();
 sg13g2_decap_8 FILLER_3_959 ();
 sg13g2_decap_8 FILLER_3_966 ();
 sg13g2_decap_8 FILLER_3_973 ();
 sg13g2_decap_8 FILLER_3_980 ();
 sg13g2_decap_8 FILLER_3_987 ();
 sg13g2_decap_8 FILLER_3_994 ();
 sg13g2_decap_8 FILLER_3_1001 ();
 sg13g2_decap_8 FILLER_3_1008 ();
 sg13g2_decap_8 FILLER_3_1015 ();
 sg13g2_decap_8 FILLER_3_1022 ();
 sg13g2_decap_8 FILLER_3_1029 ();
 sg13g2_decap_8 FILLER_3_1036 ();
 sg13g2_decap_8 FILLER_3_1043 ();
 sg13g2_decap_8 FILLER_3_1050 ();
 sg13g2_decap_8 FILLER_3_1057 ();
 sg13g2_decap_8 FILLER_3_1064 ();
 sg13g2_decap_8 FILLER_3_1071 ();
 sg13g2_decap_8 FILLER_3_1078 ();
 sg13g2_decap_8 FILLER_3_1085 ();
 sg13g2_decap_8 FILLER_3_1092 ();
 sg13g2_decap_8 FILLER_3_1099 ();
 sg13g2_decap_8 FILLER_3_1106 ();
 sg13g2_decap_8 FILLER_3_1113 ();
 sg13g2_decap_8 FILLER_3_1120 ();
 sg13g2_decap_8 FILLER_3_1127 ();
 sg13g2_decap_8 FILLER_3_1134 ();
 sg13g2_decap_8 FILLER_3_1141 ();
 sg13g2_decap_8 FILLER_3_1148 ();
 sg13g2_decap_8 FILLER_3_1155 ();
 sg13g2_decap_8 FILLER_3_1162 ();
 sg13g2_decap_8 FILLER_3_1169 ();
 sg13g2_decap_8 FILLER_3_1176 ();
 sg13g2_decap_8 FILLER_3_1183 ();
 sg13g2_decap_8 FILLER_3_1190 ();
 sg13g2_decap_8 FILLER_3_1197 ();
 sg13g2_decap_8 FILLER_3_1204 ();
 sg13g2_decap_8 FILLER_3_1211 ();
 sg13g2_decap_8 FILLER_3_1218 ();
 sg13g2_decap_8 FILLER_3_1225 ();
 sg13g2_decap_8 FILLER_3_1232 ();
 sg13g2_decap_8 FILLER_3_1239 ();
 sg13g2_decap_8 FILLER_3_1246 ();
 sg13g2_decap_8 FILLER_3_1253 ();
 sg13g2_decap_8 FILLER_3_1260 ();
 sg13g2_decap_8 FILLER_3_1267 ();
 sg13g2_decap_8 FILLER_3_1274 ();
 sg13g2_decap_8 FILLER_3_1281 ();
 sg13g2_decap_8 FILLER_3_1288 ();
 sg13g2_decap_8 FILLER_3_1295 ();
 sg13g2_decap_8 FILLER_3_1302 ();
 sg13g2_decap_8 FILLER_3_1309 ();
 sg13g2_decap_8 FILLER_3_1316 ();
 sg13g2_decap_8 FILLER_3_1323 ();
 sg13g2_decap_8 FILLER_3_1330 ();
 sg13g2_decap_8 FILLER_3_1337 ();
 sg13g2_decap_8 FILLER_3_1344 ();
 sg13g2_decap_8 FILLER_3_1351 ();
 sg13g2_decap_8 FILLER_3_1358 ();
 sg13g2_decap_8 FILLER_3_1365 ();
 sg13g2_decap_8 FILLER_3_1372 ();
 sg13g2_decap_8 FILLER_3_1379 ();
 sg13g2_decap_8 FILLER_3_1386 ();
 sg13g2_decap_8 FILLER_3_1393 ();
 sg13g2_decap_8 FILLER_3_1400 ();
 sg13g2_decap_8 FILLER_3_1407 ();
 sg13g2_decap_8 FILLER_3_1414 ();
 sg13g2_decap_8 FILLER_3_1421 ();
 sg13g2_decap_8 FILLER_3_1428 ();
 sg13g2_decap_8 FILLER_3_1435 ();
 sg13g2_decap_8 FILLER_3_1442 ();
 sg13g2_decap_8 FILLER_3_1449 ();
 sg13g2_decap_8 FILLER_3_1456 ();
 sg13g2_decap_8 FILLER_3_1463 ();
 sg13g2_decap_8 FILLER_3_1470 ();
 sg13g2_decap_8 FILLER_3_1477 ();
 sg13g2_decap_8 FILLER_3_1484 ();
 sg13g2_decap_8 FILLER_3_1491 ();
 sg13g2_decap_8 FILLER_3_1498 ();
 sg13g2_decap_8 FILLER_3_1505 ();
 sg13g2_decap_8 FILLER_3_1512 ();
 sg13g2_decap_8 FILLER_3_1519 ();
 sg13g2_decap_8 FILLER_3_1526 ();
 sg13g2_decap_8 FILLER_3_1533 ();
 sg13g2_decap_8 FILLER_3_1540 ();
 sg13g2_decap_8 FILLER_3_1547 ();
 sg13g2_decap_8 FILLER_3_1554 ();
 sg13g2_decap_8 FILLER_3_1561 ();
 sg13g2_decap_8 FILLER_3_1568 ();
 sg13g2_decap_8 FILLER_3_1575 ();
 sg13g2_decap_8 FILLER_3_1582 ();
 sg13g2_decap_8 FILLER_3_1589 ();
 sg13g2_decap_8 FILLER_3_1596 ();
 sg13g2_decap_8 FILLER_3_1603 ();
 sg13g2_decap_8 FILLER_3_1610 ();
 sg13g2_decap_8 FILLER_3_1617 ();
 sg13g2_decap_8 FILLER_3_1624 ();
 sg13g2_decap_8 FILLER_3_1631 ();
 sg13g2_decap_8 FILLER_3_1638 ();
 sg13g2_decap_8 FILLER_3_1645 ();
 sg13g2_decap_8 FILLER_3_1652 ();
 sg13g2_decap_8 FILLER_3_1659 ();
 sg13g2_decap_8 FILLER_3_1666 ();
 sg13g2_decap_8 FILLER_3_1673 ();
 sg13g2_decap_8 FILLER_3_1680 ();
 sg13g2_decap_8 FILLER_3_1687 ();
 sg13g2_decap_8 FILLER_3_1694 ();
 sg13g2_decap_8 FILLER_3_1701 ();
 sg13g2_decap_8 FILLER_3_1708 ();
 sg13g2_decap_8 FILLER_3_1715 ();
 sg13g2_decap_8 FILLER_3_1722 ();
 sg13g2_decap_8 FILLER_3_1729 ();
 sg13g2_decap_8 FILLER_3_1736 ();
 sg13g2_decap_8 FILLER_3_1743 ();
 sg13g2_decap_8 FILLER_3_1750 ();
 sg13g2_decap_8 FILLER_3_1757 ();
 sg13g2_decap_8 FILLER_3_1764 ();
 sg13g2_decap_8 FILLER_3_1771 ();
 sg13g2_decap_8 FILLER_3_1778 ();
 sg13g2_decap_8 FILLER_3_1785 ();
 sg13g2_decap_8 FILLER_3_1792 ();
 sg13g2_decap_8 FILLER_3_1799 ();
 sg13g2_decap_8 FILLER_3_1806 ();
 sg13g2_decap_8 FILLER_3_1813 ();
 sg13g2_decap_8 FILLER_3_1820 ();
 sg13g2_decap_8 FILLER_3_1827 ();
 sg13g2_decap_8 FILLER_3_1834 ();
 sg13g2_decap_8 FILLER_3_1841 ();
 sg13g2_decap_8 FILLER_3_1848 ();
 sg13g2_decap_8 FILLER_3_1855 ();
 sg13g2_decap_8 FILLER_3_1862 ();
 sg13g2_decap_8 FILLER_3_1869 ();
 sg13g2_decap_8 FILLER_3_1876 ();
 sg13g2_decap_8 FILLER_3_1883 ();
 sg13g2_decap_8 FILLER_3_1890 ();
 sg13g2_decap_8 FILLER_3_1897 ();
 sg13g2_decap_8 FILLER_3_1904 ();
 sg13g2_decap_8 FILLER_3_1911 ();
 sg13g2_decap_8 FILLER_3_1918 ();
 sg13g2_decap_8 FILLER_3_1925 ();
 sg13g2_decap_8 FILLER_3_1932 ();
 sg13g2_decap_8 FILLER_3_1939 ();
 sg13g2_decap_8 FILLER_3_1946 ();
 sg13g2_decap_8 FILLER_3_1953 ();
 sg13g2_decap_8 FILLER_3_1960 ();
 sg13g2_decap_8 FILLER_3_1967 ();
 sg13g2_decap_8 FILLER_3_1974 ();
 sg13g2_decap_8 FILLER_3_1981 ();
 sg13g2_decap_8 FILLER_3_1988 ();
 sg13g2_decap_8 FILLER_3_1995 ();
 sg13g2_decap_8 FILLER_3_2002 ();
 sg13g2_decap_8 FILLER_3_2009 ();
 sg13g2_decap_8 FILLER_3_2016 ();
 sg13g2_decap_8 FILLER_3_2023 ();
 sg13g2_decap_8 FILLER_3_2030 ();
 sg13g2_decap_8 FILLER_3_2037 ();
 sg13g2_decap_8 FILLER_3_2044 ();
 sg13g2_decap_8 FILLER_3_2051 ();
 sg13g2_decap_8 FILLER_3_2058 ();
 sg13g2_decap_8 FILLER_3_2065 ();
 sg13g2_decap_8 FILLER_3_2072 ();
 sg13g2_decap_8 FILLER_3_2079 ();
 sg13g2_decap_8 FILLER_3_2086 ();
 sg13g2_decap_8 FILLER_3_2093 ();
 sg13g2_decap_8 FILLER_3_2100 ();
 sg13g2_decap_8 FILLER_3_2107 ();
 sg13g2_decap_8 FILLER_3_2114 ();
 sg13g2_decap_8 FILLER_3_2121 ();
 sg13g2_decap_8 FILLER_3_2128 ();
 sg13g2_decap_8 FILLER_3_2135 ();
 sg13g2_decap_8 FILLER_3_2142 ();
 sg13g2_decap_8 FILLER_3_2149 ();
 sg13g2_decap_8 FILLER_3_2156 ();
 sg13g2_decap_8 FILLER_3_2163 ();
 sg13g2_decap_8 FILLER_3_2170 ();
 sg13g2_decap_8 FILLER_3_2177 ();
 sg13g2_decap_8 FILLER_3_2184 ();
 sg13g2_decap_8 FILLER_3_2191 ();
 sg13g2_decap_8 FILLER_3_2198 ();
 sg13g2_decap_8 FILLER_3_2205 ();
 sg13g2_decap_8 FILLER_3_2212 ();
 sg13g2_decap_8 FILLER_3_2219 ();
 sg13g2_decap_8 FILLER_3_2226 ();
 sg13g2_decap_8 FILLER_3_2233 ();
 sg13g2_decap_8 FILLER_3_2240 ();
 sg13g2_decap_8 FILLER_3_2247 ();
 sg13g2_decap_8 FILLER_3_2254 ();
 sg13g2_decap_8 FILLER_3_2261 ();
 sg13g2_decap_8 FILLER_3_2268 ();
 sg13g2_decap_8 FILLER_3_2275 ();
 sg13g2_decap_8 FILLER_3_2282 ();
 sg13g2_decap_8 FILLER_3_2289 ();
 sg13g2_decap_8 FILLER_3_2296 ();
 sg13g2_decap_8 FILLER_3_2303 ();
 sg13g2_decap_8 FILLER_3_2310 ();
 sg13g2_decap_8 FILLER_3_2317 ();
 sg13g2_decap_8 FILLER_3_2324 ();
 sg13g2_decap_8 FILLER_3_2331 ();
 sg13g2_decap_8 FILLER_3_2338 ();
 sg13g2_decap_8 FILLER_3_2345 ();
 sg13g2_decap_8 FILLER_3_2352 ();
 sg13g2_decap_8 FILLER_3_2359 ();
 sg13g2_decap_8 FILLER_3_2366 ();
 sg13g2_decap_8 FILLER_3_2373 ();
 sg13g2_decap_8 FILLER_3_2380 ();
 sg13g2_decap_8 FILLER_3_2387 ();
 sg13g2_decap_8 FILLER_3_2394 ();
 sg13g2_decap_8 FILLER_3_2401 ();
 sg13g2_decap_8 FILLER_3_2408 ();
 sg13g2_decap_8 FILLER_3_2415 ();
 sg13g2_decap_8 FILLER_3_2422 ();
 sg13g2_decap_8 FILLER_3_2429 ();
 sg13g2_decap_8 FILLER_3_2436 ();
 sg13g2_decap_8 FILLER_3_2443 ();
 sg13g2_decap_8 FILLER_3_2450 ();
 sg13g2_decap_8 FILLER_3_2457 ();
 sg13g2_decap_8 FILLER_3_2464 ();
 sg13g2_decap_8 FILLER_3_2471 ();
 sg13g2_decap_8 FILLER_3_2478 ();
 sg13g2_decap_8 FILLER_3_2485 ();
 sg13g2_decap_8 FILLER_3_2492 ();
 sg13g2_decap_8 FILLER_3_2499 ();
 sg13g2_decap_8 FILLER_3_2506 ();
 sg13g2_decap_8 FILLER_3_2513 ();
 sg13g2_decap_8 FILLER_3_2520 ();
 sg13g2_decap_8 FILLER_3_2527 ();
 sg13g2_decap_8 FILLER_3_2534 ();
 sg13g2_decap_8 FILLER_3_2541 ();
 sg13g2_decap_8 FILLER_3_2548 ();
 sg13g2_decap_8 FILLER_3_2555 ();
 sg13g2_decap_8 FILLER_3_2562 ();
 sg13g2_decap_8 FILLER_3_2569 ();
 sg13g2_decap_8 FILLER_3_2576 ();
 sg13g2_decap_8 FILLER_3_2583 ();
 sg13g2_decap_8 FILLER_3_2590 ();
 sg13g2_decap_8 FILLER_3_2597 ();
 sg13g2_decap_8 FILLER_3_2604 ();
 sg13g2_decap_8 FILLER_3_2611 ();
 sg13g2_decap_8 FILLER_3_2618 ();
 sg13g2_decap_8 FILLER_3_2625 ();
 sg13g2_decap_8 FILLER_3_2632 ();
 sg13g2_decap_8 FILLER_3_2639 ();
 sg13g2_decap_8 FILLER_3_2646 ();
 sg13g2_decap_8 FILLER_3_2653 ();
 sg13g2_decap_8 FILLER_3_2660 ();
 sg13g2_decap_8 FILLER_3_2667 ();
 sg13g2_decap_8 FILLER_3_2674 ();
 sg13g2_decap_8 FILLER_3_2681 ();
 sg13g2_decap_8 FILLER_3_2688 ();
 sg13g2_decap_8 FILLER_3_2695 ();
 sg13g2_decap_8 FILLER_3_2702 ();
 sg13g2_decap_8 FILLER_3_2709 ();
 sg13g2_decap_8 FILLER_3_2716 ();
 sg13g2_decap_8 FILLER_3_2723 ();
 sg13g2_decap_8 FILLER_3_2730 ();
 sg13g2_decap_8 FILLER_3_2737 ();
 sg13g2_decap_8 FILLER_3_2744 ();
 sg13g2_decap_8 FILLER_3_2751 ();
 sg13g2_decap_8 FILLER_3_2758 ();
 sg13g2_decap_8 FILLER_3_2765 ();
 sg13g2_decap_8 FILLER_3_2772 ();
 sg13g2_decap_8 FILLER_3_2779 ();
 sg13g2_decap_8 FILLER_3_2786 ();
 sg13g2_decap_8 FILLER_3_2793 ();
 sg13g2_decap_8 FILLER_3_2800 ();
 sg13g2_decap_8 FILLER_3_2807 ();
 sg13g2_decap_8 FILLER_3_2814 ();
 sg13g2_decap_8 FILLER_3_2821 ();
 sg13g2_decap_8 FILLER_3_2828 ();
 sg13g2_decap_8 FILLER_3_2835 ();
 sg13g2_decap_8 FILLER_3_2842 ();
 sg13g2_decap_8 FILLER_3_2849 ();
 sg13g2_decap_8 FILLER_3_2856 ();
 sg13g2_decap_8 FILLER_3_2863 ();
 sg13g2_decap_8 FILLER_3_2870 ();
 sg13g2_decap_8 FILLER_3_2877 ();
 sg13g2_decap_8 FILLER_3_2884 ();
 sg13g2_decap_8 FILLER_3_2891 ();
 sg13g2_decap_8 FILLER_3_2898 ();
 sg13g2_decap_8 FILLER_3_2905 ();
 sg13g2_decap_8 FILLER_3_2912 ();
 sg13g2_decap_8 FILLER_3_2919 ();
 sg13g2_decap_8 FILLER_3_2926 ();
 sg13g2_decap_8 FILLER_3_2933 ();
 sg13g2_decap_8 FILLER_3_2940 ();
 sg13g2_decap_8 FILLER_3_2947 ();
 sg13g2_decap_8 FILLER_3_2954 ();
 sg13g2_decap_8 FILLER_3_2961 ();
 sg13g2_decap_8 FILLER_3_2968 ();
 sg13g2_decap_8 FILLER_3_2975 ();
 sg13g2_decap_8 FILLER_3_2982 ();
 sg13g2_decap_8 FILLER_3_2989 ();
 sg13g2_decap_8 FILLER_3_2996 ();
 sg13g2_decap_8 FILLER_3_3003 ();
 sg13g2_decap_8 FILLER_3_3010 ();
 sg13g2_decap_8 FILLER_3_3017 ();
 sg13g2_decap_8 FILLER_3_3024 ();
 sg13g2_decap_8 FILLER_3_3031 ();
 sg13g2_decap_8 FILLER_3_3038 ();
 sg13g2_decap_8 FILLER_3_3045 ();
 sg13g2_decap_8 FILLER_3_3052 ();
 sg13g2_decap_8 FILLER_3_3059 ();
 sg13g2_decap_8 FILLER_3_3066 ();
 sg13g2_decap_8 FILLER_3_3073 ();
 sg13g2_decap_8 FILLER_3_3080 ();
 sg13g2_decap_8 FILLER_3_3087 ();
 sg13g2_decap_8 FILLER_3_3094 ();
 sg13g2_decap_8 FILLER_3_3101 ();
 sg13g2_decap_8 FILLER_3_3108 ();
 sg13g2_decap_8 FILLER_3_3115 ();
 sg13g2_decap_8 FILLER_3_3122 ();
 sg13g2_decap_8 FILLER_3_3129 ();
 sg13g2_decap_8 FILLER_3_3136 ();
 sg13g2_decap_8 FILLER_3_3143 ();
 sg13g2_decap_8 FILLER_3_3150 ();
 sg13g2_decap_8 FILLER_3_3157 ();
 sg13g2_decap_8 FILLER_3_3164 ();
 sg13g2_decap_8 FILLER_3_3171 ();
 sg13g2_decap_8 FILLER_3_3178 ();
 sg13g2_decap_8 FILLER_3_3185 ();
 sg13g2_decap_8 FILLER_3_3192 ();
 sg13g2_decap_8 FILLER_3_3199 ();
 sg13g2_decap_8 FILLER_3_3206 ();
 sg13g2_decap_8 FILLER_3_3213 ();
 sg13g2_decap_8 FILLER_3_3220 ();
 sg13g2_decap_8 FILLER_3_3227 ();
 sg13g2_decap_8 FILLER_3_3234 ();
 sg13g2_decap_8 FILLER_3_3241 ();
 sg13g2_decap_8 FILLER_3_3248 ();
 sg13g2_decap_8 FILLER_3_3255 ();
 sg13g2_decap_8 FILLER_3_3262 ();
 sg13g2_decap_8 FILLER_3_3269 ();
 sg13g2_decap_8 FILLER_3_3276 ();
 sg13g2_decap_8 FILLER_3_3283 ();
 sg13g2_decap_8 FILLER_3_3290 ();
 sg13g2_decap_8 FILLER_3_3297 ();
 sg13g2_decap_8 FILLER_3_3304 ();
 sg13g2_decap_8 FILLER_3_3311 ();
 sg13g2_decap_8 FILLER_3_3318 ();
 sg13g2_decap_8 FILLER_3_3325 ();
 sg13g2_decap_8 FILLER_3_3332 ();
 sg13g2_decap_8 FILLER_3_3339 ();
 sg13g2_decap_8 FILLER_3_3346 ();
 sg13g2_decap_8 FILLER_3_3353 ();
 sg13g2_decap_8 FILLER_3_3360 ();
 sg13g2_decap_8 FILLER_3_3367 ();
 sg13g2_decap_8 FILLER_3_3374 ();
 sg13g2_decap_8 FILLER_3_3381 ();
 sg13g2_decap_8 FILLER_3_3388 ();
 sg13g2_decap_8 FILLER_3_3395 ();
 sg13g2_decap_8 FILLER_3_3402 ();
 sg13g2_decap_8 FILLER_3_3409 ();
 sg13g2_decap_8 FILLER_3_3416 ();
 sg13g2_decap_8 FILLER_3_3423 ();
 sg13g2_decap_8 FILLER_3_3430 ();
 sg13g2_decap_8 FILLER_3_3437 ();
 sg13g2_decap_8 FILLER_3_3444 ();
 sg13g2_decap_8 FILLER_3_3451 ();
 sg13g2_decap_8 FILLER_3_3458 ();
 sg13g2_decap_8 FILLER_3_3465 ();
 sg13g2_decap_8 FILLER_3_3472 ();
 sg13g2_decap_8 FILLER_3_3479 ();
 sg13g2_decap_8 FILLER_3_3486 ();
 sg13g2_decap_8 FILLER_3_3493 ();
 sg13g2_decap_8 FILLER_3_3500 ();
 sg13g2_decap_8 FILLER_3_3507 ();
 sg13g2_decap_8 FILLER_3_3514 ();
 sg13g2_decap_8 FILLER_3_3521 ();
 sg13g2_decap_8 FILLER_3_3528 ();
 sg13g2_decap_8 FILLER_3_3535 ();
 sg13g2_decap_8 FILLER_3_3542 ();
 sg13g2_decap_8 FILLER_3_3549 ();
 sg13g2_decap_8 FILLER_3_3556 ();
 sg13g2_decap_8 FILLER_3_3563 ();
 sg13g2_decap_8 FILLER_3_3570 ();
 sg13g2_fill_2 FILLER_3_3577 ();
 sg13g2_fill_1 FILLER_3_3579 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_decap_8 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_4_868 ();
 sg13g2_decap_8 FILLER_4_875 ();
 sg13g2_decap_8 FILLER_4_882 ();
 sg13g2_decap_8 FILLER_4_889 ();
 sg13g2_decap_8 FILLER_4_896 ();
 sg13g2_decap_8 FILLER_4_903 ();
 sg13g2_decap_8 FILLER_4_910 ();
 sg13g2_decap_8 FILLER_4_917 ();
 sg13g2_decap_8 FILLER_4_924 ();
 sg13g2_decap_8 FILLER_4_931 ();
 sg13g2_decap_8 FILLER_4_938 ();
 sg13g2_decap_8 FILLER_4_945 ();
 sg13g2_decap_8 FILLER_4_952 ();
 sg13g2_decap_8 FILLER_4_959 ();
 sg13g2_decap_8 FILLER_4_966 ();
 sg13g2_decap_8 FILLER_4_973 ();
 sg13g2_decap_8 FILLER_4_980 ();
 sg13g2_decap_8 FILLER_4_987 ();
 sg13g2_decap_8 FILLER_4_994 ();
 sg13g2_decap_8 FILLER_4_1001 ();
 sg13g2_decap_8 FILLER_4_1008 ();
 sg13g2_decap_8 FILLER_4_1015 ();
 sg13g2_decap_8 FILLER_4_1022 ();
 sg13g2_decap_8 FILLER_4_1029 ();
 sg13g2_decap_8 FILLER_4_1036 ();
 sg13g2_decap_8 FILLER_4_1043 ();
 sg13g2_decap_8 FILLER_4_1050 ();
 sg13g2_decap_8 FILLER_4_1057 ();
 sg13g2_decap_8 FILLER_4_1064 ();
 sg13g2_decap_8 FILLER_4_1071 ();
 sg13g2_decap_8 FILLER_4_1078 ();
 sg13g2_decap_8 FILLER_4_1085 ();
 sg13g2_decap_8 FILLER_4_1092 ();
 sg13g2_decap_8 FILLER_4_1099 ();
 sg13g2_decap_8 FILLER_4_1106 ();
 sg13g2_decap_8 FILLER_4_1113 ();
 sg13g2_decap_8 FILLER_4_1120 ();
 sg13g2_decap_8 FILLER_4_1127 ();
 sg13g2_decap_8 FILLER_4_1134 ();
 sg13g2_decap_8 FILLER_4_1141 ();
 sg13g2_decap_8 FILLER_4_1148 ();
 sg13g2_decap_8 FILLER_4_1155 ();
 sg13g2_decap_8 FILLER_4_1162 ();
 sg13g2_decap_8 FILLER_4_1169 ();
 sg13g2_decap_8 FILLER_4_1176 ();
 sg13g2_decap_8 FILLER_4_1183 ();
 sg13g2_decap_8 FILLER_4_1190 ();
 sg13g2_decap_8 FILLER_4_1197 ();
 sg13g2_decap_8 FILLER_4_1204 ();
 sg13g2_decap_8 FILLER_4_1211 ();
 sg13g2_decap_8 FILLER_4_1218 ();
 sg13g2_decap_8 FILLER_4_1225 ();
 sg13g2_decap_8 FILLER_4_1232 ();
 sg13g2_decap_8 FILLER_4_1239 ();
 sg13g2_decap_8 FILLER_4_1246 ();
 sg13g2_decap_8 FILLER_4_1253 ();
 sg13g2_decap_8 FILLER_4_1260 ();
 sg13g2_decap_8 FILLER_4_1267 ();
 sg13g2_decap_8 FILLER_4_1274 ();
 sg13g2_decap_8 FILLER_4_1281 ();
 sg13g2_decap_8 FILLER_4_1288 ();
 sg13g2_decap_8 FILLER_4_1295 ();
 sg13g2_decap_8 FILLER_4_1302 ();
 sg13g2_decap_8 FILLER_4_1309 ();
 sg13g2_decap_8 FILLER_4_1316 ();
 sg13g2_decap_8 FILLER_4_1323 ();
 sg13g2_decap_8 FILLER_4_1330 ();
 sg13g2_decap_8 FILLER_4_1337 ();
 sg13g2_decap_8 FILLER_4_1344 ();
 sg13g2_decap_8 FILLER_4_1351 ();
 sg13g2_decap_8 FILLER_4_1358 ();
 sg13g2_decap_8 FILLER_4_1365 ();
 sg13g2_decap_8 FILLER_4_1372 ();
 sg13g2_decap_8 FILLER_4_1379 ();
 sg13g2_decap_8 FILLER_4_1386 ();
 sg13g2_decap_8 FILLER_4_1393 ();
 sg13g2_decap_8 FILLER_4_1400 ();
 sg13g2_decap_8 FILLER_4_1407 ();
 sg13g2_decap_8 FILLER_4_1414 ();
 sg13g2_decap_8 FILLER_4_1421 ();
 sg13g2_decap_8 FILLER_4_1428 ();
 sg13g2_decap_8 FILLER_4_1435 ();
 sg13g2_decap_8 FILLER_4_1442 ();
 sg13g2_decap_8 FILLER_4_1449 ();
 sg13g2_decap_8 FILLER_4_1456 ();
 sg13g2_decap_8 FILLER_4_1463 ();
 sg13g2_decap_8 FILLER_4_1470 ();
 sg13g2_decap_8 FILLER_4_1477 ();
 sg13g2_decap_8 FILLER_4_1484 ();
 sg13g2_decap_8 FILLER_4_1491 ();
 sg13g2_decap_8 FILLER_4_1498 ();
 sg13g2_decap_8 FILLER_4_1505 ();
 sg13g2_decap_8 FILLER_4_1512 ();
 sg13g2_decap_8 FILLER_4_1519 ();
 sg13g2_decap_8 FILLER_4_1526 ();
 sg13g2_decap_8 FILLER_4_1533 ();
 sg13g2_decap_8 FILLER_4_1540 ();
 sg13g2_decap_8 FILLER_4_1547 ();
 sg13g2_decap_8 FILLER_4_1554 ();
 sg13g2_decap_8 FILLER_4_1561 ();
 sg13g2_decap_8 FILLER_4_1568 ();
 sg13g2_decap_8 FILLER_4_1575 ();
 sg13g2_decap_8 FILLER_4_1582 ();
 sg13g2_decap_8 FILLER_4_1589 ();
 sg13g2_decap_8 FILLER_4_1596 ();
 sg13g2_decap_8 FILLER_4_1603 ();
 sg13g2_decap_8 FILLER_4_1610 ();
 sg13g2_decap_8 FILLER_4_1617 ();
 sg13g2_decap_8 FILLER_4_1624 ();
 sg13g2_decap_8 FILLER_4_1631 ();
 sg13g2_decap_8 FILLER_4_1638 ();
 sg13g2_decap_8 FILLER_4_1645 ();
 sg13g2_decap_8 FILLER_4_1652 ();
 sg13g2_decap_8 FILLER_4_1659 ();
 sg13g2_decap_8 FILLER_4_1666 ();
 sg13g2_decap_8 FILLER_4_1673 ();
 sg13g2_decap_8 FILLER_4_1680 ();
 sg13g2_decap_8 FILLER_4_1687 ();
 sg13g2_decap_8 FILLER_4_1694 ();
 sg13g2_decap_8 FILLER_4_1701 ();
 sg13g2_decap_8 FILLER_4_1708 ();
 sg13g2_decap_8 FILLER_4_1715 ();
 sg13g2_decap_8 FILLER_4_1722 ();
 sg13g2_decap_8 FILLER_4_1729 ();
 sg13g2_decap_8 FILLER_4_1736 ();
 sg13g2_decap_8 FILLER_4_1743 ();
 sg13g2_decap_8 FILLER_4_1750 ();
 sg13g2_decap_8 FILLER_4_1757 ();
 sg13g2_decap_8 FILLER_4_1764 ();
 sg13g2_decap_8 FILLER_4_1771 ();
 sg13g2_decap_8 FILLER_4_1778 ();
 sg13g2_decap_8 FILLER_4_1785 ();
 sg13g2_decap_8 FILLER_4_1792 ();
 sg13g2_decap_8 FILLER_4_1799 ();
 sg13g2_decap_8 FILLER_4_1806 ();
 sg13g2_decap_8 FILLER_4_1813 ();
 sg13g2_decap_8 FILLER_4_1820 ();
 sg13g2_decap_8 FILLER_4_1827 ();
 sg13g2_decap_8 FILLER_4_1834 ();
 sg13g2_decap_8 FILLER_4_1841 ();
 sg13g2_decap_8 FILLER_4_1848 ();
 sg13g2_decap_8 FILLER_4_1855 ();
 sg13g2_decap_8 FILLER_4_1862 ();
 sg13g2_decap_8 FILLER_4_1869 ();
 sg13g2_decap_8 FILLER_4_1876 ();
 sg13g2_decap_8 FILLER_4_1883 ();
 sg13g2_decap_8 FILLER_4_1890 ();
 sg13g2_decap_8 FILLER_4_1897 ();
 sg13g2_decap_8 FILLER_4_1904 ();
 sg13g2_decap_8 FILLER_4_1911 ();
 sg13g2_decap_8 FILLER_4_1918 ();
 sg13g2_decap_8 FILLER_4_1925 ();
 sg13g2_decap_8 FILLER_4_1932 ();
 sg13g2_decap_8 FILLER_4_1939 ();
 sg13g2_decap_8 FILLER_4_1946 ();
 sg13g2_decap_8 FILLER_4_1953 ();
 sg13g2_decap_8 FILLER_4_1960 ();
 sg13g2_decap_8 FILLER_4_1967 ();
 sg13g2_decap_8 FILLER_4_1974 ();
 sg13g2_decap_8 FILLER_4_1981 ();
 sg13g2_decap_8 FILLER_4_1988 ();
 sg13g2_decap_8 FILLER_4_1995 ();
 sg13g2_decap_8 FILLER_4_2002 ();
 sg13g2_decap_8 FILLER_4_2009 ();
 sg13g2_decap_8 FILLER_4_2016 ();
 sg13g2_decap_8 FILLER_4_2023 ();
 sg13g2_decap_8 FILLER_4_2030 ();
 sg13g2_decap_8 FILLER_4_2037 ();
 sg13g2_decap_8 FILLER_4_2044 ();
 sg13g2_decap_8 FILLER_4_2051 ();
 sg13g2_decap_8 FILLER_4_2058 ();
 sg13g2_decap_8 FILLER_4_2065 ();
 sg13g2_decap_8 FILLER_4_2072 ();
 sg13g2_decap_8 FILLER_4_2079 ();
 sg13g2_decap_8 FILLER_4_2086 ();
 sg13g2_decap_8 FILLER_4_2093 ();
 sg13g2_decap_8 FILLER_4_2100 ();
 sg13g2_decap_8 FILLER_4_2107 ();
 sg13g2_decap_8 FILLER_4_2114 ();
 sg13g2_decap_8 FILLER_4_2121 ();
 sg13g2_decap_8 FILLER_4_2128 ();
 sg13g2_decap_8 FILLER_4_2135 ();
 sg13g2_decap_8 FILLER_4_2142 ();
 sg13g2_decap_8 FILLER_4_2149 ();
 sg13g2_decap_8 FILLER_4_2156 ();
 sg13g2_decap_8 FILLER_4_2163 ();
 sg13g2_decap_8 FILLER_4_2170 ();
 sg13g2_decap_8 FILLER_4_2177 ();
 sg13g2_decap_8 FILLER_4_2184 ();
 sg13g2_decap_8 FILLER_4_2191 ();
 sg13g2_decap_8 FILLER_4_2198 ();
 sg13g2_decap_8 FILLER_4_2205 ();
 sg13g2_decap_8 FILLER_4_2212 ();
 sg13g2_decap_8 FILLER_4_2219 ();
 sg13g2_decap_8 FILLER_4_2226 ();
 sg13g2_decap_8 FILLER_4_2233 ();
 sg13g2_decap_8 FILLER_4_2240 ();
 sg13g2_decap_8 FILLER_4_2247 ();
 sg13g2_decap_8 FILLER_4_2254 ();
 sg13g2_decap_8 FILLER_4_2261 ();
 sg13g2_decap_8 FILLER_4_2268 ();
 sg13g2_decap_8 FILLER_4_2275 ();
 sg13g2_decap_8 FILLER_4_2282 ();
 sg13g2_decap_8 FILLER_4_2289 ();
 sg13g2_decap_8 FILLER_4_2296 ();
 sg13g2_decap_8 FILLER_4_2303 ();
 sg13g2_decap_8 FILLER_4_2310 ();
 sg13g2_decap_8 FILLER_4_2317 ();
 sg13g2_decap_8 FILLER_4_2324 ();
 sg13g2_decap_8 FILLER_4_2331 ();
 sg13g2_decap_8 FILLER_4_2338 ();
 sg13g2_decap_8 FILLER_4_2345 ();
 sg13g2_decap_8 FILLER_4_2352 ();
 sg13g2_decap_8 FILLER_4_2359 ();
 sg13g2_decap_8 FILLER_4_2366 ();
 sg13g2_decap_8 FILLER_4_2373 ();
 sg13g2_decap_8 FILLER_4_2380 ();
 sg13g2_decap_8 FILLER_4_2387 ();
 sg13g2_decap_8 FILLER_4_2394 ();
 sg13g2_decap_8 FILLER_4_2401 ();
 sg13g2_decap_8 FILLER_4_2408 ();
 sg13g2_decap_8 FILLER_4_2415 ();
 sg13g2_decap_8 FILLER_4_2422 ();
 sg13g2_decap_8 FILLER_4_2429 ();
 sg13g2_decap_8 FILLER_4_2436 ();
 sg13g2_decap_8 FILLER_4_2443 ();
 sg13g2_decap_8 FILLER_4_2450 ();
 sg13g2_decap_8 FILLER_4_2457 ();
 sg13g2_decap_8 FILLER_4_2464 ();
 sg13g2_decap_8 FILLER_4_2471 ();
 sg13g2_decap_8 FILLER_4_2478 ();
 sg13g2_decap_8 FILLER_4_2485 ();
 sg13g2_decap_8 FILLER_4_2492 ();
 sg13g2_decap_8 FILLER_4_2499 ();
 sg13g2_decap_8 FILLER_4_2506 ();
 sg13g2_decap_8 FILLER_4_2513 ();
 sg13g2_decap_8 FILLER_4_2520 ();
 sg13g2_decap_8 FILLER_4_2527 ();
 sg13g2_decap_8 FILLER_4_2534 ();
 sg13g2_decap_8 FILLER_4_2541 ();
 sg13g2_decap_8 FILLER_4_2548 ();
 sg13g2_decap_8 FILLER_4_2555 ();
 sg13g2_decap_8 FILLER_4_2562 ();
 sg13g2_decap_8 FILLER_4_2569 ();
 sg13g2_decap_8 FILLER_4_2576 ();
 sg13g2_decap_8 FILLER_4_2583 ();
 sg13g2_decap_8 FILLER_4_2590 ();
 sg13g2_decap_8 FILLER_4_2597 ();
 sg13g2_decap_8 FILLER_4_2604 ();
 sg13g2_decap_8 FILLER_4_2611 ();
 sg13g2_decap_8 FILLER_4_2618 ();
 sg13g2_decap_8 FILLER_4_2625 ();
 sg13g2_decap_8 FILLER_4_2632 ();
 sg13g2_decap_8 FILLER_4_2639 ();
 sg13g2_decap_8 FILLER_4_2646 ();
 sg13g2_decap_8 FILLER_4_2653 ();
 sg13g2_decap_8 FILLER_4_2660 ();
 sg13g2_decap_8 FILLER_4_2667 ();
 sg13g2_decap_8 FILLER_4_2674 ();
 sg13g2_decap_8 FILLER_4_2681 ();
 sg13g2_decap_8 FILLER_4_2688 ();
 sg13g2_decap_8 FILLER_4_2695 ();
 sg13g2_decap_8 FILLER_4_2702 ();
 sg13g2_decap_8 FILLER_4_2709 ();
 sg13g2_decap_8 FILLER_4_2716 ();
 sg13g2_decap_8 FILLER_4_2723 ();
 sg13g2_decap_8 FILLER_4_2730 ();
 sg13g2_decap_8 FILLER_4_2737 ();
 sg13g2_decap_8 FILLER_4_2744 ();
 sg13g2_decap_8 FILLER_4_2751 ();
 sg13g2_decap_8 FILLER_4_2758 ();
 sg13g2_decap_8 FILLER_4_2765 ();
 sg13g2_decap_8 FILLER_4_2772 ();
 sg13g2_decap_8 FILLER_4_2779 ();
 sg13g2_decap_8 FILLER_4_2786 ();
 sg13g2_decap_8 FILLER_4_2793 ();
 sg13g2_decap_8 FILLER_4_2800 ();
 sg13g2_decap_8 FILLER_4_2807 ();
 sg13g2_decap_8 FILLER_4_2814 ();
 sg13g2_decap_8 FILLER_4_2821 ();
 sg13g2_decap_8 FILLER_4_2828 ();
 sg13g2_decap_8 FILLER_4_2835 ();
 sg13g2_decap_8 FILLER_4_2842 ();
 sg13g2_decap_8 FILLER_4_2849 ();
 sg13g2_decap_8 FILLER_4_2856 ();
 sg13g2_decap_8 FILLER_4_2863 ();
 sg13g2_decap_8 FILLER_4_2870 ();
 sg13g2_decap_8 FILLER_4_2877 ();
 sg13g2_decap_8 FILLER_4_2884 ();
 sg13g2_decap_8 FILLER_4_2891 ();
 sg13g2_decap_8 FILLER_4_2898 ();
 sg13g2_decap_8 FILLER_4_2905 ();
 sg13g2_decap_8 FILLER_4_2912 ();
 sg13g2_decap_8 FILLER_4_2919 ();
 sg13g2_decap_8 FILLER_4_2926 ();
 sg13g2_decap_8 FILLER_4_2933 ();
 sg13g2_decap_8 FILLER_4_2940 ();
 sg13g2_decap_8 FILLER_4_2947 ();
 sg13g2_decap_8 FILLER_4_2954 ();
 sg13g2_decap_8 FILLER_4_2961 ();
 sg13g2_decap_8 FILLER_4_2968 ();
 sg13g2_decap_8 FILLER_4_2975 ();
 sg13g2_decap_8 FILLER_4_2982 ();
 sg13g2_decap_8 FILLER_4_2989 ();
 sg13g2_decap_8 FILLER_4_2996 ();
 sg13g2_decap_8 FILLER_4_3003 ();
 sg13g2_decap_8 FILLER_4_3010 ();
 sg13g2_decap_8 FILLER_4_3017 ();
 sg13g2_decap_8 FILLER_4_3024 ();
 sg13g2_decap_8 FILLER_4_3031 ();
 sg13g2_decap_8 FILLER_4_3038 ();
 sg13g2_decap_8 FILLER_4_3045 ();
 sg13g2_decap_8 FILLER_4_3052 ();
 sg13g2_decap_8 FILLER_4_3059 ();
 sg13g2_decap_8 FILLER_4_3066 ();
 sg13g2_decap_8 FILLER_4_3073 ();
 sg13g2_decap_8 FILLER_4_3080 ();
 sg13g2_decap_8 FILLER_4_3087 ();
 sg13g2_decap_8 FILLER_4_3094 ();
 sg13g2_decap_8 FILLER_4_3101 ();
 sg13g2_decap_8 FILLER_4_3108 ();
 sg13g2_decap_8 FILLER_4_3115 ();
 sg13g2_decap_8 FILLER_4_3122 ();
 sg13g2_decap_8 FILLER_4_3129 ();
 sg13g2_decap_8 FILLER_4_3136 ();
 sg13g2_decap_8 FILLER_4_3143 ();
 sg13g2_decap_8 FILLER_4_3150 ();
 sg13g2_decap_8 FILLER_4_3157 ();
 sg13g2_decap_8 FILLER_4_3164 ();
 sg13g2_decap_8 FILLER_4_3171 ();
 sg13g2_decap_8 FILLER_4_3178 ();
 sg13g2_decap_8 FILLER_4_3185 ();
 sg13g2_decap_8 FILLER_4_3192 ();
 sg13g2_decap_8 FILLER_4_3199 ();
 sg13g2_decap_8 FILLER_4_3206 ();
 sg13g2_decap_8 FILLER_4_3213 ();
 sg13g2_decap_8 FILLER_4_3220 ();
 sg13g2_decap_8 FILLER_4_3227 ();
 sg13g2_decap_8 FILLER_4_3234 ();
 sg13g2_decap_8 FILLER_4_3241 ();
 sg13g2_decap_8 FILLER_4_3248 ();
 sg13g2_decap_8 FILLER_4_3255 ();
 sg13g2_decap_8 FILLER_4_3262 ();
 sg13g2_decap_8 FILLER_4_3269 ();
 sg13g2_decap_8 FILLER_4_3276 ();
 sg13g2_decap_8 FILLER_4_3283 ();
 sg13g2_decap_8 FILLER_4_3290 ();
 sg13g2_decap_8 FILLER_4_3297 ();
 sg13g2_decap_8 FILLER_4_3304 ();
 sg13g2_decap_8 FILLER_4_3311 ();
 sg13g2_decap_8 FILLER_4_3318 ();
 sg13g2_decap_8 FILLER_4_3325 ();
 sg13g2_decap_8 FILLER_4_3332 ();
 sg13g2_decap_8 FILLER_4_3339 ();
 sg13g2_decap_8 FILLER_4_3346 ();
 sg13g2_decap_8 FILLER_4_3353 ();
 sg13g2_decap_8 FILLER_4_3360 ();
 sg13g2_decap_8 FILLER_4_3367 ();
 sg13g2_decap_8 FILLER_4_3374 ();
 sg13g2_decap_8 FILLER_4_3381 ();
 sg13g2_decap_8 FILLER_4_3388 ();
 sg13g2_decap_8 FILLER_4_3395 ();
 sg13g2_decap_8 FILLER_4_3402 ();
 sg13g2_decap_8 FILLER_4_3409 ();
 sg13g2_decap_8 FILLER_4_3416 ();
 sg13g2_decap_8 FILLER_4_3423 ();
 sg13g2_decap_8 FILLER_4_3430 ();
 sg13g2_decap_8 FILLER_4_3437 ();
 sg13g2_decap_8 FILLER_4_3444 ();
 sg13g2_decap_8 FILLER_4_3451 ();
 sg13g2_decap_8 FILLER_4_3458 ();
 sg13g2_decap_8 FILLER_4_3465 ();
 sg13g2_decap_8 FILLER_4_3472 ();
 sg13g2_decap_8 FILLER_4_3479 ();
 sg13g2_decap_8 FILLER_4_3486 ();
 sg13g2_decap_8 FILLER_4_3493 ();
 sg13g2_decap_8 FILLER_4_3500 ();
 sg13g2_decap_8 FILLER_4_3507 ();
 sg13g2_decap_8 FILLER_4_3514 ();
 sg13g2_decap_8 FILLER_4_3521 ();
 sg13g2_decap_8 FILLER_4_3528 ();
 sg13g2_decap_8 FILLER_4_3535 ();
 sg13g2_decap_8 FILLER_4_3542 ();
 sg13g2_decap_8 FILLER_4_3549 ();
 sg13g2_decap_8 FILLER_4_3556 ();
 sg13g2_decap_8 FILLER_4_3563 ();
 sg13g2_decap_8 FILLER_4_3570 ();
 sg13g2_fill_2 FILLER_4_3577 ();
 sg13g2_fill_1 FILLER_4_3579 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_decap_8 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_5_868 ();
 sg13g2_decap_8 FILLER_5_875 ();
 sg13g2_decap_8 FILLER_5_882 ();
 sg13g2_decap_8 FILLER_5_889 ();
 sg13g2_decap_8 FILLER_5_896 ();
 sg13g2_decap_8 FILLER_5_903 ();
 sg13g2_decap_8 FILLER_5_910 ();
 sg13g2_decap_8 FILLER_5_917 ();
 sg13g2_decap_8 FILLER_5_924 ();
 sg13g2_decap_8 FILLER_5_931 ();
 sg13g2_decap_8 FILLER_5_938 ();
 sg13g2_decap_8 FILLER_5_945 ();
 sg13g2_decap_8 FILLER_5_952 ();
 sg13g2_decap_8 FILLER_5_959 ();
 sg13g2_decap_8 FILLER_5_966 ();
 sg13g2_decap_8 FILLER_5_973 ();
 sg13g2_decap_8 FILLER_5_980 ();
 sg13g2_decap_8 FILLER_5_987 ();
 sg13g2_decap_8 FILLER_5_994 ();
 sg13g2_decap_8 FILLER_5_1001 ();
 sg13g2_decap_8 FILLER_5_1008 ();
 sg13g2_decap_8 FILLER_5_1015 ();
 sg13g2_decap_8 FILLER_5_1022 ();
 sg13g2_decap_8 FILLER_5_1029 ();
 sg13g2_decap_8 FILLER_5_1036 ();
 sg13g2_decap_8 FILLER_5_1043 ();
 sg13g2_decap_8 FILLER_5_1050 ();
 sg13g2_decap_8 FILLER_5_1057 ();
 sg13g2_decap_8 FILLER_5_1064 ();
 sg13g2_decap_8 FILLER_5_1071 ();
 sg13g2_decap_8 FILLER_5_1078 ();
 sg13g2_decap_8 FILLER_5_1085 ();
 sg13g2_decap_8 FILLER_5_1092 ();
 sg13g2_decap_8 FILLER_5_1099 ();
 sg13g2_decap_8 FILLER_5_1106 ();
 sg13g2_decap_8 FILLER_5_1113 ();
 sg13g2_decap_8 FILLER_5_1120 ();
 sg13g2_decap_8 FILLER_5_1127 ();
 sg13g2_decap_8 FILLER_5_1134 ();
 sg13g2_decap_8 FILLER_5_1141 ();
 sg13g2_decap_8 FILLER_5_1148 ();
 sg13g2_decap_8 FILLER_5_1155 ();
 sg13g2_decap_8 FILLER_5_1162 ();
 sg13g2_decap_8 FILLER_5_1169 ();
 sg13g2_decap_8 FILLER_5_1176 ();
 sg13g2_decap_8 FILLER_5_1183 ();
 sg13g2_decap_8 FILLER_5_1190 ();
 sg13g2_decap_8 FILLER_5_1197 ();
 sg13g2_decap_8 FILLER_5_1204 ();
 sg13g2_decap_8 FILLER_5_1211 ();
 sg13g2_decap_8 FILLER_5_1218 ();
 sg13g2_decap_8 FILLER_5_1225 ();
 sg13g2_decap_8 FILLER_5_1232 ();
 sg13g2_decap_8 FILLER_5_1239 ();
 sg13g2_decap_8 FILLER_5_1246 ();
 sg13g2_decap_8 FILLER_5_1253 ();
 sg13g2_decap_8 FILLER_5_1260 ();
 sg13g2_decap_8 FILLER_5_1267 ();
 sg13g2_decap_8 FILLER_5_1274 ();
 sg13g2_decap_8 FILLER_5_1281 ();
 sg13g2_decap_8 FILLER_5_1288 ();
 sg13g2_decap_8 FILLER_5_1295 ();
 sg13g2_decap_8 FILLER_5_1302 ();
 sg13g2_decap_8 FILLER_5_1309 ();
 sg13g2_decap_8 FILLER_5_1316 ();
 sg13g2_decap_8 FILLER_5_1323 ();
 sg13g2_decap_8 FILLER_5_1330 ();
 sg13g2_decap_8 FILLER_5_1337 ();
 sg13g2_decap_8 FILLER_5_1344 ();
 sg13g2_decap_8 FILLER_5_1351 ();
 sg13g2_decap_8 FILLER_5_1358 ();
 sg13g2_decap_8 FILLER_5_1365 ();
 sg13g2_decap_8 FILLER_5_1372 ();
 sg13g2_decap_8 FILLER_5_1379 ();
 sg13g2_decap_8 FILLER_5_1386 ();
 sg13g2_decap_8 FILLER_5_1393 ();
 sg13g2_decap_8 FILLER_5_1400 ();
 sg13g2_decap_8 FILLER_5_1407 ();
 sg13g2_decap_8 FILLER_5_1414 ();
 sg13g2_decap_8 FILLER_5_1421 ();
 sg13g2_decap_8 FILLER_5_1428 ();
 sg13g2_decap_8 FILLER_5_1435 ();
 sg13g2_decap_8 FILLER_5_1442 ();
 sg13g2_decap_8 FILLER_5_1449 ();
 sg13g2_decap_8 FILLER_5_1456 ();
 sg13g2_decap_8 FILLER_5_1463 ();
 sg13g2_decap_8 FILLER_5_1470 ();
 sg13g2_decap_8 FILLER_5_1477 ();
 sg13g2_decap_8 FILLER_5_1484 ();
 sg13g2_decap_8 FILLER_5_1491 ();
 sg13g2_decap_8 FILLER_5_1498 ();
 sg13g2_decap_8 FILLER_5_1505 ();
 sg13g2_decap_8 FILLER_5_1512 ();
 sg13g2_decap_8 FILLER_5_1519 ();
 sg13g2_decap_8 FILLER_5_1526 ();
 sg13g2_decap_8 FILLER_5_1533 ();
 sg13g2_decap_8 FILLER_5_1540 ();
 sg13g2_decap_8 FILLER_5_1547 ();
 sg13g2_decap_8 FILLER_5_1554 ();
 sg13g2_decap_8 FILLER_5_1561 ();
 sg13g2_decap_8 FILLER_5_1568 ();
 sg13g2_decap_8 FILLER_5_1575 ();
 sg13g2_decap_8 FILLER_5_1582 ();
 sg13g2_decap_8 FILLER_5_1589 ();
 sg13g2_decap_8 FILLER_5_1596 ();
 sg13g2_decap_8 FILLER_5_1603 ();
 sg13g2_decap_8 FILLER_5_1610 ();
 sg13g2_decap_8 FILLER_5_1617 ();
 sg13g2_decap_8 FILLER_5_1624 ();
 sg13g2_decap_8 FILLER_5_1631 ();
 sg13g2_decap_8 FILLER_5_1638 ();
 sg13g2_decap_8 FILLER_5_1645 ();
 sg13g2_decap_8 FILLER_5_1652 ();
 sg13g2_decap_8 FILLER_5_1659 ();
 sg13g2_decap_8 FILLER_5_1666 ();
 sg13g2_decap_8 FILLER_5_1673 ();
 sg13g2_decap_8 FILLER_5_1680 ();
 sg13g2_decap_8 FILLER_5_1687 ();
 sg13g2_decap_8 FILLER_5_1694 ();
 sg13g2_decap_8 FILLER_5_1701 ();
 sg13g2_decap_8 FILLER_5_1708 ();
 sg13g2_decap_8 FILLER_5_1715 ();
 sg13g2_decap_8 FILLER_5_1722 ();
 sg13g2_decap_8 FILLER_5_1729 ();
 sg13g2_decap_8 FILLER_5_1736 ();
 sg13g2_decap_8 FILLER_5_1743 ();
 sg13g2_decap_8 FILLER_5_1750 ();
 sg13g2_decap_8 FILLER_5_1757 ();
 sg13g2_decap_8 FILLER_5_1764 ();
 sg13g2_decap_8 FILLER_5_1771 ();
 sg13g2_decap_8 FILLER_5_1778 ();
 sg13g2_decap_8 FILLER_5_1785 ();
 sg13g2_decap_8 FILLER_5_1792 ();
 sg13g2_decap_8 FILLER_5_1799 ();
 sg13g2_decap_8 FILLER_5_1806 ();
 sg13g2_decap_8 FILLER_5_1813 ();
 sg13g2_decap_8 FILLER_5_1820 ();
 sg13g2_decap_8 FILLER_5_1827 ();
 sg13g2_decap_8 FILLER_5_1834 ();
 sg13g2_decap_8 FILLER_5_1841 ();
 sg13g2_decap_8 FILLER_5_1848 ();
 sg13g2_decap_8 FILLER_5_1855 ();
 sg13g2_decap_8 FILLER_5_1862 ();
 sg13g2_decap_8 FILLER_5_1869 ();
 sg13g2_decap_8 FILLER_5_1876 ();
 sg13g2_decap_8 FILLER_5_1883 ();
 sg13g2_decap_8 FILLER_5_1890 ();
 sg13g2_decap_8 FILLER_5_1897 ();
 sg13g2_decap_8 FILLER_5_1904 ();
 sg13g2_decap_8 FILLER_5_1911 ();
 sg13g2_decap_8 FILLER_5_1918 ();
 sg13g2_decap_8 FILLER_5_1925 ();
 sg13g2_decap_8 FILLER_5_1932 ();
 sg13g2_decap_8 FILLER_5_1939 ();
 sg13g2_decap_8 FILLER_5_1946 ();
 sg13g2_decap_8 FILLER_5_1953 ();
 sg13g2_decap_8 FILLER_5_1960 ();
 sg13g2_decap_8 FILLER_5_1967 ();
 sg13g2_decap_8 FILLER_5_1974 ();
 sg13g2_decap_8 FILLER_5_1981 ();
 sg13g2_decap_8 FILLER_5_1988 ();
 sg13g2_decap_8 FILLER_5_1995 ();
 sg13g2_decap_8 FILLER_5_2002 ();
 sg13g2_decap_8 FILLER_5_2009 ();
 sg13g2_decap_8 FILLER_5_2016 ();
 sg13g2_decap_8 FILLER_5_2023 ();
 sg13g2_decap_8 FILLER_5_2030 ();
 sg13g2_decap_8 FILLER_5_2037 ();
 sg13g2_decap_8 FILLER_5_2044 ();
 sg13g2_decap_8 FILLER_5_2051 ();
 sg13g2_decap_8 FILLER_5_2058 ();
 sg13g2_decap_8 FILLER_5_2065 ();
 sg13g2_decap_8 FILLER_5_2072 ();
 sg13g2_decap_8 FILLER_5_2079 ();
 sg13g2_decap_8 FILLER_5_2086 ();
 sg13g2_decap_8 FILLER_5_2093 ();
 sg13g2_decap_8 FILLER_5_2100 ();
 sg13g2_decap_8 FILLER_5_2107 ();
 sg13g2_decap_8 FILLER_5_2114 ();
 sg13g2_decap_8 FILLER_5_2121 ();
 sg13g2_decap_8 FILLER_5_2128 ();
 sg13g2_decap_8 FILLER_5_2135 ();
 sg13g2_decap_8 FILLER_5_2142 ();
 sg13g2_decap_8 FILLER_5_2149 ();
 sg13g2_decap_8 FILLER_5_2156 ();
 sg13g2_decap_8 FILLER_5_2163 ();
 sg13g2_decap_8 FILLER_5_2170 ();
 sg13g2_decap_8 FILLER_5_2177 ();
 sg13g2_decap_8 FILLER_5_2184 ();
 sg13g2_decap_8 FILLER_5_2191 ();
 sg13g2_decap_8 FILLER_5_2198 ();
 sg13g2_decap_8 FILLER_5_2205 ();
 sg13g2_decap_8 FILLER_5_2212 ();
 sg13g2_decap_8 FILLER_5_2219 ();
 sg13g2_decap_8 FILLER_5_2226 ();
 sg13g2_decap_8 FILLER_5_2233 ();
 sg13g2_decap_8 FILLER_5_2240 ();
 sg13g2_decap_8 FILLER_5_2247 ();
 sg13g2_decap_8 FILLER_5_2254 ();
 sg13g2_decap_8 FILLER_5_2261 ();
 sg13g2_decap_8 FILLER_5_2268 ();
 sg13g2_decap_8 FILLER_5_2275 ();
 sg13g2_decap_8 FILLER_5_2282 ();
 sg13g2_decap_8 FILLER_5_2289 ();
 sg13g2_decap_8 FILLER_5_2296 ();
 sg13g2_decap_8 FILLER_5_2303 ();
 sg13g2_decap_8 FILLER_5_2310 ();
 sg13g2_decap_8 FILLER_5_2317 ();
 sg13g2_decap_8 FILLER_5_2324 ();
 sg13g2_decap_8 FILLER_5_2331 ();
 sg13g2_decap_8 FILLER_5_2338 ();
 sg13g2_decap_8 FILLER_5_2345 ();
 sg13g2_decap_8 FILLER_5_2352 ();
 sg13g2_decap_8 FILLER_5_2359 ();
 sg13g2_decap_8 FILLER_5_2366 ();
 sg13g2_decap_8 FILLER_5_2373 ();
 sg13g2_decap_8 FILLER_5_2380 ();
 sg13g2_decap_8 FILLER_5_2387 ();
 sg13g2_decap_8 FILLER_5_2394 ();
 sg13g2_decap_8 FILLER_5_2401 ();
 sg13g2_decap_8 FILLER_5_2408 ();
 sg13g2_decap_8 FILLER_5_2415 ();
 sg13g2_decap_8 FILLER_5_2422 ();
 sg13g2_decap_8 FILLER_5_2429 ();
 sg13g2_decap_8 FILLER_5_2436 ();
 sg13g2_decap_8 FILLER_5_2443 ();
 sg13g2_decap_8 FILLER_5_2450 ();
 sg13g2_decap_8 FILLER_5_2457 ();
 sg13g2_decap_8 FILLER_5_2464 ();
 sg13g2_decap_8 FILLER_5_2471 ();
 sg13g2_decap_8 FILLER_5_2478 ();
 sg13g2_decap_8 FILLER_5_2485 ();
 sg13g2_decap_8 FILLER_5_2492 ();
 sg13g2_decap_8 FILLER_5_2499 ();
 sg13g2_decap_8 FILLER_5_2506 ();
 sg13g2_decap_8 FILLER_5_2513 ();
 sg13g2_decap_8 FILLER_5_2520 ();
 sg13g2_decap_8 FILLER_5_2527 ();
 sg13g2_decap_8 FILLER_5_2534 ();
 sg13g2_decap_8 FILLER_5_2541 ();
 sg13g2_decap_8 FILLER_5_2548 ();
 sg13g2_decap_8 FILLER_5_2555 ();
 sg13g2_decap_8 FILLER_5_2562 ();
 sg13g2_decap_8 FILLER_5_2569 ();
 sg13g2_decap_8 FILLER_5_2576 ();
 sg13g2_decap_8 FILLER_5_2583 ();
 sg13g2_decap_8 FILLER_5_2590 ();
 sg13g2_decap_8 FILLER_5_2597 ();
 sg13g2_decap_8 FILLER_5_2604 ();
 sg13g2_decap_8 FILLER_5_2611 ();
 sg13g2_decap_8 FILLER_5_2618 ();
 sg13g2_decap_8 FILLER_5_2625 ();
 sg13g2_decap_8 FILLER_5_2632 ();
 sg13g2_decap_8 FILLER_5_2639 ();
 sg13g2_decap_8 FILLER_5_2646 ();
 sg13g2_decap_8 FILLER_5_2653 ();
 sg13g2_decap_8 FILLER_5_2660 ();
 sg13g2_decap_8 FILLER_5_2667 ();
 sg13g2_decap_8 FILLER_5_2674 ();
 sg13g2_decap_8 FILLER_5_2681 ();
 sg13g2_decap_8 FILLER_5_2688 ();
 sg13g2_decap_8 FILLER_5_2695 ();
 sg13g2_decap_8 FILLER_5_2702 ();
 sg13g2_decap_8 FILLER_5_2709 ();
 sg13g2_decap_8 FILLER_5_2716 ();
 sg13g2_decap_8 FILLER_5_2723 ();
 sg13g2_decap_8 FILLER_5_2730 ();
 sg13g2_decap_8 FILLER_5_2737 ();
 sg13g2_decap_8 FILLER_5_2744 ();
 sg13g2_decap_8 FILLER_5_2751 ();
 sg13g2_decap_8 FILLER_5_2758 ();
 sg13g2_decap_8 FILLER_5_2765 ();
 sg13g2_decap_8 FILLER_5_2772 ();
 sg13g2_decap_8 FILLER_5_2779 ();
 sg13g2_decap_8 FILLER_5_2786 ();
 sg13g2_decap_8 FILLER_5_2793 ();
 sg13g2_decap_8 FILLER_5_2800 ();
 sg13g2_decap_8 FILLER_5_2807 ();
 sg13g2_decap_8 FILLER_5_2814 ();
 sg13g2_decap_8 FILLER_5_2821 ();
 sg13g2_decap_8 FILLER_5_2828 ();
 sg13g2_decap_8 FILLER_5_2835 ();
 sg13g2_decap_8 FILLER_5_2842 ();
 sg13g2_decap_8 FILLER_5_2849 ();
 sg13g2_decap_8 FILLER_5_2856 ();
 sg13g2_decap_8 FILLER_5_2863 ();
 sg13g2_decap_8 FILLER_5_2870 ();
 sg13g2_decap_8 FILLER_5_2877 ();
 sg13g2_decap_8 FILLER_5_2884 ();
 sg13g2_decap_8 FILLER_5_2891 ();
 sg13g2_decap_8 FILLER_5_2898 ();
 sg13g2_decap_8 FILLER_5_2905 ();
 sg13g2_decap_8 FILLER_5_2912 ();
 sg13g2_decap_8 FILLER_5_2919 ();
 sg13g2_decap_8 FILLER_5_2926 ();
 sg13g2_decap_8 FILLER_5_2933 ();
 sg13g2_decap_8 FILLER_5_2940 ();
 sg13g2_decap_8 FILLER_5_2947 ();
 sg13g2_decap_8 FILLER_5_2954 ();
 sg13g2_decap_8 FILLER_5_2961 ();
 sg13g2_decap_8 FILLER_5_2968 ();
 sg13g2_decap_8 FILLER_5_2975 ();
 sg13g2_decap_8 FILLER_5_2982 ();
 sg13g2_decap_8 FILLER_5_2989 ();
 sg13g2_decap_8 FILLER_5_2996 ();
 sg13g2_decap_8 FILLER_5_3003 ();
 sg13g2_decap_8 FILLER_5_3010 ();
 sg13g2_decap_8 FILLER_5_3017 ();
 sg13g2_decap_8 FILLER_5_3024 ();
 sg13g2_decap_8 FILLER_5_3031 ();
 sg13g2_decap_8 FILLER_5_3038 ();
 sg13g2_decap_8 FILLER_5_3045 ();
 sg13g2_decap_8 FILLER_5_3052 ();
 sg13g2_decap_8 FILLER_5_3059 ();
 sg13g2_decap_8 FILLER_5_3066 ();
 sg13g2_decap_8 FILLER_5_3073 ();
 sg13g2_decap_8 FILLER_5_3080 ();
 sg13g2_decap_8 FILLER_5_3087 ();
 sg13g2_decap_8 FILLER_5_3094 ();
 sg13g2_decap_8 FILLER_5_3101 ();
 sg13g2_decap_8 FILLER_5_3108 ();
 sg13g2_decap_8 FILLER_5_3115 ();
 sg13g2_decap_8 FILLER_5_3122 ();
 sg13g2_decap_8 FILLER_5_3129 ();
 sg13g2_decap_8 FILLER_5_3136 ();
 sg13g2_decap_8 FILLER_5_3143 ();
 sg13g2_decap_8 FILLER_5_3150 ();
 sg13g2_decap_8 FILLER_5_3157 ();
 sg13g2_decap_8 FILLER_5_3164 ();
 sg13g2_decap_8 FILLER_5_3171 ();
 sg13g2_decap_8 FILLER_5_3178 ();
 sg13g2_decap_8 FILLER_5_3185 ();
 sg13g2_decap_8 FILLER_5_3192 ();
 sg13g2_decap_8 FILLER_5_3199 ();
 sg13g2_decap_8 FILLER_5_3206 ();
 sg13g2_decap_8 FILLER_5_3213 ();
 sg13g2_decap_8 FILLER_5_3220 ();
 sg13g2_decap_8 FILLER_5_3227 ();
 sg13g2_decap_8 FILLER_5_3234 ();
 sg13g2_decap_8 FILLER_5_3241 ();
 sg13g2_decap_8 FILLER_5_3248 ();
 sg13g2_decap_8 FILLER_5_3255 ();
 sg13g2_decap_8 FILLER_5_3262 ();
 sg13g2_decap_8 FILLER_5_3269 ();
 sg13g2_decap_8 FILLER_5_3276 ();
 sg13g2_decap_8 FILLER_5_3283 ();
 sg13g2_decap_8 FILLER_5_3290 ();
 sg13g2_decap_8 FILLER_5_3297 ();
 sg13g2_decap_8 FILLER_5_3304 ();
 sg13g2_decap_8 FILLER_5_3311 ();
 sg13g2_decap_8 FILLER_5_3318 ();
 sg13g2_decap_8 FILLER_5_3325 ();
 sg13g2_decap_8 FILLER_5_3332 ();
 sg13g2_decap_8 FILLER_5_3339 ();
 sg13g2_decap_8 FILLER_5_3346 ();
 sg13g2_decap_8 FILLER_5_3353 ();
 sg13g2_decap_8 FILLER_5_3360 ();
 sg13g2_decap_8 FILLER_5_3367 ();
 sg13g2_decap_8 FILLER_5_3374 ();
 sg13g2_decap_8 FILLER_5_3381 ();
 sg13g2_decap_8 FILLER_5_3388 ();
 sg13g2_decap_8 FILLER_5_3395 ();
 sg13g2_decap_8 FILLER_5_3402 ();
 sg13g2_decap_8 FILLER_5_3409 ();
 sg13g2_decap_8 FILLER_5_3416 ();
 sg13g2_decap_8 FILLER_5_3423 ();
 sg13g2_decap_8 FILLER_5_3430 ();
 sg13g2_decap_8 FILLER_5_3437 ();
 sg13g2_decap_8 FILLER_5_3444 ();
 sg13g2_decap_8 FILLER_5_3451 ();
 sg13g2_decap_8 FILLER_5_3458 ();
 sg13g2_decap_8 FILLER_5_3465 ();
 sg13g2_decap_8 FILLER_5_3472 ();
 sg13g2_decap_8 FILLER_5_3479 ();
 sg13g2_decap_8 FILLER_5_3486 ();
 sg13g2_decap_8 FILLER_5_3493 ();
 sg13g2_decap_8 FILLER_5_3500 ();
 sg13g2_decap_8 FILLER_5_3507 ();
 sg13g2_decap_8 FILLER_5_3514 ();
 sg13g2_decap_8 FILLER_5_3521 ();
 sg13g2_decap_8 FILLER_5_3528 ();
 sg13g2_decap_8 FILLER_5_3535 ();
 sg13g2_decap_8 FILLER_5_3542 ();
 sg13g2_decap_8 FILLER_5_3549 ();
 sg13g2_decap_8 FILLER_5_3556 ();
 sg13g2_decap_8 FILLER_5_3563 ();
 sg13g2_decap_8 FILLER_5_3570 ();
 sg13g2_fill_2 FILLER_5_3577 ();
 sg13g2_fill_1 FILLER_5_3579 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_decap_8 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_6_868 ();
 sg13g2_decap_8 FILLER_6_875 ();
 sg13g2_decap_8 FILLER_6_882 ();
 sg13g2_decap_8 FILLER_6_889 ();
 sg13g2_decap_8 FILLER_6_896 ();
 sg13g2_decap_8 FILLER_6_903 ();
 sg13g2_decap_8 FILLER_6_910 ();
 sg13g2_decap_8 FILLER_6_917 ();
 sg13g2_decap_8 FILLER_6_924 ();
 sg13g2_decap_8 FILLER_6_931 ();
 sg13g2_decap_8 FILLER_6_938 ();
 sg13g2_decap_8 FILLER_6_945 ();
 sg13g2_decap_8 FILLER_6_952 ();
 sg13g2_decap_8 FILLER_6_959 ();
 sg13g2_decap_8 FILLER_6_966 ();
 sg13g2_decap_8 FILLER_6_973 ();
 sg13g2_decap_8 FILLER_6_980 ();
 sg13g2_decap_8 FILLER_6_987 ();
 sg13g2_decap_8 FILLER_6_994 ();
 sg13g2_decap_8 FILLER_6_1001 ();
 sg13g2_decap_8 FILLER_6_1008 ();
 sg13g2_decap_8 FILLER_6_1015 ();
 sg13g2_decap_8 FILLER_6_1022 ();
 sg13g2_decap_8 FILLER_6_1029 ();
 sg13g2_decap_8 FILLER_6_1036 ();
 sg13g2_decap_8 FILLER_6_1043 ();
 sg13g2_decap_8 FILLER_6_1050 ();
 sg13g2_decap_8 FILLER_6_1057 ();
 sg13g2_decap_8 FILLER_6_1064 ();
 sg13g2_decap_8 FILLER_6_1071 ();
 sg13g2_decap_8 FILLER_6_1078 ();
 sg13g2_decap_8 FILLER_6_1085 ();
 sg13g2_decap_8 FILLER_6_1092 ();
 sg13g2_decap_8 FILLER_6_1099 ();
 sg13g2_decap_8 FILLER_6_1106 ();
 sg13g2_decap_8 FILLER_6_1113 ();
 sg13g2_decap_8 FILLER_6_1120 ();
 sg13g2_decap_8 FILLER_6_1127 ();
 sg13g2_decap_8 FILLER_6_1134 ();
 sg13g2_decap_8 FILLER_6_1141 ();
 sg13g2_decap_8 FILLER_6_1148 ();
 sg13g2_decap_8 FILLER_6_1155 ();
 sg13g2_decap_8 FILLER_6_1162 ();
 sg13g2_decap_8 FILLER_6_1169 ();
 sg13g2_decap_8 FILLER_6_1176 ();
 sg13g2_decap_8 FILLER_6_1183 ();
 sg13g2_decap_8 FILLER_6_1190 ();
 sg13g2_decap_8 FILLER_6_1197 ();
 sg13g2_decap_8 FILLER_6_1204 ();
 sg13g2_decap_8 FILLER_6_1211 ();
 sg13g2_decap_8 FILLER_6_1218 ();
 sg13g2_decap_8 FILLER_6_1225 ();
 sg13g2_decap_8 FILLER_6_1232 ();
 sg13g2_decap_8 FILLER_6_1239 ();
 sg13g2_decap_8 FILLER_6_1246 ();
 sg13g2_decap_8 FILLER_6_1253 ();
 sg13g2_decap_8 FILLER_6_1260 ();
 sg13g2_decap_8 FILLER_6_1267 ();
 sg13g2_decap_8 FILLER_6_1274 ();
 sg13g2_decap_8 FILLER_6_1281 ();
 sg13g2_decap_8 FILLER_6_1288 ();
 sg13g2_decap_8 FILLER_6_1295 ();
 sg13g2_decap_8 FILLER_6_1302 ();
 sg13g2_decap_8 FILLER_6_1309 ();
 sg13g2_decap_8 FILLER_6_1316 ();
 sg13g2_decap_8 FILLER_6_1323 ();
 sg13g2_decap_8 FILLER_6_1330 ();
 sg13g2_decap_8 FILLER_6_1337 ();
 sg13g2_decap_8 FILLER_6_1344 ();
 sg13g2_decap_8 FILLER_6_1351 ();
 sg13g2_decap_8 FILLER_6_1358 ();
 sg13g2_decap_8 FILLER_6_1365 ();
 sg13g2_decap_8 FILLER_6_1372 ();
 sg13g2_decap_8 FILLER_6_1379 ();
 sg13g2_decap_8 FILLER_6_1386 ();
 sg13g2_decap_8 FILLER_6_1393 ();
 sg13g2_decap_8 FILLER_6_1400 ();
 sg13g2_decap_8 FILLER_6_1407 ();
 sg13g2_decap_8 FILLER_6_1414 ();
 sg13g2_decap_8 FILLER_6_1421 ();
 sg13g2_decap_8 FILLER_6_1428 ();
 sg13g2_decap_8 FILLER_6_1435 ();
 sg13g2_decap_8 FILLER_6_1442 ();
 sg13g2_decap_8 FILLER_6_1449 ();
 sg13g2_decap_8 FILLER_6_1456 ();
 sg13g2_decap_8 FILLER_6_1463 ();
 sg13g2_decap_8 FILLER_6_1470 ();
 sg13g2_decap_8 FILLER_6_1477 ();
 sg13g2_decap_8 FILLER_6_1484 ();
 sg13g2_decap_8 FILLER_6_1491 ();
 sg13g2_decap_8 FILLER_6_1498 ();
 sg13g2_decap_8 FILLER_6_1505 ();
 sg13g2_decap_8 FILLER_6_1512 ();
 sg13g2_decap_8 FILLER_6_1519 ();
 sg13g2_decap_8 FILLER_6_1526 ();
 sg13g2_decap_8 FILLER_6_1533 ();
 sg13g2_decap_8 FILLER_6_1540 ();
 sg13g2_decap_8 FILLER_6_1547 ();
 sg13g2_decap_8 FILLER_6_1554 ();
 sg13g2_decap_8 FILLER_6_1561 ();
 sg13g2_decap_8 FILLER_6_1568 ();
 sg13g2_decap_8 FILLER_6_1575 ();
 sg13g2_decap_8 FILLER_6_1582 ();
 sg13g2_decap_8 FILLER_6_1589 ();
 sg13g2_decap_8 FILLER_6_1596 ();
 sg13g2_decap_8 FILLER_6_1603 ();
 sg13g2_decap_8 FILLER_6_1610 ();
 sg13g2_decap_8 FILLER_6_1617 ();
 sg13g2_decap_8 FILLER_6_1624 ();
 sg13g2_decap_8 FILLER_6_1631 ();
 sg13g2_decap_8 FILLER_6_1638 ();
 sg13g2_decap_8 FILLER_6_1645 ();
 sg13g2_decap_8 FILLER_6_1652 ();
 sg13g2_decap_8 FILLER_6_1659 ();
 sg13g2_decap_8 FILLER_6_1666 ();
 sg13g2_decap_8 FILLER_6_1673 ();
 sg13g2_decap_8 FILLER_6_1680 ();
 sg13g2_decap_8 FILLER_6_1687 ();
 sg13g2_decap_8 FILLER_6_1694 ();
 sg13g2_decap_8 FILLER_6_1701 ();
 sg13g2_decap_8 FILLER_6_1708 ();
 sg13g2_decap_8 FILLER_6_1715 ();
 sg13g2_decap_8 FILLER_6_1722 ();
 sg13g2_decap_8 FILLER_6_1729 ();
 sg13g2_decap_8 FILLER_6_1736 ();
 sg13g2_decap_8 FILLER_6_1743 ();
 sg13g2_decap_8 FILLER_6_1750 ();
 sg13g2_decap_8 FILLER_6_1757 ();
 sg13g2_decap_8 FILLER_6_1764 ();
 sg13g2_decap_8 FILLER_6_1771 ();
 sg13g2_decap_8 FILLER_6_1778 ();
 sg13g2_decap_8 FILLER_6_1785 ();
 sg13g2_decap_8 FILLER_6_1792 ();
 sg13g2_decap_8 FILLER_6_1799 ();
 sg13g2_decap_8 FILLER_6_1806 ();
 sg13g2_decap_8 FILLER_6_1813 ();
 sg13g2_decap_8 FILLER_6_1820 ();
 sg13g2_decap_8 FILLER_6_1827 ();
 sg13g2_decap_8 FILLER_6_1834 ();
 sg13g2_decap_8 FILLER_6_1841 ();
 sg13g2_decap_8 FILLER_6_1848 ();
 sg13g2_decap_8 FILLER_6_1855 ();
 sg13g2_decap_8 FILLER_6_1862 ();
 sg13g2_decap_8 FILLER_6_1869 ();
 sg13g2_decap_8 FILLER_6_1876 ();
 sg13g2_decap_8 FILLER_6_1883 ();
 sg13g2_decap_8 FILLER_6_1890 ();
 sg13g2_decap_8 FILLER_6_1897 ();
 sg13g2_decap_8 FILLER_6_1904 ();
 sg13g2_decap_8 FILLER_6_1911 ();
 sg13g2_decap_8 FILLER_6_1918 ();
 sg13g2_decap_8 FILLER_6_1925 ();
 sg13g2_decap_8 FILLER_6_1932 ();
 sg13g2_decap_8 FILLER_6_1939 ();
 sg13g2_decap_8 FILLER_6_1946 ();
 sg13g2_decap_8 FILLER_6_1953 ();
 sg13g2_decap_8 FILLER_6_1960 ();
 sg13g2_decap_8 FILLER_6_1967 ();
 sg13g2_decap_8 FILLER_6_1974 ();
 sg13g2_decap_8 FILLER_6_1981 ();
 sg13g2_decap_8 FILLER_6_1988 ();
 sg13g2_decap_8 FILLER_6_1995 ();
 sg13g2_decap_8 FILLER_6_2002 ();
 sg13g2_decap_8 FILLER_6_2009 ();
 sg13g2_decap_8 FILLER_6_2016 ();
 sg13g2_decap_8 FILLER_6_2023 ();
 sg13g2_decap_8 FILLER_6_2030 ();
 sg13g2_decap_8 FILLER_6_2037 ();
 sg13g2_decap_8 FILLER_6_2044 ();
 sg13g2_decap_8 FILLER_6_2051 ();
 sg13g2_decap_8 FILLER_6_2058 ();
 sg13g2_decap_8 FILLER_6_2065 ();
 sg13g2_decap_8 FILLER_6_2072 ();
 sg13g2_decap_8 FILLER_6_2079 ();
 sg13g2_decap_8 FILLER_6_2086 ();
 sg13g2_decap_8 FILLER_6_2093 ();
 sg13g2_decap_8 FILLER_6_2100 ();
 sg13g2_decap_8 FILLER_6_2107 ();
 sg13g2_decap_8 FILLER_6_2114 ();
 sg13g2_decap_8 FILLER_6_2121 ();
 sg13g2_decap_8 FILLER_6_2128 ();
 sg13g2_decap_8 FILLER_6_2135 ();
 sg13g2_decap_8 FILLER_6_2142 ();
 sg13g2_decap_8 FILLER_6_2149 ();
 sg13g2_decap_8 FILLER_6_2156 ();
 sg13g2_decap_8 FILLER_6_2163 ();
 sg13g2_decap_8 FILLER_6_2170 ();
 sg13g2_decap_8 FILLER_6_2177 ();
 sg13g2_decap_8 FILLER_6_2184 ();
 sg13g2_decap_8 FILLER_6_2191 ();
 sg13g2_decap_8 FILLER_6_2198 ();
 sg13g2_decap_8 FILLER_6_2205 ();
 sg13g2_decap_8 FILLER_6_2212 ();
 sg13g2_decap_8 FILLER_6_2219 ();
 sg13g2_decap_8 FILLER_6_2226 ();
 sg13g2_decap_8 FILLER_6_2233 ();
 sg13g2_decap_8 FILLER_6_2240 ();
 sg13g2_decap_8 FILLER_6_2247 ();
 sg13g2_decap_8 FILLER_6_2254 ();
 sg13g2_decap_8 FILLER_6_2261 ();
 sg13g2_decap_8 FILLER_6_2268 ();
 sg13g2_decap_8 FILLER_6_2275 ();
 sg13g2_decap_8 FILLER_6_2282 ();
 sg13g2_decap_8 FILLER_6_2289 ();
 sg13g2_decap_8 FILLER_6_2296 ();
 sg13g2_decap_8 FILLER_6_2303 ();
 sg13g2_decap_8 FILLER_6_2310 ();
 sg13g2_decap_8 FILLER_6_2317 ();
 sg13g2_decap_8 FILLER_6_2324 ();
 sg13g2_decap_8 FILLER_6_2331 ();
 sg13g2_decap_8 FILLER_6_2338 ();
 sg13g2_decap_8 FILLER_6_2345 ();
 sg13g2_decap_8 FILLER_6_2352 ();
 sg13g2_decap_8 FILLER_6_2359 ();
 sg13g2_decap_8 FILLER_6_2366 ();
 sg13g2_decap_8 FILLER_6_2373 ();
 sg13g2_decap_8 FILLER_6_2380 ();
 sg13g2_decap_8 FILLER_6_2387 ();
 sg13g2_decap_8 FILLER_6_2394 ();
 sg13g2_decap_8 FILLER_6_2401 ();
 sg13g2_decap_8 FILLER_6_2408 ();
 sg13g2_decap_8 FILLER_6_2415 ();
 sg13g2_decap_8 FILLER_6_2422 ();
 sg13g2_decap_8 FILLER_6_2429 ();
 sg13g2_decap_8 FILLER_6_2436 ();
 sg13g2_decap_8 FILLER_6_2443 ();
 sg13g2_decap_8 FILLER_6_2450 ();
 sg13g2_decap_8 FILLER_6_2457 ();
 sg13g2_decap_8 FILLER_6_2464 ();
 sg13g2_decap_8 FILLER_6_2471 ();
 sg13g2_decap_8 FILLER_6_2478 ();
 sg13g2_decap_8 FILLER_6_2485 ();
 sg13g2_decap_8 FILLER_6_2492 ();
 sg13g2_decap_8 FILLER_6_2499 ();
 sg13g2_decap_8 FILLER_6_2506 ();
 sg13g2_decap_8 FILLER_6_2513 ();
 sg13g2_decap_8 FILLER_6_2520 ();
 sg13g2_decap_8 FILLER_6_2527 ();
 sg13g2_decap_8 FILLER_6_2534 ();
 sg13g2_decap_8 FILLER_6_2541 ();
 sg13g2_decap_8 FILLER_6_2548 ();
 sg13g2_decap_8 FILLER_6_2555 ();
 sg13g2_decap_8 FILLER_6_2562 ();
 sg13g2_decap_8 FILLER_6_2569 ();
 sg13g2_decap_8 FILLER_6_2576 ();
 sg13g2_decap_8 FILLER_6_2583 ();
 sg13g2_decap_8 FILLER_6_2590 ();
 sg13g2_decap_8 FILLER_6_2597 ();
 sg13g2_decap_8 FILLER_6_2604 ();
 sg13g2_decap_8 FILLER_6_2611 ();
 sg13g2_decap_8 FILLER_6_2618 ();
 sg13g2_decap_8 FILLER_6_2625 ();
 sg13g2_decap_8 FILLER_6_2632 ();
 sg13g2_decap_8 FILLER_6_2639 ();
 sg13g2_decap_8 FILLER_6_2646 ();
 sg13g2_decap_8 FILLER_6_2653 ();
 sg13g2_decap_8 FILLER_6_2660 ();
 sg13g2_decap_8 FILLER_6_2667 ();
 sg13g2_decap_8 FILLER_6_2674 ();
 sg13g2_decap_8 FILLER_6_2681 ();
 sg13g2_decap_8 FILLER_6_2688 ();
 sg13g2_decap_8 FILLER_6_2695 ();
 sg13g2_decap_8 FILLER_6_2702 ();
 sg13g2_decap_8 FILLER_6_2709 ();
 sg13g2_decap_8 FILLER_6_2716 ();
 sg13g2_decap_8 FILLER_6_2723 ();
 sg13g2_decap_8 FILLER_6_2730 ();
 sg13g2_decap_8 FILLER_6_2737 ();
 sg13g2_decap_8 FILLER_6_2744 ();
 sg13g2_decap_8 FILLER_6_2751 ();
 sg13g2_decap_8 FILLER_6_2758 ();
 sg13g2_decap_8 FILLER_6_2765 ();
 sg13g2_decap_8 FILLER_6_2772 ();
 sg13g2_decap_8 FILLER_6_2779 ();
 sg13g2_decap_8 FILLER_6_2786 ();
 sg13g2_decap_8 FILLER_6_2793 ();
 sg13g2_decap_8 FILLER_6_2800 ();
 sg13g2_decap_8 FILLER_6_2807 ();
 sg13g2_decap_8 FILLER_6_2814 ();
 sg13g2_decap_8 FILLER_6_2821 ();
 sg13g2_decap_8 FILLER_6_2828 ();
 sg13g2_decap_8 FILLER_6_2835 ();
 sg13g2_decap_8 FILLER_6_2842 ();
 sg13g2_decap_8 FILLER_6_2849 ();
 sg13g2_decap_8 FILLER_6_2856 ();
 sg13g2_decap_8 FILLER_6_2863 ();
 sg13g2_decap_8 FILLER_6_2870 ();
 sg13g2_decap_8 FILLER_6_2877 ();
 sg13g2_decap_8 FILLER_6_2884 ();
 sg13g2_decap_8 FILLER_6_2891 ();
 sg13g2_decap_8 FILLER_6_2898 ();
 sg13g2_decap_8 FILLER_6_2905 ();
 sg13g2_decap_8 FILLER_6_2912 ();
 sg13g2_decap_8 FILLER_6_2919 ();
 sg13g2_decap_8 FILLER_6_2926 ();
 sg13g2_decap_8 FILLER_6_2933 ();
 sg13g2_decap_8 FILLER_6_2940 ();
 sg13g2_decap_8 FILLER_6_2947 ();
 sg13g2_decap_8 FILLER_6_2954 ();
 sg13g2_decap_8 FILLER_6_2961 ();
 sg13g2_decap_8 FILLER_6_2968 ();
 sg13g2_decap_8 FILLER_6_2975 ();
 sg13g2_decap_8 FILLER_6_2982 ();
 sg13g2_decap_8 FILLER_6_2989 ();
 sg13g2_decap_8 FILLER_6_2996 ();
 sg13g2_decap_8 FILLER_6_3003 ();
 sg13g2_decap_8 FILLER_6_3010 ();
 sg13g2_decap_8 FILLER_6_3017 ();
 sg13g2_decap_8 FILLER_6_3024 ();
 sg13g2_decap_8 FILLER_6_3031 ();
 sg13g2_decap_8 FILLER_6_3038 ();
 sg13g2_decap_8 FILLER_6_3045 ();
 sg13g2_decap_8 FILLER_6_3052 ();
 sg13g2_decap_8 FILLER_6_3059 ();
 sg13g2_decap_8 FILLER_6_3066 ();
 sg13g2_decap_8 FILLER_6_3073 ();
 sg13g2_decap_8 FILLER_6_3080 ();
 sg13g2_decap_8 FILLER_6_3087 ();
 sg13g2_decap_8 FILLER_6_3094 ();
 sg13g2_decap_8 FILLER_6_3101 ();
 sg13g2_decap_8 FILLER_6_3108 ();
 sg13g2_decap_8 FILLER_6_3115 ();
 sg13g2_decap_8 FILLER_6_3122 ();
 sg13g2_decap_8 FILLER_6_3129 ();
 sg13g2_decap_8 FILLER_6_3136 ();
 sg13g2_decap_8 FILLER_6_3143 ();
 sg13g2_decap_8 FILLER_6_3150 ();
 sg13g2_decap_8 FILLER_6_3157 ();
 sg13g2_decap_8 FILLER_6_3164 ();
 sg13g2_decap_8 FILLER_6_3171 ();
 sg13g2_decap_8 FILLER_6_3178 ();
 sg13g2_decap_8 FILLER_6_3185 ();
 sg13g2_decap_8 FILLER_6_3192 ();
 sg13g2_decap_8 FILLER_6_3199 ();
 sg13g2_decap_8 FILLER_6_3206 ();
 sg13g2_decap_8 FILLER_6_3213 ();
 sg13g2_decap_8 FILLER_6_3220 ();
 sg13g2_decap_8 FILLER_6_3227 ();
 sg13g2_decap_8 FILLER_6_3234 ();
 sg13g2_decap_8 FILLER_6_3241 ();
 sg13g2_decap_8 FILLER_6_3248 ();
 sg13g2_decap_8 FILLER_6_3255 ();
 sg13g2_decap_8 FILLER_6_3262 ();
 sg13g2_decap_8 FILLER_6_3269 ();
 sg13g2_decap_8 FILLER_6_3276 ();
 sg13g2_decap_8 FILLER_6_3283 ();
 sg13g2_decap_8 FILLER_6_3290 ();
 sg13g2_decap_8 FILLER_6_3297 ();
 sg13g2_decap_8 FILLER_6_3304 ();
 sg13g2_decap_8 FILLER_6_3311 ();
 sg13g2_decap_8 FILLER_6_3318 ();
 sg13g2_decap_8 FILLER_6_3325 ();
 sg13g2_decap_8 FILLER_6_3332 ();
 sg13g2_decap_8 FILLER_6_3339 ();
 sg13g2_decap_8 FILLER_6_3346 ();
 sg13g2_decap_8 FILLER_6_3353 ();
 sg13g2_decap_8 FILLER_6_3360 ();
 sg13g2_decap_8 FILLER_6_3367 ();
 sg13g2_decap_8 FILLER_6_3374 ();
 sg13g2_decap_8 FILLER_6_3381 ();
 sg13g2_decap_8 FILLER_6_3388 ();
 sg13g2_decap_8 FILLER_6_3395 ();
 sg13g2_decap_8 FILLER_6_3402 ();
 sg13g2_decap_8 FILLER_6_3409 ();
 sg13g2_decap_8 FILLER_6_3416 ();
 sg13g2_decap_8 FILLER_6_3423 ();
 sg13g2_decap_8 FILLER_6_3430 ();
 sg13g2_decap_8 FILLER_6_3437 ();
 sg13g2_decap_8 FILLER_6_3444 ();
 sg13g2_decap_8 FILLER_6_3451 ();
 sg13g2_decap_8 FILLER_6_3458 ();
 sg13g2_decap_8 FILLER_6_3465 ();
 sg13g2_decap_8 FILLER_6_3472 ();
 sg13g2_decap_8 FILLER_6_3479 ();
 sg13g2_decap_8 FILLER_6_3486 ();
 sg13g2_decap_8 FILLER_6_3493 ();
 sg13g2_decap_8 FILLER_6_3500 ();
 sg13g2_decap_8 FILLER_6_3507 ();
 sg13g2_decap_8 FILLER_6_3514 ();
 sg13g2_decap_8 FILLER_6_3521 ();
 sg13g2_decap_8 FILLER_6_3528 ();
 sg13g2_decap_8 FILLER_6_3535 ();
 sg13g2_decap_8 FILLER_6_3542 ();
 sg13g2_decap_8 FILLER_6_3549 ();
 sg13g2_decap_8 FILLER_6_3556 ();
 sg13g2_decap_8 FILLER_6_3563 ();
 sg13g2_decap_8 FILLER_6_3570 ();
 sg13g2_fill_2 FILLER_6_3577 ();
 sg13g2_fill_1 FILLER_6_3579 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_decap_8 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_7_868 ();
 sg13g2_decap_8 FILLER_7_875 ();
 sg13g2_decap_8 FILLER_7_882 ();
 sg13g2_decap_8 FILLER_7_889 ();
 sg13g2_decap_8 FILLER_7_896 ();
 sg13g2_decap_8 FILLER_7_903 ();
 sg13g2_decap_8 FILLER_7_910 ();
 sg13g2_decap_8 FILLER_7_917 ();
 sg13g2_decap_8 FILLER_7_924 ();
 sg13g2_decap_8 FILLER_7_931 ();
 sg13g2_decap_8 FILLER_7_938 ();
 sg13g2_decap_8 FILLER_7_945 ();
 sg13g2_decap_8 FILLER_7_952 ();
 sg13g2_decap_8 FILLER_7_959 ();
 sg13g2_decap_8 FILLER_7_966 ();
 sg13g2_decap_8 FILLER_7_973 ();
 sg13g2_decap_8 FILLER_7_980 ();
 sg13g2_decap_8 FILLER_7_987 ();
 sg13g2_decap_8 FILLER_7_994 ();
 sg13g2_decap_8 FILLER_7_1001 ();
 sg13g2_decap_8 FILLER_7_1008 ();
 sg13g2_decap_8 FILLER_7_1015 ();
 sg13g2_decap_8 FILLER_7_1022 ();
 sg13g2_decap_8 FILLER_7_1029 ();
 sg13g2_decap_8 FILLER_7_1036 ();
 sg13g2_decap_8 FILLER_7_1043 ();
 sg13g2_decap_8 FILLER_7_1050 ();
 sg13g2_decap_8 FILLER_7_1057 ();
 sg13g2_decap_8 FILLER_7_1064 ();
 sg13g2_decap_8 FILLER_7_1071 ();
 sg13g2_decap_8 FILLER_7_1078 ();
 sg13g2_decap_8 FILLER_7_1085 ();
 sg13g2_decap_8 FILLER_7_1092 ();
 sg13g2_decap_8 FILLER_7_1099 ();
 sg13g2_decap_8 FILLER_7_1106 ();
 sg13g2_decap_8 FILLER_7_1113 ();
 sg13g2_decap_8 FILLER_7_1120 ();
 sg13g2_decap_8 FILLER_7_1127 ();
 sg13g2_decap_8 FILLER_7_1134 ();
 sg13g2_decap_8 FILLER_7_1141 ();
 sg13g2_decap_8 FILLER_7_1148 ();
 sg13g2_decap_8 FILLER_7_1155 ();
 sg13g2_decap_8 FILLER_7_1162 ();
 sg13g2_decap_8 FILLER_7_1169 ();
 sg13g2_decap_8 FILLER_7_1176 ();
 sg13g2_decap_8 FILLER_7_1183 ();
 sg13g2_decap_8 FILLER_7_1190 ();
 sg13g2_decap_8 FILLER_7_1197 ();
 sg13g2_decap_8 FILLER_7_1204 ();
 sg13g2_decap_8 FILLER_7_1211 ();
 sg13g2_decap_8 FILLER_7_1218 ();
 sg13g2_decap_8 FILLER_7_1225 ();
 sg13g2_decap_8 FILLER_7_1232 ();
 sg13g2_decap_8 FILLER_7_1239 ();
 sg13g2_decap_8 FILLER_7_1246 ();
 sg13g2_decap_8 FILLER_7_1253 ();
 sg13g2_decap_8 FILLER_7_1260 ();
 sg13g2_decap_8 FILLER_7_1267 ();
 sg13g2_decap_8 FILLER_7_1274 ();
 sg13g2_decap_8 FILLER_7_1281 ();
 sg13g2_decap_8 FILLER_7_1288 ();
 sg13g2_decap_8 FILLER_7_1295 ();
 sg13g2_decap_8 FILLER_7_1302 ();
 sg13g2_decap_8 FILLER_7_1309 ();
 sg13g2_decap_8 FILLER_7_1316 ();
 sg13g2_decap_8 FILLER_7_1323 ();
 sg13g2_decap_8 FILLER_7_1330 ();
 sg13g2_decap_8 FILLER_7_1337 ();
 sg13g2_decap_8 FILLER_7_1344 ();
 sg13g2_decap_8 FILLER_7_1351 ();
 sg13g2_decap_8 FILLER_7_1358 ();
 sg13g2_decap_8 FILLER_7_1365 ();
 sg13g2_decap_8 FILLER_7_1372 ();
 sg13g2_decap_8 FILLER_7_1379 ();
 sg13g2_decap_8 FILLER_7_1386 ();
 sg13g2_decap_8 FILLER_7_1393 ();
 sg13g2_decap_8 FILLER_7_1400 ();
 sg13g2_decap_8 FILLER_7_1407 ();
 sg13g2_decap_8 FILLER_7_1414 ();
 sg13g2_decap_8 FILLER_7_1421 ();
 sg13g2_decap_8 FILLER_7_1428 ();
 sg13g2_decap_8 FILLER_7_1435 ();
 sg13g2_decap_8 FILLER_7_1442 ();
 sg13g2_decap_8 FILLER_7_1449 ();
 sg13g2_decap_8 FILLER_7_1456 ();
 sg13g2_decap_8 FILLER_7_1463 ();
 sg13g2_decap_8 FILLER_7_1470 ();
 sg13g2_decap_8 FILLER_7_1477 ();
 sg13g2_decap_8 FILLER_7_1484 ();
 sg13g2_decap_8 FILLER_7_1491 ();
 sg13g2_decap_8 FILLER_7_1498 ();
 sg13g2_decap_8 FILLER_7_1505 ();
 sg13g2_decap_8 FILLER_7_1512 ();
 sg13g2_decap_8 FILLER_7_1519 ();
 sg13g2_decap_8 FILLER_7_1526 ();
 sg13g2_decap_8 FILLER_7_1533 ();
 sg13g2_decap_8 FILLER_7_1540 ();
 sg13g2_decap_8 FILLER_7_1547 ();
 sg13g2_decap_8 FILLER_7_1554 ();
 sg13g2_decap_8 FILLER_7_1561 ();
 sg13g2_decap_8 FILLER_7_1568 ();
 sg13g2_decap_8 FILLER_7_1575 ();
 sg13g2_decap_8 FILLER_7_1582 ();
 sg13g2_decap_8 FILLER_7_1589 ();
 sg13g2_decap_8 FILLER_7_1596 ();
 sg13g2_decap_8 FILLER_7_1603 ();
 sg13g2_decap_8 FILLER_7_1610 ();
 sg13g2_decap_8 FILLER_7_1617 ();
 sg13g2_decap_8 FILLER_7_1624 ();
 sg13g2_decap_8 FILLER_7_1631 ();
 sg13g2_decap_8 FILLER_7_1638 ();
 sg13g2_decap_8 FILLER_7_1645 ();
 sg13g2_decap_8 FILLER_7_1652 ();
 sg13g2_decap_8 FILLER_7_1659 ();
 sg13g2_decap_8 FILLER_7_1666 ();
 sg13g2_decap_8 FILLER_7_1673 ();
 sg13g2_decap_8 FILLER_7_1680 ();
 sg13g2_decap_8 FILLER_7_1687 ();
 sg13g2_decap_8 FILLER_7_1694 ();
 sg13g2_decap_8 FILLER_7_1701 ();
 sg13g2_decap_8 FILLER_7_1708 ();
 sg13g2_decap_8 FILLER_7_1715 ();
 sg13g2_decap_8 FILLER_7_1722 ();
 sg13g2_decap_8 FILLER_7_1729 ();
 sg13g2_decap_8 FILLER_7_1736 ();
 sg13g2_decap_8 FILLER_7_1743 ();
 sg13g2_decap_8 FILLER_7_1750 ();
 sg13g2_decap_8 FILLER_7_1757 ();
 sg13g2_decap_8 FILLER_7_1764 ();
 sg13g2_decap_8 FILLER_7_1771 ();
 sg13g2_decap_8 FILLER_7_1778 ();
 sg13g2_decap_8 FILLER_7_1785 ();
 sg13g2_decap_8 FILLER_7_1792 ();
 sg13g2_decap_8 FILLER_7_1799 ();
 sg13g2_decap_8 FILLER_7_1806 ();
 sg13g2_decap_8 FILLER_7_1813 ();
 sg13g2_decap_8 FILLER_7_1820 ();
 sg13g2_decap_8 FILLER_7_1827 ();
 sg13g2_decap_8 FILLER_7_1834 ();
 sg13g2_decap_8 FILLER_7_1841 ();
 sg13g2_decap_8 FILLER_7_1848 ();
 sg13g2_decap_8 FILLER_7_1855 ();
 sg13g2_decap_8 FILLER_7_1862 ();
 sg13g2_decap_8 FILLER_7_1869 ();
 sg13g2_decap_8 FILLER_7_1876 ();
 sg13g2_decap_8 FILLER_7_1883 ();
 sg13g2_decap_8 FILLER_7_1890 ();
 sg13g2_decap_8 FILLER_7_1897 ();
 sg13g2_decap_8 FILLER_7_1904 ();
 sg13g2_decap_8 FILLER_7_1911 ();
 sg13g2_decap_8 FILLER_7_1918 ();
 sg13g2_decap_8 FILLER_7_1925 ();
 sg13g2_decap_8 FILLER_7_1932 ();
 sg13g2_decap_8 FILLER_7_1939 ();
 sg13g2_decap_8 FILLER_7_1946 ();
 sg13g2_decap_8 FILLER_7_1953 ();
 sg13g2_decap_8 FILLER_7_1960 ();
 sg13g2_decap_8 FILLER_7_1967 ();
 sg13g2_decap_8 FILLER_7_1974 ();
 sg13g2_decap_8 FILLER_7_1981 ();
 sg13g2_decap_8 FILLER_7_1988 ();
 sg13g2_decap_8 FILLER_7_1995 ();
 sg13g2_decap_8 FILLER_7_2002 ();
 sg13g2_decap_8 FILLER_7_2009 ();
 sg13g2_decap_8 FILLER_7_2016 ();
 sg13g2_decap_8 FILLER_7_2023 ();
 sg13g2_decap_8 FILLER_7_2030 ();
 sg13g2_decap_8 FILLER_7_2037 ();
 sg13g2_decap_8 FILLER_7_2044 ();
 sg13g2_decap_8 FILLER_7_2051 ();
 sg13g2_decap_8 FILLER_7_2058 ();
 sg13g2_decap_8 FILLER_7_2065 ();
 sg13g2_decap_8 FILLER_7_2072 ();
 sg13g2_decap_8 FILLER_7_2079 ();
 sg13g2_decap_8 FILLER_7_2086 ();
 sg13g2_decap_8 FILLER_7_2093 ();
 sg13g2_decap_8 FILLER_7_2100 ();
 sg13g2_decap_8 FILLER_7_2107 ();
 sg13g2_decap_8 FILLER_7_2114 ();
 sg13g2_decap_8 FILLER_7_2121 ();
 sg13g2_decap_8 FILLER_7_2128 ();
 sg13g2_decap_8 FILLER_7_2135 ();
 sg13g2_decap_8 FILLER_7_2142 ();
 sg13g2_decap_8 FILLER_7_2149 ();
 sg13g2_decap_8 FILLER_7_2156 ();
 sg13g2_decap_8 FILLER_7_2163 ();
 sg13g2_decap_8 FILLER_7_2170 ();
 sg13g2_decap_8 FILLER_7_2177 ();
 sg13g2_decap_8 FILLER_7_2184 ();
 sg13g2_decap_8 FILLER_7_2191 ();
 sg13g2_decap_8 FILLER_7_2198 ();
 sg13g2_decap_8 FILLER_7_2205 ();
 sg13g2_decap_8 FILLER_7_2212 ();
 sg13g2_decap_8 FILLER_7_2219 ();
 sg13g2_decap_8 FILLER_7_2226 ();
 sg13g2_decap_8 FILLER_7_2233 ();
 sg13g2_decap_8 FILLER_7_2240 ();
 sg13g2_decap_8 FILLER_7_2247 ();
 sg13g2_decap_8 FILLER_7_2254 ();
 sg13g2_decap_8 FILLER_7_2261 ();
 sg13g2_decap_8 FILLER_7_2268 ();
 sg13g2_decap_8 FILLER_7_2275 ();
 sg13g2_decap_8 FILLER_7_2282 ();
 sg13g2_decap_8 FILLER_7_2289 ();
 sg13g2_decap_8 FILLER_7_2296 ();
 sg13g2_decap_8 FILLER_7_2303 ();
 sg13g2_decap_8 FILLER_7_2310 ();
 sg13g2_decap_8 FILLER_7_2317 ();
 sg13g2_decap_8 FILLER_7_2324 ();
 sg13g2_decap_8 FILLER_7_2331 ();
 sg13g2_decap_8 FILLER_7_2338 ();
 sg13g2_decap_8 FILLER_7_2345 ();
 sg13g2_decap_8 FILLER_7_2352 ();
 sg13g2_decap_8 FILLER_7_2359 ();
 sg13g2_decap_8 FILLER_7_2366 ();
 sg13g2_decap_8 FILLER_7_2373 ();
 sg13g2_decap_8 FILLER_7_2380 ();
 sg13g2_decap_8 FILLER_7_2387 ();
 sg13g2_decap_8 FILLER_7_2394 ();
 sg13g2_decap_8 FILLER_7_2401 ();
 sg13g2_decap_8 FILLER_7_2408 ();
 sg13g2_decap_8 FILLER_7_2415 ();
 sg13g2_decap_8 FILLER_7_2422 ();
 sg13g2_decap_8 FILLER_7_2429 ();
 sg13g2_decap_8 FILLER_7_2436 ();
 sg13g2_decap_8 FILLER_7_2443 ();
 sg13g2_decap_8 FILLER_7_2450 ();
 sg13g2_decap_8 FILLER_7_2457 ();
 sg13g2_decap_8 FILLER_7_2464 ();
 sg13g2_decap_8 FILLER_7_2471 ();
 sg13g2_decap_8 FILLER_7_2478 ();
 sg13g2_decap_8 FILLER_7_2485 ();
 sg13g2_decap_8 FILLER_7_2492 ();
 sg13g2_decap_8 FILLER_7_2499 ();
 sg13g2_decap_8 FILLER_7_2506 ();
 sg13g2_decap_8 FILLER_7_2513 ();
 sg13g2_decap_8 FILLER_7_2520 ();
 sg13g2_decap_8 FILLER_7_2527 ();
 sg13g2_decap_8 FILLER_7_2534 ();
 sg13g2_decap_8 FILLER_7_2541 ();
 sg13g2_decap_8 FILLER_7_2548 ();
 sg13g2_decap_8 FILLER_7_2555 ();
 sg13g2_decap_8 FILLER_7_2562 ();
 sg13g2_decap_8 FILLER_7_2569 ();
 sg13g2_decap_8 FILLER_7_2576 ();
 sg13g2_decap_8 FILLER_7_2583 ();
 sg13g2_decap_8 FILLER_7_2590 ();
 sg13g2_decap_8 FILLER_7_2597 ();
 sg13g2_decap_8 FILLER_7_2604 ();
 sg13g2_decap_8 FILLER_7_2611 ();
 sg13g2_decap_8 FILLER_7_2618 ();
 sg13g2_decap_8 FILLER_7_2625 ();
 sg13g2_decap_8 FILLER_7_2632 ();
 sg13g2_decap_8 FILLER_7_2639 ();
 sg13g2_decap_8 FILLER_7_2646 ();
 sg13g2_decap_8 FILLER_7_2653 ();
 sg13g2_decap_8 FILLER_7_2660 ();
 sg13g2_decap_8 FILLER_7_2667 ();
 sg13g2_decap_8 FILLER_7_2674 ();
 sg13g2_decap_8 FILLER_7_2681 ();
 sg13g2_decap_8 FILLER_7_2688 ();
 sg13g2_decap_8 FILLER_7_2695 ();
 sg13g2_decap_8 FILLER_7_2702 ();
 sg13g2_decap_8 FILLER_7_2709 ();
 sg13g2_decap_8 FILLER_7_2716 ();
 sg13g2_decap_8 FILLER_7_2723 ();
 sg13g2_decap_8 FILLER_7_2730 ();
 sg13g2_decap_8 FILLER_7_2737 ();
 sg13g2_decap_8 FILLER_7_2744 ();
 sg13g2_decap_8 FILLER_7_2751 ();
 sg13g2_decap_8 FILLER_7_2758 ();
 sg13g2_decap_8 FILLER_7_2765 ();
 sg13g2_decap_8 FILLER_7_2772 ();
 sg13g2_decap_8 FILLER_7_2779 ();
 sg13g2_decap_8 FILLER_7_2786 ();
 sg13g2_decap_8 FILLER_7_2793 ();
 sg13g2_decap_8 FILLER_7_2800 ();
 sg13g2_decap_8 FILLER_7_2807 ();
 sg13g2_decap_8 FILLER_7_2814 ();
 sg13g2_decap_8 FILLER_7_2821 ();
 sg13g2_decap_8 FILLER_7_2828 ();
 sg13g2_decap_8 FILLER_7_2835 ();
 sg13g2_decap_8 FILLER_7_2842 ();
 sg13g2_decap_8 FILLER_7_2849 ();
 sg13g2_decap_8 FILLER_7_2856 ();
 sg13g2_decap_8 FILLER_7_2863 ();
 sg13g2_decap_8 FILLER_7_2870 ();
 sg13g2_decap_8 FILLER_7_2877 ();
 sg13g2_decap_8 FILLER_7_2884 ();
 sg13g2_decap_8 FILLER_7_2891 ();
 sg13g2_decap_8 FILLER_7_2898 ();
 sg13g2_decap_8 FILLER_7_2905 ();
 sg13g2_decap_8 FILLER_7_2912 ();
 sg13g2_decap_8 FILLER_7_2919 ();
 sg13g2_decap_8 FILLER_7_2926 ();
 sg13g2_decap_8 FILLER_7_2933 ();
 sg13g2_decap_8 FILLER_7_2940 ();
 sg13g2_decap_8 FILLER_7_2947 ();
 sg13g2_decap_8 FILLER_7_2954 ();
 sg13g2_decap_8 FILLER_7_2961 ();
 sg13g2_decap_8 FILLER_7_2968 ();
 sg13g2_decap_8 FILLER_7_2975 ();
 sg13g2_decap_8 FILLER_7_2982 ();
 sg13g2_decap_8 FILLER_7_2989 ();
 sg13g2_decap_8 FILLER_7_2996 ();
 sg13g2_decap_8 FILLER_7_3003 ();
 sg13g2_decap_8 FILLER_7_3010 ();
 sg13g2_decap_8 FILLER_7_3017 ();
 sg13g2_decap_8 FILLER_7_3024 ();
 sg13g2_decap_8 FILLER_7_3031 ();
 sg13g2_decap_8 FILLER_7_3038 ();
 sg13g2_decap_8 FILLER_7_3045 ();
 sg13g2_decap_8 FILLER_7_3052 ();
 sg13g2_decap_8 FILLER_7_3059 ();
 sg13g2_decap_8 FILLER_7_3066 ();
 sg13g2_decap_8 FILLER_7_3073 ();
 sg13g2_decap_8 FILLER_7_3080 ();
 sg13g2_decap_8 FILLER_7_3087 ();
 sg13g2_decap_8 FILLER_7_3094 ();
 sg13g2_decap_8 FILLER_7_3101 ();
 sg13g2_decap_8 FILLER_7_3108 ();
 sg13g2_decap_8 FILLER_7_3115 ();
 sg13g2_decap_8 FILLER_7_3122 ();
 sg13g2_decap_8 FILLER_7_3129 ();
 sg13g2_decap_8 FILLER_7_3136 ();
 sg13g2_decap_8 FILLER_7_3143 ();
 sg13g2_decap_8 FILLER_7_3150 ();
 sg13g2_decap_8 FILLER_7_3157 ();
 sg13g2_decap_8 FILLER_7_3164 ();
 sg13g2_decap_8 FILLER_7_3171 ();
 sg13g2_decap_8 FILLER_7_3178 ();
 sg13g2_decap_8 FILLER_7_3185 ();
 sg13g2_decap_8 FILLER_7_3192 ();
 sg13g2_decap_8 FILLER_7_3199 ();
 sg13g2_decap_8 FILLER_7_3206 ();
 sg13g2_decap_8 FILLER_7_3213 ();
 sg13g2_decap_8 FILLER_7_3220 ();
 sg13g2_decap_8 FILLER_7_3227 ();
 sg13g2_decap_8 FILLER_7_3234 ();
 sg13g2_decap_8 FILLER_7_3241 ();
 sg13g2_decap_8 FILLER_7_3248 ();
 sg13g2_decap_8 FILLER_7_3255 ();
 sg13g2_decap_8 FILLER_7_3262 ();
 sg13g2_decap_8 FILLER_7_3269 ();
 sg13g2_decap_8 FILLER_7_3276 ();
 sg13g2_decap_8 FILLER_7_3283 ();
 sg13g2_decap_8 FILLER_7_3290 ();
 sg13g2_decap_8 FILLER_7_3297 ();
 sg13g2_decap_8 FILLER_7_3304 ();
 sg13g2_decap_8 FILLER_7_3311 ();
 sg13g2_decap_8 FILLER_7_3318 ();
 sg13g2_decap_8 FILLER_7_3325 ();
 sg13g2_decap_8 FILLER_7_3332 ();
 sg13g2_decap_8 FILLER_7_3339 ();
 sg13g2_decap_8 FILLER_7_3346 ();
 sg13g2_decap_8 FILLER_7_3353 ();
 sg13g2_decap_8 FILLER_7_3360 ();
 sg13g2_decap_8 FILLER_7_3367 ();
 sg13g2_decap_8 FILLER_7_3374 ();
 sg13g2_decap_8 FILLER_7_3381 ();
 sg13g2_decap_8 FILLER_7_3388 ();
 sg13g2_decap_8 FILLER_7_3395 ();
 sg13g2_decap_8 FILLER_7_3402 ();
 sg13g2_decap_8 FILLER_7_3409 ();
 sg13g2_decap_8 FILLER_7_3416 ();
 sg13g2_decap_8 FILLER_7_3423 ();
 sg13g2_decap_8 FILLER_7_3430 ();
 sg13g2_decap_8 FILLER_7_3437 ();
 sg13g2_decap_8 FILLER_7_3444 ();
 sg13g2_decap_8 FILLER_7_3451 ();
 sg13g2_decap_8 FILLER_7_3458 ();
 sg13g2_decap_8 FILLER_7_3465 ();
 sg13g2_decap_8 FILLER_7_3472 ();
 sg13g2_decap_8 FILLER_7_3479 ();
 sg13g2_decap_8 FILLER_7_3486 ();
 sg13g2_decap_8 FILLER_7_3493 ();
 sg13g2_decap_8 FILLER_7_3500 ();
 sg13g2_decap_8 FILLER_7_3507 ();
 sg13g2_decap_8 FILLER_7_3514 ();
 sg13g2_decap_8 FILLER_7_3521 ();
 sg13g2_decap_8 FILLER_7_3528 ();
 sg13g2_decap_8 FILLER_7_3535 ();
 sg13g2_decap_8 FILLER_7_3542 ();
 sg13g2_decap_8 FILLER_7_3549 ();
 sg13g2_decap_8 FILLER_7_3556 ();
 sg13g2_decap_8 FILLER_7_3563 ();
 sg13g2_decap_8 FILLER_7_3570 ();
 sg13g2_fill_2 FILLER_7_3577 ();
 sg13g2_fill_1 FILLER_7_3579 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_decap_8 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_8_868 ();
 sg13g2_decap_8 FILLER_8_875 ();
 sg13g2_decap_8 FILLER_8_882 ();
 sg13g2_decap_8 FILLER_8_889 ();
 sg13g2_decap_8 FILLER_8_896 ();
 sg13g2_decap_8 FILLER_8_903 ();
 sg13g2_decap_8 FILLER_8_910 ();
 sg13g2_decap_8 FILLER_8_917 ();
 sg13g2_decap_8 FILLER_8_924 ();
 sg13g2_decap_8 FILLER_8_931 ();
 sg13g2_decap_8 FILLER_8_938 ();
 sg13g2_decap_8 FILLER_8_945 ();
 sg13g2_decap_8 FILLER_8_952 ();
 sg13g2_decap_8 FILLER_8_959 ();
 sg13g2_decap_8 FILLER_8_966 ();
 sg13g2_decap_8 FILLER_8_973 ();
 sg13g2_decap_8 FILLER_8_980 ();
 sg13g2_decap_8 FILLER_8_987 ();
 sg13g2_decap_8 FILLER_8_994 ();
 sg13g2_decap_8 FILLER_8_1001 ();
 sg13g2_decap_8 FILLER_8_1008 ();
 sg13g2_decap_8 FILLER_8_1015 ();
 sg13g2_decap_8 FILLER_8_1022 ();
 sg13g2_decap_8 FILLER_8_1029 ();
 sg13g2_decap_8 FILLER_8_1036 ();
 sg13g2_decap_8 FILLER_8_1043 ();
 sg13g2_decap_8 FILLER_8_1050 ();
 sg13g2_decap_8 FILLER_8_1057 ();
 sg13g2_decap_8 FILLER_8_1064 ();
 sg13g2_decap_8 FILLER_8_1071 ();
 sg13g2_decap_8 FILLER_8_1078 ();
 sg13g2_decap_8 FILLER_8_1085 ();
 sg13g2_decap_8 FILLER_8_1092 ();
 sg13g2_decap_8 FILLER_8_1099 ();
 sg13g2_decap_8 FILLER_8_1106 ();
 sg13g2_decap_8 FILLER_8_1113 ();
 sg13g2_decap_8 FILLER_8_1120 ();
 sg13g2_decap_8 FILLER_8_1127 ();
 sg13g2_decap_8 FILLER_8_1134 ();
 sg13g2_decap_8 FILLER_8_1141 ();
 sg13g2_decap_8 FILLER_8_1148 ();
 sg13g2_decap_8 FILLER_8_1155 ();
 sg13g2_decap_8 FILLER_8_1162 ();
 sg13g2_decap_8 FILLER_8_1169 ();
 sg13g2_decap_8 FILLER_8_1176 ();
 sg13g2_decap_8 FILLER_8_1183 ();
 sg13g2_decap_8 FILLER_8_1190 ();
 sg13g2_decap_8 FILLER_8_1197 ();
 sg13g2_decap_8 FILLER_8_1204 ();
 sg13g2_decap_8 FILLER_8_1211 ();
 sg13g2_decap_8 FILLER_8_1218 ();
 sg13g2_decap_8 FILLER_8_1225 ();
 sg13g2_decap_8 FILLER_8_1232 ();
 sg13g2_decap_8 FILLER_8_1239 ();
 sg13g2_decap_8 FILLER_8_1246 ();
 sg13g2_decap_8 FILLER_8_1253 ();
 sg13g2_decap_8 FILLER_8_1260 ();
 sg13g2_decap_8 FILLER_8_1267 ();
 sg13g2_decap_8 FILLER_8_1274 ();
 sg13g2_decap_8 FILLER_8_1281 ();
 sg13g2_decap_8 FILLER_8_1288 ();
 sg13g2_decap_8 FILLER_8_1295 ();
 sg13g2_decap_8 FILLER_8_1302 ();
 sg13g2_decap_8 FILLER_8_1309 ();
 sg13g2_decap_8 FILLER_8_1316 ();
 sg13g2_decap_8 FILLER_8_1323 ();
 sg13g2_decap_8 FILLER_8_1330 ();
 sg13g2_decap_8 FILLER_8_1337 ();
 sg13g2_decap_8 FILLER_8_1344 ();
 sg13g2_decap_8 FILLER_8_1351 ();
 sg13g2_decap_8 FILLER_8_1358 ();
 sg13g2_decap_8 FILLER_8_1365 ();
 sg13g2_decap_8 FILLER_8_1372 ();
 sg13g2_decap_8 FILLER_8_1379 ();
 sg13g2_decap_8 FILLER_8_1386 ();
 sg13g2_decap_8 FILLER_8_1393 ();
 sg13g2_decap_8 FILLER_8_1400 ();
 sg13g2_decap_8 FILLER_8_1407 ();
 sg13g2_decap_8 FILLER_8_1414 ();
 sg13g2_decap_8 FILLER_8_1421 ();
 sg13g2_decap_8 FILLER_8_1428 ();
 sg13g2_decap_8 FILLER_8_1435 ();
 sg13g2_decap_8 FILLER_8_1442 ();
 sg13g2_decap_8 FILLER_8_1449 ();
 sg13g2_decap_8 FILLER_8_1456 ();
 sg13g2_decap_8 FILLER_8_1463 ();
 sg13g2_decap_8 FILLER_8_1470 ();
 sg13g2_decap_8 FILLER_8_1477 ();
 sg13g2_decap_8 FILLER_8_1484 ();
 sg13g2_decap_8 FILLER_8_1491 ();
 sg13g2_decap_8 FILLER_8_1498 ();
 sg13g2_decap_8 FILLER_8_1505 ();
 sg13g2_decap_8 FILLER_8_1512 ();
 sg13g2_decap_8 FILLER_8_1519 ();
 sg13g2_decap_8 FILLER_8_1526 ();
 sg13g2_decap_8 FILLER_8_1533 ();
 sg13g2_decap_8 FILLER_8_1540 ();
 sg13g2_decap_8 FILLER_8_1547 ();
 sg13g2_decap_8 FILLER_8_1554 ();
 sg13g2_decap_8 FILLER_8_1561 ();
 sg13g2_decap_8 FILLER_8_1568 ();
 sg13g2_decap_8 FILLER_8_1575 ();
 sg13g2_decap_8 FILLER_8_1582 ();
 sg13g2_decap_8 FILLER_8_1589 ();
 sg13g2_decap_8 FILLER_8_1596 ();
 sg13g2_decap_8 FILLER_8_1603 ();
 sg13g2_decap_8 FILLER_8_1610 ();
 sg13g2_decap_8 FILLER_8_1617 ();
 sg13g2_decap_8 FILLER_8_1624 ();
 sg13g2_decap_8 FILLER_8_1631 ();
 sg13g2_decap_8 FILLER_8_1638 ();
 sg13g2_decap_8 FILLER_8_1645 ();
 sg13g2_decap_8 FILLER_8_1652 ();
 sg13g2_decap_8 FILLER_8_1659 ();
 sg13g2_decap_8 FILLER_8_1666 ();
 sg13g2_decap_8 FILLER_8_1673 ();
 sg13g2_decap_8 FILLER_8_1680 ();
 sg13g2_decap_8 FILLER_8_1687 ();
 sg13g2_decap_8 FILLER_8_1694 ();
 sg13g2_decap_8 FILLER_8_1701 ();
 sg13g2_decap_8 FILLER_8_1708 ();
 sg13g2_decap_8 FILLER_8_1715 ();
 sg13g2_decap_8 FILLER_8_1722 ();
 sg13g2_decap_8 FILLER_8_1729 ();
 sg13g2_decap_8 FILLER_8_1736 ();
 sg13g2_decap_8 FILLER_8_1743 ();
 sg13g2_decap_8 FILLER_8_1750 ();
 sg13g2_decap_8 FILLER_8_1757 ();
 sg13g2_decap_8 FILLER_8_1764 ();
 sg13g2_decap_8 FILLER_8_1771 ();
 sg13g2_decap_8 FILLER_8_1778 ();
 sg13g2_decap_8 FILLER_8_1785 ();
 sg13g2_decap_8 FILLER_8_1792 ();
 sg13g2_decap_8 FILLER_8_1799 ();
 sg13g2_decap_8 FILLER_8_1806 ();
 sg13g2_decap_8 FILLER_8_1813 ();
 sg13g2_decap_8 FILLER_8_1820 ();
 sg13g2_decap_8 FILLER_8_1827 ();
 sg13g2_decap_8 FILLER_8_1834 ();
 sg13g2_decap_8 FILLER_8_1841 ();
 sg13g2_decap_8 FILLER_8_1848 ();
 sg13g2_decap_8 FILLER_8_1855 ();
 sg13g2_decap_8 FILLER_8_1862 ();
 sg13g2_decap_8 FILLER_8_1869 ();
 sg13g2_decap_8 FILLER_8_1876 ();
 sg13g2_decap_8 FILLER_8_1883 ();
 sg13g2_decap_8 FILLER_8_1890 ();
 sg13g2_decap_8 FILLER_8_1897 ();
 sg13g2_decap_8 FILLER_8_1904 ();
 sg13g2_decap_8 FILLER_8_1911 ();
 sg13g2_decap_8 FILLER_8_1918 ();
 sg13g2_decap_8 FILLER_8_1925 ();
 sg13g2_decap_8 FILLER_8_1932 ();
 sg13g2_decap_8 FILLER_8_1939 ();
 sg13g2_decap_8 FILLER_8_1946 ();
 sg13g2_decap_8 FILLER_8_1953 ();
 sg13g2_decap_8 FILLER_8_1960 ();
 sg13g2_decap_8 FILLER_8_1967 ();
 sg13g2_decap_8 FILLER_8_1974 ();
 sg13g2_decap_8 FILLER_8_1981 ();
 sg13g2_decap_8 FILLER_8_1988 ();
 sg13g2_decap_8 FILLER_8_1995 ();
 sg13g2_decap_8 FILLER_8_2002 ();
 sg13g2_decap_8 FILLER_8_2009 ();
 sg13g2_decap_8 FILLER_8_2016 ();
 sg13g2_decap_8 FILLER_8_2023 ();
 sg13g2_decap_8 FILLER_8_2030 ();
 sg13g2_decap_8 FILLER_8_2037 ();
 sg13g2_decap_8 FILLER_8_2044 ();
 sg13g2_decap_8 FILLER_8_2051 ();
 sg13g2_decap_8 FILLER_8_2058 ();
 sg13g2_decap_8 FILLER_8_2065 ();
 sg13g2_decap_8 FILLER_8_2072 ();
 sg13g2_decap_8 FILLER_8_2079 ();
 sg13g2_decap_8 FILLER_8_2086 ();
 sg13g2_decap_8 FILLER_8_2093 ();
 sg13g2_decap_8 FILLER_8_2100 ();
 sg13g2_decap_8 FILLER_8_2107 ();
 sg13g2_decap_8 FILLER_8_2114 ();
 sg13g2_decap_8 FILLER_8_2121 ();
 sg13g2_decap_8 FILLER_8_2128 ();
 sg13g2_decap_8 FILLER_8_2135 ();
 sg13g2_decap_8 FILLER_8_2142 ();
 sg13g2_decap_8 FILLER_8_2149 ();
 sg13g2_decap_8 FILLER_8_2156 ();
 sg13g2_decap_8 FILLER_8_2163 ();
 sg13g2_decap_8 FILLER_8_2170 ();
 sg13g2_decap_8 FILLER_8_2177 ();
 sg13g2_decap_8 FILLER_8_2184 ();
 sg13g2_decap_8 FILLER_8_2191 ();
 sg13g2_decap_8 FILLER_8_2198 ();
 sg13g2_decap_8 FILLER_8_2205 ();
 sg13g2_decap_8 FILLER_8_2212 ();
 sg13g2_decap_8 FILLER_8_2219 ();
 sg13g2_decap_8 FILLER_8_2226 ();
 sg13g2_decap_8 FILLER_8_2233 ();
 sg13g2_decap_8 FILLER_8_2240 ();
 sg13g2_decap_8 FILLER_8_2247 ();
 sg13g2_decap_8 FILLER_8_2254 ();
 sg13g2_decap_8 FILLER_8_2261 ();
 sg13g2_decap_8 FILLER_8_2268 ();
 sg13g2_decap_8 FILLER_8_2275 ();
 sg13g2_decap_8 FILLER_8_2282 ();
 sg13g2_decap_8 FILLER_8_2289 ();
 sg13g2_decap_8 FILLER_8_2296 ();
 sg13g2_decap_8 FILLER_8_2303 ();
 sg13g2_decap_8 FILLER_8_2310 ();
 sg13g2_decap_8 FILLER_8_2317 ();
 sg13g2_decap_8 FILLER_8_2324 ();
 sg13g2_decap_8 FILLER_8_2331 ();
 sg13g2_decap_8 FILLER_8_2338 ();
 sg13g2_decap_8 FILLER_8_2345 ();
 sg13g2_decap_8 FILLER_8_2352 ();
 sg13g2_decap_8 FILLER_8_2359 ();
 sg13g2_decap_8 FILLER_8_2366 ();
 sg13g2_decap_8 FILLER_8_2373 ();
 sg13g2_decap_8 FILLER_8_2380 ();
 sg13g2_decap_8 FILLER_8_2387 ();
 sg13g2_decap_8 FILLER_8_2394 ();
 sg13g2_decap_8 FILLER_8_2401 ();
 sg13g2_decap_8 FILLER_8_2408 ();
 sg13g2_decap_8 FILLER_8_2415 ();
 sg13g2_decap_8 FILLER_8_2422 ();
 sg13g2_decap_8 FILLER_8_2429 ();
 sg13g2_decap_8 FILLER_8_2436 ();
 sg13g2_decap_8 FILLER_8_2443 ();
 sg13g2_decap_8 FILLER_8_2450 ();
 sg13g2_decap_8 FILLER_8_2457 ();
 sg13g2_decap_8 FILLER_8_2464 ();
 sg13g2_decap_8 FILLER_8_2471 ();
 sg13g2_decap_8 FILLER_8_2478 ();
 sg13g2_decap_8 FILLER_8_2485 ();
 sg13g2_decap_8 FILLER_8_2492 ();
 sg13g2_decap_8 FILLER_8_2499 ();
 sg13g2_decap_8 FILLER_8_2506 ();
 sg13g2_decap_8 FILLER_8_2513 ();
 sg13g2_decap_8 FILLER_8_2520 ();
 sg13g2_decap_8 FILLER_8_2527 ();
 sg13g2_decap_8 FILLER_8_2534 ();
 sg13g2_decap_8 FILLER_8_2541 ();
 sg13g2_decap_8 FILLER_8_2548 ();
 sg13g2_decap_8 FILLER_8_2555 ();
 sg13g2_decap_8 FILLER_8_2562 ();
 sg13g2_decap_8 FILLER_8_2569 ();
 sg13g2_decap_8 FILLER_8_2576 ();
 sg13g2_decap_8 FILLER_8_2583 ();
 sg13g2_decap_8 FILLER_8_2590 ();
 sg13g2_decap_8 FILLER_8_2597 ();
 sg13g2_decap_8 FILLER_8_2604 ();
 sg13g2_decap_8 FILLER_8_2611 ();
 sg13g2_decap_8 FILLER_8_2618 ();
 sg13g2_decap_8 FILLER_8_2625 ();
 sg13g2_decap_8 FILLER_8_2632 ();
 sg13g2_decap_8 FILLER_8_2639 ();
 sg13g2_decap_8 FILLER_8_2646 ();
 sg13g2_decap_8 FILLER_8_2653 ();
 sg13g2_decap_8 FILLER_8_2660 ();
 sg13g2_decap_8 FILLER_8_2667 ();
 sg13g2_decap_8 FILLER_8_2674 ();
 sg13g2_decap_8 FILLER_8_2681 ();
 sg13g2_decap_8 FILLER_8_2688 ();
 sg13g2_decap_8 FILLER_8_2695 ();
 sg13g2_decap_8 FILLER_8_2702 ();
 sg13g2_decap_8 FILLER_8_2709 ();
 sg13g2_decap_8 FILLER_8_2716 ();
 sg13g2_decap_8 FILLER_8_2723 ();
 sg13g2_decap_8 FILLER_8_2730 ();
 sg13g2_decap_8 FILLER_8_2737 ();
 sg13g2_decap_8 FILLER_8_2744 ();
 sg13g2_decap_8 FILLER_8_2751 ();
 sg13g2_decap_8 FILLER_8_2758 ();
 sg13g2_decap_8 FILLER_8_2765 ();
 sg13g2_decap_8 FILLER_8_2772 ();
 sg13g2_decap_8 FILLER_8_2779 ();
 sg13g2_decap_8 FILLER_8_2786 ();
 sg13g2_decap_8 FILLER_8_2793 ();
 sg13g2_decap_8 FILLER_8_2800 ();
 sg13g2_decap_8 FILLER_8_2807 ();
 sg13g2_decap_8 FILLER_8_2814 ();
 sg13g2_decap_8 FILLER_8_2821 ();
 sg13g2_decap_8 FILLER_8_2828 ();
 sg13g2_decap_8 FILLER_8_2835 ();
 sg13g2_decap_8 FILLER_8_2842 ();
 sg13g2_decap_8 FILLER_8_2849 ();
 sg13g2_decap_8 FILLER_8_2856 ();
 sg13g2_decap_8 FILLER_8_2863 ();
 sg13g2_decap_8 FILLER_8_2870 ();
 sg13g2_decap_8 FILLER_8_2877 ();
 sg13g2_decap_8 FILLER_8_2884 ();
 sg13g2_decap_8 FILLER_8_2891 ();
 sg13g2_decap_8 FILLER_8_2898 ();
 sg13g2_decap_8 FILLER_8_2905 ();
 sg13g2_decap_8 FILLER_8_2912 ();
 sg13g2_decap_8 FILLER_8_2919 ();
 sg13g2_decap_8 FILLER_8_2926 ();
 sg13g2_decap_8 FILLER_8_2933 ();
 sg13g2_decap_8 FILLER_8_2940 ();
 sg13g2_decap_8 FILLER_8_2947 ();
 sg13g2_decap_8 FILLER_8_2954 ();
 sg13g2_decap_8 FILLER_8_2961 ();
 sg13g2_decap_8 FILLER_8_2968 ();
 sg13g2_decap_8 FILLER_8_2975 ();
 sg13g2_decap_8 FILLER_8_2982 ();
 sg13g2_decap_8 FILLER_8_2989 ();
 sg13g2_decap_8 FILLER_8_2996 ();
 sg13g2_decap_8 FILLER_8_3003 ();
 sg13g2_decap_8 FILLER_8_3010 ();
 sg13g2_decap_8 FILLER_8_3017 ();
 sg13g2_decap_8 FILLER_8_3024 ();
 sg13g2_decap_8 FILLER_8_3031 ();
 sg13g2_decap_8 FILLER_8_3038 ();
 sg13g2_decap_8 FILLER_8_3045 ();
 sg13g2_decap_8 FILLER_8_3052 ();
 sg13g2_decap_8 FILLER_8_3059 ();
 sg13g2_decap_8 FILLER_8_3066 ();
 sg13g2_decap_8 FILLER_8_3073 ();
 sg13g2_decap_8 FILLER_8_3080 ();
 sg13g2_decap_8 FILLER_8_3087 ();
 sg13g2_decap_8 FILLER_8_3094 ();
 sg13g2_decap_8 FILLER_8_3101 ();
 sg13g2_decap_8 FILLER_8_3108 ();
 sg13g2_decap_8 FILLER_8_3115 ();
 sg13g2_decap_8 FILLER_8_3122 ();
 sg13g2_decap_8 FILLER_8_3129 ();
 sg13g2_decap_8 FILLER_8_3136 ();
 sg13g2_decap_8 FILLER_8_3143 ();
 sg13g2_decap_8 FILLER_8_3150 ();
 sg13g2_decap_8 FILLER_8_3157 ();
 sg13g2_decap_8 FILLER_8_3164 ();
 sg13g2_decap_8 FILLER_8_3171 ();
 sg13g2_decap_8 FILLER_8_3178 ();
 sg13g2_decap_8 FILLER_8_3185 ();
 sg13g2_decap_8 FILLER_8_3192 ();
 sg13g2_decap_8 FILLER_8_3199 ();
 sg13g2_decap_8 FILLER_8_3206 ();
 sg13g2_decap_8 FILLER_8_3213 ();
 sg13g2_decap_8 FILLER_8_3220 ();
 sg13g2_decap_8 FILLER_8_3227 ();
 sg13g2_decap_8 FILLER_8_3234 ();
 sg13g2_decap_8 FILLER_8_3241 ();
 sg13g2_decap_8 FILLER_8_3248 ();
 sg13g2_decap_8 FILLER_8_3255 ();
 sg13g2_decap_8 FILLER_8_3262 ();
 sg13g2_decap_8 FILLER_8_3269 ();
 sg13g2_decap_8 FILLER_8_3276 ();
 sg13g2_decap_8 FILLER_8_3283 ();
 sg13g2_decap_8 FILLER_8_3290 ();
 sg13g2_decap_8 FILLER_8_3297 ();
 sg13g2_decap_8 FILLER_8_3304 ();
 sg13g2_decap_8 FILLER_8_3311 ();
 sg13g2_decap_8 FILLER_8_3318 ();
 sg13g2_decap_8 FILLER_8_3325 ();
 sg13g2_decap_8 FILLER_8_3332 ();
 sg13g2_decap_8 FILLER_8_3339 ();
 sg13g2_decap_8 FILLER_8_3346 ();
 sg13g2_decap_8 FILLER_8_3353 ();
 sg13g2_decap_8 FILLER_8_3360 ();
 sg13g2_decap_8 FILLER_8_3367 ();
 sg13g2_decap_8 FILLER_8_3374 ();
 sg13g2_decap_8 FILLER_8_3381 ();
 sg13g2_decap_8 FILLER_8_3388 ();
 sg13g2_decap_8 FILLER_8_3395 ();
 sg13g2_decap_8 FILLER_8_3402 ();
 sg13g2_decap_8 FILLER_8_3409 ();
 sg13g2_decap_8 FILLER_8_3416 ();
 sg13g2_decap_8 FILLER_8_3423 ();
 sg13g2_decap_8 FILLER_8_3430 ();
 sg13g2_decap_8 FILLER_8_3437 ();
 sg13g2_decap_8 FILLER_8_3444 ();
 sg13g2_decap_8 FILLER_8_3451 ();
 sg13g2_decap_8 FILLER_8_3458 ();
 sg13g2_decap_8 FILLER_8_3465 ();
 sg13g2_decap_8 FILLER_8_3472 ();
 sg13g2_decap_8 FILLER_8_3479 ();
 sg13g2_decap_8 FILLER_8_3486 ();
 sg13g2_decap_8 FILLER_8_3493 ();
 sg13g2_decap_8 FILLER_8_3500 ();
 sg13g2_decap_8 FILLER_8_3507 ();
 sg13g2_decap_8 FILLER_8_3514 ();
 sg13g2_decap_8 FILLER_8_3521 ();
 sg13g2_decap_8 FILLER_8_3528 ();
 sg13g2_decap_8 FILLER_8_3535 ();
 sg13g2_decap_8 FILLER_8_3542 ();
 sg13g2_decap_8 FILLER_8_3549 ();
 sg13g2_decap_8 FILLER_8_3556 ();
 sg13g2_decap_8 FILLER_8_3563 ();
 sg13g2_decap_8 FILLER_8_3570 ();
 sg13g2_fill_2 FILLER_8_3577 ();
 sg13g2_fill_1 FILLER_8_3579 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_decap_8 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_9_868 ();
 sg13g2_decap_8 FILLER_9_875 ();
 sg13g2_decap_8 FILLER_9_882 ();
 sg13g2_decap_8 FILLER_9_889 ();
 sg13g2_decap_8 FILLER_9_896 ();
 sg13g2_decap_8 FILLER_9_903 ();
 sg13g2_decap_8 FILLER_9_910 ();
 sg13g2_decap_8 FILLER_9_917 ();
 sg13g2_decap_8 FILLER_9_924 ();
 sg13g2_decap_8 FILLER_9_931 ();
 sg13g2_decap_8 FILLER_9_938 ();
 sg13g2_decap_8 FILLER_9_945 ();
 sg13g2_decap_8 FILLER_9_952 ();
 sg13g2_decap_8 FILLER_9_959 ();
 sg13g2_decap_8 FILLER_9_966 ();
 sg13g2_decap_8 FILLER_9_973 ();
 sg13g2_decap_8 FILLER_9_980 ();
 sg13g2_decap_8 FILLER_9_987 ();
 sg13g2_decap_8 FILLER_9_994 ();
 sg13g2_decap_8 FILLER_9_1001 ();
 sg13g2_decap_8 FILLER_9_1008 ();
 sg13g2_decap_8 FILLER_9_1015 ();
 sg13g2_decap_8 FILLER_9_1022 ();
 sg13g2_decap_8 FILLER_9_1029 ();
 sg13g2_decap_8 FILLER_9_1036 ();
 sg13g2_decap_8 FILLER_9_1043 ();
 sg13g2_decap_8 FILLER_9_1050 ();
 sg13g2_decap_8 FILLER_9_1057 ();
 sg13g2_decap_8 FILLER_9_1064 ();
 sg13g2_decap_8 FILLER_9_1071 ();
 sg13g2_decap_8 FILLER_9_1078 ();
 sg13g2_decap_8 FILLER_9_1085 ();
 sg13g2_decap_8 FILLER_9_1092 ();
 sg13g2_decap_8 FILLER_9_1099 ();
 sg13g2_decap_8 FILLER_9_1106 ();
 sg13g2_decap_8 FILLER_9_1113 ();
 sg13g2_decap_8 FILLER_9_1120 ();
 sg13g2_decap_8 FILLER_9_1127 ();
 sg13g2_decap_8 FILLER_9_1134 ();
 sg13g2_decap_8 FILLER_9_1141 ();
 sg13g2_decap_8 FILLER_9_1148 ();
 sg13g2_decap_8 FILLER_9_1155 ();
 sg13g2_decap_8 FILLER_9_1162 ();
 sg13g2_decap_8 FILLER_9_1169 ();
 sg13g2_decap_8 FILLER_9_1176 ();
 sg13g2_decap_8 FILLER_9_1183 ();
 sg13g2_decap_8 FILLER_9_1190 ();
 sg13g2_decap_8 FILLER_9_1197 ();
 sg13g2_decap_8 FILLER_9_1204 ();
 sg13g2_decap_8 FILLER_9_1211 ();
 sg13g2_decap_8 FILLER_9_1218 ();
 sg13g2_decap_8 FILLER_9_1225 ();
 sg13g2_decap_8 FILLER_9_1232 ();
 sg13g2_decap_8 FILLER_9_1239 ();
 sg13g2_decap_8 FILLER_9_1246 ();
 sg13g2_decap_8 FILLER_9_1253 ();
 sg13g2_decap_8 FILLER_9_1260 ();
 sg13g2_decap_8 FILLER_9_1267 ();
 sg13g2_decap_8 FILLER_9_1274 ();
 sg13g2_decap_8 FILLER_9_1281 ();
 sg13g2_decap_8 FILLER_9_1288 ();
 sg13g2_decap_8 FILLER_9_1295 ();
 sg13g2_decap_8 FILLER_9_1302 ();
 sg13g2_decap_8 FILLER_9_1309 ();
 sg13g2_decap_8 FILLER_9_1316 ();
 sg13g2_decap_8 FILLER_9_1323 ();
 sg13g2_decap_8 FILLER_9_1330 ();
 sg13g2_decap_8 FILLER_9_1337 ();
 sg13g2_decap_8 FILLER_9_1344 ();
 sg13g2_decap_8 FILLER_9_1351 ();
 sg13g2_decap_8 FILLER_9_1358 ();
 sg13g2_decap_8 FILLER_9_1365 ();
 sg13g2_decap_8 FILLER_9_1372 ();
 sg13g2_decap_8 FILLER_9_1379 ();
 sg13g2_decap_8 FILLER_9_1386 ();
 sg13g2_decap_8 FILLER_9_1393 ();
 sg13g2_decap_8 FILLER_9_1400 ();
 sg13g2_decap_8 FILLER_9_1407 ();
 sg13g2_decap_8 FILLER_9_1414 ();
 sg13g2_decap_8 FILLER_9_1421 ();
 sg13g2_decap_8 FILLER_9_1428 ();
 sg13g2_decap_8 FILLER_9_1435 ();
 sg13g2_decap_8 FILLER_9_1442 ();
 sg13g2_decap_8 FILLER_9_1449 ();
 sg13g2_decap_8 FILLER_9_1456 ();
 sg13g2_decap_8 FILLER_9_1463 ();
 sg13g2_decap_8 FILLER_9_1470 ();
 sg13g2_decap_8 FILLER_9_1477 ();
 sg13g2_decap_8 FILLER_9_1484 ();
 sg13g2_decap_8 FILLER_9_1491 ();
 sg13g2_decap_8 FILLER_9_1498 ();
 sg13g2_decap_8 FILLER_9_1505 ();
 sg13g2_decap_8 FILLER_9_1512 ();
 sg13g2_decap_8 FILLER_9_1519 ();
 sg13g2_decap_8 FILLER_9_1526 ();
 sg13g2_decap_8 FILLER_9_1533 ();
 sg13g2_decap_8 FILLER_9_1540 ();
 sg13g2_decap_8 FILLER_9_1547 ();
 sg13g2_decap_8 FILLER_9_1554 ();
 sg13g2_decap_8 FILLER_9_1561 ();
 sg13g2_decap_8 FILLER_9_1568 ();
 sg13g2_decap_8 FILLER_9_1575 ();
 sg13g2_decap_8 FILLER_9_1582 ();
 sg13g2_decap_8 FILLER_9_1589 ();
 sg13g2_decap_8 FILLER_9_1596 ();
 sg13g2_decap_8 FILLER_9_1603 ();
 sg13g2_decap_8 FILLER_9_1610 ();
 sg13g2_decap_8 FILLER_9_1617 ();
 sg13g2_decap_8 FILLER_9_1624 ();
 sg13g2_decap_8 FILLER_9_1631 ();
 sg13g2_decap_8 FILLER_9_1638 ();
 sg13g2_decap_8 FILLER_9_1645 ();
 sg13g2_decap_8 FILLER_9_1652 ();
 sg13g2_decap_8 FILLER_9_1659 ();
 sg13g2_decap_8 FILLER_9_1666 ();
 sg13g2_decap_8 FILLER_9_1673 ();
 sg13g2_decap_8 FILLER_9_1680 ();
 sg13g2_decap_8 FILLER_9_1687 ();
 sg13g2_decap_8 FILLER_9_1694 ();
 sg13g2_decap_8 FILLER_9_1701 ();
 sg13g2_decap_8 FILLER_9_1708 ();
 sg13g2_decap_8 FILLER_9_1715 ();
 sg13g2_decap_8 FILLER_9_1722 ();
 sg13g2_decap_8 FILLER_9_1729 ();
 sg13g2_decap_8 FILLER_9_1736 ();
 sg13g2_decap_8 FILLER_9_1743 ();
 sg13g2_decap_8 FILLER_9_1750 ();
 sg13g2_decap_8 FILLER_9_1757 ();
 sg13g2_decap_8 FILLER_9_1764 ();
 sg13g2_decap_8 FILLER_9_1771 ();
 sg13g2_decap_8 FILLER_9_1778 ();
 sg13g2_decap_8 FILLER_9_1785 ();
 sg13g2_decap_8 FILLER_9_1792 ();
 sg13g2_decap_8 FILLER_9_1799 ();
 sg13g2_decap_8 FILLER_9_1806 ();
 sg13g2_decap_8 FILLER_9_1813 ();
 sg13g2_decap_8 FILLER_9_1820 ();
 sg13g2_decap_8 FILLER_9_1827 ();
 sg13g2_decap_8 FILLER_9_1834 ();
 sg13g2_decap_8 FILLER_9_1841 ();
 sg13g2_decap_8 FILLER_9_1848 ();
 sg13g2_decap_8 FILLER_9_1855 ();
 sg13g2_decap_8 FILLER_9_1862 ();
 sg13g2_decap_8 FILLER_9_1869 ();
 sg13g2_decap_8 FILLER_9_1876 ();
 sg13g2_decap_8 FILLER_9_1883 ();
 sg13g2_decap_8 FILLER_9_1890 ();
 sg13g2_decap_8 FILLER_9_1897 ();
 sg13g2_decap_8 FILLER_9_1904 ();
 sg13g2_decap_8 FILLER_9_1911 ();
 sg13g2_decap_8 FILLER_9_1918 ();
 sg13g2_decap_8 FILLER_9_1925 ();
 sg13g2_decap_8 FILLER_9_1932 ();
 sg13g2_decap_8 FILLER_9_1939 ();
 sg13g2_decap_8 FILLER_9_1946 ();
 sg13g2_decap_8 FILLER_9_1953 ();
 sg13g2_decap_8 FILLER_9_1960 ();
 sg13g2_decap_8 FILLER_9_1967 ();
 sg13g2_decap_8 FILLER_9_1974 ();
 sg13g2_decap_8 FILLER_9_1981 ();
 sg13g2_decap_8 FILLER_9_1988 ();
 sg13g2_decap_8 FILLER_9_1995 ();
 sg13g2_decap_8 FILLER_9_2002 ();
 sg13g2_decap_8 FILLER_9_2009 ();
 sg13g2_decap_8 FILLER_9_2016 ();
 sg13g2_decap_8 FILLER_9_2023 ();
 sg13g2_decap_8 FILLER_9_2030 ();
 sg13g2_decap_8 FILLER_9_2037 ();
 sg13g2_decap_8 FILLER_9_2044 ();
 sg13g2_decap_8 FILLER_9_2051 ();
 sg13g2_decap_8 FILLER_9_2058 ();
 sg13g2_decap_8 FILLER_9_2065 ();
 sg13g2_decap_8 FILLER_9_2072 ();
 sg13g2_decap_8 FILLER_9_2079 ();
 sg13g2_decap_8 FILLER_9_2086 ();
 sg13g2_decap_8 FILLER_9_2093 ();
 sg13g2_decap_8 FILLER_9_2100 ();
 sg13g2_decap_8 FILLER_9_2107 ();
 sg13g2_decap_8 FILLER_9_2114 ();
 sg13g2_decap_8 FILLER_9_2121 ();
 sg13g2_decap_8 FILLER_9_2128 ();
 sg13g2_decap_8 FILLER_9_2135 ();
 sg13g2_decap_8 FILLER_9_2142 ();
 sg13g2_decap_8 FILLER_9_2149 ();
 sg13g2_decap_8 FILLER_9_2156 ();
 sg13g2_decap_8 FILLER_9_2163 ();
 sg13g2_decap_8 FILLER_9_2170 ();
 sg13g2_decap_8 FILLER_9_2177 ();
 sg13g2_decap_8 FILLER_9_2184 ();
 sg13g2_decap_8 FILLER_9_2191 ();
 sg13g2_decap_8 FILLER_9_2198 ();
 sg13g2_decap_8 FILLER_9_2205 ();
 sg13g2_decap_8 FILLER_9_2212 ();
 sg13g2_decap_8 FILLER_9_2219 ();
 sg13g2_decap_8 FILLER_9_2226 ();
 sg13g2_decap_8 FILLER_9_2233 ();
 sg13g2_decap_8 FILLER_9_2240 ();
 sg13g2_decap_8 FILLER_9_2247 ();
 sg13g2_decap_8 FILLER_9_2254 ();
 sg13g2_decap_8 FILLER_9_2261 ();
 sg13g2_decap_8 FILLER_9_2268 ();
 sg13g2_decap_8 FILLER_9_2275 ();
 sg13g2_decap_8 FILLER_9_2282 ();
 sg13g2_decap_8 FILLER_9_2289 ();
 sg13g2_decap_8 FILLER_9_2296 ();
 sg13g2_decap_8 FILLER_9_2303 ();
 sg13g2_decap_8 FILLER_9_2310 ();
 sg13g2_decap_8 FILLER_9_2317 ();
 sg13g2_decap_8 FILLER_9_2324 ();
 sg13g2_decap_8 FILLER_9_2331 ();
 sg13g2_decap_8 FILLER_9_2338 ();
 sg13g2_decap_8 FILLER_9_2345 ();
 sg13g2_decap_8 FILLER_9_2352 ();
 sg13g2_decap_8 FILLER_9_2359 ();
 sg13g2_decap_8 FILLER_9_2366 ();
 sg13g2_decap_8 FILLER_9_2373 ();
 sg13g2_decap_8 FILLER_9_2380 ();
 sg13g2_decap_8 FILLER_9_2387 ();
 sg13g2_decap_8 FILLER_9_2394 ();
 sg13g2_decap_8 FILLER_9_2401 ();
 sg13g2_decap_8 FILLER_9_2408 ();
 sg13g2_decap_8 FILLER_9_2415 ();
 sg13g2_decap_8 FILLER_9_2422 ();
 sg13g2_decap_8 FILLER_9_2429 ();
 sg13g2_decap_8 FILLER_9_2436 ();
 sg13g2_decap_8 FILLER_9_2443 ();
 sg13g2_decap_8 FILLER_9_2450 ();
 sg13g2_decap_8 FILLER_9_2457 ();
 sg13g2_decap_8 FILLER_9_2464 ();
 sg13g2_decap_8 FILLER_9_2471 ();
 sg13g2_decap_8 FILLER_9_2478 ();
 sg13g2_decap_8 FILLER_9_2485 ();
 sg13g2_decap_8 FILLER_9_2492 ();
 sg13g2_decap_8 FILLER_9_2499 ();
 sg13g2_decap_8 FILLER_9_2506 ();
 sg13g2_decap_8 FILLER_9_2513 ();
 sg13g2_decap_8 FILLER_9_2520 ();
 sg13g2_decap_8 FILLER_9_2527 ();
 sg13g2_decap_8 FILLER_9_2534 ();
 sg13g2_decap_8 FILLER_9_2541 ();
 sg13g2_decap_8 FILLER_9_2548 ();
 sg13g2_decap_8 FILLER_9_2555 ();
 sg13g2_decap_8 FILLER_9_2562 ();
 sg13g2_decap_8 FILLER_9_2569 ();
 sg13g2_decap_8 FILLER_9_2576 ();
 sg13g2_decap_8 FILLER_9_2583 ();
 sg13g2_decap_8 FILLER_9_2590 ();
 sg13g2_decap_8 FILLER_9_2597 ();
 sg13g2_decap_8 FILLER_9_2604 ();
 sg13g2_decap_8 FILLER_9_2611 ();
 sg13g2_decap_8 FILLER_9_2618 ();
 sg13g2_decap_8 FILLER_9_2625 ();
 sg13g2_decap_8 FILLER_9_2632 ();
 sg13g2_decap_8 FILLER_9_2639 ();
 sg13g2_decap_8 FILLER_9_2646 ();
 sg13g2_decap_8 FILLER_9_2653 ();
 sg13g2_decap_8 FILLER_9_2660 ();
 sg13g2_decap_8 FILLER_9_2667 ();
 sg13g2_decap_8 FILLER_9_2674 ();
 sg13g2_decap_8 FILLER_9_2681 ();
 sg13g2_decap_8 FILLER_9_2688 ();
 sg13g2_decap_8 FILLER_9_2695 ();
 sg13g2_decap_8 FILLER_9_2702 ();
 sg13g2_decap_8 FILLER_9_2709 ();
 sg13g2_decap_8 FILLER_9_2716 ();
 sg13g2_decap_8 FILLER_9_2723 ();
 sg13g2_decap_8 FILLER_9_2730 ();
 sg13g2_decap_8 FILLER_9_2737 ();
 sg13g2_decap_8 FILLER_9_2744 ();
 sg13g2_decap_8 FILLER_9_2751 ();
 sg13g2_decap_8 FILLER_9_2758 ();
 sg13g2_decap_8 FILLER_9_2765 ();
 sg13g2_decap_8 FILLER_9_2772 ();
 sg13g2_decap_8 FILLER_9_2779 ();
 sg13g2_decap_8 FILLER_9_2786 ();
 sg13g2_decap_8 FILLER_9_2793 ();
 sg13g2_decap_8 FILLER_9_2800 ();
 sg13g2_decap_8 FILLER_9_2807 ();
 sg13g2_decap_8 FILLER_9_2814 ();
 sg13g2_decap_8 FILLER_9_2821 ();
 sg13g2_decap_8 FILLER_9_2828 ();
 sg13g2_decap_8 FILLER_9_2835 ();
 sg13g2_decap_8 FILLER_9_2842 ();
 sg13g2_decap_8 FILLER_9_2849 ();
 sg13g2_decap_8 FILLER_9_2856 ();
 sg13g2_decap_8 FILLER_9_2863 ();
 sg13g2_decap_8 FILLER_9_2870 ();
 sg13g2_decap_8 FILLER_9_2877 ();
 sg13g2_decap_8 FILLER_9_2884 ();
 sg13g2_decap_8 FILLER_9_2891 ();
 sg13g2_decap_8 FILLER_9_2898 ();
 sg13g2_decap_8 FILLER_9_2905 ();
 sg13g2_decap_8 FILLER_9_2912 ();
 sg13g2_decap_8 FILLER_9_2919 ();
 sg13g2_decap_8 FILLER_9_2926 ();
 sg13g2_decap_8 FILLER_9_2933 ();
 sg13g2_decap_8 FILLER_9_2940 ();
 sg13g2_decap_8 FILLER_9_2947 ();
 sg13g2_decap_8 FILLER_9_2954 ();
 sg13g2_decap_8 FILLER_9_2961 ();
 sg13g2_decap_8 FILLER_9_2968 ();
 sg13g2_decap_8 FILLER_9_2975 ();
 sg13g2_decap_8 FILLER_9_2982 ();
 sg13g2_decap_8 FILLER_9_2989 ();
 sg13g2_decap_8 FILLER_9_2996 ();
 sg13g2_decap_8 FILLER_9_3003 ();
 sg13g2_decap_8 FILLER_9_3010 ();
 sg13g2_decap_8 FILLER_9_3017 ();
 sg13g2_decap_8 FILLER_9_3024 ();
 sg13g2_decap_8 FILLER_9_3031 ();
 sg13g2_decap_8 FILLER_9_3038 ();
 sg13g2_decap_8 FILLER_9_3045 ();
 sg13g2_decap_8 FILLER_9_3052 ();
 sg13g2_decap_8 FILLER_9_3059 ();
 sg13g2_decap_8 FILLER_9_3066 ();
 sg13g2_decap_8 FILLER_9_3073 ();
 sg13g2_decap_8 FILLER_9_3080 ();
 sg13g2_decap_8 FILLER_9_3087 ();
 sg13g2_decap_8 FILLER_9_3094 ();
 sg13g2_decap_8 FILLER_9_3101 ();
 sg13g2_decap_8 FILLER_9_3108 ();
 sg13g2_decap_8 FILLER_9_3115 ();
 sg13g2_decap_8 FILLER_9_3122 ();
 sg13g2_decap_8 FILLER_9_3129 ();
 sg13g2_decap_8 FILLER_9_3136 ();
 sg13g2_decap_8 FILLER_9_3143 ();
 sg13g2_decap_8 FILLER_9_3150 ();
 sg13g2_decap_8 FILLER_9_3157 ();
 sg13g2_decap_8 FILLER_9_3164 ();
 sg13g2_decap_8 FILLER_9_3171 ();
 sg13g2_decap_8 FILLER_9_3178 ();
 sg13g2_decap_8 FILLER_9_3185 ();
 sg13g2_decap_8 FILLER_9_3192 ();
 sg13g2_decap_8 FILLER_9_3199 ();
 sg13g2_decap_8 FILLER_9_3206 ();
 sg13g2_decap_8 FILLER_9_3213 ();
 sg13g2_decap_8 FILLER_9_3220 ();
 sg13g2_decap_8 FILLER_9_3227 ();
 sg13g2_decap_8 FILLER_9_3234 ();
 sg13g2_decap_8 FILLER_9_3241 ();
 sg13g2_decap_8 FILLER_9_3248 ();
 sg13g2_decap_8 FILLER_9_3255 ();
 sg13g2_decap_8 FILLER_9_3262 ();
 sg13g2_decap_8 FILLER_9_3269 ();
 sg13g2_decap_8 FILLER_9_3276 ();
 sg13g2_decap_8 FILLER_9_3283 ();
 sg13g2_decap_8 FILLER_9_3290 ();
 sg13g2_decap_8 FILLER_9_3297 ();
 sg13g2_decap_8 FILLER_9_3304 ();
 sg13g2_decap_8 FILLER_9_3311 ();
 sg13g2_decap_8 FILLER_9_3318 ();
 sg13g2_decap_8 FILLER_9_3325 ();
 sg13g2_decap_8 FILLER_9_3332 ();
 sg13g2_decap_8 FILLER_9_3339 ();
 sg13g2_decap_8 FILLER_9_3346 ();
 sg13g2_decap_8 FILLER_9_3353 ();
 sg13g2_decap_8 FILLER_9_3360 ();
 sg13g2_decap_8 FILLER_9_3367 ();
 sg13g2_decap_8 FILLER_9_3374 ();
 sg13g2_decap_8 FILLER_9_3381 ();
 sg13g2_decap_8 FILLER_9_3388 ();
 sg13g2_decap_8 FILLER_9_3395 ();
 sg13g2_decap_8 FILLER_9_3402 ();
 sg13g2_decap_8 FILLER_9_3409 ();
 sg13g2_decap_8 FILLER_9_3416 ();
 sg13g2_decap_8 FILLER_9_3423 ();
 sg13g2_decap_8 FILLER_9_3430 ();
 sg13g2_decap_8 FILLER_9_3437 ();
 sg13g2_decap_8 FILLER_9_3444 ();
 sg13g2_decap_8 FILLER_9_3451 ();
 sg13g2_decap_8 FILLER_9_3458 ();
 sg13g2_decap_8 FILLER_9_3465 ();
 sg13g2_decap_8 FILLER_9_3472 ();
 sg13g2_decap_8 FILLER_9_3479 ();
 sg13g2_decap_8 FILLER_9_3486 ();
 sg13g2_decap_8 FILLER_9_3493 ();
 sg13g2_decap_8 FILLER_9_3500 ();
 sg13g2_decap_8 FILLER_9_3507 ();
 sg13g2_decap_8 FILLER_9_3514 ();
 sg13g2_decap_8 FILLER_9_3521 ();
 sg13g2_decap_8 FILLER_9_3528 ();
 sg13g2_decap_8 FILLER_9_3535 ();
 sg13g2_decap_8 FILLER_9_3542 ();
 sg13g2_decap_8 FILLER_9_3549 ();
 sg13g2_decap_8 FILLER_9_3556 ();
 sg13g2_decap_8 FILLER_9_3563 ();
 sg13g2_decap_8 FILLER_9_3570 ();
 sg13g2_fill_2 FILLER_9_3577 ();
 sg13g2_fill_1 FILLER_9_3579 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_decap_8 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_10_868 ();
 sg13g2_decap_8 FILLER_10_875 ();
 sg13g2_decap_8 FILLER_10_882 ();
 sg13g2_decap_8 FILLER_10_889 ();
 sg13g2_decap_8 FILLER_10_896 ();
 sg13g2_decap_8 FILLER_10_903 ();
 sg13g2_decap_8 FILLER_10_910 ();
 sg13g2_decap_8 FILLER_10_917 ();
 sg13g2_decap_8 FILLER_10_924 ();
 sg13g2_decap_8 FILLER_10_931 ();
 sg13g2_decap_8 FILLER_10_938 ();
 sg13g2_decap_8 FILLER_10_945 ();
 sg13g2_decap_8 FILLER_10_952 ();
 sg13g2_decap_8 FILLER_10_959 ();
 sg13g2_decap_8 FILLER_10_966 ();
 sg13g2_decap_8 FILLER_10_973 ();
 sg13g2_decap_8 FILLER_10_980 ();
 sg13g2_decap_8 FILLER_10_987 ();
 sg13g2_decap_8 FILLER_10_994 ();
 sg13g2_decap_8 FILLER_10_1001 ();
 sg13g2_decap_8 FILLER_10_1008 ();
 sg13g2_decap_8 FILLER_10_1015 ();
 sg13g2_decap_8 FILLER_10_1022 ();
 sg13g2_decap_8 FILLER_10_1029 ();
 sg13g2_decap_8 FILLER_10_1036 ();
 sg13g2_decap_8 FILLER_10_1043 ();
 sg13g2_decap_8 FILLER_10_1050 ();
 sg13g2_decap_8 FILLER_10_1057 ();
 sg13g2_decap_8 FILLER_10_1064 ();
 sg13g2_decap_8 FILLER_10_1071 ();
 sg13g2_decap_8 FILLER_10_1078 ();
 sg13g2_decap_8 FILLER_10_1085 ();
 sg13g2_decap_8 FILLER_10_1092 ();
 sg13g2_decap_8 FILLER_10_1099 ();
 sg13g2_decap_8 FILLER_10_1106 ();
 sg13g2_decap_8 FILLER_10_1113 ();
 sg13g2_decap_8 FILLER_10_1120 ();
 sg13g2_decap_8 FILLER_10_1127 ();
 sg13g2_decap_8 FILLER_10_1134 ();
 sg13g2_decap_8 FILLER_10_1141 ();
 sg13g2_decap_8 FILLER_10_1148 ();
 sg13g2_decap_8 FILLER_10_1155 ();
 sg13g2_decap_8 FILLER_10_1162 ();
 sg13g2_decap_8 FILLER_10_1169 ();
 sg13g2_decap_8 FILLER_10_1176 ();
 sg13g2_decap_8 FILLER_10_1183 ();
 sg13g2_decap_8 FILLER_10_1190 ();
 sg13g2_decap_8 FILLER_10_1197 ();
 sg13g2_decap_8 FILLER_10_1204 ();
 sg13g2_decap_8 FILLER_10_1211 ();
 sg13g2_decap_8 FILLER_10_1218 ();
 sg13g2_decap_8 FILLER_10_1225 ();
 sg13g2_decap_8 FILLER_10_1232 ();
 sg13g2_decap_8 FILLER_10_1239 ();
 sg13g2_decap_8 FILLER_10_1246 ();
 sg13g2_decap_8 FILLER_10_1253 ();
 sg13g2_decap_8 FILLER_10_1260 ();
 sg13g2_decap_8 FILLER_10_1267 ();
 sg13g2_decap_8 FILLER_10_1274 ();
 sg13g2_decap_8 FILLER_10_1281 ();
 sg13g2_decap_8 FILLER_10_1288 ();
 sg13g2_decap_8 FILLER_10_1295 ();
 sg13g2_decap_8 FILLER_10_1302 ();
 sg13g2_decap_8 FILLER_10_1309 ();
 sg13g2_decap_8 FILLER_10_1316 ();
 sg13g2_decap_8 FILLER_10_1323 ();
 sg13g2_decap_8 FILLER_10_1330 ();
 sg13g2_decap_8 FILLER_10_1337 ();
 sg13g2_decap_8 FILLER_10_1344 ();
 sg13g2_decap_8 FILLER_10_1351 ();
 sg13g2_decap_8 FILLER_10_1358 ();
 sg13g2_decap_8 FILLER_10_1365 ();
 sg13g2_decap_8 FILLER_10_1372 ();
 sg13g2_decap_8 FILLER_10_1379 ();
 sg13g2_decap_8 FILLER_10_1386 ();
 sg13g2_decap_8 FILLER_10_1393 ();
 sg13g2_decap_8 FILLER_10_1400 ();
 sg13g2_decap_8 FILLER_10_1407 ();
 sg13g2_decap_8 FILLER_10_1414 ();
 sg13g2_decap_8 FILLER_10_1421 ();
 sg13g2_decap_8 FILLER_10_1428 ();
 sg13g2_decap_8 FILLER_10_1435 ();
 sg13g2_decap_8 FILLER_10_1442 ();
 sg13g2_decap_8 FILLER_10_1449 ();
 sg13g2_decap_8 FILLER_10_1456 ();
 sg13g2_decap_8 FILLER_10_1463 ();
 sg13g2_decap_8 FILLER_10_1470 ();
 sg13g2_decap_8 FILLER_10_1477 ();
 sg13g2_decap_8 FILLER_10_1484 ();
 sg13g2_decap_8 FILLER_10_1491 ();
 sg13g2_decap_8 FILLER_10_1498 ();
 sg13g2_decap_8 FILLER_10_1505 ();
 sg13g2_decap_8 FILLER_10_1512 ();
 sg13g2_decap_8 FILLER_10_1519 ();
 sg13g2_decap_8 FILLER_10_1526 ();
 sg13g2_decap_8 FILLER_10_1533 ();
 sg13g2_decap_8 FILLER_10_1540 ();
 sg13g2_decap_8 FILLER_10_1547 ();
 sg13g2_decap_8 FILLER_10_1554 ();
 sg13g2_decap_8 FILLER_10_1561 ();
 sg13g2_decap_8 FILLER_10_1568 ();
 sg13g2_decap_8 FILLER_10_1575 ();
 sg13g2_decap_8 FILLER_10_1582 ();
 sg13g2_decap_8 FILLER_10_1589 ();
 sg13g2_decap_8 FILLER_10_1596 ();
 sg13g2_decap_8 FILLER_10_1603 ();
 sg13g2_decap_8 FILLER_10_1610 ();
 sg13g2_decap_8 FILLER_10_1617 ();
 sg13g2_decap_8 FILLER_10_1624 ();
 sg13g2_decap_8 FILLER_10_1631 ();
 sg13g2_decap_8 FILLER_10_1638 ();
 sg13g2_decap_8 FILLER_10_1645 ();
 sg13g2_decap_8 FILLER_10_1652 ();
 sg13g2_decap_8 FILLER_10_1659 ();
 sg13g2_decap_8 FILLER_10_1666 ();
 sg13g2_decap_8 FILLER_10_1673 ();
 sg13g2_decap_8 FILLER_10_1680 ();
 sg13g2_decap_8 FILLER_10_1687 ();
 sg13g2_decap_8 FILLER_10_1694 ();
 sg13g2_decap_8 FILLER_10_1701 ();
 sg13g2_decap_8 FILLER_10_1708 ();
 sg13g2_decap_8 FILLER_10_1715 ();
 sg13g2_decap_8 FILLER_10_1722 ();
 sg13g2_decap_8 FILLER_10_1729 ();
 sg13g2_decap_8 FILLER_10_1736 ();
 sg13g2_decap_8 FILLER_10_1743 ();
 sg13g2_decap_8 FILLER_10_1750 ();
 sg13g2_decap_8 FILLER_10_1757 ();
 sg13g2_decap_8 FILLER_10_1764 ();
 sg13g2_decap_8 FILLER_10_1771 ();
 sg13g2_decap_8 FILLER_10_1778 ();
 sg13g2_decap_8 FILLER_10_1785 ();
 sg13g2_decap_8 FILLER_10_1792 ();
 sg13g2_decap_8 FILLER_10_1799 ();
 sg13g2_decap_8 FILLER_10_1806 ();
 sg13g2_decap_8 FILLER_10_1813 ();
 sg13g2_decap_8 FILLER_10_1820 ();
 sg13g2_decap_8 FILLER_10_1827 ();
 sg13g2_decap_8 FILLER_10_1834 ();
 sg13g2_decap_8 FILLER_10_1841 ();
 sg13g2_decap_8 FILLER_10_1848 ();
 sg13g2_decap_8 FILLER_10_1855 ();
 sg13g2_decap_8 FILLER_10_1862 ();
 sg13g2_decap_8 FILLER_10_1869 ();
 sg13g2_decap_8 FILLER_10_1876 ();
 sg13g2_decap_8 FILLER_10_1883 ();
 sg13g2_decap_8 FILLER_10_1890 ();
 sg13g2_decap_8 FILLER_10_1897 ();
 sg13g2_decap_8 FILLER_10_1904 ();
 sg13g2_decap_8 FILLER_10_1911 ();
 sg13g2_decap_8 FILLER_10_1918 ();
 sg13g2_decap_8 FILLER_10_1925 ();
 sg13g2_decap_8 FILLER_10_1932 ();
 sg13g2_decap_8 FILLER_10_1939 ();
 sg13g2_decap_8 FILLER_10_1946 ();
 sg13g2_decap_8 FILLER_10_1953 ();
 sg13g2_decap_8 FILLER_10_1960 ();
 sg13g2_decap_8 FILLER_10_1967 ();
 sg13g2_decap_8 FILLER_10_1974 ();
 sg13g2_decap_8 FILLER_10_1981 ();
 sg13g2_decap_8 FILLER_10_1988 ();
 sg13g2_decap_8 FILLER_10_1995 ();
 sg13g2_decap_8 FILLER_10_2002 ();
 sg13g2_decap_8 FILLER_10_2009 ();
 sg13g2_decap_8 FILLER_10_2016 ();
 sg13g2_decap_8 FILLER_10_2023 ();
 sg13g2_decap_8 FILLER_10_2030 ();
 sg13g2_decap_8 FILLER_10_2037 ();
 sg13g2_decap_8 FILLER_10_2044 ();
 sg13g2_decap_8 FILLER_10_2051 ();
 sg13g2_decap_8 FILLER_10_2058 ();
 sg13g2_decap_8 FILLER_10_2065 ();
 sg13g2_decap_8 FILLER_10_2072 ();
 sg13g2_decap_8 FILLER_10_2079 ();
 sg13g2_decap_8 FILLER_10_2086 ();
 sg13g2_decap_8 FILLER_10_2093 ();
 sg13g2_decap_8 FILLER_10_2100 ();
 sg13g2_decap_8 FILLER_10_2107 ();
 sg13g2_decap_8 FILLER_10_2114 ();
 sg13g2_decap_8 FILLER_10_2121 ();
 sg13g2_decap_8 FILLER_10_2128 ();
 sg13g2_decap_8 FILLER_10_2135 ();
 sg13g2_decap_8 FILLER_10_2142 ();
 sg13g2_decap_8 FILLER_10_2149 ();
 sg13g2_decap_8 FILLER_10_2156 ();
 sg13g2_decap_8 FILLER_10_2163 ();
 sg13g2_decap_8 FILLER_10_2170 ();
 sg13g2_decap_8 FILLER_10_2177 ();
 sg13g2_decap_8 FILLER_10_2184 ();
 sg13g2_decap_8 FILLER_10_2191 ();
 sg13g2_decap_8 FILLER_10_2198 ();
 sg13g2_decap_8 FILLER_10_2205 ();
 sg13g2_decap_8 FILLER_10_2212 ();
 sg13g2_decap_8 FILLER_10_2219 ();
 sg13g2_decap_8 FILLER_10_2226 ();
 sg13g2_decap_8 FILLER_10_2233 ();
 sg13g2_decap_8 FILLER_10_2240 ();
 sg13g2_decap_8 FILLER_10_2247 ();
 sg13g2_decap_8 FILLER_10_2254 ();
 sg13g2_decap_8 FILLER_10_2261 ();
 sg13g2_decap_8 FILLER_10_2268 ();
 sg13g2_decap_8 FILLER_10_2275 ();
 sg13g2_decap_8 FILLER_10_2282 ();
 sg13g2_decap_8 FILLER_10_2289 ();
 sg13g2_decap_8 FILLER_10_2296 ();
 sg13g2_decap_8 FILLER_10_2303 ();
 sg13g2_decap_8 FILLER_10_2310 ();
 sg13g2_decap_8 FILLER_10_2317 ();
 sg13g2_decap_8 FILLER_10_2324 ();
 sg13g2_decap_8 FILLER_10_2331 ();
 sg13g2_decap_8 FILLER_10_2338 ();
 sg13g2_decap_8 FILLER_10_2345 ();
 sg13g2_decap_8 FILLER_10_2352 ();
 sg13g2_decap_8 FILLER_10_2359 ();
 sg13g2_decap_8 FILLER_10_2366 ();
 sg13g2_decap_8 FILLER_10_2373 ();
 sg13g2_decap_8 FILLER_10_2380 ();
 sg13g2_decap_8 FILLER_10_2387 ();
 sg13g2_decap_8 FILLER_10_2394 ();
 sg13g2_decap_8 FILLER_10_2401 ();
 sg13g2_decap_8 FILLER_10_2408 ();
 sg13g2_decap_8 FILLER_10_2415 ();
 sg13g2_decap_8 FILLER_10_2422 ();
 sg13g2_decap_8 FILLER_10_2429 ();
 sg13g2_decap_8 FILLER_10_2436 ();
 sg13g2_decap_8 FILLER_10_2443 ();
 sg13g2_decap_8 FILLER_10_2450 ();
 sg13g2_decap_8 FILLER_10_2457 ();
 sg13g2_decap_8 FILLER_10_2464 ();
 sg13g2_decap_8 FILLER_10_2471 ();
 sg13g2_decap_8 FILLER_10_2478 ();
 sg13g2_decap_8 FILLER_10_2485 ();
 sg13g2_decap_8 FILLER_10_2492 ();
 sg13g2_decap_8 FILLER_10_2499 ();
 sg13g2_decap_8 FILLER_10_2506 ();
 sg13g2_decap_8 FILLER_10_2513 ();
 sg13g2_decap_8 FILLER_10_2520 ();
 sg13g2_decap_8 FILLER_10_2527 ();
 sg13g2_decap_8 FILLER_10_2534 ();
 sg13g2_decap_8 FILLER_10_2541 ();
 sg13g2_decap_8 FILLER_10_2548 ();
 sg13g2_decap_8 FILLER_10_2555 ();
 sg13g2_decap_8 FILLER_10_2562 ();
 sg13g2_decap_8 FILLER_10_2569 ();
 sg13g2_decap_8 FILLER_10_2576 ();
 sg13g2_decap_8 FILLER_10_2583 ();
 sg13g2_decap_8 FILLER_10_2590 ();
 sg13g2_decap_8 FILLER_10_2597 ();
 sg13g2_decap_8 FILLER_10_2604 ();
 sg13g2_decap_8 FILLER_10_2611 ();
 sg13g2_decap_8 FILLER_10_2618 ();
 sg13g2_decap_8 FILLER_10_2625 ();
 sg13g2_decap_8 FILLER_10_2632 ();
 sg13g2_decap_8 FILLER_10_2639 ();
 sg13g2_decap_8 FILLER_10_2646 ();
 sg13g2_decap_8 FILLER_10_2653 ();
 sg13g2_decap_8 FILLER_10_2660 ();
 sg13g2_decap_8 FILLER_10_2667 ();
 sg13g2_decap_8 FILLER_10_2674 ();
 sg13g2_decap_8 FILLER_10_2681 ();
 sg13g2_decap_8 FILLER_10_2688 ();
 sg13g2_decap_8 FILLER_10_2695 ();
 sg13g2_decap_8 FILLER_10_2702 ();
 sg13g2_decap_8 FILLER_10_2709 ();
 sg13g2_decap_8 FILLER_10_2716 ();
 sg13g2_decap_8 FILLER_10_2723 ();
 sg13g2_decap_8 FILLER_10_2730 ();
 sg13g2_decap_8 FILLER_10_2737 ();
 sg13g2_decap_8 FILLER_10_2744 ();
 sg13g2_decap_8 FILLER_10_2751 ();
 sg13g2_decap_8 FILLER_10_2758 ();
 sg13g2_decap_8 FILLER_10_2765 ();
 sg13g2_decap_8 FILLER_10_2772 ();
 sg13g2_decap_8 FILLER_10_2779 ();
 sg13g2_decap_8 FILLER_10_2786 ();
 sg13g2_decap_8 FILLER_10_2793 ();
 sg13g2_decap_8 FILLER_10_2800 ();
 sg13g2_decap_8 FILLER_10_2807 ();
 sg13g2_decap_8 FILLER_10_2814 ();
 sg13g2_decap_8 FILLER_10_2821 ();
 sg13g2_decap_8 FILLER_10_2828 ();
 sg13g2_decap_8 FILLER_10_2835 ();
 sg13g2_decap_8 FILLER_10_2842 ();
 sg13g2_decap_8 FILLER_10_2849 ();
 sg13g2_decap_8 FILLER_10_2856 ();
 sg13g2_decap_8 FILLER_10_2863 ();
 sg13g2_decap_8 FILLER_10_2870 ();
 sg13g2_decap_8 FILLER_10_2877 ();
 sg13g2_decap_8 FILLER_10_2884 ();
 sg13g2_decap_8 FILLER_10_2891 ();
 sg13g2_decap_8 FILLER_10_2898 ();
 sg13g2_decap_8 FILLER_10_2905 ();
 sg13g2_decap_8 FILLER_10_2912 ();
 sg13g2_decap_8 FILLER_10_2919 ();
 sg13g2_decap_8 FILLER_10_2926 ();
 sg13g2_decap_8 FILLER_10_2933 ();
 sg13g2_decap_8 FILLER_10_2940 ();
 sg13g2_decap_8 FILLER_10_2947 ();
 sg13g2_decap_8 FILLER_10_2954 ();
 sg13g2_decap_8 FILLER_10_2961 ();
 sg13g2_decap_8 FILLER_10_2968 ();
 sg13g2_decap_8 FILLER_10_2975 ();
 sg13g2_decap_8 FILLER_10_2982 ();
 sg13g2_decap_8 FILLER_10_2989 ();
 sg13g2_decap_8 FILLER_10_2996 ();
 sg13g2_decap_8 FILLER_10_3003 ();
 sg13g2_decap_8 FILLER_10_3010 ();
 sg13g2_decap_8 FILLER_10_3017 ();
 sg13g2_decap_8 FILLER_10_3024 ();
 sg13g2_decap_8 FILLER_10_3031 ();
 sg13g2_decap_8 FILLER_10_3038 ();
 sg13g2_decap_8 FILLER_10_3045 ();
 sg13g2_decap_8 FILLER_10_3052 ();
 sg13g2_decap_8 FILLER_10_3059 ();
 sg13g2_decap_8 FILLER_10_3066 ();
 sg13g2_decap_8 FILLER_10_3073 ();
 sg13g2_decap_8 FILLER_10_3080 ();
 sg13g2_decap_8 FILLER_10_3087 ();
 sg13g2_decap_8 FILLER_10_3094 ();
 sg13g2_decap_8 FILLER_10_3101 ();
 sg13g2_decap_8 FILLER_10_3108 ();
 sg13g2_decap_8 FILLER_10_3115 ();
 sg13g2_decap_8 FILLER_10_3122 ();
 sg13g2_decap_8 FILLER_10_3129 ();
 sg13g2_decap_8 FILLER_10_3136 ();
 sg13g2_decap_8 FILLER_10_3143 ();
 sg13g2_decap_8 FILLER_10_3150 ();
 sg13g2_decap_8 FILLER_10_3157 ();
 sg13g2_decap_8 FILLER_10_3164 ();
 sg13g2_decap_8 FILLER_10_3171 ();
 sg13g2_decap_8 FILLER_10_3178 ();
 sg13g2_decap_8 FILLER_10_3185 ();
 sg13g2_decap_8 FILLER_10_3192 ();
 sg13g2_decap_8 FILLER_10_3199 ();
 sg13g2_decap_8 FILLER_10_3206 ();
 sg13g2_decap_8 FILLER_10_3213 ();
 sg13g2_decap_8 FILLER_10_3220 ();
 sg13g2_decap_8 FILLER_10_3227 ();
 sg13g2_decap_8 FILLER_10_3234 ();
 sg13g2_decap_8 FILLER_10_3241 ();
 sg13g2_decap_8 FILLER_10_3248 ();
 sg13g2_decap_8 FILLER_10_3255 ();
 sg13g2_decap_8 FILLER_10_3262 ();
 sg13g2_decap_8 FILLER_10_3269 ();
 sg13g2_decap_8 FILLER_10_3276 ();
 sg13g2_decap_8 FILLER_10_3283 ();
 sg13g2_decap_8 FILLER_10_3290 ();
 sg13g2_decap_8 FILLER_10_3297 ();
 sg13g2_decap_8 FILLER_10_3304 ();
 sg13g2_decap_8 FILLER_10_3311 ();
 sg13g2_decap_8 FILLER_10_3318 ();
 sg13g2_decap_8 FILLER_10_3325 ();
 sg13g2_decap_8 FILLER_10_3332 ();
 sg13g2_decap_8 FILLER_10_3339 ();
 sg13g2_decap_8 FILLER_10_3346 ();
 sg13g2_decap_8 FILLER_10_3353 ();
 sg13g2_decap_8 FILLER_10_3360 ();
 sg13g2_decap_8 FILLER_10_3367 ();
 sg13g2_decap_8 FILLER_10_3374 ();
 sg13g2_decap_8 FILLER_10_3381 ();
 sg13g2_decap_8 FILLER_10_3388 ();
 sg13g2_decap_8 FILLER_10_3395 ();
 sg13g2_decap_8 FILLER_10_3402 ();
 sg13g2_decap_8 FILLER_10_3409 ();
 sg13g2_decap_8 FILLER_10_3416 ();
 sg13g2_decap_8 FILLER_10_3423 ();
 sg13g2_decap_8 FILLER_10_3430 ();
 sg13g2_decap_8 FILLER_10_3437 ();
 sg13g2_decap_8 FILLER_10_3444 ();
 sg13g2_decap_8 FILLER_10_3451 ();
 sg13g2_decap_8 FILLER_10_3458 ();
 sg13g2_decap_8 FILLER_10_3465 ();
 sg13g2_decap_8 FILLER_10_3472 ();
 sg13g2_decap_8 FILLER_10_3479 ();
 sg13g2_decap_8 FILLER_10_3486 ();
 sg13g2_decap_8 FILLER_10_3493 ();
 sg13g2_decap_8 FILLER_10_3500 ();
 sg13g2_decap_8 FILLER_10_3507 ();
 sg13g2_decap_8 FILLER_10_3514 ();
 sg13g2_decap_8 FILLER_10_3521 ();
 sg13g2_decap_8 FILLER_10_3528 ();
 sg13g2_decap_8 FILLER_10_3535 ();
 sg13g2_decap_8 FILLER_10_3542 ();
 sg13g2_decap_8 FILLER_10_3549 ();
 sg13g2_decap_8 FILLER_10_3556 ();
 sg13g2_decap_8 FILLER_10_3563 ();
 sg13g2_decap_8 FILLER_10_3570 ();
 sg13g2_fill_2 FILLER_10_3577 ();
 sg13g2_fill_1 FILLER_10_3579 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_decap_8 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_11_868 ();
 sg13g2_decap_8 FILLER_11_875 ();
 sg13g2_decap_8 FILLER_11_882 ();
 sg13g2_decap_8 FILLER_11_889 ();
 sg13g2_decap_8 FILLER_11_896 ();
 sg13g2_decap_8 FILLER_11_903 ();
 sg13g2_decap_8 FILLER_11_910 ();
 sg13g2_decap_8 FILLER_11_917 ();
 sg13g2_decap_8 FILLER_11_924 ();
 sg13g2_decap_8 FILLER_11_931 ();
 sg13g2_decap_8 FILLER_11_938 ();
 sg13g2_decap_8 FILLER_11_945 ();
 sg13g2_decap_8 FILLER_11_952 ();
 sg13g2_decap_8 FILLER_11_959 ();
 sg13g2_decap_8 FILLER_11_966 ();
 sg13g2_decap_8 FILLER_11_973 ();
 sg13g2_decap_8 FILLER_11_980 ();
 sg13g2_decap_8 FILLER_11_987 ();
 sg13g2_decap_8 FILLER_11_994 ();
 sg13g2_decap_8 FILLER_11_1001 ();
 sg13g2_decap_8 FILLER_11_1008 ();
 sg13g2_decap_8 FILLER_11_1015 ();
 sg13g2_decap_8 FILLER_11_1022 ();
 sg13g2_decap_8 FILLER_11_1029 ();
 sg13g2_decap_8 FILLER_11_1036 ();
 sg13g2_decap_8 FILLER_11_1043 ();
 sg13g2_decap_8 FILLER_11_1050 ();
 sg13g2_decap_8 FILLER_11_1057 ();
 sg13g2_decap_8 FILLER_11_1064 ();
 sg13g2_decap_8 FILLER_11_1071 ();
 sg13g2_decap_8 FILLER_11_1078 ();
 sg13g2_decap_8 FILLER_11_1085 ();
 sg13g2_decap_8 FILLER_11_1092 ();
 sg13g2_decap_8 FILLER_11_1099 ();
 sg13g2_decap_8 FILLER_11_1106 ();
 sg13g2_decap_8 FILLER_11_1113 ();
 sg13g2_decap_8 FILLER_11_1120 ();
 sg13g2_decap_8 FILLER_11_1127 ();
 sg13g2_decap_8 FILLER_11_1134 ();
 sg13g2_decap_8 FILLER_11_1141 ();
 sg13g2_decap_8 FILLER_11_1148 ();
 sg13g2_decap_8 FILLER_11_1155 ();
 sg13g2_decap_8 FILLER_11_1162 ();
 sg13g2_decap_8 FILLER_11_1169 ();
 sg13g2_decap_8 FILLER_11_1176 ();
 sg13g2_decap_8 FILLER_11_1183 ();
 sg13g2_decap_8 FILLER_11_1190 ();
 sg13g2_decap_8 FILLER_11_1197 ();
 sg13g2_decap_8 FILLER_11_1204 ();
 sg13g2_decap_8 FILLER_11_1211 ();
 sg13g2_decap_8 FILLER_11_1218 ();
 sg13g2_decap_8 FILLER_11_1225 ();
 sg13g2_decap_8 FILLER_11_1232 ();
 sg13g2_decap_8 FILLER_11_1239 ();
 sg13g2_decap_8 FILLER_11_1246 ();
 sg13g2_decap_8 FILLER_11_1253 ();
 sg13g2_decap_8 FILLER_11_1260 ();
 sg13g2_decap_8 FILLER_11_1267 ();
 sg13g2_decap_8 FILLER_11_1274 ();
 sg13g2_decap_8 FILLER_11_1281 ();
 sg13g2_decap_8 FILLER_11_1288 ();
 sg13g2_decap_8 FILLER_11_1295 ();
 sg13g2_decap_8 FILLER_11_1302 ();
 sg13g2_decap_8 FILLER_11_1309 ();
 sg13g2_decap_8 FILLER_11_1316 ();
 sg13g2_decap_8 FILLER_11_1323 ();
 sg13g2_decap_8 FILLER_11_1330 ();
 sg13g2_decap_8 FILLER_11_1337 ();
 sg13g2_decap_8 FILLER_11_1344 ();
 sg13g2_decap_8 FILLER_11_1351 ();
 sg13g2_decap_8 FILLER_11_1358 ();
 sg13g2_decap_8 FILLER_11_1365 ();
 sg13g2_decap_8 FILLER_11_1372 ();
 sg13g2_decap_8 FILLER_11_1379 ();
 sg13g2_decap_8 FILLER_11_1386 ();
 sg13g2_decap_8 FILLER_11_1393 ();
 sg13g2_decap_8 FILLER_11_1400 ();
 sg13g2_decap_8 FILLER_11_1407 ();
 sg13g2_decap_8 FILLER_11_1414 ();
 sg13g2_decap_8 FILLER_11_1421 ();
 sg13g2_decap_8 FILLER_11_1428 ();
 sg13g2_decap_8 FILLER_11_1435 ();
 sg13g2_decap_8 FILLER_11_1442 ();
 sg13g2_decap_8 FILLER_11_1449 ();
 sg13g2_decap_8 FILLER_11_1456 ();
 sg13g2_decap_8 FILLER_11_1463 ();
 sg13g2_decap_8 FILLER_11_1470 ();
 sg13g2_decap_8 FILLER_11_1477 ();
 sg13g2_decap_8 FILLER_11_1484 ();
 sg13g2_decap_8 FILLER_11_1491 ();
 sg13g2_decap_8 FILLER_11_1498 ();
 sg13g2_decap_8 FILLER_11_1505 ();
 sg13g2_decap_8 FILLER_11_1512 ();
 sg13g2_decap_8 FILLER_11_1519 ();
 sg13g2_decap_8 FILLER_11_1526 ();
 sg13g2_decap_8 FILLER_11_1533 ();
 sg13g2_decap_8 FILLER_11_1540 ();
 sg13g2_decap_8 FILLER_11_1547 ();
 sg13g2_decap_8 FILLER_11_1554 ();
 sg13g2_decap_8 FILLER_11_1561 ();
 sg13g2_decap_8 FILLER_11_1568 ();
 sg13g2_decap_8 FILLER_11_1575 ();
 sg13g2_decap_8 FILLER_11_1582 ();
 sg13g2_decap_8 FILLER_11_1589 ();
 sg13g2_decap_8 FILLER_11_1596 ();
 sg13g2_decap_8 FILLER_11_1603 ();
 sg13g2_decap_8 FILLER_11_1610 ();
 sg13g2_decap_8 FILLER_11_1617 ();
 sg13g2_decap_8 FILLER_11_1624 ();
 sg13g2_decap_8 FILLER_11_1631 ();
 sg13g2_decap_8 FILLER_11_1638 ();
 sg13g2_decap_8 FILLER_11_1645 ();
 sg13g2_decap_8 FILLER_11_1652 ();
 sg13g2_decap_8 FILLER_11_1659 ();
 sg13g2_decap_8 FILLER_11_1666 ();
 sg13g2_decap_8 FILLER_11_1673 ();
 sg13g2_decap_8 FILLER_11_1680 ();
 sg13g2_decap_8 FILLER_11_1687 ();
 sg13g2_decap_8 FILLER_11_1694 ();
 sg13g2_decap_8 FILLER_11_1701 ();
 sg13g2_decap_8 FILLER_11_1708 ();
 sg13g2_decap_8 FILLER_11_1715 ();
 sg13g2_decap_8 FILLER_11_1722 ();
 sg13g2_decap_8 FILLER_11_1729 ();
 sg13g2_decap_8 FILLER_11_1736 ();
 sg13g2_decap_8 FILLER_11_1743 ();
 sg13g2_decap_8 FILLER_11_1750 ();
 sg13g2_decap_8 FILLER_11_1757 ();
 sg13g2_decap_8 FILLER_11_1764 ();
 sg13g2_decap_8 FILLER_11_1771 ();
 sg13g2_decap_8 FILLER_11_1778 ();
 sg13g2_decap_8 FILLER_11_1785 ();
 sg13g2_decap_8 FILLER_11_1792 ();
 sg13g2_decap_8 FILLER_11_1799 ();
 sg13g2_decap_8 FILLER_11_1806 ();
 sg13g2_decap_8 FILLER_11_1813 ();
 sg13g2_decap_8 FILLER_11_1820 ();
 sg13g2_decap_8 FILLER_11_1827 ();
 sg13g2_decap_8 FILLER_11_1834 ();
 sg13g2_decap_8 FILLER_11_1841 ();
 sg13g2_decap_8 FILLER_11_1848 ();
 sg13g2_decap_8 FILLER_11_1855 ();
 sg13g2_decap_8 FILLER_11_1862 ();
 sg13g2_decap_8 FILLER_11_1869 ();
 sg13g2_decap_8 FILLER_11_1876 ();
 sg13g2_decap_8 FILLER_11_1883 ();
 sg13g2_decap_8 FILLER_11_1890 ();
 sg13g2_decap_8 FILLER_11_1897 ();
 sg13g2_decap_8 FILLER_11_1904 ();
 sg13g2_decap_8 FILLER_11_1911 ();
 sg13g2_decap_8 FILLER_11_1918 ();
 sg13g2_decap_8 FILLER_11_1925 ();
 sg13g2_decap_8 FILLER_11_1932 ();
 sg13g2_decap_8 FILLER_11_1939 ();
 sg13g2_decap_8 FILLER_11_1946 ();
 sg13g2_decap_8 FILLER_11_1953 ();
 sg13g2_decap_8 FILLER_11_1960 ();
 sg13g2_decap_8 FILLER_11_1967 ();
 sg13g2_decap_8 FILLER_11_1974 ();
 sg13g2_decap_8 FILLER_11_1981 ();
 sg13g2_decap_8 FILLER_11_1988 ();
 sg13g2_decap_8 FILLER_11_1995 ();
 sg13g2_decap_8 FILLER_11_2002 ();
 sg13g2_decap_8 FILLER_11_2009 ();
 sg13g2_decap_8 FILLER_11_2016 ();
 sg13g2_decap_8 FILLER_11_2023 ();
 sg13g2_decap_8 FILLER_11_2030 ();
 sg13g2_decap_8 FILLER_11_2037 ();
 sg13g2_decap_8 FILLER_11_2044 ();
 sg13g2_decap_8 FILLER_11_2051 ();
 sg13g2_decap_8 FILLER_11_2058 ();
 sg13g2_decap_8 FILLER_11_2065 ();
 sg13g2_decap_8 FILLER_11_2072 ();
 sg13g2_decap_8 FILLER_11_2079 ();
 sg13g2_decap_8 FILLER_11_2086 ();
 sg13g2_decap_8 FILLER_11_2093 ();
 sg13g2_decap_8 FILLER_11_2100 ();
 sg13g2_decap_8 FILLER_11_2107 ();
 sg13g2_decap_8 FILLER_11_2114 ();
 sg13g2_decap_8 FILLER_11_2121 ();
 sg13g2_decap_8 FILLER_11_2128 ();
 sg13g2_decap_8 FILLER_11_2135 ();
 sg13g2_decap_8 FILLER_11_2142 ();
 sg13g2_decap_8 FILLER_11_2149 ();
 sg13g2_decap_8 FILLER_11_2156 ();
 sg13g2_decap_8 FILLER_11_2163 ();
 sg13g2_decap_8 FILLER_11_2170 ();
 sg13g2_decap_8 FILLER_11_2177 ();
 sg13g2_decap_8 FILLER_11_2184 ();
 sg13g2_decap_8 FILLER_11_2191 ();
 sg13g2_decap_8 FILLER_11_2198 ();
 sg13g2_decap_8 FILLER_11_2205 ();
 sg13g2_decap_8 FILLER_11_2212 ();
 sg13g2_decap_8 FILLER_11_2219 ();
 sg13g2_decap_8 FILLER_11_2226 ();
 sg13g2_decap_8 FILLER_11_2233 ();
 sg13g2_decap_8 FILLER_11_2240 ();
 sg13g2_decap_8 FILLER_11_2247 ();
 sg13g2_decap_8 FILLER_11_2254 ();
 sg13g2_decap_8 FILLER_11_2261 ();
 sg13g2_decap_8 FILLER_11_2268 ();
 sg13g2_decap_8 FILLER_11_2275 ();
 sg13g2_decap_8 FILLER_11_2282 ();
 sg13g2_decap_8 FILLER_11_2289 ();
 sg13g2_decap_8 FILLER_11_2296 ();
 sg13g2_decap_8 FILLER_11_2303 ();
 sg13g2_decap_8 FILLER_11_2310 ();
 sg13g2_decap_8 FILLER_11_2317 ();
 sg13g2_decap_8 FILLER_11_2324 ();
 sg13g2_decap_8 FILLER_11_2331 ();
 sg13g2_decap_8 FILLER_11_2338 ();
 sg13g2_decap_8 FILLER_11_2345 ();
 sg13g2_decap_8 FILLER_11_2352 ();
 sg13g2_decap_8 FILLER_11_2359 ();
 sg13g2_decap_8 FILLER_11_2366 ();
 sg13g2_decap_8 FILLER_11_2373 ();
 sg13g2_decap_8 FILLER_11_2380 ();
 sg13g2_decap_8 FILLER_11_2387 ();
 sg13g2_decap_8 FILLER_11_2394 ();
 sg13g2_decap_8 FILLER_11_2401 ();
 sg13g2_decap_8 FILLER_11_2408 ();
 sg13g2_decap_8 FILLER_11_2415 ();
 sg13g2_decap_8 FILLER_11_2422 ();
 sg13g2_decap_8 FILLER_11_2429 ();
 sg13g2_decap_8 FILLER_11_2436 ();
 sg13g2_decap_8 FILLER_11_2443 ();
 sg13g2_decap_8 FILLER_11_2450 ();
 sg13g2_decap_8 FILLER_11_2457 ();
 sg13g2_decap_8 FILLER_11_2464 ();
 sg13g2_decap_8 FILLER_11_2471 ();
 sg13g2_decap_8 FILLER_11_2478 ();
 sg13g2_decap_8 FILLER_11_2485 ();
 sg13g2_decap_8 FILLER_11_2492 ();
 sg13g2_decap_8 FILLER_11_2499 ();
 sg13g2_decap_8 FILLER_11_2506 ();
 sg13g2_decap_8 FILLER_11_2513 ();
 sg13g2_decap_8 FILLER_11_2520 ();
 sg13g2_decap_8 FILLER_11_2527 ();
 sg13g2_decap_8 FILLER_11_2534 ();
 sg13g2_decap_8 FILLER_11_2541 ();
 sg13g2_decap_8 FILLER_11_2548 ();
 sg13g2_decap_8 FILLER_11_2555 ();
 sg13g2_decap_8 FILLER_11_2562 ();
 sg13g2_decap_8 FILLER_11_2569 ();
 sg13g2_decap_8 FILLER_11_2576 ();
 sg13g2_decap_8 FILLER_11_2583 ();
 sg13g2_decap_8 FILLER_11_2590 ();
 sg13g2_decap_8 FILLER_11_2597 ();
 sg13g2_decap_8 FILLER_11_2604 ();
 sg13g2_decap_8 FILLER_11_2611 ();
 sg13g2_decap_8 FILLER_11_2618 ();
 sg13g2_decap_8 FILLER_11_2625 ();
 sg13g2_decap_8 FILLER_11_2632 ();
 sg13g2_decap_8 FILLER_11_2639 ();
 sg13g2_decap_8 FILLER_11_2646 ();
 sg13g2_decap_8 FILLER_11_2653 ();
 sg13g2_decap_8 FILLER_11_2660 ();
 sg13g2_decap_8 FILLER_11_2667 ();
 sg13g2_decap_8 FILLER_11_2674 ();
 sg13g2_decap_8 FILLER_11_2681 ();
 sg13g2_decap_8 FILLER_11_2688 ();
 sg13g2_decap_8 FILLER_11_2695 ();
 sg13g2_decap_8 FILLER_11_2702 ();
 sg13g2_decap_8 FILLER_11_2709 ();
 sg13g2_decap_8 FILLER_11_2716 ();
 sg13g2_decap_8 FILLER_11_2723 ();
 sg13g2_decap_8 FILLER_11_2730 ();
 sg13g2_decap_8 FILLER_11_2737 ();
 sg13g2_decap_8 FILLER_11_2744 ();
 sg13g2_decap_8 FILLER_11_2751 ();
 sg13g2_decap_8 FILLER_11_2758 ();
 sg13g2_decap_8 FILLER_11_2765 ();
 sg13g2_decap_8 FILLER_11_2772 ();
 sg13g2_decap_8 FILLER_11_2779 ();
 sg13g2_decap_8 FILLER_11_2786 ();
 sg13g2_decap_8 FILLER_11_2793 ();
 sg13g2_decap_8 FILLER_11_2800 ();
 sg13g2_decap_8 FILLER_11_2807 ();
 sg13g2_decap_8 FILLER_11_2814 ();
 sg13g2_decap_8 FILLER_11_2821 ();
 sg13g2_decap_8 FILLER_11_2828 ();
 sg13g2_decap_8 FILLER_11_2835 ();
 sg13g2_decap_8 FILLER_11_2842 ();
 sg13g2_decap_8 FILLER_11_2849 ();
 sg13g2_decap_8 FILLER_11_2856 ();
 sg13g2_decap_8 FILLER_11_2863 ();
 sg13g2_decap_8 FILLER_11_2870 ();
 sg13g2_decap_8 FILLER_11_2877 ();
 sg13g2_decap_8 FILLER_11_2884 ();
 sg13g2_decap_8 FILLER_11_2891 ();
 sg13g2_decap_8 FILLER_11_2898 ();
 sg13g2_decap_8 FILLER_11_2905 ();
 sg13g2_decap_8 FILLER_11_2912 ();
 sg13g2_decap_8 FILLER_11_2919 ();
 sg13g2_decap_8 FILLER_11_2926 ();
 sg13g2_decap_8 FILLER_11_2933 ();
 sg13g2_decap_8 FILLER_11_2940 ();
 sg13g2_decap_8 FILLER_11_2947 ();
 sg13g2_decap_8 FILLER_11_2954 ();
 sg13g2_decap_8 FILLER_11_2961 ();
 sg13g2_decap_8 FILLER_11_2968 ();
 sg13g2_decap_8 FILLER_11_2975 ();
 sg13g2_decap_8 FILLER_11_2982 ();
 sg13g2_decap_8 FILLER_11_2989 ();
 sg13g2_decap_8 FILLER_11_2996 ();
 sg13g2_decap_8 FILLER_11_3003 ();
 sg13g2_decap_8 FILLER_11_3010 ();
 sg13g2_decap_8 FILLER_11_3017 ();
 sg13g2_decap_8 FILLER_11_3024 ();
 sg13g2_decap_8 FILLER_11_3031 ();
 sg13g2_decap_8 FILLER_11_3038 ();
 sg13g2_decap_8 FILLER_11_3045 ();
 sg13g2_decap_8 FILLER_11_3052 ();
 sg13g2_decap_8 FILLER_11_3059 ();
 sg13g2_decap_8 FILLER_11_3066 ();
 sg13g2_decap_8 FILLER_11_3073 ();
 sg13g2_decap_8 FILLER_11_3080 ();
 sg13g2_decap_8 FILLER_11_3087 ();
 sg13g2_decap_8 FILLER_11_3094 ();
 sg13g2_decap_8 FILLER_11_3101 ();
 sg13g2_decap_8 FILLER_11_3108 ();
 sg13g2_decap_8 FILLER_11_3115 ();
 sg13g2_decap_8 FILLER_11_3122 ();
 sg13g2_decap_8 FILLER_11_3129 ();
 sg13g2_decap_8 FILLER_11_3136 ();
 sg13g2_decap_8 FILLER_11_3143 ();
 sg13g2_decap_8 FILLER_11_3150 ();
 sg13g2_decap_8 FILLER_11_3157 ();
 sg13g2_decap_8 FILLER_11_3164 ();
 sg13g2_decap_8 FILLER_11_3171 ();
 sg13g2_decap_8 FILLER_11_3178 ();
 sg13g2_decap_8 FILLER_11_3185 ();
 sg13g2_decap_8 FILLER_11_3192 ();
 sg13g2_decap_8 FILLER_11_3199 ();
 sg13g2_decap_8 FILLER_11_3206 ();
 sg13g2_decap_8 FILLER_11_3213 ();
 sg13g2_decap_8 FILLER_11_3220 ();
 sg13g2_decap_8 FILLER_11_3227 ();
 sg13g2_decap_8 FILLER_11_3234 ();
 sg13g2_decap_8 FILLER_11_3241 ();
 sg13g2_decap_8 FILLER_11_3248 ();
 sg13g2_decap_8 FILLER_11_3255 ();
 sg13g2_decap_8 FILLER_11_3262 ();
 sg13g2_decap_8 FILLER_11_3269 ();
 sg13g2_decap_8 FILLER_11_3276 ();
 sg13g2_decap_8 FILLER_11_3283 ();
 sg13g2_decap_8 FILLER_11_3290 ();
 sg13g2_decap_8 FILLER_11_3297 ();
 sg13g2_decap_8 FILLER_11_3304 ();
 sg13g2_decap_8 FILLER_11_3311 ();
 sg13g2_decap_8 FILLER_11_3318 ();
 sg13g2_decap_8 FILLER_11_3325 ();
 sg13g2_decap_8 FILLER_11_3332 ();
 sg13g2_decap_8 FILLER_11_3339 ();
 sg13g2_decap_8 FILLER_11_3346 ();
 sg13g2_decap_8 FILLER_11_3353 ();
 sg13g2_decap_8 FILLER_11_3360 ();
 sg13g2_decap_8 FILLER_11_3367 ();
 sg13g2_decap_8 FILLER_11_3374 ();
 sg13g2_decap_8 FILLER_11_3381 ();
 sg13g2_decap_8 FILLER_11_3388 ();
 sg13g2_decap_8 FILLER_11_3395 ();
 sg13g2_decap_8 FILLER_11_3402 ();
 sg13g2_decap_8 FILLER_11_3409 ();
 sg13g2_decap_8 FILLER_11_3416 ();
 sg13g2_decap_8 FILLER_11_3423 ();
 sg13g2_decap_8 FILLER_11_3430 ();
 sg13g2_decap_8 FILLER_11_3437 ();
 sg13g2_decap_8 FILLER_11_3444 ();
 sg13g2_decap_8 FILLER_11_3451 ();
 sg13g2_decap_8 FILLER_11_3458 ();
 sg13g2_decap_8 FILLER_11_3465 ();
 sg13g2_decap_8 FILLER_11_3472 ();
 sg13g2_decap_8 FILLER_11_3479 ();
 sg13g2_decap_8 FILLER_11_3486 ();
 sg13g2_decap_8 FILLER_11_3493 ();
 sg13g2_decap_8 FILLER_11_3500 ();
 sg13g2_decap_8 FILLER_11_3507 ();
 sg13g2_decap_8 FILLER_11_3514 ();
 sg13g2_decap_8 FILLER_11_3521 ();
 sg13g2_decap_8 FILLER_11_3528 ();
 sg13g2_decap_8 FILLER_11_3535 ();
 sg13g2_decap_8 FILLER_11_3542 ();
 sg13g2_decap_8 FILLER_11_3549 ();
 sg13g2_decap_8 FILLER_11_3556 ();
 sg13g2_decap_8 FILLER_11_3563 ();
 sg13g2_decap_8 FILLER_11_3570 ();
 sg13g2_fill_2 FILLER_11_3577 ();
 sg13g2_fill_1 FILLER_11_3579 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_448 ();
 sg13g2_decap_8 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_469 ();
 sg13g2_decap_8 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_518 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_8 FILLER_12_595 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_decap_8 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_12_868 ();
 sg13g2_decap_8 FILLER_12_875 ();
 sg13g2_decap_8 FILLER_12_882 ();
 sg13g2_decap_8 FILLER_12_889 ();
 sg13g2_decap_8 FILLER_12_896 ();
 sg13g2_decap_8 FILLER_12_903 ();
 sg13g2_decap_8 FILLER_12_910 ();
 sg13g2_decap_8 FILLER_12_917 ();
 sg13g2_decap_8 FILLER_12_924 ();
 sg13g2_decap_8 FILLER_12_931 ();
 sg13g2_decap_8 FILLER_12_938 ();
 sg13g2_decap_8 FILLER_12_945 ();
 sg13g2_decap_8 FILLER_12_952 ();
 sg13g2_decap_8 FILLER_12_959 ();
 sg13g2_decap_8 FILLER_12_966 ();
 sg13g2_decap_8 FILLER_12_973 ();
 sg13g2_decap_8 FILLER_12_980 ();
 sg13g2_decap_8 FILLER_12_987 ();
 sg13g2_decap_8 FILLER_12_994 ();
 sg13g2_decap_8 FILLER_12_1001 ();
 sg13g2_decap_8 FILLER_12_1008 ();
 sg13g2_decap_8 FILLER_12_1015 ();
 sg13g2_decap_8 FILLER_12_1022 ();
 sg13g2_decap_8 FILLER_12_1029 ();
 sg13g2_decap_8 FILLER_12_1036 ();
 sg13g2_decap_8 FILLER_12_1043 ();
 sg13g2_decap_8 FILLER_12_1050 ();
 sg13g2_decap_8 FILLER_12_1057 ();
 sg13g2_decap_8 FILLER_12_1064 ();
 sg13g2_decap_8 FILLER_12_1071 ();
 sg13g2_decap_8 FILLER_12_1078 ();
 sg13g2_decap_8 FILLER_12_1085 ();
 sg13g2_decap_8 FILLER_12_1092 ();
 sg13g2_decap_8 FILLER_12_1099 ();
 sg13g2_decap_8 FILLER_12_1106 ();
 sg13g2_decap_8 FILLER_12_1113 ();
 sg13g2_decap_8 FILLER_12_1120 ();
 sg13g2_decap_8 FILLER_12_1127 ();
 sg13g2_decap_8 FILLER_12_1134 ();
 sg13g2_decap_8 FILLER_12_1141 ();
 sg13g2_decap_8 FILLER_12_1148 ();
 sg13g2_decap_8 FILLER_12_1155 ();
 sg13g2_decap_8 FILLER_12_1162 ();
 sg13g2_decap_8 FILLER_12_1169 ();
 sg13g2_decap_8 FILLER_12_1176 ();
 sg13g2_decap_8 FILLER_12_1183 ();
 sg13g2_decap_8 FILLER_12_1190 ();
 sg13g2_decap_8 FILLER_12_1197 ();
 sg13g2_decap_8 FILLER_12_1204 ();
 sg13g2_decap_8 FILLER_12_1211 ();
 sg13g2_decap_8 FILLER_12_1218 ();
 sg13g2_decap_8 FILLER_12_1225 ();
 sg13g2_decap_8 FILLER_12_1232 ();
 sg13g2_decap_8 FILLER_12_1239 ();
 sg13g2_decap_8 FILLER_12_1246 ();
 sg13g2_decap_8 FILLER_12_1253 ();
 sg13g2_decap_8 FILLER_12_1260 ();
 sg13g2_decap_8 FILLER_12_1267 ();
 sg13g2_decap_8 FILLER_12_1274 ();
 sg13g2_decap_8 FILLER_12_1281 ();
 sg13g2_decap_8 FILLER_12_1288 ();
 sg13g2_decap_8 FILLER_12_1295 ();
 sg13g2_decap_8 FILLER_12_1302 ();
 sg13g2_decap_8 FILLER_12_1309 ();
 sg13g2_decap_8 FILLER_12_1316 ();
 sg13g2_decap_8 FILLER_12_1323 ();
 sg13g2_decap_8 FILLER_12_1330 ();
 sg13g2_decap_8 FILLER_12_1337 ();
 sg13g2_decap_8 FILLER_12_1344 ();
 sg13g2_decap_8 FILLER_12_1351 ();
 sg13g2_decap_8 FILLER_12_1358 ();
 sg13g2_decap_8 FILLER_12_1365 ();
 sg13g2_decap_8 FILLER_12_1372 ();
 sg13g2_decap_8 FILLER_12_1379 ();
 sg13g2_decap_8 FILLER_12_1386 ();
 sg13g2_decap_8 FILLER_12_1393 ();
 sg13g2_decap_8 FILLER_12_1400 ();
 sg13g2_decap_8 FILLER_12_1407 ();
 sg13g2_decap_8 FILLER_12_1414 ();
 sg13g2_decap_8 FILLER_12_1421 ();
 sg13g2_decap_8 FILLER_12_1428 ();
 sg13g2_decap_8 FILLER_12_1435 ();
 sg13g2_decap_8 FILLER_12_1442 ();
 sg13g2_decap_8 FILLER_12_1449 ();
 sg13g2_decap_8 FILLER_12_1456 ();
 sg13g2_decap_8 FILLER_12_1463 ();
 sg13g2_decap_8 FILLER_12_1470 ();
 sg13g2_decap_8 FILLER_12_1477 ();
 sg13g2_decap_8 FILLER_12_1484 ();
 sg13g2_decap_8 FILLER_12_1491 ();
 sg13g2_decap_8 FILLER_12_1498 ();
 sg13g2_decap_8 FILLER_12_1505 ();
 sg13g2_decap_8 FILLER_12_1512 ();
 sg13g2_decap_8 FILLER_12_1519 ();
 sg13g2_decap_8 FILLER_12_1526 ();
 sg13g2_decap_8 FILLER_12_1533 ();
 sg13g2_decap_8 FILLER_12_1540 ();
 sg13g2_decap_8 FILLER_12_1547 ();
 sg13g2_decap_8 FILLER_12_1554 ();
 sg13g2_decap_8 FILLER_12_1561 ();
 sg13g2_decap_8 FILLER_12_1568 ();
 sg13g2_decap_8 FILLER_12_1575 ();
 sg13g2_decap_8 FILLER_12_1582 ();
 sg13g2_decap_8 FILLER_12_1589 ();
 sg13g2_decap_8 FILLER_12_1596 ();
 sg13g2_decap_8 FILLER_12_1603 ();
 sg13g2_decap_8 FILLER_12_1610 ();
 sg13g2_decap_8 FILLER_12_1617 ();
 sg13g2_decap_8 FILLER_12_1624 ();
 sg13g2_decap_8 FILLER_12_1631 ();
 sg13g2_decap_8 FILLER_12_1638 ();
 sg13g2_decap_8 FILLER_12_1645 ();
 sg13g2_decap_8 FILLER_12_1652 ();
 sg13g2_decap_8 FILLER_12_1659 ();
 sg13g2_decap_8 FILLER_12_1666 ();
 sg13g2_decap_8 FILLER_12_1673 ();
 sg13g2_decap_8 FILLER_12_1680 ();
 sg13g2_decap_8 FILLER_12_1687 ();
 sg13g2_decap_8 FILLER_12_1694 ();
 sg13g2_decap_8 FILLER_12_1701 ();
 sg13g2_decap_8 FILLER_12_1708 ();
 sg13g2_decap_8 FILLER_12_1715 ();
 sg13g2_decap_8 FILLER_12_1722 ();
 sg13g2_decap_8 FILLER_12_1729 ();
 sg13g2_decap_8 FILLER_12_1736 ();
 sg13g2_decap_8 FILLER_12_1743 ();
 sg13g2_decap_8 FILLER_12_1750 ();
 sg13g2_decap_8 FILLER_12_1757 ();
 sg13g2_decap_8 FILLER_12_1764 ();
 sg13g2_decap_8 FILLER_12_1771 ();
 sg13g2_decap_8 FILLER_12_1778 ();
 sg13g2_decap_8 FILLER_12_1785 ();
 sg13g2_decap_8 FILLER_12_1792 ();
 sg13g2_decap_8 FILLER_12_1799 ();
 sg13g2_decap_8 FILLER_12_1806 ();
 sg13g2_decap_8 FILLER_12_1813 ();
 sg13g2_decap_8 FILLER_12_1820 ();
 sg13g2_decap_8 FILLER_12_1827 ();
 sg13g2_decap_8 FILLER_12_1834 ();
 sg13g2_decap_8 FILLER_12_1841 ();
 sg13g2_decap_8 FILLER_12_1848 ();
 sg13g2_decap_8 FILLER_12_1855 ();
 sg13g2_decap_8 FILLER_12_1862 ();
 sg13g2_decap_8 FILLER_12_1869 ();
 sg13g2_decap_8 FILLER_12_1876 ();
 sg13g2_decap_8 FILLER_12_1883 ();
 sg13g2_decap_8 FILLER_12_1890 ();
 sg13g2_decap_8 FILLER_12_1897 ();
 sg13g2_decap_8 FILLER_12_1904 ();
 sg13g2_decap_8 FILLER_12_1911 ();
 sg13g2_decap_8 FILLER_12_1918 ();
 sg13g2_decap_8 FILLER_12_1925 ();
 sg13g2_decap_8 FILLER_12_1932 ();
 sg13g2_decap_8 FILLER_12_1939 ();
 sg13g2_decap_8 FILLER_12_1946 ();
 sg13g2_decap_8 FILLER_12_1953 ();
 sg13g2_decap_8 FILLER_12_1960 ();
 sg13g2_decap_8 FILLER_12_1967 ();
 sg13g2_decap_8 FILLER_12_1974 ();
 sg13g2_decap_8 FILLER_12_1981 ();
 sg13g2_decap_8 FILLER_12_1988 ();
 sg13g2_decap_8 FILLER_12_1995 ();
 sg13g2_decap_8 FILLER_12_2002 ();
 sg13g2_decap_8 FILLER_12_2009 ();
 sg13g2_decap_8 FILLER_12_2016 ();
 sg13g2_decap_8 FILLER_12_2023 ();
 sg13g2_decap_8 FILLER_12_2030 ();
 sg13g2_decap_8 FILLER_12_2037 ();
 sg13g2_decap_8 FILLER_12_2044 ();
 sg13g2_decap_8 FILLER_12_2051 ();
 sg13g2_decap_8 FILLER_12_2058 ();
 sg13g2_decap_8 FILLER_12_2065 ();
 sg13g2_decap_8 FILLER_12_2072 ();
 sg13g2_decap_8 FILLER_12_2079 ();
 sg13g2_decap_8 FILLER_12_2086 ();
 sg13g2_decap_8 FILLER_12_2093 ();
 sg13g2_decap_8 FILLER_12_2100 ();
 sg13g2_decap_8 FILLER_12_2107 ();
 sg13g2_decap_8 FILLER_12_2114 ();
 sg13g2_decap_8 FILLER_12_2121 ();
 sg13g2_decap_8 FILLER_12_2128 ();
 sg13g2_decap_8 FILLER_12_2135 ();
 sg13g2_decap_8 FILLER_12_2142 ();
 sg13g2_decap_8 FILLER_12_2149 ();
 sg13g2_decap_8 FILLER_12_2156 ();
 sg13g2_decap_8 FILLER_12_2163 ();
 sg13g2_decap_8 FILLER_12_2170 ();
 sg13g2_decap_8 FILLER_12_2177 ();
 sg13g2_decap_8 FILLER_12_2184 ();
 sg13g2_decap_8 FILLER_12_2191 ();
 sg13g2_decap_8 FILLER_12_2198 ();
 sg13g2_decap_8 FILLER_12_2205 ();
 sg13g2_decap_8 FILLER_12_2212 ();
 sg13g2_decap_8 FILLER_12_2219 ();
 sg13g2_decap_8 FILLER_12_2226 ();
 sg13g2_decap_8 FILLER_12_2233 ();
 sg13g2_decap_8 FILLER_12_2240 ();
 sg13g2_decap_8 FILLER_12_2247 ();
 sg13g2_decap_8 FILLER_12_2254 ();
 sg13g2_decap_8 FILLER_12_2261 ();
 sg13g2_decap_8 FILLER_12_2268 ();
 sg13g2_decap_8 FILLER_12_2275 ();
 sg13g2_decap_8 FILLER_12_2282 ();
 sg13g2_decap_8 FILLER_12_2289 ();
 sg13g2_decap_8 FILLER_12_2296 ();
 sg13g2_decap_8 FILLER_12_2303 ();
 sg13g2_decap_8 FILLER_12_2310 ();
 sg13g2_decap_8 FILLER_12_2317 ();
 sg13g2_decap_8 FILLER_12_2324 ();
 sg13g2_decap_8 FILLER_12_2331 ();
 sg13g2_decap_8 FILLER_12_2338 ();
 sg13g2_decap_8 FILLER_12_2345 ();
 sg13g2_decap_8 FILLER_12_2352 ();
 sg13g2_decap_8 FILLER_12_2359 ();
 sg13g2_decap_8 FILLER_12_2366 ();
 sg13g2_decap_8 FILLER_12_2373 ();
 sg13g2_decap_8 FILLER_12_2380 ();
 sg13g2_decap_8 FILLER_12_2387 ();
 sg13g2_decap_8 FILLER_12_2394 ();
 sg13g2_decap_8 FILLER_12_2401 ();
 sg13g2_decap_8 FILLER_12_2408 ();
 sg13g2_decap_8 FILLER_12_2415 ();
 sg13g2_decap_8 FILLER_12_2422 ();
 sg13g2_decap_8 FILLER_12_2429 ();
 sg13g2_decap_8 FILLER_12_2436 ();
 sg13g2_decap_8 FILLER_12_2443 ();
 sg13g2_decap_8 FILLER_12_2450 ();
 sg13g2_decap_8 FILLER_12_2457 ();
 sg13g2_decap_8 FILLER_12_2464 ();
 sg13g2_decap_8 FILLER_12_2471 ();
 sg13g2_decap_8 FILLER_12_2478 ();
 sg13g2_decap_8 FILLER_12_2485 ();
 sg13g2_decap_8 FILLER_12_2492 ();
 sg13g2_decap_8 FILLER_12_2499 ();
 sg13g2_decap_8 FILLER_12_2506 ();
 sg13g2_decap_8 FILLER_12_2513 ();
 sg13g2_decap_8 FILLER_12_2520 ();
 sg13g2_decap_8 FILLER_12_2527 ();
 sg13g2_decap_8 FILLER_12_2534 ();
 sg13g2_decap_8 FILLER_12_2541 ();
 sg13g2_decap_8 FILLER_12_2548 ();
 sg13g2_decap_8 FILLER_12_2555 ();
 sg13g2_decap_8 FILLER_12_2562 ();
 sg13g2_decap_8 FILLER_12_2569 ();
 sg13g2_decap_8 FILLER_12_2576 ();
 sg13g2_decap_8 FILLER_12_2583 ();
 sg13g2_decap_8 FILLER_12_2590 ();
 sg13g2_decap_8 FILLER_12_2597 ();
 sg13g2_decap_8 FILLER_12_2604 ();
 sg13g2_decap_8 FILLER_12_2611 ();
 sg13g2_decap_8 FILLER_12_2618 ();
 sg13g2_decap_8 FILLER_12_2625 ();
 sg13g2_decap_8 FILLER_12_2632 ();
 sg13g2_decap_8 FILLER_12_2639 ();
 sg13g2_decap_8 FILLER_12_2646 ();
 sg13g2_decap_8 FILLER_12_2653 ();
 sg13g2_decap_8 FILLER_12_2660 ();
 sg13g2_decap_8 FILLER_12_2667 ();
 sg13g2_decap_8 FILLER_12_2674 ();
 sg13g2_decap_8 FILLER_12_2681 ();
 sg13g2_decap_8 FILLER_12_2688 ();
 sg13g2_decap_8 FILLER_12_2695 ();
 sg13g2_decap_8 FILLER_12_2702 ();
 sg13g2_decap_8 FILLER_12_2709 ();
 sg13g2_decap_8 FILLER_12_2716 ();
 sg13g2_decap_8 FILLER_12_2723 ();
 sg13g2_decap_8 FILLER_12_2730 ();
 sg13g2_decap_8 FILLER_12_2737 ();
 sg13g2_decap_8 FILLER_12_2744 ();
 sg13g2_decap_8 FILLER_12_2751 ();
 sg13g2_decap_8 FILLER_12_2758 ();
 sg13g2_decap_8 FILLER_12_2765 ();
 sg13g2_decap_8 FILLER_12_2772 ();
 sg13g2_decap_8 FILLER_12_2779 ();
 sg13g2_decap_8 FILLER_12_2786 ();
 sg13g2_decap_8 FILLER_12_2793 ();
 sg13g2_decap_8 FILLER_12_2800 ();
 sg13g2_decap_8 FILLER_12_2807 ();
 sg13g2_decap_8 FILLER_12_2814 ();
 sg13g2_decap_8 FILLER_12_2821 ();
 sg13g2_decap_8 FILLER_12_2828 ();
 sg13g2_decap_8 FILLER_12_2835 ();
 sg13g2_decap_8 FILLER_12_2842 ();
 sg13g2_decap_8 FILLER_12_2849 ();
 sg13g2_decap_8 FILLER_12_2856 ();
 sg13g2_decap_8 FILLER_12_2863 ();
 sg13g2_decap_8 FILLER_12_2870 ();
 sg13g2_decap_8 FILLER_12_2877 ();
 sg13g2_decap_8 FILLER_12_2884 ();
 sg13g2_decap_8 FILLER_12_2891 ();
 sg13g2_decap_8 FILLER_12_2898 ();
 sg13g2_decap_8 FILLER_12_2905 ();
 sg13g2_decap_8 FILLER_12_2912 ();
 sg13g2_decap_8 FILLER_12_2919 ();
 sg13g2_decap_8 FILLER_12_2926 ();
 sg13g2_decap_8 FILLER_12_2933 ();
 sg13g2_decap_8 FILLER_12_2940 ();
 sg13g2_decap_8 FILLER_12_2947 ();
 sg13g2_decap_8 FILLER_12_2954 ();
 sg13g2_decap_8 FILLER_12_2961 ();
 sg13g2_decap_8 FILLER_12_2968 ();
 sg13g2_decap_8 FILLER_12_2975 ();
 sg13g2_decap_8 FILLER_12_2982 ();
 sg13g2_decap_8 FILLER_12_2989 ();
 sg13g2_decap_8 FILLER_12_2996 ();
 sg13g2_decap_8 FILLER_12_3003 ();
 sg13g2_decap_8 FILLER_12_3010 ();
 sg13g2_decap_8 FILLER_12_3017 ();
 sg13g2_decap_8 FILLER_12_3024 ();
 sg13g2_decap_8 FILLER_12_3031 ();
 sg13g2_decap_8 FILLER_12_3038 ();
 sg13g2_decap_8 FILLER_12_3045 ();
 sg13g2_decap_8 FILLER_12_3052 ();
 sg13g2_decap_8 FILLER_12_3059 ();
 sg13g2_decap_8 FILLER_12_3066 ();
 sg13g2_decap_8 FILLER_12_3073 ();
 sg13g2_decap_8 FILLER_12_3080 ();
 sg13g2_decap_8 FILLER_12_3087 ();
 sg13g2_decap_8 FILLER_12_3094 ();
 sg13g2_decap_8 FILLER_12_3101 ();
 sg13g2_decap_8 FILLER_12_3108 ();
 sg13g2_decap_8 FILLER_12_3115 ();
 sg13g2_decap_8 FILLER_12_3122 ();
 sg13g2_decap_8 FILLER_12_3129 ();
 sg13g2_decap_8 FILLER_12_3136 ();
 sg13g2_decap_8 FILLER_12_3143 ();
 sg13g2_decap_8 FILLER_12_3150 ();
 sg13g2_decap_8 FILLER_12_3157 ();
 sg13g2_decap_8 FILLER_12_3164 ();
 sg13g2_decap_8 FILLER_12_3171 ();
 sg13g2_decap_8 FILLER_12_3178 ();
 sg13g2_decap_8 FILLER_12_3185 ();
 sg13g2_decap_8 FILLER_12_3192 ();
 sg13g2_decap_8 FILLER_12_3199 ();
 sg13g2_decap_8 FILLER_12_3206 ();
 sg13g2_decap_8 FILLER_12_3213 ();
 sg13g2_decap_8 FILLER_12_3220 ();
 sg13g2_decap_8 FILLER_12_3227 ();
 sg13g2_decap_8 FILLER_12_3234 ();
 sg13g2_decap_8 FILLER_12_3241 ();
 sg13g2_decap_8 FILLER_12_3248 ();
 sg13g2_decap_8 FILLER_12_3255 ();
 sg13g2_decap_8 FILLER_12_3262 ();
 sg13g2_decap_8 FILLER_12_3269 ();
 sg13g2_decap_8 FILLER_12_3276 ();
 sg13g2_decap_8 FILLER_12_3283 ();
 sg13g2_decap_8 FILLER_12_3290 ();
 sg13g2_decap_8 FILLER_12_3297 ();
 sg13g2_decap_8 FILLER_12_3304 ();
 sg13g2_decap_8 FILLER_12_3311 ();
 sg13g2_decap_8 FILLER_12_3318 ();
 sg13g2_decap_8 FILLER_12_3325 ();
 sg13g2_decap_8 FILLER_12_3332 ();
 sg13g2_decap_8 FILLER_12_3339 ();
 sg13g2_decap_8 FILLER_12_3346 ();
 sg13g2_decap_8 FILLER_12_3353 ();
 sg13g2_decap_8 FILLER_12_3360 ();
 sg13g2_decap_8 FILLER_12_3367 ();
 sg13g2_decap_8 FILLER_12_3374 ();
 sg13g2_decap_8 FILLER_12_3381 ();
 sg13g2_decap_8 FILLER_12_3388 ();
 sg13g2_decap_8 FILLER_12_3395 ();
 sg13g2_decap_8 FILLER_12_3402 ();
 sg13g2_decap_8 FILLER_12_3409 ();
 sg13g2_decap_8 FILLER_12_3416 ();
 sg13g2_decap_8 FILLER_12_3423 ();
 sg13g2_decap_8 FILLER_12_3430 ();
 sg13g2_decap_8 FILLER_12_3437 ();
 sg13g2_decap_8 FILLER_12_3444 ();
 sg13g2_decap_8 FILLER_12_3451 ();
 sg13g2_decap_8 FILLER_12_3458 ();
 sg13g2_decap_8 FILLER_12_3465 ();
 sg13g2_decap_8 FILLER_12_3472 ();
 sg13g2_decap_8 FILLER_12_3479 ();
 sg13g2_decap_8 FILLER_12_3486 ();
 sg13g2_decap_8 FILLER_12_3493 ();
 sg13g2_decap_8 FILLER_12_3500 ();
 sg13g2_decap_8 FILLER_12_3507 ();
 sg13g2_decap_8 FILLER_12_3514 ();
 sg13g2_decap_8 FILLER_12_3521 ();
 sg13g2_decap_8 FILLER_12_3528 ();
 sg13g2_decap_8 FILLER_12_3535 ();
 sg13g2_decap_8 FILLER_12_3542 ();
 sg13g2_decap_8 FILLER_12_3549 ();
 sg13g2_decap_8 FILLER_12_3556 ();
 sg13g2_decap_8 FILLER_12_3563 ();
 sg13g2_decap_8 FILLER_12_3570 ();
 sg13g2_fill_2 FILLER_12_3577 ();
 sg13g2_fill_1 FILLER_12_3579 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_8 FILLER_13_462 ();
 sg13g2_decap_8 FILLER_13_469 ();
 sg13g2_decap_8 FILLER_13_476 ();
 sg13g2_decap_8 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_490 ();
 sg13g2_decap_8 FILLER_13_497 ();
 sg13g2_decap_8 FILLER_13_504 ();
 sg13g2_decap_8 FILLER_13_511 ();
 sg13g2_decap_8 FILLER_13_518 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_decap_8 FILLER_13_532 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_decap_8 FILLER_13_546 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_560 ();
 sg13g2_decap_8 FILLER_13_567 ();
 sg13g2_decap_8 FILLER_13_574 ();
 sg13g2_decap_8 FILLER_13_581 ();
 sg13g2_decap_8 FILLER_13_588 ();
 sg13g2_decap_8 FILLER_13_595 ();
 sg13g2_decap_8 FILLER_13_602 ();
 sg13g2_decap_8 FILLER_13_609 ();
 sg13g2_decap_8 FILLER_13_616 ();
 sg13g2_decap_8 FILLER_13_623 ();
 sg13g2_decap_8 FILLER_13_630 ();
 sg13g2_decap_8 FILLER_13_637 ();
 sg13g2_decap_8 FILLER_13_644 ();
 sg13g2_decap_8 FILLER_13_651 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_679 ();
 sg13g2_decap_8 FILLER_13_686 ();
 sg13g2_decap_8 FILLER_13_693 ();
 sg13g2_decap_8 FILLER_13_700 ();
 sg13g2_decap_8 FILLER_13_707 ();
 sg13g2_decap_8 FILLER_13_714 ();
 sg13g2_decap_8 FILLER_13_721 ();
 sg13g2_decap_8 FILLER_13_728 ();
 sg13g2_decap_8 FILLER_13_735 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_763 ();
 sg13g2_decap_8 FILLER_13_770 ();
 sg13g2_decap_8 FILLER_13_777 ();
 sg13g2_decap_8 FILLER_13_784 ();
 sg13g2_decap_8 FILLER_13_791 ();
 sg13g2_decap_8 FILLER_13_798 ();
 sg13g2_decap_8 FILLER_13_805 ();
 sg13g2_decap_8 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_819 ();
 sg13g2_decap_8 FILLER_13_826 ();
 sg13g2_decap_8 FILLER_13_833 ();
 sg13g2_decap_8 FILLER_13_840 ();
 sg13g2_decap_8 FILLER_13_847 ();
 sg13g2_decap_8 FILLER_13_854 ();
 sg13g2_decap_8 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_13_868 ();
 sg13g2_decap_8 FILLER_13_875 ();
 sg13g2_decap_8 FILLER_13_882 ();
 sg13g2_decap_8 FILLER_13_889 ();
 sg13g2_decap_8 FILLER_13_896 ();
 sg13g2_decap_8 FILLER_13_903 ();
 sg13g2_decap_8 FILLER_13_910 ();
 sg13g2_decap_8 FILLER_13_917 ();
 sg13g2_decap_8 FILLER_13_924 ();
 sg13g2_decap_8 FILLER_13_931 ();
 sg13g2_decap_8 FILLER_13_938 ();
 sg13g2_decap_8 FILLER_13_945 ();
 sg13g2_decap_8 FILLER_13_952 ();
 sg13g2_decap_8 FILLER_13_959 ();
 sg13g2_decap_8 FILLER_13_966 ();
 sg13g2_decap_8 FILLER_13_973 ();
 sg13g2_decap_8 FILLER_13_980 ();
 sg13g2_decap_8 FILLER_13_987 ();
 sg13g2_decap_8 FILLER_13_994 ();
 sg13g2_decap_8 FILLER_13_1001 ();
 sg13g2_decap_8 FILLER_13_1008 ();
 sg13g2_decap_8 FILLER_13_1015 ();
 sg13g2_decap_8 FILLER_13_1022 ();
 sg13g2_decap_8 FILLER_13_1029 ();
 sg13g2_decap_8 FILLER_13_1036 ();
 sg13g2_decap_8 FILLER_13_1043 ();
 sg13g2_decap_8 FILLER_13_1050 ();
 sg13g2_decap_8 FILLER_13_1057 ();
 sg13g2_decap_8 FILLER_13_1064 ();
 sg13g2_decap_8 FILLER_13_1071 ();
 sg13g2_decap_8 FILLER_13_1078 ();
 sg13g2_decap_8 FILLER_13_1085 ();
 sg13g2_decap_8 FILLER_13_1092 ();
 sg13g2_decap_8 FILLER_13_1099 ();
 sg13g2_decap_8 FILLER_13_1106 ();
 sg13g2_decap_8 FILLER_13_1113 ();
 sg13g2_decap_8 FILLER_13_1120 ();
 sg13g2_decap_8 FILLER_13_1127 ();
 sg13g2_decap_8 FILLER_13_1134 ();
 sg13g2_decap_8 FILLER_13_1141 ();
 sg13g2_decap_8 FILLER_13_1148 ();
 sg13g2_decap_8 FILLER_13_1155 ();
 sg13g2_decap_8 FILLER_13_1162 ();
 sg13g2_decap_8 FILLER_13_1169 ();
 sg13g2_decap_8 FILLER_13_1176 ();
 sg13g2_decap_8 FILLER_13_1183 ();
 sg13g2_decap_8 FILLER_13_1190 ();
 sg13g2_decap_8 FILLER_13_1197 ();
 sg13g2_decap_8 FILLER_13_1204 ();
 sg13g2_decap_8 FILLER_13_1211 ();
 sg13g2_decap_8 FILLER_13_1218 ();
 sg13g2_decap_8 FILLER_13_1225 ();
 sg13g2_decap_8 FILLER_13_1232 ();
 sg13g2_decap_8 FILLER_13_1239 ();
 sg13g2_decap_8 FILLER_13_1246 ();
 sg13g2_decap_8 FILLER_13_1253 ();
 sg13g2_decap_8 FILLER_13_1260 ();
 sg13g2_decap_8 FILLER_13_1267 ();
 sg13g2_decap_8 FILLER_13_1274 ();
 sg13g2_decap_8 FILLER_13_1281 ();
 sg13g2_decap_8 FILLER_13_1288 ();
 sg13g2_decap_8 FILLER_13_1295 ();
 sg13g2_decap_8 FILLER_13_1302 ();
 sg13g2_decap_8 FILLER_13_1309 ();
 sg13g2_decap_8 FILLER_13_1316 ();
 sg13g2_decap_8 FILLER_13_1323 ();
 sg13g2_decap_8 FILLER_13_1330 ();
 sg13g2_decap_8 FILLER_13_1337 ();
 sg13g2_decap_8 FILLER_13_1344 ();
 sg13g2_decap_8 FILLER_13_1351 ();
 sg13g2_decap_8 FILLER_13_1358 ();
 sg13g2_decap_8 FILLER_13_1365 ();
 sg13g2_decap_8 FILLER_13_1372 ();
 sg13g2_decap_8 FILLER_13_1379 ();
 sg13g2_decap_8 FILLER_13_1386 ();
 sg13g2_decap_8 FILLER_13_1393 ();
 sg13g2_decap_8 FILLER_13_1400 ();
 sg13g2_decap_8 FILLER_13_1407 ();
 sg13g2_decap_8 FILLER_13_1414 ();
 sg13g2_decap_8 FILLER_13_1421 ();
 sg13g2_decap_8 FILLER_13_1428 ();
 sg13g2_decap_8 FILLER_13_1435 ();
 sg13g2_decap_8 FILLER_13_1442 ();
 sg13g2_decap_8 FILLER_13_1449 ();
 sg13g2_decap_8 FILLER_13_1456 ();
 sg13g2_decap_8 FILLER_13_1463 ();
 sg13g2_decap_8 FILLER_13_1470 ();
 sg13g2_decap_8 FILLER_13_1477 ();
 sg13g2_decap_8 FILLER_13_1484 ();
 sg13g2_decap_8 FILLER_13_1491 ();
 sg13g2_decap_8 FILLER_13_1498 ();
 sg13g2_decap_8 FILLER_13_1505 ();
 sg13g2_decap_8 FILLER_13_1512 ();
 sg13g2_decap_8 FILLER_13_1519 ();
 sg13g2_decap_8 FILLER_13_1526 ();
 sg13g2_decap_8 FILLER_13_1533 ();
 sg13g2_decap_8 FILLER_13_1540 ();
 sg13g2_decap_8 FILLER_13_1547 ();
 sg13g2_decap_8 FILLER_13_1554 ();
 sg13g2_decap_8 FILLER_13_1561 ();
 sg13g2_decap_8 FILLER_13_1568 ();
 sg13g2_decap_8 FILLER_13_1575 ();
 sg13g2_decap_8 FILLER_13_1582 ();
 sg13g2_decap_8 FILLER_13_1589 ();
 sg13g2_decap_8 FILLER_13_1596 ();
 sg13g2_decap_8 FILLER_13_1603 ();
 sg13g2_decap_8 FILLER_13_1610 ();
 sg13g2_decap_8 FILLER_13_1617 ();
 sg13g2_decap_8 FILLER_13_1624 ();
 sg13g2_decap_8 FILLER_13_1631 ();
 sg13g2_decap_8 FILLER_13_1638 ();
 sg13g2_decap_8 FILLER_13_1645 ();
 sg13g2_decap_8 FILLER_13_1652 ();
 sg13g2_decap_8 FILLER_13_1659 ();
 sg13g2_decap_8 FILLER_13_1666 ();
 sg13g2_decap_8 FILLER_13_1673 ();
 sg13g2_decap_8 FILLER_13_1680 ();
 sg13g2_decap_8 FILLER_13_1687 ();
 sg13g2_decap_8 FILLER_13_1694 ();
 sg13g2_decap_8 FILLER_13_1701 ();
 sg13g2_decap_8 FILLER_13_1708 ();
 sg13g2_decap_8 FILLER_13_1715 ();
 sg13g2_decap_8 FILLER_13_1722 ();
 sg13g2_decap_8 FILLER_13_1729 ();
 sg13g2_decap_8 FILLER_13_1736 ();
 sg13g2_decap_8 FILLER_13_1743 ();
 sg13g2_decap_8 FILLER_13_1750 ();
 sg13g2_decap_8 FILLER_13_1757 ();
 sg13g2_decap_8 FILLER_13_1764 ();
 sg13g2_decap_8 FILLER_13_1771 ();
 sg13g2_decap_8 FILLER_13_1778 ();
 sg13g2_decap_8 FILLER_13_1785 ();
 sg13g2_decap_8 FILLER_13_1792 ();
 sg13g2_decap_8 FILLER_13_1799 ();
 sg13g2_decap_8 FILLER_13_1806 ();
 sg13g2_decap_8 FILLER_13_1813 ();
 sg13g2_decap_8 FILLER_13_1820 ();
 sg13g2_decap_8 FILLER_13_1827 ();
 sg13g2_decap_8 FILLER_13_1834 ();
 sg13g2_decap_8 FILLER_13_1841 ();
 sg13g2_decap_8 FILLER_13_1848 ();
 sg13g2_decap_8 FILLER_13_1855 ();
 sg13g2_decap_8 FILLER_13_1862 ();
 sg13g2_decap_8 FILLER_13_1869 ();
 sg13g2_decap_8 FILLER_13_1876 ();
 sg13g2_decap_8 FILLER_13_1883 ();
 sg13g2_decap_8 FILLER_13_1890 ();
 sg13g2_decap_8 FILLER_13_1897 ();
 sg13g2_decap_8 FILLER_13_1904 ();
 sg13g2_decap_8 FILLER_13_1911 ();
 sg13g2_decap_8 FILLER_13_1918 ();
 sg13g2_decap_8 FILLER_13_1925 ();
 sg13g2_decap_8 FILLER_13_1932 ();
 sg13g2_decap_8 FILLER_13_1939 ();
 sg13g2_decap_8 FILLER_13_1946 ();
 sg13g2_decap_8 FILLER_13_1953 ();
 sg13g2_decap_8 FILLER_13_1960 ();
 sg13g2_decap_8 FILLER_13_1967 ();
 sg13g2_decap_8 FILLER_13_1974 ();
 sg13g2_decap_8 FILLER_13_1981 ();
 sg13g2_decap_8 FILLER_13_1988 ();
 sg13g2_decap_8 FILLER_13_1995 ();
 sg13g2_decap_8 FILLER_13_2002 ();
 sg13g2_decap_8 FILLER_13_2009 ();
 sg13g2_decap_8 FILLER_13_2016 ();
 sg13g2_decap_8 FILLER_13_2023 ();
 sg13g2_decap_8 FILLER_13_2030 ();
 sg13g2_decap_8 FILLER_13_2037 ();
 sg13g2_decap_8 FILLER_13_2044 ();
 sg13g2_decap_8 FILLER_13_2051 ();
 sg13g2_decap_8 FILLER_13_2058 ();
 sg13g2_decap_8 FILLER_13_2065 ();
 sg13g2_decap_8 FILLER_13_2072 ();
 sg13g2_decap_8 FILLER_13_2079 ();
 sg13g2_decap_8 FILLER_13_2086 ();
 sg13g2_decap_8 FILLER_13_2093 ();
 sg13g2_decap_8 FILLER_13_2100 ();
 sg13g2_decap_8 FILLER_13_2107 ();
 sg13g2_decap_8 FILLER_13_2114 ();
 sg13g2_decap_8 FILLER_13_2121 ();
 sg13g2_decap_8 FILLER_13_2128 ();
 sg13g2_decap_8 FILLER_13_2135 ();
 sg13g2_decap_8 FILLER_13_2142 ();
 sg13g2_decap_8 FILLER_13_2149 ();
 sg13g2_decap_8 FILLER_13_2156 ();
 sg13g2_decap_8 FILLER_13_2163 ();
 sg13g2_decap_8 FILLER_13_2170 ();
 sg13g2_decap_8 FILLER_13_2177 ();
 sg13g2_decap_8 FILLER_13_2184 ();
 sg13g2_decap_8 FILLER_13_2191 ();
 sg13g2_decap_8 FILLER_13_2198 ();
 sg13g2_decap_8 FILLER_13_2205 ();
 sg13g2_decap_8 FILLER_13_2212 ();
 sg13g2_decap_8 FILLER_13_2219 ();
 sg13g2_decap_8 FILLER_13_2226 ();
 sg13g2_decap_8 FILLER_13_2233 ();
 sg13g2_decap_8 FILLER_13_2240 ();
 sg13g2_decap_8 FILLER_13_2247 ();
 sg13g2_decap_8 FILLER_13_2254 ();
 sg13g2_decap_8 FILLER_13_2261 ();
 sg13g2_decap_8 FILLER_13_2268 ();
 sg13g2_decap_8 FILLER_13_2275 ();
 sg13g2_decap_8 FILLER_13_2282 ();
 sg13g2_decap_8 FILLER_13_2289 ();
 sg13g2_decap_8 FILLER_13_2296 ();
 sg13g2_decap_8 FILLER_13_2303 ();
 sg13g2_decap_8 FILLER_13_2310 ();
 sg13g2_decap_8 FILLER_13_2317 ();
 sg13g2_decap_8 FILLER_13_2324 ();
 sg13g2_decap_8 FILLER_13_2331 ();
 sg13g2_decap_8 FILLER_13_2338 ();
 sg13g2_decap_8 FILLER_13_2345 ();
 sg13g2_decap_8 FILLER_13_2352 ();
 sg13g2_decap_8 FILLER_13_2359 ();
 sg13g2_decap_8 FILLER_13_2366 ();
 sg13g2_decap_8 FILLER_13_2373 ();
 sg13g2_decap_8 FILLER_13_2380 ();
 sg13g2_decap_8 FILLER_13_2387 ();
 sg13g2_decap_8 FILLER_13_2394 ();
 sg13g2_decap_8 FILLER_13_2401 ();
 sg13g2_decap_8 FILLER_13_2408 ();
 sg13g2_decap_8 FILLER_13_2415 ();
 sg13g2_decap_8 FILLER_13_2422 ();
 sg13g2_decap_8 FILLER_13_2429 ();
 sg13g2_decap_8 FILLER_13_2436 ();
 sg13g2_decap_8 FILLER_13_2443 ();
 sg13g2_decap_8 FILLER_13_2450 ();
 sg13g2_decap_8 FILLER_13_2457 ();
 sg13g2_decap_8 FILLER_13_2464 ();
 sg13g2_decap_8 FILLER_13_2471 ();
 sg13g2_decap_8 FILLER_13_2478 ();
 sg13g2_decap_8 FILLER_13_2485 ();
 sg13g2_decap_8 FILLER_13_2492 ();
 sg13g2_decap_8 FILLER_13_2499 ();
 sg13g2_decap_8 FILLER_13_2506 ();
 sg13g2_decap_8 FILLER_13_2513 ();
 sg13g2_decap_8 FILLER_13_2520 ();
 sg13g2_decap_8 FILLER_13_2527 ();
 sg13g2_decap_8 FILLER_13_2534 ();
 sg13g2_decap_8 FILLER_13_2541 ();
 sg13g2_decap_8 FILLER_13_2548 ();
 sg13g2_decap_8 FILLER_13_2555 ();
 sg13g2_decap_8 FILLER_13_2562 ();
 sg13g2_decap_8 FILLER_13_2569 ();
 sg13g2_decap_8 FILLER_13_2576 ();
 sg13g2_decap_8 FILLER_13_2583 ();
 sg13g2_decap_8 FILLER_13_2590 ();
 sg13g2_decap_8 FILLER_13_2597 ();
 sg13g2_decap_8 FILLER_13_2604 ();
 sg13g2_decap_8 FILLER_13_2611 ();
 sg13g2_decap_8 FILLER_13_2618 ();
 sg13g2_decap_8 FILLER_13_2625 ();
 sg13g2_decap_8 FILLER_13_2632 ();
 sg13g2_decap_8 FILLER_13_2639 ();
 sg13g2_decap_8 FILLER_13_2646 ();
 sg13g2_decap_8 FILLER_13_2653 ();
 sg13g2_decap_8 FILLER_13_2660 ();
 sg13g2_decap_8 FILLER_13_2667 ();
 sg13g2_decap_8 FILLER_13_2674 ();
 sg13g2_decap_8 FILLER_13_2681 ();
 sg13g2_decap_8 FILLER_13_2688 ();
 sg13g2_decap_8 FILLER_13_2695 ();
 sg13g2_decap_8 FILLER_13_2702 ();
 sg13g2_decap_8 FILLER_13_2709 ();
 sg13g2_decap_8 FILLER_13_2716 ();
 sg13g2_decap_8 FILLER_13_2723 ();
 sg13g2_decap_8 FILLER_13_2730 ();
 sg13g2_decap_8 FILLER_13_2737 ();
 sg13g2_decap_8 FILLER_13_2744 ();
 sg13g2_decap_8 FILLER_13_2751 ();
 sg13g2_decap_8 FILLER_13_2758 ();
 sg13g2_decap_8 FILLER_13_2765 ();
 sg13g2_decap_8 FILLER_13_2772 ();
 sg13g2_decap_8 FILLER_13_2779 ();
 sg13g2_decap_8 FILLER_13_2786 ();
 sg13g2_decap_8 FILLER_13_2793 ();
 sg13g2_decap_8 FILLER_13_2800 ();
 sg13g2_decap_8 FILLER_13_2807 ();
 sg13g2_decap_8 FILLER_13_2814 ();
 sg13g2_decap_8 FILLER_13_2821 ();
 sg13g2_decap_8 FILLER_13_2828 ();
 sg13g2_decap_8 FILLER_13_2835 ();
 sg13g2_decap_8 FILLER_13_2842 ();
 sg13g2_decap_8 FILLER_13_2849 ();
 sg13g2_decap_8 FILLER_13_2856 ();
 sg13g2_decap_8 FILLER_13_2863 ();
 sg13g2_decap_8 FILLER_13_2870 ();
 sg13g2_decap_8 FILLER_13_2877 ();
 sg13g2_decap_8 FILLER_13_2884 ();
 sg13g2_decap_8 FILLER_13_2891 ();
 sg13g2_decap_8 FILLER_13_2898 ();
 sg13g2_decap_8 FILLER_13_2905 ();
 sg13g2_decap_8 FILLER_13_2912 ();
 sg13g2_decap_8 FILLER_13_2919 ();
 sg13g2_decap_8 FILLER_13_2926 ();
 sg13g2_decap_8 FILLER_13_2933 ();
 sg13g2_decap_8 FILLER_13_2940 ();
 sg13g2_decap_8 FILLER_13_2947 ();
 sg13g2_decap_8 FILLER_13_2954 ();
 sg13g2_decap_8 FILLER_13_2961 ();
 sg13g2_decap_8 FILLER_13_2968 ();
 sg13g2_decap_8 FILLER_13_2975 ();
 sg13g2_decap_8 FILLER_13_2982 ();
 sg13g2_decap_8 FILLER_13_2989 ();
 sg13g2_decap_8 FILLER_13_2996 ();
 sg13g2_decap_8 FILLER_13_3003 ();
 sg13g2_decap_8 FILLER_13_3010 ();
 sg13g2_decap_8 FILLER_13_3017 ();
 sg13g2_decap_8 FILLER_13_3024 ();
 sg13g2_decap_8 FILLER_13_3031 ();
 sg13g2_decap_8 FILLER_13_3038 ();
 sg13g2_decap_8 FILLER_13_3045 ();
 sg13g2_decap_8 FILLER_13_3052 ();
 sg13g2_decap_8 FILLER_13_3059 ();
 sg13g2_decap_8 FILLER_13_3066 ();
 sg13g2_decap_8 FILLER_13_3073 ();
 sg13g2_decap_8 FILLER_13_3080 ();
 sg13g2_decap_8 FILLER_13_3087 ();
 sg13g2_decap_8 FILLER_13_3094 ();
 sg13g2_decap_8 FILLER_13_3101 ();
 sg13g2_decap_8 FILLER_13_3108 ();
 sg13g2_decap_8 FILLER_13_3115 ();
 sg13g2_decap_8 FILLER_13_3122 ();
 sg13g2_decap_8 FILLER_13_3129 ();
 sg13g2_decap_8 FILLER_13_3136 ();
 sg13g2_decap_8 FILLER_13_3143 ();
 sg13g2_decap_8 FILLER_13_3150 ();
 sg13g2_decap_8 FILLER_13_3157 ();
 sg13g2_decap_8 FILLER_13_3164 ();
 sg13g2_decap_8 FILLER_13_3171 ();
 sg13g2_decap_8 FILLER_13_3178 ();
 sg13g2_decap_8 FILLER_13_3185 ();
 sg13g2_decap_8 FILLER_13_3192 ();
 sg13g2_decap_8 FILLER_13_3199 ();
 sg13g2_decap_8 FILLER_13_3206 ();
 sg13g2_decap_8 FILLER_13_3213 ();
 sg13g2_decap_8 FILLER_13_3220 ();
 sg13g2_decap_8 FILLER_13_3227 ();
 sg13g2_decap_8 FILLER_13_3234 ();
 sg13g2_decap_8 FILLER_13_3241 ();
 sg13g2_decap_8 FILLER_13_3248 ();
 sg13g2_decap_8 FILLER_13_3255 ();
 sg13g2_decap_8 FILLER_13_3262 ();
 sg13g2_decap_8 FILLER_13_3269 ();
 sg13g2_decap_8 FILLER_13_3276 ();
 sg13g2_decap_8 FILLER_13_3283 ();
 sg13g2_decap_8 FILLER_13_3290 ();
 sg13g2_decap_8 FILLER_13_3297 ();
 sg13g2_decap_8 FILLER_13_3304 ();
 sg13g2_decap_8 FILLER_13_3311 ();
 sg13g2_decap_8 FILLER_13_3318 ();
 sg13g2_decap_8 FILLER_13_3325 ();
 sg13g2_decap_8 FILLER_13_3332 ();
 sg13g2_decap_8 FILLER_13_3339 ();
 sg13g2_decap_8 FILLER_13_3346 ();
 sg13g2_decap_8 FILLER_13_3353 ();
 sg13g2_decap_8 FILLER_13_3360 ();
 sg13g2_decap_8 FILLER_13_3367 ();
 sg13g2_decap_8 FILLER_13_3374 ();
 sg13g2_decap_8 FILLER_13_3381 ();
 sg13g2_decap_8 FILLER_13_3388 ();
 sg13g2_decap_8 FILLER_13_3395 ();
 sg13g2_decap_8 FILLER_13_3402 ();
 sg13g2_decap_8 FILLER_13_3409 ();
 sg13g2_decap_8 FILLER_13_3416 ();
 sg13g2_decap_8 FILLER_13_3423 ();
 sg13g2_decap_8 FILLER_13_3430 ();
 sg13g2_decap_8 FILLER_13_3437 ();
 sg13g2_decap_8 FILLER_13_3444 ();
 sg13g2_decap_8 FILLER_13_3451 ();
 sg13g2_decap_8 FILLER_13_3458 ();
 sg13g2_decap_8 FILLER_13_3465 ();
 sg13g2_decap_8 FILLER_13_3472 ();
 sg13g2_decap_8 FILLER_13_3479 ();
 sg13g2_decap_8 FILLER_13_3486 ();
 sg13g2_decap_8 FILLER_13_3493 ();
 sg13g2_decap_8 FILLER_13_3500 ();
 sg13g2_decap_8 FILLER_13_3507 ();
 sg13g2_decap_8 FILLER_13_3514 ();
 sg13g2_decap_8 FILLER_13_3521 ();
 sg13g2_decap_8 FILLER_13_3528 ();
 sg13g2_decap_8 FILLER_13_3535 ();
 sg13g2_decap_8 FILLER_13_3542 ();
 sg13g2_decap_8 FILLER_13_3549 ();
 sg13g2_decap_8 FILLER_13_3556 ();
 sg13g2_decap_8 FILLER_13_3563 ();
 sg13g2_decap_8 FILLER_13_3570 ();
 sg13g2_fill_2 FILLER_13_3577 ();
 sg13g2_fill_1 FILLER_13_3579 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_decap_8 FILLER_14_483 ();
 sg13g2_decap_8 FILLER_14_490 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_decap_8 FILLER_14_504 ();
 sg13g2_decap_8 FILLER_14_511 ();
 sg13g2_decap_8 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_525 ();
 sg13g2_decap_8 FILLER_14_532 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_decap_8 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_decap_8 FILLER_14_560 ();
 sg13g2_decap_8 FILLER_14_567 ();
 sg13g2_decap_8 FILLER_14_574 ();
 sg13g2_decap_8 FILLER_14_581 ();
 sg13g2_decap_8 FILLER_14_588 ();
 sg13g2_decap_8 FILLER_14_595 ();
 sg13g2_decap_8 FILLER_14_602 ();
 sg13g2_decap_8 FILLER_14_609 ();
 sg13g2_decap_8 FILLER_14_616 ();
 sg13g2_decap_8 FILLER_14_623 ();
 sg13g2_decap_8 FILLER_14_630 ();
 sg13g2_decap_8 FILLER_14_637 ();
 sg13g2_decap_8 FILLER_14_644 ();
 sg13g2_decap_8 FILLER_14_651 ();
 sg13g2_decap_8 FILLER_14_658 ();
 sg13g2_decap_8 FILLER_14_665 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_decap_8 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_686 ();
 sg13g2_decap_8 FILLER_14_693 ();
 sg13g2_decap_8 FILLER_14_700 ();
 sg13g2_decap_8 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_714 ();
 sg13g2_decap_8 FILLER_14_721 ();
 sg13g2_decap_8 FILLER_14_728 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_decap_8 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_8 FILLER_14_777 ();
 sg13g2_decap_8 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_8 FILLER_14_805 ();
 sg13g2_decap_8 FILLER_14_812 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_decap_8 FILLER_14_826 ();
 sg13g2_decap_8 FILLER_14_833 ();
 sg13g2_decap_8 FILLER_14_840 ();
 sg13g2_decap_8 FILLER_14_847 ();
 sg13g2_decap_8 FILLER_14_854 ();
 sg13g2_decap_8 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_14_868 ();
 sg13g2_decap_8 FILLER_14_875 ();
 sg13g2_decap_8 FILLER_14_882 ();
 sg13g2_decap_8 FILLER_14_889 ();
 sg13g2_decap_8 FILLER_14_896 ();
 sg13g2_decap_8 FILLER_14_903 ();
 sg13g2_decap_8 FILLER_14_910 ();
 sg13g2_decap_8 FILLER_14_917 ();
 sg13g2_decap_8 FILLER_14_924 ();
 sg13g2_decap_8 FILLER_14_931 ();
 sg13g2_decap_8 FILLER_14_938 ();
 sg13g2_decap_8 FILLER_14_945 ();
 sg13g2_decap_8 FILLER_14_952 ();
 sg13g2_decap_8 FILLER_14_959 ();
 sg13g2_decap_8 FILLER_14_966 ();
 sg13g2_decap_8 FILLER_14_973 ();
 sg13g2_decap_8 FILLER_14_980 ();
 sg13g2_decap_8 FILLER_14_987 ();
 sg13g2_decap_8 FILLER_14_994 ();
 sg13g2_decap_8 FILLER_14_1001 ();
 sg13g2_decap_8 FILLER_14_1008 ();
 sg13g2_decap_8 FILLER_14_1015 ();
 sg13g2_decap_8 FILLER_14_1022 ();
 sg13g2_decap_8 FILLER_14_1029 ();
 sg13g2_decap_8 FILLER_14_1036 ();
 sg13g2_decap_8 FILLER_14_1043 ();
 sg13g2_decap_8 FILLER_14_1050 ();
 sg13g2_decap_8 FILLER_14_1057 ();
 sg13g2_decap_8 FILLER_14_1064 ();
 sg13g2_decap_8 FILLER_14_1071 ();
 sg13g2_decap_8 FILLER_14_1078 ();
 sg13g2_decap_8 FILLER_14_1085 ();
 sg13g2_decap_8 FILLER_14_1092 ();
 sg13g2_decap_8 FILLER_14_1099 ();
 sg13g2_decap_8 FILLER_14_1106 ();
 sg13g2_decap_8 FILLER_14_1113 ();
 sg13g2_decap_8 FILLER_14_1120 ();
 sg13g2_decap_8 FILLER_14_1127 ();
 sg13g2_decap_8 FILLER_14_1134 ();
 sg13g2_decap_8 FILLER_14_1141 ();
 sg13g2_decap_8 FILLER_14_1148 ();
 sg13g2_decap_8 FILLER_14_1155 ();
 sg13g2_decap_8 FILLER_14_1162 ();
 sg13g2_decap_8 FILLER_14_1169 ();
 sg13g2_decap_8 FILLER_14_1176 ();
 sg13g2_decap_8 FILLER_14_1183 ();
 sg13g2_decap_8 FILLER_14_1190 ();
 sg13g2_decap_8 FILLER_14_1197 ();
 sg13g2_decap_8 FILLER_14_1204 ();
 sg13g2_decap_8 FILLER_14_1211 ();
 sg13g2_decap_8 FILLER_14_1218 ();
 sg13g2_decap_8 FILLER_14_1225 ();
 sg13g2_decap_8 FILLER_14_1232 ();
 sg13g2_decap_8 FILLER_14_1239 ();
 sg13g2_decap_8 FILLER_14_1246 ();
 sg13g2_decap_8 FILLER_14_1253 ();
 sg13g2_decap_8 FILLER_14_1260 ();
 sg13g2_decap_8 FILLER_14_1267 ();
 sg13g2_decap_8 FILLER_14_1274 ();
 sg13g2_decap_8 FILLER_14_1281 ();
 sg13g2_decap_8 FILLER_14_1288 ();
 sg13g2_decap_8 FILLER_14_1295 ();
 sg13g2_decap_8 FILLER_14_1302 ();
 sg13g2_decap_8 FILLER_14_1309 ();
 sg13g2_decap_8 FILLER_14_1316 ();
 sg13g2_decap_8 FILLER_14_1323 ();
 sg13g2_decap_8 FILLER_14_1330 ();
 sg13g2_decap_8 FILLER_14_1337 ();
 sg13g2_decap_8 FILLER_14_1344 ();
 sg13g2_decap_8 FILLER_14_1351 ();
 sg13g2_decap_8 FILLER_14_1358 ();
 sg13g2_decap_8 FILLER_14_1365 ();
 sg13g2_decap_8 FILLER_14_1372 ();
 sg13g2_decap_8 FILLER_14_1379 ();
 sg13g2_decap_8 FILLER_14_1386 ();
 sg13g2_decap_8 FILLER_14_1393 ();
 sg13g2_decap_8 FILLER_14_1400 ();
 sg13g2_decap_8 FILLER_14_1407 ();
 sg13g2_decap_8 FILLER_14_1414 ();
 sg13g2_decap_8 FILLER_14_1421 ();
 sg13g2_decap_8 FILLER_14_1428 ();
 sg13g2_decap_8 FILLER_14_1435 ();
 sg13g2_decap_8 FILLER_14_1442 ();
 sg13g2_decap_8 FILLER_14_1449 ();
 sg13g2_decap_8 FILLER_14_1456 ();
 sg13g2_decap_8 FILLER_14_1463 ();
 sg13g2_decap_8 FILLER_14_1470 ();
 sg13g2_decap_8 FILLER_14_1477 ();
 sg13g2_decap_8 FILLER_14_1484 ();
 sg13g2_decap_8 FILLER_14_1491 ();
 sg13g2_decap_8 FILLER_14_1498 ();
 sg13g2_decap_8 FILLER_14_1505 ();
 sg13g2_decap_8 FILLER_14_1512 ();
 sg13g2_decap_8 FILLER_14_1519 ();
 sg13g2_decap_8 FILLER_14_1526 ();
 sg13g2_decap_8 FILLER_14_1533 ();
 sg13g2_decap_8 FILLER_14_1540 ();
 sg13g2_decap_8 FILLER_14_1547 ();
 sg13g2_decap_8 FILLER_14_1554 ();
 sg13g2_decap_8 FILLER_14_1561 ();
 sg13g2_decap_8 FILLER_14_1568 ();
 sg13g2_decap_8 FILLER_14_1575 ();
 sg13g2_decap_8 FILLER_14_1582 ();
 sg13g2_decap_8 FILLER_14_1589 ();
 sg13g2_decap_8 FILLER_14_1596 ();
 sg13g2_decap_8 FILLER_14_1603 ();
 sg13g2_decap_8 FILLER_14_1610 ();
 sg13g2_decap_8 FILLER_14_1617 ();
 sg13g2_decap_8 FILLER_14_1624 ();
 sg13g2_decap_8 FILLER_14_1631 ();
 sg13g2_decap_8 FILLER_14_1638 ();
 sg13g2_decap_8 FILLER_14_1645 ();
 sg13g2_decap_8 FILLER_14_1652 ();
 sg13g2_decap_8 FILLER_14_1659 ();
 sg13g2_decap_8 FILLER_14_1666 ();
 sg13g2_decap_8 FILLER_14_1673 ();
 sg13g2_decap_8 FILLER_14_1680 ();
 sg13g2_decap_8 FILLER_14_1687 ();
 sg13g2_decap_8 FILLER_14_1694 ();
 sg13g2_decap_8 FILLER_14_1701 ();
 sg13g2_decap_8 FILLER_14_1708 ();
 sg13g2_decap_8 FILLER_14_1715 ();
 sg13g2_decap_8 FILLER_14_1722 ();
 sg13g2_decap_8 FILLER_14_1729 ();
 sg13g2_decap_8 FILLER_14_1736 ();
 sg13g2_decap_8 FILLER_14_1743 ();
 sg13g2_decap_8 FILLER_14_1750 ();
 sg13g2_decap_8 FILLER_14_1757 ();
 sg13g2_decap_8 FILLER_14_1764 ();
 sg13g2_decap_8 FILLER_14_1771 ();
 sg13g2_decap_8 FILLER_14_1778 ();
 sg13g2_decap_8 FILLER_14_1785 ();
 sg13g2_decap_8 FILLER_14_1792 ();
 sg13g2_decap_8 FILLER_14_1799 ();
 sg13g2_decap_8 FILLER_14_1806 ();
 sg13g2_decap_8 FILLER_14_1813 ();
 sg13g2_decap_8 FILLER_14_1820 ();
 sg13g2_decap_8 FILLER_14_1827 ();
 sg13g2_decap_8 FILLER_14_1834 ();
 sg13g2_decap_8 FILLER_14_1841 ();
 sg13g2_decap_8 FILLER_14_1848 ();
 sg13g2_decap_8 FILLER_14_1855 ();
 sg13g2_decap_8 FILLER_14_1862 ();
 sg13g2_decap_8 FILLER_14_1869 ();
 sg13g2_decap_8 FILLER_14_1876 ();
 sg13g2_decap_8 FILLER_14_1883 ();
 sg13g2_decap_8 FILLER_14_1890 ();
 sg13g2_decap_8 FILLER_14_1897 ();
 sg13g2_decap_8 FILLER_14_1904 ();
 sg13g2_decap_8 FILLER_14_1911 ();
 sg13g2_decap_8 FILLER_14_1918 ();
 sg13g2_decap_8 FILLER_14_1925 ();
 sg13g2_decap_8 FILLER_14_1932 ();
 sg13g2_decap_8 FILLER_14_1939 ();
 sg13g2_decap_8 FILLER_14_1946 ();
 sg13g2_decap_8 FILLER_14_1953 ();
 sg13g2_decap_8 FILLER_14_1960 ();
 sg13g2_decap_8 FILLER_14_1967 ();
 sg13g2_decap_8 FILLER_14_1974 ();
 sg13g2_decap_8 FILLER_14_1981 ();
 sg13g2_decap_8 FILLER_14_1988 ();
 sg13g2_decap_8 FILLER_14_1995 ();
 sg13g2_decap_8 FILLER_14_2002 ();
 sg13g2_decap_8 FILLER_14_2009 ();
 sg13g2_decap_8 FILLER_14_2016 ();
 sg13g2_decap_8 FILLER_14_2023 ();
 sg13g2_decap_8 FILLER_14_2030 ();
 sg13g2_decap_8 FILLER_14_2037 ();
 sg13g2_decap_8 FILLER_14_2044 ();
 sg13g2_decap_8 FILLER_14_2051 ();
 sg13g2_decap_8 FILLER_14_2058 ();
 sg13g2_decap_8 FILLER_14_2065 ();
 sg13g2_decap_8 FILLER_14_2072 ();
 sg13g2_decap_8 FILLER_14_2079 ();
 sg13g2_decap_8 FILLER_14_2086 ();
 sg13g2_decap_8 FILLER_14_2093 ();
 sg13g2_decap_8 FILLER_14_2100 ();
 sg13g2_decap_8 FILLER_14_2107 ();
 sg13g2_decap_8 FILLER_14_2114 ();
 sg13g2_decap_8 FILLER_14_2121 ();
 sg13g2_decap_8 FILLER_14_2128 ();
 sg13g2_decap_8 FILLER_14_2135 ();
 sg13g2_decap_8 FILLER_14_2142 ();
 sg13g2_decap_8 FILLER_14_2149 ();
 sg13g2_decap_8 FILLER_14_2156 ();
 sg13g2_decap_8 FILLER_14_2163 ();
 sg13g2_decap_8 FILLER_14_2170 ();
 sg13g2_decap_8 FILLER_14_2177 ();
 sg13g2_decap_8 FILLER_14_2184 ();
 sg13g2_decap_8 FILLER_14_2191 ();
 sg13g2_decap_8 FILLER_14_2198 ();
 sg13g2_decap_8 FILLER_14_2205 ();
 sg13g2_decap_8 FILLER_14_2212 ();
 sg13g2_decap_8 FILLER_14_2219 ();
 sg13g2_decap_8 FILLER_14_2226 ();
 sg13g2_decap_8 FILLER_14_2233 ();
 sg13g2_decap_8 FILLER_14_2240 ();
 sg13g2_decap_8 FILLER_14_2247 ();
 sg13g2_decap_8 FILLER_14_2254 ();
 sg13g2_decap_8 FILLER_14_2261 ();
 sg13g2_decap_8 FILLER_14_2268 ();
 sg13g2_decap_8 FILLER_14_2275 ();
 sg13g2_decap_8 FILLER_14_2282 ();
 sg13g2_decap_8 FILLER_14_2289 ();
 sg13g2_decap_8 FILLER_14_2296 ();
 sg13g2_decap_8 FILLER_14_2303 ();
 sg13g2_decap_8 FILLER_14_2310 ();
 sg13g2_decap_8 FILLER_14_2317 ();
 sg13g2_decap_8 FILLER_14_2324 ();
 sg13g2_decap_8 FILLER_14_2331 ();
 sg13g2_decap_8 FILLER_14_2338 ();
 sg13g2_decap_8 FILLER_14_2345 ();
 sg13g2_decap_8 FILLER_14_2352 ();
 sg13g2_decap_8 FILLER_14_2359 ();
 sg13g2_decap_8 FILLER_14_2366 ();
 sg13g2_decap_8 FILLER_14_2373 ();
 sg13g2_decap_8 FILLER_14_2380 ();
 sg13g2_decap_8 FILLER_14_2387 ();
 sg13g2_decap_8 FILLER_14_2394 ();
 sg13g2_decap_8 FILLER_14_2401 ();
 sg13g2_decap_8 FILLER_14_2408 ();
 sg13g2_decap_8 FILLER_14_2415 ();
 sg13g2_decap_8 FILLER_14_2422 ();
 sg13g2_decap_8 FILLER_14_2429 ();
 sg13g2_decap_8 FILLER_14_2436 ();
 sg13g2_decap_8 FILLER_14_2443 ();
 sg13g2_decap_8 FILLER_14_2450 ();
 sg13g2_decap_8 FILLER_14_2457 ();
 sg13g2_decap_8 FILLER_14_2464 ();
 sg13g2_decap_8 FILLER_14_2471 ();
 sg13g2_decap_8 FILLER_14_2478 ();
 sg13g2_decap_8 FILLER_14_2485 ();
 sg13g2_decap_8 FILLER_14_2492 ();
 sg13g2_decap_8 FILLER_14_2499 ();
 sg13g2_decap_8 FILLER_14_2506 ();
 sg13g2_decap_8 FILLER_14_2513 ();
 sg13g2_decap_8 FILLER_14_2520 ();
 sg13g2_decap_8 FILLER_14_2527 ();
 sg13g2_decap_8 FILLER_14_2534 ();
 sg13g2_decap_8 FILLER_14_2541 ();
 sg13g2_decap_8 FILLER_14_2548 ();
 sg13g2_decap_8 FILLER_14_2555 ();
 sg13g2_decap_8 FILLER_14_2562 ();
 sg13g2_decap_8 FILLER_14_2569 ();
 sg13g2_decap_8 FILLER_14_2576 ();
 sg13g2_decap_8 FILLER_14_2583 ();
 sg13g2_decap_8 FILLER_14_2590 ();
 sg13g2_decap_8 FILLER_14_2597 ();
 sg13g2_decap_8 FILLER_14_2604 ();
 sg13g2_decap_8 FILLER_14_2611 ();
 sg13g2_decap_8 FILLER_14_2618 ();
 sg13g2_decap_8 FILLER_14_2625 ();
 sg13g2_decap_8 FILLER_14_2632 ();
 sg13g2_decap_8 FILLER_14_2639 ();
 sg13g2_decap_8 FILLER_14_2646 ();
 sg13g2_decap_8 FILLER_14_2653 ();
 sg13g2_decap_8 FILLER_14_2660 ();
 sg13g2_decap_8 FILLER_14_2667 ();
 sg13g2_decap_8 FILLER_14_2674 ();
 sg13g2_decap_8 FILLER_14_2681 ();
 sg13g2_decap_8 FILLER_14_2688 ();
 sg13g2_decap_8 FILLER_14_2695 ();
 sg13g2_decap_8 FILLER_14_2702 ();
 sg13g2_decap_8 FILLER_14_2709 ();
 sg13g2_decap_8 FILLER_14_2716 ();
 sg13g2_decap_8 FILLER_14_2723 ();
 sg13g2_decap_8 FILLER_14_2730 ();
 sg13g2_decap_8 FILLER_14_2737 ();
 sg13g2_decap_8 FILLER_14_2744 ();
 sg13g2_decap_8 FILLER_14_2751 ();
 sg13g2_decap_8 FILLER_14_2758 ();
 sg13g2_decap_8 FILLER_14_2765 ();
 sg13g2_decap_8 FILLER_14_2772 ();
 sg13g2_decap_8 FILLER_14_2779 ();
 sg13g2_decap_8 FILLER_14_2786 ();
 sg13g2_decap_8 FILLER_14_2793 ();
 sg13g2_decap_8 FILLER_14_2800 ();
 sg13g2_decap_8 FILLER_14_2807 ();
 sg13g2_decap_8 FILLER_14_2814 ();
 sg13g2_decap_8 FILLER_14_2821 ();
 sg13g2_decap_8 FILLER_14_2828 ();
 sg13g2_decap_8 FILLER_14_2835 ();
 sg13g2_decap_8 FILLER_14_2842 ();
 sg13g2_decap_8 FILLER_14_2849 ();
 sg13g2_decap_8 FILLER_14_2856 ();
 sg13g2_decap_8 FILLER_14_2863 ();
 sg13g2_decap_8 FILLER_14_2870 ();
 sg13g2_decap_8 FILLER_14_2877 ();
 sg13g2_decap_8 FILLER_14_2884 ();
 sg13g2_decap_8 FILLER_14_2891 ();
 sg13g2_decap_8 FILLER_14_2898 ();
 sg13g2_decap_8 FILLER_14_2905 ();
 sg13g2_decap_8 FILLER_14_2912 ();
 sg13g2_decap_8 FILLER_14_2919 ();
 sg13g2_decap_8 FILLER_14_2926 ();
 sg13g2_decap_8 FILLER_14_2933 ();
 sg13g2_decap_8 FILLER_14_2940 ();
 sg13g2_decap_8 FILLER_14_2947 ();
 sg13g2_decap_8 FILLER_14_2954 ();
 sg13g2_decap_8 FILLER_14_2961 ();
 sg13g2_decap_8 FILLER_14_2968 ();
 sg13g2_decap_8 FILLER_14_2975 ();
 sg13g2_decap_8 FILLER_14_2982 ();
 sg13g2_decap_8 FILLER_14_2989 ();
 sg13g2_decap_8 FILLER_14_2996 ();
 sg13g2_decap_8 FILLER_14_3003 ();
 sg13g2_decap_8 FILLER_14_3010 ();
 sg13g2_decap_8 FILLER_14_3017 ();
 sg13g2_decap_8 FILLER_14_3024 ();
 sg13g2_decap_8 FILLER_14_3031 ();
 sg13g2_decap_8 FILLER_14_3038 ();
 sg13g2_decap_8 FILLER_14_3045 ();
 sg13g2_decap_8 FILLER_14_3052 ();
 sg13g2_decap_8 FILLER_14_3059 ();
 sg13g2_decap_8 FILLER_14_3066 ();
 sg13g2_decap_8 FILLER_14_3073 ();
 sg13g2_decap_8 FILLER_14_3080 ();
 sg13g2_decap_8 FILLER_14_3087 ();
 sg13g2_decap_8 FILLER_14_3094 ();
 sg13g2_decap_8 FILLER_14_3101 ();
 sg13g2_decap_8 FILLER_14_3108 ();
 sg13g2_decap_8 FILLER_14_3115 ();
 sg13g2_decap_8 FILLER_14_3122 ();
 sg13g2_decap_8 FILLER_14_3129 ();
 sg13g2_decap_8 FILLER_14_3136 ();
 sg13g2_decap_8 FILLER_14_3143 ();
 sg13g2_decap_8 FILLER_14_3150 ();
 sg13g2_decap_8 FILLER_14_3157 ();
 sg13g2_decap_8 FILLER_14_3164 ();
 sg13g2_decap_8 FILLER_14_3171 ();
 sg13g2_decap_8 FILLER_14_3178 ();
 sg13g2_decap_8 FILLER_14_3185 ();
 sg13g2_decap_8 FILLER_14_3192 ();
 sg13g2_decap_8 FILLER_14_3199 ();
 sg13g2_decap_8 FILLER_14_3206 ();
 sg13g2_decap_8 FILLER_14_3213 ();
 sg13g2_decap_8 FILLER_14_3220 ();
 sg13g2_decap_8 FILLER_14_3227 ();
 sg13g2_decap_8 FILLER_14_3234 ();
 sg13g2_decap_8 FILLER_14_3241 ();
 sg13g2_decap_8 FILLER_14_3248 ();
 sg13g2_decap_8 FILLER_14_3255 ();
 sg13g2_decap_8 FILLER_14_3262 ();
 sg13g2_decap_8 FILLER_14_3269 ();
 sg13g2_decap_8 FILLER_14_3276 ();
 sg13g2_decap_8 FILLER_14_3283 ();
 sg13g2_decap_8 FILLER_14_3290 ();
 sg13g2_decap_8 FILLER_14_3297 ();
 sg13g2_decap_8 FILLER_14_3304 ();
 sg13g2_decap_8 FILLER_14_3311 ();
 sg13g2_decap_8 FILLER_14_3318 ();
 sg13g2_decap_8 FILLER_14_3325 ();
 sg13g2_decap_8 FILLER_14_3332 ();
 sg13g2_decap_8 FILLER_14_3339 ();
 sg13g2_decap_8 FILLER_14_3346 ();
 sg13g2_decap_8 FILLER_14_3353 ();
 sg13g2_decap_8 FILLER_14_3360 ();
 sg13g2_decap_8 FILLER_14_3367 ();
 sg13g2_decap_8 FILLER_14_3374 ();
 sg13g2_decap_8 FILLER_14_3381 ();
 sg13g2_decap_8 FILLER_14_3388 ();
 sg13g2_decap_8 FILLER_14_3395 ();
 sg13g2_decap_8 FILLER_14_3402 ();
 sg13g2_decap_8 FILLER_14_3409 ();
 sg13g2_decap_8 FILLER_14_3416 ();
 sg13g2_decap_8 FILLER_14_3423 ();
 sg13g2_decap_8 FILLER_14_3430 ();
 sg13g2_decap_8 FILLER_14_3437 ();
 sg13g2_decap_8 FILLER_14_3444 ();
 sg13g2_decap_8 FILLER_14_3451 ();
 sg13g2_decap_8 FILLER_14_3458 ();
 sg13g2_decap_8 FILLER_14_3465 ();
 sg13g2_decap_8 FILLER_14_3472 ();
 sg13g2_decap_8 FILLER_14_3479 ();
 sg13g2_decap_8 FILLER_14_3486 ();
 sg13g2_decap_8 FILLER_14_3493 ();
 sg13g2_decap_8 FILLER_14_3500 ();
 sg13g2_decap_8 FILLER_14_3507 ();
 sg13g2_decap_8 FILLER_14_3514 ();
 sg13g2_decap_8 FILLER_14_3521 ();
 sg13g2_decap_8 FILLER_14_3528 ();
 sg13g2_decap_8 FILLER_14_3535 ();
 sg13g2_decap_8 FILLER_14_3542 ();
 sg13g2_decap_8 FILLER_14_3549 ();
 sg13g2_decap_8 FILLER_14_3556 ();
 sg13g2_decap_8 FILLER_14_3563 ();
 sg13g2_decap_8 FILLER_14_3570 ();
 sg13g2_fill_2 FILLER_14_3577 ();
 sg13g2_fill_1 FILLER_14_3579 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_decap_8 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_434 ();
 sg13g2_decap_8 FILLER_15_441 ();
 sg13g2_decap_8 FILLER_15_448 ();
 sg13g2_decap_8 FILLER_15_455 ();
 sg13g2_decap_8 FILLER_15_462 ();
 sg13g2_decap_8 FILLER_15_469 ();
 sg13g2_decap_8 FILLER_15_476 ();
 sg13g2_decap_8 FILLER_15_483 ();
 sg13g2_decap_8 FILLER_15_490 ();
 sg13g2_decap_8 FILLER_15_497 ();
 sg13g2_decap_8 FILLER_15_504 ();
 sg13g2_decap_8 FILLER_15_511 ();
 sg13g2_decap_8 FILLER_15_518 ();
 sg13g2_decap_8 FILLER_15_525 ();
 sg13g2_decap_8 FILLER_15_532 ();
 sg13g2_decap_8 FILLER_15_539 ();
 sg13g2_decap_8 FILLER_15_546 ();
 sg13g2_decap_8 FILLER_15_553 ();
 sg13g2_decap_8 FILLER_15_560 ();
 sg13g2_decap_8 FILLER_15_567 ();
 sg13g2_decap_8 FILLER_15_574 ();
 sg13g2_decap_8 FILLER_15_581 ();
 sg13g2_decap_8 FILLER_15_588 ();
 sg13g2_decap_8 FILLER_15_595 ();
 sg13g2_decap_8 FILLER_15_602 ();
 sg13g2_decap_8 FILLER_15_609 ();
 sg13g2_decap_8 FILLER_15_616 ();
 sg13g2_decap_8 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_630 ();
 sg13g2_decap_8 FILLER_15_637 ();
 sg13g2_decap_8 FILLER_15_644 ();
 sg13g2_decap_8 FILLER_15_651 ();
 sg13g2_decap_8 FILLER_15_658 ();
 sg13g2_decap_8 FILLER_15_665 ();
 sg13g2_decap_8 FILLER_15_672 ();
 sg13g2_decap_8 FILLER_15_679 ();
 sg13g2_decap_8 FILLER_15_686 ();
 sg13g2_decap_8 FILLER_15_693 ();
 sg13g2_decap_8 FILLER_15_700 ();
 sg13g2_decap_8 FILLER_15_707 ();
 sg13g2_decap_8 FILLER_15_714 ();
 sg13g2_decap_8 FILLER_15_721 ();
 sg13g2_decap_8 FILLER_15_728 ();
 sg13g2_decap_8 FILLER_15_735 ();
 sg13g2_decap_8 FILLER_15_742 ();
 sg13g2_decap_8 FILLER_15_749 ();
 sg13g2_decap_8 FILLER_15_756 ();
 sg13g2_decap_8 FILLER_15_763 ();
 sg13g2_decap_8 FILLER_15_770 ();
 sg13g2_decap_8 FILLER_15_777 ();
 sg13g2_decap_8 FILLER_15_784 ();
 sg13g2_decap_8 FILLER_15_791 ();
 sg13g2_decap_8 FILLER_15_798 ();
 sg13g2_decap_8 FILLER_15_805 ();
 sg13g2_decap_8 FILLER_15_812 ();
 sg13g2_decap_8 FILLER_15_819 ();
 sg13g2_decap_8 FILLER_15_826 ();
 sg13g2_decap_8 FILLER_15_833 ();
 sg13g2_decap_8 FILLER_15_840 ();
 sg13g2_decap_8 FILLER_15_847 ();
 sg13g2_decap_8 FILLER_15_854 ();
 sg13g2_decap_8 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_15_868 ();
 sg13g2_decap_8 FILLER_15_875 ();
 sg13g2_decap_8 FILLER_15_882 ();
 sg13g2_decap_8 FILLER_15_889 ();
 sg13g2_decap_8 FILLER_15_896 ();
 sg13g2_decap_8 FILLER_15_903 ();
 sg13g2_decap_8 FILLER_15_910 ();
 sg13g2_decap_8 FILLER_15_917 ();
 sg13g2_decap_8 FILLER_15_924 ();
 sg13g2_decap_8 FILLER_15_931 ();
 sg13g2_decap_8 FILLER_15_938 ();
 sg13g2_decap_8 FILLER_15_945 ();
 sg13g2_decap_8 FILLER_15_952 ();
 sg13g2_decap_8 FILLER_15_959 ();
 sg13g2_decap_8 FILLER_15_966 ();
 sg13g2_decap_8 FILLER_15_973 ();
 sg13g2_decap_8 FILLER_15_980 ();
 sg13g2_decap_8 FILLER_15_987 ();
 sg13g2_decap_8 FILLER_15_994 ();
 sg13g2_decap_8 FILLER_15_1001 ();
 sg13g2_decap_8 FILLER_15_1008 ();
 sg13g2_decap_8 FILLER_15_1015 ();
 sg13g2_decap_8 FILLER_15_1022 ();
 sg13g2_decap_8 FILLER_15_1029 ();
 sg13g2_decap_8 FILLER_15_1036 ();
 sg13g2_decap_8 FILLER_15_1043 ();
 sg13g2_decap_8 FILLER_15_1050 ();
 sg13g2_decap_8 FILLER_15_1057 ();
 sg13g2_decap_8 FILLER_15_1064 ();
 sg13g2_decap_8 FILLER_15_1071 ();
 sg13g2_decap_8 FILLER_15_1078 ();
 sg13g2_decap_8 FILLER_15_1085 ();
 sg13g2_decap_8 FILLER_15_1092 ();
 sg13g2_decap_8 FILLER_15_1099 ();
 sg13g2_decap_8 FILLER_15_1106 ();
 sg13g2_decap_8 FILLER_15_1113 ();
 sg13g2_decap_8 FILLER_15_1120 ();
 sg13g2_decap_8 FILLER_15_1127 ();
 sg13g2_decap_8 FILLER_15_1134 ();
 sg13g2_decap_8 FILLER_15_1141 ();
 sg13g2_decap_8 FILLER_15_1148 ();
 sg13g2_decap_8 FILLER_15_1155 ();
 sg13g2_decap_8 FILLER_15_1162 ();
 sg13g2_decap_8 FILLER_15_1169 ();
 sg13g2_decap_8 FILLER_15_1176 ();
 sg13g2_decap_8 FILLER_15_1183 ();
 sg13g2_decap_8 FILLER_15_1190 ();
 sg13g2_decap_8 FILLER_15_1197 ();
 sg13g2_decap_8 FILLER_15_1204 ();
 sg13g2_decap_8 FILLER_15_1211 ();
 sg13g2_decap_8 FILLER_15_1218 ();
 sg13g2_decap_8 FILLER_15_1225 ();
 sg13g2_decap_8 FILLER_15_1232 ();
 sg13g2_decap_8 FILLER_15_1239 ();
 sg13g2_decap_8 FILLER_15_1246 ();
 sg13g2_decap_8 FILLER_15_1253 ();
 sg13g2_decap_8 FILLER_15_1260 ();
 sg13g2_decap_8 FILLER_15_1267 ();
 sg13g2_decap_8 FILLER_15_1274 ();
 sg13g2_decap_8 FILLER_15_1281 ();
 sg13g2_decap_8 FILLER_15_1288 ();
 sg13g2_decap_8 FILLER_15_1295 ();
 sg13g2_decap_8 FILLER_15_1302 ();
 sg13g2_decap_8 FILLER_15_1309 ();
 sg13g2_decap_8 FILLER_15_1316 ();
 sg13g2_decap_8 FILLER_15_1323 ();
 sg13g2_decap_8 FILLER_15_1330 ();
 sg13g2_decap_8 FILLER_15_1337 ();
 sg13g2_decap_8 FILLER_15_1344 ();
 sg13g2_decap_8 FILLER_15_1351 ();
 sg13g2_decap_8 FILLER_15_1358 ();
 sg13g2_decap_8 FILLER_15_1365 ();
 sg13g2_decap_8 FILLER_15_1372 ();
 sg13g2_decap_8 FILLER_15_1379 ();
 sg13g2_decap_8 FILLER_15_1386 ();
 sg13g2_decap_8 FILLER_15_1393 ();
 sg13g2_decap_8 FILLER_15_1400 ();
 sg13g2_decap_8 FILLER_15_1407 ();
 sg13g2_decap_8 FILLER_15_1414 ();
 sg13g2_decap_8 FILLER_15_1421 ();
 sg13g2_decap_8 FILLER_15_1428 ();
 sg13g2_decap_8 FILLER_15_1435 ();
 sg13g2_decap_8 FILLER_15_1442 ();
 sg13g2_decap_8 FILLER_15_1449 ();
 sg13g2_decap_8 FILLER_15_1456 ();
 sg13g2_decap_8 FILLER_15_1463 ();
 sg13g2_decap_8 FILLER_15_1470 ();
 sg13g2_decap_8 FILLER_15_1477 ();
 sg13g2_decap_8 FILLER_15_1484 ();
 sg13g2_decap_8 FILLER_15_1491 ();
 sg13g2_decap_8 FILLER_15_1498 ();
 sg13g2_decap_8 FILLER_15_1505 ();
 sg13g2_decap_8 FILLER_15_1512 ();
 sg13g2_decap_8 FILLER_15_1519 ();
 sg13g2_decap_8 FILLER_15_1526 ();
 sg13g2_decap_8 FILLER_15_1533 ();
 sg13g2_decap_8 FILLER_15_1540 ();
 sg13g2_decap_8 FILLER_15_1547 ();
 sg13g2_decap_8 FILLER_15_1554 ();
 sg13g2_decap_8 FILLER_15_1561 ();
 sg13g2_decap_8 FILLER_15_1568 ();
 sg13g2_decap_8 FILLER_15_1575 ();
 sg13g2_decap_8 FILLER_15_1582 ();
 sg13g2_decap_8 FILLER_15_1589 ();
 sg13g2_decap_8 FILLER_15_1596 ();
 sg13g2_decap_8 FILLER_15_1603 ();
 sg13g2_decap_8 FILLER_15_1610 ();
 sg13g2_decap_8 FILLER_15_1617 ();
 sg13g2_decap_8 FILLER_15_1624 ();
 sg13g2_decap_8 FILLER_15_1631 ();
 sg13g2_decap_8 FILLER_15_1638 ();
 sg13g2_decap_8 FILLER_15_1645 ();
 sg13g2_decap_8 FILLER_15_1652 ();
 sg13g2_decap_8 FILLER_15_1659 ();
 sg13g2_decap_8 FILLER_15_1666 ();
 sg13g2_decap_8 FILLER_15_1673 ();
 sg13g2_decap_8 FILLER_15_1680 ();
 sg13g2_decap_8 FILLER_15_1687 ();
 sg13g2_decap_8 FILLER_15_1694 ();
 sg13g2_decap_8 FILLER_15_1701 ();
 sg13g2_decap_8 FILLER_15_1708 ();
 sg13g2_decap_8 FILLER_15_1715 ();
 sg13g2_decap_8 FILLER_15_1722 ();
 sg13g2_decap_8 FILLER_15_1729 ();
 sg13g2_decap_8 FILLER_15_1736 ();
 sg13g2_decap_8 FILLER_15_1743 ();
 sg13g2_decap_8 FILLER_15_1750 ();
 sg13g2_decap_8 FILLER_15_1757 ();
 sg13g2_decap_8 FILLER_15_1764 ();
 sg13g2_decap_8 FILLER_15_1771 ();
 sg13g2_decap_8 FILLER_15_1778 ();
 sg13g2_decap_8 FILLER_15_1785 ();
 sg13g2_decap_8 FILLER_15_1792 ();
 sg13g2_decap_8 FILLER_15_1799 ();
 sg13g2_decap_8 FILLER_15_1806 ();
 sg13g2_decap_8 FILLER_15_1813 ();
 sg13g2_decap_8 FILLER_15_1820 ();
 sg13g2_decap_8 FILLER_15_1827 ();
 sg13g2_decap_8 FILLER_15_1834 ();
 sg13g2_decap_8 FILLER_15_1841 ();
 sg13g2_decap_8 FILLER_15_1848 ();
 sg13g2_decap_8 FILLER_15_1855 ();
 sg13g2_decap_8 FILLER_15_1862 ();
 sg13g2_decap_8 FILLER_15_1869 ();
 sg13g2_decap_8 FILLER_15_1876 ();
 sg13g2_decap_8 FILLER_15_1883 ();
 sg13g2_decap_8 FILLER_15_1890 ();
 sg13g2_decap_8 FILLER_15_1897 ();
 sg13g2_decap_8 FILLER_15_1904 ();
 sg13g2_decap_8 FILLER_15_1911 ();
 sg13g2_decap_8 FILLER_15_1918 ();
 sg13g2_decap_8 FILLER_15_1925 ();
 sg13g2_decap_8 FILLER_15_1932 ();
 sg13g2_decap_8 FILLER_15_1939 ();
 sg13g2_decap_8 FILLER_15_1946 ();
 sg13g2_decap_8 FILLER_15_1953 ();
 sg13g2_decap_8 FILLER_15_1960 ();
 sg13g2_decap_8 FILLER_15_1967 ();
 sg13g2_decap_8 FILLER_15_1974 ();
 sg13g2_decap_8 FILLER_15_1981 ();
 sg13g2_decap_8 FILLER_15_1988 ();
 sg13g2_decap_8 FILLER_15_1995 ();
 sg13g2_decap_8 FILLER_15_2002 ();
 sg13g2_decap_8 FILLER_15_2009 ();
 sg13g2_decap_8 FILLER_15_2016 ();
 sg13g2_decap_8 FILLER_15_2023 ();
 sg13g2_decap_8 FILLER_15_2030 ();
 sg13g2_decap_8 FILLER_15_2037 ();
 sg13g2_decap_8 FILLER_15_2044 ();
 sg13g2_decap_8 FILLER_15_2051 ();
 sg13g2_decap_8 FILLER_15_2058 ();
 sg13g2_decap_8 FILLER_15_2065 ();
 sg13g2_decap_8 FILLER_15_2072 ();
 sg13g2_decap_8 FILLER_15_2079 ();
 sg13g2_decap_8 FILLER_15_2086 ();
 sg13g2_decap_8 FILLER_15_2093 ();
 sg13g2_decap_8 FILLER_15_2100 ();
 sg13g2_decap_8 FILLER_15_2107 ();
 sg13g2_decap_8 FILLER_15_2114 ();
 sg13g2_decap_8 FILLER_15_2121 ();
 sg13g2_decap_8 FILLER_15_2128 ();
 sg13g2_decap_8 FILLER_15_2135 ();
 sg13g2_decap_8 FILLER_15_2142 ();
 sg13g2_decap_8 FILLER_15_2149 ();
 sg13g2_decap_8 FILLER_15_2156 ();
 sg13g2_decap_8 FILLER_15_2163 ();
 sg13g2_decap_8 FILLER_15_2170 ();
 sg13g2_decap_8 FILLER_15_2177 ();
 sg13g2_decap_8 FILLER_15_2184 ();
 sg13g2_decap_8 FILLER_15_2191 ();
 sg13g2_decap_8 FILLER_15_2198 ();
 sg13g2_decap_8 FILLER_15_2205 ();
 sg13g2_decap_8 FILLER_15_2212 ();
 sg13g2_decap_8 FILLER_15_2219 ();
 sg13g2_decap_8 FILLER_15_2226 ();
 sg13g2_decap_8 FILLER_15_2233 ();
 sg13g2_decap_8 FILLER_15_2240 ();
 sg13g2_decap_8 FILLER_15_2247 ();
 sg13g2_decap_8 FILLER_15_2254 ();
 sg13g2_decap_8 FILLER_15_2261 ();
 sg13g2_decap_8 FILLER_15_2268 ();
 sg13g2_decap_8 FILLER_15_2275 ();
 sg13g2_decap_8 FILLER_15_2282 ();
 sg13g2_decap_8 FILLER_15_2289 ();
 sg13g2_decap_8 FILLER_15_2296 ();
 sg13g2_decap_8 FILLER_15_2303 ();
 sg13g2_decap_8 FILLER_15_2310 ();
 sg13g2_decap_8 FILLER_15_2317 ();
 sg13g2_decap_8 FILLER_15_2324 ();
 sg13g2_decap_8 FILLER_15_2331 ();
 sg13g2_decap_8 FILLER_15_2338 ();
 sg13g2_decap_8 FILLER_15_2345 ();
 sg13g2_decap_8 FILLER_15_2352 ();
 sg13g2_decap_8 FILLER_15_2359 ();
 sg13g2_decap_8 FILLER_15_2366 ();
 sg13g2_decap_8 FILLER_15_2373 ();
 sg13g2_decap_8 FILLER_15_2380 ();
 sg13g2_decap_8 FILLER_15_2387 ();
 sg13g2_decap_8 FILLER_15_2394 ();
 sg13g2_decap_8 FILLER_15_2401 ();
 sg13g2_decap_8 FILLER_15_2408 ();
 sg13g2_decap_8 FILLER_15_2415 ();
 sg13g2_decap_8 FILLER_15_2422 ();
 sg13g2_decap_8 FILLER_15_2429 ();
 sg13g2_decap_8 FILLER_15_2436 ();
 sg13g2_decap_8 FILLER_15_2443 ();
 sg13g2_decap_8 FILLER_15_2450 ();
 sg13g2_decap_8 FILLER_15_2457 ();
 sg13g2_decap_8 FILLER_15_2464 ();
 sg13g2_decap_8 FILLER_15_2471 ();
 sg13g2_decap_8 FILLER_15_2478 ();
 sg13g2_decap_8 FILLER_15_2485 ();
 sg13g2_decap_8 FILLER_15_2492 ();
 sg13g2_decap_8 FILLER_15_2499 ();
 sg13g2_decap_8 FILLER_15_2506 ();
 sg13g2_decap_8 FILLER_15_2513 ();
 sg13g2_decap_8 FILLER_15_2520 ();
 sg13g2_decap_8 FILLER_15_2527 ();
 sg13g2_decap_8 FILLER_15_2534 ();
 sg13g2_decap_8 FILLER_15_2541 ();
 sg13g2_decap_8 FILLER_15_2548 ();
 sg13g2_decap_8 FILLER_15_2555 ();
 sg13g2_decap_8 FILLER_15_2562 ();
 sg13g2_decap_8 FILLER_15_2569 ();
 sg13g2_decap_8 FILLER_15_2576 ();
 sg13g2_decap_8 FILLER_15_2583 ();
 sg13g2_decap_8 FILLER_15_2590 ();
 sg13g2_decap_8 FILLER_15_2597 ();
 sg13g2_decap_8 FILLER_15_2604 ();
 sg13g2_decap_8 FILLER_15_2611 ();
 sg13g2_decap_8 FILLER_15_2618 ();
 sg13g2_decap_8 FILLER_15_2625 ();
 sg13g2_decap_8 FILLER_15_2632 ();
 sg13g2_decap_8 FILLER_15_2639 ();
 sg13g2_decap_8 FILLER_15_2646 ();
 sg13g2_decap_8 FILLER_15_2653 ();
 sg13g2_decap_8 FILLER_15_2660 ();
 sg13g2_decap_8 FILLER_15_2667 ();
 sg13g2_decap_8 FILLER_15_2674 ();
 sg13g2_decap_8 FILLER_15_2681 ();
 sg13g2_decap_8 FILLER_15_2688 ();
 sg13g2_decap_8 FILLER_15_2695 ();
 sg13g2_decap_8 FILLER_15_2702 ();
 sg13g2_decap_8 FILLER_15_2709 ();
 sg13g2_decap_8 FILLER_15_2716 ();
 sg13g2_decap_8 FILLER_15_2723 ();
 sg13g2_decap_8 FILLER_15_2730 ();
 sg13g2_decap_8 FILLER_15_2737 ();
 sg13g2_decap_8 FILLER_15_2744 ();
 sg13g2_decap_8 FILLER_15_2751 ();
 sg13g2_decap_8 FILLER_15_2758 ();
 sg13g2_decap_8 FILLER_15_2765 ();
 sg13g2_decap_8 FILLER_15_2772 ();
 sg13g2_decap_8 FILLER_15_2779 ();
 sg13g2_decap_8 FILLER_15_2786 ();
 sg13g2_decap_8 FILLER_15_2793 ();
 sg13g2_decap_8 FILLER_15_2800 ();
 sg13g2_decap_8 FILLER_15_2807 ();
 sg13g2_decap_8 FILLER_15_2814 ();
 sg13g2_decap_8 FILLER_15_2821 ();
 sg13g2_decap_8 FILLER_15_2828 ();
 sg13g2_decap_8 FILLER_15_2835 ();
 sg13g2_decap_8 FILLER_15_2842 ();
 sg13g2_decap_8 FILLER_15_2849 ();
 sg13g2_decap_8 FILLER_15_2856 ();
 sg13g2_decap_8 FILLER_15_2863 ();
 sg13g2_decap_8 FILLER_15_2870 ();
 sg13g2_decap_8 FILLER_15_2877 ();
 sg13g2_decap_8 FILLER_15_2884 ();
 sg13g2_decap_8 FILLER_15_2891 ();
 sg13g2_decap_8 FILLER_15_2898 ();
 sg13g2_decap_8 FILLER_15_2905 ();
 sg13g2_decap_8 FILLER_15_2912 ();
 sg13g2_decap_8 FILLER_15_2919 ();
 sg13g2_decap_8 FILLER_15_2926 ();
 sg13g2_decap_8 FILLER_15_2933 ();
 sg13g2_decap_8 FILLER_15_2940 ();
 sg13g2_decap_8 FILLER_15_2947 ();
 sg13g2_decap_8 FILLER_15_2954 ();
 sg13g2_decap_8 FILLER_15_2961 ();
 sg13g2_decap_8 FILLER_15_2968 ();
 sg13g2_decap_8 FILLER_15_2975 ();
 sg13g2_decap_8 FILLER_15_2982 ();
 sg13g2_decap_8 FILLER_15_2989 ();
 sg13g2_decap_8 FILLER_15_2996 ();
 sg13g2_decap_8 FILLER_15_3003 ();
 sg13g2_decap_8 FILLER_15_3010 ();
 sg13g2_decap_8 FILLER_15_3017 ();
 sg13g2_decap_8 FILLER_15_3024 ();
 sg13g2_decap_8 FILLER_15_3031 ();
 sg13g2_decap_8 FILLER_15_3038 ();
 sg13g2_decap_8 FILLER_15_3045 ();
 sg13g2_decap_8 FILLER_15_3052 ();
 sg13g2_decap_8 FILLER_15_3059 ();
 sg13g2_decap_8 FILLER_15_3066 ();
 sg13g2_decap_8 FILLER_15_3073 ();
 sg13g2_decap_8 FILLER_15_3080 ();
 sg13g2_decap_8 FILLER_15_3087 ();
 sg13g2_decap_8 FILLER_15_3094 ();
 sg13g2_decap_8 FILLER_15_3101 ();
 sg13g2_decap_8 FILLER_15_3108 ();
 sg13g2_decap_8 FILLER_15_3115 ();
 sg13g2_decap_8 FILLER_15_3122 ();
 sg13g2_decap_8 FILLER_15_3129 ();
 sg13g2_decap_8 FILLER_15_3136 ();
 sg13g2_decap_8 FILLER_15_3143 ();
 sg13g2_decap_8 FILLER_15_3150 ();
 sg13g2_decap_8 FILLER_15_3157 ();
 sg13g2_decap_8 FILLER_15_3164 ();
 sg13g2_decap_8 FILLER_15_3171 ();
 sg13g2_decap_8 FILLER_15_3178 ();
 sg13g2_decap_8 FILLER_15_3185 ();
 sg13g2_decap_8 FILLER_15_3192 ();
 sg13g2_decap_8 FILLER_15_3199 ();
 sg13g2_decap_8 FILLER_15_3206 ();
 sg13g2_decap_8 FILLER_15_3213 ();
 sg13g2_decap_8 FILLER_15_3220 ();
 sg13g2_decap_8 FILLER_15_3227 ();
 sg13g2_decap_8 FILLER_15_3234 ();
 sg13g2_decap_8 FILLER_15_3241 ();
 sg13g2_decap_8 FILLER_15_3248 ();
 sg13g2_decap_8 FILLER_15_3255 ();
 sg13g2_decap_8 FILLER_15_3262 ();
 sg13g2_decap_8 FILLER_15_3269 ();
 sg13g2_decap_8 FILLER_15_3276 ();
 sg13g2_decap_8 FILLER_15_3283 ();
 sg13g2_decap_8 FILLER_15_3290 ();
 sg13g2_decap_8 FILLER_15_3297 ();
 sg13g2_decap_8 FILLER_15_3304 ();
 sg13g2_decap_8 FILLER_15_3311 ();
 sg13g2_decap_8 FILLER_15_3318 ();
 sg13g2_decap_8 FILLER_15_3325 ();
 sg13g2_decap_8 FILLER_15_3332 ();
 sg13g2_decap_8 FILLER_15_3339 ();
 sg13g2_decap_8 FILLER_15_3346 ();
 sg13g2_decap_8 FILLER_15_3353 ();
 sg13g2_decap_8 FILLER_15_3360 ();
 sg13g2_decap_8 FILLER_15_3367 ();
 sg13g2_decap_8 FILLER_15_3374 ();
 sg13g2_decap_8 FILLER_15_3381 ();
 sg13g2_decap_8 FILLER_15_3388 ();
 sg13g2_decap_8 FILLER_15_3395 ();
 sg13g2_decap_8 FILLER_15_3402 ();
 sg13g2_decap_8 FILLER_15_3409 ();
 sg13g2_decap_8 FILLER_15_3416 ();
 sg13g2_decap_8 FILLER_15_3423 ();
 sg13g2_decap_8 FILLER_15_3430 ();
 sg13g2_decap_8 FILLER_15_3437 ();
 sg13g2_decap_8 FILLER_15_3444 ();
 sg13g2_decap_8 FILLER_15_3451 ();
 sg13g2_decap_8 FILLER_15_3458 ();
 sg13g2_decap_8 FILLER_15_3465 ();
 sg13g2_decap_8 FILLER_15_3472 ();
 sg13g2_decap_8 FILLER_15_3479 ();
 sg13g2_decap_8 FILLER_15_3486 ();
 sg13g2_decap_8 FILLER_15_3493 ();
 sg13g2_decap_8 FILLER_15_3500 ();
 sg13g2_decap_8 FILLER_15_3507 ();
 sg13g2_decap_8 FILLER_15_3514 ();
 sg13g2_decap_8 FILLER_15_3521 ();
 sg13g2_decap_8 FILLER_15_3528 ();
 sg13g2_decap_8 FILLER_15_3535 ();
 sg13g2_decap_8 FILLER_15_3542 ();
 sg13g2_decap_8 FILLER_15_3549 ();
 sg13g2_decap_8 FILLER_15_3556 ();
 sg13g2_decap_8 FILLER_15_3563 ();
 sg13g2_decap_8 FILLER_15_3570 ();
 sg13g2_fill_2 FILLER_15_3577 ();
 sg13g2_fill_1 FILLER_15_3579 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_decap_8 FILLER_16_427 ();
 sg13g2_decap_8 FILLER_16_434 ();
 sg13g2_decap_8 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_448 ();
 sg13g2_decap_8 FILLER_16_455 ();
 sg13g2_decap_8 FILLER_16_462 ();
 sg13g2_decap_8 FILLER_16_469 ();
 sg13g2_decap_8 FILLER_16_476 ();
 sg13g2_decap_8 FILLER_16_483 ();
 sg13g2_decap_8 FILLER_16_490 ();
 sg13g2_decap_8 FILLER_16_497 ();
 sg13g2_decap_8 FILLER_16_504 ();
 sg13g2_decap_8 FILLER_16_511 ();
 sg13g2_decap_8 FILLER_16_518 ();
 sg13g2_decap_8 FILLER_16_525 ();
 sg13g2_decap_8 FILLER_16_532 ();
 sg13g2_decap_8 FILLER_16_539 ();
 sg13g2_decap_8 FILLER_16_546 ();
 sg13g2_decap_8 FILLER_16_553 ();
 sg13g2_decap_8 FILLER_16_560 ();
 sg13g2_decap_8 FILLER_16_567 ();
 sg13g2_decap_8 FILLER_16_574 ();
 sg13g2_decap_8 FILLER_16_581 ();
 sg13g2_decap_8 FILLER_16_588 ();
 sg13g2_decap_8 FILLER_16_595 ();
 sg13g2_decap_8 FILLER_16_602 ();
 sg13g2_decap_8 FILLER_16_609 ();
 sg13g2_decap_8 FILLER_16_616 ();
 sg13g2_decap_8 FILLER_16_623 ();
 sg13g2_decap_8 FILLER_16_630 ();
 sg13g2_decap_8 FILLER_16_637 ();
 sg13g2_decap_8 FILLER_16_644 ();
 sg13g2_decap_8 FILLER_16_651 ();
 sg13g2_decap_8 FILLER_16_658 ();
 sg13g2_decap_8 FILLER_16_665 ();
 sg13g2_decap_8 FILLER_16_672 ();
 sg13g2_decap_8 FILLER_16_679 ();
 sg13g2_decap_8 FILLER_16_686 ();
 sg13g2_decap_8 FILLER_16_693 ();
 sg13g2_decap_8 FILLER_16_700 ();
 sg13g2_decap_8 FILLER_16_707 ();
 sg13g2_decap_8 FILLER_16_714 ();
 sg13g2_decap_8 FILLER_16_721 ();
 sg13g2_decap_8 FILLER_16_728 ();
 sg13g2_decap_8 FILLER_16_735 ();
 sg13g2_decap_8 FILLER_16_742 ();
 sg13g2_decap_8 FILLER_16_749 ();
 sg13g2_decap_8 FILLER_16_756 ();
 sg13g2_decap_8 FILLER_16_763 ();
 sg13g2_decap_8 FILLER_16_770 ();
 sg13g2_decap_8 FILLER_16_777 ();
 sg13g2_decap_8 FILLER_16_784 ();
 sg13g2_decap_8 FILLER_16_791 ();
 sg13g2_decap_8 FILLER_16_798 ();
 sg13g2_decap_8 FILLER_16_805 ();
 sg13g2_decap_8 FILLER_16_812 ();
 sg13g2_decap_8 FILLER_16_819 ();
 sg13g2_decap_8 FILLER_16_826 ();
 sg13g2_decap_8 FILLER_16_833 ();
 sg13g2_decap_8 FILLER_16_840 ();
 sg13g2_decap_8 FILLER_16_847 ();
 sg13g2_decap_8 FILLER_16_854 ();
 sg13g2_decap_8 FILLER_16_861 ();
 sg13g2_decap_8 FILLER_16_868 ();
 sg13g2_decap_8 FILLER_16_875 ();
 sg13g2_decap_8 FILLER_16_882 ();
 sg13g2_decap_8 FILLER_16_889 ();
 sg13g2_decap_8 FILLER_16_896 ();
 sg13g2_decap_8 FILLER_16_903 ();
 sg13g2_decap_8 FILLER_16_910 ();
 sg13g2_decap_8 FILLER_16_917 ();
 sg13g2_decap_8 FILLER_16_924 ();
 sg13g2_decap_8 FILLER_16_931 ();
 sg13g2_decap_8 FILLER_16_938 ();
 sg13g2_decap_8 FILLER_16_945 ();
 sg13g2_decap_8 FILLER_16_952 ();
 sg13g2_decap_8 FILLER_16_959 ();
 sg13g2_decap_8 FILLER_16_966 ();
 sg13g2_decap_8 FILLER_16_973 ();
 sg13g2_decap_8 FILLER_16_980 ();
 sg13g2_decap_8 FILLER_16_987 ();
 sg13g2_decap_8 FILLER_16_994 ();
 sg13g2_decap_8 FILLER_16_1001 ();
 sg13g2_decap_8 FILLER_16_1008 ();
 sg13g2_decap_8 FILLER_16_1015 ();
 sg13g2_decap_8 FILLER_16_1022 ();
 sg13g2_decap_8 FILLER_16_1029 ();
 sg13g2_decap_8 FILLER_16_1036 ();
 sg13g2_decap_8 FILLER_16_1043 ();
 sg13g2_decap_8 FILLER_16_1050 ();
 sg13g2_decap_8 FILLER_16_1057 ();
 sg13g2_decap_8 FILLER_16_1064 ();
 sg13g2_decap_8 FILLER_16_1071 ();
 sg13g2_decap_8 FILLER_16_1078 ();
 sg13g2_decap_8 FILLER_16_1085 ();
 sg13g2_decap_8 FILLER_16_1092 ();
 sg13g2_decap_8 FILLER_16_1099 ();
 sg13g2_decap_8 FILLER_16_1106 ();
 sg13g2_decap_8 FILLER_16_1113 ();
 sg13g2_decap_8 FILLER_16_1120 ();
 sg13g2_decap_8 FILLER_16_1127 ();
 sg13g2_decap_8 FILLER_16_1134 ();
 sg13g2_decap_8 FILLER_16_1141 ();
 sg13g2_decap_8 FILLER_16_1148 ();
 sg13g2_decap_8 FILLER_16_1155 ();
 sg13g2_decap_8 FILLER_16_1162 ();
 sg13g2_decap_8 FILLER_16_1169 ();
 sg13g2_decap_8 FILLER_16_1176 ();
 sg13g2_decap_8 FILLER_16_1183 ();
 sg13g2_decap_8 FILLER_16_1190 ();
 sg13g2_decap_8 FILLER_16_1197 ();
 sg13g2_decap_8 FILLER_16_1204 ();
 sg13g2_decap_8 FILLER_16_1211 ();
 sg13g2_decap_8 FILLER_16_1218 ();
 sg13g2_decap_8 FILLER_16_1225 ();
 sg13g2_decap_8 FILLER_16_1232 ();
 sg13g2_decap_8 FILLER_16_1239 ();
 sg13g2_decap_8 FILLER_16_1246 ();
 sg13g2_decap_8 FILLER_16_1253 ();
 sg13g2_decap_8 FILLER_16_1260 ();
 sg13g2_decap_8 FILLER_16_1267 ();
 sg13g2_decap_8 FILLER_16_1274 ();
 sg13g2_decap_8 FILLER_16_1281 ();
 sg13g2_decap_8 FILLER_16_1288 ();
 sg13g2_decap_8 FILLER_16_1295 ();
 sg13g2_decap_8 FILLER_16_1302 ();
 sg13g2_decap_8 FILLER_16_1309 ();
 sg13g2_decap_8 FILLER_16_1316 ();
 sg13g2_decap_8 FILLER_16_1323 ();
 sg13g2_decap_8 FILLER_16_1330 ();
 sg13g2_decap_8 FILLER_16_1337 ();
 sg13g2_decap_8 FILLER_16_1344 ();
 sg13g2_decap_8 FILLER_16_1351 ();
 sg13g2_decap_8 FILLER_16_1358 ();
 sg13g2_decap_8 FILLER_16_1365 ();
 sg13g2_decap_8 FILLER_16_1372 ();
 sg13g2_decap_8 FILLER_16_1379 ();
 sg13g2_decap_8 FILLER_16_1386 ();
 sg13g2_decap_8 FILLER_16_1393 ();
 sg13g2_decap_8 FILLER_16_1400 ();
 sg13g2_decap_8 FILLER_16_1407 ();
 sg13g2_decap_8 FILLER_16_1414 ();
 sg13g2_decap_8 FILLER_16_1421 ();
 sg13g2_decap_8 FILLER_16_1428 ();
 sg13g2_decap_8 FILLER_16_1435 ();
 sg13g2_decap_8 FILLER_16_1442 ();
 sg13g2_decap_8 FILLER_16_1449 ();
 sg13g2_decap_8 FILLER_16_1456 ();
 sg13g2_decap_8 FILLER_16_1463 ();
 sg13g2_decap_8 FILLER_16_1470 ();
 sg13g2_decap_8 FILLER_16_1477 ();
 sg13g2_decap_8 FILLER_16_1484 ();
 sg13g2_decap_8 FILLER_16_1491 ();
 sg13g2_decap_8 FILLER_16_1498 ();
 sg13g2_decap_8 FILLER_16_1505 ();
 sg13g2_decap_8 FILLER_16_1512 ();
 sg13g2_decap_8 FILLER_16_1519 ();
 sg13g2_decap_8 FILLER_16_1526 ();
 sg13g2_decap_8 FILLER_16_1533 ();
 sg13g2_decap_8 FILLER_16_1540 ();
 sg13g2_decap_8 FILLER_16_1547 ();
 sg13g2_decap_8 FILLER_16_1554 ();
 sg13g2_decap_8 FILLER_16_1561 ();
 sg13g2_decap_8 FILLER_16_1568 ();
 sg13g2_decap_8 FILLER_16_1575 ();
 sg13g2_decap_8 FILLER_16_1582 ();
 sg13g2_decap_8 FILLER_16_1589 ();
 sg13g2_decap_8 FILLER_16_1596 ();
 sg13g2_decap_8 FILLER_16_1603 ();
 sg13g2_decap_8 FILLER_16_1610 ();
 sg13g2_decap_8 FILLER_16_1617 ();
 sg13g2_decap_8 FILLER_16_1624 ();
 sg13g2_decap_8 FILLER_16_1631 ();
 sg13g2_decap_8 FILLER_16_1638 ();
 sg13g2_decap_8 FILLER_16_1645 ();
 sg13g2_decap_8 FILLER_16_1652 ();
 sg13g2_decap_8 FILLER_16_1659 ();
 sg13g2_decap_8 FILLER_16_1666 ();
 sg13g2_decap_8 FILLER_16_1673 ();
 sg13g2_decap_8 FILLER_16_1680 ();
 sg13g2_decap_8 FILLER_16_1687 ();
 sg13g2_decap_8 FILLER_16_1694 ();
 sg13g2_decap_8 FILLER_16_1701 ();
 sg13g2_decap_8 FILLER_16_1708 ();
 sg13g2_decap_8 FILLER_16_1715 ();
 sg13g2_decap_8 FILLER_16_1722 ();
 sg13g2_decap_8 FILLER_16_1729 ();
 sg13g2_decap_8 FILLER_16_1736 ();
 sg13g2_decap_8 FILLER_16_1743 ();
 sg13g2_decap_8 FILLER_16_1750 ();
 sg13g2_decap_8 FILLER_16_1757 ();
 sg13g2_decap_8 FILLER_16_1764 ();
 sg13g2_decap_8 FILLER_16_1771 ();
 sg13g2_decap_8 FILLER_16_1778 ();
 sg13g2_decap_8 FILLER_16_1785 ();
 sg13g2_decap_8 FILLER_16_1792 ();
 sg13g2_decap_8 FILLER_16_1799 ();
 sg13g2_decap_8 FILLER_16_1806 ();
 sg13g2_decap_8 FILLER_16_1813 ();
 sg13g2_decap_8 FILLER_16_1820 ();
 sg13g2_decap_8 FILLER_16_1827 ();
 sg13g2_decap_8 FILLER_16_1834 ();
 sg13g2_decap_8 FILLER_16_1841 ();
 sg13g2_decap_8 FILLER_16_1848 ();
 sg13g2_decap_8 FILLER_16_1855 ();
 sg13g2_decap_8 FILLER_16_1862 ();
 sg13g2_decap_8 FILLER_16_1869 ();
 sg13g2_decap_8 FILLER_16_1876 ();
 sg13g2_decap_8 FILLER_16_1883 ();
 sg13g2_decap_8 FILLER_16_1890 ();
 sg13g2_decap_8 FILLER_16_1897 ();
 sg13g2_decap_8 FILLER_16_1904 ();
 sg13g2_decap_8 FILLER_16_1911 ();
 sg13g2_decap_8 FILLER_16_1918 ();
 sg13g2_decap_8 FILLER_16_1925 ();
 sg13g2_decap_8 FILLER_16_1932 ();
 sg13g2_decap_8 FILLER_16_1939 ();
 sg13g2_decap_8 FILLER_16_1946 ();
 sg13g2_decap_8 FILLER_16_1953 ();
 sg13g2_decap_8 FILLER_16_1960 ();
 sg13g2_decap_8 FILLER_16_1967 ();
 sg13g2_decap_8 FILLER_16_1974 ();
 sg13g2_decap_8 FILLER_16_1981 ();
 sg13g2_decap_8 FILLER_16_1988 ();
 sg13g2_decap_8 FILLER_16_1995 ();
 sg13g2_decap_8 FILLER_16_2002 ();
 sg13g2_decap_8 FILLER_16_2009 ();
 sg13g2_decap_8 FILLER_16_2016 ();
 sg13g2_decap_8 FILLER_16_2023 ();
 sg13g2_decap_8 FILLER_16_2030 ();
 sg13g2_decap_8 FILLER_16_2037 ();
 sg13g2_decap_8 FILLER_16_2044 ();
 sg13g2_decap_8 FILLER_16_2051 ();
 sg13g2_decap_8 FILLER_16_2058 ();
 sg13g2_decap_8 FILLER_16_2065 ();
 sg13g2_decap_8 FILLER_16_2072 ();
 sg13g2_decap_8 FILLER_16_2079 ();
 sg13g2_decap_8 FILLER_16_2086 ();
 sg13g2_decap_8 FILLER_16_2093 ();
 sg13g2_decap_8 FILLER_16_2100 ();
 sg13g2_decap_8 FILLER_16_2107 ();
 sg13g2_decap_8 FILLER_16_2114 ();
 sg13g2_decap_8 FILLER_16_2121 ();
 sg13g2_decap_8 FILLER_16_2128 ();
 sg13g2_decap_8 FILLER_16_2135 ();
 sg13g2_decap_8 FILLER_16_2142 ();
 sg13g2_decap_8 FILLER_16_2149 ();
 sg13g2_decap_8 FILLER_16_2156 ();
 sg13g2_decap_8 FILLER_16_2163 ();
 sg13g2_decap_8 FILLER_16_2170 ();
 sg13g2_decap_8 FILLER_16_2177 ();
 sg13g2_decap_8 FILLER_16_2184 ();
 sg13g2_decap_8 FILLER_16_2191 ();
 sg13g2_decap_8 FILLER_16_2198 ();
 sg13g2_decap_8 FILLER_16_2205 ();
 sg13g2_decap_8 FILLER_16_2212 ();
 sg13g2_decap_8 FILLER_16_2219 ();
 sg13g2_decap_8 FILLER_16_2226 ();
 sg13g2_decap_8 FILLER_16_2233 ();
 sg13g2_decap_8 FILLER_16_2240 ();
 sg13g2_decap_8 FILLER_16_2247 ();
 sg13g2_decap_8 FILLER_16_2254 ();
 sg13g2_decap_8 FILLER_16_2261 ();
 sg13g2_decap_8 FILLER_16_2268 ();
 sg13g2_decap_8 FILLER_16_2275 ();
 sg13g2_decap_8 FILLER_16_2282 ();
 sg13g2_decap_8 FILLER_16_2289 ();
 sg13g2_decap_8 FILLER_16_2296 ();
 sg13g2_decap_8 FILLER_16_2303 ();
 sg13g2_decap_8 FILLER_16_2310 ();
 sg13g2_decap_8 FILLER_16_2317 ();
 sg13g2_decap_8 FILLER_16_2324 ();
 sg13g2_decap_8 FILLER_16_2331 ();
 sg13g2_decap_8 FILLER_16_2338 ();
 sg13g2_decap_8 FILLER_16_2345 ();
 sg13g2_decap_8 FILLER_16_2352 ();
 sg13g2_decap_8 FILLER_16_2359 ();
 sg13g2_decap_8 FILLER_16_2366 ();
 sg13g2_decap_8 FILLER_16_2373 ();
 sg13g2_decap_8 FILLER_16_2380 ();
 sg13g2_decap_8 FILLER_16_2387 ();
 sg13g2_decap_8 FILLER_16_2394 ();
 sg13g2_decap_8 FILLER_16_2401 ();
 sg13g2_decap_8 FILLER_16_2408 ();
 sg13g2_decap_8 FILLER_16_2415 ();
 sg13g2_decap_8 FILLER_16_2422 ();
 sg13g2_decap_8 FILLER_16_2429 ();
 sg13g2_decap_8 FILLER_16_2436 ();
 sg13g2_decap_8 FILLER_16_2443 ();
 sg13g2_decap_8 FILLER_16_2450 ();
 sg13g2_decap_8 FILLER_16_2457 ();
 sg13g2_decap_8 FILLER_16_2464 ();
 sg13g2_decap_8 FILLER_16_2471 ();
 sg13g2_decap_8 FILLER_16_2478 ();
 sg13g2_decap_8 FILLER_16_2485 ();
 sg13g2_decap_8 FILLER_16_2492 ();
 sg13g2_decap_8 FILLER_16_2499 ();
 sg13g2_decap_8 FILLER_16_2506 ();
 sg13g2_decap_8 FILLER_16_2513 ();
 sg13g2_decap_8 FILLER_16_2520 ();
 sg13g2_decap_8 FILLER_16_2527 ();
 sg13g2_decap_8 FILLER_16_2534 ();
 sg13g2_decap_8 FILLER_16_2541 ();
 sg13g2_decap_8 FILLER_16_2548 ();
 sg13g2_decap_8 FILLER_16_2555 ();
 sg13g2_decap_8 FILLER_16_2562 ();
 sg13g2_decap_8 FILLER_16_2569 ();
 sg13g2_decap_8 FILLER_16_2576 ();
 sg13g2_decap_8 FILLER_16_2583 ();
 sg13g2_decap_8 FILLER_16_2590 ();
 sg13g2_decap_8 FILLER_16_2597 ();
 sg13g2_decap_8 FILLER_16_2604 ();
 sg13g2_decap_8 FILLER_16_2611 ();
 sg13g2_decap_8 FILLER_16_2618 ();
 sg13g2_decap_8 FILLER_16_2625 ();
 sg13g2_decap_8 FILLER_16_2632 ();
 sg13g2_decap_8 FILLER_16_2639 ();
 sg13g2_decap_8 FILLER_16_2646 ();
 sg13g2_decap_8 FILLER_16_2653 ();
 sg13g2_decap_8 FILLER_16_2660 ();
 sg13g2_decap_8 FILLER_16_2667 ();
 sg13g2_decap_8 FILLER_16_2674 ();
 sg13g2_decap_8 FILLER_16_2681 ();
 sg13g2_decap_8 FILLER_16_2688 ();
 sg13g2_decap_8 FILLER_16_2695 ();
 sg13g2_decap_8 FILLER_16_2702 ();
 sg13g2_decap_8 FILLER_16_2709 ();
 sg13g2_decap_8 FILLER_16_2716 ();
 sg13g2_decap_8 FILLER_16_2723 ();
 sg13g2_decap_8 FILLER_16_2730 ();
 sg13g2_decap_8 FILLER_16_2737 ();
 sg13g2_decap_8 FILLER_16_2744 ();
 sg13g2_decap_8 FILLER_16_2751 ();
 sg13g2_decap_8 FILLER_16_2758 ();
 sg13g2_decap_8 FILLER_16_2765 ();
 sg13g2_decap_8 FILLER_16_2772 ();
 sg13g2_decap_8 FILLER_16_2779 ();
 sg13g2_decap_8 FILLER_16_2786 ();
 sg13g2_decap_8 FILLER_16_2793 ();
 sg13g2_decap_8 FILLER_16_2800 ();
 sg13g2_decap_8 FILLER_16_2807 ();
 sg13g2_decap_8 FILLER_16_2814 ();
 sg13g2_decap_8 FILLER_16_2821 ();
 sg13g2_decap_8 FILLER_16_2828 ();
 sg13g2_decap_8 FILLER_16_2835 ();
 sg13g2_decap_8 FILLER_16_2842 ();
 sg13g2_decap_8 FILLER_16_2849 ();
 sg13g2_decap_8 FILLER_16_2856 ();
 sg13g2_decap_8 FILLER_16_2863 ();
 sg13g2_decap_8 FILLER_16_2870 ();
 sg13g2_decap_8 FILLER_16_2877 ();
 sg13g2_decap_8 FILLER_16_2884 ();
 sg13g2_decap_8 FILLER_16_2891 ();
 sg13g2_decap_8 FILLER_16_2898 ();
 sg13g2_decap_8 FILLER_16_2905 ();
 sg13g2_decap_8 FILLER_16_2912 ();
 sg13g2_decap_8 FILLER_16_2919 ();
 sg13g2_decap_8 FILLER_16_2926 ();
 sg13g2_decap_8 FILLER_16_2933 ();
 sg13g2_decap_8 FILLER_16_2940 ();
 sg13g2_decap_8 FILLER_16_2947 ();
 sg13g2_decap_8 FILLER_16_2954 ();
 sg13g2_decap_8 FILLER_16_2961 ();
 sg13g2_decap_8 FILLER_16_2968 ();
 sg13g2_decap_8 FILLER_16_2975 ();
 sg13g2_decap_8 FILLER_16_2982 ();
 sg13g2_decap_8 FILLER_16_2989 ();
 sg13g2_decap_8 FILLER_16_2996 ();
 sg13g2_decap_8 FILLER_16_3003 ();
 sg13g2_decap_8 FILLER_16_3010 ();
 sg13g2_decap_8 FILLER_16_3017 ();
 sg13g2_decap_8 FILLER_16_3024 ();
 sg13g2_decap_8 FILLER_16_3031 ();
 sg13g2_decap_8 FILLER_16_3038 ();
 sg13g2_decap_8 FILLER_16_3045 ();
 sg13g2_decap_8 FILLER_16_3052 ();
 sg13g2_decap_8 FILLER_16_3059 ();
 sg13g2_decap_8 FILLER_16_3066 ();
 sg13g2_decap_8 FILLER_16_3073 ();
 sg13g2_decap_8 FILLER_16_3080 ();
 sg13g2_decap_8 FILLER_16_3087 ();
 sg13g2_decap_8 FILLER_16_3094 ();
 sg13g2_decap_8 FILLER_16_3101 ();
 sg13g2_decap_8 FILLER_16_3108 ();
 sg13g2_decap_8 FILLER_16_3115 ();
 sg13g2_decap_8 FILLER_16_3122 ();
 sg13g2_decap_8 FILLER_16_3129 ();
 sg13g2_decap_8 FILLER_16_3136 ();
 sg13g2_decap_8 FILLER_16_3143 ();
 sg13g2_decap_8 FILLER_16_3150 ();
 sg13g2_decap_8 FILLER_16_3157 ();
 sg13g2_decap_8 FILLER_16_3164 ();
 sg13g2_decap_8 FILLER_16_3171 ();
 sg13g2_decap_8 FILLER_16_3178 ();
 sg13g2_decap_8 FILLER_16_3185 ();
 sg13g2_decap_8 FILLER_16_3192 ();
 sg13g2_decap_8 FILLER_16_3199 ();
 sg13g2_decap_8 FILLER_16_3206 ();
 sg13g2_decap_8 FILLER_16_3213 ();
 sg13g2_decap_8 FILLER_16_3220 ();
 sg13g2_decap_8 FILLER_16_3227 ();
 sg13g2_decap_8 FILLER_16_3234 ();
 sg13g2_decap_8 FILLER_16_3241 ();
 sg13g2_decap_8 FILLER_16_3248 ();
 sg13g2_decap_8 FILLER_16_3255 ();
 sg13g2_decap_8 FILLER_16_3262 ();
 sg13g2_decap_8 FILLER_16_3269 ();
 sg13g2_decap_8 FILLER_16_3276 ();
 sg13g2_decap_8 FILLER_16_3283 ();
 sg13g2_decap_8 FILLER_16_3290 ();
 sg13g2_decap_8 FILLER_16_3297 ();
 sg13g2_decap_8 FILLER_16_3304 ();
 sg13g2_decap_8 FILLER_16_3311 ();
 sg13g2_decap_8 FILLER_16_3318 ();
 sg13g2_decap_8 FILLER_16_3325 ();
 sg13g2_decap_8 FILLER_16_3332 ();
 sg13g2_decap_8 FILLER_16_3339 ();
 sg13g2_decap_8 FILLER_16_3346 ();
 sg13g2_decap_8 FILLER_16_3353 ();
 sg13g2_decap_8 FILLER_16_3360 ();
 sg13g2_decap_8 FILLER_16_3367 ();
 sg13g2_decap_8 FILLER_16_3374 ();
 sg13g2_decap_8 FILLER_16_3381 ();
 sg13g2_decap_8 FILLER_16_3388 ();
 sg13g2_decap_8 FILLER_16_3395 ();
 sg13g2_decap_8 FILLER_16_3402 ();
 sg13g2_decap_8 FILLER_16_3409 ();
 sg13g2_decap_8 FILLER_16_3416 ();
 sg13g2_decap_8 FILLER_16_3423 ();
 sg13g2_decap_8 FILLER_16_3430 ();
 sg13g2_decap_8 FILLER_16_3437 ();
 sg13g2_decap_8 FILLER_16_3444 ();
 sg13g2_decap_8 FILLER_16_3451 ();
 sg13g2_decap_8 FILLER_16_3458 ();
 sg13g2_decap_8 FILLER_16_3465 ();
 sg13g2_decap_8 FILLER_16_3472 ();
 sg13g2_decap_8 FILLER_16_3479 ();
 sg13g2_decap_8 FILLER_16_3486 ();
 sg13g2_decap_8 FILLER_16_3493 ();
 sg13g2_decap_8 FILLER_16_3500 ();
 sg13g2_decap_8 FILLER_16_3507 ();
 sg13g2_decap_8 FILLER_16_3514 ();
 sg13g2_decap_8 FILLER_16_3521 ();
 sg13g2_decap_8 FILLER_16_3528 ();
 sg13g2_decap_8 FILLER_16_3535 ();
 sg13g2_decap_8 FILLER_16_3542 ();
 sg13g2_decap_8 FILLER_16_3549 ();
 sg13g2_decap_8 FILLER_16_3556 ();
 sg13g2_decap_8 FILLER_16_3563 ();
 sg13g2_decap_8 FILLER_16_3570 ();
 sg13g2_fill_2 FILLER_16_3577 ();
 sg13g2_fill_1 FILLER_16_3579 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_8 FILLER_17_427 ();
 sg13g2_decap_8 FILLER_17_434 ();
 sg13g2_decap_8 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_448 ();
 sg13g2_decap_8 FILLER_17_455 ();
 sg13g2_decap_8 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_decap_8 FILLER_17_483 ();
 sg13g2_decap_8 FILLER_17_490 ();
 sg13g2_decap_8 FILLER_17_497 ();
 sg13g2_decap_8 FILLER_17_504 ();
 sg13g2_decap_8 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_518 ();
 sg13g2_decap_8 FILLER_17_525 ();
 sg13g2_decap_8 FILLER_17_532 ();
 sg13g2_decap_8 FILLER_17_539 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_decap_8 FILLER_17_567 ();
 sg13g2_decap_8 FILLER_17_574 ();
 sg13g2_decap_8 FILLER_17_581 ();
 sg13g2_decap_8 FILLER_17_588 ();
 sg13g2_decap_8 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_decap_8 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_644 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_679 ();
 sg13g2_decap_8 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_693 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_8 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_8 FILLER_17_854 ();
 sg13g2_decap_8 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_17_868 ();
 sg13g2_decap_8 FILLER_17_875 ();
 sg13g2_decap_8 FILLER_17_882 ();
 sg13g2_decap_8 FILLER_17_889 ();
 sg13g2_decap_8 FILLER_17_896 ();
 sg13g2_decap_8 FILLER_17_903 ();
 sg13g2_decap_8 FILLER_17_910 ();
 sg13g2_decap_8 FILLER_17_917 ();
 sg13g2_decap_8 FILLER_17_924 ();
 sg13g2_decap_8 FILLER_17_931 ();
 sg13g2_decap_8 FILLER_17_938 ();
 sg13g2_decap_8 FILLER_17_945 ();
 sg13g2_decap_8 FILLER_17_952 ();
 sg13g2_decap_8 FILLER_17_959 ();
 sg13g2_decap_8 FILLER_17_966 ();
 sg13g2_decap_8 FILLER_17_973 ();
 sg13g2_decap_8 FILLER_17_980 ();
 sg13g2_decap_8 FILLER_17_987 ();
 sg13g2_decap_8 FILLER_17_994 ();
 sg13g2_decap_8 FILLER_17_1001 ();
 sg13g2_decap_8 FILLER_17_1008 ();
 sg13g2_decap_8 FILLER_17_1015 ();
 sg13g2_decap_8 FILLER_17_1022 ();
 sg13g2_decap_8 FILLER_17_1029 ();
 sg13g2_decap_8 FILLER_17_1036 ();
 sg13g2_decap_8 FILLER_17_1043 ();
 sg13g2_decap_8 FILLER_17_1050 ();
 sg13g2_decap_8 FILLER_17_1057 ();
 sg13g2_decap_8 FILLER_17_1064 ();
 sg13g2_decap_8 FILLER_17_1071 ();
 sg13g2_decap_8 FILLER_17_1078 ();
 sg13g2_decap_8 FILLER_17_1085 ();
 sg13g2_decap_8 FILLER_17_1092 ();
 sg13g2_decap_8 FILLER_17_1099 ();
 sg13g2_decap_8 FILLER_17_1106 ();
 sg13g2_decap_8 FILLER_17_1113 ();
 sg13g2_decap_8 FILLER_17_1120 ();
 sg13g2_decap_8 FILLER_17_1127 ();
 sg13g2_decap_8 FILLER_17_1134 ();
 sg13g2_decap_8 FILLER_17_1141 ();
 sg13g2_decap_8 FILLER_17_1148 ();
 sg13g2_decap_8 FILLER_17_1155 ();
 sg13g2_decap_8 FILLER_17_1162 ();
 sg13g2_decap_8 FILLER_17_1169 ();
 sg13g2_decap_8 FILLER_17_1176 ();
 sg13g2_decap_8 FILLER_17_1183 ();
 sg13g2_decap_8 FILLER_17_1190 ();
 sg13g2_decap_8 FILLER_17_1197 ();
 sg13g2_decap_8 FILLER_17_1204 ();
 sg13g2_decap_8 FILLER_17_1211 ();
 sg13g2_decap_8 FILLER_17_1218 ();
 sg13g2_decap_8 FILLER_17_1225 ();
 sg13g2_decap_8 FILLER_17_1232 ();
 sg13g2_decap_8 FILLER_17_1239 ();
 sg13g2_decap_8 FILLER_17_1246 ();
 sg13g2_decap_8 FILLER_17_1253 ();
 sg13g2_decap_8 FILLER_17_1260 ();
 sg13g2_decap_8 FILLER_17_1267 ();
 sg13g2_decap_8 FILLER_17_1274 ();
 sg13g2_decap_8 FILLER_17_1281 ();
 sg13g2_decap_8 FILLER_17_1288 ();
 sg13g2_decap_8 FILLER_17_1295 ();
 sg13g2_decap_8 FILLER_17_1302 ();
 sg13g2_decap_8 FILLER_17_1309 ();
 sg13g2_decap_8 FILLER_17_1316 ();
 sg13g2_decap_8 FILLER_17_1323 ();
 sg13g2_decap_8 FILLER_17_1330 ();
 sg13g2_decap_8 FILLER_17_1337 ();
 sg13g2_decap_8 FILLER_17_1344 ();
 sg13g2_decap_8 FILLER_17_1351 ();
 sg13g2_decap_8 FILLER_17_1358 ();
 sg13g2_decap_8 FILLER_17_1365 ();
 sg13g2_decap_8 FILLER_17_1372 ();
 sg13g2_decap_8 FILLER_17_1379 ();
 sg13g2_decap_8 FILLER_17_1386 ();
 sg13g2_decap_8 FILLER_17_1393 ();
 sg13g2_decap_8 FILLER_17_1400 ();
 sg13g2_decap_8 FILLER_17_1407 ();
 sg13g2_decap_8 FILLER_17_1414 ();
 sg13g2_decap_8 FILLER_17_1421 ();
 sg13g2_decap_8 FILLER_17_1428 ();
 sg13g2_decap_8 FILLER_17_1435 ();
 sg13g2_decap_8 FILLER_17_1442 ();
 sg13g2_decap_8 FILLER_17_1449 ();
 sg13g2_decap_8 FILLER_17_1456 ();
 sg13g2_decap_8 FILLER_17_1463 ();
 sg13g2_decap_8 FILLER_17_1470 ();
 sg13g2_decap_8 FILLER_17_1477 ();
 sg13g2_decap_8 FILLER_17_1484 ();
 sg13g2_decap_8 FILLER_17_1491 ();
 sg13g2_decap_8 FILLER_17_1498 ();
 sg13g2_decap_8 FILLER_17_1505 ();
 sg13g2_decap_8 FILLER_17_1512 ();
 sg13g2_decap_8 FILLER_17_1519 ();
 sg13g2_decap_8 FILLER_17_1526 ();
 sg13g2_decap_8 FILLER_17_1533 ();
 sg13g2_decap_8 FILLER_17_1540 ();
 sg13g2_decap_8 FILLER_17_1547 ();
 sg13g2_decap_8 FILLER_17_1554 ();
 sg13g2_decap_8 FILLER_17_1561 ();
 sg13g2_decap_8 FILLER_17_1568 ();
 sg13g2_decap_8 FILLER_17_1575 ();
 sg13g2_decap_8 FILLER_17_1582 ();
 sg13g2_decap_8 FILLER_17_1589 ();
 sg13g2_decap_8 FILLER_17_1596 ();
 sg13g2_decap_8 FILLER_17_1603 ();
 sg13g2_decap_8 FILLER_17_1610 ();
 sg13g2_decap_8 FILLER_17_1617 ();
 sg13g2_decap_8 FILLER_17_1624 ();
 sg13g2_decap_8 FILLER_17_1631 ();
 sg13g2_decap_8 FILLER_17_1638 ();
 sg13g2_decap_8 FILLER_17_1645 ();
 sg13g2_decap_8 FILLER_17_1652 ();
 sg13g2_decap_8 FILLER_17_1659 ();
 sg13g2_decap_8 FILLER_17_1666 ();
 sg13g2_decap_8 FILLER_17_1673 ();
 sg13g2_decap_8 FILLER_17_1680 ();
 sg13g2_decap_8 FILLER_17_1687 ();
 sg13g2_decap_8 FILLER_17_1694 ();
 sg13g2_decap_8 FILLER_17_1701 ();
 sg13g2_decap_8 FILLER_17_1708 ();
 sg13g2_decap_8 FILLER_17_1715 ();
 sg13g2_decap_8 FILLER_17_1722 ();
 sg13g2_decap_8 FILLER_17_1729 ();
 sg13g2_decap_8 FILLER_17_1736 ();
 sg13g2_decap_8 FILLER_17_1743 ();
 sg13g2_decap_8 FILLER_17_1750 ();
 sg13g2_decap_8 FILLER_17_1757 ();
 sg13g2_decap_8 FILLER_17_1764 ();
 sg13g2_decap_8 FILLER_17_1771 ();
 sg13g2_decap_8 FILLER_17_1778 ();
 sg13g2_decap_8 FILLER_17_1785 ();
 sg13g2_decap_8 FILLER_17_1792 ();
 sg13g2_decap_8 FILLER_17_1799 ();
 sg13g2_decap_8 FILLER_17_1806 ();
 sg13g2_decap_8 FILLER_17_1813 ();
 sg13g2_decap_8 FILLER_17_1820 ();
 sg13g2_decap_8 FILLER_17_1827 ();
 sg13g2_decap_8 FILLER_17_1834 ();
 sg13g2_decap_8 FILLER_17_1841 ();
 sg13g2_decap_8 FILLER_17_1848 ();
 sg13g2_decap_8 FILLER_17_1855 ();
 sg13g2_decap_8 FILLER_17_1862 ();
 sg13g2_decap_8 FILLER_17_1869 ();
 sg13g2_decap_8 FILLER_17_1876 ();
 sg13g2_decap_8 FILLER_17_1883 ();
 sg13g2_decap_8 FILLER_17_1890 ();
 sg13g2_decap_8 FILLER_17_1897 ();
 sg13g2_decap_8 FILLER_17_1904 ();
 sg13g2_decap_8 FILLER_17_1911 ();
 sg13g2_decap_8 FILLER_17_1918 ();
 sg13g2_decap_8 FILLER_17_1925 ();
 sg13g2_decap_8 FILLER_17_1932 ();
 sg13g2_decap_8 FILLER_17_1939 ();
 sg13g2_decap_8 FILLER_17_1946 ();
 sg13g2_decap_8 FILLER_17_1953 ();
 sg13g2_decap_8 FILLER_17_1960 ();
 sg13g2_decap_8 FILLER_17_1967 ();
 sg13g2_decap_8 FILLER_17_1974 ();
 sg13g2_decap_8 FILLER_17_1981 ();
 sg13g2_decap_8 FILLER_17_1988 ();
 sg13g2_decap_8 FILLER_17_1995 ();
 sg13g2_decap_8 FILLER_17_2002 ();
 sg13g2_decap_8 FILLER_17_2009 ();
 sg13g2_decap_8 FILLER_17_2016 ();
 sg13g2_decap_8 FILLER_17_2023 ();
 sg13g2_decap_8 FILLER_17_2030 ();
 sg13g2_decap_8 FILLER_17_2037 ();
 sg13g2_decap_8 FILLER_17_2044 ();
 sg13g2_decap_8 FILLER_17_2051 ();
 sg13g2_decap_8 FILLER_17_2058 ();
 sg13g2_decap_8 FILLER_17_2065 ();
 sg13g2_decap_8 FILLER_17_2072 ();
 sg13g2_decap_8 FILLER_17_2079 ();
 sg13g2_decap_8 FILLER_17_2086 ();
 sg13g2_decap_8 FILLER_17_2093 ();
 sg13g2_decap_8 FILLER_17_2100 ();
 sg13g2_decap_8 FILLER_17_2107 ();
 sg13g2_decap_8 FILLER_17_2114 ();
 sg13g2_decap_8 FILLER_17_2121 ();
 sg13g2_decap_8 FILLER_17_2128 ();
 sg13g2_decap_8 FILLER_17_2135 ();
 sg13g2_decap_8 FILLER_17_2142 ();
 sg13g2_decap_8 FILLER_17_2149 ();
 sg13g2_decap_8 FILLER_17_2156 ();
 sg13g2_decap_8 FILLER_17_2163 ();
 sg13g2_decap_8 FILLER_17_2170 ();
 sg13g2_decap_8 FILLER_17_2177 ();
 sg13g2_decap_8 FILLER_17_2184 ();
 sg13g2_decap_8 FILLER_17_2191 ();
 sg13g2_decap_8 FILLER_17_2198 ();
 sg13g2_decap_8 FILLER_17_2205 ();
 sg13g2_decap_8 FILLER_17_2212 ();
 sg13g2_decap_8 FILLER_17_2219 ();
 sg13g2_decap_8 FILLER_17_2226 ();
 sg13g2_decap_8 FILLER_17_2233 ();
 sg13g2_decap_8 FILLER_17_2240 ();
 sg13g2_decap_8 FILLER_17_2247 ();
 sg13g2_decap_8 FILLER_17_2254 ();
 sg13g2_decap_8 FILLER_17_2261 ();
 sg13g2_decap_8 FILLER_17_2268 ();
 sg13g2_decap_8 FILLER_17_2275 ();
 sg13g2_decap_8 FILLER_17_2282 ();
 sg13g2_decap_8 FILLER_17_2289 ();
 sg13g2_decap_8 FILLER_17_2296 ();
 sg13g2_decap_8 FILLER_17_2303 ();
 sg13g2_decap_8 FILLER_17_2310 ();
 sg13g2_decap_8 FILLER_17_2317 ();
 sg13g2_decap_8 FILLER_17_2324 ();
 sg13g2_decap_8 FILLER_17_2331 ();
 sg13g2_decap_8 FILLER_17_2338 ();
 sg13g2_decap_8 FILLER_17_2345 ();
 sg13g2_decap_8 FILLER_17_2352 ();
 sg13g2_decap_8 FILLER_17_2359 ();
 sg13g2_decap_8 FILLER_17_2366 ();
 sg13g2_decap_8 FILLER_17_2373 ();
 sg13g2_decap_8 FILLER_17_2380 ();
 sg13g2_decap_8 FILLER_17_2387 ();
 sg13g2_decap_8 FILLER_17_2394 ();
 sg13g2_decap_8 FILLER_17_2401 ();
 sg13g2_decap_8 FILLER_17_2408 ();
 sg13g2_decap_8 FILLER_17_2415 ();
 sg13g2_decap_8 FILLER_17_2422 ();
 sg13g2_decap_8 FILLER_17_2429 ();
 sg13g2_decap_8 FILLER_17_2436 ();
 sg13g2_decap_8 FILLER_17_2443 ();
 sg13g2_decap_8 FILLER_17_2450 ();
 sg13g2_decap_8 FILLER_17_2457 ();
 sg13g2_decap_8 FILLER_17_2464 ();
 sg13g2_decap_8 FILLER_17_2471 ();
 sg13g2_decap_8 FILLER_17_2478 ();
 sg13g2_decap_8 FILLER_17_2485 ();
 sg13g2_decap_8 FILLER_17_2492 ();
 sg13g2_decap_8 FILLER_17_2499 ();
 sg13g2_decap_8 FILLER_17_2506 ();
 sg13g2_decap_8 FILLER_17_2513 ();
 sg13g2_decap_8 FILLER_17_2520 ();
 sg13g2_decap_8 FILLER_17_2527 ();
 sg13g2_decap_8 FILLER_17_2534 ();
 sg13g2_decap_8 FILLER_17_2541 ();
 sg13g2_decap_8 FILLER_17_2548 ();
 sg13g2_decap_8 FILLER_17_2555 ();
 sg13g2_decap_8 FILLER_17_2562 ();
 sg13g2_decap_8 FILLER_17_2569 ();
 sg13g2_decap_8 FILLER_17_2576 ();
 sg13g2_decap_8 FILLER_17_2583 ();
 sg13g2_decap_8 FILLER_17_2590 ();
 sg13g2_decap_8 FILLER_17_2597 ();
 sg13g2_decap_8 FILLER_17_2604 ();
 sg13g2_decap_8 FILLER_17_2611 ();
 sg13g2_decap_8 FILLER_17_2618 ();
 sg13g2_decap_8 FILLER_17_2625 ();
 sg13g2_decap_8 FILLER_17_2632 ();
 sg13g2_decap_8 FILLER_17_2639 ();
 sg13g2_decap_8 FILLER_17_2646 ();
 sg13g2_decap_8 FILLER_17_2653 ();
 sg13g2_decap_8 FILLER_17_2660 ();
 sg13g2_decap_8 FILLER_17_2667 ();
 sg13g2_decap_8 FILLER_17_2674 ();
 sg13g2_decap_8 FILLER_17_2681 ();
 sg13g2_decap_8 FILLER_17_2688 ();
 sg13g2_decap_8 FILLER_17_2695 ();
 sg13g2_decap_8 FILLER_17_2702 ();
 sg13g2_decap_8 FILLER_17_2709 ();
 sg13g2_decap_8 FILLER_17_2716 ();
 sg13g2_decap_8 FILLER_17_2723 ();
 sg13g2_decap_8 FILLER_17_2730 ();
 sg13g2_decap_8 FILLER_17_2737 ();
 sg13g2_decap_8 FILLER_17_2744 ();
 sg13g2_decap_8 FILLER_17_2751 ();
 sg13g2_decap_8 FILLER_17_2758 ();
 sg13g2_decap_8 FILLER_17_2765 ();
 sg13g2_decap_8 FILLER_17_2772 ();
 sg13g2_decap_8 FILLER_17_2779 ();
 sg13g2_decap_8 FILLER_17_2786 ();
 sg13g2_decap_8 FILLER_17_2793 ();
 sg13g2_decap_8 FILLER_17_2800 ();
 sg13g2_decap_8 FILLER_17_2807 ();
 sg13g2_decap_8 FILLER_17_2814 ();
 sg13g2_decap_8 FILLER_17_2821 ();
 sg13g2_decap_8 FILLER_17_2828 ();
 sg13g2_decap_8 FILLER_17_2835 ();
 sg13g2_decap_8 FILLER_17_2842 ();
 sg13g2_decap_8 FILLER_17_2849 ();
 sg13g2_decap_8 FILLER_17_2856 ();
 sg13g2_decap_8 FILLER_17_2863 ();
 sg13g2_decap_8 FILLER_17_2870 ();
 sg13g2_decap_8 FILLER_17_2877 ();
 sg13g2_decap_8 FILLER_17_2884 ();
 sg13g2_decap_8 FILLER_17_2891 ();
 sg13g2_decap_8 FILLER_17_2898 ();
 sg13g2_decap_8 FILLER_17_2905 ();
 sg13g2_decap_8 FILLER_17_2912 ();
 sg13g2_decap_8 FILLER_17_2919 ();
 sg13g2_decap_8 FILLER_17_2926 ();
 sg13g2_decap_8 FILLER_17_2933 ();
 sg13g2_decap_8 FILLER_17_2940 ();
 sg13g2_decap_8 FILLER_17_2947 ();
 sg13g2_decap_8 FILLER_17_2954 ();
 sg13g2_decap_8 FILLER_17_2961 ();
 sg13g2_decap_8 FILLER_17_2968 ();
 sg13g2_decap_8 FILLER_17_2975 ();
 sg13g2_decap_8 FILLER_17_2982 ();
 sg13g2_decap_8 FILLER_17_2989 ();
 sg13g2_decap_8 FILLER_17_2996 ();
 sg13g2_decap_8 FILLER_17_3003 ();
 sg13g2_decap_8 FILLER_17_3010 ();
 sg13g2_decap_8 FILLER_17_3017 ();
 sg13g2_decap_8 FILLER_17_3024 ();
 sg13g2_decap_8 FILLER_17_3031 ();
 sg13g2_decap_8 FILLER_17_3038 ();
 sg13g2_decap_8 FILLER_17_3045 ();
 sg13g2_decap_8 FILLER_17_3052 ();
 sg13g2_decap_8 FILLER_17_3059 ();
 sg13g2_decap_8 FILLER_17_3066 ();
 sg13g2_decap_8 FILLER_17_3073 ();
 sg13g2_decap_8 FILLER_17_3080 ();
 sg13g2_decap_8 FILLER_17_3087 ();
 sg13g2_decap_8 FILLER_17_3094 ();
 sg13g2_decap_8 FILLER_17_3101 ();
 sg13g2_decap_8 FILLER_17_3108 ();
 sg13g2_decap_8 FILLER_17_3115 ();
 sg13g2_decap_8 FILLER_17_3122 ();
 sg13g2_decap_8 FILLER_17_3129 ();
 sg13g2_decap_8 FILLER_17_3136 ();
 sg13g2_decap_8 FILLER_17_3143 ();
 sg13g2_decap_8 FILLER_17_3150 ();
 sg13g2_decap_8 FILLER_17_3157 ();
 sg13g2_decap_8 FILLER_17_3164 ();
 sg13g2_decap_8 FILLER_17_3171 ();
 sg13g2_decap_8 FILLER_17_3178 ();
 sg13g2_decap_8 FILLER_17_3185 ();
 sg13g2_decap_8 FILLER_17_3192 ();
 sg13g2_decap_8 FILLER_17_3199 ();
 sg13g2_decap_8 FILLER_17_3206 ();
 sg13g2_decap_8 FILLER_17_3213 ();
 sg13g2_decap_8 FILLER_17_3220 ();
 sg13g2_decap_8 FILLER_17_3227 ();
 sg13g2_decap_8 FILLER_17_3234 ();
 sg13g2_decap_8 FILLER_17_3241 ();
 sg13g2_decap_8 FILLER_17_3248 ();
 sg13g2_decap_8 FILLER_17_3255 ();
 sg13g2_decap_8 FILLER_17_3262 ();
 sg13g2_decap_8 FILLER_17_3269 ();
 sg13g2_decap_8 FILLER_17_3276 ();
 sg13g2_decap_8 FILLER_17_3283 ();
 sg13g2_decap_8 FILLER_17_3290 ();
 sg13g2_decap_8 FILLER_17_3297 ();
 sg13g2_decap_8 FILLER_17_3304 ();
 sg13g2_decap_8 FILLER_17_3311 ();
 sg13g2_decap_8 FILLER_17_3318 ();
 sg13g2_decap_8 FILLER_17_3325 ();
 sg13g2_decap_8 FILLER_17_3332 ();
 sg13g2_decap_8 FILLER_17_3339 ();
 sg13g2_decap_8 FILLER_17_3346 ();
 sg13g2_decap_8 FILLER_17_3353 ();
 sg13g2_decap_8 FILLER_17_3360 ();
 sg13g2_decap_8 FILLER_17_3367 ();
 sg13g2_decap_8 FILLER_17_3374 ();
 sg13g2_decap_8 FILLER_17_3381 ();
 sg13g2_decap_8 FILLER_17_3388 ();
 sg13g2_decap_8 FILLER_17_3395 ();
 sg13g2_decap_8 FILLER_17_3402 ();
 sg13g2_decap_8 FILLER_17_3409 ();
 sg13g2_decap_8 FILLER_17_3416 ();
 sg13g2_decap_8 FILLER_17_3423 ();
 sg13g2_decap_8 FILLER_17_3430 ();
 sg13g2_decap_8 FILLER_17_3437 ();
 sg13g2_decap_8 FILLER_17_3444 ();
 sg13g2_decap_8 FILLER_17_3451 ();
 sg13g2_decap_8 FILLER_17_3458 ();
 sg13g2_decap_8 FILLER_17_3465 ();
 sg13g2_decap_8 FILLER_17_3472 ();
 sg13g2_decap_8 FILLER_17_3479 ();
 sg13g2_decap_8 FILLER_17_3486 ();
 sg13g2_decap_8 FILLER_17_3493 ();
 sg13g2_decap_8 FILLER_17_3500 ();
 sg13g2_decap_8 FILLER_17_3507 ();
 sg13g2_decap_8 FILLER_17_3514 ();
 sg13g2_decap_8 FILLER_17_3521 ();
 sg13g2_decap_8 FILLER_17_3528 ();
 sg13g2_decap_8 FILLER_17_3535 ();
 sg13g2_decap_8 FILLER_17_3542 ();
 sg13g2_decap_8 FILLER_17_3549 ();
 sg13g2_decap_8 FILLER_17_3556 ();
 sg13g2_decap_8 FILLER_17_3563 ();
 sg13g2_decap_8 FILLER_17_3570 ();
 sg13g2_fill_2 FILLER_17_3577 ();
 sg13g2_fill_1 FILLER_17_3579 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_8 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_decap_8 FILLER_18_427 ();
 sg13g2_decap_8 FILLER_18_434 ();
 sg13g2_decap_8 FILLER_18_441 ();
 sg13g2_decap_8 FILLER_18_448 ();
 sg13g2_decap_8 FILLER_18_455 ();
 sg13g2_decap_8 FILLER_18_462 ();
 sg13g2_decap_8 FILLER_18_469 ();
 sg13g2_decap_8 FILLER_18_476 ();
 sg13g2_decap_8 FILLER_18_483 ();
 sg13g2_decap_8 FILLER_18_490 ();
 sg13g2_decap_8 FILLER_18_497 ();
 sg13g2_decap_8 FILLER_18_504 ();
 sg13g2_decap_8 FILLER_18_511 ();
 sg13g2_decap_8 FILLER_18_518 ();
 sg13g2_decap_8 FILLER_18_525 ();
 sg13g2_decap_8 FILLER_18_532 ();
 sg13g2_decap_8 FILLER_18_539 ();
 sg13g2_decap_8 FILLER_18_546 ();
 sg13g2_decap_8 FILLER_18_553 ();
 sg13g2_decap_8 FILLER_18_560 ();
 sg13g2_decap_8 FILLER_18_567 ();
 sg13g2_decap_8 FILLER_18_574 ();
 sg13g2_decap_8 FILLER_18_581 ();
 sg13g2_decap_8 FILLER_18_588 ();
 sg13g2_decap_8 FILLER_18_595 ();
 sg13g2_decap_8 FILLER_18_602 ();
 sg13g2_decap_8 FILLER_18_609 ();
 sg13g2_decap_8 FILLER_18_616 ();
 sg13g2_decap_8 FILLER_18_623 ();
 sg13g2_decap_8 FILLER_18_630 ();
 sg13g2_decap_8 FILLER_18_637 ();
 sg13g2_decap_8 FILLER_18_644 ();
 sg13g2_decap_8 FILLER_18_651 ();
 sg13g2_decap_8 FILLER_18_658 ();
 sg13g2_decap_8 FILLER_18_665 ();
 sg13g2_decap_8 FILLER_18_672 ();
 sg13g2_decap_8 FILLER_18_679 ();
 sg13g2_decap_8 FILLER_18_686 ();
 sg13g2_decap_8 FILLER_18_693 ();
 sg13g2_decap_8 FILLER_18_700 ();
 sg13g2_decap_8 FILLER_18_707 ();
 sg13g2_decap_8 FILLER_18_714 ();
 sg13g2_decap_8 FILLER_18_721 ();
 sg13g2_decap_8 FILLER_18_728 ();
 sg13g2_decap_8 FILLER_18_735 ();
 sg13g2_decap_8 FILLER_18_742 ();
 sg13g2_decap_8 FILLER_18_749 ();
 sg13g2_decap_8 FILLER_18_756 ();
 sg13g2_decap_8 FILLER_18_763 ();
 sg13g2_decap_8 FILLER_18_770 ();
 sg13g2_decap_8 FILLER_18_777 ();
 sg13g2_decap_8 FILLER_18_784 ();
 sg13g2_decap_8 FILLER_18_791 ();
 sg13g2_decap_8 FILLER_18_798 ();
 sg13g2_decap_8 FILLER_18_805 ();
 sg13g2_decap_8 FILLER_18_812 ();
 sg13g2_decap_8 FILLER_18_819 ();
 sg13g2_decap_8 FILLER_18_826 ();
 sg13g2_decap_8 FILLER_18_833 ();
 sg13g2_decap_8 FILLER_18_840 ();
 sg13g2_decap_8 FILLER_18_847 ();
 sg13g2_decap_8 FILLER_18_854 ();
 sg13g2_decap_8 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_18_868 ();
 sg13g2_decap_8 FILLER_18_875 ();
 sg13g2_decap_8 FILLER_18_882 ();
 sg13g2_decap_8 FILLER_18_889 ();
 sg13g2_decap_8 FILLER_18_896 ();
 sg13g2_decap_8 FILLER_18_903 ();
 sg13g2_decap_8 FILLER_18_910 ();
 sg13g2_decap_8 FILLER_18_917 ();
 sg13g2_decap_8 FILLER_18_924 ();
 sg13g2_decap_8 FILLER_18_931 ();
 sg13g2_decap_8 FILLER_18_938 ();
 sg13g2_decap_8 FILLER_18_945 ();
 sg13g2_decap_8 FILLER_18_952 ();
 sg13g2_decap_8 FILLER_18_959 ();
 sg13g2_decap_8 FILLER_18_966 ();
 sg13g2_decap_8 FILLER_18_973 ();
 sg13g2_decap_8 FILLER_18_980 ();
 sg13g2_decap_8 FILLER_18_987 ();
 sg13g2_decap_8 FILLER_18_994 ();
 sg13g2_decap_8 FILLER_18_1001 ();
 sg13g2_decap_8 FILLER_18_1008 ();
 sg13g2_decap_8 FILLER_18_1015 ();
 sg13g2_decap_8 FILLER_18_1022 ();
 sg13g2_decap_8 FILLER_18_1029 ();
 sg13g2_decap_8 FILLER_18_1036 ();
 sg13g2_decap_8 FILLER_18_1043 ();
 sg13g2_decap_8 FILLER_18_1050 ();
 sg13g2_decap_8 FILLER_18_1057 ();
 sg13g2_decap_8 FILLER_18_1064 ();
 sg13g2_decap_8 FILLER_18_1071 ();
 sg13g2_decap_8 FILLER_18_1078 ();
 sg13g2_decap_8 FILLER_18_1085 ();
 sg13g2_decap_8 FILLER_18_1092 ();
 sg13g2_decap_8 FILLER_18_1099 ();
 sg13g2_decap_8 FILLER_18_1106 ();
 sg13g2_decap_8 FILLER_18_1113 ();
 sg13g2_decap_8 FILLER_18_1120 ();
 sg13g2_decap_8 FILLER_18_1127 ();
 sg13g2_decap_8 FILLER_18_1134 ();
 sg13g2_decap_8 FILLER_18_1141 ();
 sg13g2_decap_8 FILLER_18_1148 ();
 sg13g2_decap_8 FILLER_18_1155 ();
 sg13g2_decap_8 FILLER_18_1162 ();
 sg13g2_decap_8 FILLER_18_1169 ();
 sg13g2_decap_8 FILLER_18_1176 ();
 sg13g2_decap_8 FILLER_18_1183 ();
 sg13g2_decap_8 FILLER_18_1190 ();
 sg13g2_decap_8 FILLER_18_1197 ();
 sg13g2_decap_8 FILLER_18_1204 ();
 sg13g2_decap_8 FILLER_18_1211 ();
 sg13g2_decap_8 FILLER_18_1218 ();
 sg13g2_decap_8 FILLER_18_1225 ();
 sg13g2_decap_8 FILLER_18_1232 ();
 sg13g2_decap_8 FILLER_18_1239 ();
 sg13g2_decap_8 FILLER_18_1246 ();
 sg13g2_decap_8 FILLER_18_1253 ();
 sg13g2_decap_8 FILLER_18_1260 ();
 sg13g2_decap_8 FILLER_18_1267 ();
 sg13g2_decap_8 FILLER_18_1274 ();
 sg13g2_decap_8 FILLER_18_1281 ();
 sg13g2_decap_8 FILLER_18_1288 ();
 sg13g2_decap_8 FILLER_18_1295 ();
 sg13g2_decap_8 FILLER_18_1302 ();
 sg13g2_decap_8 FILLER_18_1309 ();
 sg13g2_decap_8 FILLER_18_1316 ();
 sg13g2_decap_8 FILLER_18_1323 ();
 sg13g2_decap_8 FILLER_18_1330 ();
 sg13g2_decap_8 FILLER_18_1337 ();
 sg13g2_decap_8 FILLER_18_1344 ();
 sg13g2_decap_8 FILLER_18_1351 ();
 sg13g2_decap_8 FILLER_18_1358 ();
 sg13g2_decap_8 FILLER_18_1365 ();
 sg13g2_decap_8 FILLER_18_1372 ();
 sg13g2_decap_8 FILLER_18_1379 ();
 sg13g2_decap_8 FILLER_18_1386 ();
 sg13g2_decap_8 FILLER_18_1393 ();
 sg13g2_decap_8 FILLER_18_1400 ();
 sg13g2_decap_8 FILLER_18_1407 ();
 sg13g2_decap_8 FILLER_18_1414 ();
 sg13g2_decap_8 FILLER_18_1421 ();
 sg13g2_decap_8 FILLER_18_1428 ();
 sg13g2_decap_8 FILLER_18_1435 ();
 sg13g2_decap_8 FILLER_18_1442 ();
 sg13g2_decap_8 FILLER_18_1449 ();
 sg13g2_decap_8 FILLER_18_1456 ();
 sg13g2_decap_8 FILLER_18_1463 ();
 sg13g2_decap_8 FILLER_18_1470 ();
 sg13g2_decap_8 FILLER_18_1477 ();
 sg13g2_decap_8 FILLER_18_1484 ();
 sg13g2_decap_8 FILLER_18_1491 ();
 sg13g2_decap_8 FILLER_18_1498 ();
 sg13g2_decap_8 FILLER_18_1505 ();
 sg13g2_decap_8 FILLER_18_1512 ();
 sg13g2_decap_8 FILLER_18_1519 ();
 sg13g2_decap_8 FILLER_18_1526 ();
 sg13g2_decap_8 FILLER_18_1533 ();
 sg13g2_decap_8 FILLER_18_1540 ();
 sg13g2_decap_8 FILLER_18_1547 ();
 sg13g2_decap_8 FILLER_18_1554 ();
 sg13g2_decap_8 FILLER_18_1561 ();
 sg13g2_decap_8 FILLER_18_1568 ();
 sg13g2_decap_8 FILLER_18_1575 ();
 sg13g2_decap_8 FILLER_18_1582 ();
 sg13g2_decap_8 FILLER_18_1589 ();
 sg13g2_decap_8 FILLER_18_1596 ();
 sg13g2_decap_8 FILLER_18_1603 ();
 sg13g2_decap_8 FILLER_18_1610 ();
 sg13g2_decap_8 FILLER_18_1617 ();
 sg13g2_decap_8 FILLER_18_1624 ();
 sg13g2_decap_8 FILLER_18_1631 ();
 sg13g2_decap_8 FILLER_18_1638 ();
 sg13g2_decap_8 FILLER_18_1645 ();
 sg13g2_decap_8 FILLER_18_1652 ();
 sg13g2_decap_8 FILLER_18_1659 ();
 sg13g2_decap_8 FILLER_18_1666 ();
 sg13g2_decap_8 FILLER_18_1673 ();
 sg13g2_decap_8 FILLER_18_1680 ();
 sg13g2_decap_8 FILLER_18_1687 ();
 sg13g2_decap_8 FILLER_18_1694 ();
 sg13g2_decap_8 FILLER_18_1701 ();
 sg13g2_decap_8 FILLER_18_1708 ();
 sg13g2_decap_8 FILLER_18_1715 ();
 sg13g2_decap_8 FILLER_18_1722 ();
 sg13g2_decap_8 FILLER_18_1729 ();
 sg13g2_decap_8 FILLER_18_1736 ();
 sg13g2_decap_8 FILLER_18_1743 ();
 sg13g2_decap_8 FILLER_18_1750 ();
 sg13g2_decap_8 FILLER_18_1757 ();
 sg13g2_decap_8 FILLER_18_1764 ();
 sg13g2_decap_8 FILLER_18_1771 ();
 sg13g2_decap_8 FILLER_18_1778 ();
 sg13g2_decap_8 FILLER_18_1785 ();
 sg13g2_decap_8 FILLER_18_1792 ();
 sg13g2_decap_8 FILLER_18_1799 ();
 sg13g2_decap_8 FILLER_18_1806 ();
 sg13g2_decap_8 FILLER_18_1813 ();
 sg13g2_decap_8 FILLER_18_1820 ();
 sg13g2_decap_8 FILLER_18_1827 ();
 sg13g2_decap_8 FILLER_18_1834 ();
 sg13g2_decap_8 FILLER_18_1841 ();
 sg13g2_decap_8 FILLER_18_1848 ();
 sg13g2_decap_8 FILLER_18_1855 ();
 sg13g2_decap_8 FILLER_18_1862 ();
 sg13g2_decap_8 FILLER_18_1869 ();
 sg13g2_decap_8 FILLER_18_1876 ();
 sg13g2_decap_8 FILLER_18_1883 ();
 sg13g2_decap_8 FILLER_18_1890 ();
 sg13g2_decap_8 FILLER_18_1897 ();
 sg13g2_decap_8 FILLER_18_1904 ();
 sg13g2_decap_8 FILLER_18_1911 ();
 sg13g2_decap_8 FILLER_18_1918 ();
 sg13g2_decap_8 FILLER_18_1925 ();
 sg13g2_decap_8 FILLER_18_1932 ();
 sg13g2_decap_8 FILLER_18_1939 ();
 sg13g2_decap_8 FILLER_18_1946 ();
 sg13g2_decap_8 FILLER_18_1953 ();
 sg13g2_decap_8 FILLER_18_1960 ();
 sg13g2_decap_8 FILLER_18_1967 ();
 sg13g2_decap_8 FILLER_18_1974 ();
 sg13g2_decap_8 FILLER_18_1981 ();
 sg13g2_decap_8 FILLER_18_1988 ();
 sg13g2_decap_8 FILLER_18_1995 ();
 sg13g2_decap_8 FILLER_18_2002 ();
 sg13g2_decap_8 FILLER_18_2009 ();
 sg13g2_decap_8 FILLER_18_2016 ();
 sg13g2_decap_8 FILLER_18_2023 ();
 sg13g2_decap_8 FILLER_18_2030 ();
 sg13g2_decap_8 FILLER_18_2037 ();
 sg13g2_decap_8 FILLER_18_2044 ();
 sg13g2_decap_8 FILLER_18_2051 ();
 sg13g2_decap_8 FILLER_18_2058 ();
 sg13g2_decap_8 FILLER_18_2065 ();
 sg13g2_decap_8 FILLER_18_2072 ();
 sg13g2_decap_8 FILLER_18_2079 ();
 sg13g2_decap_8 FILLER_18_2086 ();
 sg13g2_decap_8 FILLER_18_2093 ();
 sg13g2_decap_8 FILLER_18_2100 ();
 sg13g2_decap_8 FILLER_18_2107 ();
 sg13g2_decap_8 FILLER_18_2114 ();
 sg13g2_decap_8 FILLER_18_2121 ();
 sg13g2_decap_8 FILLER_18_2128 ();
 sg13g2_decap_8 FILLER_18_2135 ();
 sg13g2_decap_8 FILLER_18_2142 ();
 sg13g2_decap_8 FILLER_18_2149 ();
 sg13g2_decap_8 FILLER_18_2156 ();
 sg13g2_decap_8 FILLER_18_2163 ();
 sg13g2_decap_8 FILLER_18_2170 ();
 sg13g2_decap_8 FILLER_18_2177 ();
 sg13g2_decap_8 FILLER_18_2184 ();
 sg13g2_decap_8 FILLER_18_2191 ();
 sg13g2_decap_8 FILLER_18_2198 ();
 sg13g2_decap_8 FILLER_18_2205 ();
 sg13g2_decap_8 FILLER_18_2212 ();
 sg13g2_decap_8 FILLER_18_2219 ();
 sg13g2_decap_8 FILLER_18_2226 ();
 sg13g2_decap_8 FILLER_18_2233 ();
 sg13g2_decap_8 FILLER_18_2240 ();
 sg13g2_decap_8 FILLER_18_2247 ();
 sg13g2_decap_8 FILLER_18_2254 ();
 sg13g2_decap_8 FILLER_18_2261 ();
 sg13g2_decap_8 FILLER_18_2268 ();
 sg13g2_decap_8 FILLER_18_2275 ();
 sg13g2_decap_8 FILLER_18_2282 ();
 sg13g2_decap_8 FILLER_18_2289 ();
 sg13g2_decap_8 FILLER_18_2296 ();
 sg13g2_decap_8 FILLER_18_2303 ();
 sg13g2_decap_8 FILLER_18_2310 ();
 sg13g2_decap_8 FILLER_18_2317 ();
 sg13g2_decap_8 FILLER_18_2324 ();
 sg13g2_decap_8 FILLER_18_2331 ();
 sg13g2_decap_8 FILLER_18_2338 ();
 sg13g2_decap_8 FILLER_18_2345 ();
 sg13g2_decap_8 FILLER_18_2352 ();
 sg13g2_decap_8 FILLER_18_2359 ();
 sg13g2_decap_8 FILLER_18_2366 ();
 sg13g2_decap_8 FILLER_18_2373 ();
 sg13g2_decap_8 FILLER_18_2380 ();
 sg13g2_decap_8 FILLER_18_2387 ();
 sg13g2_decap_8 FILLER_18_2394 ();
 sg13g2_decap_8 FILLER_18_2401 ();
 sg13g2_decap_8 FILLER_18_2408 ();
 sg13g2_decap_8 FILLER_18_2415 ();
 sg13g2_decap_8 FILLER_18_2422 ();
 sg13g2_decap_8 FILLER_18_2429 ();
 sg13g2_decap_8 FILLER_18_2436 ();
 sg13g2_decap_8 FILLER_18_2443 ();
 sg13g2_decap_8 FILLER_18_2450 ();
 sg13g2_decap_8 FILLER_18_2457 ();
 sg13g2_decap_8 FILLER_18_2464 ();
 sg13g2_decap_8 FILLER_18_2471 ();
 sg13g2_decap_8 FILLER_18_2478 ();
 sg13g2_decap_8 FILLER_18_2485 ();
 sg13g2_decap_8 FILLER_18_2492 ();
 sg13g2_decap_8 FILLER_18_2499 ();
 sg13g2_decap_8 FILLER_18_2506 ();
 sg13g2_decap_8 FILLER_18_2513 ();
 sg13g2_decap_8 FILLER_18_2520 ();
 sg13g2_decap_8 FILLER_18_2527 ();
 sg13g2_decap_8 FILLER_18_2534 ();
 sg13g2_decap_8 FILLER_18_2541 ();
 sg13g2_decap_8 FILLER_18_2548 ();
 sg13g2_decap_8 FILLER_18_2555 ();
 sg13g2_decap_8 FILLER_18_2562 ();
 sg13g2_decap_8 FILLER_18_2569 ();
 sg13g2_decap_8 FILLER_18_2576 ();
 sg13g2_decap_8 FILLER_18_2583 ();
 sg13g2_decap_8 FILLER_18_2590 ();
 sg13g2_decap_8 FILLER_18_2597 ();
 sg13g2_decap_8 FILLER_18_2604 ();
 sg13g2_decap_8 FILLER_18_2611 ();
 sg13g2_decap_8 FILLER_18_2618 ();
 sg13g2_decap_8 FILLER_18_2625 ();
 sg13g2_decap_8 FILLER_18_2632 ();
 sg13g2_decap_8 FILLER_18_2639 ();
 sg13g2_decap_8 FILLER_18_2646 ();
 sg13g2_decap_8 FILLER_18_2653 ();
 sg13g2_decap_8 FILLER_18_2660 ();
 sg13g2_decap_8 FILLER_18_2667 ();
 sg13g2_decap_8 FILLER_18_2674 ();
 sg13g2_decap_8 FILLER_18_2681 ();
 sg13g2_decap_8 FILLER_18_2688 ();
 sg13g2_decap_8 FILLER_18_2695 ();
 sg13g2_decap_8 FILLER_18_2702 ();
 sg13g2_decap_8 FILLER_18_2709 ();
 sg13g2_decap_8 FILLER_18_2716 ();
 sg13g2_decap_8 FILLER_18_2723 ();
 sg13g2_decap_8 FILLER_18_2730 ();
 sg13g2_decap_8 FILLER_18_2737 ();
 sg13g2_decap_8 FILLER_18_2744 ();
 sg13g2_decap_8 FILLER_18_2751 ();
 sg13g2_decap_8 FILLER_18_2758 ();
 sg13g2_decap_8 FILLER_18_2765 ();
 sg13g2_decap_8 FILLER_18_2772 ();
 sg13g2_decap_8 FILLER_18_2779 ();
 sg13g2_decap_8 FILLER_18_2786 ();
 sg13g2_decap_8 FILLER_18_2793 ();
 sg13g2_decap_8 FILLER_18_2800 ();
 sg13g2_decap_8 FILLER_18_2807 ();
 sg13g2_decap_8 FILLER_18_2814 ();
 sg13g2_decap_8 FILLER_18_2821 ();
 sg13g2_decap_8 FILLER_18_2828 ();
 sg13g2_decap_8 FILLER_18_2835 ();
 sg13g2_decap_8 FILLER_18_2842 ();
 sg13g2_decap_8 FILLER_18_2849 ();
 sg13g2_decap_8 FILLER_18_2856 ();
 sg13g2_decap_8 FILLER_18_2863 ();
 sg13g2_decap_8 FILLER_18_2870 ();
 sg13g2_decap_8 FILLER_18_2877 ();
 sg13g2_decap_8 FILLER_18_2884 ();
 sg13g2_decap_8 FILLER_18_2891 ();
 sg13g2_decap_8 FILLER_18_2898 ();
 sg13g2_decap_8 FILLER_18_2905 ();
 sg13g2_decap_8 FILLER_18_2912 ();
 sg13g2_decap_8 FILLER_18_2919 ();
 sg13g2_decap_8 FILLER_18_2926 ();
 sg13g2_decap_8 FILLER_18_2933 ();
 sg13g2_decap_8 FILLER_18_2940 ();
 sg13g2_decap_8 FILLER_18_2947 ();
 sg13g2_decap_8 FILLER_18_2954 ();
 sg13g2_decap_8 FILLER_18_2961 ();
 sg13g2_decap_8 FILLER_18_2968 ();
 sg13g2_decap_8 FILLER_18_2975 ();
 sg13g2_decap_8 FILLER_18_2982 ();
 sg13g2_decap_8 FILLER_18_2989 ();
 sg13g2_decap_8 FILLER_18_2996 ();
 sg13g2_decap_8 FILLER_18_3003 ();
 sg13g2_decap_8 FILLER_18_3010 ();
 sg13g2_decap_8 FILLER_18_3017 ();
 sg13g2_decap_8 FILLER_18_3024 ();
 sg13g2_decap_8 FILLER_18_3031 ();
 sg13g2_decap_8 FILLER_18_3038 ();
 sg13g2_decap_8 FILLER_18_3045 ();
 sg13g2_decap_8 FILLER_18_3052 ();
 sg13g2_decap_8 FILLER_18_3059 ();
 sg13g2_decap_8 FILLER_18_3066 ();
 sg13g2_decap_8 FILLER_18_3073 ();
 sg13g2_decap_8 FILLER_18_3080 ();
 sg13g2_decap_8 FILLER_18_3087 ();
 sg13g2_decap_8 FILLER_18_3094 ();
 sg13g2_decap_8 FILLER_18_3101 ();
 sg13g2_decap_8 FILLER_18_3108 ();
 sg13g2_decap_8 FILLER_18_3115 ();
 sg13g2_decap_8 FILLER_18_3122 ();
 sg13g2_decap_8 FILLER_18_3129 ();
 sg13g2_decap_8 FILLER_18_3136 ();
 sg13g2_decap_8 FILLER_18_3143 ();
 sg13g2_decap_8 FILLER_18_3150 ();
 sg13g2_decap_8 FILLER_18_3157 ();
 sg13g2_decap_8 FILLER_18_3164 ();
 sg13g2_decap_8 FILLER_18_3171 ();
 sg13g2_decap_8 FILLER_18_3178 ();
 sg13g2_decap_8 FILLER_18_3185 ();
 sg13g2_decap_8 FILLER_18_3192 ();
 sg13g2_decap_8 FILLER_18_3199 ();
 sg13g2_decap_8 FILLER_18_3206 ();
 sg13g2_decap_8 FILLER_18_3213 ();
 sg13g2_decap_8 FILLER_18_3220 ();
 sg13g2_decap_8 FILLER_18_3227 ();
 sg13g2_decap_8 FILLER_18_3234 ();
 sg13g2_decap_8 FILLER_18_3241 ();
 sg13g2_decap_8 FILLER_18_3248 ();
 sg13g2_decap_8 FILLER_18_3255 ();
 sg13g2_decap_8 FILLER_18_3262 ();
 sg13g2_decap_8 FILLER_18_3269 ();
 sg13g2_decap_8 FILLER_18_3276 ();
 sg13g2_decap_8 FILLER_18_3283 ();
 sg13g2_decap_8 FILLER_18_3290 ();
 sg13g2_decap_8 FILLER_18_3297 ();
 sg13g2_decap_8 FILLER_18_3304 ();
 sg13g2_decap_8 FILLER_18_3311 ();
 sg13g2_decap_8 FILLER_18_3318 ();
 sg13g2_decap_8 FILLER_18_3325 ();
 sg13g2_decap_8 FILLER_18_3332 ();
 sg13g2_decap_8 FILLER_18_3339 ();
 sg13g2_decap_8 FILLER_18_3346 ();
 sg13g2_decap_8 FILLER_18_3353 ();
 sg13g2_decap_8 FILLER_18_3360 ();
 sg13g2_decap_8 FILLER_18_3367 ();
 sg13g2_decap_8 FILLER_18_3374 ();
 sg13g2_decap_8 FILLER_18_3381 ();
 sg13g2_decap_8 FILLER_18_3388 ();
 sg13g2_decap_8 FILLER_18_3395 ();
 sg13g2_decap_8 FILLER_18_3402 ();
 sg13g2_decap_8 FILLER_18_3409 ();
 sg13g2_decap_8 FILLER_18_3416 ();
 sg13g2_decap_8 FILLER_18_3423 ();
 sg13g2_decap_8 FILLER_18_3430 ();
 sg13g2_decap_8 FILLER_18_3437 ();
 sg13g2_decap_8 FILLER_18_3444 ();
 sg13g2_decap_8 FILLER_18_3451 ();
 sg13g2_decap_8 FILLER_18_3458 ();
 sg13g2_decap_8 FILLER_18_3465 ();
 sg13g2_decap_8 FILLER_18_3472 ();
 sg13g2_decap_8 FILLER_18_3479 ();
 sg13g2_decap_8 FILLER_18_3486 ();
 sg13g2_decap_8 FILLER_18_3493 ();
 sg13g2_decap_8 FILLER_18_3500 ();
 sg13g2_decap_8 FILLER_18_3507 ();
 sg13g2_decap_8 FILLER_18_3514 ();
 sg13g2_decap_8 FILLER_18_3521 ();
 sg13g2_decap_8 FILLER_18_3528 ();
 sg13g2_decap_8 FILLER_18_3535 ();
 sg13g2_decap_8 FILLER_18_3542 ();
 sg13g2_decap_8 FILLER_18_3549 ();
 sg13g2_decap_8 FILLER_18_3556 ();
 sg13g2_decap_8 FILLER_18_3563 ();
 sg13g2_decap_8 FILLER_18_3570 ();
 sg13g2_fill_2 FILLER_18_3577 ();
 sg13g2_fill_1 FILLER_18_3579 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_decap_8 FILLER_19_427 ();
 sg13g2_decap_8 FILLER_19_434 ();
 sg13g2_decap_8 FILLER_19_441 ();
 sg13g2_decap_8 FILLER_19_448 ();
 sg13g2_decap_8 FILLER_19_455 ();
 sg13g2_decap_8 FILLER_19_462 ();
 sg13g2_decap_8 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_476 ();
 sg13g2_decap_8 FILLER_19_483 ();
 sg13g2_decap_8 FILLER_19_490 ();
 sg13g2_decap_8 FILLER_19_497 ();
 sg13g2_decap_8 FILLER_19_504 ();
 sg13g2_decap_8 FILLER_19_511 ();
 sg13g2_decap_8 FILLER_19_518 ();
 sg13g2_decap_8 FILLER_19_525 ();
 sg13g2_decap_8 FILLER_19_532 ();
 sg13g2_decap_8 FILLER_19_539 ();
 sg13g2_decap_8 FILLER_19_546 ();
 sg13g2_decap_8 FILLER_19_553 ();
 sg13g2_decap_8 FILLER_19_560 ();
 sg13g2_decap_8 FILLER_19_567 ();
 sg13g2_decap_8 FILLER_19_574 ();
 sg13g2_decap_8 FILLER_19_581 ();
 sg13g2_decap_8 FILLER_19_588 ();
 sg13g2_decap_8 FILLER_19_595 ();
 sg13g2_decap_8 FILLER_19_602 ();
 sg13g2_decap_8 FILLER_19_609 ();
 sg13g2_decap_8 FILLER_19_616 ();
 sg13g2_decap_8 FILLER_19_623 ();
 sg13g2_decap_8 FILLER_19_630 ();
 sg13g2_decap_8 FILLER_19_637 ();
 sg13g2_decap_8 FILLER_19_644 ();
 sg13g2_decap_8 FILLER_19_651 ();
 sg13g2_decap_8 FILLER_19_658 ();
 sg13g2_decap_8 FILLER_19_665 ();
 sg13g2_decap_8 FILLER_19_672 ();
 sg13g2_decap_8 FILLER_19_679 ();
 sg13g2_decap_8 FILLER_19_686 ();
 sg13g2_decap_8 FILLER_19_693 ();
 sg13g2_decap_8 FILLER_19_700 ();
 sg13g2_decap_8 FILLER_19_707 ();
 sg13g2_decap_8 FILLER_19_714 ();
 sg13g2_decap_8 FILLER_19_721 ();
 sg13g2_decap_8 FILLER_19_728 ();
 sg13g2_decap_8 FILLER_19_735 ();
 sg13g2_decap_8 FILLER_19_742 ();
 sg13g2_decap_8 FILLER_19_749 ();
 sg13g2_decap_8 FILLER_19_756 ();
 sg13g2_decap_8 FILLER_19_763 ();
 sg13g2_decap_8 FILLER_19_770 ();
 sg13g2_decap_8 FILLER_19_777 ();
 sg13g2_decap_8 FILLER_19_784 ();
 sg13g2_decap_8 FILLER_19_791 ();
 sg13g2_decap_8 FILLER_19_798 ();
 sg13g2_decap_8 FILLER_19_805 ();
 sg13g2_decap_8 FILLER_19_812 ();
 sg13g2_decap_8 FILLER_19_819 ();
 sg13g2_decap_8 FILLER_19_826 ();
 sg13g2_decap_8 FILLER_19_833 ();
 sg13g2_decap_8 FILLER_19_840 ();
 sg13g2_decap_8 FILLER_19_847 ();
 sg13g2_decap_8 FILLER_19_854 ();
 sg13g2_decap_8 FILLER_19_861 ();
 sg13g2_decap_8 FILLER_19_868 ();
 sg13g2_decap_8 FILLER_19_875 ();
 sg13g2_decap_8 FILLER_19_882 ();
 sg13g2_decap_8 FILLER_19_889 ();
 sg13g2_decap_8 FILLER_19_896 ();
 sg13g2_decap_8 FILLER_19_903 ();
 sg13g2_decap_8 FILLER_19_910 ();
 sg13g2_decap_8 FILLER_19_917 ();
 sg13g2_decap_8 FILLER_19_924 ();
 sg13g2_decap_8 FILLER_19_931 ();
 sg13g2_decap_8 FILLER_19_938 ();
 sg13g2_decap_8 FILLER_19_945 ();
 sg13g2_decap_8 FILLER_19_952 ();
 sg13g2_decap_8 FILLER_19_959 ();
 sg13g2_decap_8 FILLER_19_966 ();
 sg13g2_decap_8 FILLER_19_973 ();
 sg13g2_decap_8 FILLER_19_980 ();
 sg13g2_decap_8 FILLER_19_987 ();
 sg13g2_decap_8 FILLER_19_994 ();
 sg13g2_decap_8 FILLER_19_1001 ();
 sg13g2_decap_8 FILLER_19_1008 ();
 sg13g2_decap_8 FILLER_19_1015 ();
 sg13g2_decap_8 FILLER_19_1022 ();
 sg13g2_decap_8 FILLER_19_1029 ();
 sg13g2_decap_8 FILLER_19_1036 ();
 sg13g2_decap_8 FILLER_19_1043 ();
 sg13g2_decap_8 FILLER_19_1050 ();
 sg13g2_decap_8 FILLER_19_1057 ();
 sg13g2_decap_8 FILLER_19_1064 ();
 sg13g2_decap_8 FILLER_19_1071 ();
 sg13g2_decap_8 FILLER_19_1078 ();
 sg13g2_decap_8 FILLER_19_1085 ();
 sg13g2_decap_8 FILLER_19_1092 ();
 sg13g2_decap_8 FILLER_19_1099 ();
 sg13g2_decap_8 FILLER_19_1106 ();
 sg13g2_decap_8 FILLER_19_1113 ();
 sg13g2_decap_8 FILLER_19_1120 ();
 sg13g2_decap_8 FILLER_19_1127 ();
 sg13g2_decap_8 FILLER_19_1134 ();
 sg13g2_decap_8 FILLER_19_1141 ();
 sg13g2_decap_8 FILLER_19_1148 ();
 sg13g2_decap_8 FILLER_19_1155 ();
 sg13g2_decap_8 FILLER_19_1162 ();
 sg13g2_decap_8 FILLER_19_1169 ();
 sg13g2_decap_8 FILLER_19_1176 ();
 sg13g2_decap_8 FILLER_19_1183 ();
 sg13g2_decap_8 FILLER_19_1190 ();
 sg13g2_decap_8 FILLER_19_1197 ();
 sg13g2_decap_8 FILLER_19_1204 ();
 sg13g2_decap_8 FILLER_19_1211 ();
 sg13g2_decap_8 FILLER_19_1218 ();
 sg13g2_decap_8 FILLER_19_1225 ();
 sg13g2_decap_8 FILLER_19_1232 ();
 sg13g2_decap_8 FILLER_19_1239 ();
 sg13g2_decap_8 FILLER_19_1246 ();
 sg13g2_decap_8 FILLER_19_1253 ();
 sg13g2_decap_8 FILLER_19_1260 ();
 sg13g2_decap_8 FILLER_19_1267 ();
 sg13g2_decap_8 FILLER_19_1274 ();
 sg13g2_decap_8 FILLER_19_1281 ();
 sg13g2_decap_8 FILLER_19_1288 ();
 sg13g2_decap_8 FILLER_19_1295 ();
 sg13g2_decap_8 FILLER_19_1302 ();
 sg13g2_decap_8 FILLER_19_1309 ();
 sg13g2_decap_8 FILLER_19_1316 ();
 sg13g2_decap_8 FILLER_19_1323 ();
 sg13g2_decap_8 FILLER_19_1330 ();
 sg13g2_decap_8 FILLER_19_1337 ();
 sg13g2_decap_8 FILLER_19_1344 ();
 sg13g2_decap_8 FILLER_19_1351 ();
 sg13g2_decap_8 FILLER_19_1358 ();
 sg13g2_decap_8 FILLER_19_1365 ();
 sg13g2_decap_8 FILLER_19_1372 ();
 sg13g2_decap_8 FILLER_19_1379 ();
 sg13g2_decap_8 FILLER_19_1386 ();
 sg13g2_decap_8 FILLER_19_1393 ();
 sg13g2_decap_8 FILLER_19_1400 ();
 sg13g2_decap_8 FILLER_19_1407 ();
 sg13g2_decap_8 FILLER_19_1414 ();
 sg13g2_decap_8 FILLER_19_1421 ();
 sg13g2_decap_8 FILLER_19_1428 ();
 sg13g2_decap_8 FILLER_19_1435 ();
 sg13g2_decap_8 FILLER_19_1442 ();
 sg13g2_decap_8 FILLER_19_1449 ();
 sg13g2_decap_8 FILLER_19_1456 ();
 sg13g2_decap_8 FILLER_19_1463 ();
 sg13g2_decap_8 FILLER_19_1470 ();
 sg13g2_decap_8 FILLER_19_1477 ();
 sg13g2_decap_8 FILLER_19_1484 ();
 sg13g2_decap_8 FILLER_19_1491 ();
 sg13g2_decap_8 FILLER_19_1498 ();
 sg13g2_decap_8 FILLER_19_1505 ();
 sg13g2_decap_8 FILLER_19_1512 ();
 sg13g2_decap_8 FILLER_19_1519 ();
 sg13g2_decap_8 FILLER_19_1526 ();
 sg13g2_decap_8 FILLER_19_1533 ();
 sg13g2_decap_8 FILLER_19_1540 ();
 sg13g2_decap_8 FILLER_19_1547 ();
 sg13g2_decap_8 FILLER_19_1554 ();
 sg13g2_decap_8 FILLER_19_1561 ();
 sg13g2_decap_8 FILLER_19_1568 ();
 sg13g2_decap_8 FILLER_19_1575 ();
 sg13g2_decap_8 FILLER_19_1582 ();
 sg13g2_decap_8 FILLER_19_1589 ();
 sg13g2_decap_8 FILLER_19_1596 ();
 sg13g2_decap_8 FILLER_19_1603 ();
 sg13g2_decap_8 FILLER_19_1610 ();
 sg13g2_decap_8 FILLER_19_1617 ();
 sg13g2_decap_8 FILLER_19_1624 ();
 sg13g2_decap_8 FILLER_19_1631 ();
 sg13g2_decap_8 FILLER_19_1638 ();
 sg13g2_decap_8 FILLER_19_1645 ();
 sg13g2_decap_8 FILLER_19_1652 ();
 sg13g2_decap_8 FILLER_19_1659 ();
 sg13g2_decap_8 FILLER_19_1666 ();
 sg13g2_decap_8 FILLER_19_1673 ();
 sg13g2_decap_8 FILLER_19_1680 ();
 sg13g2_decap_8 FILLER_19_1687 ();
 sg13g2_decap_8 FILLER_19_1694 ();
 sg13g2_decap_8 FILLER_19_1701 ();
 sg13g2_decap_8 FILLER_19_1708 ();
 sg13g2_decap_8 FILLER_19_1715 ();
 sg13g2_decap_8 FILLER_19_1722 ();
 sg13g2_decap_8 FILLER_19_1729 ();
 sg13g2_decap_8 FILLER_19_1736 ();
 sg13g2_decap_8 FILLER_19_1743 ();
 sg13g2_decap_8 FILLER_19_1750 ();
 sg13g2_decap_8 FILLER_19_1757 ();
 sg13g2_decap_8 FILLER_19_1764 ();
 sg13g2_decap_8 FILLER_19_1771 ();
 sg13g2_decap_8 FILLER_19_1778 ();
 sg13g2_decap_8 FILLER_19_1785 ();
 sg13g2_decap_8 FILLER_19_1792 ();
 sg13g2_decap_8 FILLER_19_1799 ();
 sg13g2_decap_8 FILLER_19_1806 ();
 sg13g2_decap_8 FILLER_19_1813 ();
 sg13g2_decap_8 FILLER_19_1820 ();
 sg13g2_decap_8 FILLER_19_1827 ();
 sg13g2_decap_8 FILLER_19_1834 ();
 sg13g2_decap_8 FILLER_19_1841 ();
 sg13g2_decap_8 FILLER_19_1848 ();
 sg13g2_decap_8 FILLER_19_1855 ();
 sg13g2_decap_8 FILLER_19_1862 ();
 sg13g2_decap_8 FILLER_19_1869 ();
 sg13g2_decap_8 FILLER_19_1876 ();
 sg13g2_decap_8 FILLER_19_1883 ();
 sg13g2_decap_8 FILLER_19_1890 ();
 sg13g2_decap_8 FILLER_19_1897 ();
 sg13g2_decap_8 FILLER_19_1904 ();
 sg13g2_decap_8 FILLER_19_1911 ();
 sg13g2_decap_8 FILLER_19_1918 ();
 sg13g2_decap_8 FILLER_19_1925 ();
 sg13g2_decap_8 FILLER_19_1932 ();
 sg13g2_decap_8 FILLER_19_1939 ();
 sg13g2_decap_8 FILLER_19_1946 ();
 sg13g2_decap_8 FILLER_19_1953 ();
 sg13g2_decap_8 FILLER_19_1960 ();
 sg13g2_decap_8 FILLER_19_1967 ();
 sg13g2_decap_8 FILLER_19_1974 ();
 sg13g2_decap_8 FILLER_19_1981 ();
 sg13g2_decap_8 FILLER_19_1988 ();
 sg13g2_decap_8 FILLER_19_1995 ();
 sg13g2_decap_8 FILLER_19_2002 ();
 sg13g2_decap_8 FILLER_19_2009 ();
 sg13g2_decap_8 FILLER_19_2016 ();
 sg13g2_decap_8 FILLER_19_2023 ();
 sg13g2_decap_8 FILLER_19_2030 ();
 sg13g2_decap_8 FILLER_19_2037 ();
 sg13g2_decap_8 FILLER_19_2044 ();
 sg13g2_decap_8 FILLER_19_2051 ();
 sg13g2_decap_8 FILLER_19_2058 ();
 sg13g2_decap_8 FILLER_19_2065 ();
 sg13g2_decap_8 FILLER_19_2072 ();
 sg13g2_decap_8 FILLER_19_2079 ();
 sg13g2_decap_8 FILLER_19_2086 ();
 sg13g2_decap_8 FILLER_19_2093 ();
 sg13g2_decap_8 FILLER_19_2100 ();
 sg13g2_decap_8 FILLER_19_2107 ();
 sg13g2_decap_8 FILLER_19_2114 ();
 sg13g2_decap_8 FILLER_19_2121 ();
 sg13g2_decap_8 FILLER_19_2128 ();
 sg13g2_decap_8 FILLER_19_2135 ();
 sg13g2_decap_8 FILLER_19_2142 ();
 sg13g2_decap_8 FILLER_19_2149 ();
 sg13g2_decap_8 FILLER_19_2156 ();
 sg13g2_decap_8 FILLER_19_2163 ();
 sg13g2_decap_8 FILLER_19_2170 ();
 sg13g2_decap_8 FILLER_19_2177 ();
 sg13g2_decap_8 FILLER_19_2184 ();
 sg13g2_decap_8 FILLER_19_2191 ();
 sg13g2_decap_8 FILLER_19_2198 ();
 sg13g2_decap_8 FILLER_19_2205 ();
 sg13g2_decap_8 FILLER_19_2212 ();
 sg13g2_decap_8 FILLER_19_2219 ();
 sg13g2_decap_8 FILLER_19_2226 ();
 sg13g2_decap_8 FILLER_19_2233 ();
 sg13g2_decap_8 FILLER_19_2240 ();
 sg13g2_decap_8 FILLER_19_2247 ();
 sg13g2_decap_8 FILLER_19_2254 ();
 sg13g2_decap_8 FILLER_19_2261 ();
 sg13g2_decap_8 FILLER_19_2268 ();
 sg13g2_decap_8 FILLER_19_2275 ();
 sg13g2_decap_8 FILLER_19_2282 ();
 sg13g2_decap_8 FILLER_19_2289 ();
 sg13g2_decap_8 FILLER_19_2296 ();
 sg13g2_decap_8 FILLER_19_2303 ();
 sg13g2_decap_8 FILLER_19_2310 ();
 sg13g2_decap_8 FILLER_19_2317 ();
 sg13g2_decap_8 FILLER_19_2324 ();
 sg13g2_decap_8 FILLER_19_2331 ();
 sg13g2_decap_8 FILLER_19_2338 ();
 sg13g2_decap_8 FILLER_19_2345 ();
 sg13g2_decap_8 FILLER_19_2352 ();
 sg13g2_decap_8 FILLER_19_2359 ();
 sg13g2_decap_8 FILLER_19_2366 ();
 sg13g2_decap_8 FILLER_19_2373 ();
 sg13g2_decap_8 FILLER_19_2380 ();
 sg13g2_decap_8 FILLER_19_2387 ();
 sg13g2_decap_8 FILLER_19_2394 ();
 sg13g2_decap_8 FILLER_19_2401 ();
 sg13g2_decap_8 FILLER_19_2408 ();
 sg13g2_decap_8 FILLER_19_2415 ();
 sg13g2_decap_8 FILLER_19_2422 ();
 sg13g2_decap_8 FILLER_19_2429 ();
 sg13g2_decap_8 FILLER_19_2436 ();
 sg13g2_decap_8 FILLER_19_2443 ();
 sg13g2_decap_8 FILLER_19_2450 ();
 sg13g2_decap_8 FILLER_19_2457 ();
 sg13g2_decap_8 FILLER_19_2464 ();
 sg13g2_decap_8 FILLER_19_2471 ();
 sg13g2_decap_8 FILLER_19_2478 ();
 sg13g2_decap_8 FILLER_19_2485 ();
 sg13g2_decap_8 FILLER_19_2492 ();
 sg13g2_decap_8 FILLER_19_2499 ();
 sg13g2_decap_8 FILLER_19_2506 ();
 sg13g2_decap_8 FILLER_19_2513 ();
 sg13g2_decap_8 FILLER_19_2520 ();
 sg13g2_decap_8 FILLER_19_2527 ();
 sg13g2_decap_8 FILLER_19_2534 ();
 sg13g2_decap_8 FILLER_19_2541 ();
 sg13g2_decap_8 FILLER_19_2548 ();
 sg13g2_decap_8 FILLER_19_2555 ();
 sg13g2_decap_8 FILLER_19_2562 ();
 sg13g2_decap_8 FILLER_19_2569 ();
 sg13g2_decap_8 FILLER_19_2576 ();
 sg13g2_decap_8 FILLER_19_2583 ();
 sg13g2_decap_8 FILLER_19_2590 ();
 sg13g2_decap_8 FILLER_19_2597 ();
 sg13g2_decap_8 FILLER_19_2604 ();
 sg13g2_decap_8 FILLER_19_2611 ();
 sg13g2_decap_8 FILLER_19_2618 ();
 sg13g2_decap_8 FILLER_19_2625 ();
 sg13g2_decap_8 FILLER_19_2632 ();
 sg13g2_decap_8 FILLER_19_2639 ();
 sg13g2_decap_8 FILLER_19_2646 ();
 sg13g2_decap_8 FILLER_19_2653 ();
 sg13g2_decap_8 FILLER_19_2660 ();
 sg13g2_decap_8 FILLER_19_2667 ();
 sg13g2_decap_8 FILLER_19_2674 ();
 sg13g2_decap_8 FILLER_19_2681 ();
 sg13g2_decap_8 FILLER_19_2688 ();
 sg13g2_decap_8 FILLER_19_2695 ();
 sg13g2_decap_8 FILLER_19_2702 ();
 sg13g2_decap_8 FILLER_19_2709 ();
 sg13g2_decap_8 FILLER_19_2716 ();
 sg13g2_decap_8 FILLER_19_2723 ();
 sg13g2_decap_8 FILLER_19_2730 ();
 sg13g2_decap_8 FILLER_19_2737 ();
 sg13g2_decap_8 FILLER_19_2744 ();
 sg13g2_decap_8 FILLER_19_2751 ();
 sg13g2_decap_8 FILLER_19_2758 ();
 sg13g2_decap_8 FILLER_19_2765 ();
 sg13g2_decap_8 FILLER_19_2772 ();
 sg13g2_decap_8 FILLER_19_2779 ();
 sg13g2_decap_8 FILLER_19_2786 ();
 sg13g2_decap_8 FILLER_19_2793 ();
 sg13g2_decap_8 FILLER_19_2800 ();
 sg13g2_decap_8 FILLER_19_2807 ();
 sg13g2_decap_8 FILLER_19_2814 ();
 sg13g2_decap_8 FILLER_19_2821 ();
 sg13g2_decap_8 FILLER_19_2828 ();
 sg13g2_decap_8 FILLER_19_2835 ();
 sg13g2_decap_8 FILLER_19_2842 ();
 sg13g2_decap_8 FILLER_19_2849 ();
 sg13g2_decap_8 FILLER_19_2856 ();
 sg13g2_decap_8 FILLER_19_2863 ();
 sg13g2_decap_8 FILLER_19_2870 ();
 sg13g2_decap_8 FILLER_19_2877 ();
 sg13g2_decap_8 FILLER_19_2884 ();
 sg13g2_decap_8 FILLER_19_2891 ();
 sg13g2_decap_8 FILLER_19_2898 ();
 sg13g2_decap_8 FILLER_19_2905 ();
 sg13g2_decap_8 FILLER_19_2912 ();
 sg13g2_decap_8 FILLER_19_2919 ();
 sg13g2_decap_8 FILLER_19_2926 ();
 sg13g2_decap_8 FILLER_19_2933 ();
 sg13g2_decap_8 FILLER_19_2940 ();
 sg13g2_decap_8 FILLER_19_2947 ();
 sg13g2_decap_8 FILLER_19_2954 ();
 sg13g2_decap_8 FILLER_19_2961 ();
 sg13g2_decap_8 FILLER_19_2968 ();
 sg13g2_decap_8 FILLER_19_2975 ();
 sg13g2_decap_8 FILLER_19_2982 ();
 sg13g2_decap_8 FILLER_19_2989 ();
 sg13g2_decap_8 FILLER_19_2996 ();
 sg13g2_decap_8 FILLER_19_3003 ();
 sg13g2_decap_8 FILLER_19_3010 ();
 sg13g2_decap_8 FILLER_19_3017 ();
 sg13g2_decap_8 FILLER_19_3024 ();
 sg13g2_decap_8 FILLER_19_3031 ();
 sg13g2_decap_8 FILLER_19_3038 ();
 sg13g2_decap_8 FILLER_19_3045 ();
 sg13g2_decap_8 FILLER_19_3052 ();
 sg13g2_decap_8 FILLER_19_3059 ();
 sg13g2_decap_8 FILLER_19_3066 ();
 sg13g2_decap_8 FILLER_19_3073 ();
 sg13g2_decap_8 FILLER_19_3080 ();
 sg13g2_decap_8 FILLER_19_3087 ();
 sg13g2_decap_8 FILLER_19_3094 ();
 sg13g2_decap_8 FILLER_19_3101 ();
 sg13g2_decap_8 FILLER_19_3108 ();
 sg13g2_decap_8 FILLER_19_3115 ();
 sg13g2_decap_8 FILLER_19_3122 ();
 sg13g2_decap_8 FILLER_19_3129 ();
 sg13g2_decap_8 FILLER_19_3136 ();
 sg13g2_decap_8 FILLER_19_3143 ();
 sg13g2_decap_8 FILLER_19_3150 ();
 sg13g2_decap_8 FILLER_19_3157 ();
 sg13g2_decap_8 FILLER_19_3164 ();
 sg13g2_decap_8 FILLER_19_3171 ();
 sg13g2_decap_8 FILLER_19_3178 ();
 sg13g2_decap_8 FILLER_19_3185 ();
 sg13g2_decap_8 FILLER_19_3192 ();
 sg13g2_decap_8 FILLER_19_3199 ();
 sg13g2_decap_8 FILLER_19_3206 ();
 sg13g2_decap_8 FILLER_19_3213 ();
 sg13g2_decap_8 FILLER_19_3220 ();
 sg13g2_decap_8 FILLER_19_3227 ();
 sg13g2_decap_8 FILLER_19_3234 ();
 sg13g2_decap_8 FILLER_19_3241 ();
 sg13g2_decap_8 FILLER_19_3248 ();
 sg13g2_decap_8 FILLER_19_3255 ();
 sg13g2_decap_8 FILLER_19_3262 ();
 sg13g2_decap_8 FILLER_19_3269 ();
 sg13g2_decap_8 FILLER_19_3276 ();
 sg13g2_decap_8 FILLER_19_3283 ();
 sg13g2_decap_8 FILLER_19_3290 ();
 sg13g2_decap_8 FILLER_19_3297 ();
 sg13g2_decap_8 FILLER_19_3304 ();
 sg13g2_decap_8 FILLER_19_3311 ();
 sg13g2_decap_8 FILLER_19_3318 ();
 sg13g2_decap_8 FILLER_19_3325 ();
 sg13g2_decap_8 FILLER_19_3332 ();
 sg13g2_decap_8 FILLER_19_3339 ();
 sg13g2_decap_8 FILLER_19_3346 ();
 sg13g2_decap_8 FILLER_19_3353 ();
 sg13g2_decap_8 FILLER_19_3360 ();
 sg13g2_decap_8 FILLER_19_3367 ();
 sg13g2_decap_8 FILLER_19_3374 ();
 sg13g2_decap_8 FILLER_19_3381 ();
 sg13g2_decap_8 FILLER_19_3388 ();
 sg13g2_decap_8 FILLER_19_3395 ();
 sg13g2_decap_8 FILLER_19_3402 ();
 sg13g2_decap_8 FILLER_19_3409 ();
 sg13g2_decap_8 FILLER_19_3416 ();
 sg13g2_decap_8 FILLER_19_3423 ();
 sg13g2_decap_8 FILLER_19_3430 ();
 sg13g2_decap_8 FILLER_19_3437 ();
 sg13g2_decap_8 FILLER_19_3444 ();
 sg13g2_decap_8 FILLER_19_3451 ();
 sg13g2_decap_8 FILLER_19_3458 ();
 sg13g2_decap_8 FILLER_19_3465 ();
 sg13g2_decap_8 FILLER_19_3472 ();
 sg13g2_decap_8 FILLER_19_3479 ();
 sg13g2_decap_8 FILLER_19_3486 ();
 sg13g2_decap_8 FILLER_19_3493 ();
 sg13g2_decap_8 FILLER_19_3500 ();
 sg13g2_decap_8 FILLER_19_3507 ();
 sg13g2_decap_8 FILLER_19_3514 ();
 sg13g2_decap_8 FILLER_19_3521 ();
 sg13g2_decap_8 FILLER_19_3528 ();
 sg13g2_decap_8 FILLER_19_3535 ();
 sg13g2_decap_8 FILLER_19_3542 ();
 sg13g2_decap_8 FILLER_19_3549 ();
 sg13g2_decap_8 FILLER_19_3556 ();
 sg13g2_decap_8 FILLER_19_3563 ();
 sg13g2_decap_8 FILLER_19_3570 ();
 sg13g2_fill_2 FILLER_19_3577 ();
 sg13g2_fill_1 FILLER_19_3579 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_406 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_decap_8 FILLER_20_427 ();
 sg13g2_decap_8 FILLER_20_434 ();
 sg13g2_decap_8 FILLER_20_441 ();
 sg13g2_decap_8 FILLER_20_448 ();
 sg13g2_decap_8 FILLER_20_455 ();
 sg13g2_decap_8 FILLER_20_462 ();
 sg13g2_decap_8 FILLER_20_469 ();
 sg13g2_decap_8 FILLER_20_476 ();
 sg13g2_decap_8 FILLER_20_483 ();
 sg13g2_decap_8 FILLER_20_490 ();
 sg13g2_decap_8 FILLER_20_497 ();
 sg13g2_decap_8 FILLER_20_504 ();
 sg13g2_decap_8 FILLER_20_511 ();
 sg13g2_decap_8 FILLER_20_518 ();
 sg13g2_decap_8 FILLER_20_525 ();
 sg13g2_decap_8 FILLER_20_532 ();
 sg13g2_decap_8 FILLER_20_539 ();
 sg13g2_decap_8 FILLER_20_546 ();
 sg13g2_decap_8 FILLER_20_553 ();
 sg13g2_decap_8 FILLER_20_560 ();
 sg13g2_decap_8 FILLER_20_567 ();
 sg13g2_decap_8 FILLER_20_574 ();
 sg13g2_decap_8 FILLER_20_581 ();
 sg13g2_decap_8 FILLER_20_588 ();
 sg13g2_decap_8 FILLER_20_595 ();
 sg13g2_decap_8 FILLER_20_602 ();
 sg13g2_decap_8 FILLER_20_609 ();
 sg13g2_decap_8 FILLER_20_616 ();
 sg13g2_decap_8 FILLER_20_623 ();
 sg13g2_decap_8 FILLER_20_630 ();
 sg13g2_decap_8 FILLER_20_637 ();
 sg13g2_decap_8 FILLER_20_644 ();
 sg13g2_decap_8 FILLER_20_651 ();
 sg13g2_decap_8 FILLER_20_658 ();
 sg13g2_decap_8 FILLER_20_665 ();
 sg13g2_decap_8 FILLER_20_672 ();
 sg13g2_decap_8 FILLER_20_679 ();
 sg13g2_decap_8 FILLER_20_686 ();
 sg13g2_decap_8 FILLER_20_693 ();
 sg13g2_decap_8 FILLER_20_700 ();
 sg13g2_decap_8 FILLER_20_707 ();
 sg13g2_decap_8 FILLER_20_714 ();
 sg13g2_decap_8 FILLER_20_721 ();
 sg13g2_decap_8 FILLER_20_728 ();
 sg13g2_decap_8 FILLER_20_735 ();
 sg13g2_decap_8 FILLER_20_742 ();
 sg13g2_decap_8 FILLER_20_749 ();
 sg13g2_decap_8 FILLER_20_756 ();
 sg13g2_decap_8 FILLER_20_763 ();
 sg13g2_decap_8 FILLER_20_770 ();
 sg13g2_decap_8 FILLER_20_777 ();
 sg13g2_decap_8 FILLER_20_784 ();
 sg13g2_decap_8 FILLER_20_791 ();
 sg13g2_decap_8 FILLER_20_798 ();
 sg13g2_decap_8 FILLER_20_805 ();
 sg13g2_decap_8 FILLER_20_812 ();
 sg13g2_decap_8 FILLER_20_819 ();
 sg13g2_decap_8 FILLER_20_826 ();
 sg13g2_decap_8 FILLER_20_833 ();
 sg13g2_decap_8 FILLER_20_840 ();
 sg13g2_decap_8 FILLER_20_847 ();
 sg13g2_decap_8 FILLER_20_854 ();
 sg13g2_decap_8 FILLER_20_861 ();
 sg13g2_decap_8 FILLER_20_868 ();
 sg13g2_decap_8 FILLER_20_875 ();
 sg13g2_decap_8 FILLER_20_882 ();
 sg13g2_decap_8 FILLER_20_889 ();
 sg13g2_decap_8 FILLER_20_896 ();
 sg13g2_decap_8 FILLER_20_903 ();
 sg13g2_decap_8 FILLER_20_910 ();
 sg13g2_decap_8 FILLER_20_917 ();
 sg13g2_decap_8 FILLER_20_924 ();
 sg13g2_decap_8 FILLER_20_931 ();
 sg13g2_decap_8 FILLER_20_938 ();
 sg13g2_decap_8 FILLER_20_945 ();
 sg13g2_decap_8 FILLER_20_952 ();
 sg13g2_decap_8 FILLER_20_959 ();
 sg13g2_decap_8 FILLER_20_966 ();
 sg13g2_decap_8 FILLER_20_973 ();
 sg13g2_decap_8 FILLER_20_980 ();
 sg13g2_decap_8 FILLER_20_987 ();
 sg13g2_decap_8 FILLER_20_994 ();
 sg13g2_decap_8 FILLER_20_1001 ();
 sg13g2_decap_8 FILLER_20_1008 ();
 sg13g2_decap_8 FILLER_20_1015 ();
 sg13g2_decap_8 FILLER_20_1022 ();
 sg13g2_decap_8 FILLER_20_1029 ();
 sg13g2_decap_8 FILLER_20_1036 ();
 sg13g2_decap_8 FILLER_20_1043 ();
 sg13g2_decap_8 FILLER_20_1050 ();
 sg13g2_decap_8 FILLER_20_1057 ();
 sg13g2_decap_8 FILLER_20_1064 ();
 sg13g2_decap_8 FILLER_20_1071 ();
 sg13g2_decap_8 FILLER_20_1078 ();
 sg13g2_decap_8 FILLER_20_1085 ();
 sg13g2_decap_8 FILLER_20_1092 ();
 sg13g2_decap_8 FILLER_20_1099 ();
 sg13g2_decap_8 FILLER_20_1106 ();
 sg13g2_decap_8 FILLER_20_1113 ();
 sg13g2_decap_8 FILLER_20_1120 ();
 sg13g2_decap_8 FILLER_20_1127 ();
 sg13g2_decap_8 FILLER_20_1134 ();
 sg13g2_decap_8 FILLER_20_1141 ();
 sg13g2_decap_8 FILLER_20_1148 ();
 sg13g2_decap_8 FILLER_20_1155 ();
 sg13g2_decap_8 FILLER_20_1162 ();
 sg13g2_decap_8 FILLER_20_1169 ();
 sg13g2_decap_8 FILLER_20_1176 ();
 sg13g2_decap_8 FILLER_20_1183 ();
 sg13g2_decap_8 FILLER_20_1190 ();
 sg13g2_decap_8 FILLER_20_1197 ();
 sg13g2_decap_8 FILLER_20_1204 ();
 sg13g2_decap_8 FILLER_20_1211 ();
 sg13g2_decap_8 FILLER_20_1218 ();
 sg13g2_decap_8 FILLER_20_1225 ();
 sg13g2_decap_8 FILLER_20_1232 ();
 sg13g2_decap_8 FILLER_20_1239 ();
 sg13g2_decap_8 FILLER_20_1246 ();
 sg13g2_decap_8 FILLER_20_1253 ();
 sg13g2_decap_8 FILLER_20_1260 ();
 sg13g2_decap_8 FILLER_20_1267 ();
 sg13g2_decap_8 FILLER_20_1274 ();
 sg13g2_decap_8 FILLER_20_1281 ();
 sg13g2_decap_8 FILLER_20_1288 ();
 sg13g2_decap_8 FILLER_20_1295 ();
 sg13g2_decap_8 FILLER_20_1302 ();
 sg13g2_decap_8 FILLER_20_1309 ();
 sg13g2_decap_8 FILLER_20_1316 ();
 sg13g2_decap_8 FILLER_20_1323 ();
 sg13g2_decap_8 FILLER_20_1330 ();
 sg13g2_decap_8 FILLER_20_1337 ();
 sg13g2_decap_8 FILLER_20_1344 ();
 sg13g2_decap_8 FILLER_20_1351 ();
 sg13g2_decap_8 FILLER_20_1358 ();
 sg13g2_decap_8 FILLER_20_1365 ();
 sg13g2_decap_8 FILLER_20_1372 ();
 sg13g2_decap_8 FILLER_20_1379 ();
 sg13g2_decap_8 FILLER_20_1386 ();
 sg13g2_decap_8 FILLER_20_1393 ();
 sg13g2_decap_8 FILLER_20_1400 ();
 sg13g2_decap_8 FILLER_20_1407 ();
 sg13g2_decap_8 FILLER_20_1414 ();
 sg13g2_decap_8 FILLER_20_1421 ();
 sg13g2_decap_8 FILLER_20_1428 ();
 sg13g2_decap_8 FILLER_20_1435 ();
 sg13g2_decap_8 FILLER_20_1442 ();
 sg13g2_decap_8 FILLER_20_1449 ();
 sg13g2_decap_8 FILLER_20_1456 ();
 sg13g2_decap_8 FILLER_20_1463 ();
 sg13g2_decap_8 FILLER_20_1470 ();
 sg13g2_decap_8 FILLER_20_1477 ();
 sg13g2_decap_8 FILLER_20_1484 ();
 sg13g2_decap_8 FILLER_20_1491 ();
 sg13g2_decap_8 FILLER_20_1498 ();
 sg13g2_decap_8 FILLER_20_1505 ();
 sg13g2_decap_8 FILLER_20_1512 ();
 sg13g2_decap_8 FILLER_20_1519 ();
 sg13g2_decap_8 FILLER_20_1526 ();
 sg13g2_decap_8 FILLER_20_1533 ();
 sg13g2_decap_8 FILLER_20_1540 ();
 sg13g2_decap_8 FILLER_20_1547 ();
 sg13g2_decap_8 FILLER_20_1554 ();
 sg13g2_decap_8 FILLER_20_1561 ();
 sg13g2_decap_8 FILLER_20_1568 ();
 sg13g2_decap_8 FILLER_20_1575 ();
 sg13g2_decap_8 FILLER_20_1582 ();
 sg13g2_decap_8 FILLER_20_1589 ();
 sg13g2_decap_8 FILLER_20_1596 ();
 sg13g2_decap_8 FILLER_20_1603 ();
 sg13g2_decap_8 FILLER_20_1610 ();
 sg13g2_decap_8 FILLER_20_1617 ();
 sg13g2_decap_8 FILLER_20_1624 ();
 sg13g2_decap_8 FILLER_20_1631 ();
 sg13g2_decap_8 FILLER_20_1638 ();
 sg13g2_decap_8 FILLER_20_1645 ();
 sg13g2_decap_8 FILLER_20_1652 ();
 sg13g2_decap_8 FILLER_20_1659 ();
 sg13g2_decap_8 FILLER_20_1666 ();
 sg13g2_decap_8 FILLER_20_1673 ();
 sg13g2_decap_8 FILLER_20_1680 ();
 sg13g2_decap_8 FILLER_20_1687 ();
 sg13g2_decap_8 FILLER_20_1694 ();
 sg13g2_decap_8 FILLER_20_1701 ();
 sg13g2_decap_8 FILLER_20_1708 ();
 sg13g2_decap_8 FILLER_20_1715 ();
 sg13g2_decap_8 FILLER_20_1722 ();
 sg13g2_decap_8 FILLER_20_1729 ();
 sg13g2_decap_8 FILLER_20_1736 ();
 sg13g2_decap_8 FILLER_20_1743 ();
 sg13g2_decap_8 FILLER_20_1750 ();
 sg13g2_decap_8 FILLER_20_1757 ();
 sg13g2_decap_8 FILLER_20_1764 ();
 sg13g2_decap_8 FILLER_20_1771 ();
 sg13g2_decap_8 FILLER_20_1778 ();
 sg13g2_decap_8 FILLER_20_1785 ();
 sg13g2_decap_8 FILLER_20_1792 ();
 sg13g2_decap_8 FILLER_20_1799 ();
 sg13g2_decap_8 FILLER_20_1806 ();
 sg13g2_decap_8 FILLER_20_1813 ();
 sg13g2_decap_8 FILLER_20_1820 ();
 sg13g2_decap_8 FILLER_20_1827 ();
 sg13g2_decap_8 FILLER_20_1834 ();
 sg13g2_decap_8 FILLER_20_1841 ();
 sg13g2_decap_8 FILLER_20_1848 ();
 sg13g2_decap_8 FILLER_20_1855 ();
 sg13g2_decap_8 FILLER_20_1862 ();
 sg13g2_decap_8 FILLER_20_1869 ();
 sg13g2_decap_8 FILLER_20_1876 ();
 sg13g2_decap_8 FILLER_20_1883 ();
 sg13g2_decap_8 FILLER_20_1890 ();
 sg13g2_decap_8 FILLER_20_1897 ();
 sg13g2_decap_8 FILLER_20_1904 ();
 sg13g2_decap_8 FILLER_20_1911 ();
 sg13g2_decap_8 FILLER_20_1918 ();
 sg13g2_decap_8 FILLER_20_1925 ();
 sg13g2_decap_8 FILLER_20_1932 ();
 sg13g2_decap_8 FILLER_20_1939 ();
 sg13g2_decap_8 FILLER_20_1946 ();
 sg13g2_decap_8 FILLER_20_1953 ();
 sg13g2_decap_8 FILLER_20_1960 ();
 sg13g2_decap_8 FILLER_20_1967 ();
 sg13g2_decap_8 FILLER_20_1974 ();
 sg13g2_decap_8 FILLER_20_1981 ();
 sg13g2_decap_8 FILLER_20_1988 ();
 sg13g2_decap_8 FILLER_20_1995 ();
 sg13g2_decap_8 FILLER_20_2002 ();
 sg13g2_decap_8 FILLER_20_2009 ();
 sg13g2_decap_8 FILLER_20_2016 ();
 sg13g2_decap_8 FILLER_20_2023 ();
 sg13g2_decap_8 FILLER_20_2030 ();
 sg13g2_decap_8 FILLER_20_2037 ();
 sg13g2_decap_8 FILLER_20_2044 ();
 sg13g2_decap_8 FILLER_20_2051 ();
 sg13g2_decap_8 FILLER_20_2058 ();
 sg13g2_decap_8 FILLER_20_2065 ();
 sg13g2_decap_8 FILLER_20_2072 ();
 sg13g2_decap_8 FILLER_20_2079 ();
 sg13g2_decap_8 FILLER_20_2086 ();
 sg13g2_decap_8 FILLER_20_2093 ();
 sg13g2_decap_8 FILLER_20_2100 ();
 sg13g2_decap_8 FILLER_20_2107 ();
 sg13g2_decap_8 FILLER_20_2114 ();
 sg13g2_decap_8 FILLER_20_2121 ();
 sg13g2_decap_8 FILLER_20_2128 ();
 sg13g2_decap_8 FILLER_20_2135 ();
 sg13g2_decap_8 FILLER_20_2142 ();
 sg13g2_decap_8 FILLER_20_2149 ();
 sg13g2_decap_8 FILLER_20_2156 ();
 sg13g2_decap_8 FILLER_20_2163 ();
 sg13g2_decap_8 FILLER_20_2170 ();
 sg13g2_decap_8 FILLER_20_2177 ();
 sg13g2_decap_8 FILLER_20_2184 ();
 sg13g2_decap_8 FILLER_20_2191 ();
 sg13g2_decap_8 FILLER_20_2198 ();
 sg13g2_decap_8 FILLER_20_2205 ();
 sg13g2_decap_8 FILLER_20_2212 ();
 sg13g2_decap_8 FILLER_20_2219 ();
 sg13g2_decap_8 FILLER_20_2226 ();
 sg13g2_decap_8 FILLER_20_2233 ();
 sg13g2_decap_8 FILLER_20_2240 ();
 sg13g2_decap_8 FILLER_20_2247 ();
 sg13g2_decap_8 FILLER_20_2254 ();
 sg13g2_decap_8 FILLER_20_2261 ();
 sg13g2_decap_8 FILLER_20_2268 ();
 sg13g2_decap_8 FILLER_20_2275 ();
 sg13g2_decap_8 FILLER_20_2282 ();
 sg13g2_decap_8 FILLER_20_2289 ();
 sg13g2_decap_8 FILLER_20_2296 ();
 sg13g2_decap_8 FILLER_20_2303 ();
 sg13g2_decap_8 FILLER_20_2310 ();
 sg13g2_decap_8 FILLER_20_2317 ();
 sg13g2_decap_8 FILLER_20_2324 ();
 sg13g2_decap_8 FILLER_20_2331 ();
 sg13g2_decap_8 FILLER_20_2338 ();
 sg13g2_decap_8 FILLER_20_2345 ();
 sg13g2_decap_8 FILLER_20_2352 ();
 sg13g2_decap_8 FILLER_20_2359 ();
 sg13g2_decap_8 FILLER_20_2366 ();
 sg13g2_decap_8 FILLER_20_2373 ();
 sg13g2_decap_8 FILLER_20_2380 ();
 sg13g2_decap_8 FILLER_20_2387 ();
 sg13g2_decap_8 FILLER_20_2394 ();
 sg13g2_decap_8 FILLER_20_2401 ();
 sg13g2_decap_8 FILLER_20_2408 ();
 sg13g2_decap_8 FILLER_20_2415 ();
 sg13g2_decap_8 FILLER_20_2422 ();
 sg13g2_decap_8 FILLER_20_2429 ();
 sg13g2_decap_8 FILLER_20_2436 ();
 sg13g2_decap_8 FILLER_20_2443 ();
 sg13g2_decap_8 FILLER_20_2450 ();
 sg13g2_decap_8 FILLER_20_2457 ();
 sg13g2_decap_8 FILLER_20_2464 ();
 sg13g2_decap_8 FILLER_20_2471 ();
 sg13g2_decap_8 FILLER_20_2478 ();
 sg13g2_decap_8 FILLER_20_2485 ();
 sg13g2_decap_8 FILLER_20_2492 ();
 sg13g2_decap_8 FILLER_20_2499 ();
 sg13g2_decap_8 FILLER_20_2506 ();
 sg13g2_decap_8 FILLER_20_2513 ();
 sg13g2_decap_8 FILLER_20_2520 ();
 sg13g2_decap_8 FILLER_20_2527 ();
 sg13g2_decap_8 FILLER_20_2534 ();
 sg13g2_decap_8 FILLER_20_2541 ();
 sg13g2_decap_8 FILLER_20_2548 ();
 sg13g2_decap_8 FILLER_20_2555 ();
 sg13g2_decap_8 FILLER_20_2562 ();
 sg13g2_decap_8 FILLER_20_2569 ();
 sg13g2_decap_8 FILLER_20_2576 ();
 sg13g2_decap_8 FILLER_20_2583 ();
 sg13g2_decap_8 FILLER_20_2590 ();
 sg13g2_decap_8 FILLER_20_2597 ();
 sg13g2_decap_8 FILLER_20_2604 ();
 sg13g2_decap_8 FILLER_20_2611 ();
 sg13g2_decap_8 FILLER_20_2618 ();
 sg13g2_decap_8 FILLER_20_2625 ();
 sg13g2_decap_8 FILLER_20_2632 ();
 sg13g2_decap_8 FILLER_20_2639 ();
 sg13g2_decap_8 FILLER_20_2646 ();
 sg13g2_decap_8 FILLER_20_2653 ();
 sg13g2_decap_8 FILLER_20_2660 ();
 sg13g2_decap_8 FILLER_20_2667 ();
 sg13g2_decap_8 FILLER_20_2674 ();
 sg13g2_decap_8 FILLER_20_2681 ();
 sg13g2_decap_8 FILLER_20_2688 ();
 sg13g2_decap_8 FILLER_20_2695 ();
 sg13g2_decap_8 FILLER_20_2702 ();
 sg13g2_decap_8 FILLER_20_2709 ();
 sg13g2_decap_8 FILLER_20_2716 ();
 sg13g2_decap_8 FILLER_20_2723 ();
 sg13g2_decap_8 FILLER_20_2730 ();
 sg13g2_decap_8 FILLER_20_2737 ();
 sg13g2_decap_8 FILLER_20_2744 ();
 sg13g2_decap_8 FILLER_20_2751 ();
 sg13g2_decap_8 FILLER_20_2758 ();
 sg13g2_decap_8 FILLER_20_2765 ();
 sg13g2_decap_8 FILLER_20_2772 ();
 sg13g2_decap_8 FILLER_20_2779 ();
 sg13g2_decap_8 FILLER_20_2786 ();
 sg13g2_decap_8 FILLER_20_2793 ();
 sg13g2_decap_8 FILLER_20_2800 ();
 sg13g2_decap_8 FILLER_20_2807 ();
 sg13g2_decap_8 FILLER_20_2814 ();
 sg13g2_decap_8 FILLER_20_2821 ();
 sg13g2_decap_8 FILLER_20_2828 ();
 sg13g2_decap_8 FILLER_20_2835 ();
 sg13g2_decap_8 FILLER_20_2842 ();
 sg13g2_decap_8 FILLER_20_2849 ();
 sg13g2_decap_8 FILLER_20_2856 ();
 sg13g2_decap_8 FILLER_20_2863 ();
 sg13g2_decap_8 FILLER_20_2870 ();
 sg13g2_decap_8 FILLER_20_2877 ();
 sg13g2_decap_8 FILLER_20_2884 ();
 sg13g2_decap_8 FILLER_20_2891 ();
 sg13g2_decap_8 FILLER_20_2898 ();
 sg13g2_decap_8 FILLER_20_2905 ();
 sg13g2_decap_8 FILLER_20_2912 ();
 sg13g2_decap_8 FILLER_20_2919 ();
 sg13g2_decap_8 FILLER_20_2926 ();
 sg13g2_decap_8 FILLER_20_2933 ();
 sg13g2_decap_8 FILLER_20_2940 ();
 sg13g2_decap_8 FILLER_20_2947 ();
 sg13g2_decap_8 FILLER_20_2954 ();
 sg13g2_decap_8 FILLER_20_2961 ();
 sg13g2_decap_8 FILLER_20_2968 ();
 sg13g2_decap_8 FILLER_20_2975 ();
 sg13g2_decap_8 FILLER_20_2982 ();
 sg13g2_decap_8 FILLER_20_2989 ();
 sg13g2_decap_8 FILLER_20_2996 ();
 sg13g2_decap_8 FILLER_20_3003 ();
 sg13g2_decap_8 FILLER_20_3010 ();
 sg13g2_decap_8 FILLER_20_3017 ();
 sg13g2_decap_8 FILLER_20_3024 ();
 sg13g2_decap_8 FILLER_20_3031 ();
 sg13g2_decap_8 FILLER_20_3038 ();
 sg13g2_decap_8 FILLER_20_3045 ();
 sg13g2_decap_8 FILLER_20_3052 ();
 sg13g2_decap_8 FILLER_20_3059 ();
 sg13g2_decap_8 FILLER_20_3066 ();
 sg13g2_decap_8 FILLER_20_3073 ();
 sg13g2_decap_8 FILLER_20_3080 ();
 sg13g2_decap_8 FILLER_20_3087 ();
 sg13g2_decap_8 FILLER_20_3094 ();
 sg13g2_decap_8 FILLER_20_3101 ();
 sg13g2_decap_8 FILLER_20_3108 ();
 sg13g2_decap_8 FILLER_20_3115 ();
 sg13g2_decap_8 FILLER_20_3122 ();
 sg13g2_decap_8 FILLER_20_3129 ();
 sg13g2_decap_8 FILLER_20_3136 ();
 sg13g2_decap_8 FILLER_20_3143 ();
 sg13g2_decap_8 FILLER_20_3150 ();
 sg13g2_decap_8 FILLER_20_3157 ();
 sg13g2_decap_8 FILLER_20_3164 ();
 sg13g2_decap_8 FILLER_20_3171 ();
 sg13g2_decap_8 FILLER_20_3178 ();
 sg13g2_decap_8 FILLER_20_3185 ();
 sg13g2_decap_8 FILLER_20_3192 ();
 sg13g2_decap_8 FILLER_20_3199 ();
 sg13g2_decap_8 FILLER_20_3206 ();
 sg13g2_decap_8 FILLER_20_3213 ();
 sg13g2_decap_8 FILLER_20_3220 ();
 sg13g2_decap_8 FILLER_20_3227 ();
 sg13g2_decap_8 FILLER_20_3234 ();
 sg13g2_decap_8 FILLER_20_3241 ();
 sg13g2_decap_8 FILLER_20_3248 ();
 sg13g2_decap_8 FILLER_20_3255 ();
 sg13g2_decap_8 FILLER_20_3262 ();
 sg13g2_decap_8 FILLER_20_3269 ();
 sg13g2_decap_8 FILLER_20_3276 ();
 sg13g2_decap_8 FILLER_20_3283 ();
 sg13g2_decap_8 FILLER_20_3290 ();
 sg13g2_decap_8 FILLER_20_3297 ();
 sg13g2_decap_8 FILLER_20_3304 ();
 sg13g2_decap_8 FILLER_20_3311 ();
 sg13g2_decap_8 FILLER_20_3318 ();
 sg13g2_decap_8 FILLER_20_3325 ();
 sg13g2_decap_8 FILLER_20_3332 ();
 sg13g2_decap_8 FILLER_20_3339 ();
 sg13g2_decap_8 FILLER_20_3346 ();
 sg13g2_decap_8 FILLER_20_3353 ();
 sg13g2_decap_8 FILLER_20_3360 ();
 sg13g2_decap_8 FILLER_20_3367 ();
 sg13g2_decap_8 FILLER_20_3374 ();
 sg13g2_decap_8 FILLER_20_3381 ();
 sg13g2_decap_8 FILLER_20_3388 ();
 sg13g2_decap_8 FILLER_20_3395 ();
 sg13g2_decap_8 FILLER_20_3402 ();
 sg13g2_decap_8 FILLER_20_3409 ();
 sg13g2_decap_8 FILLER_20_3416 ();
 sg13g2_decap_8 FILLER_20_3423 ();
 sg13g2_decap_8 FILLER_20_3430 ();
 sg13g2_decap_8 FILLER_20_3437 ();
 sg13g2_decap_8 FILLER_20_3444 ();
 sg13g2_decap_8 FILLER_20_3451 ();
 sg13g2_decap_8 FILLER_20_3458 ();
 sg13g2_decap_8 FILLER_20_3465 ();
 sg13g2_decap_8 FILLER_20_3472 ();
 sg13g2_decap_8 FILLER_20_3479 ();
 sg13g2_decap_8 FILLER_20_3486 ();
 sg13g2_decap_8 FILLER_20_3493 ();
 sg13g2_decap_8 FILLER_20_3500 ();
 sg13g2_decap_8 FILLER_20_3507 ();
 sg13g2_decap_8 FILLER_20_3514 ();
 sg13g2_decap_8 FILLER_20_3521 ();
 sg13g2_decap_8 FILLER_20_3528 ();
 sg13g2_decap_8 FILLER_20_3535 ();
 sg13g2_decap_8 FILLER_20_3542 ();
 sg13g2_decap_8 FILLER_20_3549 ();
 sg13g2_decap_8 FILLER_20_3556 ();
 sg13g2_decap_8 FILLER_20_3563 ();
 sg13g2_decap_8 FILLER_20_3570 ();
 sg13g2_fill_2 FILLER_20_3577 ();
 sg13g2_fill_1 FILLER_20_3579 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_406 ();
 sg13g2_decap_8 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_420 ();
 sg13g2_decap_8 FILLER_21_427 ();
 sg13g2_decap_8 FILLER_21_434 ();
 sg13g2_decap_8 FILLER_21_441 ();
 sg13g2_decap_8 FILLER_21_448 ();
 sg13g2_decap_8 FILLER_21_455 ();
 sg13g2_decap_8 FILLER_21_462 ();
 sg13g2_decap_8 FILLER_21_469 ();
 sg13g2_decap_8 FILLER_21_476 ();
 sg13g2_decap_8 FILLER_21_483 ();
 sg13g2_decap_8 FILLER_21_490 ();
 sg13g2_decap_8 FILLER_21_497 ();
 sg13g2_decap_8 FILLER_21_504 ();
 sg13g2_decap_8 FILLER_21_511 ();
 sg13g2_decap_8 FILLER_21_518 ();
 sg13g2_decap_8 FILLER_21_525 ();
 sg13g2_decap_8 FILLER_21_532 ();
 sg13g2_decap_8 FILLER_21_539 ();
 sg13g2_decap_8 FILLER_21_546 ();
 sg13g2_decap_8 FILLER_21_553 ();
 sg13g2_decap_8 FILLER_21_560 ();
 sg13g2_decap_8 FILLER_21_567 ();
 sg13g2_decap_8 FILLER_21_574 ();
 sg13g2_decap_8 FILLER_21_581 ();
 sg13g2_decap_8 FILLER_21_588 ();
 sg13g2_decap_8 FILLER_21_595 ();
 sg13g2_decap_8 FILLER_21_602 ();
 sg13g2_decap_8 FILLER_21_609 ();
 sg13g2_decap_8 FILLER_21_616 ();
 sg13g2_decap_8 FILLER_21_623 ();
 sg13g2_decap_8 FILLER_21_630 ();
 sg13g2_decap_8 FILLER_21_637 ();
 sg13g2_decap_8 FILLER_21_644 ();
 sg13g2_decap_8 FILLER_21_651 ();
 sg13g2_decap_8 FILLER_21_658 ();
 sg13g2_decap_8 FILLER_21_665 ();
 sg13g2_decap_8 FILLER_21_672 ();
 sg13g2_decap_8 FILLER_21_679 ();
 sg13g2_decap_8 FILLER_21_686 ();
 sg13g2_decap_8 FILLER_21_693 ();
 sg13g2_decap_8 FILLER_21_700 ();
 sg13g2_decap_8 FILLER_21_707 ();
 sg13g2_decap_8 FILLER_21_714 ();
 sg13g2_decap_8 FILLER_21_721 ();
 sg13g2_decap_8 FILLER_21_728 ();
 sg13g2_decap_8 FILLER_21_735 ();
 sg13g2_decap_8 FILLER_21_742 ();
 sg13g2_decap_8 FILLER_21_749 ();
 sg13g2_decap_8 FILLER_21_756 ();
 sg13g2_decap_8 FILLER_21_763 ();
 sg13g2_decap_8 FILLER_21_770 ();
 sg13g2_decap_8 FILLER_21_777 ();
 sg13g2_decap_8 FILLER_21_784 ();
 sg13g2_decap_8 FILLER_21_791 ();
 sg13g2_decap_8 FILLER_21_798 ();
 sg13g2_decap_8 FILLER_21_805 ();
 sg13g2_decap_8 FILLER_21_812 ();
 sg13g2_decap_8 FILLER_21_819 ();
 sg13g2_decap_8 FILLER_21_826 ();
 sg13g2_decap_8 FILLER_21_833 ();
 sg13g2_decap_8 FILLER_21_840 ();
 sg13g2_decap_8 FILLER_21_847 ();
 sg13g2_decap_8 FILLER_21_854 ();
 sg13g2_decap_8 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_21_868 ();
 sg13g2_decap_8 FILLER_21_875 ();
 sg13g2_decap_8 FILLER_21_882 ();
 sg13g2_decap_8 FILLER_21_889 ();
 sg13g2_decap_8 FILLER_21_896 ();
 sg13g2_decap_8 FILLER_21_903 ();
 sg13g2_decap_8 FILLER_21_910 ();
 sg13g2_decap_8 FILLER_21_917 ();
 sg13g2_decap_8 FILLER_21_924 ();
 sg13g2_decap_8 FILLER_21_931 ();
 sg13g2_decap_8 FILLER_21_938 ();
 sg13g2_decap_8 FILLER_21_945 ();
 sg13g2_decap_8 FILLER_21_952 ();
 sg13g2_decap_8 FILLER_21_959 ();
 sg13g2_decap_8 FILLER_21_966 ();
 sg13g2_decap_8 FILLER_21_973 ();
 sg13g2_decap_8 FILLER_21_980 ();
 sg13g2_decap_8 FILLER_21_987 ();
 sg13g2_decap_8 FILLER_21_994 ();
 sg13g2_decap_8 FILLER_21_1001 ();
 sg13g2_decap_8 FILLER_21_1008 ();
 sg13g2_decap_8 FILLER_21_1015 ();
 sg13g2_decap_8 FILLER_21_1022 ();
 sg13g2_decap_8 FILLER_21_1029 ();
 sg13g2_decap_8 FILLER_21_1036 ();
 sg13g2_decap_8 FILLER_21_1043 ();
 sg13g2_decap_8 FILLER_21_1050 ();
 sg13g2_decap_8 FILLER_21_1057 ();
 sg13g2_decap_8 FILLER_21_1064 ();
 sg13g2_decap_8 FILLER_21_1071 ();
 sg13g2_decap_8 FILLER_21_1078 ();
 sg13g2_decap_8 FILLER_21_1085 ();
 sg13g2_decap_8 FILLER_21_1092 ();
 sg13g2_decap_8 FILLER_21_1099 ();
 sg13g2_decap_8 FILLER_21_1106 ();
 sg13g2_decap_8 FILLER_21_1113 ();
 sg13g2_decap_8 FILLER_21_1120 ();
 sg13g2_decap_8 FILLER_21_1127 ();
 sg13g2_decap_8 FILLER_21_1134 ();
 sg13g2_decap_8 FILLER_21_1141 ();
 sg13g2_decap_8 FILLER_21_1148 ();
 sg13g2_decap_8 FILLER_21_1155 ();
 sg13g2_decap_8 FILLER_21_1162 ();
 sg13g2_decap_8 FILLER_21_1169 ();
 sg13g2_decap_8 FILLER_21_1176 ();
 sg13g2_decap_8 FILLER_21_1183 ();
 sg13g2_decap_8 FILLER_21_1190 ();
 sg13g2_decap_8 FILLER_21_1197 ();
 sg13g2_decap_8 FILLER_21_1204 ();
 sg13g2_decap_8 FILLER_21_1211 ();
 sg13g2_decap_8 FILLER_21_1218 ();
 sg13g2_decap_8 FILLER_21_1225 ();
 sg13g2_decap_8 FILLER_21_1232 ();
 sg13g2_decap_8 FILLER_21_1239 ();
 sg13g2_decap_8 FILLER_21_1246 ();
 sg13g2_decap_8 FILLER_21_1253 ();
 sg13g2_decap_8 FILLER_21_1260 ();
 sg13g2_decap_8 FILLER_21_1267 ();
 sg13g2_decap_8 FILLER_21_1274 ();
 sg13g2_decap_8 FILLER_21_1281 ();
 sg13g2_decap_8 FILLER_21_1288 ();
 sg13g2_decap_8 FILLER_21_1295 ();
 sg13g2_decap_8 FILLER_21_1302 ();
 sg13g2_decap_8 FILLER_21_1309 ();
 sg13g2_decap_8 FILLER_21_1316 ();
 sg13g2_decap_8 FILLER_21_1323 ();
 sg13g2_decap_8 FILLER_21_1330 ();
 sg13g2_decap_8 FILLER_21_1337 ();
 sg13g2_decap_8 FILLER_21_1344 ();
 sg13g2_decap_8 FILLER_21_1351 ();
 sg13g2_decap_8 FILLER_21_1358 ();
 sg13g2_decap_8 FILLER_21_1365 ();
 sg13g2_decap_8 FILLER_21_1372 ();
 sg13g2_decap_8 FILLER_21_1379 ();
 sg13g2_decap_8 FILLER_21_1386 ();
 sg13g2_decap_8 FILLER_21_1393 ();
 sg13g2_decap_8 FILLER_21_1400 ();
 sg13g2_decap_8 FILLER_21_1407 ();
 sg13g2_decap_8 FILLER_21_1414 ();
 sg13g2_decap_8 FILLER_21_1421 ();
 sg13g2_decap_8 FILLER_21_1428 ();
 sg13g2_decap_8 FILLER_21_1435 ();
 sg13g2_decap_8 FILLER_21_1442 ();
 sg13g2_decap_8 FILLER_21_1449 ();
 sg13g2_decap_8 FILLER_21_1456 ();
 sg13g2_decap_8 FILLER_21_1463 ();
 sg13g2_decap_8 FILLER_21_1470 ();
 sg13g2_decap_8 FILLER_21_1477 ();
 sg13g2_decap_8 FILLER_21_1484 ();
 sg13g2_decap_8 FILLER_21_1491 ();
 sg13g2_decap_8 FILLER_21_1498 ();
 sg13g2_decap_8 FILLER_21_1505 ();
 sg13g2_decap_8 FILLER_21_1512 ();
 sg13g2_decap_8 FILLER_21_1519 ();
 sg13g2_decap_8 FILLER_21_1526 ();
 sg13g2_decap_8 FILLER_21_1533 ();
 sg13g2_decap_8 FILLER_21_1540 ();
 sg13g2_decap_8 FILLER_21_1547 ();
 sg13g2_decap_8 FILLER_21_1554 ();
 sg13g2_decap_8 FILLER_21_1561 ();
 sg13g2_decap_8 FILLER_21_1568 ();
 sg13g2_decap_8 FILLER_21_1575 ();
 sg13g2_decap_8 FILLER_21_1582 ();
 sg13g2_decap_8 FILLER_21_1589 ();
 sg13g2_decap_8 FILLER_21_1596 ();
 sg13g2_decap_8 FILLER_21_1603 ();
 sg13g2_decap_8 FILLER_21_1610 ();
 sg13g2_decap_8 FILLER_21_1617 ();
 sg13g2_decap_8 FILLER_21_1624 ();
 sg13g2_decap_8 FILLER_21_1631 ();
 sg13g2_decap_8 FILLER_21_1638 ();
 sg13g2_decap_8 FILLER_21_1645 ();
 sg13g2_decap_8 FILLER_21_1652 ();
 sg13g2_decap_8 FILLER_21_1659 ();
 sg13g2_decap_8 FILLER_21_1666 ();
 sg13g2_decap_8 FILLER_21_1673 ();
 sg13g2_decap_8 FILLER_21_1680 ();
 sg13g2_decap_8 FILLER_21_1687 ();
 sg13g2_decap_8 FILLER_21_1694 ();
 sg13g2_decap_8 FILLER_21_1701 ();
 sg13g2_decap_8 FILLER_21_1708 ();
 sg13g2_decap_8 FILLER_21_1715 ();
 sg13g2_decap_8 FILLER_21_1722 ();
 sg13g2_decap_8 FILLER_21_1729 ();
 sg13g2_decap_8 FILLER_21_1736 ();
 sg13g2_decap_8 FILLER_21_1743 ();
 sg13g2_decap_8 FILLER_21_1750 ();
 sg13g2_decap_8 FILLER_21_1757 ();
 sg13g2_decap_8 FILLER_21_1764 ();
 sg13g2_decap_8 FILLER_21_1771 ();
 sg13g2_decap_8 FILLER_21_1778 ();
 sg13g2_decap_8 FILLER_21_1785 ();
 sg13g2_decap_8 FILLER_21_1792 ();
 sg13g2_decap_8 FILLER_21_1799 ();
 sg13g2_decap_8 FILLER_21_1806 ();
 sg13g2_decap_8 FILLER_21_1813 ();
 sg13g2_decap_8 FILLER_21_1820 ();
 sg13g2_decap_8 FILLER_21_1827 ();
 sg13g2_decap_8 FILLER_21_1834 ();
 sg13g2_decap_8 FILLER_21_1841 ();
 sg13g2_decap_8 FILLER_21_1848 ();
 sg13g2_decap_8 FILLER_21_1855 ();
 sg13g2_decap_8 FILLER_21_1862 ();
 sg13g2_decap_8 FILLER_21_1869 ();
 sg13g2_decap_8 FILLER_21_1876 ();
 sg13g2_decap_8 FILLER_21_1883 ();
 sg13g2_decap_8 FILLER_21_1890 ();
 sg13g2_decap_8 FILLER_21_1897 ();
 sg13g2_decap_8 FILLER_21_1904 ();
 sg13g2_decap_8 FILLER_21_1911 ();
 sg13g2_decap_8 FILLER_21_1918 ();
 sg13g2_decap_8 FILLER_21_1925 ();
 sg13g2_decap_8 FILLER_21_1932 ();
 sg13g2_decap_8 FILLER_21_1939 ();
 sg13g2_decap_8 FILLER_21_1946 ();
 sg13g2_decap_8 FILLER_21_1953 ();
 sg13g2_decap_8 FILLER_21_1960 ();
 sg13g2_decap_8 FILLER_21_1967 ();
 sg13g2_decap_8 FILLER_21_1974 ();
 sg13g2_decap_8 FILLER_21_1981 ();
 sg13g2_decap_8 FILLER_21_1988 ();
 sg13g2_decap_8 FILLER_21_1995 ();
 sg13g2_decap_8 FILLER_21_2002 ();
 sg13g2_decap_8 FILLER_21_2009 ();
 sg13g2_decap_8 FILLER_21_2016 ();
 sg13g2_decap_8 FILLER_21_2023 ();
 sg13g2_decap_8 FILLER_21_2030 ();
 sg13g2_decap_8 FILLER_21_2037 ();
 sg13g2_decap_8 FILLER_21_2044 ();
 sg13g2_decap_8 FILLER_21_2051 ();
 sg13g2_decap_8 FILLER_21_2058 ();
 sg13g2_decap_8 FILLER_21_2065 ();
 sg13g2_decap_8 FILLER_21_2072 ();
 sg13g2_decap_8 FILLER_21_2079 ();
 sg13g2_decap_8 FILLER_21_2086 ();
 sg13g2_decap_8 FILLER_21_2093 ();
 sg13g2_decap_8 FILLER_21_2100 ();
 sg13g2_decap_8 FILLER_21_2107 ();
 sg13g2_decap_8 FILLER_21_2114 ();
 sg13g2_decap_8 FILLER_21_2121 ();
 sg13g2_decap_8 FILLER_21_2128 ();
 sg13g2_decap_8 FILLER_21_2135 ();
 sg13g2_decap_8 FILLER_21_2142 ();
 sg13g2_decap_8 FILLER_21_2149 ();
 sg13g2_decap_8 FILLER_21_2156 ();
 sg13g2_decap_8 FILLER_21_2163 ();
 sg13g2_decap_8 FILLER_21_2170 ();
 sg13g2_decap_8 FILLER_21_2177 ();
 sg13g2_decap_8 FILLER_21_2184 ();
 sg13g2_decap_8 FILLER_21_2191 ();
 sg13g2_decap_8 FILLER_21_2198 ();
 sg13g2_decap_8 FILLER_21_2205 ();
 sg13g2_decap_8 FILLER_21_2212 ();
 sg13g2_decap_8 FILLER_21_2219 ();
 sg13g2_decap_8 FILLER_21_2226 ();
 sg13g2_decap_8 FILLER_21_2233 ();
 sg13g2_decap_8 FILLER_21_2240 ();
 sg13g2_decap_8 FILLER_21_2247 ();
 sg13g2_decap_8 FILLER_21_2254 ();
 sg13g2_decap_8 FILLER_21_2261 ();
 sg13g2_decap_8 FILLER_21_2268 ();
 sg13g2_decap_8 FILLER_21_2275 ();
 sg13g2_decap_8 FILLER_21_2282 ();
 sg13g2_decap_8 FILLER_21_2289 ();
 sg13g2_decap_8 FILLER_21_2296 ();
 sg13g2_decap_8 FILLER_21_2303 ();
 sg13g2_decap_8 FILLER_21_2310 ();
 sg13g2_decap_8 FILLER_21_2317 ();
 sg13g2_decap_8 FILLER_21_2324 ();
 sg13g2_decap_8 FILLER_21_2331 ();
 sg13g2_decap_8 FILLER_21_2338 ();
 sg13g2_decap_8 FILLER_21_2345 ();
 sg13g2_decap_8 FILLER_21_2352 ();
 sg13g2_decap_8 FILLER_21_2359 ();
 sg13g2_decap_8 FILLER_21_2366 ();
 sg13g2_decap_8 FILLER_21_2373 ();
 sg13g2_decap_8 FILLER_21_2380 ();
 sg13g2_decap_8 FILLER_21_2387 ();
 sg13g2_decap_8 FILLER_21_2394 ();
 sg13g2_decap_8 FILLER_21_2401 ();
 sg13g2_decap_8 FILLER_21_2408 ();
 sg13g2_decap_8 FILLER_21_2415 ();
 sg13g2_decap_8 FILLER_21_2422 ();
 sg13g2_decap_8 FILLER_21_2429 ();
 sg13g2_decap_8 FILLER_21_2436 ();
 sg13g2_decap_8 FILLER_21_2443 ();
 sg13g2_decap_8 FILLER_21_2450 ();
 sg13g2_decap_8 FILLER_21_2457 ();
 sg13g2_decap_8 FILLER_21_2464 ();
 sg13g2_decap_8 FILLER_21_2471 ();
 sg13g2_decap_8 FILLER_21_2478 ();
 sg13g2_decap_8 FILLER_21_2485 ();
 sg13g2_decap_8 FILLER_21_2492 ();
 sg13g2_decap_8 FILLER_21_2499 ();
 sg13g2_decap_8 FILLER_21_2506 ();
 sg13g2_decap_8 FILLER_21_2513 ();
 sg13g2_decap_8 FILLER_21_2520 ();
 sg13g2_decap_8 FILLER_21_2527 ();
 sg13g2_decap_8 FILLER_21_2534 ();
 sg13g2_decap_8 FILLER_21_2541 ();
 sg13g2_decap_8 FILLER_21_2548 ();
 sg13g2_decap_8 FILLER_21_2555 ();
 sg13g2_decap_8 FILLER_21_2562 ();
 sg13g2_decap_8 FILLER_21_2569 ();
 sg13g2_decap_8 FILLER_21_2576 ();
 sg13g2_decap_8 FILLER_21_2583 ();
 sg13g2_decap_8 FILLER_21_2590 ();
 sg13g2_decap_8 FILLER_21_2597 ();
 sg13g2_decap_8 FILLER_21_2604 ();
 sg13g2_decap_8 FILLER_21_2611 ();
 sg13g2_decap_8 FILLER_21_2618 ();
 sg13g2_decap_8 FILLER_21_2625 ();
 sg13g2_decap_8 FILLER_21_2632 ();
 sg13g2_decap_8 FILLER_21_2639 ();
 sg13g2_decap_8 FILLER_21_2646 ();
 sg13g2_decap_8 FILLER_21_2653 ();
 sg13g2_decap_8 FILLER_21_2660 ();
 sg13g2_decap_8 FILLER_21_2667 ();
 sg13g2_decap_8 FILLER_21_2674 ();
 sg13g2_decap_8 FILLER_21_2681 ();
 sg13g2_decap_8 FILLER_21_2688 ();
 sg13g2_decap_8 FILLER_21_2695 ();
 sg13g2_decap_8 FILLER_21_2702 ();
 sg13g2_decap_8 FILLER_21_2709 ();
 sg13g2_decap_8 FILLER_21_2716 ();
 sg13g2_decap_8 FILLER_21_2723 ();
 sg13g2_decap_8 FILLER_21_2730 ();
 sg13g2_decap_8 FILLER_21_2737 ();
 sg13g2_decap_8 FILLER_21_2744 ();
 sg13g2_decap_8 FILLER_21_2751 ();
 sg13g2_decap_8 FILLER_21_2758 ();
 sg13g2_decap_8 FILLER_21_2765 ();
 sg13g2_decap_8 FILLER_21_2772 ();
 sg13g2_decap_8 FILLER_21_2779 ();
 sg13g2_decap_8 FILLER_21_2786 ();
 sg13g2_decap_8 FILLER_21_2793 ();
 sg13g2_decap_8 FILLER_21_2800 ();
 sg13g2_decap_8 FILLER_21_2807 ();
 sg13g2_decap_8 FILLER_21_2814 ();
 sg13g2_decap_8 FILLER_21_2821 ();
 sg13g2_decap_8 FILLER_21_2828 ();
 sg13g2_decap_8 FILLER_21_2835 ();
 sg13g2_decap_8 FILLER_21_2842 ();
 sg13g2_decap_8 FILLER_21_2849 ();
 sg13g2_decap_8 FILLER_21_2856 ();
 sg13g2_decap_8 FILLER_21_2863 ();
 sg13g2_decap_8 FILLER_21_2870 ();
 sg13g2_decap_8 FILLER_21_2877 ();
 sg13g2_decap_8 FILLER_21_2884 ();
 sg13g2_decap_8 FILLER_21_2891 ();
 sg13g2_decap_8 FILLER_21_2898 ();
 sg13g2_decap_8 FILLER_21_2905 ();
 sg13g2_decap_8 FILLER_21_2912 ();
 sg13g2_decap_8 FILLER_21_2919 ();
 sg13g2_decap_8 FILLER_21_2926 ();
 sg13g2_decap_8 FILLER_21_2933 ();
 sg13g2_decap_8 FILLER_21_2940 ();
 sg13g2_decap_8 FILLER_21_2947 ();
 sg13g2_decap_8 FILLER_21_2954 ();
 sg13g2_decap_8 FILLER_21_2961 ();
 sg13g2_decap_8 FILLER_21_2968 ();
 sg13g2_decap_8 FILLER_21_2975 ();
 sg13g2_decap_8 FILLER_21_2982 ();
 sg13g2_decap_8 FILLER_21_2989 ();
 sg13g2_decap_8 FILLER_21_2996 ();
 sg13g2_decap_8 FILLER_21_3003 ();
 sg13g2_decap_8 FILLER_21_3010 ();
 sg13g2_decap_8 FILLER_21_3017 ();
 sg13g2_decap_8 FILLER_21_3024 ();
 sg13g2_decap_8 FILLER_21_3031 ();
 sg13g2_decap_8 FILLER_21_3038 ();
 sg13g2_decap_8 FILLER_21_3045 ();
 sg13g2_decap_8 FILLER_21_3052 ();
 sg13g2_decap_8 FILLER_21_3059 ();
 sg13g2_decap_8 FILLER_21_3066 ();
 sg13g2_decap_8 FILLER_21_3073 ();
 sg13g2_decap_8 FILLER_21_3080 ();
 sg13g2_decap_8 FILLER_21_3087 ();
 sg13g2_decap_8 FILLER_21_3094 ();
 sg13g2_decap_8 FILLER_21_3101 ();
 sg13g2_decap_8 FILLER_21_3108 ();
 sg13g2_decap_8 FILLER_21_3115 ();
 sg13g2_decap_8 FILLER_21_3122 ();
 sg13g2_decap_8 FILLER_21_3129 ();
 sg13g2_decap_8 FILLER_21_3136 ();
 sg13g2_decap_8 FILLER_21_3143 ();
 sg13g2_decap_8 FILLER_21_3150 ();
 sg13g2_decap_8 FILLER_21_3157 ();
 sg13g2_decap_8 FILLER_21_3164 ();
 sg13g2_decap_8 FILLER_21_3171 ();
 sg13g2_decap_8 FILLER_21_3178 ();
 sg13g2_decap_8 FILLER_21_3185 ();
 sg13g2_decap_8 FILLER_21_3192 ();
 sg13g2_decap_8 FILLER_21_3199 ();
 sg13g2_decap_8 FILLER_21_3206 ();
 sg13g2_decap_8 FILLER_21_3213 ();
 sg13g2_decap_8 FILLER_21_3220 ();
 sg13g2_decap_8 FILLER_21_3227 ();
 sg13g2_decap_8 FILLER_21_3234 ();
 sg13g2_decap_8 FILLER_21_3241 ();
 sg13g2_decap_8 FILLER_21_3248 ();
 sg13g2_decap_8 FILLER_21_3255 ();
 sg13g2_decap_8 FILLER_21_3262 ();
 sg13g2_decap_8 FILLER_21_3269 ();
 sg13g2_decap_8 FILLER_21_3276 ();
 sg13g2_decap_8 FILLER_21_3283 ();
 sg13g2_decap_8 FILLER_21_3290 ();
 sg13g2_decap_8 FILLER_21_3297 ();
 sg13g2_decap_8 FILLER_21_3304 ();
 sg13g2_decap_8 FILLER_21_3311 ();
 sg13g2_decap_8 FILLER_21_3318 ();
 sg13g2_decap_8 FILLER_21_3325 ();
 sg13g2_decap_8 FILLER_21_3332 ();
 sg13g2_decap_8 FILLER_21_3339 ();
 sg13g2_decap_8 FILLER_21_3346 ();
 sg13g2_decap_8 FILLER_21_3353 ();
 sg13g2_decap_8 FILLER_21_3360 ();
 sg13g2_decap_8 FILLER_21_3367 ();
 sg13g2_decap_8 FILLER_21_3374 ();
 sg13g2_decap_8 FILLER_21_3381 ();
 sg13g2_decap_8 FILLER_21_3388 ();
 sg13g2_decap_8 FILLER_21_3395 ();
 sg13g2_decap_8 FILLER_21_3402 ();
 sg13g2_decap_8 FILLER_21_3409 ();
 sg13g2_decap_8 FILLER_21_3416 ();
 sg13g2_decap_8 FILLER_21_3423 ();
 sg13g2_decap_8 FILLER_21_3430 ();
 sg13g2_decap_8 FILLER_21_3437 ();
 sg13g2_decap_8 FILLER_21_3444 ();
 sg13g2_decap_8 FILLER_21_3451 ();
 sg13g2_decap_8 FILLER_21_3458 ();
 sg13g2_decap_8 FILLER_21_3465 ();
 sg13g2_decap_8 FILLER_21_3472 ();
 sg13g2_decap_8 FILLER_21_3479 ();
 sg13g2_decap_8 FILLER_21_3486 ();
 sg13g2_decap_8 FILLER_21_3493 ();
 sg13g2_decap_8 FILLER_21_3500 ();
 sg13g2_decap_8 FILLER_21_3507 ();
 sg13g2_decap_8 FILLER_21_3514 ();
 sg13g2_decap_8 FILLER_21_3521 ();
 sg13g2_decap_8 FILLER_21_3528 ();
 sg13g2_decap_8 FILLER_21_3535 ();
 sg13g2_decap_8 FILLER_21_3542 ();
 sg13g2_decap_8 FILLER_21_3549 ();
 sg13g2_decap_8 FILLER_21_3556 ();
 sg13g2_decap_8 FILLER_21_3563 ();
 sg13g2_decap_8 FILLER_21_3570 ();
 sg13g2_fill_2 FILLER_21_3577 ();
 sg13g2_fill_1 FILLER_21_3579 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_decap_8 FILLER_22_406 ();
 sg13g2_decap_8 FILLER_22_413 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_decap_8 FILLER_22_427 ();
 sg13g2_decap_8 FILLER_22_434 ();
 sg13g2_decap_8 FILLER_22_441 ();
 sg13g2_decap_8 FILLER_22_448 ();
 sg13g2_decap_8 FILLER_22_455 ();
 sg13g2_decap_8 FILLER_22_462 ();
 sg13g2_decap_8 FILLER_22_469 ();
 sg13g2_decap_8 FILLER_22_476 ();
 sg13g2_decap_8 FILLER_22_483 ();
 sg13g2_decap_8 FILLER_22_490 ();
 sg13g2_decap_8 FILLER_22_497 ();
 sg13g2_decap_8 FILLER_22_504 ();
 sg13g2_decap_8 FILLER_22_511 ();
 sg13g2_decap_8 FILLER_22_518 ();
 sg13g2_decap_8 FILLER_22_525 ();
 sg13g2_decap_8 FILLER_22_532 ();
 sg13g2_decap_8 FILLER_22_539 ();
 sg13g2_decap_8 FILLER_22_546 ();
 sg13g2_decap_8 FILLER_22_553 ();
 sg13g2_decap_8 FILLER_22_560 ();
 sg13g2_decap_8 FILLER_22_567 ();
 sg13g2_decap_8 FILLER_22_574 ();
 sg13g2_decap_8 FILLER_22_581 ();
 sg13g2_decap_8 FILLER_22_588 ();
 sg13g2_decap_8 FILLER_22_595 ();
 sg13g2_decap_8 FILLER_22_602 ();
 sg13g2_decap_8 FILLER_22_609 ();
 sg13g2_decap_8 FILLER_22_616 ();
 sg13g2_decap_8 FILLER_22_623 ();
 sg13g2_decap_8 FILLER_22_630 ();
 sg13g2_decap_8 FILLER_22_637 ();
 sg13g2_decap_8 FILLER_22_644 ();
 sg13g2_decap_8 FILLER_22_651 ();
 sg13g2_decap_8 FILLER_22_658 ();
 sg13g2_decap_8 FILLER_22_665 ();
 sg13g2_decap_8 FILLER_22_672 ();
 sg13g2_decap_8 FILLER_22_679 ();
 sg13g2_decap_8 FILLER_22_686 ();
 sg13g2_decap_8 FILLER_22_693 ();
 sg13g2_decap_8 FILLER_22_700 ();
 sg13g2_decap_8 FILLER_22_707 ();
 sg13g2_decap_8 FILLER_22_714 ();
 sg13g2_decap_8 FILLER_22_721 ();
 sg13g2_decap_8 FILLER_22_728 ();
 sg13g2_decap_8 FILLER_22_735 ();
 sg13g2_decap_8 FILLER_22_742 ();
 sg13g2_decap_8 FILLER_22_749 ();
 sg13g2_decap_8 FILLER_22_756 ();
 sg13g2_decap_8 FILLER_22_763 ();
 sg13g2_decap_8 FILLER_22_770 ();
 sg13g2_decap_8 FILLER_22_777 ();
 sg13g2_decap_8 FILLER_22_784 ();
 sg13g2_decap_8 FILLER_22_791 ();
 sg13g2_decap_8 FILLER_22_798 ();
 sg13g2_decap_8 FILLER_22_805 ();
 sg13g2_decap_8 FILLER_22_812 ();
 sg13g2_decap_8 FILLER_22_819 ();
 sg13g2_decap_8 FILLER_22_826 ();
 sg13g2_decap_8 FILLER_22_833 ();
 sg13g2_decap_8 FILLER_22_840 ();
 sg13g2_decap_8 FILLER_22_847 ();
 sg13g2_decap_8 FILLER_22_854 ();
 sg13g2_decap_8 FILLER_22_861 ();
 sg13g2_decap_8 FILLER_22_868 ();
 sg13g2_decap_8 FILLER_22_875 ();
 sg13g2_decap_8 FILLER_22_882 ();
 sg13g2_decap_8 FILLER_22_889 ();
 sg13g2_decap_8 FILLER_22_896 ();
 sg13g2_decap_8 FILLER_22_903 ();
 sg13g2_decap_8 FILLER_22_910 ();
 sg13g2_decap_8 FILLER_22_917 ();
 sg13g2_decap_8 FILLER_22_924 ();
 sg13g2_decap_8 FILLER_22_931 ();
 sg13g2_decap_8 FILLER_22_938 ();
 sg13g2_decap_8 FILLER_22_945 ();
 sg13g2_decap_8 FILLER_22_952 ();
 sg13g2_decap_8 FILLER_22_959 ();
 sg13g2_decap_8 FILLER_22_966 ();
 sg13g2_decap_8 FILLER_22_973 ();
 sg13g2_decap_8 FILLER_22_980 ();
 sg13g2_decap_8 FILLER_22_987 ();
 sg13g2_decap_8 FILLER_22_994 ();
 sg13g2_decap_8 FILLER_22_1001 ();
 sg13g2_decap_8 FILLER_22_1008 ();
 sg13g2_decap_8 FILLER_22_1015 ();
 sg13g2_decap_8 FILLER_22_1022 ();
 sg13g2_decap_8 FILLER_22_1029 ();
 sg13g2_decap_8 FILLER_22_1036 ();
 sg13g2_decap_8 FILLER_22_1043 ();
 sg13g2_decap_8 FILLER_22_1050 ();
 sg13g2_decap_8 FILLER_22_1057 ();
 sg13g2_decap_8 FILLER_22_1064 ();
 sg13g2_decap_8 FILLER_22_1071 ();
 sg13g2_decap_8 FILLER_22_1078 ();
 sg13g2_decap_8 FILLER_22_1085 ();
 sg13g2_decap_8 FILLER_22_1092 ();
 sg13g2_decap_8 FILLER_22_1099 ();
 sg13g2_decap_8 FILLER_22_1106 ();
 sg13g2_decap_8 FILLER_22_1113 ();
 sg13g2_decap_8 FILLER_22_1120 ();
 sg13g2_decap_8 FILLER_22_1127 ();
 sg13g2_decap_8 FILLER_22_1134 ();
 sg13g2_decap_8 FILLER_22_1141 ();
 sg13g2_decap_8 FILLER_22_1148 ();
 sg13g2_decap_8 FILLER_22_1155 ();
 sg13g2_decap_8 FILLER_22_1162 ();
 sg13g2_decap_8 FILLER_22_1169 ();
 sg13g2_decap_8 FILLER_22_1176 ();
 sg13g2_decap_8 FILLER_22_1183 ();
 sg13g2_decap_8 FILLER_22_1190 ();
 sg13g2_decap_8 FILLER_22_1197 ();
 sg13g2_decap_8 FILLER_22_1204 ();
 sg13g2_decap_8 FILLER_22_1211 ();
 sg13g2_decap_8 FILLER_22_1218 ();
 sg13g2_decap_8 FILLER_22_1225 ();
 sg13g2_decap_8 FILLER_22_1232 ();
 sg13g2_decap_8 FILLER_22_1239 ();
 sg13g2_decap_8 FILLER_22_1246 ();
 sg13g2_decap_8 FILLER_22_1253 ();
 sg13g2_decap_8 FILLER_22_1260 ();
 sg13g2_decap_8 FILLER_22_1267 ();
 sg13g2_decap_8 FILLER_22_1274 ();
 sg13g2_decap_8 FILLER_22_1281 ();
 sg13g2_decap_8 FILLER_22_1288 ();
 sg13g2_decap_8 FILLER_22_1295 ();
 sg13g2_decap_8 FILLER_22_1302 ();
 sg13g2_decap_8 FILLER_22_1309 ();
 sg13g2_decap_8 FILLER_22_1316 ();
 sg13g2_decap_8 FILLER_22_1323 ();
 sg13g2_decap_8 FILLER_22_1330 ();
 sg13g2_decap_8 FILLER_22_1337 ();
 sg13g2_decap_8 FILLER_22_1344 ();
 sg13g2_decap_8 FILLER_22_1351 ();
 sg13g2_decap_8 FILLER_22_1358 ();
 sg13g2_decap_8 FILLER_22_1365 ();
 sg13g2_decap_8 FILLER_22_1372 ();
 sg13g2_decap_8 FILLER_22_1379 ();
 sg13g2_decap_8 FILLER_22_1386 ();
 sg13g2_decap_8 FILLER_22_1393 ();
 sg13g2_decap_8 FILLER_22_1400 ();
 sg13g2_decap_8 FILLER_22_1407 ();
 sg13g2_decap_8 FILLER_22_1414 ();
 sg13g2_decap_8 FILLER_22_1421 ();
 sg13g2_decap_8 FILLER_22_1428 ();
 sg13g2_decap_8 FILLER_22_1435 ();
 sg13g2_decap_8 FILLER_22_1442 ();
 sg13g2_decap_8 FILLER_22_1449 ();
 sg13g2_decap_8 FILLER_22_1456 ();
 sg13g2_decap_8 FILLER_22_1463 ();
 sg13g2_decap_8 FILLER_22_1470 ();
 sg13g2_decap_8 FILLER_22_1477 ();
 sg13g2_decap_8 FILLER_22_1484 ();
 sg13g2_decap_8 FILLER_22_1491 ();
 sg13g2_decap_8 FILLER_22_1498 ();
 sg13g2_decap_8 FILLER_22_1505 ();
 sg13g2_decap_8 FILLER_22_1512 ();
 sg13g2_decap_8 FILLER_22_1519 ();
 sg13g2_decap_8 FILLER_22_1526 ();
 sg13g2_decap_8 FILLER_22_1533 ();
 sg13g2_decap_8 FILLER_22_1540 ();
 sg13g2_decap_8 FILLER_22_1547 ();
 sg13g2_decap_8 FILLER_22_1554 ();
 sg13g2_decap_8 FILLER_22_1561 ();
 sg13g2_decap_8 FILLER_22_1568 ();
 sg13g2_decap_8 FILLER_22_1575 ();
 sg13g2_decap_8 FILLER_22_1582 ();
 sg13g2_decap_8 FILLER_22_1589 ();
 sg13g2_decap_8 FILLER_22_1596 ();
 sg13g2_decap_8 FILLER_22_1603 ();
 sg13g2_decap_8 FILLER_22_1610 ();
 sg13g2_decap_8 FILLER_22_1617 ();
 sg13g2_decap_8 FILLER_22_1624 ();
 sg13g2_decap_8 FILLER_22_1631 ();
 sg13g2_decap_8 FILLER_22_1638 ();
 sg13g2_decap_8 FILLER_22_1645 ();
 sg13g2_decap_8 FILLER_22_1652 ();
 sg13g2_decap_8 FILLER_22_1659 ();
 sg13g2_decap_8 FILLER_22_1666 ();
 sg13g2_decap_8 FILLER_22_1673 ();
 sg13g2_decap_8 FILLER_22_1680 ();
 sg13g2_decap_8 FILLER_22_1687 ();
 sg13g2_decap_8 FILLER_22_1694 ();
 sg13g2_decap_8 FILLER_22_1701 ();
 sg13g2_decap_8 FILLER_22_1708 ();
 sg13g2_decap_8 FILLER_22_1715 ();
 sg13g2_decap_8 FILLER_22_1722 ();
 sg13g2_decap_8 FILLER_22_1729 ();
 sg13g2_decap_8 FILLER_22_1736 ();
 sg13g2_decap_8 FILLER_22_1743 ();
 sg13g2_decap_8 FILLER_22_1750 ();
 sg13g2_decap_8 FILLER_22_1757 ();
 sg13g2_decap_8 FILLER_22_1764 ();
 sg13g2_decap_8 FILLER_22_1771 ();
 sg13g2_decap_8 FILLER_22_1778 ();
 sg13g2_decap_8 FILLER_22_1785 ();
 sg13g2_decap_8 FILLER_22_1792 ();
 sg13g2_decap_8 FILLER_22_1799 ();
 sg13g2_decap_8 FILLER_22_1806 ();
 sg13g2_decap_8 FILLER_22_1813 ();
 sg13g2_decap_8 FILLER_22_1820 ();
 sg13g2_decap_8 FILLER_22_1827 ();
 sg13g2_decap_8 FILLER_22_1834 ();
 sg13g2_decap_8 FILLER_22_1841 ();
 sg13g2_decap_8 FILLER_22_1848 ();
 sg13g2_decap_8 FILLER_22_1855 ();
 sg13g2_decap_8 FILLER_22_1862 ();
 sg13g2_decap_8 FILLER_22_1869 ();
 sg13g2_decap_8 FILLER_22_1876 ();
 sg13g2_decap_8 FILLER_22_1883 ();
 sg13g2_decap_8 FILLER_22_1890 ();
 sg13g2_decap_8 FILLER_22_1897 ();
 sg13g2_decap_8 FILLER_22_1904 ();
 sg13g2_decap_8 FILLER_22_1911 ();
 sg13g2_decap_8 FILLER_22_1918 ();
 sg13g2_decap_8 FILLER_22_1925 ();
 sg13g2_decap_8 FILLER_22_1932 ();
 sg13g2_decap_8 FILLER_22_1939 ();
 sg13g2_decap_8 FILLER_22_1946 ();
 sg13g2_decap_8 FILLER_22_1953 ();
 sg13g2_decap_8 FILLER_22_1960 ();
 sg13g2_decap_8 FILLER_22_1967 ();
 sg13g2_decap_8 FILLER_22_1974 ();
 sg13g2_decap_8 FILLER_22_1981 ();
 sg13g2_decap_8 FILLER_22_1988 ();
 sg13g2_decap_8 FILLER_22_1995 ();
 sg13g2_decap_8 FILLER_22_2002 ();
 sg13g2_decap_8 FILLER_22_2009 ();
 sg13g2_decap_8 FILLER_22_2016 ();
 sg13g2_decap_8 FILLER_22_2023 ();
 sg13g2_decap_8 FILLER_22_2030 ();
 sg13g2_decap_8 FILLER_22_2037 ();
 sg13g2_decap_8 FILLER_22_2044 ();
 sg13g2_decap_8 FILLER_22_2051 ();
 sg13g2_decap_8 FILLER_22_2058 ();
 sg13g2_decap_8 FILLER_22_2065 ();
 sg13g2_decap_8 FILLER_22_2072 ();
 sg13g2_decap_8 FILLER_22_2079 ();
 sg13g2_decap_8 FILLER_22_2086 ();
 sg13g2_decap_8 FILLER_22_2093 ();
 sg13g2_decap_8 FILLER_22_2100 ();
 sg13g2_decap_8 FILLER_22_2107 ();
 sg13g2_decap_8 FILLER_22_2114 ();
 sg13g2_decap_8 FILLER_22_2121 ();
 sg13g2_decap_8 FILLER_22_2128 ();
 sg13g2_decap_8 FILLER_22_2135 ();
 sg13g2_decap_8 FILLER_22_2142 ();
 sg13g2_decap_8 FILLER_22_2149 ();
 sg13g2_decap_8 FILLER_22_2156 ();
 sg13g2_decap_8 FILLER_22_2163 ();
 sg13g2_decap_8 FILLER_22_2170 ();
 sg13g2_decap_8 FILLER_22_2177 ();
 sg13g2_decap_8 FILLER_22_2184 ();
 sg13g2_decap_8 FILLER_22_2191 ();
 sg13g2_decap_8 FILLER_22_2198 ();
 sg13g2_decap_8 FILLER_22_2205 ();
 sg13g2_decap_8 FILLER_22_2212 ();
 sg13g2_decap_8 FILLER_22_2219 ();
 sg13g2_decap_8 FILLER_22_2226 ();
 sg13g2_decap_8 FILLER_22_2233 ();
 sg13g2_decap_8 FILLER_22_2240 ();
 sg13g2_decap_8 FILLER_22_2247 ();
 sg13g2_decap_8 FILLER_22_2254 ();
 sg13g2_decap_8 FILLER_22_2261 ();
 sg13g2_decap_8 FILLER_22_2268 ();
 sg13g2_decap_8 FILLER_22_2275 ();
 sg13g2_decap_8 FILLER_22_2282 ();
 sg13g2_decap_8 FILLER_22_2289 ();
 sg13g2_decap_8 FILLER_22_2296 ();
 sg13g2_decap_8 FILLER_22_2303 ();
 sg13g2_decap_8 FILLER_22_2310 ();
 sg13g2_decap_8 FILLER_22_2317 ();
 sg13g2_decap_8 FILLER_22_2324 ();
 sg13g2_decap_8 FILLER_22_2331 ();
 sg13g2_decap_8 FILLER_22_2338 ();
 sg13g2_decap_8 FILLER_22_2345 ();
 sg13g2_decap_8 FILLER_22_2352 ();
 sg13g2_decap_8 FILLER_22_2359 ();
 sg13g2_decap_8 FILLER_22_2366 ();
 sg13g2_decap_8 FILLER_22_2373 ();
 sg13g2_decap_8 FILLER_22_2380 ();
 sg13g2_decap_8 FILLER_22_2387 ();
 sg13g2_decap_8 FILLER_22_2394 ();
 sg13g2_decap_8 FILLER_22_2401 ();
 sg13g2_decap_8 FILLER_22_2408 ();
 sg13g2_decap_8 FILLER_22_2415 ();
 sg13g2_decap_8 FILLER_22_2422 ();
 sg13g2_decap_8 FILLER_22_2429 ();
 sg13g2_decap_8 FILLER_22_2436 ();
 sg13g2_decap_8 FILLER_22_2443 ();
 sg13g2_decap_8 FILLER_22_2450 ();
 sg13g2_decap_8 FILLER_22_2457 ();
 sg13g2_decap_8 FILLER_22_2464 ();
 sg13g2_decap_8 FILLER_22_2471 ();
 sg13g2_decap_8 FILLER_22_2478 ();
 sg13g2_decap_8 FILLER_22_2485 ();
 sg13g2_decap_8 FILLER_22_2492 ();
 sg13g2_decap_8 FILLER_22_2499 ();
 sg13g2_decap_8 FILLER_22_2506 ();
 sg13g2_decap_8 FILLER_22_2513 ();
 sg13g2_decap_8 FILLER_22_2520 ();
 sg13g2_decap_8 FILLER_22_2527 ();
 sg13g2_decap_8 FILLER_22_2534 ();
 sg13g2_decap_8 FILLER_22_2541 ();
 sg13g2_decap_8 FILLER_22_2548 ();
 sg13g2_decap_8 FILLER_22_2555 ();
 sg13g2_decap_8 FILLER_22_2562 ();
 sg13g2_decap_8 FILLER_22_2569 ();
 sg13g2_decap_8 FILLER_22_2576 ();
 sg13g2_decap_8 FILLER_22_2583 ();
 sg13g2_decap_8 FILLER_22_2590 ();
 sg13g2_decap_8 FILLER_22_2597 ();
 sg13g2_decap_8 FILLER_22_2604 ();
 sg13g2_decap_8 FILLER_22_2611 ();
 sg13g2_decap_8 FILLER_22_2618 ();
 sg13g2_decap_8 FILLER_22_2625 ();
 sg13g2_decap_8 FILLER_22_2632 ();
 sg13g2_decap_8 FILLER_22_2639 ();
 sg13g2_decap_8 FILLER_22_2646 ();
 sg13g2_decap_8 FILLER_22_2653 ();
 sg13g2_decap_8 FILLER_22_2660 ();
 sg13g2_decap_8 FILLER_22_2667 ();
 sg13g2_decap_8 FILLER_22_2674 ();
 sg13g2_decap_8 FILLER_22_2681 ();
 sg13g2_decap_8 FILLER_22_2688 ();
 sg13g2_decap_8 FILLER_22_2695 ();
 sg13g2_decap_8 FILLER_22_2702 ();
 sg13g2_decap_8 FILLER_22_2709 ();
 sg13g2_decap_8 FILLER_22_2716 ();
 sg13g2_decap_8 FILLER_22_2723 ();
 sg13g2_decap_8 FILLER_22_2730 ();
 sg13g2_decap_8 FILLER_22_2737 ();
 sg13g2_decap_8 FILLER_22_2744 ();
 sg13g2_decap_8 FILLER_22_2751 ();
 sg13g2_decap_8 FILLER_22_2758 ();
 sg13g2_decap_8 FILLER_22_2765 ();
 sg13g2_decap_8 FILLER_22_2772 ();
 sg13g2_decap_8 FILLER_22_2779 ();
 sg13g2_decap_8 FILLER_22_2786 ();
 sg13g2_decap_8 FILLER_22_2793 ();
 sg13g2_decap_8 FILLER_22_2800 ();
 sg13g2_decap_8 FILLER_22_2807 ();
 sg13g2_decap_8 FILLER_22_2814 ();
 sg13g2_decap_8 FILLER_22_2821 ();
 sg13g2_decap_8 FILLER_22_2828 ();
 sg13g2_decap_8 FILLER_22_2835 ();
 sg13g2_decap_8 FILLER_22_2842 ();
 sg13g2_decap_8 FILLER_22_2849 ();
 sg13g2_decap_8 FILLER_22_2856 ();
 sg13g2_decap_8 FILLER_22_2863 ();
 sg13g2_decap_8 FILLER_22_2870 ();
 sg13g2_decap_8 FILLER_22_2877 ();
 sg13g2_decap_8 FILLER_22_2884 ();
 sg13g2_decap_8 FILLER_22_2891 ();
 sg13g2_decap_8 FILLER_22_2898 ();
 sg13g2_decap_8 FILLER_22_2905 ();
 sg13g2_decap_8 FILLER_22_2912 ();
 sg13g2_decap_8 FILLER_22_2919 ();
 sg13g2_decap_8 FILLER_22_2926 ();
 sg13g2_decap_8 FILLER_22_2933 ();
 sg13g2_decap_8 FILLER_22_2940 ();
 sg13g2_decap_8 FILLER_22_2947 ();
 sg13g2_decap_8 FILLER_22_2954 ();
 sg13g2_decap_8 FILLER_22_2961 ();
 sg13g2_decap_8 FILLER_22_2968 ();
 sg13g2_decap_8 FILLER_22_2975 ();
 sg13g2_decap_8 FILLER_22_2982 ();
 sg13g2_decap_8 FILLER_22_2989 ();
 sg13g2_decap_8 FILLER_22_2996 ();
 sg13g2_decap_8 FILLER_22_3003 ();
 sg13g2_decap_8 FILLER_22_3010 ();
 sg13g2_decap_8 FILLER_22_3017 ();
 sg13g2_decap_8 FILLER_22_3024 ();
 sg13g2_decap_8 FILLER_22_3031 ();
 sg13g2_decap_8 FILLER_22_3038 ();
 sg13g2_decap_8 FILLER_22_3045 ();
 sg13g2_decap_8 FILLER_22_3052 ();
 sg13g2_decap_8 FILLER_22_3059 ();
 sg13g2_decap_8 FILLER_22_3066 ();
 sg13g2_decap_8 FILLER_22_3073 ();
 sg13g2_decap_8 FILLER_22_3080 ();
 sg13g2_decap_8 FILLER_22_3087 ();
 sg13g2_decap_8 FILLER_22_3094 ();
 sg13g2_decap_8 FILLER_22_3101 ();
 sg13g2_decap_8 FILLER_22_3108 ();
 sg13g2_decap_8 FILLER_22_3115 ();
 sg13g2_decap_8 FILLER_22_3122 ();
 sg13g2_decap_8 FILLER_22_3129 ();
 sg13g2_decap_8 FILLER_22_3136 ();
 sg13g2_decap_8 FILLER_22_3143 ();
 sg13g2_decap_8 FILLER_22_3150 ();
 sg13g2_decap_8 FILLER_22_3157 ();
 sg13g2_decap_8 FILLER_22_3164 ();
 sg13g2_decap_8 FILLER_22_3171 ();
 sg13g2_decap_8 FILLER_22_3178 ();
 sg13g2_decap_8 FILLER_22_3185 ();
 sg13g2_decap_8 FILLER_22_3192 ();
 sg13g2_decap_8 FILLER_22_3199 ();
 sg13g2_decap_8 FILLER_22_3206 ();
 sg13g2_decap_8 FILLER_22_3213 ();
 sg13g2_decap_8 FILLER_22_3220 ();
 sg13g2_decap_8 FILLER_22_3227 ();
 sg13g2_decap_8 FILLER_22_3234 ();
 sg13g2_decap_8 FILLER_22_3241 ();
 sg13g2_decap_8 FILLER_22_3248 ();
 sg13g2_decap_8 FILLER_22_3255 ();
 sg13g2_decap_8 FILLER_22_3262 ();
 sg13g2_decap_8 FILLER_22_3269 ();
 sg13g2_decap_8 FILLER_22_3276 ();
 sg13g2_decap_8 FILLER_22_3283 ();
 sg13g2_decap_8 FILLER_22_3290 ();
 sg13g2_decap_8 FILLER_22_3297 ();
 sg13g2_decap_8 FILLER_22_3304 ();
 sg13g2_decap_8 FILLER_22_3311 ();
 sg13g2_decap_8 FILLER_22_3318 ();
 sg13g2_decap_8 FILLER_22_3325 ();
 sg13g2_decap_8 FILLER_22_3332 ();
 sg13g2_decap_8 FILLER_22_3339 ();
 sg13g2_decap_8 FILLER_22_3346 ();
 sg13g2_decap_8 FILLER_22_3353 ();
 sg13g2_decap_8 FILLER_22_3360 ();
 sg13g2_decap_8 FILLER_22_3367 ();
 sg13g2_decap_8 FILLER_22_3374 ();
 sg13g2_decap_8 FILLER_22_3381 ();
 sg13g2_decap_8 FILLER_22_3388 ();
 sg13g2_decap_8 FILLER_22_3395 ();
 sg13g2_decap_8 FILLER_22_3402 ();
 sg13g2_decap_8 FILLER_22_3409 ();
 sg13g2_decap_8 FILLER_22_3416 ();
 sg13g2_decap_8 FILLER_22_3423 ();
 sg13g2_decap_8 FILLER_22_3430 ();
 sg13g2_decap_8 FILLER_22_3437 ();
 sg13g2_decap_8 FILLER_22_3444 ();
 sg13g2_decap_8 FILLER_22_3451 ();
 sg13g2_decap_8 FILLER_22_3458 ();
 sg13g2_decap_8 FILLER_22_3465 ();
 sg13g2_decap_8 FILLER_22_3472 ();
 sg13g2_decap_8 FILLER_22_3479 ();
 sg13g2_decap_8 FILLER_22_3486 ();
 sg13g2_decap_8 FILLER_22_3493 ();
 sg13g2_decap_8 FILLER_22_3500 ();
 sg13g2_decap_8 FILLER_22_3507 ();
 sg13g2_decap_8 FILLER_22_3514 ();
 sg13g2_decap_8 FILLER_22_3521 ();
 sg13g2_decap_8 FILLER_22_3528 ();
 sg13g2_decap_8 FILLER_22_3535 ();
 sg13g2_decap_8 FILLER_22_3542 ();
 sg13g2_decap_8 FILLER_22_3549 ();
 sg13g2_decap_8 FILLER_22_3556 ();
 sg13g2_decap_8 FILLER_22_3563 ();
 sg13g2_decap_8 FILLER_22_3570 ();
 sg13g2_fill_2 FILLER_22_3577 ();
 sg13g2_fill_1 FILLER_22_3579 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_decap_8 FILLER_23_406 ();
 sg13g2_decap_8 FILLER_23_413 ();
 sg13g2_decap_8 FILLER_23_420 ();
 sg13g2_decap_8 FILLER_23_427 ();
 sg13g2_decap_8 FILLER_23_434 ();
 sg13g2_decap_8 FILLER_23_441 ();
 sg13g2_decap_8 FILLER_23_448 ();
 sg13g2_decap_8 FILLER_23_455 ();
 sg13g2_decap_8 FILLER_23_462 ();
 sg13g2_decap_8 FILLER_23_469 ();
 sg13g2_decap_8 FILLER_23_476 ();
 sg13g2_decap_8 FILLER_23_483 ();
 sg13g2_decap_8 FILLER_23_490 ();
 sg13g2_decap_8 FILLER_23_497 ();
 sg13g2_decap_8 FILLER_23_504 ();
 sg13g2_decap_8 FILLER_23_511 ();
 sg13g2_decap_8 FILLER_23_518 ();
 sg13g2_decap_8 FILLER_23_525 ();
 sg13g2_decap_8 FILLER_23_532 ();
 sg13g2_decap_8 FILLER_23_539 ();
 sg13g2_decap_8 FILLER_23_546 ();
 sg13g2_decap_8 FILLER_23_553 ();
 sg13g2_decap_8 FILLER_23_560 ();
 sg13g2_decap_8 FILLER_23_567 ();
 sg13g2_decap_8 FILLER_23_574 ();
 sg13g2_decap_8 FILLER_23_581 ();
 sg13g2_decap_8 FILLER_23_588 ();
 sg13g2_decap_8 FILLER_23_595 ();
 sg13g2_decap_8 FILLER_23_602 ();
 sg13g2_decap_8 FILLER_23_609 ();
 sg13g2_decap_8 FILLER_23_616 ();
 sg13g2_decap_8 FILLER_23_623 ();
 sg13g2_decap_8 FILLER_23_630 ();
 sg13g2_decap_8 FILLER_23_637 ();
 sg13g2_decap_8 FILLER_23_644 ();
 sg13g2_decap_8 FILLER_23_651 ();
 sg13g2_decap_8 FILLER_23_658 ();
 sg13g2_decap_8 FILLER_23_665 ();
 sg13g2_decap_8 FILLER_23_672 ();
 sg13g2_decap_8 FILLER_23_679 ();
 sg13g2_decap_8 FILLER_23_686 ();
 sg13g2_decap_8 FILLER_23_693 ();
 sg13g2_decap_8 FILLER_23_700 ();
 sg13g2_decap_8 FILLER_23_707 ();
 sg13g2_decap_8 FILLER_23_714 ();
 sg13g2_decap_8 FILLER_23_721 ();
 sg13g2_decap_8 FILLER_23_728 ();
 sg13g2_decap_8 FILLER_23_735 ();
 sg13g2_decap_8 FILLER_23_742 ();
 sg13g2_decap_8 FILLER_23_749 ();
 sg13g2_decap_8 FILLER_23_756 ();
 sg13g2_decap_8 FILLER_23_763 ();
 sg13g2_decap_8 FILLER_23_770 ();
 sg13g2_decap_8 FILLER_23_777 ();
 sg13g2_decap_8 FILLER_23_784 ();
 sg13g2_decap_8 FILLER_23_791 ();
 sg13g2_decap_8 FILLER_23_798 ();
 sg13g2_decap_8 FILLER_23_805 ();
 sg13g2_decap_8 FILLER_23_812 ();
 sg13g2_decap_8 FILLER_23_819 ();
 sg13g2_decap_8 FILLER_23_826 ();
 sg13g2_decap_8 FILLER_23_833 ();
 sg13g2_decap_8 FILLER_23_840 ();
 sg13g2_decap_8 FILLER_23_847 ();
 sg13g2_decap_8 FILLER_23_854 ();
 sg13g2_decap_8 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_23_868 ();
 sg13g2_decap_8 FILLER_23_875 ();
 sg13g2_decap_8 FILLER_23_882 ();
 sg13g2_decap_8 FILLER_23_889 ();
 sg13g2_decap_8 FILLER_23_896 ();
 sg13g2_decap_8 FILLER_23_903 ();
 sg13g2_decap_8 FILLER_23_910 ();
 sg13g2_decap_8 FILLER_23_917 ();
 sg13g2_decap_8 FILLER_23_924 ();
 sg13g2_decap_8 FILLER_23_931 ();
 sg13g2_decap_8 FILLER_23_938 ();
 sg13g2_decap_8 FILLER_23_945 ();
 sg13g2_decap_8 FILLER_23_952 ();
 sg13g2_decap_8 FILLER_23_959 ();
 sg13g2_decap_8 FILLER_23_966 ();
 sg13g2_decap_8 FILLER_23_973 ();
 sg13g2_decap_8 FILLER_23_980 ();
 sg13g2_decap_8 FILLER_23_987 ();
 sg13g2_decap_8 FILLER_23_994 ();
 sg13g2_decap_8 FILLER_23_1001 ();
 sg13g2_decap_8 FILLER_23_1008 ();
 sg13g2_decap_8 FILLER_23_1015 ();
 sg13g2_decap_8 FILLER_23_1022 ();
 sg13g2_decap_8 FILLER_23_1029 ();
 sg13g2_decap_8 FILLER_23_1036 ();
 sg13g2_decap_8 FILLER_23_1043 ();
 sg13g2_decap_8 FILLER_23_1050 ();
 sg13g2_decap_8 FILLER_23_1057 ();
 sg13g2_decap_8 FILLER_23_1064 ();
 sg13g2_decap_8 FILLER_23_1071 ();
 sg13g2_decap_8 FILLER_23_1078 ();
 sg13g2_decap_8 FILLER_23_1085 ();
 sg13g2_decap_8 FILLER_23_1092 ();
 sg13g2_decap_8 FILLER_23_1099 ();
 sg13g2_decap_8 FILLER_23_1106 ();
 sg13g2_decap_8 FILLER_23_1113 ();
 sg13g2_decap_8 FILLER_23_1120 ();
 sg13g2_decap_8 FILLER_23_1127 ();
 sg13g2_decap_8 FILLER_23_1134 ();
 sg13g2_decap_8 FILLER_23_1141 ();
 sg13g2_decap_8 FILLER_23_1148 ();
 sg13g2_decap_8 FILLER_23_1155 ();
 sg13g2_decap_8 FILLER_23_1162 ();
 sg13g2_decap_8 FILLER_23_1169 ();
 sg13g2_decap_8 FILLER_23_1176 ();
 sg13g2_decap_8 FILLER_23_1183 ();
 sg13g2_decap_8 FILLER_23_1190 ();
 sg13g2_decap_8 FILLER_23_1197 ();
 sg13g2_decap_8 FILLER_23_1204 ();
 sg13g2_decap_8 FILLER_23_1211 ();
 sg13g2_decap_8 FILLER_23_1218 ();
 sg13g2_decap_8 FILLER_23_1225 ();
 sg13g2_decap_8 FILLER_23_1232 ();
 sg13g2_decap_8 FILLER_23_1239 ();
 sg13g2_decap_8 FILLER_23_1246 ();
 sg13g2_decap_8 FILLER_23_1253 ();
 sg13g2_decap_8 FILLER_23_1260 ();
 sg13g2_decap_8 FILLER_23_1267 ();
 sg13g2_decap_8 FILLER_23_1274 ();
 sg13g2_decap_8 FILLER_23_1281 ();
 sg13g2_decap_8 FILLER_23_1288 ();
 sg13g2_decap_8 FILLER_23_1295 ();
 sg13g2_decap_8 FILLER_23_1302 ();
 sg13g2_decap_8 FILLER_23_1309 ();
 sg13g2_decap_8 FILLER_23_1316 ();
 sg13g2_decap_8 FILLER_23_1323 ();
 sg13g2_decap_8 FILLER_23_1330 ();
 sg13g2_decap_8 FILLER_23_1337 ();
 sg13g2_decap_8 FILLER_23_1344 ();
 sg13g2_decap_8 FILLER_23_1351 ();
 sg13g2_decap_8 FILLER_23_1358 ();
 sg13g2_decap_8 FILLER_23_1365 ();
 sg13g2_decap_8 FILLER_23_1372 ();
 sg13g2_decap_8 FILLER_23_1379 ();
 sg13g2_decap_8 FILLER_23_1386 ();
 sg13g2_decap_8 FILLER_23_1393 ();
 sg13g2_decap_8 FILLER_23_1400 ();
 sg13g2_decap_8 FILLER_23_1407 ();
 sg13g2_decap_8 FILLER_23_1414 ();
 sg13g2_decap_8 FILLER_23_1421 ();
 sg13g2_decap_8 FILLER_23_1428 ();
 sg13g2_decap_8 FILLER_23_1435 ();
 sg13g2_decap_8 FILLER_23_1442 ();
 sg13g2_decap_8 FILLER_23_1449 ();
 sg13g2_decap_8 FILLER_23_1456 ();
 sg13g2_decap_8 FILLER_23_1463 ();
 sg13g2_decap_8 FILLER_23_1470 ();
 sg13g2_decap_8 FILLER_23_1477 ();
 sg13g2_decap_8 FILLER_23_1484 ();
 sg13g2_decap_8 FILLER_23_1491 ();
 sg13g2_decap_8 FILLER_23_1498 ();
 sg13g2_decap_8 FILLER_23_1505 ();
 sg13g2_decap_8 FILLER_23_1512 ();
 sg13g2_decap_8 FILLER_23_1519 ();
 sg13g2_decap_8 FILLER_23_1526 ();
 sg13g2_decap_8 FILLER_23_1533 ();
 sg13g2_decap_8 FILLER_23_1540 ();
 sg13g2_decap_8 FILLER_23_1547 ();
 sg13g2_decap_8 FILLER_23_1554 ();
 sg13g2_decap_8 FILLER_23_1561 ();
 sg13g2_decap_8 FILLER_23_1568 ();
 sg13g2_decap_8 FILLER_23_1575 ();
 sg13g2_decap_8 FILLER_23_1582 ();
 sg13g2_decap_8 FILLER_23_1589 ();
 sg13g2_decap_8 FILLER_23_1596 ();
 sg13g2_decap_8 FILLER_23_1603 ();
 sg13g2_decap_8 FILLER_23_1610 ();
 sg13g2_decap_8 FILLER_23_1617 ();
 sg13g2_decap_8 FILLER_23_1624 ();
 sg13g2_decap_8 FILLER_23_1631 ();
 sg13g2_decap_8 FILLER_23_1638 ();
 sg13g2_decap_8 FILLER_23_1645 ();
 sg13g2_decap_8 FILLER_23_1652 ();
 sg13g2_decap_8 FILLER_23_1659 ();
 sg13g2_decap_8 FILLER_23_1666 ();
 sg13g2_decap_8 FILLER_23_1673 ();
 sg13g2_decap_8 FILLER_23_1680 ();
 sg13g2_decap_8 FILLER_23_1687 ();
 sg13g2_decap_8 FILLER_23_1694 ();
 sg13g2_decap_8 FILLER_23_1701 ();
 sg13g2_decap_8 FILLER_23_1708 ();
 sg13g2_decap_8 FILLER_23_1715 ();
 sg13g2_decap_8 FILLER_23_1722 ();
 sg13g2_decap_8 FILLER_23_1729 ();
 sg13g2_decap_8 FILLER_23_1736 ();
 sg13g2_decap_8 FILLER_23_1743 ();
 sg13g2_decap_8 FILLER_23_1750 ();
 sg13g2_decap_8 FILLER_23_1757 ();
 sg13g2_decap_8 FILLER_23_1764 ();
 sg13g2_decap_8 FILLER_23_1771 ();
 sg13g2_decap_8 FILLER_23_1778 ();
 sg13g2_decap_8 FILLER_23_1785 ();
 sg13g2_decap_8 FILLER_23_1792 ();
 sg13g2_decap_8 FILLER_23_1799 ();
 sg13g2_decap_8 FILLER_23_1806 ();
 sg13g2_decap_8 FILLER_23_1813 ();
 sg13g2_decap_8 FILLER_23_1820 ();
 sg13g2_decap_8 FILLER_23_1827 ();
 sg13g2_decap_8 FILLER_23_1834 ();
 sg13g2_decap_8 FILLER_23_1841 ();
 sg13g2_decap_8 FILLER_23_1848 ();
 sg13g2_decap_8 FILLER_23_1855 ();
 sg13g2_decap_8 FILLER_23_1862 ();
 sg13g2_decap_8 FILLER_23_1869 ();
 sg13g2_decap_8 FILLER_23_1876 ();
 sg13g2_decap_8 FILLER_23_1883 ();
 sg13g2_decap_8 FILLER_23_1890 ();
 sg13g2_decap_8 FILLER_23_1897 ();
 sg13g2_decap_8 FILLER_23_1904 ();
 sg13g2_decap_8 FILLER_23_1911 ();
 sg13g2_decap_8 FILLER_23_1918 ();
 sg13g2_decap_8 FILLER_23_1925 ();
 sg13g2_decap_8 FILLER_23_1932 ();
 sg13g2_decap_8 FILLER_23_1939 ();
 sg13g2_decap_8 FILLER_23_1946 ();
 sg13g2_decap_8 FILLER_23_1953 ();
 sg13g2_decap_8 FILLER_23_1960 ();
 sg13g2_decap_8 FILLER_23_1967 ();
 sg13g2_decap_8 FILLER_23_1974 ();
 sg13g2_decap_8 FILLER_23_1981 ();
 sg13g2_decap_8 FILLER_23_1988 ();
 sg13g2_decap_8 FILLER_23_1995 ();
 sg13g2_decap_8 FILLER_23_2002 ();
 sg13g2_decap_8 FILLER_23_2009 ();
 sg13g2_decap_8 FILLER_23_2016 ();
 sg13g2_decap_8 FILLER_23_2023 ();
 sg13g2_decap_8 FILLER_23_2030 ();
 sg13g2_decap_8 FILLER_23_2037 ();
 sg13g2_decap_8 FILLER_23_2044 ();
 sg13g2_decap_8 FILLER_23_2051 ();
 sg13g2_decap_8 FILLER_23_2058 ();
 sg13g2_decap_8 FILLER_23_2065 ();
 sg13g2_decap_8 FILLER_23_2072 ();
 sg13g2_decap_8 FILLER_23_2079 ();
 sg13g2_decap_8 FILLER_23_2086 ();
 sg13g2_decap_8 FILLER_23_2093 ();
 sg13g2_decap_8 FILLER_23_2100 ();
 sg13g2_decap_8 FILLER_23_2107 ();
 sg13g2_decap_8 FILLER_23_2114 ();
 sg13g2_decap_8 FILLER_23_2121 ();
 sg13g2_decap_8 FILLER_23_2128 ();
 sg13g2_decap_8 FILLER_23_2135 ();
 sg13g2_decap_8 FILLER_23_2142 ();
 sg13g2_decap_8 FILLER_23_2149 ();
 sg13g2_decap_8 FILLER_23_2156 ();
 sg13g2_decap_8 FILLER_23_2163 ();
 sg13g2_decap_8 FILLER_23_2170 ();
 sg13g2_decap_8 FILLER_23_2177 ();
 sg13g2_decap_8 FILLER_23_2184 ();
 sg13g2_decap_8 FILLER_23_2191 ();
 sg13g2_decap_8 FILLER_23_2198 ();
 sg13g2_decap_8 FILLER_23_2205 ();
 sg13g2_decap_8 FILLER_23_2212 ();
 sg13g2_decap_8 FILLER_23_2219 ();
 sg13g2_decap_8 FILLER_23_2226 ();
 sg13g2_decap_8 FILLER_23_2233 ();
 sg13g2_decap_8 FILLER_23_2240 ();
 sg13g2_decap_8 FILLER_23_2247 ();
 sg13g2_decap_8 FILLER_23_2254 ();
 sg13g2_decap_8 FILLER_23_2261 ();
 sg13g2_decap_8 FILLER_23_2268 ();
 sg13g2_decap_8 FILLER_23_2275 ();
 sg13g2_decap_8 FILLER_23_2282 ();
 sg13g2_decap_8 FILLER_23_2289 ();
 sg13g2_decap_8 FILLER_23_2296 ();
 sg13g2_decap_8 FILLER_23_2303 ();
 sg13g2_decap_8 FILLER_23_2310 ();
 sg13g2_decap_8 FILLER_23_2317 ();
 sg13g2_decap_8 FILLER_23_2324 ();
 sg13g2_decap_8 FILLER_23_2331 ();
 sg13g2_decap_8 FILLER_23_2338 ();
 sg13g2_decap_8 FILLER_23_2345 ();
 sg13g2_decap_8 FILLER_23_2352 ();
 sg13g2_decap_8 FILLER_23_2359 ();
 sg13g2_decap_8 FILLER_23_2366 ();
 sg13g2_decap_8 FILLER_23_2373 ();
 sg13g2_decap_8 FILLER_23_2380 ();
 sg13g2_decap_8 FILLER_23_2387 ();
 sg13g2_decap_8 FILLER_23_2394 ();
 sg13g2_decap_8 FILLER_23_2401 ();
 sg13g2_decap_8 FILLER_23_2408 ();
 sg13g2_decap_8 FILLER_23_2415 ();
 sg13g2_decap_8 FILLER_23_2422 ();
 sg13g2_decap_8 FILLER_23_2429 ();
 sg13g2_decap_8 FILLER_23_2436 ();
 sg13g2_decap_8 FILLER_23_2443 ();
 sg13g2_decap_8 FILLER_23_2450 ();
 sg13g2_decap_8 FILLER_23_2457 ();
 sg13g2_decap_8 FILLER_23_2464 ();
 sg13g2_decap_8 FILLER_23_2471 ();
 sg13g2_decap_8 FILLER_23_2478 ();
 sg13g2_decap_8 FILLER_23_2485 ();
 sg13g2_decap_8 FILLER_23_2492 ();
 sg13g2_decap_8 FILLER_23_2499 ();
 sg13g2_decap_8 FILLER_23_2506 ();
 sg13g2_decap_8 FILLER_23_2513 ();
 sg13g2_decap_8 FILLER_23_2520 ();
 sg13g2_decap_8 FILLER_23_2527 ();
 sg13g2_decap_8 FILLER_23_2534 ();
 sg13g2_decap_8 FILLER_23_2541 ();
 sg13g2_decap_8 FILLER_23_2548 ();
 sg13g2_decap_8 FILLER_23_2555 ();
 sg13g2_decap_8 FILLER_23_2562 ();
 sg13g2_decap_8 FILLER_23_2569 ();
 sg13g2_decap_8 FILLER_23_2576 ();
 sg13g2_decap_8 FILLER_23_2583 ();
 sg13g2_decap_8 FILLER_23_2590 ();
 sg13g2_decap_8 FILLER_23_2597 ();
 sg13g2_decap_8 FILLER_23_2604 ();
 sg13g2_decap_8 FILLER_23_2611 ();
 sg13g2_decap_8 FILLER_23_2618 ();
 sg13g2_decap_8 FILLER_23_2625 ();
 sg13g2_decap_8 FILLER_23_2632 ();
 sg13g2_decap_8 FILLER_23_2639 ();
 sg13g2_decap_8 FILLER_23_2646 ();
 sg13g2_decap_8 FILLER_23_2653 ();
 sg13g2_decap_8 FILLER_23_2660 ();
 sg13g2_decap_8 FILLER_23_2667 ();
 sg13g2_decap_8 FILLER_23_2674 ();
 sg13g2_decap_8 FILLER_23_2681 ();
 sg13g2_decap_8 FILLER_23_2688 ();
 sg13g2_decap_8 FILLER_23_2695 ();
 sg13g2_decap_8 FILLER_23_2702 ();
 sg13g2_decap_8 FILLER_23_2709 ();
 sg13g2_decap_8 FILLER_23_2716 ();
 sg13g2_decap_8 FILLER_23_2723 ();
 sg13g2_decap_8 FILLER_23_2730 ();
 sg13g2_decap_8 FILLER_23_2737 ();
 sg13g2_decap_8 FILLER_23_2744 ();
 sg13g2_decap_8 FILLER_23_2751 ();
 sg13g2_decap_8 FILLER_23_2758 ();
 sg13g2_decap_8 FILLER_23_2765 ();
 sg13g2_decap_8 FILLER_23_2772 ();
 sg13g2_decap_8 FILLER_23_2779 ();
 sg13g2_decap_8 FILLER_23_2786 ();
 sg13g2_decap_8 FILLER_23_2793 ();
 sg13g2_decap_8 FILLER_23_2800 ();
 sg13g2_decap_8 FILLER_23_2807 ();
 sg13g2_decap_8 FILLER_23_2814 ();
 sg13g2_decap_8 FILLER_23_2821 ();
 sg13g2_decap_8 FILLER_23_2828 ();
 sg13g2_decap_8 FILLER_23_2835 ();
 sg13g2_decap_8 FILLER_23_2842 ();
 sg13g2_decap_8 FILLER_23_2849 ();
 sg13g2_decap_8 FILLER_23_2856 ();
 sg13g2_decap_8 FILLER_23_2863 ();
 sg13g2_decap_8 FILLER_23_2870 ();
 sg13g2_decap_8 FILLER_23_2877 ();
 sg13g2_decap_8 FILLER_23_2884 ();
 sg13g2_decap_8 FILLER_23_2891 ();
 sg13g2_decap_8 FILLER_23_2898 ();
 sg13g2_decap_8 FILLER_23_2905 ();
 sg13g2_decap_8 FILLER_23_2912 ();
 sg13g2_decap_8 FILLER_23_2919 ();
 sg13g2_decap_8 FILLER_23_2926 ();
 sg13g2_decap_8 FILLER_23_2933 ();
 sg13g2_decap_8 FILLER_23_2940 ();
 sg13g2_decap_8 FILLER_23_2947 ();
 sg13g2_decap_8 FILLER_23_2954 ();
 sg13g2_decap_8 FILLER_23_2961 ();
 sg13g2_decap_8 FILLER_23_2968 ();
 sg13g2_decap_8 FILLER_23_2975 ();
 sg13g2_decap_8 FILLER_23_2982 ();
 sg13g2_decap_8 FILLER_23_2989 ();
 sg13g2_decap_8 FILLER_23_2996 ();
 sg13g2_decap_8 FILLER_23_3003 ();
 sg13g2_decap_8 FILLER_23_3010 ();
 sg13g2_decap_8 FILLER_23_3017 ();
 sg13g2_decap_8 FILLER_23_3024 ();
 sg13g2_decap_8 FILLER_23_3031 ();
 sg13g2_decap_8 FILLER_23_3038 ();
 sg13g2_decap_8 FILLER_23_3045 ();
 sg13g2_decap_8 FILLER_23_3052 ();
 sg13g2_decap_8 FILLER_23_3059 ();
 sg13g2_decap_8 FILLER_23_3066 ();
 sg13g2_decap_8 FILLER_23_3073 ();
 sg13g2_decap_8 FILLER_23_3080 ();
 sg13g2_decap_8 FILLER_23_3087 ();
 sg13g2_decap_8 FILLER_23_3094 ();
 sg13g2_decap_8 FILLER_23_3101 ();
 sg13g2_decap_8 FILLER_23_3108 ();
 sg13g2_decap_8 FILLER_23_3115 ();
 sg13g2_decap_8 FILLER_23_3122 ();
 sg13g2_decap_8 FILLER_23_3129 ();
 sg13g2_decap_8 FILLER_23_3136 ();
 sg13g2_decap_8 FILLER_23_3143 ();
 sg13g2_decap_8 FILLER_23_3150 ();
 sg13g2_decap_8 FILLER_23_3157 ();
 sg13g2_decap_8 FILLER_23_3164 ();
 sg13g2_decap_8 FILLER_23_3171 ();
 sg13g2_decap_8 FILLER_23_3178 ();
 sg13g2_decap_8 FILLER_23_3185 ();
 sg13g2_decap_8 FILLER_23_3192 ();
 sg13g2_decap_8 FILLER_23_3199 ();
 sg13g2_decap_8 FILLER_23_3206 ();
 sg13g2_decap_8 FILLER_23_3213 ();
 sg13g2_decap_8 FILLER_23_3220 ();
 sg13g2_decap_8 FILLER_23_3227 ();
 sg13g2_decap_8 FILLER_23_3234 ();
 sg13g2_decap_8 FILLER_23_3241 ();
 sg13g2_decap_8 FILLER_23_3248 ();
 sg13g2_decap_8 FILLER_23_3255 ();
 sg13g2_decap_8 FILLER_23_3262 ();
 sg13g2_decap_8 FILLER_23_3269 ();
 sg13g2_decap_8 FILLER_23_3276 ();
 sg13g2_decap_8 FILLER_23_3283 ();
 sg13g2_decap_8 FILLER_23_3290 ();
 sg13g2_decap_8 FILLER_23_3297 ();
 sg13g2_decap_8 FILLER_23_3304 ();
 sg13g2_decap_8 FILLER_23_3311 ();
 sg13g2_decap_8 FILLER_23_3318 ();
 sg13g2_decap_8 FILLER_23_3325 ();
 sg13g2_decap_8 FILLER_23_3332 ();
 sg13g2_decap_8 FILLER_23_3339 ();
 sg13g2_decap_8 FILLER_23_3346 ();
 sg13g2_decap_8 FILLER_23_3353 ();
 sg13g2_decap_8 FILLER_23_3360 ();
 sg13g2_decap_8 FILLER_23_3367 ();
 sg13g2_decap_8 FILLER_23_3374 ();
 sg13g2_decap_8 FILLER_23_3381 ();
 sg13g2_decap_8 FILLER_23_3388 ();
 sg13g2_decap_8 FILLER_23_3395 ();
 sg13g2_decap_8 FILLER_23_3402 ();
 sg13g2_decap_8 FILLER_23_3409 ();
 sg13g2_decap_8 FILLER_23_3416 ();
 sg13g2_decap_8 FILLER_23_3423 ();
 sg13g2_decap_8 FILLER_23_3430 ();
 sg13g2_decap_8 FILLER_23_3437 ();
 sg13g2_decap_8 FILLER_23_3444 ();
 sg13g2_decap_8 FILLER_23_3451 ();
 sg13g2_decap_8 FILLER_23_3458 ();
 sg13g2_decap_8 FILLER_23_3465 ();
 sg13g2_decap_8 FILLER_23_3472 ();
 sg13g2_decap_8 FILLER_23_3479 ();
 sg13g2_decap_8 FILLER_23_3486 ();
 sg13g2_decap_8 FILLER_23_3493 ();
 sg13g2_decap_8 FILLER_23_3500 ();
 sg13g2_decap_8 FILLER_23_3507 ();
 sg13g2_decap_8 FILLER_23_3514 ();
 sg13g2_decap_8 FILLER_23_3521 ();
 sg13g2_decap_8 FILLER_23_3528 ();
 sg13g2_decap_8 FILLER_23_3535 ();
 sg13g2_decap_8 FILLER_23_3542 ();
 sg13g2_decap_8 FILLER_23_3549 ();
 sg13g2_decap_8 FILLER_23_3556 ();
 sg13g2_decap_8 FILLER_23_3563 ();
 sg13g2_decap_8 FILLER_23_3570 ();
 sg13g2_fill_2 FILLER_23_3577 ();
 sg13g2_fill_1 FILLER_23_3579 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_decap_8 FILLER_24_406 ();
 sg13g2_decap_8 FILLER_24_413 ();
 sg13g2_decap_8 FILLER_24_420 ();
 sg13g2_decap_8 FILLER_24_427 ();
 sg13g2_decap_8 FILLER_24_434 ();
 sg13g2_decap_8 FILLER_24_441 ();
 sg13g2_decap_8 FILLER_24_448 ();
 sg13g2_decap_8 FILLER_24_455 ();
 sg13g2_decap_8 FILLER_24_462 ();
 sg13g2_decap_8 FILLER_24_469 ();
 sg13g2_decap_8 FILLER_24_476 ();
 sg13g2_decap_8 FILLER_24_483 ();
 sg13g2_decap_8 FILLER_24_490 ();
 sg13g2_decap_8 FILLER_24_497 ();
 sg13g2_decap_8 FILLER_24_504 ();
 sg13g2_decap_8 FILLER_24_511 ();
 sg13g2_decap_8 FILLER_24_518 ();
 sg13g2_decap_8 FILLER_24_525 ();
 sg13g2_decap_8 FILLER_24_532 ();
 sg13g2_decap_8 FILLER_24_539 ();
 sg13g2_decap_8 FILLER_24_546 ();
 sg13g2_decap_8 FILLER_24_553 ();
 sg13g2_decap_8 FILLER_24_560 ();
 sg13g2_decap_8 FILLER_24_567 ();
 sg13g2_decap_8 FILLER_24_574 ();
 sg13g2_decap_8 FILLER_24_581 ();
 sg13g2_decap_8 FILLER_24_588 ();
 sg13g2_decap_8 FILLER_24_595 ();
 sg13g2_decap_8 FILLER_24_602 ();
 sg13g2_decap_8 FILLER_24_609 ();
 sg13g2_decap_8 FILLER_24_616 ();
 sg13g2_decap_8 FILLER_24_623 ();
 sg13g2_decap_8 FILLER_24_630 ();
 sg13g2_decap_8 FILLER_24_637 ();
 sg13g2_decap_8 FILLER_24_644 ();
 sg13g2_decap_8 FILLER_24_651 ();
 sg13g2_decap_8 FILLER_24_658 ();
 sg13g2_decap_8 FILLER_24_665 ();
 sg13g2_decap_8 FILLER_24_672 ();
 sg13g2_decap_8 FILLER_24_679 ();
 sg13g2_decap_8 FILLER_24_686 ();
 sg13g2_decap_8 FILLER_24_693 ();
 sg13g2_decap_8 FILLER_24_700 ();
 sg13g2_decap_8 FILLER_24_707 ();
 sg13g2_decap_8 FILLER_24_714 ();
 sg13g2_decap_8 FILLER_24_721 ();
 sg13g2_decap_8 FILLER_24_728 ();
 sg13g2_decap_8 FILLER_24_735 ();
 sg13g2_decap_8 FILLER_24_742 ();
 sg13g2_decap_8 FILLER_24_749 ();
 sg13g2_decap_8 FILLER_24_756 ();
 sg13g2_decap_8 FILLER_24_763 ();
 sg13g2_decap_8 FILLER_24_770 ();
 sg13g2_decap_8 FILLER_24_777 ();
 sg13g2_decap_8 FILLER_24_784 ();
 sg13g2_decap_8 FILLER_24_791 ();
 sg13g2_decap_8 FILLER_24_798 ();
 sg13g2_decap_8 FILLER_24_805 ();
 sg13g2_decap_8 FILLER_24_812 ();
 sg13g2_decap_8 FILLER_24_819 ();
 sg13g2_decap_8 FILLER_24_826 ();
 sg13g2_decap_8 FILLER_24_833 ();
 sg13g2_decap_8 FILLER_24_840 ();
 sg13g2_decap_8 FILLER_24_847 ();
 sg13g2_decap_8 FILLER_24_854 ();
 sg13g2_decap_8 FILLER_24_861 ();
 sg13g2_decap_8 FILLER_24_868 ();
 sg13g2_decap_8 FILLER_24_875 ();
 sg13g2_decap_8 FILLER_24_882 ();
 sg13g2_decap_8 FILLER_24_889 ();
 sg13g2_decap_8 FILLER_24_896 ();
 sg13g2_decap_8 FILLER_24_903 ();
 sg13g2_decap_8 FILLER_24_910 ();
 sg13g2_decap_8 FILLER_24_917 ();
 sg13g2_decap_8 FILLER_24_924 ();
 sg13g2_decap_8 FILLER_24_931 ();
 sg13g2_decap_8 FILLER_24_938 ();
 sg13g2_decap_8 FILLER_24_945 ();
 sg13g2_decap_8 FILLER_24_952 ();
 sg13g2_decap_8 FILLER_24_959 ();
 sg13g2_decap_8 FILLER_24_966 ();
 sg13g2_decap_8 FILLER_24_973 ();
 sg13g2_decap_8 FILLER_24_980 ();
 sg13g2_decap_8 FILLER_24_987 ();
 sg13g2_decap_8 FILLER_24_994 ();
 sg13g2_decap_8 FILLER_24_1001 ();
 sg13g2_decap_8 FILLER_24_1008 ();
 sg13g2_decap_8 FILLER_24_1015 ();
 sg13g2_decap_8 FILLER_24_1022 ();
 sg13g2_decap_8 FILLER_24_1029 ();
 sg13g2_decap_8 FILLER_24_1036 ();
 sg13g2_decap_8 FILLER_24_1043 ();
 sg13g2_decap_8 FILLER_24_1050 ();
 sg13g2_decap_8 FILLER_24_1057 ();
 sg13g2_decap_8 FILLER_24_1064 ();
 sg13g2_decap_8 FILLER_24_1071 ();
 sg13g2_decap_8 FILLER_24_1078 ();
 sg13g2_decap_8 FILLER_24_1085 ();
 sg13g2_decap_8 FILLER_24_1092 ();
 sg13g2_decap_8 FILLER_24_1099 ();
 sg13g2_decap_8 FILLER_24_1106 ();
 sg13g2_decap_8 FILLER_24_1113 ();
 sg13g2_decap_8 FILLER_24_1120 ();
 sg13g2_decap_8 FILLER_24_1127 ();
 sg13g2_decap_8 FILLER_24_1134 ();
 sg13g2_decap_8 FILLER_24_1141 ();
 sg13g2_decap_8 FILLER_24_1148 ();
 sg13g2_decap_8 FILLER_24_1155 ();
 sg13g2_decap_8 FILLER_24_1162 ();
 sg13g2_decap_8 FILLER_24_1169 ();
 sg13g2_decap_8 FILLER_24_1176 ();
 sg13g2_decap_8 FILLER_24_1183 ();
 sg13g2_decap_8 FILLER_24_1190 ();
 sg13g2_decap_8 FILLER_24_1197 ();
 sg13g2_decap_8 FILLER_24_1204 ();
 sg13g2_decap_8 FILLER_24_1211 ();
 sg13g2_decap_8 FILLER_24_1218 ();
 sg13g2_decap_8 FILLER_24_1225 ();
 sg13g2_decap_8 FILLER_24_1232 ();
 sg13g2_decap_8 FILLER_24_1239 ();
 sg13g2_decap_8 FILLER_24_1246 ();
 sg13g2_decap_8 FILLER_24_1253 ();
 sg13g2_decap_8 FILLER_24_1260 ();
 sg13g2_decap_8 FILLER_24_1267 ();
 sg13g2_decap_8 FILLER_24_1274 ();
 sg13g2_decap_8 FILLER_24_1281 ();
 sg13g2_decap_8 FILLER_24_1288 ();
 sg13g2_decap_8 FILLER_24_1295 ();
 sg13g2_decap_8 FILLER_24_1302 ();
 sg13g2_decap_8 FILLER_24_1309 ();
 sg13g2_decap_8 FILLER_24_1316 ();
 sg13g2_decap_8 FILLER_24_1323 ();
 sg13g2_decap_8 FILLER_24_1330 ();
 sg13g2_decap_8 FILLER_24_1337 ();
 sg13g2_decap_8 FILLER_24_1344 ();
 sg13g2_decap_8 FILLER_24_1351 ();
 sg13g2_decap_8 FILLER_24_1358 ();
 sg13g2_decap_8 FILLER_24_1365 ();
 sg13g2_decap_8 FILLER_24_1372 ();
 sg13g2_decap_8 FILLER_24_1379 ();
 sg13g2_decap_8 FILLER_24_1386 ();
 sg13g2_decap_8 FILLER_24_1393 ();
 sg13g2_decap_8 FILLER_24_1400 ();
 sg13g2_decap_8 FILLER_24_1407 ();
 sg13g2_decap_8 FILLER_24_1414 ();
 sg13g2_decap_8 FILLER_24_1421 ();
 sg13g2_decap_8 FILLER_24_1428 ();
 sg13g2_decap_8 FILLER_24_1435 ();
 sg13g2_decap_8 FILLER_24_1442 ();
 sg13g2_decap_8 FILLER_24_1449 ();
 sg13g2_decap_8 FILLER_24_1456 ();
 sg13g2_decap_8 FILLER_24_1463 ();
 sg13g2_decap_8 FILLER_24_1470 ();
 sg13g2_decap_8 FILLER_24_1477 ();
 sg13g2_decap_8 FILLER_24_1484 ();
 sg13g2_decap_8 FILLER_24_1491 ();
 sg13g2_decap_8 FILLER_24_1498 ();
 sg13g2_decap_8 FILLER_24_1505 ();
 sg13g2_decap_8 FILLER_24_1512 ();
 sg13g2_decap_8 FILLER_24_1519 ();
 sg13g2_decap_8 FILLER_24_1526 ();
 sg13g2_decap_8 FILLER_24_1533 ();
 sg13g2_decap_8 FILLER_24_1540 ();
 sg13g2_decap_8 FILLER_24_1547 ();
 sg13g2_decap_8 FILLER_24_1554 ();
 sg13g2_decap_8 FILLER_24_1561 ();
 sg13g2_decap_8 FILLER_24_1568 ();
 sg13g2_decap_8 FILLER_24_1575 ();
 sg13g2_decap_8 FILLER_24_1582 ();
 sg13g2_decap_8 FILLER_24_1589 ();
 sg13g2_decap_8 FILLER_24_1596 ();
 sg13g2_decap_8 FILLER_24_1603 ();
 sg13g2_decap_8 FILLER_24_1610 ();
 sg13g2_decap_8 FILLER_24_1617 ();
 sg13g2_decap_8 FILLER_24_1624 ();
 sg13g2_decap_8 FILLER_24_1631 ();
 sg13g2_decap_8 FILLER_24_1638 ();
 sg13g2_decap_8 FILLER_24_1645 ();
 sg13g2_decap_8 FILLER_24_1652 ();
 sg13g2_decap_8 FILLER_24_1659 ();
 sg13g2_decap_8 FILLER_24_1666 ();
 sg13g2_decap_8 FILLER_24_1673 ();
 sg13g2_decap_8 FILLER_24_1680 ();
 sg13g2_decap_8 FILLER_24_1687 ();
 sg13g2_decap_8 FILLER_24_1694 ();
 sg13g2_decap_8 FILLER_24_1701 ();
 sg13g2_decap_8 FILLER_24_1708 ();
 sg13g2_decap_8 FILLER_24_1715 ();
 sg13g2_decap_8 FILLER_24_1722 ();
 sg13g2_decap_8 FILLER_24_1729 ();
 sg13g2_decap_8 FILLER_24_1736 ();
 sg13g2_decap_8 FILLER_24_1743 ();
 sg13g2_decap_8 FILLER_24_1750 ();
 sg13g2_decap_8 FILLER_24_1757 ();
 sg13g2_decap_8 FILLER_24_1764 ();
 sg13g2_decap_8 FILLER_24_1771 ();
 sg13g2_decap_8 FILLER_24_1778 ();
 sg13g2_decap_8 FILLER_24_1785 ();
 sg13g2_decap_8 FILLER_24_1792 ();
 sg13g2_decap_8 FILLER_24_1799 ();
 sg13g2_decap_8 FILLER_24_1806 ();
 sg13g2_decap_8 FILLER_24_1813 ();
 sg13g2_decap_8 FILLER_24_1820 ();
 sg13g2_decap_8 FILLER_24_1827 ();
 sg13g2_decap_8 FILLER_24_1834 ();
 sg13g2_decap_8 FILLER_24_1841 ();
 sg13g2_decap_8 FILLER_24_1848 ();
 sg13g2_decap_8 FILLER_24_1855 ();
 sg13g2_decap_8 FILLER_24_1862 ();
 sg13g2_decap_8 FILLER_24_1869 ();
 sg13g2_decap_8 FILLER_24_1876 ();
 sg13g2_decap_8 FILLER_24_1883 ();
 sg13g2_decap_8 FILLER_24_1890 ();
 sg13g2_decap_8 FILLER_24_1897 ();
 sg13g2_decap_8 FILLER_24_1904 ();
 sg13g2_decap_8 FILLER_24_1911 ();
 sg13g2_decap_8 FILLER_24_1918 ();
 sg13g2_decap_8 FILLER_24_1925 ();
 sg13g2_decap_8 FILLER_24_1932 ();
 sg13g2_decap_8 FILLER_24_1939 ();
 sg13g2_decap_8 FILLER_24_1946 ();
 sg13g2_decap_8 FILLER_24_1953 ();
 sg13g2_decap_8 FILLER_24_1960 ();
 sg13g2_decap_8 FILLER_24_1967 ();
 sg13g2_decap_8 FILLER_24_1974 ();
 sg13g2_decap_8 FILLER_24_1981 ();
 sg13g2_decap_8 FILLER_24_1988 ();
 sg13g2_decap_8 FILLER_24_1995 ();
 sg13g2_decap_8 FILLER_24_2002 ();
 sg13g2_decap_8 FILLER_24_2009 ();
 sg13g2_decap_8 FILLER_24_2016 ();
 sg13g2_decap_8 FILLER_24_2023 ();
 sg13g2_decap_8 FILLER_24_2030 ();
 sg13g2_decap_8 FILLER_24_2037 ();
 sg13g2_decap_8 FILLER_24_2044 ();
 sg13g2_decap_8 FILLER_24_2051 ();
 sg13g2_decap_8 FILLER_24_2058 ();
 sg13g2_decap_8 FILLER_24_2065 ();
 sg13g2_decap_8 FILLER_24_2072 ();
 sg13g2_decap_8 FILLER_24_2079 ();
 sg13g2_decap_8 FILLER_24_2086 ();
 sg13g2_decap_8 FILLER_24_2093 ();
 sg13g2_decap_8 FILLER_24_2100 ();
 sg13g2_decap_8 FILLER_24_2107 ();
 sg13g2_decap_8 FILLER_24_2114 ();
 sg13g2_decap_8 FILLER_24_2121 ();
 sg13g2_decap_8 FILLER_24_2128 ();
 sg13g2_decap_8 FILLER_24_2135 ();
 sg13g2_decap_8 FILLER_24_2142 ();
 sg13g2_decap_8 FILLER_24_2149 ();
 sg13g2_decap_8 FILLER_24_2156 ();
 sg13g2_decap_8 FILLER_24_2163 ();
 sg13g2_decap_8 FILLER_24_2170 ();
 sg13g2_decap_8 FILLER_24_2177 ();
 sg13g2_decap_8 FILLER_24_2184 ();
 sg13g2_decap_8 FILLER_24_2191 ();
 sg13g2_decap_8 FILLER_24_2198 ();
 sg13g2_decap_8 FILLER_24_2205 ();
 sg13g2_decap_8 FILLER_24_2212 ();
 sg13g2_decap_8 FILLER_24_2219 ();
 sg13g2_decap_8 FILLER_24_2226 ();
 sg13g2_decap_8 FILLER_24_2233 ();
 sg13g2_decap_8 FILLER_24_2240 ();
 sg13g2_decap_8 FILLER_24_2247 ();
 sg13g2_decap_8 FILLER_24_2254 ();
 sg13g2_decap_8 FILLER_24_2261 ();
 sg13g2_decap_8 FILLER_24_2268 ();
 sg13g2_decap_8 FILLER_24_2275 ();
 sg13g2_decap_8 FILLER_24_2282 ();
 sg13g2_decap_8 FILLER_24_2289 ();
 sg13g2_decap_8 FILLER_24_2296 ();
 sg13g2_decap_8 FILLER_24_2303 ();
 sg13g2_decap_8 FILLER_24_2310 ();
 sg13g2_decap_8 FILLER_24_2317 ();
 sg13g2_decap_8 FILLER_24_2324 ();
 sg13g2_decap_8 FILLER_24_2331 ();
 sg13g2_decap_8 FILLER_24_2338 ();
 sg13g2_decap_8 FILLER_24_2345 ();
 sg13g2_decap_8 FILLER_24_2352 ();
 sg13g2_decap_8 FILLER_24_2359 ();
 sg13g2_decap_8 FILLER_24_2366 ();
 sg13g2_decap_8 FILLER_24_2373 ();
 sg13g2_decap_8 FILLER_24_2380 ();
 sg13g2_decap_8 FILLER_24_2387 ();
 sg13g2_decap_8 FILLER_24_2394 ();
 sg13g2_decap_8 FILLER_24_2401 ();
 sg13g2_decap_8 FILLER_24_2408 ();
 sg13g2_decap_8 FILLER_24_2415 ();
 sg13g2_decap_8 FILLER_24_2422 ();
 sg13g2_decap_8 FILLER_24_2429 ();
 sg13g2_decap_8 FILLER_24_2436 ();
 sg13g2_decap_8 FILLER_24_2443 ();
 sg13g2_decap_8 FILLER_24_2450 ();
 sg13g2_decap_8 FILLER_24_2457 ();
 sg13g2_decap_8 FILLER_24_2464 ();
 sg13g2_decap_8 FILLER_24_2471 ();
 sg13g2_decap_8 FILLER_24_2478 ();
 sg13g2_decap_8 FILLER_24_2485 ();
 sg13g2_decap_8 FILLER_24_2492 ();
 sg13g2_decap_8 FILLER_24_2499 ();
 sg13g2_decap_8 FILLER_24_2506 ();
 sg13g2_decap_8 FILLER_24_2513 ();
 sg13g2_decap_8 FILLER_24_2520 ();
 sg13g2_decap_8 FILLER_24_2527 ();
 sg13g2_decap_8 FILLER_24_2534 ();
 sg13g2_decap_8 FILLER_24_2541 ();
 sg13g2_decap_8 FILLER_24_2548 ();
 sg13g2_decap_8 FILLER_24_2555 ();
 sg13g2_decap_8 FILLER_24_2562 ();
 sg13g2_decap_8 FILLER_24_2569 ();
 sg13g2_decap_8 FILLER_24_2576 ();
 sg13g2_decap_8 FILLER_24_2583 ();
 sg13g2_decap_8 FILLER_24_2590 ();
 sg13g2_decap_8 FILLER_24_2597 ();
 sg13g2_decap_8 FILLER_24_2604 ();
 sg13g2_decap_8 FILLER_24_2611 ();
 sg13g2_decap_8 FILLER_24_2618 ();
 sg13g2_decap_8 FILLER_24_2625 ();
 sg13g2_decap_8 FILLER_24_2632 ();
 sg13g2_decap_8 FILLER_24_2639 ();
 sg13g2_decap_8 FILLER_24_2646 ();
 sg13g2_decap_8 FILLER_24_2653 ();
 sg13g2_decap_8 FILLER_24_2660 ();
 sg13g2_decap_8 FILLER_24_2667 ();
 sg13g2_decap_8 FILLER_24_2674 ();
 sg13g2_decap_8 FILLER_24_2681 ();
 sg13g2_decap_8 FILLER_24_2688 ();
 sg13g2_decap_8 FILLER_24_2695 ();
 sg13g2_decap_8 FILLER_24_2702 ();
 sg13g2_decap_8 FILLER_24_2709 ();
 sg13g2_decap_8 FILLER_24_2716 ();
 sg13g2_decap_8 FILLER_24_2723 ();
 sg13g2_decap_8 FILLER_24_2730 ();
 sg13g2_decap_8 FILLER_24_2737 ();
 sg13g2_decap_8 FILLER_24_2744 ();
 sg13g2_decap_8 FILLER_24_2751 ();
 sg13g2_decap_8 FILLER_24_2758 ();
 sg13g2_decap_8 FILLER_24_2765 ();
 sg13g2_decap_8 FILLER_24_2772 ();
 sg13g2_decap_8 FILLER_24_2779 ();
 sg13g2_decap_8 FILLER_24_2786 ();
 sg13g2_decap_8 FILLER_24_2793 ();
 sg13g2_decap_8 FILLER_24_2800 ();
 sg13g2_decap_8 FILLER_24_2807 ();
 sg13g2_decap_8 FILLER_24_2814 ();
 sg13g2_decap_8 FILLER_24_2821 ();
 sg13g2_decap_8 FILLER_24_2828 ();
 sg13g2_decap_8 FILLER_24_2835 ();
 sg13g2_decap_8 FILLER_24_2842 ();
 sg13g2_decap_8 FILLER_24_2849 ();
 sg13g2_decap_8 FILLER_24_2856 ();
 sg13g2_decap_8 FILLER_24_2863 ();
 sg13g2_decap_8 FILLER_24_2870 ();
 sg13g2_decap_8 FILLER_24_2877 ();
 sg13g2_decap_8 FILLER_24_2884 ();
 sg13g2_decap_8 FILLER_24_2891 ();
 sg13g2_decap_8 FILLER_24_2898 ();
 sg13g2_decap_8 FILLER_24_2905 ();
 sg13g2_decap_8 FILLER_24_2912 ();
 sg13g2_decap_8 FILLER_24_2919 ();
 sg13g2_decap_8 FILLER_24_2926 ();
 sg13g2_decap_8 FILLER_24_2933 ();
 sg13g2_decap_8 FILLER_24_2940 ();
 sg13g2_decap_8 FILLER_24_2947 ();
 sg13g2_decap_8 FILLER_24_2954 ();
 sg13g2_decap_8 FILLER_24_2961 ();
 sg13g2_decap_8 FILLER_24_2968 ();
 sg13g2_decap_8 FILLER_24_2975 ();
 sg13g2_decap_8 FILLER_24_2982 ();
 sg13g2_decap_8 FILLER_24_2989 ();
 sg13g2_decap_8 FILLER_24_2996 ();
 sg13g2_decap_8 FILLER_24_3003 ();
 sg13g2_decap_8 FILLER_24_3010 ();
 sg13g2_decap_8 FILLER_24_3017 ();
 sg13g2_decap_8 FILLER_24_3024 ();
 sg13g2_decap_8 FILLER_24_3031 ();
 sg13g2_decap_8 FILLER_24_3038 ();
 sg13g2_decap_8 FILLER_24_3045 ();
 sg13g2_decap_8 FILLER_24_3052 ();
 sg13g2_decap_8 FILLER_24_3059 ();
 sg13g2_decap_8 FILLER_24_3066 ();
 sg13g2_decap_8 FILLER_24_3073 ();
 sg13g2_decap_8 FILLER_24_3080 ();
 sg13g2_decap_8 FILLER_24_3087 ();
 sg13g2_decap_8 FILLER_24_3094 ();
 sg13g2_decap_8 FILLER_24_3101 ();
 sg13g2_decap_8 FILLER_24_3108 ();
 sg13g2_decap_8 FILLER_24_3115 ();
 sg13g2_decap_8 FILLER_24_3122 ();
 sg13g2_decap_8 FILLER_24_3129 ();
 sg13g2_decap_8 FILLER_24_3136 ();
 sg13g2_decap_8 FILLER_24_3143 ();
 sg13g2_decap_8 FILLER_24_3150 ();
 sg13g2_decap_8 FILLER_24_3157 ();
 sg13g2_decap_8 FILLER_24_3164 ();
 sg13g2_decap_8 FILLER_24_3171 ();
 sg13g2_decap_8 FILLER_24_3178 ();
 sg13g2_decap_8 FILLER_24_3185 ();
 sg13g2_decap_8 FILLER_24_3192 ();
 sg13g2_decap_8 FILLER_24_3199 ();
 sg13g2_decap_8 FILLER_24_3206 ();
 sg13g2_decap_8 FILLER_24_3213 ();
 sg13g2_decap_8 FILLER_24_3220 ();
 sg13g2_decap_8 FILLER_24_3227 ();
 sg13g2_decap_8 FILLER_24_3234 ();
 sg13g2_decap_8 FILLER_24_3241 ();
 sg13g2_decap_8 FILLER_24_3248 ();
 sg13g2_decap_8 FILLER_24_3255 ();
 sg13g2_decap_8 FILLER_24_3262 ();
 sg13g2_decap_8 FILLER_24_3269 ();
 sg13g2_decap_8 FILLER_24_3276 ();
 sg13g2_decap_8 FILLER_24_3283 ();
 sg13g2_decap_8 FILLER_24_3290 ();
 sg13g2_decap_8 FILLER_24_3297 ();
 sg13g2_decap_8 FILLER_24_3304 ();
 sg13g2_decap_8 FILLER_24_3311 ();
 sg13g2_decap_8 FILLER_24_3318 ();
 sg13g2_decap_8 FILLER_24_3325 ();
 sg13g2_decap_8 FILLER_24_3332 ();
 sg13g2_decap_8 FILLER_24_3339 ();
 sg13g2_decap_8 FILLER_24_3346 ();
 sg13g2_decap_8 FILLER_24_3353 ();
 sg13g2_decap_8 FILLER_24_3360 ();
 sg13g2_decap_8 FILLER_24_3367 ();
 sg13g2_decap_8 FILLER_24_3374 ();
 sg13g2_decap_8 FILLER_24_3381 ();
 sg13g2_decap_8 FILLER_24_3388 ();
 sg13g2_decap_8 FILLER_24_3395 ();
 sg13g2_decap_8 FILLER_24_3402 ();
 sg13g2_decap_8 FILLER_24_3409 ();
 sg13g2_decap_8 FILLER_24_3416 ();
 sg13g2_decap_8 FILLER_24_3423 ();
 sg13g2_decap_8 FILLER_24_3430 ();
 sg13g2_decap_8 FILLER_24_3437 ();
 sg13g2_decap_8 FILLER_24_3444 ();
 sg13g2_decap_8 FILLER_24_3451 ();
 sg13g2_decap_8 FILLER_24_3458 ();
 sg13g2_decap_8 FILLER_24_3465 ();
 sg13g2_decap_8 FILLER_24_3472 ();
 sg13g2_decap_8 FILLER_24_3479 ();
 sg13g2_decap_8 FILLER_24_3486 ();
 sg13g2_decap_8 FILLER_24_3493 ();
 sg13g2_decap_8 FILLER_24_3500 ();
 sg13g2_decap_8 FILLER_24_3507 ();
 sg13g2_decap_8 FILLER_24_3514 ();
 sg13g2_decap_8 FILLER_24_3521 ();
 sg13g2_decap_8 FILLER_24_3528 ();
 sg13g2_decap_8 FILLER_24_3535 ();
 sg13g2_decap_8 FILLER_24_3542 ();
 sg13g2_decap_8 FILLER_24_3549 ();
 sg13g2_decap_8 FILLER_24_3556 ();
 sg13g2_decap_8 FILLER_24_3563 ();
 sg13g2_decap_8 FILLER_24_3570 ();
 sg13g2_fill_2 FILLER_24_3577 ();
 sg13g2_fill_1 FILLER_24_3579 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_decap_8 FILLER_25_406 ();
 sg13g2_decap_8 FILLER_25_413 ();
 sg13g2_decap_8 FILLER_25_420 ();
 sg13g2_decap_8 FILLER_25_427 ();
 sg13g2_decap_8 FILLER_25_434 ();
 sg13g2_decap_8 FILLER_25_441 ();
 sg13g2_decap_8 FILLER_25_448 ();
 sg13g2_decap_8 FILLER_25_455 ();
 sg13g2_decap_8 FILLER_25_462 ();
 sg13g2_decap_8 FILLER_25_469 ();
 sg13g2_decap_8 FILLER_25_476 ();
 sg13g2_decap_8 FILLER_25_483 ();
 sg13g2_decap_8 FILLER_25_490 ();
 sg13g2_decap_8 FILLER_25_497 ();
 sg13g2_decap_8 FILLER_25_504 ();
 sg13g2_decap_8 FILLER_25_511 ();
 sg13g2_decap_8 FILLER_25_518 ();
 sg13g2_decap_8 FILLER_25_525 ();
 sg13g2_decap_8 FILLER_25_532 ();
 sg13g2_decap_8 FILLER_25_539 ();
 sg13g2_decap_8 FILLER_25_546 ();
 sg13g2_decap_8 FILLER_25_553 ();
 sg13g2_decap_8 FILLER_25_560 ();
 sg13g2_decap_8 FILLER_25_567 ();
 sg13g2_decap_8 FILLER_25_574 ();
 sg13g2_decap_8 FILLER_25_581 ();
 sg13g2_decap_8 FILLER_25_588 ();
 sg13g2_decap_8 FILLER_25_595 ();
 sg13g2_decap_8 FILLER_25_602 ();
 sg13g2_decap_8 FILLER_25_609 ();
 sg13g2_decap_8 FILLER_25_616 ();
 sg13g2_decap_8 FILLER_25_623 ();
 sg13g2_decap_8 FILLER_25_630 ();
 sg13g2_decap_8 FILLER_25_637 ();
 sg13g2_decap_8 FILLER_25_644 ();
 sg13g2_decap_8 FILLER_25_651 ();
 sg13g2_decap_8 FILLER_25_658 ();
 sg13g2_decap_8 FILLER_25_665 ();
 sg13g2_decap_8 FILLER_25_672 ();
 sg13g2_decap_8 FILLER_25_679 ();
 sg13g2_decap_8 FILLER_25_686 ();
 sg13g2_decap_8 FILLER_25_693 ();
 sg13g2_decap_8 FILLER_25_700 ();
 sg13g2_decap_8 FILLER_25_707 ();
 sg13g2_decap_8 FILLER_25_714 ();
 sg13g2_decap_8 FILLER_25_721 ();
 sg13g2_decap_8 FILLER_25_728 ();
 sg13g2_decap_8 FILLER_25_735 ();
 sg13g2_decap_8 FILLER_25_742 ();
 sg13g2_decap_8 FILLER_25_749 ();
 sg13g2_decap_8 FILLER_25_756 ();
 sg13g2_decap_8 FILLER_25_763 ();
 sg13g2_decap_8 FILLER_25_770 ();
 sg13g2_decap_8 FILLER_25_777 ();
 sg13g2_decap_8 FILLER_25_784 ();
 sg13g2_decap_8 FILLER_25_791 ();
 sg13g2_decap_8 FILLER_25_798 ();
 sg13g2_decap_8 FILLER_25_805 ();
 sg13g2_decap_8 FILLER_25_812 ();
 sg13g2_decap_8 FILLER_25_819 ();
 sg13g2_decap_8 FILLER_25_826 ();
 sg13g2_decap_8 FILLER_25_833 ();
 sg13g2_decap_8 FILLER_25_840 ();
 sg13g2_decap_8 FILLER_25_847 ();
 sg13g2_decap_8 FILLER_25_854 ();
 sg13g2_decap_8 FILLER_25_861 ();
 sg13g2_decap_8 FILLER_25_868 ();
 sg13g2_decap_8 FILLER_25_875 ();
 sg13g2_decap_8 FILLER_25_882 ();
 sg13g2_decap_8 FILLER_25_889 ();
 sg13g2_decap_8 FILLER_25_896 ();
 sg13g2_decap_8 FILLER_25_903 ();
 sg13g2_decap_8 FILLER_25_910 ();
 sg13g2_decap_8 FILLER_25_917 ();
 sg13g2_decap_8 FILLER_25_924 ();
 sg13g2_decap_8 FILLER_25_931 ();
 sg13g2_decap_8 FILLER_25_938 ();
 sg13g2_decap_8 FILLER_25_945 ();
 sg13g2_decap_8 FILLER_25_952 ();
 sg13g2_decap_8 FILLER_25_959 ();
 sg13g2_decap_8 FILLER_25_966 ();
 sg13g2_decap_8 FILLER_25_973 ();
 sg13g2_decap_8 FILLER_25_980 ();
 sg13g2_decap_8 FILLER_25_987 ();
 sg13g2_decap_8 FILLER_25_994 ();
 sg13g2_decap_8 FILLER_25_1001 ();
 sg13g2_decap_8 FILLER_25_1008 ();
 sg13g2_decap_8 FILLER_25_1015 ();
 sg13g2_decap_8 FILLER_25_1022 ();
 sg13g2_decap_8 FILLER_25_1029 ();
 sg13g2_decap_8 FILLER_25_1036 ();
 sg13g2_decap_8 FILLER_25_1043 ();
 sg13g2_decap_8 FILLER_25_1050 ();
 sg13g2_decap_8 FILLER_25_1057 ();
 sg13g2_decap_8 FILLER_25_1064 ();
 sg13g2_decap_8 FILLER_25_1071 ();
 sg13g2_decap_8 FILLER_25_1078 ();
 sg13g2_decap_8 FILLER_25_1085 ();
 sg13g2_decap_8 FILLER_25_1092 ();
 sg13g2_decap_8 FILLER_25_1099 ();
 sg13g2_decap_8 FILLER_25_1106 ();
 sg13g2_decap_8 FILLER_25_1113 ();
 sg13g2_decap_8 FILLER_25_1120 ();
 sg13g2_decap_8 FILLER_25_1127 ();
 sg13g2_decap_8 FILLER_25_1134 ();
 sg13g2_decap_8 FILLER_25_1141 ();
 sg13g2_decap_8 FILLER_25_1148 ();
 sg13g2_decap_8 FILLER_25_1155 ();
 sg13g2_decap_8 FILLER_25_1162 ();
 sg13g2_decap_8 FILLER_25_1169 ();
 sg13g2_decap_8 FILLER_25_1176 ();
 sg13g2_decap_8 FILLER_25_1183 ();
 sg13g2_decap_8 FILLER_25_1190 ();
 sg13g2_decap_8 FILLER_25_1197 ();
 sg13g2_decap_8 FILLER_25_1204 ();
 sg13g2_decap_8 FILLER_25_1211 ();
 sg13g2_decap_8 FILLER_25_1218 ();
 sg13g2_decap_8 FILLER_25_1225 ();
 sg13g2_decap_8 FILLER_25_1232 ();
 sg13g2_decap_8 FILLER_25_1239 ();
 sg13g2_decap_8 FILLER_25_1246 ();
 sg13g2_decap_8 FILLER_25_1253 ();
 sg13g2_decap_8 FILLER_25_1260 ();
 sg13g2_decap_8 FILLER_25_1267 ();
 sg13g2_decap_8 FILLER_25_1274 ();
 sg13g2_decap_8 FILLER_25_1281 ();
 sg13g2_decap_8 FILLER_25_1288 ();
 sg13g2_decap_8 FILLER_25_1295 ();
 sg13g2_decap_8 FILLER_25_1302 ();
 sg13g2_decap_8 FILLER_25_1309 ();
 sg13g2_decap_8 FILLER_25_1316 ();
 sg13g2_decap_8 FILLER_25_1323 ();
 sg13g2_decap_8 FILLER_25_1330 ();
 sg13g2_decap_8 FILLER_25_1337 ();
 sg13g2_decap_8 FILLER_25_1344 ();
 sg13g2_decap_8 FILLER_25_1351 ();
 sg13g2_decap_8 FILLER_25_1358 ();
 sg13g2_decap_8 FILLER_25_1365 ();
 sg13g2_decap_8 FILLER_25_1372 ();
 sg13g2_decap_8 FILLER_25_1379 ();
 sg13g2_decap_8 FILLER_25_1386 ();
 sg13g2_decap_8 FILLER_25_1393 ();
 sg13g2_decap_8 FILLER_25_1400 ();
 sg13g2_decap_8 FILLER_25_1407 ();
 sg13g2_decap_8 FILLER_25_1414 ();
 sg13g2_decap_8 FILLER_25_1421 ();
 sg13g2_decap_8 FILLER_25_1428 ();
 sg13g2_decap_8 FILLER_25_1435 ();
 sg13g2_decap_8 FILLER_25_1442 ();
 sg13g2_decap_8 FILLER_25_1449 ();
 sg13g2_decap_8 FILLER_25_1456 ();
 sg13g2_decap_8 FILLER_25_1463 ();
 sg13g2_decap_8 FILLER_25_1470 ();
 sg13g2_decap_8 FILLER_25_1477 ();
 sg13g2_decap_8 FILLER_25_1484 ();
 sg13g2_decap_8 FILLER_25_1491 ();
 sg13g2_decap_8 FILLER_25_1498 ();
 sg13g2_decap_8 FILLER_25_1505 ();
 sg13g2_decap_8 FILLER_25_1512 ();
 sg13g2_decap_8 FILLER_25_1519 ();
 sg13g2_decap_8 FILLER_25_1526 ();
 sg13g2_decap_8 FILLER_25_1533 ();
 sg13g2_decap_8 FILLER_25_1540 ();
 sg13g2_decap_8 FILLER_25_1547 ();
 sg13g2_decap_8 FILLER_25_1554 ();
 sg13g2_decap_8 FILLER_25_1561 ();
 sg13g2_decap_8 FILLER_25_1568 ();
 sg13g2_decap_8 FILLER_25_1575 ();
 sg13g2_decap_8 FILLER_25_1582 ();
 sg13g2_decap_8 FILLER_25_1589 ();
 sg13g2_decap_8 FILLER_25_1596 ();
 sg13g2_decap_8 FILLER_25_1603 ();
 sg13g2_decap_8 FILLER_25_1610 ();
 sg13g2_decap_8 FILLER_25_1617 ();
 sg13g2_decap_8 FILLER_25_1624 ();
 sg13g2_decap_8 FILLER_25_1631 ();
 sg13g2_decap_8 FILLER_25_1638 ();
 sg13g2_decap_8 FILLER_25_1645 ();
 sg13g2_decap_8 FILLER_25_1652 ();
 sg13g2_decap_8 FILLER_25_1659 ();
 sg13g2_decap_8 FILLER_25_1666 ();
 sg13g2_decap_8 FILLER_25_1673 ();
 sg13g2_decap_8 FILLER_25_1680 ();
 sg13g2_decap_8 FILLER_25_1687 ();
 sg13g2_decap_8 FILLER_25_1694 ();
 sg13g2_decap_8 FILLER_25_1701 ();
 sg13g2_decap_8 FILLER_25_1708 ();
 sg13g2_decap_8 FILLER_25_1715 ();
 sg13g2_decap_8 FILLER_25_1722 ();
 sg13g2_decap_8 FILLER_25_1729 ();
 sg13g2_decap_8 FILLER_25_1736 ();
 sg13g2_decap_8 FILLER_25_1743 ();
 sg13g2_decap_8 FILLER_25_1750 ();
 sg13g2_decap_8 FILLER_25_1757 ();
 sg13g2_decap_8 FILLER_25_1764 ();
 sg13g2_decap_8 FILLER_25_1771 ();
 sg13g2_decap_8 FILLER_25_1778 ();
 sg13g2_decap_8 FILLER_25_1785 ();
 sg13g2_decap_8 FILLER_25_1792 ();
 sg13g2_decap_8 FILLER_25_1799 ();
 sg13g2_decap_8 FILLER_25_1806 ();
 sg13g2_decap_8 FILLER_25_1813 ();
 sg13g2_decap_8 FILLER_25_1820 ();
 sg13g2_decap_8 FILLER_25_1827 ();
 sg13g2_decap_8 FILLER_25_1834 ();
 sg13g2_decap_8 FILLER_25_1841 ();
 sg13g2_decap_8 FILLER_25_1848 ();
 sg13g2_decap_8 FILLER_25_1855 ();
 sg13g2_decap_8 FILLER_25_1862 ();
 sg13g2_decap_8 FILLER_25_1869 ();
 sg13g2_decap_8 FILLER_25_1876 ();
 sg13g2_decap_8 FILLER_25_1883 ();
 sg13g2_decap_8 FILLER_25_1890 ();
 sg13g2_decap_8 FILLER_25_1897 ();
 sg13g2_decap_8 FILLER_25_1904 ();
 sg13g2_decap_8 FILLER_25_1911 ();
 sg13g2_decap_8 FILLER_25_1918 ();
 sg13g2_decap_8 FILLER_25_1925 ();
 sg13g2_decap_8 FILLER_25_1932 ();
 sg13g2_decap_8 FILLER_25_1939 ();
 sg13g2_decap_8 FILLER_25_1946 ();
 sg13g2_decap_8 FILLER_25_1953 ();
 sg13g2_decap_8 FILLER_25_1960 ();
 sg13g2_decap_8 FILLER_25_1967 ();
 sg13g2_decap_8 FILLER_25_1974 ();
 sg13g2_decap_8 FILLER_25_1981 ();
 sg13g2_decap_8 FILLER_25_1988 ();
 sg13g2_decap_8 FILLER_25_1995 ();
 sg13g2_decap_8 FILLER_25_2002 ();
 sg13g2_decap_8 FILLER_25_2009 ();
 sg13g2_decap_8 FILLER_25_2016 ();
 sg13g2_decap_8 FILLER_25_2023 ();
 sg13g2_decap_8 FILLER_25_2030 ();
 sg13g2_decap_8 FILLER_25_2037 ();
 sg13g2_decap_8 FILLER_25_2044 ();
 sg13g2_decap_8 FILLER_25_2051 ();
 sg13g2_decap_8 FILLER_25_2058 ();
 sg13g2_decap_8 FILLER_25_2065 ();
 sg13g2_decap_8 FILLER_25_2072 ();
 sg13g2_decap_8 FILLER_25_2079 ();
 sg13g2_decap_8 FILLER_25_2086 ();
 sg13g2_decap_8 FILLER_25_2093 ();
 sg13g2_decap_8 FILLER_25_2100 ();
 sg13g2_decap_8 FILLER_25_2107 ();
 sg13g2_decap_8 FILLER_25_2114 ();
 sg13g2_decap_8 FILLER_25_2121 ();
 sg13g2_decap_8 FILLER_25_2128 ();
 sg13g2_decap_8 FILLER_25_2135 ();
 sg13g2_decap_8 FILLER_25_2142 ();
 sg13g2_decap_8 FILLER_25_2149 ();
 sg13g2_decap_8 FILLER_25_2156 ();
 sg13g2_decap_8 FILLER_25_2163 ();
 sg13g2_decap_8 FILLER_25_2170 ();
 sg13g2_decap_8 FILLER_25_2177 ();
 sg13g2_decap_8 FILLER_25_2184 ();
 sg13g2_decap_8 FILLER_25_2191 ();
 sg13g2_decap_8 FILLER_25_2198 ();
 sg13g2_decap_8 FILLER_25_2205 ();
 sg13g2_decap_8 FILLER_25_2212 ();
 sg13g2_decap_8 FILLER_25_2219 ();
 sg13g2_decap_8 FILLER_25_2226 ();
 sg13g2_decap_8 FILLER_25_2233 ();
 sg13g2_decap_8 FILLER_25_2240 ();
 sg13g2_decap_8 FILLER_25_2247 ();
 sg13g2_decap_8 FILLER_25_2254 ();
 sg13g2_decap_8 FILLER_25_2261 ();
 sg13g2_decap_8 FILLER_25_2268 ();
 sg13g2_decap_8 FILLER_25_2275 ();
 sg13g2_decap_8 FILLER_25_2282 ();
 sg13g2_decap_8 FILLER_25_2289 ();
 sg13g2_decap_8 FILLER_25_2296 ();
 sg13g2_decap_8 FILLER_25_2303 ();
 sg13g2_decap_8 FILLER_25_2310 ();
 sg13g2_decap_8 FILLER_25_2317 ();
 sg13g2_decap_8 FILLER_25_2324 ();
 sg13g2_decap_8 FILLER_25_2331 ();
 sg13g2_decap_8 FILLER_25_2338 ();
 sg13g2_decap_8 FILLER_25_2345 ();
 sg13g2_decap_8 FILLER_25_2352 ();
 sg13g2_decap_8 FILLER_25_2359 ();
 sg13g2_decap_8 FILLER_25_2366 ();
 sg13g2_decap_8 FILLER_25_2373 ();
 sg13g2_decap_8 FILLER_25_2380 ();
 sg13g2_decap_8 FILLER_25_2387 ();
 sg13g2_decap_8 FILLER_25_2394 ();
 sg13g2_decap_8 FILLER_25_2401 ();
 sg13g2_decap_8 FILLER_25_2408 ();
 sg13g2_decap_8 FILLER_25_2415 ();
 sg13g2_decap_8 FILLER_25_2422 ();
 sg13g2_decap_8 FILLER_25_2429 ();
 sg13g2_decap_8 FILLER_25_2436 ();
 sg13g2_decap_8 FILLER_25_2443 ();
 sg13g2_decap_8 FILLER_25_2450 ();
 sg13g2_decap_8 FILLER_25_2457 ();
 sg13g2_decap_8 FILLER_25_2464 ();
 sg13g2_decap_8 FILLER_25_2471 ();
 sg13g2_decap_8 FILLER_25_2478 ();
 sg13g2_decap_8 FILLER_25_2485 ();
 sg13g2_decap_8 FILLER_25_2492 ();
 sg13g2_decap_8 FILLER_25_2499 ();
 sg13g2_decap_8 FILLER_25_2506 ();
 sg13g2_decap_8 FILLER_25_2513 ();
 sg13g2_decap_8 FILLER_25_2520 ();
 sg13g2_decap_8 FILLER_25_2527 ();
 sg13g2_decap_8 FILLER_25_2534 ();
 sg13g2_decap_8 FILLER_25_2541 ();
 sg13g2_decap_8 FILLER_25_2548 ();
 sg13g2_decap_8 FILLER_25_2555 ();
 sg13g2_decap_8 FILLER_25_2562 ();
 sg13g2_decap_8 FILLER_25_2569 ();
 sg13g2_decap_8 FILLER_25_2576 ();
 sg13g2_decap_8 FILLER_25_2583 ();
 sg13g2_decap_8 FILLER_25_2590 ();
 sg13g2_decap_8 FILLER_25_2597 ();
 sg13g2_decap_8 FILLER_25_2604 ();
 sg13g2_decap_8 FILLER_25_2611 ();
 sg13g2_decap_8 FILLER_25_2618 ();
 sg13g2_decap_8 FILLER_25_2625 ();
 sg13g2_decap_8 FILLER_25_2632 ();
 sg13g2_decap_8 FILLER_25_2639 ();
 sg13g2_decap_8 FILLER_25_2646 ();
 sg13g2_decap_8 FILLER_25_2653 ();
 sg13g2_decap_8 FILLER_25_2660 ();
 sg13g2_decap_8 FILLER_25_2667 ();
 sg13g2_decap_8 FILLER_25_2674 ();
 sg13g2_decap_8 FILLER_25_2681 ();
 sg13g2_decap_8 FILLER_25_2688 ();
 sg13g2_decap_8 FILLER_25_2695 ();
 sg13g2_decap_8 FILLER_25_2702 ();
 sg13g2_decap_8 FILLER_25_2709 ();
 sg13g2_decap_8 FILLER_25_2716 ();
 sg13g2_decap_8 FILLER_25_2723 ();
 sg13g2_decap_8 FILLER_25_2730 ();
 sg13g2_decap_8 FILLER_25_2737 ();
 sg13g2_decap_8 FILLER_25_2744 ();
 sg13g2_decap_8 FILLER_25_2751 ();
 sg13g2_decap_8 FILLER_25_2758 ();
 sg13g2_decap_8 FILLER_25_2765 ();
 sg13g2_decap_8 FILLER_25_2772 ();
 sg13g2_decap_8 FILLER_25_2779 ();
 sg13g2_decap_8 FILLER_25_2786 ();
 sg13g2_decap_8 FILLER_25_2793 ();
 sg13g2_decap_8 FILLER_25_2800 ();
 sg13g2_decap_8 FILLER_25_2807 ();
 sg13g2_decap_8 FILLER_25_2814 ();
 sg13g2_decap_8 FILLER_25_2821 ();
 sg13g2_decap_8 FILLER_25_2828 ();
 sg13g2_decap_8 FILLER_25_2835 ();
 sg13g2_decap_8 FILLER_25_2842 ();
 sg13g2_decap_8 FILLER_25_2849 ();
 sg13g2_decap_8 FILLER_25_2856 ();
 sg13g2_decap_8 FILLER_25_2863 ();
 sg13g2_decap_8 FILLER_25_2870 ();
 sg13g2_decap_8 FILLER_25_2877 ();
 sg13g2_decap_8 FILLER_25_2884 ();
 sg13g2_decap_8 FILLER_25_2891 ();
 sg13g2_decap_8 FILLER_25_2898 ();
 sg13g2_decap_8 FILLER_25_2905 ();
 sg13g2_decap_8 FILLER_25_2912 ();
 sg13g2_decap_8 FILLER_25_2919 ();
 sg13g2_decap_8 FILLER_25_2926 ();
 sg13g2_decap_8 FILLER_25_2933 ();
 sg13g2_decap_8 FILLER_25_2940 ();
 sg13g2_decap_8 FILLER_25_2947 ();
 sg13g2_decap_8 FILLER_25_2954 ();
 sg13g2_decap_8 FILLER_25_2961 ();
 sg13g2_decap_8 FILLER_25_2968 ();
 sg13g2_decap_8 FILLER_25_2975 ();
 sg13g2_decap_8 FILLER_25_2982 ();
 sg13g2_decap_8 FILLER_25_2989 ();
 sg13g2_decap_8 FILLER_25_2996 ();
 sg13g2_decap_8 FILLER_25_3003 ();
 sg13g2_decap_8 FILLER_25_3010 ();
 sg13g2_decap_8 FILLER_25_3017 ();
 sg13g2_decap_8 FILLER_25_3024 ();
 sg13g2_decap_8 FILLER_25_3031 ();
 sg13g2_decap_8 FILLER_25_3038 ();
 sg13g2_decap_8 FILLER_25_3045 ();
 sg13g2_decap_8 FILLER_25_3052 ();
 sg13g2_decap_8 FILLER_25_3059 ();
 sg13g2_decap_8 FILLER_25_3066 ();
 sg13g2_decap_8 FILLER_25_3073 ();
 sg13g2_decap_8 FILLER_25_3080 ();
 sg13g2_decap_8 FILLER_25_3087 ();
 sg13g2_decap_8 FILLER_25_3094 ();
 sg13g2_decap_8 FILLER_25_3101 ();
 sg13g2_decap_8 FILLER_25_3108 ();
 sg13g2_decap_8 FILLER_25_3115 ();
 sg13g2_decap_8 FILLER_25_3122 ();
 sg13g2_decap_8 FILLER_25_3129 ();
 sg13g2_decap_8 FILLER_25_3136 ();
 sg13g2_decap_8 FILLER_25_3143 ();
 sg13g2_decap_8 FILLER_25_3150 ();
 sg13g2_decap_8 FILLER_25_3157 ();
 sg13g2_decap_8 FILLER_25_3164 ();
 sg13g2_decap_8 FILLER_25_3171 ();
 sg13g2_decap_8 FILLER_25_3178 ();
 sg13g2_decap_8 FILLER_25_3185 ();
 sg13g2_decap_8 FILLER_25_3192 ();
 sg13g2_decap_8 FILLER_25_3199 ();
 sg13g2_decap_8 FILLER_25_3206 ();
 sg13g2_decap_8 FILLER_25_3213 ();
 sg13g2_decap_8 FILLER_25_3220 ();
 sg13g2_decap_8 FILLER_25_3227 ();
 sg13g2_decap_8 FILLER_25_3234 ();
 sg13g2_decap_8 FILLER_25_3241 ();
 sg13g2_decap_8 FILLER_25_3248 ();
 sg13g2_decap_8 FILLER_25_3255 ();
 sg13g2_decap_8 FILLER_25_3262 ();
 sg13g2_decap_8 FILLER_25_3269 ();
 sg13g2_decap_8 FILLER_25_3276 ();
 sg13g2_decap_8 FILLER_25_3283 ();
 sg13g2_decap_8 FILLER_25_3290 ();
 sg13g2_decap_8 FILLER_25_3297 ();
 sg13g2_decap_8 FILLER_25_3304 ();
 sg13g2_decap_8 FILLER_25_3311 ();
 sg13g2_decap_8 FILLER_25_3318 ();
 sg13g2_decap_8 FILLER_25_3325 ();
 sg13g2_decap_8 FILLER_25_3332 ();
 sg13g2_decap_8 FILLER_25_3339 ();
 sg13g2_decap_8 FILLER_25_3346 ();
 sg13g2_decap_8 FILLER_25_3353 ();
 sg13g2_decap_8 FILLER_25_3360 ();
 sg13g2_decap_8 FILLER_25_3367 ();
 sg13g2_decap_8 FILLER_25_3374 ();
 sg13g2_decap_8 FILLER_25_3381 ();
 sg13g2_decap_8 FILLER_25_3388 ();
 sg13g2_decap_8 FILLER_25_3395 ();
 sg13g2_decap_8 FILLER_25_3402 ();
 sg13g2_decap_8 FILLER_25_3409 ();
 sg13g2_decap_8 FILLER_25_3416 ();
 sg13g2_decap_8 FILLER_25_3423 ();
 sg13g2_decap_8 FILLER_25_3430 ();
 sg13g2_decap_8 FILLER_25_3437 ();
 sg13g2_decap_8 FILLER_25_3444 ();
 sg13g2_decap_8 FILLER_25_3451 ();
 sg13g2_decap_8 FILLER_25_3458 ();
 sg13g2_decap_8 FILLER_25_3465 ();
 sg13g2_decap_8 FILLER_25_3472 ();
 sg13g2_decap_8 FILLER_25_3479 ();
 sg13g2_decap_8 FILLER_25_3486 ();
 sg13g2_decap_8 FILLER_25_3493 ();
 sg13g2_decap_8 FILLER_25_3500 ();
 sg13g2_decap_8 FILLER_25_3507 ();
 sg13g2_decap_8 FILLER_25_3514 ();
 sg13g2_decap_8 FILLER_25_3521 ();
 sg13g2_decap_8 FILLER_25_3528 ();
 sg13g2_decap_8 FILLER_25_3535 ();
 sg13g2_decap_8 FILLER_25_3542 ();
 sg13g2_decap_8 FILLER_25_3549 ();
 sg13g2_decap_8 FILLER_25_3556 ();
 sg13g2_decap_8 FILLER_25_3563 ();
 sg13g2_decap_8 FILLER_25_3570 ();
 sg13g2_fill_2 FILLER_25_3577 ();
 sg13g2_fill_1 FILLER_25_3579 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_329 ();
 sg13g2_decap_8 FILLER_26_336 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_8 FILLER_26_357 ();
 sg13g2_decap_8 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_decap_8 FILLER_26_406 ();
 sg13g2_decap_8 FILLER_26_413 ();
 sg13g2_decap_8 FILLER_26_420 ();
 sg13g2_decap_8 FILLER_26_427 ();
 sg13g2_decap_8 FILLER_26_434 ();
 sg13g2_decap_8 FILLER_26_441 ();
 sg13g2_decap_8 FILLER_26_448 ();
 sg13g2_decap_8 FILLER_26_455 ();
 sg13g2_decap_8 FILLER_26_462 ();
 sg13g2_decap_8 FILLER_26_469 ();
 sg13g2_decap_8 FILLER_26_476 ();
 sg13g2_decap_8 FILLER_26_483 ();
 sg13g2_decap_8 FILLER_26_490 ();
 sg13g2_decap_8 FILLER_26_497 ();
 sg13g2_decap_8 FILLER_26_504 ();
 sg13g2_decap_8 FILLER_26_511 ();
 sg13g2_decap_8 FILLER_26_518 ();
 sg13g2_decap_8 FILLER_26_525 ();
 sg13g2_decap_8 FILLER_26_532 ();
 sg13g2_decap_8 FILLER_26_539 ();
 sg13g2_decap_8 FILLER_26_546 ();
 sg13g2_decap_8 FILLER_26_553 ();
 sg13g2_decap_8 FILLER_26_560 ();
 sg13g2_decap_8 FILLER_26_567 ();
 sg13g2_decap_8 FILLER_26_574 ();
 sg13g2_decap_8 FILLER_26_581 ();
 sg13g2_decap_8 FILLER_26_588 ();
 sg13g2_decap_8 FILLER_26_595 ();
 sg13g2_decap_8 FILLER_26_602 ();
 sg13g2_decap_8 FILLER_26_609 ();
 sg13g2_decap_8 FILLER_26_616 ();
 sg13g2_decap_8 FILLER_26_623 ();
 sg13g2_decap_8 FILLER_26_630 ();
 sg13g2_decap_8 FILLER_26_637 ();
 sg13g2_decap_8 FILLER_26_644 ();
 sg13g2_decap_8 FILLER_26_651 ();
 sg13g2_decap_8 FILLER_26_658 ();
 sg13g2_decap_8 FILLER_26_665 ();
 sg13g2_decap_8 FILLER_26_672 ();
 sg13g2_decap_8 FILLER_26_679 ();
 sg13g2_decap_8 FILLER_26_686 ();
 sg13g2_decap_8 FILLER_26_693 ();
 sg13g2_decap_8 FILLER_26_700 ();
 sg13g2_decap_8 FILLER_26_707 ();
 sg13g2_decap_8 FILLER_26_714 ();
 sg13g2_decap_8 FILLER_26_721 ();
 sg13g2_decap_8 FILLER_26_728 ();
 sg13g2_decap_8 FILLER_26_735 ();
 sg13g2_decap_8 FILLER_26_742 ();
 sg13g2_decap_8 FILLER_26_749 ();
 sg13g2_decap_8 FILLER_26_756 ();
 sg13g2_decap_8 FILLER_26_763 ();
 sg13g2_decap_8 FILLER_26_770 ();
 sg13g2_decap_8 FILLER_26_777 ();
 sg13g2_decap_8 FILLER_26_784 ();
 sg13g2_decap_8 FILLER_26_791 ();
 sg13g2_decap_8 FILLER_26_798 ();
 sg13g2_decap_8 FILLER_26_805 ();
 sg13g2_decap_8 FILLER_26_812 ();
 sg13g2_decap_8 FILLER_26_819 ();
 sg13g2_decap_8 FILLER_26_826 ();
 sg13g2_decap_8 FILLER_26_833 ();
 sg13g2_decap_8 FILLER_26_840 ();
 sg13g2_decap_8 FILLER_26_847 ();
 sg13g2_decap_8 FILLER_26_854 ();
 sg13g2_decap_8 FILLER_26_861 ();
 sg13g2_decap_8 FILLER_26_868 ();
 sg13g2_decap_8 FILLER_26_875 ();
 sg13g2_decap_8 FILLER_26_882 ();
 sg13g2_decap_8 FILLER_26_889 ();
 sg13g2_decap_8 FILLER_26_896 ();
 sg13g2_decap_8 FILLER_26_903 ();
 sg13g2_decap_8 FILLER_26_910 ();
 sg13g2_decap_8 FILLER_26_917 ();
 sg13g2_decap_8 FILLER_26_924 ();
 sg13g2_decap_8 FILLER_26_931 ();
 sg13g2_decap_8 FILLER_26_938 ();
 sg13g2_decap_8 FILLER_26_945 ();
 sg13g2_decap_8 FILLER_26_952 ();
 sg13g2_decap_8 FILLER_26_959 ();
 sg13g2_decap_8 FILLER_26_966 ();
 sg13g2_decap_8 FILLER_26_973 ();
 sg13g2_decap_8 FILLER_26_980 ();
 sg13g2_decap_8 FILLER_26_987 ();
 sg13g2_decap_8 FILLER_26_994 ();
 sg13g2_decap_8 FILLER_26_1001 ();
 sg13g2_decap_8 FILLER_26_1008 ();
 sg13g2_decap_8 FILLER_26_1015 ();
 sg13g2_decap_8 FILLER_26_1022 ();
 sg13g2_decap_8 FILLER_26_1029 ();
 sg13g2_decap_8 FILLER_26_1036 ();
 sg13g2_decap_8 FILLER_26_1043 ();
 sg13g2_decap_8 FILLER_26_1050 ();
 sg13g2_decap_8 FILLER_26_1057 ();
 sg13g2_decap_8 FILLER_26_1064 ();
 sg13g2_decap_8 FILLER_26_1071 ();
 sg13g2_decap_8 FILLER_26_1078 ();
 sg13g2_decap_8 FILLER_26_1085 ();
 sg13g2_decap_8 FILLER_26_1092 ();
 sg13g2_decap_8 FILLER_26_1099 ();
 sg13g2_decap_8 FILLER_26_1106 ();
 sg13g2_decap_8 FILLER_26_1113 ();
 sg13g2_decap_8 FILLER_26_1120 ();
 sg13g2_decap_8 FILLER_26_1127 ();
 sg13g2_decap_8 FILLER_26_1134 ();
 sg13g2_decap_8 FILLER_26_1141 ();
 sg13g2_decap_8 FILLER_26_1148 ();
 sg13g2_decap_8 FILLER_26_1155 ();
 sg13g2_decap_8 FILLER_26_1162 ();
 sg13g2_decap_8 FILLER_26_1169 ();
 sg13g2_decap_8 FILLER_26_1176 ();
 sg13g2_decap_8 FILLER_26_1183 ();
 sg13g2_decap_8 FILLER_26_1190 ();
 sg13g2_decap_8 FILLER_26_1197 ();
 sg13g2_decap_8 FILLER_26_1204 ();
 sg13g2_decap_8 FILLER_26_1211 ();
 sg13g2_decap_8 FILLER_26_1218 ();
 sg13g2_decap_8 FILLER_26_1225 ();
 sg13g2_decap_8 FILLER_26_1232 ();
 sg13g2_decap_8 FILLER_26_1239 ();
 sg13g2_decap_8 FILLER_26_1246 ();
 sg13g2_decap_8 FILLER_26_1253 ();
 sg13g2_decap_8 FILLER_26_1260 ();
 sg13g2_decap_8 FILLER_26_1267 ();
 sg13g2_decap_8 FILLER_26_1274 ();
 sg13g2_decap_8 FILLER_26_1281 ();
 sg13g2_decap_8 FILLER_26_1288 ();
 sg13g2_decap_8 FILLER_26_1295 ();
 sg13g2_decap_8 FILLER_26_1302 ();
 sg13g2_decap_8 FILLER_26_1309 ();
 sg13g2_decap_8 FILLER_26_1316 ();
 sg13g2_decap_8 FILLER_26_1323 ();
 sg13g2_decap_8 FILLER_26_1330 ();
 sg13g2_decap_8 FILLER_26_1337 ();
 sg13g2_decap_8 FILLER_26_1344 ();
 sg13g2_decap_8 FILLER_26_1351 ();
 sg13g2_decap_8 FILLER_26_1358 ();
 sg13g2_decap_8 FILLER_26_1365 ();
 sg13g2_decap_8 FILLER_26_1372 ();
 sg13g2_decap_8 FILLER_26_1379 ();
 sg13g2_decap_8 FILLER_26_1386 ();
 sg13g2_decap_8 FILLER_26_1393 ();
 sg13g2_decap_8 FILLER_26_1400 ();
 sg13g2_decap_8 FILLER_26_1407 ();
 sg13g2_decap_8 FILLER_26_1414 ();
 sg13g2_decap_8 FILLER_26_1421 ();
 sg13g2_decap_8 FILLER_26_1428 ();
 sg13g2_decap_8 FILLER_26_1435 ();
 sg13g2_decap_8 FILLER_26_1442 ();
 sg13g2_decap_8 FILLER_26_1449 ();
 sg13g2_decap_8 FILLER_26_1456 ();
 sg13g2_decap_8 FILLER_26_1463 ();
 sg13g2_decap_8 FILLER_26_1470 ();
 sg13g2_decap_8 FILLER_26_1477 ();
 sg13g2_decap_8 FILLER_26_1484 ();
 sg13g2_decap_8 FILLER_26_1491 ();
 sg13g2_decap_8 FILLER_26_1498 ();
 sg13g2_decap_8 FILLER_26_1505 ();
 sg13g2_decap_8 FILLER_26_1512 ();
 sg13g2_decap_8 FILLER_26_1519 ();
 sg13g2_decap_8 FILLER_26_1526 ();
 sg13g2_decap_8 FILLER_26_1533 ();
 sg13g2_decap_8 FILLER_26_1540 ();
 sg13g2_decap_8 FILLER_26_1547 ();
 sg13g2_decap_8 FILLER_26_1554 ();
 sg13g2_decap_8 FILLER_26_1561 ();
 sg13g2_decap_8 FILLER_26_1568 ();
 sg13g2_decap_8 FILLER_26_1575 ();
 sg13g2_decap_8 FILLER_26_1582 ();
 sg13g2_decap_8 FILLER_26_1589 ();
 sg13g2_decap_8 FILLER_26_1596 ();
 sg13g2_decap_8 FILLER_26_1603 ();
 sg13g2_decap_8 FILLER_26_1610 ();
 sg13g2_decap_8 FILLER_26_1617 ();
 sg13g2_decap_8 FILLER_26_1624 ();
 sg13g2_decap_8 FILLER_26_1631 ();
 sg13g2_decap_8 FILLER_26_1638 ();
 sg13g2_decap_8 FILLER_26_1645 ();
 sg13g2_decap_8 FILLER_26_1652 ();
 sg13g2_decap_8 FILLER_26_1659 ();
 sg13g2_decap_8 FILLER_26_1666 ();
 sg13g2_decap_8 FILLER_26_1673 ();
 sg13g2_decap_8 FILLER_26_1680 ();
 sg13g2_decap_8 FILLER_26_1687 ();
 sg13g2_decap_8 FILLER_26_1694 ();
 sg13g2_decap_8 FILLER_26_1701 ();
 sg13g2_decap_8 FILLER_26_1708 ();
 sg13g2_decap_8 FILLER_26_1715 ();
 sg13g2_decap_8 FILLER_26_1722 ();
 sg13g2_decap_8 FILLER_26_1729 ();
 sg13g2_decap_8 FILLER_26_1736 ();
 sg13g2_decap_8 FILLER_26_1743 ();
 sg13g2_decap_8 FILLER_26_1750 ();
 sg13g2_decap_8 FILLER_26_1757 ();
 sg13g2_decap_8 FILLER_26_1764 ();
 sg13g2_decap_8 FILLER_26_1771 ();
 sg13g2_decap_8 FILLER_26_1778 ();
 sg13g2_decap_8 FILLER_26_1785 ();
 sg13g2_decap_8 FILLER_26_1792 ();
 sg13g2_decap_8 FILLER_26_1799 ();
 sg13g2_decap_8 FILLER_26_1806 ();
 sg13g2_decap_8 FILLER_26_1813 ();
 sg13g2_decap_8 FILLER_26_1820 ();
 sg13g2_decap_8 FILLER_26_1827 ();
 sg13g2_decap_8 FILLER_26_1834 ();
 sg13g2_decap_8 FILLER_26_1841 ();
 sg13g2_decap_8 FILLER_26_1848 ();
 sg13g2_decap_8 FILLER_26_1855 ();
 sg13g2_decap_8 FILLER_26_1862 ();
 sg13g2_decap_8 FILLER_26_1869 ();
 sg13g2_decap_8 FILLER_26_1876 ();
 sg13g2_decap_8 FILLER_26_1883 ();
 sg13g2_decap_8 FILLER_26_1890 ();
 sg13g2_decap_8 FILLER_26_1897 ();
 sg13g2_decap_8 FILLER_26_1904 ();
 sg13g2_decap_8 FILLER_26_1911 ();
 sg13g2_decap_8 FILLER_26_1918 ();
 sg13g2_decap_8 FILLER_26_1925 ();
 sg13g2_decap_8 FILLER_26_1932 ();
 sg13g2_decap_8 FILLER_26_1939 ();
 sg13g2_decap_8 FILLER_26_1946 ();
 sg13g2_decap_8 FILLER_26_1953 ();
 sg13g2_decap_8 FILLER_26_1960 ();
 sg13g2_decap_8 FILLER_26_1967 ();
 sg13g2_decap_8 FILLER_26_1974 ();
 sg13g2_decap_8 FILLER_26_1981 ();
 sg13g2_decap_8 FILLER_26_1988 ();
 sg13g2_decap_8 FILLER_26_1995 ();
 sg13g2_decap_8 FILLER_26_2002 ();
 sg13g2_decap_8 FILLER_26_2009 ();
 sg13g2_decap_8 FILLER_26_2016 ();
 sg13g2_decap_8 FILLER_26_2023 ();
 sg13g2_decap_8 FILLER_26_2030 ();
 sg13g2_decap_8 FILLER_26_2037 ();
 sg13g2_decap_8 FILLER_26_2044 ();
 sg13g2_decap_8 FILLER_26_2051 ();
 sg13g2_decap_8 FILLER_26_2058 ();
 sg13g2_decap_8 FILLER_26_2065 ();
 sg13g2_decap_8 FILLER_26_2072 ();
 sg13g2_decap_8 FILLER_26_2079 ();
 sg13g2_decap_8 FILLER_26_2086 ();
 sg13g2_decap_8 FILLER_26_2093 ();
 sg13g2_decap_8 FILLER_26_2100 ();
 sg13g2_decap_8 FILLER_26_2107 ();
 sg13g2_decap_8 FILLER_26_2114 ();
 sg13g2_decap_8 FILLER_26_2121 ();
 sg13g2_decap_8 FILLER_26_2128 ();
 sg13g2_decap_8 FILLER_26_2135 ();
 sg13g2_decap_8 FILLER_26_2142 ();
 sg13g2_decap_8 FILLER_26_2149 ();
 sg13g2_decap_8 FILLER_26_2156 ();
 sg13g2_decap_8 FILLER_26_2163 ();
 sg13g2_decap_8 FILLER_26_2170 ();
 sg13g2_decap_8 FILLER_26_2177 ();
 sg13g2_decap_8 FILLER_26_2184 ();
 sg13g2_decap_8 FILLER_26_2191 ();
 sg13g2_decap_8 FILLER_26_2198 ();
 sg13g2_decap_8 FILLER_26_2205 ();
 sg13g2_decap_8 FILLER_26_2212 ();
 sg13g2_decap_8 FILLER_26_2219 ();
 sg13g2_decap_8 FILLER_26_2226 ();
 sg13g2_decap_8 FILLER_26_2233 ();
 sg13g2_decap_8 FILLER_26_2240 ();
 sg13g2_decap_8 FILLER_26_2247 ();
 sg13g2_decap_8 FILLER_26_2254 ();
 sg13g2_decap_8 FILLER_26_2261 ();
 sg13g2_decap_8 FILLER_26_2268 ();
 sg13g2_decap_8 FILLER_26_2275 ();
 sg13g2_decap_8 FILLER_26_2282 ();
 sg13g2_decap_8 FILLER_26_2289 ();
 sg13g2_decap_8 FILLER_26_2296 ();
 sg13g2_decap_8 FILLER_26_2303 ();
 sg13g2_decap_8 FILLER_26_2310 ();
 sg13g2_decap_8 FILLER_26_2317 ();
 sg13g2_decap_8 FILLER_26_2324 ();
 sg13g2_decap_8 FILLER_26_2331 ();
 sg13g2_decap_8 FILLER_26_2338 ();
 sg13g2_decap_8 FILLER_26_2345 ();
 sg13g2_decap_8 FILLER_26_2352 ();
 sg13g2_decap_8 FILLER_26_2359 ();
 sg13g2_decap_8 FILLER_26_2366 ();
 sg13g2_decap_8 FILLER_26_2373 ();
 sg13g2_decap_8 FILLER_26_2380 ();
 sg13g2_decap_8 FILLER_26_2387 ();
 sg13g2_decap_8 FILLER_26_2394 ();
 sg13g2_decap_8 FILLER_26_2401 ();
 sg13g2_decap_8 FILLER_26_2408 ();
 sg13g2_decap_8 FILLER_26_2415 ();
 sg13g2_decap_8 FILLER_26_2422 ();
 sg13g2_decap_8 FILLER_26_2429 ();
 sg13g2_decap_8 FILLER_26_2436 ();
 sg13g2_decap_8 FILLER_26_2443 ();
 sg13g2_decap_8 FILLER_26_2450 ();
 sg13g2_decap_8 FILLER_26_2457 ();
 sg13g2_decap_8 FILLER_26_2464 ();
 sg13g2_decap_8 FILLER_26_2471 ();
 sg13g2_decap_8 FILLER_26_2478 ();
 sg13g2_decap_8 FILLER_26_2485 ();
 sg13g2_decap_8 FILLER_26_2492 ();
 sg13g2_decap_8 FILLER_26_2499 ();
 sg13g2_decap_8 FILLER_26_2506 ();
 sg13g2_decap_8 FILLER_26_2513 ();
 sg13g2_decap_8 FILLER_26_2520 ();
 sg13g2_decap_8 FILLER_26_2527 ();
 sg13g2_decap_8 FILLER_26_2534 ();
 sg13g2_decap_8 FILLER_26_2541 ();
 sg13g2_decap_8 FILLER_26_2548 ();
 sg13g2_decap_8 FILLER_26_2555 ();
 sg13g2_decap_8 FILLER_26_2562 ();
 sg13g2_decap_8 FILLER_26_2569 ();
 sg13g2_decap_8 FILLER_26_2576 ();
 sg13g2_decap_8 FILLER_26_2583 ();
 sg13g2_decap_8 FILLER_26_2590 ();
 sg13g2_decap_8 FILLER_26_2597 ();
 sg13g2_decap_8 FILLER_26_2604 ();
 sg13g2_decap_8 FILLER_26_2611 ();
 sg13g2_decap_8 FILLER_26_2618 ();
 sg13g2_decap_8 FILLER_26_2625 ();
 sg13g2_decap_8 FILLER_26_2632 ();
 sg13g2_decap_8 FILLER_26_2639 ();
 sg13g2_decap_8 FILLER_26_2646 ();
 sg13g2_decap_8 FILLER_26_2653 ();
 sg13g2_decap_8 FILLER_26_2660 ();
 sg13g2_decap_8 FILLER_26_2667 ();
 sg13g2_decap_8 FILLER_26_2674 ();
 sg13g2_decap_8 FILLER_26_2681 ();
 sg13g2_decap_8 FILLER_26_2688 ();
 sg13g2_decap_8 FILLER_26_2695 ();
 sg13g2_decap_8 FILLER_26_2702 ();
 sg13g2_decap_8 FILLER_26_2709 ();
 sg13g2_decap_8 FILLER_26_2716 ();
 sg13g2_decap_8 FILLER_26_2723 ();
 sg13g2_decap_8 FILLER_26_2730 ();
 sg13g2_decap_8 FILLER_26_2737 ();
 sg13g2_decap_8 FILLER_26_2744 ();
 sg13g2_decap_8 FILLER_26_2751 ();
 sg13g2_decap_8 FILLER_26_2758 ();
 sg13g2_decap_8 FILLER_26_2765 ();
 sg13g2_decap_8 FILLER_26_2772 ();
 sg13g2_decap_8 FILLER_26_2779 ();
 sg13g2_decap_8 FILLER_26_2786 ();
 sg13g2_decap_8 FILLER_26_2793 ();
 sg13g2_decap_8 FILLER_26_2800 ();
 sg13g2_decap_8 FILLER_26_2807 ();
 sg13g2_decap_8 FILLER_26_2814 ();
 sg13g2_decap_8 FILLER_26_2821 ();
 sg13g2_decap_8 FILLER_26_2828 ();
 sg13g2_decap_8 FILLER_26_2835 ();
 sg13g2_decap_8 FILLER_26_2842 ();
 sg13g2_decap_8 FILLER_26_2849 ();
 sg13g2_decap_8 FILLER_26_2856 ();
 sg13g2_decap_8 FILLER_26_2863 ();
 sg13g2_decap_8 FILLER_26_2870 ();
 sg13g2_decap_8 FILLER_26_2877 ();
 sg13g2_decap_8 FILLER_26_2884 ();
 sg13g2_decap_8 FILLER_26_2891 ();
 sg13g2_decap_8 FILLER_26_2898 ();
 sg13g2_decap_8 FILLER_26_2905 ();
 sg13g2_decap_8 FILLER_26_2912 ();
 sg13g2_decap_8 FILLER_26_2919 ();
 sg13g2_decap_8 FILLER_26_2926 ();
 sg13g2_decap_8 FILLER_26_2933 ();
 sg13g2_decap_8 FILLER_26_2940 ();
 sg13g2_decap_8 FILLER_26_2947 ();
 sg13g2_decap_8 FILLER_26_2954 ();
 sg13g2_decap_8 FILLER_26_2961 ();
 sg13g2_decap_8 FILLER_26_2968 ();
 sg13g2_decap_8 FILLER_26_2975 ();
 sg13g2_decap_8 FILLER_26_2982 ();
 sg13g2_decap_8 FILLER_26_2989 ();
 sg13g2_decap_8 FILLER_26_2996 ();
 sg13g2_decap_8 FILLER_26_3003 ();
 sg13g2_decap_8 FILLER_26_3010 ();
 sg13g2_decap_8 FILLER_26_3017 ();
 sg13g2_decap_8 FILLER_26_3024 ();
 sg13g2_decap_8 FILLER_26_3031 ();
 sg13g2_decap_8 FILLER_26_3038 ();
 sg13g2_decap_8 FILLER_26_3045 ();
 sg13g2_decap_8 FILLER_26_3052 ();
 sg13g2_decap_8 FILLER_26_3059 ();
 sg13g2_decap_8 FILLER_26_3066 ();
 sg13g2_decap_8 FILLER_26_3073 ();
 sg13g2_decap_8 FILLER_26_3080 ();
 sg13g2_decap_8 FILLER_26_3087 ();
 sg13g2_decap_8 FILLER_26_3094 ();
 sg13g2_decap_8 FILLER_26_3101 ();
 sg13g2_decap_8 FILLER_26_3108 ();
 sg13g2_decap_8 FILLER_26_3115 ();
 sg13g2_decap_8 FILLER_26_3122 ();
 sg13g2_decap_8 FILLER_26_3129 ();
 sg13g2_decap_8 FILLER_26_3136 ();
 sg13g2_decap_8 FILLER_26_3143 ();
 sg13g2_decap_8 FILLER_26_3150 ();
 sg13g2_decap_8 FILLER_26_3157 ();
 sg13g2_decap_8 FILLER_26_3164 ();
 sg13g2_decap_8 FILLER_26_3171 ();
 sg13g2_decap_8 FILLER_26_3178 ();
 sg13g2_decap_8 FILLER_26_3185 ();
 sg13g2_decap_8 FILLER_26_3192 ();
 sg13g2_decap_8 FILLER_26_3199 ();
 sg13g2_decap_8 FILLER_26_3206 ();
 sg13g2_decap_8 FILLER_26_3213 ();
 sg13g2_decap_8 FILLER_26_3220 ();
 sg13g2_decap_8 FILLER_26_3227 ();
 sg13g2_decap_8 FILLER_26_3234 ();
 sg13g2_decap_8 FILLER_26_3241 ();
 sg13g2_decap_8 FILLER_26_3248 ();
 sg13g2_decap_8 FILLER_26_3255 ();
 sg13g2_decap_8 FILLER_26_3262 ();
 sg13g2_decap_8 FILLER_26_3269 ();
 sg13g2_decap_8 FILLER_26_3276 ();
 sg13g2_decap_8 FILLER_26_3283 ();
 sg13g2_decap_8 FILLER_26_3290 ();
 sg13g2_decap_8 FILLER_26_3297 ();
 sg13g2_decap_8 FILLER_26_3304 ();
 sg13g2_decap_8 FILLER_26_3311 ();
 sg13g2_decap_8 FILLER_26_3318 ();
 sg13g2_decap_8 FILLER_26_3325 ();
 sg13g2_decap_8 FILLER_26_3332 ();
 sg13g2_decap_8 FILLER_26_3339 ();
 sg13g2_decap_8 FILLER_26_3346 ();
 sg13g2_decap_8 FILLER_26_3353 ();
 sg13g2_decap_8 FILLER_26_3360 ();
 sg13g2_decap_8 FILLER_26_3367 ();
 sg13g2_decap_8 FILLER_26_3374 ();
 sg13g2_decap_8 FILLER_26_3381 ();
 sg13g2_decap_8 FILLER_26_3388 ();
 sg13g2_decap_8 FILLER_26_3395 ();
 sg13g2_decap_8 FILLER_26_3402 ();
 sg13g2_decap_8 FILLER_26_3409 ();
 sg13g2_decap_8 FILLER_26_3416 ();
 sg13g2_decap_8 FILLER_26_3423 ();
 sg13g2_decap_8 FILLER_26_3430 ();
 sg13g2_decap_8 FILLER_26_3437 ();
 sg13g2_decap_8 FILLER_26_3444 ();
 sg13g2_decap_8 FILLER_26_3451 ();
 sg13g2_decap_8 FILLER_26_3458 ();
 sg13g2_decap_8 FILLER_26_3465 ();
 sg13g2_decap_8 FILLER_26_3472 ();
 sg13g2_decap_8 FILLER_26_3479 ();
 sg13g2_decap_8 FILLER_26_3486 ();
 sg13g2_decap_8 FILLER_26_3493 ();
 sg13g2_decap_8 FILLER_26_3500 ();
 sg13g2_decap_8 FILLER_26_3507 ();
 sg13g2_decap_8 FILLER_26_3514 ();
 sg13g2_decap_8 FILLER_26_3521 ();
 sg13g2_decap_8 FILLER_26_3528 ();
 sg13g2_decap_8 FILLER_26_3535 ();
 sg13g2_decap_8 FILLER_26_3542 ();
 sg13g2_decap_8 FILLER_26_3549 ();
 sg13g2_decap_8 FILLER_26_3556 ();
 sg13g2_decap_8 FILLER_26_3563 ();
 sg13g2_decap_8 FILLER_26_3570 ();
 sg13g2_fill_2 FILLER_26_3577 ();
 sg13g2_fill_1 FILLER_26_3579 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_decap_8 FILLER_27_287 ();
 sg13g2_decap_8 FILLER_27_294 ();
 sg13g2_decap_8 FILLER_27_301 ();
 sg13g2_decap_8 FILLER_27_308 ();
 sg13g2_decap_8 FILLER_27_315 ();
 sg13g2_decap_8 FILLER_27_322 ();
 sg13g2_decap_8 FILLER_27_329 ();
 sg13g2_decap_8 FILLER_27_336 ();
 sg13g2_decap_8 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_350 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_decap_8 FILLER_27_406 ();
 sg13g2_decap_8 FILLER_27_413 ();
 sg13g2_decap_8 FILLER_27_420 ();
 sg13g2_decap_8 FILLER_27_427 ();
 sg13g2_decap_8 FILLER_27_434 ();
 sg13g2_decap_8 FILLER_27_441 ();
 sg13g2_decap_8 FILLER_27_448 ();
 sg13g2_decap_8 FILLER_27_455 ();
 sg13g2_decap_8 FILLER_27_462 ();
 sg13g2_decap_8 FILLER_27_469 ();
 sg13g2_decap_8 FILLER_27_476 ();
 sg13g2_decap_8 FILLER_27_483 ();
 sg13g2_decap_8 FILLER_27_490 ();
 sg13g2_decap_8 FILLER_27_497 ();
 sg13g2_decap_8 FILLER_27_504 ();
 sg13g2_decap_8 FILLER_27_511 ();
 sg13g2_decap_8 FILLER_27_518 ();
 sg13g2_decap_8 FILLER_27_525 ();
 sg13g2_decap_8 FILLER_27_532 ();
 sg13g2_decap_8 FILLER_27_539 ();
 sg13g2_decap_8 FILLER_27_546 ();
 sg13g2_decap_8 FILLER_27_553 ();
 sg13g2_decap_8 FILLER_27_560 ();
 sg13g2_decap_8 FILLER_27_567 ();
 sg13g2_decap_8 FILLER_27_574 ();
 sg13g2_decap_8 FILLER_27_581 ();
 sg13g2_decap_8 FILLER_27_588 ();
 sg13g2_decap_8 FILLER_27_595 ();
 sg13g2_decap_8 FILLER_27_602 ();
 sg13g2_decap_8 FILLER_27_609 ();
 sg13g2_decap_8 FILLER_27_616 ();
 sg13g2_decap_8 FILLER_27_623 ();
 sg13g2_decap_8 FILLER_27_630 ();
 sg13g2_decap_8 FILLER_27_637 ();
 sg13g2_decap_8 FILLER_27_644 ();
 sg13g2_decap_8 FILLER_27_651 ();
 sg13g2_decap_8 FILLER_27_658 ();
 sg13g2_decap_8 FILLER_27_665 ();
 sg13g2_decap_8 FILLER_27_672 ();
 sg13g2_decap_8 FILLER_27_679 ();
 sg13g2_decap_8 FILLER_27_686 ();
 sg13g2_decap_8 FILLER_27_693 ();
 sg13g2_decap_8 FILLER_27_700 ();
 sg13g2_decap_8 FILLER_27_707 ();
 sg13g2_decap_8 FILLER_27_714 ();
 sg13g2_decap_8 FILLER_27_721 ();
 sg13g2_decap_8 FILLER_27_728 ();
 sg13g2_decap_8 FILLER_27_735 ();
 sg13g2_decap_8 FILLER_27_742 ();
 sg13g2_decap_8 FILLER_27_749 ();
 sg13g2_decap_8 FILLER_27_756 ();
 sg13g2_decap_8 FILLER_27_763 ();
 sg13g2_decap_8 FILLER_27_770 ();
 sg13g2_decap_8 FILLER_27_777 ();
 sg13g2_decap_8 FILLER_27_784 ();
 sg13g2_decap_8 FILLER_27_791 ();
 sg13g2_decap_8 FILLER_27_798 ();
 sg13g2_decap_8 FILLER_27_805 ();
 sg13g2_decap_8 FILLER_27_812 ();
 sg13g2_decap_8 FILLER_27_819 ();
 sg13g2_decap_8 FILLER_27_826 ();
 sg13g2_decap_8 FILLER_27_833 ();
 sg13g2_decap_8 FILLER_27_840 ();
 sg13g2_decap_8 FILLER_27_847 ();
 sg13g2_decap_8 FILLER_27_854 ();
 sg13g2_decap_8 FILLER_27_861 ();
 sg13g2_decap_8 FILLER_27_868 ();
 sg13g2_decap_8 FILLER_27_875 ();
 sg13g2_decap_8 FILLER_27_882 ();
 sg13g2_decap_8 FILLER_27_889 ();
 sg13g2_decap_8 FILLER_27_896 ();
 sg13g2_decap_8 FILLER_27_903 ();
 sg13g2_decap_8 FILLER_27_910 ();
 sg13g2_decap_8 FILLER_27_917 ();
 sg13g2_decap_8 FILLER_27_924 ();
 sg13g2_decap_8 FILLER_27_931 ();
 sg13g2_decap_8 FILLER_27_938 ();
 sg13g2_decap_8 FILLER_27_945 ();
 sg13g2_decap_8 FILLER_27_952 ();
 sg13g2_decap_8 FILLER_27_959 ();
 sg13g2_decap_8 FILLER_27_966 ();
 sg13g2_decap_8 FILLER_27_973 ();
 sg13g2_decap_8 FILLER_27_980 ();
 sg13g2_decap_8 FILLER_27_987 ();
 sg13g2_decap_8 FILLER_27_994 ();
 sg13g2_decap_8 FILLER_27_1001 ();
 sg13g2_decap_8 FILLER_27_1008 ();
 sg13g2_decap_8 FILLER_27_1015 ();
 sg13g2_decap_8 FILLER_27_1022 ();
 sg13g2_decap_8 FILLER_27_1029 ();
 sg13g2_decap_8 FILLER_27_1036 ();
 sg13g2_decap_8 FILLER_27_1043 ();
 sg13g2_decap_8 FILLER_27_1050 ();
 sg13g2_decap_8 FILLER_27_1057 ();
 sg13g2_decap_8 FILLER_27_1064 ();
 sg13g2_decap_8 FILLER_27_1071 ();
 sg13g2_decap_8 FILLER_27_1078 ();
 sg13g2_decap_8 FILLER_27_1085 ();
 sg13g2_decap_8 FILLER_27_1092 ();
 sg13g2_decap_8 FILLER_27_1099 ();
 sg13g2_decap_8 FILLER_27_1106 ();
 sg13g2_decap_8 FILLER_27_1113 ();
 sg13g2_decap_8 FILLER_27_1120 ();
 sg13g2_decap_8 FILLER_27_1127 ();
 sg13g2_decap_8 FILLER_27_1134 ();
 sg13g2_decap_8 FILLER_27_1141 ();
 sg13g2_decap_8 FILLER_27_1148 ();
 sg13g2_decap_8 FILLER_27_1155 ();
 sg13g2_decap_8 FILLER_27_1162 ();
 sg13g2_decap_8 FILLER_27_1169 ();
 sg13g2_decap_8 FILLER_27_1176 ();
 sg13g2_decap_8 FILLER_27_1183 ();
 sg13g2_decap_8 FILLER_27_1190 ();
 sg13g2_decap_8 FILLER_27_1197 ();
 sg13g2_decap_8 FILLER_27_1204 ();
 sg13g2_decap_8 FILLER_27_1211 ();
 sg13g2_decap_8 FILLER_27_1218 ();
 sg13g2_decap_8 FILLER_27_1225 ();
 sg13g2_decap_8 FILLER_27_1232 ();
 sg13g2_decap_8 FILLER_27_1239 ();
 sg13g2_decap_8 FILLER_27_1246 ();
 sg13g2_decap_8 FILLER_27_1253 ();
 sg13g2_decap_8 FILLER_27_1260 ();
 sg13g2_decap_8 FILLER_27_1267 ();
 sg13g2_decap_8 FILLER_27_1274 ();
 sg13g2_decap_8 FILLER_27_1281 ();
 sg13g2_decap_8 FILLER_27_1288 ();
 sg13g2_decap_8 FILLER_27_1295 ();
 sg13g2_decap_8 FILLER_27_1302 ();
 sg13g2_decap_8 FILLER_27_1309 ();
 sg13g2_decap_8 FILLER_27_1316 ();
 sg13g2_decap_8 FILLER_27_1323 ();
 sg13g2_decap_8 FILLER_27_1330 ();
 sg13g2_decap_8 FILLER_27_1337 ();
 sg13g2_decap_8 FILLER_27_1344 ();
 sg13g2_decap_8 FILLER_27_1351 ();
 sg13g2_decap_8 FILLER_27_1358 ();
 sg13g2_decap_8 FILLER_27_1365 ();
 sg13g2_decap_8 FILLER_27_1372 ();
 sg13g2_decap_8 FILLER_27_1379 ();
 sg13g2_decap_8 FILLER_27_1386 ();
 sg13g2_decap_8 FILLER_27_1393 ();
 sg13g2_decap_8 FILLER_27_1400 ();
 sg13g2_decap_8 FILLER_27_1407 ();
 sg13g2_decap_8 FILLER_27_1414 ();
 sg13g2_decap_8 FILLER_27_1421 ();
 sg13g2_decap_8 FILLER_27_1428 ();
 sg13g2_decap_8 FILLER_27_1435 ();
 sg13g2_decap_8 FILLER_27_1442 ();
 sg13g2_decap_8 FILLER_27_1449 ();
 sg13g2_decap_8 FILLER_27_1456 ();
 sg13g2_decap_8 FILLER_27_1463 ();
 sg13g2_decap_8 FILLER_27_1470 ();
 sg13g2_decap_8 FILLER_27_1477 ();
 sg13g2_decap_8 FILLER_27_1484 ();
 sg13g2_decap_8 FILLER_27_1491 ();
 sg13g2_decap_8 FILLER_27_1498 ();
 sg13g2_decap_8 FILLER_27_1505 ();
 sg13g2_decap_8 FILLER_27_1512 ();
 sg13g2_decap_8 FILLER_27_1519 ();
 sg13g2_decap_8 FILLER_27_1526 ();
 sg13g2_decap_8 FILLER_27_1533 ();
 sg13g2_decap_8 FILLER_27_1540 ();
 sg13g2_decap_8 FILLER_27_1547 ();
 sg13g2_decap_8 FILLER_27_1554 ();
 sg13g2_decap_8 FILLER_27_1561 ();
 sg13g2_decap_8 FILLER_27_1568 ();
 sg13g2_decap_8 FILLER_27_1575 ();
 sg13g2_decap_8 FILLER_27_1582 ();
 sg13g2_decap_8 FILLER_27_1589 ();
 sg13g2_decap_8 FILLER_27_1596 ();
 sg13g2_decap_8 FILLER_27_1603 ();
 sg13g2_decap_8 FILLER_27_1610 ();
 sg13g2_decap_8 FILLER_27_1617 ();
 sg13g2_decap_8 FILLER_27_1624 ();
 sg13g2_decap_8 FILLER_27_1631 ();
 sg13g2_decap_8 FILLER_27_1638 ();
 sg13g2_decap_8 FILLER_27_1645 ();
 sg13g2_decap_8 FILLER_27_1652 ();
 sg13g2_decap_8 FILLER_27_1659 ();
 sg13g2_decap_8 FILLER_27_1666 ();
 sg13g2_decap_8 FILLER_27_1673 ();
 sg13g2_decap_8 FILLER_27_1680 ();
 sg13g2_decap_8 FILLER_27_1687 ();
 sg13g2_decap_8 FILLER_27_1694 ();
 sg13g2_decap_8 FILLER_27_1701 ();
 sg13g2_decap_8 FILLER_27_1708 ();
 sg13g2_decap_8 FILLER_27_1715 ();
 sg13g2_decap_8 FILLER_27_1722 ();
 sg13g2_decap_8 FILLER_27_1729 ();
 sg13g2_decap_8 FILLER_27_1736 ();
 sg13g2_decap_8 FILLER_27_1743 ();
 sg13g2_decap_8 FILLER_27_1750 ();
 sg13g2_decap_8 FILLER_27_1757 ();
 sg13g2_decap_8 FILLER_27_1764 ();
 sg13g2_decap_8 FILLER_27_1771 ();
 sg13g2_decap_8 FILLER_27_1778 ();
 sg13g2_decap_8 FILLER_27_1785 ();
 sg13g2_decap_8 FILLER_27_1792 ();
 sg13g2_decap_8 FILLER_27_1799 ();
 sg13g2_decap_8 FILLER_27_1806 ();
 sg13g2_decap_8 FILLER_27_1813 ();
 sg13g2_decap_8 FILLER_27_1820 ();
 sg13g2_decap_8 FILLER_27_1827 ();
 sg13g2_decap_8 FILLER_27_1834 ();
 sg13g2_decap_8 FILLER_27_1841 ();
 sg13g2_decap_8 FILLER_27_1848 ();
 sg13g2_decap_8 FILLER_27_1855 ();
 sg13g2_decap_8 FILLER_27_1862 ();
 sg13g2_decap_8 FILLER_27_1869 ();
 sg13g2_decap_8 FILLER_27_1876 ();
 sg13g2_decap_8 FILLER_27_1883 ();
 sg13g2_decap_8 FILLER_27_1890 ();
 sg13g2_decap_8 FILLER_27_1897 ();
 sg13g2_decap_8 FILLER_27_1904 ();
 sg13g2_decap_8 FILLER_27_1911 ();
 sg13g2_decap_8 FILLER_27_1918 ();
 sg13g2_decap_8 FILLER_27_1925 ();
 sg13g2_decap_8 FILLER_27_1932 ();
 sg13g2_decap_8 FILLER_27_1939 ();
 sg13g2_decap_8 FILLER_27_1946 ();
 sg13g2_decap_8 FILLER_27_1953 ();
 sg13g2_decap_8 FILLER_27_1960 ();
 sg13g2_decap_8 FILLER_27_1967 ();
 sg13g2_decap_8 FILLER_27_1974 ();
 sg13g2_decap_8 FILLER_27_1981 ();
 sg13g2_decap_8 FILLER_27_1988 ();
 sg13g2_decap_8 FILLER_27_1995 ();
 sg13g2_decap_8 FILLER_27_2002 ();
 sg13g2_decap_8 FILLER_27_2009 ();
 sg13g2_decap_8 FILLER_27_2016 ();
 sg13g2_decap_8 FILLER_27_2023 ();
 sg13g2_decap_8 FILLER_27_2030 ();
 sg13g2_decap_8 FILLER_27_2037 ();
 sg13g2_decap_8 FILLER_27_2044 ();
 sg13g2_decap_8 FILLER_27_2051 ();
 sg13g2_decap_8 FILLER_27_2058 ();
 sg13g2_decap_8 FILLER_27_2065 ();
 sg13g2_decap_8 FILLER_27_2072 ();
 sg13g2_decap_8 FILLER_27_2079 ();
 sg13g2_decap_8 FILLER_27_2086 ();
 sg13g2_decap_8 FILLER_27_2093 ();
 sg13g2_decap_8 FILLER_27_2100 ();
 sg13g2_decap_8 FILLER_27_2107 ();
 sg13g2_decap_8 FILLER_27_2114 ();
 sg13g2_decap_8 FILLER_27_2121 ();
 sg13g2_decap_8 FILLER_27_2128 ();
 sg13g2_decap_8 FILLER_27_2135 ();
 sg13g2_decap_8 FILLER_27_2142 ();
 sg13g2_decap_8 FILLER_27_2149 ();
 sg13g2_decap_8 FILLER_27_2156 ();
 sg13g2_decap_8 FILLER_27_2163 ();
 sg13g2_decap_8 FILLER_27_2170 ();
 sg13g2_decap_8 FILLER_27_2177 ();
 sg13g2_decap_8 FILLER_27_2184 ();
 sg13g2_decap_8 FILLER_27_2191 ();
 sg13g2_decap_8 FILLER_27_2198 ();
 sg13g2_decap_8 FILLER_27_2205 ();
 sg13g2_decap_8 FILLER_27_2212 ();
 sg13g2_decap_8 FILLER_27_2219 ();
 sg13g2_decap_8 FILLER_27_2226 ();
 sg13g2_decap_8 FILLER_27_2233 ();
 sg13g2_decap_8 FILLER_27_2240 ();
 sg13g2_decap_8 FILLER_27_2247 ();
 sg13g2_decap_8 FILLER_27_2254 ();
 sg13g2_decap_8 FILLER_27_2261 ();
 sg13g2_decap_8 FILLER_27_2268 ();
 sg13g2_decap_8 FILLER_27_2275 ();
 sg13g2_decap_8 FILLER_27_2282 ();
 sg13g2_decap_8 FILLER_27_2289 ();
 sg13g2_decap_8 FILLER_27_2296 ();
 sg13g2_decap_8 FILLER_27_2303 ();
 sg13g2_decap_8 FILLER_27_2310 ();
 sg13g2_decap_8 FILLER_27_2317 ();
 sg13g2_decap_8 FILLER_27_2324 ();
 sg13g2_decap_8 FILLER_27_2331 ();
 sg13g2_decap_8 FILLER_27_2338 ();
 sg13g2_decap_8 FILLER_27_2345 ();
 sg13g2_decap_8 FILLER_27_2352 ();
 sg13g2_decap_8 FILLER_27_2359 ();
 sg13g2_decap_8 FILLER_27_2366 ();
 sg13g2_decap_8 FILLER_27_2373 ();
 sg13g2_decap_8 FILLER_27_2380 ();
 sg13g2_decap_8 FILLER_27_2387 ();
 sg13g2_decap_8 FILLER_27_2394 ();
 sg13g2_decap_8 FILLER_27_2401 ();
 sg13g2_decap_8 FILLER_27_2408 ();
 sg13g2_decap_8 FILLER_27_2415 ();
 sg13g2_decap_8 FILLER_27_2422 ();
 sg13g2_decap_8 FILLER_27_2429 ();
 sg13g2_decap_8 FILLER_27_2436 ();
 sg13g2_decap_8 FILLER_27_2443 ();
 sg13g2_decap_8 FILLER_27_2450 ();
 sg13g2_decap_8 FILLER_27_2457 ();
 sg13g2_decap_8 FILLER_27_2464 ();
 sg13g2_decap_8 FILLER_27_2471 ();
 sg13g2_decap_8 FILLER_27_2478 ();
 sg13g2_decap_8 FILLER_27_2485 ();
 sg13g2_decap_8 FILLER_27_2492 ();
 sg13g2_decap_8 FILLER_27_2499 ();
 sg13g2_decap_8 FILLER_27_2506 ();
 sg13g2_decap_8 FILLER_27_2513 ();
 sg13g2_decap_8 FILLER_27_2520 ();
 sg13g2_decap_8 FILLER_27_2527 ();
 sg13g2_decap_8 FILLER_27_2534 ();
 sg13g2_decap_8 FILLER_27_2541 ();
 sg13g2_decap_8 FILLER_27_2548 ();
 sg13g2_decap_8 FILLER_27_2555 ();
 sg13g2_decap_8 FILLER_27_2562 ();
 sg13g2_decap_8 FILLER_27_2569 ();
 sg13g2_decap_8 FILLER_27_2576 ();
 sg13g2_decap_8 FILLER_27_2583 ();
 sg13g2_decap_8 FILLER_27_2590 ();
 sg13g2_decap_8 FILLER_27_2597 ();
 sg13g2_decap_8 FILLER_27_2604 ();
 sg13g2_decap_8 FILLER_27_2611 ();
 sg13g2_decap_8 FILLER_27_2618 ();
 sg13g2_decap_8 FILLER_27_2625 ();
 sg13g2_decap_8 FILLER_27_2632 ();
 sg13g2_decap_8 FILLER_27_2639 ();
 sg13g2_decap_8 FILLER_27_2646 ();
 sg13g2_decap_8 FILLER_27_2653 ();
 sg13g2_decap_8 FILLER_27_2660 ();
 sg13g2_decap_8 FILLER_27_2667 ();
 sg13g2_decap_8 FILLER_27_2674 ();
 sg13g2_decap_8 FILLER_27_2681 ();
 sg13g2_decap_8 FILLER_27_2688 ();
 sg13g2_decap_8 FILLER_27_2695 ();
 sg13g2_decap_8 FILLER_27_2702 ();
 sg13g2_decap_8 FILLER_27_2709 ();
 sg13g2_decap_8 FILLER_27_2716 ();
 sg13g2_decap_8 FILLER_27_2723 ();
 sg13g2_decap_8 FILLER_27_2730 ();
 sg13g2_decap_8 FILLER_27_2737 ();
 sg13g2_decap_8 FILLER_27_2744 ();
 sg13g2_decap_8 FILLER_27_2751 ();
 sg13g2_decap_8 FILLER_27_2758 ();
 sg13g2_decap_8 FILLER_27_2765 ();
 sg13g2_decap_8 FILLER_27_2772 ();
 sg13g2_decap_8 FILLER_27_2779 ();
 sg13g2_decap_8 FILLER_27_2786 ();
 sg13g2_decap_8 FILLER_27_2793 ();
 sg13g2_decap_8 FILLER_27_2800 ();
 sg13g2_decap_8 FILLER_27_2807 ();
 sg13g2_decap_8 FILLER_27_2814 ();
 sg13g2_decap_8 FILLER_27_2821 ();
 sg13g2_decap_8 FILLER_27_2828 ();
 sg13g2_decap_8 FILLER_27_2835 ();
 sg13g2_decap_8 FILLER_27_2842 ();
 sg13g2_decap_8 FILLER_27_2849 ();
 sg13g2_decap_8 FILLER_27_2856 ();
 sg13g2_decap_8 FILLER_27_2863 ();
 sg13g2_decap_8 FILLER_27_2870 ();
 sg13g2_decap_8 FILLER_27_2877 ();
 sg13g2_decap_8 FILLER_27_2884 ();
 sg13g2_decap_8 FILLER_27_2891 ();
 sg13g2_decap_8 FILLER_27_2898 ();
 sg13g2_decap_8 FILLER_27_2905 ();
 sg13g2_decap_8 FILLER_27_2912 ();
 sg13g2_decap_8 FILLER_27_2919 ();
 sg13g2_decap_8 FILLER_27_2926 ();
 sg13g2_decap_8 FILLER_27_2933 ();
 sg13g2_decap_8 FILLER_27_2940 ();
 sg13g2_decap_8 FILLER_27_2947 ();
 sg13g2_decap_8 FILLER_27_2954 ();
 sg13g2_decap_8 FILLER_27_2961 ();
 sg13g2_decap_8 FILLER_27_2968 ();
 sg13g2_decap_8 FILLER_27_2975 ();
 sg13g2_decap_8 FILLER_27_2982 ();
 sg13g2_decap_8 FILLER_27_2989 ();
 sg13g2_decap_8 FILLER_27_2996 ();
 sg13g2_decap_8 FILLER_27_3003 ();
 sg13g2_decap_8 FILLER_27_3010 ();
 sg13g2_decap_8 FILLER_27_3017 ();
 sg13g2_decap_8 FILLER_27_3024 ();
 sg13g2_decap_8 FILLER_27_3031 ();
 sg13g2_decap_8 FILLER_27_3038 ();
 sg13g2_decap_8 FILLER_27_3045 ();
 sg13g2_decap_8 FILLER_27_3052 ();
 sg13g2_decap_8 FILLER_27_3059 ();
 sg13g2_decap_8 FILLER_27_3066 ();
 sg13g2_decap_8 FILLER_27_3073 ();
 sg13g2_decap_8 FILLER_27_3080 ();
 sg13g2_decap_8 FILLER_27_3087 ();
 sg13g2_decap_8 FILLER_27_3094 ();
 sg13g2_decap_8 FILLER_27_3101 ();
 sg13g2_decap_8 FILLER_27_3108 ();
 sg13g2_decap_8 FILLER_27_3115 ();
 sg13g2_decap_8 FILLER_27_3122 ();
 sg13g2_decap_8 FILLER_27_3129 ();
 sg13g2_decap_8 FILLER_27_3136 ();
 sg13g2_decap_8 FILLER_27_3143 ();
 sg13g2_decap_8 FILLER_27_3150 ();
 sg13g2_decap_8 FILLER_27_3157 ();
 sg13g2_decap_8 FILLER_27_3164 ();
 sg13g2_decap_8 FILLER_27_3171 ();
 sg13g2_decap_8 FILLER_27_3178 ();
 sg13g2_decap_8 FILLER_27_3185 ();
 sg13g2_decap_8 FILLER_27_3192 ();
 sg13g2_decap_8 FILLER_27_3199 ();
 sg13g2_decap_8 FILLER_27_3206 ();
 sg13g2_decap_8 FILLER_27_3213 ();
 sg13g2_decap_8 FILLER_27_3220 ();
 sg13g2_decap_8 FILLER_27_3227 ();
 sg13g2_decap_8 FILLER_27_3234 ();
 sg13g2_decap_8 FILLER_27_3241 ();
 sg13g2_decap_8 FILLER_27_3248 ();
 sg13g2_decap_8 FILLER_27_3255 ();
 sg13g2_decap_8 FILLER_27_3262 ();
 sg13g2_decap_8 FILLER_27_3269 ();
 sg13g2_decap_8 FILLER_27_3276 ();
 sg13g2_decap_8 FILLER_27_3283 ();
 sg13g2_decap_8 FILLER_27_3290 ();
 sg13g2_decap_8 FILLER_27_3297 ();
 sg13g2_decap_8 FILLER_27_3304 ();
 sg13g2_decap_8 FILLER_27_3311 ();
 sg13g2_decap_8 FILLER_27_3318 ();
 sg13g2_decap_8 FILLER_27_3325 ();
 sg13g2_decap_8 FILLER_27_3332 ();
 sg13g2_decap_8 FILLER_27_3339 ();
 sg13g2_decap_8 FILLER_27_3346 ();
 sg13g2_decap_8 FILLER_27_3353 ();
 sg13g2_decap_8 FILLER_27_3360 ();
 sg13g2_decap_8 FILLER_27_3367 ();
 sg13g2_decap_8 FILLER_27_3374 ();
 sg13g2_decap_8 FILLER_27_3381 ();
 sg13g2_decap_8 FILLER_27_3388 ();
 sg13g2_decap_8 FILLER_27_3395 ();
 sg13g2_decap_8 FILLER_27_3402 ();
 sg13g2_decap_8 FILLER_27_3409 ();
 sg13g2_decap_8 FILLER_27_3416 ();
 sg13g2_decap_8 FILLER_27_3423 ();
 sg13g2_decap_8 FILLER_27_3430 ();
 sg13g2_decap_8 FILLER_27_3437 ();
 sg13g2_decap_8 FILLER_27_3444 ();
 sg13g2_decap_8 FILLER_27_3451 ();
 sg13g2_decap_8 FILLER_27_3458 ();
 sg13g2_decap_8 FILLER_27_3465 ();
 sg13g2_decap_8 FILLER_27_3472 ();
 sg13g2_decap_8 FILLER_27_3479 ();
 sg13g2_decap_8 FILLER_27_3486 ();
 sg13g2_decap_8 FILLER_27_3493 ();
 sg13g2_decap_8 FILLER_27_3500 ();
 sg13g2_decap_8 FILLER_27_3507 ();
 sg13g2_decap_8 FILLER_27_3514 ();
 sg13g2_decap_8 FILLER_27_3521 ();
 sg13g2_decap_8 FILLER_27_3528 ();
 sg13g2_decap_8 FILLER_27_3535 ();
 sg13g2_decap_8 FILLER_27_3542 ();
 sg13g2_decap_8 FILLER_27_3549 ();
 sg13g2_decap_8 FILLER_27_3556 ();
 sg13g2_decap_8 FILLER_27_3563 ();
 sg13g2_decap_8 FILLER_27_3570 ();
 sg13g2_fill_2 FILLER_27_3577 ();
 sg13g2_fill_1 FILLER_27_3579 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_8 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_decap_8 FILLER_28_245 ();
 sg13g2_decap_8 FILLER_28_252 ();
 sg13g2_decap_8 FILLER_28_259 ();
 sg13g2_decap_8 FILLER_28_266 ();
 sg13g2_decap_8 FILLER_28_273 ();
 sg13g2_decap_8 FILLER_28_280 ();
 sg13g2_decap_8 FILLER_28_287 ();
 sg13g2_decap_8 FILLER_28_294 ();
 sg13g2_decap_8 FILLER_28_301 ();
 sg13g2_decap_8 FILLER_28_308 ();
 sg13g2_decap_8 FILLER_28_315 ();
 sg13g2_decap_8 FILLER_28_322 ();
 sg13g2_decap_8 FILLER_28_329 ();
 sg13g2_decap_8 FILLER_28_336 ();
 sg13g2_decap_8 FILLER_28_343 ();
 sg13g2_decap_8 FILLER_28_350 ();
 sg13g2_decap_8 FILLER_28_357 ();
 sg13g2_decap_8 FILLER_28_364 ();
 sg13g2_decap_8 FILLER_28_371 ();
 sg13g2_decap_8 FILLER_28_378 ();
 sg13g2_decap_8 FILLER_28_385 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_decap_8 FILLER_28_406 ();
 sg13g2_decap_8 FILLER_28_413 ();
 sg13g2_decap_8 FILLER_28_420 ();
 sg13g2_decap_8 FILLER_28_427 ();
 sg13g2_decap_8 FILLER_28_434 ();
 sg13g2_decap_8 FILLER_28_441 ();
 sg13g2_decap_8 FILLER_28_448 ();
 sg13g2_decap_8 FILLER_28_455 ();
 sg13g2_decap_8 FILLER_28_462 ();
 sg13g2_decap_8 FILLER_28_469 ();
 sg13g2_decap_8 FILLER_28_476 ();
 sg13g2_decap_8 FILLER_28_483 ();
 sg13g2_decap_8 FILLER_28_490 ();
 sg13g2_decap_8 FILLER_28_497 ();
 sg13g2_decap_8 FILLER_28_504 ();
 sg13g2_decap_8 FILLER_28_511 ();
 sg13g2_decap_8 FILLER_28_518 ();
 sg13g2_decap_8 FILLER_28_525 ();
 sg13g2_decap_8 FILLER_28_532 ();
 sg13g2_decap_8 FILLER_28_539 ();
 sg13g2_decap_8 FILLER_28_546 ();
 sg13g2_decap_8 FILLER_28_553 ();
 sg13g2_decap_8 FILLER_28_560 ();
 sg13g2_decap_8 FILLER_28_567 ();
 sg13g2_decap_8 FILLER_28_574 ();
 sg13g2_decap_8 FILLER_28_581 ();
 sg13g2_decap_8 FILLER_28_588 ();
 sg13g2_decap_8 FILLER_28_595 ();
 sg13g2_decap_8 FILLER_28_602 ();
 sg13g2_decap_8 FILLER_28_609 ();
 sg13g2_decap_8 FILLER_28_616 ();
 sg13g2_decap_8 FILLER_28_623 ();
 sg13g2_decap_8 FILLER_28_630 ();
 sg13g2_decap_8 FILLER_28_637 ();
 sg13g2_decap_8 FILLER_28_644 ();
 sg13g2_decap_8 FILLER_28_651 ();
 sg13g2_decap_8 FILLER_28_658 ();
 sg13g2_decap_8 FILLER_28_665 ();
 sg13g2_decap_8 FILLER_28_672 ();
 sg13g2_decap_8 FILLER_28_679 ();
 sg13g2_decap_8 FILLER_28_686 ();
 sg13g2_decap_8 FILLER_28_693 ();
 sg13g2_decap_8 FILLER_28_700 ();
 sg13g2_decap_8 FILLER_28_707 ();
 sg13g2_decap_8 FILLER_28_714 ();
 sg13g2_decap_8 FILLER_28_721 ();
 sg13g2_decap_8 FILLER_28_728 ();
 sg13g2_decap_8 FILLER_28_735 ();
 sg13g2_decap_8 FILLER_28_742 ();
 sg13g2_decap_8 FILLER_28_749 ();
 sg13g2_decap_8 FILLER_28_756 ();
 sg13g2_decap_8 FILLER_28_763 ();
 sg13g2_decap_8 FILLER_28_770 ();
 sg13g2_decap_8 FILLER_28_777 ();
 sg13g2_decap_8 FILLER_28_784 ();
 sg13g2_decap_8 FILLER_28_791 ();
 sg13g2_decap_8 FILLER_28_798 ();
 sg13g2_decap_8 FILLER_28_805 ();
 sg13g2_decap_8 FILLER_28_812 ();
 sg13g2_decap_8 FILLER_28_819 ();
 sg13g2_decap_8 FILLER_28_826 ();
 sg13g2_decap_8 FILLER_28_833 ();
 sg13g2_decap_8 FILLER_28_840 ();
 sg13g2_decap_8 FILLER_28_847 ();
 sg13g2_decap_8 FILLER_28_854 ();
 sg13g2_decap_8 FILLER_28_861 ();
 sg13g2_decap_8 FILLER_28_868 ();
 sg13g2_decap_8 FILLER_28_875 ();
 sg13g2_decap_8 FILLER_28_882 ();
 sg13g2_decap_8 FILLER_28_889 ();
 sg13g2_decap_8 FILLER_28_896 ();
 sg13g2_decap_8 FILLER_28_903 ();
 sg13g2_decap_8 FILLER_28_910 ();
 sg13g2_decap_8 FILLER_28_917 ();
 sg13g2_decap_8 FILLER_28_924 ();
 sg13g2_decap_8 FILLER_28_931 ();
 sg13g2_decap_8 FILLER_28_938 ();
 sg13g2_decap_8 FILLER_28_945 ();
 sg13g2_decap_8 FILLER_28_952 ();
 sg13g2_decap_8 FILLER_28_959 ();
 sg13g2_decap_8 FILLER_28_966 ();
 sg13g2_decap_8 FILLER_28_973 ();
 sg13g2_decap_8 FILLER_28_980 ();
 sg13g2_decap_8 FILLER_28_987 ();
 sg13g2_decap_8 FILLER_28_994 ();
 sg13g2_decap_8 FILLER_28_1001 ();
 sg13g2_decap_8 FILLER_28_1008 ();
 sg13g2_decap_8 FILLER_28_1015 ();
 sg13g2_decap_8 FILLER_28_1022 ();
 sg13g2_decap_8 FILLER_28_1029 ();
 sg13g2_decap_8 FILLER_28_1036 ();
 sg13g2_decap_8 FILLER_28_1043 ();
 sg13g2_decap_8 FILLER_28_1050 ();
 sg13g2_decap_8 FILLER_28_1057 ();
 sg13g2_decap_8 FILLER_28_1064 ();
 sg13g2_decap_8 FILLER_28_1071 ();
 sg13g2_decap_8 FILLER_28_1078 ();
 sg13g2_decap_8 FILLER_28_1085 ();
 sg13g2_decap_8 FILLER_28_1092 ();
 sg13g2_decap_8 FILLER_28_1099 ();
 sg13g2_decap_8 FILLER_28_1106 ();
 sg13g2_decap_8 FILLER_28_1113 ();
 sg13g2_decap_8 FILLER_28_1120 ();
 sg13g2_decap_8 FILLER_28_1127 ();
 sg13g2_decap_8 FILLER_28_1134 ();
 sg13g2_decap_8 FILLER_28_1141 ();
 sg13g2_decap_8 FILLER_28_1148 ();
 sg13g2_decap_8 FILLER_28_1155 ();
 sg13g2_decap_8 FILLER_28_1162 ();
 sg13g2_decap_8 FILLER_28_1169 ();
 sg13g2_decap_8 FILLER_28_1176 ();
 sg13g2_decap_8 FILLER_28_1183 ();
 sg13g2_decap_8 FILLER_28_1190 ();
 sg13g2_decap_8 FILLER_28_1197 ();
 sg13g2_decap_8 FILLER_28_1204 ();
 sg13g2_decap_8 FILLER_28_1211 ();
 sg13g2_decap_8 FILLER_28_1218 ();
 sg13g2_decap_8 FILLER_28_1225 ();
 sg13g2_decap_8 FILLER_28_1232 ();
 sg13g2_decap_8 FILLER_28_1239 ();
 sg13g2_decap_8 FILLER_28_1246 ();
 sg13g2_decap_8 FILLER_28_1253 ();
 sg13g2_decap_8 FILLER_28_1260 ();
 sg13g2_decap_8 FILLER_28_1267 ();
 sg13g2_decap_8 FILLER_28_1274 ();
 sg13g2_decap_8 FILLER_28_1281 ();
 sg13g2_decap_8 FILLER_28_1288 ();
 sg13g2_decap_8 FILLER_28_1295 ();
 sg13g2_decap_8 FILLER_28_1302 ();
 sg13g2_decap_8 FILLER_28_1309 ();
 sg13g2_decap_8 FILLER_28_1316 ();
 sg13g2_decap_8 FILLER_28_1323 ();
 sg13g2_decap_8 FILLER_28_1330 ();
 sg13g2_decap_8 FILLER_28_1337 ();
 sg13g2_decap_8 FILLER_28_1344 ();
 sg13g2_decap_8 FILLER_28_1351 ();
 sg13g2_decap_8 FILLER_28_1358 ();
 sg13g2_decap_8 FILLER_28_1365 ();
 sg13g2_decap_8 FILLER_28_1372 ();
 sg13g2_decap_8 FILLER_28_1379 ();
 sg13g2_decap_8 FILLER_28_1386 ();
 sg13g2_decap_8 FILLER_28_1393 ();
 sg13g2_decap_8 FILLER_28_1400 ();
 sg13g2_decap_8 FILLER_28_1407 ();
 sg13g2_decap_8 FILLER_28_1414 ();
 sg13g2_decap_8 FILLER_28_1421 ();
 sg13g2_decap_8 FILLER_28_1428 ();
 sg13g2_decap_8 FILLER_28_1435 ();
 sg13g2_decap_8 FILLER_28_1442 ();
 sg13g2_decap_8 FILLER_28_1449 ();
 sg13g2_decap_8 FILLER_28_1456 ();
 sg13g2_decap_8 FILLER_28_1463 ();
 sg13g2_decap_8 FILLER_28_1470 ();
 sg13g2_decap_8 FILLER_28_1477 ();
 sg13g2_decap_8 FILLER_28_1484 ();
 sg13g2_decap_8 FILLER_28_1491 ();
 sg13g2_decap_8 FILLER_28_1498 ();
 sg13g2_decap_8 FILLER_28_1505 ();
 sg13g2_decap_8 FILLER_28_1512 ();
 sg13g2_decap_8 FILLER_28_1519 ();
 sg13g2_decap_8 FILLER_28_1526 ();
 sg13g2_decap_8 FILLER_28_1533 ();
 sg13g2_decap_8 FILLER_28_1540 ();
 sg13g2_decap_8 FILLER_28_1547 ();
 sg13g2_decap_8 FILLER_28_1554 ();
 sg13g2_decap_8 FILLER_28_1561 ();
 sg13g2_decap_8 FILLER_28_1568 ();
 sg13g2_decap_8 FILLER_28_1575 ();
 sg13g2_decap_8 FILLER_28_1582 ();
 sg13g2_decap_8 FILLER_28_1589 ();
 sg13g2_decap_8 FILLER_28_1596 ();
 sg13g2_decap_8 FILLER_28_1603 ();
 sg13g2_decap_8 FILLER_28_1610 ();
 sg13g2_decap_8 FILLER_28_1617 ();
 sg13g2_decap_8 FILLER_28_1624 ();
 sg13g2_decap_8 FILLER_28_1631 ();
 sg13g2_decap_8 FILLER_28_1638 ();
 sg13g2_decap_8 FILLER_28_1645 ();
 sg13g2_decap_8 FILLER_28_1652 ();
 sg13g2_decap_8 FILLER_28_1659 ();
 sg13g2_decap_8 FILLER_28_1666 ();
 sg13g2_decap_8 FILLER_28_1673 ();
 sg13g2_decap_8 FILLER_28_1680 ();
 sg13g2_decap_8 FILLER_28_1687 ();
 sg13g2_decap_8 FILLER_28_1694 ();
 sg13g2_decap_8 FILLER_28_1701 ();
 sg13g2_decap_8 FILLER_28_1708 ();
 sg13g2_decap_8 FILLER_28_1715 ();
 sg13g2_decap_8 FILLER_28_1722 ();
 sg13g2_decap_8 FILLER_28_1729 ();
 sg13g2_decap_8 FILLER_28_1736 ();
 sg13g2_decap_8 FILLER_28_1743 ();
 sg13g2_decap_8 FILLER_28_1750 ();
 sg13g2_decap_8 FILLER_28_1757 ();
 sg13g2_decap_8 FILLER_28_1764 ();
 sg13g2_decap_8 FILLER_28_1771 ();
 sg13g2_decap_8 FILLER_28_1778 ();
 sg13g2_decap_8 FILLER_28_1785 ();
 sg13g2_decap_8 FILLER_28_1792 ();
 sg13g2_decap_8 FILLER_28_1799 ();
 sg13g2_decap_8 FILLER_28_1806 ();
 sg13g2_decap_8 FILLER_28_1813 ();
 sg13g2_decap_8 FILLER_28_1820 ();
 sg13g2_decap_8 FILLER_28_1827 ();
 sg13g2_decap_8 FILLER_28_1834 ();
 sg13g2_decap_8 FILLER_28_1841 ();
 sg13g2_decap_8 FILLER_28_1848 ();
 sg13g2_decap_8 FILLER_28_1855 ();
 sg13g2_decap_8 FILLER_28_1862 ();
 sg13g2_decap_8 FILLER_28_1869 ();
 sg13g2_decap_8 FILLER_28_1876 ();
 sg13g2_decap_8 FILLER_28_1883 ();
 sg13g2_decap_8 FILLER_28_1890 ();
 sg13g2_decap_8 FILLER_28_1897 ();
 sg13g2_decap_8 FILLER_28_1904 ();
 sg13g2_decap_8 FILLER_28_1911 ();
 sg13g2_decap_8 FILLER_28_1918 ();
 sg13g2_decap_8 FILLER_28_1925 ();
 sg13g2_decap_8 FILLER_28_1932 ();
 sg13g2_decap_8 FILLER_28_1939 ();
 sg13g2_decap_8 FILLER_28_1946 ();
 sg13g2_decap_8 FILLER_28_1953 ();
 sg13g2_decap_8 FILLER_28_1960 ();
 sg13g2_decap_8 FILLER_28_1967 ();
 sg13g2_decap_8 FILLER_28_1974 ();
 sg13g2_decap_8 FILLER_28_1981 ();
 sg13g2_decap_8 FILLER_28_1988 ();
 sg13g2_decap_8 FILLER_28_1995 ();
 sg13g2_decap_8 FILLER_28_2002 ();
 sg13g2_decap_8 FILLER_28_2009 ();
 sg13g2_decap_8 FILLER_28_2016 ();
 sg13g2_decap_8 FILLER_28_2023 ();
 sg13g2_decap_8 FILLER_28_2030 ();
 sg13g2_decap_8 FILLER_28_2037 ();
 sg13g2_decap_8 FILLER_28_2044 ();
 sg13g2_decap_8 FILLER_28_2051 ();
 sg13g2_decap_8 FILLER_28_2058 ();
 sg13g2_decap_8 FILLER_28_2065 ();
 sg13g2_decap_8 FILLER_28_2072 ();
 sg13g2_decap_8 FILLER_28_2079 ();
 sg13g2_decap_8 FILLER_28_2086 ();
 sg13g2_decap_8 FILLER_28_2093 ();
 sg13g2_decap_8 FILLER_28_2100 ();
 sg13g2_decap_8 FILLER_28_2107 ();
 sg13g2_decap_8 FILLER_28_2114 ();
 sg13g2_decap_8 FILLER_28_2121 ();
 sg13g2_decap_8 FILLER_28_2128 ();
 sg13g2_decap_8 FILLER_28_2135 ();
 sg13g2_decap_8 FILLER_28_2142 ();
 sg13g2_decap_8 FILLER_28_2149 ();
 sg13g2_decap_8 FILLER_28_2156 ();
 sg13g2_decap_8 FILLER_28_2163 ();
 sg13g2_decap_8 FILLER_28_2170 ();
 sg13g2_decap_8 FILLER_28_2177 ();
 sg13g2_decap_8 FILLER_28_2184 ();
 sg13g2_decap_8 FILLER_28_2191 ();
 sg13g2_decap_8 FILLER_28_2198 ();
 sg13g2_decap_8 FILLER_28_2205 ();
 sg13g2_decap_8 FILLER_28_2212 ();
 sg13g2_decap_8 FILLER_28_2219 ();
 sg13g2_decap_8 FILLER_28_2226 ();
 sg13g2_decap_8 FILLER_28_2233 ();
 sg13g2_decap_8 FILLER_28_2240 ();
 sg13g2_decap_8 FILLER_28_2247 ();
 sg13g2_decap_8 FILLER_28_2254 ();
 sg13g2_decap_8 FILLER_28_2261 ();
 sg13g2_decap_8 FILLER_28_2268 ();
 sg13g2_decap_8 FILLER_28_2275 ();
 sg13g2_decap_8 FILLER_28_2282 ();
 sg13g2_decap_8 FILLER_28_2289 ();
 sg13g2_decap_8 FILLER_28_2296 ();
 sg13g2_decap_8 FILLER_28_2303 ();
 sg13g2_decap_8 FILLER_28_2310 ();
 sg13g2_decap_8 FILLER_28_2317 ();
 sg13g2_decap_8 FILLER_28_2324 ();
 sg13g2_decap_8 FILLER_28_2331 ();
 sg13g2_decap_8 FILLER_28_2338 ();
 sg13g2_decap_8 FILLER_28_2345 ();
 sg13g2_decap_8 FILLER_28_2352 ();
 sg13g2_decap_8 FILLER_28_2359 ();
 sg13g2_decap_8 FILLER_28_2366 ();
 sg13g2_decap_8 FILLER_28_2373 ();
 sg13g2_decap_8 FILLER_28_2380 ();
 sg13g2_decap_8 FILLER_28_2387 ();
 sg13g2_decap_8 FILLER_28_2394 ();
 sg13g2_decap_8 FILLER_28_2401 ();
 sg13g2_decap_8 FILLER_28_2408 ();
 sg13g2_decap_8 FILLER_28_2415 ();
 sg13g2_decap_8 FILLER_28_2422 ();
 sg13g2_decap_8 FILLER_28_2429 ();
 sg13g2_decap_8 FILLER_28_2436 ();
 sg13g2_decap_8 FILLER_28_2443 ();
 sg13g2_decap_8 FILLER_28_2450 ();
 sg13g2_decap_8 FILLER_28_2457 ();
 sg13g2_decap_8 FILLER_28_2464 ();
 sg13g2_decap_8 FILLER_28_2471 ();
 sg13g2_decap_8 FILLER_28_2478 ();
 sg13g2_decap_8 FILLER_28_2485 ();
 sg13g2_decap_8 FILLER_28_2492 ();
 sg13g2_decap_8 FILLER_28_2499 ();
 sg13g2_decap_8 FILLER_28_2506 ();
 sg13g2_decap_8 FILLER_28_2513 ();
 sg13g2_decap_8 FILLER_28_2520 ();
 sg13g2_decap_8 FILLER_28_2527 ();
 sg13g2_decap_8 FILLER_28_2534 ();
 sg13g2_decap_8 FILLER_28_2541 ();
 sg13g2_decap_8 FILLER_28_2548 ();
 sg13g2_decap_8 FILLER_28_2555 ();
 sg13g2_decap_8 FILLER_28_2562 ();
 sg13g2_decap_8 FILLER_28_2569 ();
 sg13g2_decap_8 FILLER_28_2576 ();
 sg13g2_decap_8 FILLER_28_2583 ();
 sg13g2_decap_8 FILLER_28_2590 ();
 sg13g2_decap_8 FILLER_28_2597 ();
 sg13g2_decap_8 FILLER_28_2604 ();
 sg13g2_decap_8 FILLER_28_2611 ();
 sg13g2_decap_8 FILLER_28_2618 ();
 sg13g2_decap_8 FILLER_28_2625 ();
 sg13g2_decap_8 FILLER_28_2632 ();
 sg13g2_decap_8 FILLER_28_2639 ();
 sg13g2_decap_8 FILLER_28_2646 ();
 sg13g2_decap_8 FILLER_28_2653 ();
 sg13g2_decap_8 FILLER_28_2660 ();
 sg13g2_decap_8 FILLER_28_2667 ();
 sg13g2_decap_8 FILLER_28_2674 ();
 sg13g2_decap_8 FILLER_28_2681 ();
 sg13g2_decap_8 FILLER_28_2688 ();
 sg13g2_decap_8 FILLER_28_2695 ();
 sg13g2_decap_8 FILLER_28_2702 ();
 sg13g2_decap_8 FILLER_28_2709 ();
 sg13g2_decap_8 FILLER_28_2716 ();
 sg13g2_decap_8 FILLER_28_2723 ();
 sg13g2_decap_8 FILLER_28_2730 ();
 sg13g2_decap_8 FILLER_28_2737 ();
 sg13g2_decap_8 FILLER_28_2744 ();
 sg13g2_decap_8 FILLER_28_2751 ();
 sg13g2_decap_8 FILLER_28_2758 ();
 sg13g2_decap_8 FILLER_28_2765 ();
 sg13g2_decap_8 FILLER_28_2772 ();
 sg13g2_decap_8 FILLER_28_2779 ();
 sg13g2_decap_8 FILLER_28_2786 ();
 sg13g2_decap_8 FILLER_28_2793 ();
 sg13g2_decap_8 FILLER_28_2800 ();
 sg13g2_decap_8 FILLER_28_2807 ();
 sg13g2_decap_8 FILLER_28_2814 ();
 sg13g2_decap_8 FILLER_28_2821 ();
 sg13g2_decap_8 FILLER_28_2828 ();
 sg13g2_decap_8 FILLER_28_2835 ();
 sg13g2_decap_8 FILLER_28_2842 ();
 sg13g2_decap_8 FILLER_28_2849 ();
 sg13g2_decap_8 FILLER_28_2856 ();
 sg13g2_decap_8 FILLER_28_2863 ();
 sg13g2_decap_8 FILLER_28_2870 ();
 sg13g2_decap_8 FILLER_28_2877 ();
 sg13g2_decap_8 FILLER_28_2884 ();
 sg13g2_decap_8 FILLER_28_2891 ();
 sg13g2_decap_8 FILLER_28_2898 ();
 sg13g2_decap_8 FILLER_28_2905 ();
 sg13g2_decap_8 FILLER_28_2912 ();
 sg13g2_decap_8 FILLER_28_2919 ();
 sg13g2_decap_8 FILLER_28_2926 ();
 sg13g2_decap_8 FILLER_28_2933 ();
 sg13g2_decap_8 FILLER_28_2940 ();
 sg13g2_decap_8 FILLER_28_2947 ();
 sg13g2_decap_8 FILLER_28_2954 ();
 sg13g2_decap_8 FILLER_28_2961 ();
 sg13g2_decap_8 FILLER_28_2968 ();
 sg13g2_decap_8 FILLER_28_2975 ();
 sg13g2_decap_8 FILLER_28_2982 ();
 sg13g2_decap_8 FILLER_28_2989 ();
 sg13g2_decap_8 FILLER_28_2996 ();
 sg13g2_decap_8 FILLER_28_3003 ();
 sg13g2_decap_8 FILLER_28_3010 ();
 sg13g2_decap_8 FILLER_28_3017 ();
 sg13g2_decap_8 FILLER_28_3024 ();
 sg13g2_decap_8 FILLER_28_3031 ();
 sg13g2_decap_8 FILLER_28_3038 ();
 sg13g2_decap_8 FILLER_28_3045 ();
 sg13g2_decap_8 FILLER_28_3052 ();
 sg13g2_decap_8 FILLER_28_3059 ();
 sg13g2_decap_8 FILLER_28_3066 ();
 sg13g2_decap_8 FILLER_28_3073 ();
 sg13g2_decap_8 FILLER_28_3080 ();
 sg13g2_decap_8 FILLER_28_3087 ();
 sg13g2_decap_8 FILLER_28_3094 ();
 sg13g2_decap_8 FILLER_28_3101 ();
 sg13g2_decap_8 FILLER_28_3108 ();
 sg13g2_decap_8 FILLER_28_3115 ();
 sg13g2_decap_8 FILLER_28_3122 ();
 sg13g2_decap_8 FILLER_28_3129 ();
 sg13g2_decap_8 FILLER_28_3136 ();
 sg13g2_decap_8 FILLER_28_3143 ();
 sg13g2_decap_8 FILLER_28_3150 ();
 sg13g2_decap_8 FILLER_28_3157 ();
 sg13g2_decap_8 FILLER_28_3164 ();
 sg13g2_decap_8 FILLER_28_3171 ();
 sg13g2_decap_8 FILLER_28_3178 ();
 sg13g2_decap_8 FILLER_28_3185 ();
 sg13g2_decap_8 FILLER_28_3192 ();
 sg13g2_decap_8 FILLER_28_3199 ();
 sg13g2_decap_8 FILLER_28_3206 ();
 sg13g2_decap_8 FILLER_28_3213 ();
 sg13g2_decap_8 FILLER_28_3220 ();
 sg13g2_decap_8 FILLER_28_3227 ();
 sg13g2_decap_8 FILLER_28_3234 ();
 sg13g2_decap_8 FILLER_28_3241 ();
 sg13g2_decap_8 FILLER_28_3248 ();
 sg13g2_decap_8 FILLER_28_3255 ();
 sg13g2_decap_8 FILLER_28_3262 ();
 sg13g2_decap_8 FILLER_28_3269 ();
 sg13g2_decap_8 FILLER_28_3276 ();
 sg13g2_decap_8 FILLER_28_3283 ();
 sg13g2_decap_8 FILLER_28_3290 ();
 sg13g2_decap_8 FILLER_28_3297 ();
 sg13g2_decap_8 FILLER_28_3304 ();
 sg13g2_decap_8 FILLER_28_3311 ();
 sg13g2_decap_8 FILLER_28_3318 ();
 sg13g2_decap_8 FILLER_28_3325 ();
 sg13g2_decap_8 FILLER_28_3332 ();
 sg13g2_decap_8 FILLER_28_3339 ();
 sg13g2_decap_8 FILLER_28_3346 ();
 sg13g2_decap_8 FILLER_28_3353 ();
 sg13g2_decap_8 FILLER_28_3360 ();
 sg13g2_decap_8 FILLER_28_3367 ();
 sg13g2_decap_8 FILLER_28_3374 ();
 sg13g2_decap_8 FILLER_28_3381 ();
 sg13g2_decap_8 FILLER_28_3388 ();
 sg13g2_decap_8 FILLER_28_3395 ();
 sg13g2_decap_8 FILLER_28_3402 ();
 sg13g2_decap_8 FILLER_28_3409 ();
 sg13g2_decap_8 FILLER_28_3416 ();
 sg13g2_decap_8 FILLER_28_3423 ();
 sg13g2_decap_8 FILLER_28_3430 ();
 sg13g2_decap_8 FILLER_28_3437 ();
 sg13g2_decap_8 FILLER_28_3444 ();
 sg13g2_decap_8 FILLER_28_3451 ();
 sg13g2_decap_8 FILLER_28_3458 ();
 sg13g2_decap_8 FILLER_28_3465 ();
 sg13g2_decap_8 FILLER_28_3472 ();
 sg13g2_decap_8 FILLER_28_3479 ();
 sg13g2_decap_8 FILLER_28_3486 ();
 sg13g2_decap_8 FILLER_28_3493 ();
 sg13g2_decap_8 FILLER_28_3500 ();
 sg13g2_decap_8 FILLER_28_3507 ();
 sg13g2_decap_8 FILLER_28_3514 ();
 sg13g2_decap_8 FILLER_28_3521 ();
 sg13g2_decap_8 FILLER_28_3528 ();
 sg13g2_decap_8 FILLER_28_3535 ();
 sg13g2_decap_8 FILLER_28_3542 ();
 sg13g2_decap_8 FILLER_28_3549 ();
 sg13g2_decap_8 FILLER_28_3556 ();
 sg13g2_decap_8 FILLER_28_3563 ();
 sg13g2_decap_8 FILLER_28_3570 ();
 sg13g2_fill_2 FILLER_28_3577 ();
 sg13g2_fill_1 FILLER_28_3579 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_decap_8 FILLER_29_224 ();
 sg13g2_decap_8 FILLER_29_231 ();
 sg13g2_decap_8 FILLER_29_238 ();
 sg13g2_decap_8 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_252 ();
 sg13g2_decap_8 FILLER_29_259 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_decap_8 FILLER_29_273 ();
 sg13g2_decap_8 FILLER_29_280 ();
 sg13g2_decap_8 FILLER_29_287 ();
 sg13g2_decap_8 FILLER_29_294 ();
 sg13g2_decap_8 FILLER_29_301 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_decap_8 FILLER_29_315 ();
 sg13g2_decap_8 FILLER_29_322 ();
 sg13g2_decap_8 FILLER_29_329 ();
 sg13g2_decap_8 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_343 ();
 sg13g2_decap_8 FILLER_29_350 ();
 sg13g2_decap_8 FILLER_29_357 ();
 sg13g2_decap_8 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_29_371 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_decap_8 FILLER_29_406 ();
 sg13g2_decap_8 FILLER_29_413 ();
 sg13g2_decap_8 FILLER_29_420 ();
 sg13g2_decap_8 FILLER_29_427 ();
 sg13g2_decap_8 FILLER_29_434 ();
 sg13g2_decap_8 FILLER_29_441 ();
 sg13g2_decap_8 FILLER_29_448 ();
 sg13g2_decap_8 FILLER_29_455 ();
 sg13g2_decap_8 FILLER_29_462 ();
 sg13g2_decap_8 FILLER_29_469 ();
 sg13g2_decap_8 FILLER_29_476 ();
 sg13g2_decap_8 FILLER_29_483 ();
 sg13g2_decap_8 FILLER_29_490 ();
 sg13g2_decap_8 FILLER_29_497 ();
 sg13g2_decap_8 FILLER_29_504 ();
 sg13g2_decap_8 FILLER_29_511 ();
 sg13g2_decap_8 FILLER_29_518 ();
 sg13g2_decap_8 FILLER_29_525 ();
 sg13g2_decap_8 FILLER_29_532 ();
 sg13g2_decap_8 FILLER_29_539 ();
 sg13g2_decap_8 FILLER_29_546 ();
 sg13g2_decap_8 FILLER_29_553 ();
 sg13g2_decap_8 FILLER_29_560 ();
 sg13g2_decap_8 FILLER_29_567 ();
 sg13g2_decap_8 FILLER_29_574 ();
 sg13g2_decap_8 FILLER_29_581 ();
 sg13g2_decap_8 FILLER_29_588 ();
 sg13g2_decap_8 FILLER_29_595 ();
 sg13g2_decap_8 FILLER_29_602 ();
 sg13g2_decap_8 FILLER_29_609 ();
 sg13g2_decap_8 FILLER_29_616 ();
 sg13g2_decap_8 FILLER_29_623 ();
 sg13g2_decap_8 FILLER_29_630 ();
 sg13g2_decap_8 FILLER_29_637 ();
 sg13g2_decap_8 FILLER_29_644 ();
 sg13g2_decap_8 FILLER_29_651 ();
 sg13g2_decap_8 FILLER_29_658 ();
 sg13g2_decap_8 FILLER_29_665 ();
 sg13g2_decap_8 FILLER_29_672 ();
 sg13g2_decap_8 FILLER_29_679 ();
 sg13g2_decap_8 FILLER_29_686 ();
 sg13g2_decap_8 FILLER_29_693 ();
 sg13g2_decap_8 FILLER_29_700 ();
 sg13g2_decap_8 FILLER_29_707 ();
 sg13g2_decap_8 FILLER_29_714 ();
 sg13g2_decap_8 FILLER_29_721 ();
 sg13g2_decap_8 FILLER_29_728 ();
 sg13g2_decap_8 FILLER_29_735 ();
 sg13g2_decap_8 FILLER_29_742 ();
 sg13g2_decap_8 FILLER_29_749 ();
 sg13g2_decap_8 FILLER_29_756 ();
 sg13g2_decap_8 FILLER_29_763 ();
 sg13g2_decap_8 FILLER_29_770 ();
 sg13g2_decap_8 FILLER_29_777 ();
 sg13g2_decap_8 FILLER_29_784 ();
 sg13g2_decap_8 FILLER_29_791 ();
 sg13g2_decap_8 FILLER_29_798 ();
 sg13g2_decap_8 FILLER_29_805 ();
 sg13g2_decap_8 FILLER_29_812 ();
 sg13g2_decap_8 FILLER_29_819 ();
 sg13g2_decap_8 FILLER_29_826 ();
 sg13g2_decap_8 FILLER_29_833 ();
 sg13g2_decap_8 FILLER_29_840 ();
 sg13g2_decap_8 FILLER_29_847 ();
 sg13g2_decap_8 FILLER_29_854 ();
 sg13g2_decap_8 FILLER_29_861 ();
 sg13g2_decap_8 FILLER_29_868 ();
 sg13g2_decap_8 FILLER_29_875 ();
 sg13g2_decap_8 FILLER_29_882 ();
 sg13g2_decap_8 FILLER_29_889 ();
 sg13g2_decap_8 FILLER_29_896 ();
 sg13g2_decap_8 FILLER_29_903 ();
 sg13g2_decap_8 FILLER_29_910 ();
 sg13g2_decap_8 FILLER_29_917 ();
 sg13g2_decap_8 FILLER_29_924 ();
 sg13g2_decap_8 FILLER_29_931 ();
 sg13g2_decap_8 FILLER_29_938 ();
 sg13g2_decap_8 FILLER_29_945 ();
 sg13g2_decap_8 FILLER_29_952 ();
 sg13g2_decap_8 FILLER_29_959 ();
 sg13g2_decap_8 FILLER_29_966 ();
 sg13g2_decap_8 FILLER_29_973 ();
 sg13g2_decap_8 FILLER_29_980 ();
 sg13g2_decap_8 FILLER_29_987 ();
 sg13g2_decap_8 FILLER_29_994 ();
 sg13g2_decap_8 FILLER_29_1001 ();
 sg13g2_decap_8 FILLER_29_1008 ();
 sg13g2_decap_8 FILLER_29_1015 ();
 sg13g2_decap_8 FILLER_29_1022 ();
 sg13g2_decap_8 FILLER_29_1029 ();
 sg13g2_decap_8 FILLER_29_1036 ();
 sg13g2_decap_8 FILLER_29_1043 ();
 sg13g2_decap_8 FILLER_29_1050 ();
 sg13g2_decap_8 FILLER_29_1057 ();
 sg13g2_decap_8 FILLER_29_1064 ();
 sg13g2_decap_8 FILLER_29_1071 ();
 sg13g2_decap_8 FILLER_29_1078 ();
 sg13g2_decap_8 FILLER_29_1085 ();
 sg13g2_decap_8 FILLER_29_1092 ();
 sg13g2_decap_8 FILLER_29_1099 ();
 sg13g2_decap_8 FILLER_29_1106 ();
 sg13g2_decap_8 FILLER_29_1113 ();
 sg13g2_decap_8 FILLER_29_1120 ();
 sg13g2_decap_8 FILLER_29_1127 ();
 sg13g2_decap_8 FILLER_29_1134 ();
 sg13g2_decap_8 FILLER_29_1141 ();
 sg13g2_decap_8 FILLER_29_1148 ();
 sg13g2_decap_8 FILLER_29_1155 ();
 sg13g2_decap_8 FILLER_29_1162 ();
 sg13g2_decap_8 FILLER_29_1169 ();
 sg13g2_decap_8 FILLER_29_1176 ();
 sg13g2_decap_8 FILLER_29_1183 ();
 sg13g2_decap_8 FILLER_29_1190 ();
 sg13g2_decap_8 FILLER_29_1197 ();
 sg13g2_decap_8 FILLER_29_1204 ();
 sg13g2_decap_8 FILLER_29_1211 ();
 sg13g2_decap_8 FILLER_29_1218 ();
 sg13g2_decap_8 FILLER_29_1225 ();
 sg13g2_decap_8 FILLER_29_1232 ();
 sg13g2_decap_8 FILLER_29_1239 ();
 sg13g2_decap_8 FILLER_29_1246 ();
 sg13g2_decap_8 FILLER_29_1253 ();
 sg13g2_decap_8 FILLER_29_1260 ();
 sg13g2_decap_8 FILLER_29_1267 ();
 sg13g2_decap_8 FILLER_29_1274 ();
 sg13g2_decap_8 FILLER_29_1281 ();
 sg13g2_decap_8 FILLER_29_1288 ();
 sg13g2_decap_8 FILLER_29_1295 ();
 sg13g2_decap_8 FILLER_29_1302 ();
 sg13g2_decap_8 FILLER_29_1309 ();
 sg13g2_decap_8 FILLER_29_1316 ();
 sg13g2_decap_8 FILLER_29_1323 ();
 sg13g2_decap_8 FILLER_29_1330 ();
 sg13g2_decap_8 FILLER_29_1337 ();
 sg13g2_decap_8 FILLER_29_1344 ();
 sg13g2_decap_8 FILLER_29_1351 ();
 sg13g2_decap_8 FILLER_29_1358 ();
 sg13g2_decap_8 FILLER_29_1365 ();
 sg13g2_decap_8 FILLER_29_1372 ();
 sg13g2_decap_8 FILLER_29_1379 ();
 sg13g2_decap_8 FILLER_29_1386 ();
 sg13g2_decap_8 FILLER_29_1393 ();
 sg13g2_decap_8 FILLER_29_1400 ();
 sg13g2_decap_8 FILLER_29_1407 ();
 sg13g2_decap_8 FILLER_29_1414 ();
 sg13g2_decap_8 FILLER_29_1421 ();
 sg13g2_decap_8 FILLER_29_1428 ();
 sg13g2_decap_8 FILLER_29_1435 ();
 sg13g2_decap_8 FILLER_29_1442 ();
 sg13g2_decap_8 FILLER_29_1449 ();
 sg13g2_decap_8 FILLER_29_1456 ();
 sg13g2_decap_8 FILLER_29_1463 ();
 sg13g2_decap_8 FILLER_29_1470 ();
 sg13g2_decap_8 FILLER_29_1477 ();
 sg13g2_decap_8 FILLER_29_1484 ();
 sg13g2_decap_8 FILLER_29_1491 ();
 sg13g2_decap_8 FILLER_29_1498 ();
 sg13g2_decap_8 FILLER_29_1505 ();
 sg13g2_decap_8 FILLER_29_1512 ();
 sg13g2_decap_8 FILLER_29_1519 ();
 sg13g2_decap_8 FILLER_29_1526 ();
 sg13g2_decap_8 FILLER_29_1533 ();
 sg13g2_decap_8 FILLER_29_1540 ();
 sg13g2_decap_8 FILLER_29_1547 ();
 sg13g2_decap_8 FILLER_29_1554 ();
 sg13g2_decap_8 FILLER_29_1561 ();
 sg13g2_decap_8 FILLER_29_1568 ();
 sg13g2_decap_8 FILLER_29_1575 ();
 sg13g2_decap_8 FILLER_29_1582 ();
 sg13g2_decap_8 FILLER_29_1589 ();
 sg13g2_decap_8 FILLER_29_1596 ();
 sg13g2_decap_8 FILLER_29_1603 ();
 sg13g2_decap_8 FILLER_29_1610 ();
 sg13g2_decap_8 FILLER_29_1617 ();
 sg13g2_decap_8 FILLER_29_1624 ();
 sg13g2_decap_8 FILLER_29_1631 ();
 sg13g2_decap_8 FILLER_29_1638 ();
 sg13g2_decap_8 FILLER_29_1645 ();
 sg13g2_decap_8 FILLER_29_1652 ();
 sg13g2_decap_8 FILLER_29_1659 ();
 sg13g2_decap_8 FILLER_29_1666 ();
 sg13g2_decap_8 FILLER_29_1673 ();
 sg13g2_decap_8 FILLER_29_1680 ();
 sg13g2_decap_8 FILLER_29_1687 ();
 sg13g2_decap_8 FILLER_29_1694 ();
 sg13g2_decap_8 FILLER_29_1701 ();
 sg13g2_decap_8 FILLER_29_1708 ();
 sg13g2_decap_8 FILLER_29_1715 ();
 sg13g2_decap_8 FILLER_29_1722 ();
 sg13g2_decap_8 FILLER_29_1729 ();
 sg13g2_decap_8 FILLER_29_1736 ();
 sg13g2_decap_8 FILLER_29_1743 ();
 sg13g2_decap_8 FILLER_29_1750 ();
 sg13g2_decap_8 FILLER_29_1757 ();
 sg13g2_decap_8 FILLER_29_1764 ();
 sg13g2_decap_8 FILLER_29_1771 ();
 sg13g2_decap_8 FILLER_29_1778 ();
 sg13g2_decap_8 FILLER_29_1785 ();
 sg13g2_decap_8 FILLER_29_1792 ();
 sg13g2_decap_8 FILLER_29_1799 ();
 sg13g2_decap_8 FILLER_29_1806 ();
 sg13g2_decap_8 FILLER_29_1813 ();
 sg13g2_decap_8 FILLER_29_1820 ();
 sg13g2_decap_8 FILLER_29_1827 ();
 sg13g2_decap_8 FILLER_29_1834 ();
 sg13g2_decap_8 FILLER_29_1841 ();
 sg13g2_decap_8 FILLER_29_1848 ();
 sg13g2_decap_8 FILLER_29_1855 ();
 sg13g2_decap_8 FILLER_29_1862 ();
 sg13g2_decap_8 FILLER_29_1869 ();
 sg13g2_decap_8 FILLER_29_1876 ();
 sg13g2_decap_8 FILLER_29_1883 ();
 sg13g2_decap_8 FILLER_29_1890 ();
 sg13g2_decap_8 FILLER_29_1897 ();
 sg13g2_decap_8 FILLER_29_1904 ();
 sg13g2_decap_8 FILLER_29_1911 ();
 sg13g2_decap_8 FILLER_29_1918 ();
 sg13g2_decap_8 FILLER_29_1925 ();
 sg13g2_decap_8 FILLER_29_1932 ();
 sg13g2_decap_8 FILLER_29_1939 ();
 sg13g2_decap_8 FILLER_29_1946 ();
 sg13g2_decap_8 FILLER_29_1953 ();
 sg13g2_decap_8 FILLER_29_1960 ();
 sg13g2_decap_8 FILLER_29_1967 ();
 sg13g2_decap_8 FILLER_29_1974 ();
 sg13g2_decap_8 FILLER_29_1981 ();
 sg13g2_decap_8 FILLER_29_1988 ();
 sg13g2_decap_8 FILLER_29_1995 ();
 sg13g2_decap_8 FILLER_29_2002 ();
 sg13g2_decap_8 FILLER_29_2009 ();
 sg13g2_decap_8 FILLER_29_2016 ();
 sg13g2_decap_8 FILLER_29_2023 ();
 sg13g2_decap_8 FILLER_29_2030 ();
 sg13g2_decap_8 FILLER_29_2037 ();
 sg13g2_decap_8 FILLER_29_2044 ();
 sg13g2_decap_8 FILLER_29_2051 ();
 sg13g2_decap_8 FILLER_29_2058 ();
 sg13g2_decap_8 FILLER_29_2065 ();
 sg13g2_decap_8 FILLER_29_2072 ();
 sg13g2_decap_8 FILLER_29_2079 ();
 sg13g2_decap_8 FILLER_29_2086 ();
 sg13g2_decap_8 FILLER_29_2093 ();
 sg13g2_decap_8 FILLER_29_2100 ();
 sg13g2_decap_8 FILLER_29_2107 ();
 sg13g2_decap_8 FILLER_29_2114 ();
 sg13g2_decap_8 FILLER_29_2121 ();
 sg13g2_decap_8 FILLER_29_2128 ();
 sg13g2_decap_8 FILLER_29_2135 ();
 sg13g2_decap_8 FILLER_29_2142 ();
 sg13g2_decap_8 FILLER_29_2149 ();
 sg13g2_decap_8 FILLER_29_2156 ();
 sg13g2_decap_8 FILLER_29_2163 ();
 sg13g2_decap_8 FILLER_29_2170 ();
 sg13g2_decap_8 FILLER_29_2177 ();
 sg13g2_decap_8 FILLER_29_2184 ();
 sg13g2_decap_8 FILLER_29_2191 ();
 sg13g2_decap_8 FILLER_29_2198 ();
 sg13g2_decap_8 FILLER_29_2205 ();
 sg13g2_decap_8 FILLER_29_2212 ();
 sg13g2_decap_8 FILLER_29_2219 ();
 sg13g2_decap_8 FILLER_29_2226 ();
 sg13g2_decap_8 FILLER_29_2233 ();
 sg13g2_decap_8 FILLER_29_2240 ();
 sg13g2_decap_8 FILLER_29_2247 ();
 sg13g2_decap_8 FILLER_29_2254 ();
 sg13g2_decap_8 FILLER_29_2261 ();
 sg13g2_decap_8 FILLER_29_2268 ();
 sg13g2_decap_8 FILLER_29_2275 ();
 sg13g2_decap_8 FILLER_29_2282 ();
 sg13g2_decap_8 FILLER_29_2289 ();
 sg13g2_decap_8 FILLER_29_2296 ();
 sg13g2_decap_8 FILLER_29_2303 ();
 sg13g2_decap_8 FILLER_29_2310 ();
 sg13g2_decap_8 FILLER_29_2317 ();
 sg13g2_decap_8 FILLER_29_2324 ();
 sg13g2_decap_8 FILLER_29_2331 ();
 sg13g2_decap_8 FILLER_29_2338 ();
 sg13g2_decap_8 FILLER_29_2345 ();
 sg13g2_decap_8 FILLER_29_2352 ();
 sg13g2_decap_8 FILLER_29_2359 ();
 sg13g2_decap_8 FILLER_29_2366 ();
 sg13g2_decap_8 FILLER_29_2373 ();
 sg13g2_decap_8 FILLER_29_2380 ();
 sg13g2_decap_8 FILLER_29_2387 ();
 sg13g2_decap_8 FILLER_29_2394 ();
 sg13g2_decap_8 FILLER_29_2401 ();
 sg13g2_decap_8 FILLER_29_2408 ();
 sg13g2_decap_8 FILLER_29_2415 ();
 sg13g2_decap_8 FILLER_29_2422 ();
 sg13g2_decap_8 FILLER_29_2429 ();
 sg13g2_decap_8 FILLER_29_2436 ();
 sg13g2_decap_8 FILLER_29_2443 ();
 sg13g2_decap_8 FILLER_29_2450 ();
 sg13g2_decap_8 FILLER_29_2457 ();
 sg13g2_decap_8 FILLER_29_2464 ();
 sg13g2_decap_8 FILLER_29_2471 ();
 sg13g2_decap_8 FILLER_29_2478 ();
 sg13g2_decap_8 FILLER_29_2485 ();
 sg13g2_decap_8 FILLER_29_2492 ();
 sg13g2_decap_8 FILLER_29_2499 ();
 sg13g2_decap_8 FILLER_29_2506 ();
 sg13g2_decap_8 FILLER_29_2513 ();
 sg13g2_decap_8 FILLER_29_2520 ();
 sg13g2_decap_8 FILLER_29_2527 ();
 sg13g2_decap_8 FILLER_29_2534 ();
 sg13g2_decap_8 FILLER_29_2541 ();
 sg13g2_decap_8 FILLER_29_2548 ();
 sg13g2_decap_8 FILLER_29_2555 ();
 sg13g2_decap_8 FILLER_29_2562 ();
 sg13g2_decap_8 FILLER_29_2569 ();
 sg13g2_decap_8 FILLER_29_2576 ();
 sg13g2_decap_8 FILLER_29_2583 ();
 sg13g2_decap_8 FILLER_29_2590 ();
 sg13g2_decap_8 FILLER_29_2597 ();
 sg13g2_decap_8 FILLER_29_2604 ();
 sg13g2_decap_8 FILLER_29_2611 ();
 sg13g2_decap_8 FILLER_29_2618 ();
 sg13g2_decap_8 FILLER_29_2625 ();
 sg13g2_decap_8 FILLER_29_2632 ();
 sg13g2_decap_8 FILLER_29_2639 ();
 sg13g2_decap_8 FILLER_29_2646 ();
 sg13g2_decap_8 FILLER_29_2653 ();
 sg13g2_decap_8 FILLER_29_2660 ();
 sg13g2_decap_8 FILLER_29_2667 ();
 sg13g2_decap_8 FILLER_29_2674 ();
 sg13g2_decap_8 FILLER_29_2681 ();
 sg13g2_decap_8 FILLER_29_2688 ();
 sg13g2_decap_8 FILLER_29_2695 ();
 sg13g2_decap_8 FILLER_29_2702 ();
 sg13g2_decap_8 FILLER_29_2709 ();
 sg13g2_decap_8 FILLER_29_2716 ();
 sg13g2_decap_8 FILLER_29_2723 ();
 sg13g2_decap_8 FILLER_29_2730 ();
 sg13g2_decap_8 FILLER_29_2737 ();
 sg13g2_decap_8 FILLER_29_2744 ();
 sg13g2_decap_8 FILLER_29_2751 ();
 sg13g2_decap_8 FILLER_29_2758 ();
 sg13g2_decap_8 FILLER_29_2765 ();
 sg13g2_decap_8 FILLER_29_2772 ();
 sg13g2_decap_8 FILLER_29_2779 ();
 sg13g2_decap_8 FILLER_29_2786 ();
 sg13g2_decap_8 FILLER_29_2793 ();
 sg13g2_decap_8 FILLER_29_2800 ();
 sg13g2_decap_8 FILLER_29_2807 ();
 sg13g2_decap_8 FILLER_29_2814 ();
 sg13g2_decap_8 FILLER_29_2821 ();
 sg13g2_decap_8 FILLER_29_2828 ();
 sg13g2_decap_8 FILLER_29_2835 ();
 sg13g2_decap_8 FILLER_29_2842 ();
 sg13g2_decap_8 FILLER_29_2849 ();
 sg13g2_decap_8 FILLER_29_2856 ();
 sg13g2_decap_8 FILLER_29_2863 ();
 sg13g2_decap_8 FILLER_29_2870 ();
 sg13g2_decap_8 FILLER_29_2877 ();
 sg13g2_decap_8 FILLER_29_2884 ();
 sg13g2_decap_8 FILLER_29_2891 ();
 sg13g2_decap_8 FILLER_29_2898 ();
 sg13g2_decap_8 FILLER_29_2905 ();
 sg13g2_decap_8 FILLER_29_2912 ();
 sg13g2_decap_8 FILLER_29_2919 ();
 sg13g2_decap_8 FILLER_29_2926 ();
 sg13g2_decap_8 FILLER_29_2933 ();
 sg13g2_decap_8 FILLER_29_2940 ();
 sg13g2_decap_8 FILLER_29_2947 ();
 sg13g2_decap_8 FILLER_29_2954 ();
 sg13g2_decap_8 FILLER_29_2961 ();
 sg13g2_decap_8 FILLER_29_2968 ();
 sg13g2_decap_8 FILLER_29_2975 ();
 sg13g2_decap_8 FILLER_29_2982 ();
 sg13g2_decap_8 FILLER_29_2989 ();
 sg13g2_decap_8 FILLER_29_2996 ();
 sg13g2_decap_8 FILLER_29_3003 ();
 sg13g2_decap_8 FILLER_29_3010 ();
 sg13g2_decap_8 FILLER_29_3017 ();
 sg13g2_decap_8 FILLER_29_3024 ();
 sg13g2_decap_8 FILLER_29_3031 ();
 sg13g2_decap_8 FILLER_29_3038 ();
 sg13g2_decap_8 FILLER_29_3045 ();
 sg13g2_decap_8 FILLER_29_3052 ();
 sg13g2_decap_8 FILLER_29_3059 ();
 sg13g2_decap_8 FILLER_29_3066 ();
 sg13g2_decap_8 FILLER_29_3073 ();
 sg13g2_decap_8 FILLER_29_3080 ();
 sg13g2_decap_8 FILLER_29_3087 ();
 sg13g2_decap_8 FILLER_29_3094 ();
 sg13g2_decap_8 FILLER_29_3101 ();
 sg13g2_decap_8 FILLER_29_3108 ();
 sg13g2_decap_8 FILLER_29_3115 ();
 sg13g2_decap_8 FILLER_29_3122 ();
 sg13g2_decap_8 FILLER_29_3129 ();
 sg13g2_decap_8 FILLER_29_3136 ();
 sg13g2_decap_8 FILLER_29_3143 ();
 sg13g2_decap_8 FILLER_29_3150 ();
 sg13g2_decap_8 FILLER_29_3157 ();
 sg13g2_decap_8 FILLER_29_3164 ();
 sg13g2_decap_8 FILLER_29_3171 ();
 sg13g2_decap_8 FILLER_29_3178 ();
 sg13g2_decap_8 FILLER_29_3185 ();
 sg13g2_decap_8 FILLER_29_3192 ();
 sg13g2_decap_8 FILLER_29_3199 ();
 sg13g2_decap_8 FILLER_29_3206 ();
 sg13g2_decap_8 FILLER_29_3213 ();
 sg13g2_decap_8 FILLER_29_3220 ();
 sg13g2_decap_8 FILLER_29_3227 ();
 sg13g2_decap_8 FILLER_29_3234 ();
 sg13g2_decap_8 FILLER_29_3241 ();
 sg13g2_decap_8 FILLER_29_3248 ();
 sg13g2_decap_8 FILLER_29_3255 ();
 sg13g2_decap_8 FILLER_29_3262 ();
 sg13g2_decap_8 FILLER_29_3269 ();
 sg13g2_decap_8 FILLER_29_3276 ();
 sg13g2_decap_8 FILLER_29_3283 ();
 sg13g2_decap_8 FILLER_29_3290 ();
 sg13g2_decap_8 FILLER_29_3297 ();
 sg13g2_decap_8 FILLER_29_3304 ();
 sg13g2_decap_8 FILLER_29_3311 ();
 sg13g2_decap_8 FILLER_29_3318 ();
 sg13g2_decap_8 FILLER_29_3325 ();
 sg13g2_decap_8 FILLER_29_3332 ();
 sg13g2_decap_8 FILLER_29_3339 ();
 sg13g2_decap_8 FILLER_29_3346 ();
 sg13g2_decap_8 FILLER_29_3353 ();
 sg13g2_decap_8 FILLER_29_3360 ();
 sg13g2_decap_8 FILLER_29_3367 ();
 sg13g2_decap_8 FILLER_29_3374 ();
 sg13g2_decap_8 FILLER_29_3381 ();
 sg13g2_decap_8 FILLER_29_3388 ();
 sg13g2_decap_8 FILLER_29_3395 ();
 sg13g2_decap_8 FILLER_29_3402 ();
 sg13g2_decap_8 FILLER_29_3409 ();
 sg13g2_decap_8 FILLER_29_3416 ();
 sg13g2_decap_8 FILLER_29_3423 ();
 sg13g2_decap_8 FILLER_29_3430 ();
 sg13g2_decap_8 FILLER_29_3437 ();
 sg13g2_decap_8 FILLER_29_3444 ();
 sg13g2_decap_8 FILLER_29_3451 ();
 sg13g2_decap_8 FILLER_29_3458 ();
 sg13g2_decap_8 FILLER_29_3465 ();
 sg13g2_decap_8 FILLER_29_3472 ();
 sg13g2_decap_8 FILLER_29_3479 ();
 sg13g2_decap_8 FILLER_29_3486 ();
 sg13g2_decap_8 FILLER_29_3493 ();
 sg13g2_decap_8 FILLER_29_3500 ();
 sg13g2_decap_8 FILLER_29_3507 ();
 sg13g2_decap_8 FILLER_29_3514 ();
 sg13g2_decap_8 FILLER_29_3521 ();
 sg13g2_decap_8 FILLER_29_3528 ();
 sg13g2_decap_8 FILLER_29_3535 ();
 sg13g2_decap_8 FILLER_29_3542 ();
 sg13g2_decap_8 FILLER_29_3549 ();
 sg13g2_decap_8 FILLER_29_3556 ();
 sg13g2_decap_8 FILLER_29_3563 ();
 sg13g2_decap_8 FILLER_29_3570 ();
 sg13g2_fill_2 FILLER_29_3577 ();
 sg13g2_fill_1 FILLER_29_3579 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_decap_8 FILLER_30_266 ();
 sg13g2_decap_8 FILLER_30_273 ();
 sg13g2_decap_8 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_decap_8 FILLER_30_294 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_decap_8 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_decap_8 FILLER_30_343 ();
 sg13g2_decap_8 FILLER_30_350 ();
 sg13g2_decap_8 FILLER_30_357 ();
 sg13g2_decap_8 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_30_371 ();
 sg13g2_decap_8 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_decap_8 FILLER_30_406 ();
 sg13g2_decap_8 FILLER_30_413 ();
 sg13g2_decap_8 FILLER_30_420 ();
 sg13g2_decap_8 FILLER_30_427 ();
 sg13g2_decap_8 FILLER_30_434 ();
 sg13g2_decap_8 FILLER_30_441 ();
 sg13g2_decap_8 FILLER_30_448 ();
 sg13g2_decap_8 FILLER_30_455 ();
 sg13g2_decap_8 FILLER_30_462 ();
 sg13g2_decap_8 FILLER_30_469 ();
 sg13g2_decap_8 FILLER_30_476 ();
 sg13g2_decap_8 FILLER_30_483 ();
 sg13g2_decap_8 FILLER_30_490 ();
 sg13g2_decap_8 FILLER_30_497 ();
 sg13g2_decap_8 FILLER_30_504 ();
 sg13g2_decap_8 FILLER_30_511 ();
 sg13g2_decap_8 FILLER_30_518 ();
 sg13g2_decap_8 FILLER_30_525 ();
 sg13g2_decap_8 FILLER_30_532 ();
 sg13g2_decap_8 FILLER_30_539 ();
 sg13g2_decap_8 FILLER_30_546 ();
 sg13g2_decap_8 FILLER_30_553 ();
 sg13g2_decap_8 FILLER_30_560 ();
 sg13g2_decap_8 FILLER_30_567 ();
 sg13g2_decap_8 FILLER_30_574 ();
 sg13g2_decap_8 FILLER_30_581 ();
 sg13g2_decap_8 FILLER_30_588 ();
 sg13g2_decap_8 FILLER_30_595 ();
 sg13g2_decap_8 FILLER_30_602 ();
 sg13g2_decap_8 FILLER_30_609 ();
 sg13g2_decap_8 FILLER_30_616 ();
 sg13g2_decap_8 FILLER_30_623 ();
 sg13g2_decap_8 FILLER_30_630 ();
 sg13g2_decap_8 FILLER_30_637 ();
 sg13g2_decap_8 FILLER_30_644 ();
 sg13g2_decap_8 FILLER_30_651 ();
 sg13g2_decap_8 FILLER_30_658 ();
 sg13g2_decap_8 FILLER_30_665 ();
 sg13g2_decap_8 FILLER_30_672 ();
 sg13g2_decap_8 FILLER_30_679 ();
 sg13g2_decap_8 FILLER_30_686 ();
 sg13g2_decap_8 FILLER_30_693 ();
 sg13g2_decap_8 FILLER_30_700 ();
 sg13g2_decap_8 FILLER_30_707 ();
 sg13g2_decap_8 FILLER_30_714 ();
 sg13g2_decap_8 FILLER_30_721 ();
 sg13g2_decap_8 FILLER_30_728 ();
 sg13g2_decap_8 FILLER_30_735 ();
 sg13g2_decap_8 FILLER_30_742 ();
 sg13g2_decap_8 FILLER_30_749 ();
 sg13g2_decap_8 FILLER_30_756 ();
 sg13g2_decap_8 FILLER_30_763 ();
 sg13g2_decap_8 FILLER_30_770 ();
 sg13g2_decap_8 FILLER_30_777 ();
 sg13g2_decap_8 FILLER_30_784 ();
 sg13g2_decap_8 FILLER_30_791 ();
 sg13g2_decap_8 FILLER_30_798 ();
 sg13g2_decap_8 FILLER_30_805 ();
 sg13g2_decap_8 FILLER_30_812 ();
 sg13g2_decap_8 FILLER_30_819 ();
 sg13g2_decap_8 FILLER_30_826 ();
 sg13g2_decap_8 FILLER_30_833 ();
 sg13g2_decap_8 FILLER_30_840 ();
 sg13g2_decap_8 FILLER_30_847 ();
 sg13g2_decap_8 FILLER_30_854 ();
 sg13g2_decap_8 FILLER_30_861 ();
 sg13g2_decap_8 FILLER_30_868 ();
 sg13g2_decap_8 FILLER_30_875 ();
 sg13g2_decap_8 FILLER_30_882 ();
 sg13g2_decap_8 FILLER_30_889 ();
 sg13g2_decap_8 FILLER_30_896 ();
 sg13g2_decap_8 FILLER_30_903 ();
 sg13g2_decap_8 FILLER_30_910 ();
 sg13g2_decap_8 FILLER_30_917 ();
 sg13g2_decap_8 FILLER_30_924 ();
 sg13g2_decap_8 FILLER_30_931 ();
 sg13g2_decap_8 FILLER_30_938 ();
 sg13g2_decap_8 FILLER_30_945 ();
 sg13g2_decap_8 FILLER_30_952 ();
 sg13g2_decap_8 FILLER_30_959 ();
 sg13g2_decap_8 FILLER_30_966 ();
 sg13g2_decap_8 FILLER_30_973 ();
 sg13g2_decap_8 FILLER_30_980 ();
 sg13g2_decap_8 FILLER_30_987 ();
 sg13g2_decap_8 FILLER_30_994 ();
 sg13g2_decap_8 FILLER_30_1001 ();
 sg13g2_decap_8 FILLER_30_1008 ();
 sg13g2_decap_8 FILLER_30_1015 ();
 sg13g2_decap_8 FILLER_30_1022 ();
 sg13g2_decap_8 FILLER_30_1029 ();
 sg13g2_decap_8 FILLER_30_1036 ();
 sg13g2_decap_8 FILLER_30_1043 ();
 sg13g2_decap_8 FILLER_30_1050 ();
 sg13g2_decap_8 FILLER_30_1057 ();
 sg13g2_decap_8 FILLER_30_1064 ();
 sg13g2_decap_8 FILLER_30_1071 ();
 sg13g2_decap_8 FILLER_30_1078 ();
 sg13g2_decap_8 FILLER_30_1085 ();
 sg13g2_decap_8 FILLER_30_1092 ();
 sg13g2_decap_8 FILLER_30_1099 ();
 sg13g2_decap_8 FILLER_30_1106 ();
 sg13g2_decap_8 FILLER_30_1113 ();
 sg13g2_decap_8 FILLER_30_1120 ();
 sg13g2_decap_8 FILLER_30_1127 ();
 sg13g2_decap_8 FILLER_30_1134 ();
 sg13g2_decap_8 FILLER_30_1141 ();
 sg13g2_decap_8 FILLER_30_1148 ();
 sg13g2_decap_8 FILLER_30_1155 ();
 sg13g2_decap_8 FILLER_30_1162 ();
 sg13g2_decap_8 FILLER_30_1169 ();
 sg13g2_decap_8 FILLER_30_1176 ();
 sg13g2_decap_8 FILLER_30_1183 ();
 sg13g2_decap_8 FILLER_30_1190 ();
 sg13g2_decap_8 FILLER_30_1197 ();
 sg13g2_decap_8 FILLER_30_1204 ();
 sg13g2_decap_8 FILLER_30_1211 ();
 sg13g2_decap_8 FILLER_30_1218 ();
 sg13g2_decap_8 FILLER_30_1225 ();
 sg13g2_decap_8 FILLER_30_1232 ();
 sg13g2_decap_8 FILLER_30_1239 ();
 sg13g2_decap_8 FILLER_30_1246 ();
 sg13g2_decap_8 FILLER_30_1253 ();
 sg13g2_decap_8 FILLER_30_1260 ();
 sg13g2_decap_8 FILLER_30_1267 ();
 sg13g2_decap_8 FILLER_30_1274 ();
 sg13g2_decap_8 FILLER_30_1281 ();
 sg13g2_decap_8 FILLER_30_1288 ();
 sg13g2_decap_8 FILLER_30_1295 ();
 sg13g2_decap_8 FILLER_30_1302 ();
 sg13g2_decap_8 FILLER_30_1309 ();
 sg13g2_decap_8 FILLER_30_1316 ();
 sg13g2_decap_8 FILLER_30_1323 ();
 sg13g2_decap_8 FILLER_30_1330 ();
 sg13g2_decap_8 FILLER_30_1337 ();
 sg13g2_decap_8 FILLER_30_1344 ();
 sg13g2_decap_8 FILLER_30_1351 ();
 sg13g2_decap_8 FILLER_30_1358 ();
 sg13g2_decap_8 FILLER_30_1365 ();
 sg13g2_decap_8 FILLER_30_1372 ();
 sg13g2_decap_8 FILLER_30_1379 ();
 sg13g2_decap_8 FILLER_30_1386 ();
 sg13g2_decap_8 FILLER_30_1393 ();
 sg13g2_decap_8 FILLER_30_1400 ();
 sg13g2_decap_8 FILLER_30_1407 ();
 sg13g2_decap_8 FILLER_30_1414 ();
 sg13g2_decap_8 FILLER_30_1421 ();
 sg13g2_decap_8 FILLER_30_1428 ();
 sg13g2_decap_8 FILLER_30_1435 ();
 sg13g2_decap_8 FILLER_30_1442 ();
 sg13g2_decap_8 FILLER_30_1449 ();
 sg13g2_decap_8 FILLER_30_1456 ();
 sg13g2_decap_8 FILLER_30_1463 ();
 sg13g2_decap_8 FILLER_30_1470 ();
 sg13g2_decap_8 FILLER_30_1477 ();
 sg13g2_decap_8 FILLER_30_1484 ();
 sg13g2_decap_8 FILLER_30_1491 ();
 sg13g2_decap_8 FILLER_30_1498 ();
 sg13g2_decap_8 FILLER_30_1505 ();
 sg13g2_decap_8 FILLER_30_1512 ();
 sg13g2_decap_8 FILLER_30_1519 ();
 sg13g2_decap_8 FILLER_30_1526 ();
 sg13g2_decap_8 FILLER_30_1533 ();
 sg13g2_decap_8 FILLER_30_1540 ();
 sg13g2_decap_8 FILLER_30_1547 ();
 sg13g2_decap_8 FILLER_30_1554 ();
 sg13g2_decap_8 FILLER_30_1561 ();
 sg13g2_decap_8 FILLER_30_1568 ();
 sg13g2_decap_8 FILLER_30_1575 ();
 sg13g2_decap_8 FILLER_30_1582 ();
 sg13g2_decap_8 FILLER_30_1589 ();
 sg13g2_decap_8 FILLER_30_1596 ();
 sg13g2_decap_8 FILLER_30_1603 ();
 sg13g2_decap_8 FILLER_30_1610 ();
 sg13g2_decap_8 FILLER_30_1617 ();
 sg13g2_decap_8 FILLER_30_1624 ();
 sg13g2_decap_8 FILLER_30_1631 ();
 sg13g2_decap_8 FILLER_30_1638 ();
 sg13g2_decap_8 FILLER_30_1645 ();
 sg13g2_decap_8 FILLER_30_1652 ();
 sg13g2_decap_8 FILLER_30_1659 ();
 sg13g2_decap_8 FILLER_30_1666 ();
 sg13g2_decap_8 FILLER_30_1673 ();
 sg13g2_decap_8 FILLER_30_1680 ();
 sg13g2_decap_8 FILLER_30_1687 ();
 sg13g2_decap_8 FILLER_30_1694 ();
 sg13g2_decap_8 FILLER_30_1701 ();
 sg13g2_decap_8 FILLER_30_1708 ();
 sg13g2_decap_8 FILLER_30_1715 ();
 sg13g2_decap_8 FILLER_30_1722 ();
 sg13g2_decap_8 FILLER_30_1729 ();
 sg13g2_decap_8 FILLER_30_1736 ();
 sg13g2_decap_8 FILLER_30_1743 ();
 sg13g2_decap_8 FILLER_30_1750 ();
 sg13g2_decap_8 FILLER_30_1757 ();
 sg13g2_decap_8 FILLER_30_1764 ();
 sg13g2_decap_8 FILLER_30_1771 ();
 sg13g2_decap_8 FILLER_30_1778 ();
 sg13g2_decap_8 FILLER_30_1785 ();
 sg13g2_decap_8 FILLER_30_1792 ();
 sg13g2_decap_8 FILLER_30_1799 ();
 sg13g2_decap_8 FILLER_30_1806 ();
 sg13g2_decap_8 FILLER_30_1813 ();
 sg13g2_decap_8 FILLER_30_1820 ();
 sg13g2_decap_8 FILLER_30_1827 ();
 sg13g2_decap_8 FILLER_30_1834 ();
 sg13g2_decap_8 FILLER_30_1841 ();
 sg13g2_decap_8 FILLER_30_1848 ();
 sg13g2_decap_8 FILLER_30_1855 ();
 sg13g2_decap_8 FILLER_30_1862 ();
 sg13g2_decap_8 FILLER_30_1869 ();
 sg13g2_decap_8 FILLER_30_1876 ();
 sg13g2_decap_8 FILLER_30_1883 ();
 sg13g2_decap_8 FILLER_30_1890 ();
 sg13g2_decap_8 FILLER_30_1897 ();
 sg13g2_decap_8 FILLER_30_1904 ();
 sg13g2_decap_8 FILLER_30_1911 ();
 sg13g2_decap_8 FILLER_30_1918 ();
 sg13g2_decap_8 FILLER_30_1925 ();
 sg13g2_decap_8 FILLER_30_1932 ();
 sg13g2_decap_8 FILLER_30_1939 ();
 sg13g2_decap_8 FILLER_30_1946 ();
 sg13g2_decap_8 FILLER_30_1953 ();
 sg13g2_decap_8 FILLER_30_1960 ();
 sg13g2_decap_8 FILLER_30_1967 ();
 sg13g2_decap_8 FILLER_30_1974 ();
 sg13g2_decap_8 FILLER_30_1981 ();
 sg13g2_decap_8 FILLER_30_1988 ();
 sg13g2_decap_8 FILLER_30_1995 ();
 sg13g2_decap_8 FILLER_30_2002 ();
 sg13g2_decap_8 FILLER_30_2009 ();
 sg13g2_decap_8 FILLER_30_2016 ();
 sg13g2_decap_8 FILLER_30_2023 ();
 sg13g2_decap_8 FILLER_30_2030 ();
 sg13g2_decap_8 FILLER_30_2037 ();
 sg13g2_decap_8 FILLER_30_2044 ();
 sg13g2_decap_8 FILLER_30_2051 ();
 sg13g2_decap_8 FILLER_30_2058 ();
 sg13g2_decap_8 FILLER_30_2065 ();
 sg13g2_decap_8 FILLER_30_2072 ();
 sg13g2_decap_8 FILLER_30_2079 ();
 sg13g2_decap_8 FILLER_30_2086 ();
 sg13g2_decap_8 FILLER_30_2093 ();
 sg13g2_decap_8 FILLER_30_2100 ();
 sg13g2_decap_8 FILLER_30_2107 ();
 sg13g2_decap_8 FILLER_30_2114 ();
 sg13g2_decap_8 FILLER_30_2121 ();
 sg13g2_decap_8 FILLER_30_2128 ();
 sg13g2_decap_8 FILLER_30_2135 ();
 sg13g2_decap_8 FILLER_30_2142 ();
 sg13g2_decap_8 FILLER_30_2149 ();
 sg13g2_decap_8 FILLER_30_2156 ();
 sg13g2_decap_8 FILLER_30_2163 ();
 sg13g2_decap_8 FILLER_30_2170 ();
 sg13g2_decap_8 FILLER_30_2177 ();
 sg13g2_decap_8 FILLER_30_2184 ();
 sg13g2_decap_8 FILLER_30_2191 ();
 sg13g2_decap_8 FILLER_30_2198 ();
 sg13g2_decap_8 FILLER_30_2205 ();
 sg13g2_decap_8 FILLER_30_2212 ();
 sg13g2_decap_8 FILLER_30_2219 ();
 sg13g2_decap_8 FILLER_30_2226 ();
 sg13g2_decap_8 FILLER_30_2233 ();
 sg13g2_decap_8 FILLER_30_2240 ();
 sg13g2_decap_8 FILLER_30_2247 ();
 sg13g2_decap_8 FILLER_30_2254 ();
 sg13g2_decap_8 FILLER_30_2261 ();
 sg13g2_decap_8 FILLER_30_2268 ();
 sg13g2_decap_8 FILLER_30_2275 ();
 sg13g2_decap_8 FILLER_30_2282 ();
 sg13g2_decap_8 FILLER_30_2289 ();
 sg13g2_decap_8 FILLER_30_2296 ();
 sg13g2_decap_8 FILLER_30_2303 ();
 sg13g2_decap_8 FILLER_30_2310 ();
 sg13g2_decap_8 FILLER_30_2317 ();
 sg13g2_decap_8 FILLER_30_2324 ();
 sg13g2_decap_8 FILLER_30_2331 ();
 sg13g2_decap_8 FILLER_30_2338 ();
 sg13g2_decap_8 FILLER_30_2345 ();
 sg13g2_decap_8 FILLER_30_2352 ();
 sg13g2_decap_8 FILLER_30_2359 ();
 sg13g2_decap_8 FILLER_30_2366 ();
 sg13g2_decap_8 FILLER_30_2373 ();
 sg13g2_decap_8 FILLER_30_2380 ();
 sg13g2_decap_8 FILLER_30_2387 ();
 sg13g2_decap_8 FILLER_30_2394 ();
 sg13g2_decap_8 FILLER_30_2401 ();
 sg13g2_decap_8 FILLER_30_2408 ();
 sg13g2_decap_8 FILLER_30_2415 ();
 sg13g2_decap_8 FILLER_30_2422 ();
 sg13g2_decap_8 FILLER_30_2429 ();
 sg13g2_decap_8 FILLER_30_2436 ();
 sg13g2_decap_8 FILLER_30_2443 ();
 sg13g2_decap_8 FILLER_30_2450 ();
 sg13g2_decap_8 FILLER_30_2457 ();
 sg13g2_decap_8 FILLER_30_2464 ();
 sg13g2_decap_8 FILLER_30_2471 ();
 sg13g2_decap_8 FILLER_30_2478 ();
 sg13g2_decap_8 FILLER_30_2485 ();
 sg13g2_decap_8 FILLER_30_2492 ();
 sg13g2_decap_8 FILLER_30_2499 ();
 sg13g2_decap_8 FILLER_30_2506 ();
 sg13g2_decap_8 FILLER_30_2513 ();
 sg13g2_decap_8 FILLER_30_2520 ();
 sg13g2_decap_8 FILLER_30_2527 ();
 sg13g2_decap_8 FILLER_30_2534 ();
 sg13g2_decap_8 FILLER_30_2541 ();
 sg13g2_decap_8 FILLER_30_2548 ();
 sg13g2_decap_8 FILLER_30_2555 ();
 sg13g2_decap_8 FILLER_30_2562 ();
 sg13g2_decap_8 FILLER_30_2569 ();
 sg13g2_decap_8 FILLER_30_2576 ();
 sg13g2_decap_8 FILLER_30_2583 ();
 sg13g2_decap_8 FILLER_30_2590 ();
 sg13g2_decap_8 FILLER_30_2597 ();
 sg13g2_decap_8 FILLER_30_2604 ();
 sg13g2_decap_8 FILLER_30_2611 ();
 sg13g2_decap_8 FILLER_30_2618 ();
 sg13g2_decap_8 FILLER_30_2625 ();
 sg13g2_decap_8 FILLER_30_2632 ();
 sg13g2_decap_8 FILLER_30_2639 ();
 sg13g2_decap_8 FILLER_30_2646 ();
 sg13g2_decap_8 FILLER_30_2653 ();
 sg13g2_decap_8 FILLER_30_2660 ();
 sg13g2_decap_8 FILLER_30_2667 ();
 sg13g2_decap_8 FILLER_30_2674 ();
 sg13g2_decap_8 FILLER_30_2681 ();
 sg13g2_decap_8 FILLER_30_2688 ();
 sg13g2_decap_8 FILLER_30_2695 ();
 sg13g2_decap_8 FILLER_30_2702 ();
 sg13g2_decap_8 FILLER_30_2709 ();
 sg13g2_decap_8 FILLER_30_2716 ();
 sg13g2_decap_8 FILLER_30_2723 ();
 sg13g2_decap_8 FILLER_30_2730 ();
 sg13g2_decap_8 FILLER_30_2737 ();
 sg13g2_decap_8 FILLER_30_2744 ();
 sg13g2_decap_8 FILLER_30_2751 ();
 sg13g2_decap_8 FILLER_30_2758 ();
 sg13g2_decap_8 FILLER_30_2765 ();
 sg13g2_decap_8 FILLER_30_2772 ();
 sg13g2_decap_8 FILLER_30_2779 ();
 sg13g2_decap_8 FILLER_30_2786 ();
 sg13g2_decap_8 FILLER_30_2793 ();
 sg13g2_decap_8 FILLER_30_2800 ();
 sg13g2_decap_8 FILLER_30_2807 ();
 sg13g2_decap_8 FILLER_30_2814 ();
 sg13g2_decap_8 FILLER_30_2821 ();
 sg13g2_decap_8 FILLER_30_2828 ();
 sg13g2_decap_8 FILLER_30_2835 ();
 sg13g2_decap_8 FILLER_30_2842 ();
 sg13g2_decap_8 FILLER_30_2849 ();
 sg13g2_decap_8 FILLER_30_2856 ();
 sg13g2_decap_8 FILLER_30_2863 ();
 sg13g2_decap_8 FILLER_30_2870 ();
 sg13g2_decap_8 FILLER_30_2877 ();
 sg13g2_decap_8 FILLER_30_2884 ();
 sg13g2_decap_8 FILLER_30_2891 ();
 sg13g2_decap_8 FILLER_30_2898 ();
 sg13g2_decap_8 FILLER_30_2905 ();
 sg13g2_decap_8 FILLER_30_2912 ();
 sg13g2_decap_8 FILLER_30_2919 ();
 sg13g2_decap_8 FILLER_30_2926 ();
 sg13g2_decap_8 FILLER_30_2933 ();
 sg13g2_decap_8 FILLER_30_2940 ();
 sg13g2_decap_8 FILLER_30_2947 ();
 sg13g2_decap_8 FILLER_30_2954 ();
 sg13g2_decap_8 FILLER_30_2961 ();
 sg13g2_decap_8 FILLER_30_2968 ();
 sg13g2_decap_8 FILLER_30_2975 ();
 sg13g2_decap_8 FILLER_30_2982 ();
 sg13g2_decap_8 FILLER_30_2989 ();
 sg13g2_decap_8 FILLER_30_2996 ();
 sg13g2_decap_8 FILLER_30_3003 ();
 sg13g2_decap_8 FILLER_30_3010 ();
 sg13g2_decap_8 FILLER_30_3017 ();
 sg13g2_decap_8 FILLER_30_3024 ();
 sg13g2_decap_8 FILLER_30_3031 ();
 sg13g2_decap_8 FILLER_30_3038 ();
 sg13g2_decap_8 FILLER_30_3045 ();
 sg13g2_decap_8 FILLER_30_3052 ();
 sg13g2_decap_8 FILLER_30_3059 ();
 sg13g2_decap_8 FILLER_30_3066 ();
 sg13g2_decap_8 FILLER_30_3073 ();
 sg13g2_decap_8 FILLER_30_3080 ();
 sg13g2_decap_8 FILLER_30_3087 ();
 sg13g2_decap_8 FILLER_30_3094 ();
 sg13g2_decap_8 FILLER_30_3101 ();
 sg13g2_decap_8 FILLER_30_3108 ();
 sg13g2_decap_8 FILLER_30_3115 ();
 sg13g2_decap_8 FILLER_30_3122 ();
 sg13g2_decap_8 FILLER_30_3129 ();
 sg13g2_decap_8 FILLER_30_3136 ();
 sg13g2_decap_8 FILLER_30_3143 ();
 sg13g2_decap_8 FILLER_30_3150 ();
 sg13g2_decap_8 FILLER_30_3157 ();
 sg13g2_decap_8 FILLER_30_3164 ();
 sg13g2_decap_8 FILLER_30_3171 ();
 sg13g2_decap_8 FILLER_30_3178 ();
 sg13g2_decap_8 FILLER_30_3185 ();
 sg13g2_decap_8 FILLER_30_3192 ();
 sg13g2_decap_8 FILLER_30_3199 ();
 sg13g2_decap_8 FILLER_30_3206 ();
 sg13g2_decap_8 FILLER_30_3213 ();
 sg13g2_decap_8 FILLER_30_3220 ();
 sg13g2_decap_8 FILLER_30_3227 ();
 sg13g2_decap_8 FILLER_30_3234 ();
 sg13g2_decap_8 FILLER_30_3241 ();
 sg13g2_decap_8 FILLER_30_3248 ();
 sg13g2_decap_8 FILLER_30_3255 ();
 sg13g2_decap_8 FILLER_30_3262 ();
 sg13g2_decap_8 FILLER_30_3269 ();
 sg13g2_decap_8 FILLER_30_3276 ();
 sg13g2_decap_8 FILLER_30_3283 ();
 sg13g2_decap_8 FILLER_30_3290 ();
 sg13g2_decap_8 FILLER_30_3297 ();
 sg13g2_decap_8 FILLER_30_3304 ();
 sg13g2_decap_8 FILLER_30_3311 ();
 sg13g2_decap_8 FILLER_30_3318 ();
 sg13g2_decap_8 FILLER_30_3325 ();
 sg13g2_decap_8 FILLER_30_3332 ();
 sg13g2_decap_8 FILLER_30_3339 ();
 sg13g2_decap_8 FILLER_30_3346 ();
 sg13g2_decap_8 FILLER_30_3353 ();
 sg13g2_decap_8 FILLER_30_3360 ();
 sg13g2_decap_8 FILLER_30_3367 ();
 sg13g2_decap_8 FILLER_30_3374 ();
 sg13g2_decap_8 FILLER_30_3381 ();
 sg13g2_decap_8 FILLER_30_3388 ();
 sg13g2_decap_8 FILLER_30_3395 ();
 sg13g2_decap_8 FILLER_30_3402 ();
 sg13g2_decap_8 FILLER_30_3409 ();
 sg13g2_decap_8 FILLER_30_3416 ();
 sg13g2_decap_8 FILLER_30_3423 ();
 sg13g2_decap_8 FILLER_30_3430 ();
 sg13g2_decap_8 FILLER_30_3437 ();
 sg13g2_decap_8 FILLER_30_3444 ();
 sg13g2_decap_8 FILLER_30_3451 ();
 sg13g2_decap_8 FILLER_30_3458 ();
 sg13g2_decap_8 FILLER_30_3465 ();
 sg13g2_decap_8 FILLER_30_3472 ();
 sg13g2_decap_8 FILLER_30_3479 ();
 sg13g2_decap_8 FILLER_30_3486 ();
 sg13g2_decap_8 FILLER_30_3493 ();
 sg13g2_decap_8 FILLER_30_3500 ();
 sg13g2_decap_8 FILLER_30_3507 ();
 sg13g2_decap_8 FILLER_30_3514 ();
 sg13g2_decap_8 FILLER_30_3521 ();
 sg13g2_decap_8 FILLER_30_3528 ();
 sg13g2_decap_8 FILLER_30_3535 ();
 sg13g2_decap_8 FILLER_30_3542 ();
 sg13g2_decap_8 FILLER_30_3549 ();
 sg13g2_decap_8 FILLER_30_3556 ();
 sg13g2_decap_8 FILLER_30_3563 ();
 sg13g2_decap_8 FILLER_30_3570 ();
 sg13g2_fill_2 FILLER_30_3577 ();
 sg13g2_fill_1 FILLER_30_3579 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_245 ();
 sg13g2_decap_8 FILLER_31_252 ();
 sg13g2_decap_8 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_266 ();
 sg13g2_decap_8 FILLER_31_273 ();
 sg13g2_decap_8 FILLER_31_280 ();
 sg13g2_decap_8 FILLER_31_287 ();
 sg13g2_decap_8 FILLER_31_294 ();
 sg13g2_decap_8 FILLER_31_301 ();
 sg13g2_decap_8 FILLER_31_308 ();
 sg13g2_decap_8 FILLER_31_315 ();
 sg13g2_decap_8 FILLER_31_322 ();
 sg13g2_decap_8 FILLER_31_329 ();
 sg13g2_decap_8 FILLER_31_336 ();
 sg13g2_decap_8 FILLER_31_343 ();
 sg13g2_decap_8 FILLER_31_350 ();
 sg13g2_decap_8 FILLER_31_357 ();
 sg13g2_decap_8 FILLER_31_364 ();
 sg13g2_decap_8 FILLER_31_371 ();
 sg13g2_decap_8 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_385 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_decap_8 FILLER_31_406 ();
 sg13g2_decap_8 FILLER_31_413 ();
 sg13g2_decap_8 FILLER_31_420 ();
 sg13g2_decap_8 FILLER_31_427 ();
 sg13g2_decap_8 FILLER_31_434 ();
 sg13g2_decap_8 FILLER_31_441 ();
 sg13g2_decap_8 FILLER_31_448 ();
 sg13g2_decap_8 FILLER_31_455 ();
 sg13g2_decap_8 FILLER_31_462 ();
 sg13g2_decap_8 FILLER_31_469 ();
 sg13g2_decap_8 FILLER_31_476 ();
 sg13g2_decap_8 FILLER_31_483 ();
 sg13g2_decap_8 FILLER_31_490 ();
 sg13g2_decap_8 FILLER_31_497 ();
 sg13g2_decap_8 FILLER_31_504 ();
 sg13g2_decap_8 FILLER_31_511 ();
 sg13g2_decap_8 FILLER_31_518 ();
 sg13g2_decap_8 FILLER_31_525 ();
 sg13g2_decap_8 FILLER_31_532 ();
 sg13g2_decap_8 FILLER_31_539 ();
 sg13g2_decap_8 FILLER_31_546 ();
 sg13g2_decap_8 FILLER_31_553 ();
 sg13g2_decap_8 FILLER_31_560 ();
 sg13g2_decap_8 FILLER_31_567 ();
 sg13g2_decap_8 FILLER_31_574 ();
 sg13g2_decap_8 FILLER_31_581 ();
 sg13g2_decap_8 FILLER_31_588 ();
 sg13g2_decap_8 FILLER_31_595 ();
 sg13g2_decap_8 FILLER_31_602 ();
 sg13g2_decap_8 FILLER_31_609 ();
 sg13g2_decap_8 FILLER_31_616 ();
 sg13g2_decap_8 FILLER_31_623 ();
 sg13g2_decap_8 FILLER_31_630 ();
 sg13g2_decap_8 FILLER_31_637 ();
 sg13g2_decap_8 FILLER_31_644 ();
 sg13g2_decap_8 FILLER_31_651 ();
 sg13g2_decap_8 FILLER_31_658 ();
 sg13g2_decap_8 FILLER_31_665 ();
 sg13g2_decap_8 FILLER_31_672 ();
 sg13g2_decap_8 FILLER_31_679 ();
 sg13g2_decap_8 FILLER_31_686 ();
 sg13g2_decap_8 FILLER_31_693 ();
 sg13g2_decap_8 FILLER_31_700 ();
 sg13g2_decap_8 FILLER_31_707 ();
 sg13g2_decap_8 FILLER_31_714 ();
 sg13g2_decap_8 FILLER_31_721 ();
 sg13g2_decap_8 FILLER_31_728 ();
 sg13g2_decap_8 FILLER_31_735 ();
 sg13g2_decap_8 FILLER_31_742 ();
 sg13g2_decap_8 FILLER_31_749 ();
 sg13g2_decap_8 FILLER_31_756 ();
 sg13g2_decap_8 FILLER_31_763 ();
 sg13g2_decap_8 FILLER_31_770 ();
 sg13g2_decap_8 FILLER_31_777 ();
 sg13g2_decap_8 FILLER_31_784 ();
 sg13g2_decap_8 FILLER_31_791 ();
 sg13g2_decap_8 FILLER_31_798 ();
 sg13g2_decap_8 FILLER_31_805 ();
 sg13g2_decap_8 FILLER_31_812 ();
 sg13g2_decap_8 FILLER_31_819 ();
 sg13g2_decap_8 FILLER_31_826 ();
 sg13g2_decap_8 FILLER_31_833 ();
 sg13g2_decap_8 FILLER_31_840 ();
 sg13g2_decap_8 FILLER_31_847 ();
 sg13g2_decap_8 FILLER_31_854 ();
 sg13g2_decap_8 FILLER_31_861 ();
 sg13g2_decap_8 FILLER_31_868 ();
 sg13g2_decap_8 FILLER_31_875 ();
 sg13g2_decap_8 FILLER_31_882 ();
 sg13g2_decap_8 FILLER_31_889 ();
 sg13g2_decap_8 FILLER_31_896 ();
 sg13g2_decap_8 FILLER_31_903 ();
 sg13g2_decap_8 FILLER_31_910 ();
 sg13g2_decap_8 FILLER_31_917 ();
 sg13g2_decap_8 FILLER_31_924 ();
 sg13g2_decap_8 FILLER_31_931 ();
 sg13g2_decap_8 FILLER_31_938 ();
 sg13g2_decap_8 FILLER_31_945 ();
 sg13g2_decap_8 FILLER_31_952 ();
 sg13g2_decap_8 FILLER_31_959 ();
 sg13g2_decap_8 FILLER_31_966 ();
 sg13g2_decap_8 FILLER_31_973 ();
 sg13g2_decap_8 FILLER_31_980 ();
 sg13g2_decap_8 FILLER_31_987 ();
 sg13g2_decap_8 FILLER_31_994 ();
 sg13g2_decap_8 FILLER_31_1001 ();
 sg13g2_decap_8 FILLER_31_1008 ();
 sg13g2_decap_8 FILLER_31_1015 ();
 sg13g2_decap_8 FILLER_31_1022 ();
 sg13g2_decap_8 FILLER_31_1029 ();
 sg13g2_decap_8 FILLER_31_1036 ();
 sg13g2_decap_8 FILLER_31_1043 ();
 sg13g2_decap_8 FILLER_31_1050 ();
 sg13g2_decap_8 FILLER_31_1057 ();
 sg13g2_decap_8 FILLER_31_1064 ();
 sg13g2_decap_8 FILLER_31_1071 ();
 sg13g2_decap_8 FILLER_31_1078 ();
 sg13g2_decap_8 FILLER_31_1085 ();
 sg13g2_decap_8 FILLER_31_1092 ();
 sg13g2_decap_8 FILLER_31_1099 ();
 sg13g2_decap_8 FILLER_31_1106 ();
 sg13g2_decap_8 FILLER_31_1113 ();
 sg13g2_decap_8 FILLER_31_1120 ();
 sg13g2_decap_8 FILLER_31_1127 ();
 sg13g2_decap_8 FILLER_31_1134 ();
 sg13g2_decap_8 FILLER_31_1141 ();
 sg13g2_decap_8 FILLER_31_1148 ();
 sg13g2_decap_8 FILLER_31_1155 ();
 sg13g2_decap_8 FILLER_31_1162 ();
 sg13g2_decap_8 FILLER_31_1169 ();
 sg13g2_decap_8 FILLER_31_1176 ();
 sg13g2_decap_8 FILLER_31_1183 ();
 sg13g2_decap_8 FILLER_31_1190 ();
 sg13g2_decap_8 FILLER_31_1197 ();
 sg13g2_decap_8 FILLER_31_1204 ();
 sg13g2_decap_8 FILLER_31_1211 ();
 sg13g2_decap_8 FILLER_31_1218 ();
 sg13g2_decap_8 FILLER_31_1225 ();
 sg13g2_decap_8 FILLER_31_1232 ();
 sg13g2_decap_8 FILLER_31_1239 ();
 sg13g2_decap_8 FILLER_31_1246 ();
 sg13g2_decap_8 FILLER_31_1253 ();
 sg13g2_decap_8 FILLER_31_1260 ();
 sg13g2_decap_8 FILLER_31_1267 ();
 sg13g2_decap_8 FILLER_31_1274 ();
 sg13g2_decap_8 FILLER_31_1281 ();
 sg13g2_decap_8 FILLER_31_1288 ();
 sg13g2_decap_8 FILLER_31_1295 ();
 sg13g2_decap_8 FILLER_31_1302 ();
 sg13g2_decap_8 FILLER_31_1309 ();
 sg13g2_decap_8 FILLER_31_1316 ();
 sg13g2_decap_8 FILLER_31_1323 ();
 sg13g2_decap_8 FILLER_31_1330 ();
 sg13g2_decap_8 FILLER_31_1337 ();
 sg13g2_decap_8 FILLER_31_1344 ();
 sg13g2_decap_8 FILLER_31_1351 ();
 sg13g2_decap_8 FILLER_31_1358 ();
 sg13g2_decap_8 FILLER_31_1365 ();
 sg13g2_decap_8 FILLER_31_1372 ();
 sg13g2_decap_8 FILLER_31_1379 ();
 sg13g2_decap_8 FILLER_31_1386 ();
 sg13g2_decap_8 FILLER_31_1393 ();
 sg13g2_decap_8 FILLER_31_1400 ();
 sg13g2_decap_8 FILLER_31_1407 ();
 sg13g2_decap_8 FILLER_31_1414 ();
 sg13g2_decap_8 FILLER_31_1421 ();
 sg13g2_decap_8 FILLER_31_1428 ();
 sg13g2_decap_8 FILLER_31_1435 ();
 sg13g2_decap_8 FILLER_31_1442 ();
 sg13g2_decap_8 FILLER_31_1449 ();
 sg13g2_decap_8 FILLER_31_1456 ();
 sg13g2_decap_8 FILLER_31_1463 ();
 sg13g2_decap_8 FILLER_31_1470 ();
 sg13g2_decap_8 FILLER_31_1477 ();
 sg13g2_decap_8 FILLER_31_1484 ();
 sg13g2_decap_8 FILLER_31_1491 ();
 sg13g2_decap_8 FILLER_31_1498 ();
 sg13g2_decap_8 FILLER_31_1505 ();
 sg13g2_decap_8 FILLER_31_1512 ();
 sg13g2_decap_8 FILLER_31_1519 ();
 sg13g2_decap_8 FILLER_31_1526 ();
 sg13g2_decap_8 FILLER_31_1533 ();
 sg13g2_decap_8 FILLER_31_1540 ();
 sg13g2_decap_8 FILLER_31_1547 ();
 sg13g2_decap_8 FILLER_31_1554 ();
 sg13g2_decap_8 FILLER_31_1561 ();
 sg13g2_decap_8 FILLER_31_1568 ();
 sg13g2_decap_8 FILLER_31_1575 ();
 sg13g2_decap_8 FILLER_31_1582 ();
 sg13g2_decap_8 FILLER_31_1589 ();
 sg13g2_decap_8 FILLER_31_1596 ();
 sg13g2_decap_8 FILLER_31_1603 ();
 sg13g2_decap_8 FILLER_31_1610 ();
 sg13g2_decap_8 FILLER_31_1617 ();
 sg13g2_decap_8 FILLER_31_1624 ();
 sg13g2_decap_8 FILLER_31_1631 ();
 sg13g2_decap_8 FILLER_31_1638 ();
 sg13g2_decap_8 FILLER_31_1645 ();
 sg13g2_decap_8 FILLER_31_1652 ();
 sg13g2_decap_8 FILLER_31_1659 ();
 sg13g2_decap_8 FILLER_31_1666 ();
 sg13g2_decap_8 FILLER_31_1673 ();
 sg13g2_decap_8 FILLER_31_1680 ();
 sg13g2_decap_8 FILLER_31_1687 ();
 sg13g2_decap_8 FILLER_31_1694 ();
 sg13g2_decap_8 FILLER_31_1701 ();
 sg13g2_decap_8 FILLER_31_1708 ();
 sg13g2_decap_8 FILLER_31_1715 ();
 sg13g2_decap_8 FILLER_31_1722 ();
 sg13g2_decap_8 FILLER_31_1729 ();
 sg13g2_decap_8 FILLER_31_1736 ();
 sg13g2_decap_8 FILLER_31_1743 ();
 sg13g2_decap_8 FILLER_31_1750 ();
 sg13g2_decap_8 FILLER_31_1757 ();
 sg13g2_decap_8 FILLER_31_1764 ();
 sg13g2_decap_8 FILLER_31_1771 ();
 sg13g2_decap_8 FILLER_31_1778 ();
 sg13g2_decap_8 FILLER_31_1785 ();
 sg13g2_decap_8 FILLER_31_1792 ();
 sg13g2_decap_8 FILLER_31_1799 ();
 sg13g2_decap_8 FILLER_31_1806 ();
 sg13g2_decap_8 FILLER_31_1813 ();
 sg13g2_decap_8 FILLER_31_1820 ();
 sg13g2_decap_8 FILLER_31_1827 ();
 sg13g2_decap_8 FILLER_31_1834 ();
 sg13g2_decap_8 FILLER_31_1841 ();
 sg13g2_decap_8 FILLER_31_1848 ();
 sg13g2_decap_8 FILLER_31_1855 ();
 sg13g2_decap_8 FILLER_31_1862 ();
 sg13g2_decap_8 FILLER_31_1869 ();
 sg13g2_decap_8 FILLER_31_1876 ();
 sg13g2_decap_8 FILLER_31_1883 ();
 sg13g2_decap_8 FILLER_31_1890 ();
 sg13g2_decap_8 FILLER_31_1897 ();
 sg13g2_decap_8 FILLER_31_1904 ();
 sg13g2_decap_8 FILLER_31_1911 ();
 sg13g2_decap_8 FILLER_31_1918 ();
 sg13g2_decap_8 FILLER_31_1925 ();
 sg13g2_decap_8 FILLER_31_1932 ();
 sg13g2_decap_8 FILLER_31_1939 ();
 sg13g2_decap_8 FILLER_31_1946 ();
 sg13g2_decap_8 FILLER_31_1953 ();
 sg13g2_decap_8 FILLER_31_1960 ();
 sg13g2_decap_8 FILLER_31_1967 ();
 sg13g2_decap_8 FILLER_31_1974 ();
 sg13g2_decap_8 FILLER_31_1981 ();
 sg13g2_decap_8 FILLER_31_1988 ();
 sg13g2_decap_8 FILLER_31_1995 ();
 sg13g2_decap_8 FILLER_31_2002 ();
 sg13g2_decap_8 FILLER_31_2009 ();
 sg13g2_decap_8 FILLER_31_2016 ();
 sg13g2_decap_8 FILLER_31_2023 ();
 sg13g2_decap_8 FILLER_31_2030 ();
 sg13g2_decap_8 FILLER_31_2037 ();
 sg13g2_decap_8 FILLER_31_2044 ();
 sg13g2_decap_8 FILLER_31_2051 ();
 sg13g2_decap_8 FILLER_31_2058 ();
 sg13g2_decap_8 FILLER_31_2065 ();
 sg13g2_decap_8 FILLER_31_2072 ();
 sg13g2_decap_8 FILLER_31_2079 ();
 sg13g2_decap_8 FILLER_31_2086 ();
 sg13g2_decap_8 FILLER_31_2093 ();
 sg13g2_decap_8 FILLER_31_2100 ();
 sg13g2_decap_8 FILLER_31_2107 ();
 sg13g2_decap_8 FILLER_31_2114 ();
 sg13g2_decap_8 FILLER_31_2121 ();
 sg13g2_decap_8 FILLER_31_2128 ();
 sg13g2_decap_8 FILLER_31_2135 ();
 sg13g2_decap_8 FILLER_31_2142 ();
 sg13g2_decap_8 FILLER_31_2149 ();
 sg13g2_decap_8 FILLER_31_2156 ();
 sg13g2_decap_8 FILLER_31_2163 ();
 sg13g2_decap_8 FILLER_31_2170 ();
 sg13g2_decap_8 FILLER_31_2177 ();
 sg13g2_decap_8 FILLER_31_2184 ();
 sg13g2_decap_8 FILLER_31_2191 ();
 sg13g2_decap_8 FILLER_31_2198 ();
 sg13g2_decap_8 FILLER_31_2205 ();
 sg13g2_decap_8 FILLER_31_2212 ();
 sg13g2_decap_8 FILLER_31_2219 ();
 sg13g2_decap_8 FILLER_31_2226 ();
 sg13g2_decap_8 FILLER_31_2233 ();
 sg13g2_decap_8 FILLER_31_2240 ();
 sg13g2_decap_8 FILLER_31_2247 ();
 sg13g2_decap_8 FILLER_31_2254 ();
 sg13g2_decap_8 FILLER_31_2261 ();
 sg13g2_decap_8 FILLER_31_2268 ();
 sg13g2_decap_8 FILLER_31_2275 ();
 sg13g2_decap_8 FILLER_31_2282 ();
 sg13g2_decap_8 FILLER_31_2289 ();
 sg13g2_decap_8 FILLER_31_2296 ();
 sg13g2_decap_8 FILLER_31_2303 ();
 sg13g2_decap_8 FILLER_31_2310 ();
 sg13g2_decap_8 FILLER_31_2317 ();
 sg13g2_decap_8 FILLER_31_2324 ();
 sg13g2_decap_8 FILLER_31_2331 ();
 sg13g2_decap_8 FILLER_31_2338 ();
 sg13g2_decap_8 FILLER_31_2345 ();
 sg13g2_decap_8 FILLER_31_2352 ();
 sg13g2_decap_8 FILLER_31_2359 ();
 sg13g2_decap_8 FILLER_31_2366 ();
 sg13g2_decap_8 FILLER_31_2373 ();
 sg13g2_decap_8 FILLER_31_2380 ();
 sg13g2_decap_8 FILLER_31_2387 ();
 sg13g2_decap_8 FILLER_31_2394 ();
 sg13g2_decap_8 FILLER_31_2401 ();
 sg13g2_decap_8 FILLER_31_2408 ();
 sg13g2_decap_8 FILLER_31_2415 ();
 sg13g2_decap_8 FILLER_31_2422 ();
 sg13g2_decap_8 FILLER_31_2429 ();
 sg13g2_decap_8 FILLER_31_2436 ();
 sg13g2_decap_8 FILLER_31_2443 ();
 sg13g2_decap_8 FILLER_31_2450 ();
 sg13g2_decap_8 FILLER_31_2457 ();
 sg13g2_decap_8 FILLER_31_2464 ();
 sg13g2_decap_8 FILLER_31_2471 ();
 sg13g2_decap_8 FILLER_31_2478 ();
 sg13g2_decap_8 FILLER_31_2485 ();
 sg13g2_decap_8 FILLER_31_2492 ();
 sg13g2_decap_8 FILLER_31_2499 ();
 sg13g2_decap_8 FILLER_31_2506 ();
 sg13g2_decap_8 FILLER_31_2513 ();
 sg13g2_decap_8 FILLER_31_2520 ();
 sg13g2_decap_8 FILLER_31_2527 ();
 sg13g2_decap_8 FILLER_31_2534 ();
 sg13g2_decap_8 FILLER_31_2541 ();
 sg13g2_decap_8 FILLER_31_2548 ();
 sg13g2_decap_8 FILLER_31_2555 ();
 sg13g2_decap_8 FILLER_31_2562 ();
 sg13g2_decap_8 FILLER_31_2569 ();
 sg13g2_decap_8 FILLER_31_2576 ();
 sg13g2_decap_8 FILLER_31_2583 ();
 sg13g2_decap_8 FILLER_31_2590 ();
 sg13g2_decap_8 FILLER_31_2597 ();
 sg13g2_decap_8 FILLER_31_2604 ();
 sg13g2_decap_8 FILLER_31_2611 ();
 sg13g2_decap_8 FILLER_31_2618 ();
 sg13g2_decap_8 FILLER_31_2625 ();
 sg13g2_decap_8 FILLER_31_2632 ();
 sg13g2_decap_8 FILLER_31_2639 ();
 sg13g2_decap_8 FILLER_31_2646 ();
 sg13g2_decap_8 FILLER_31_2653 ();
 sg13g2_decap_8 FILLER_31_2660 ();
 sg13g2_decap_8 FILLER_31_2667 ();
 sg13g2_decap_8 FILLER_31_2674 ();
 sg13g2_decap_8 FILLER_31_2681 ();
 sg13g2_decap_8 FILLER_31_2688 ();
 sg13g2_decap_8 FILLER_31_2695 ();
 sg13g2_decap_8 FILLER_31_2702 ();
 sg13g2_decap_8 FILLER_31_2709 ();
 sg13g2_decap_8 FILLER_31_2716 ();
 sg13g2_decap_8 FILLER_31_2723 ();
 sg13g2_decap_8 FILLER_31_2730 ();
 sg13g2_decap_8 FILLER_31_2737 ();
 sg13g2_decap_8 FILLER_31_2744 ();
 sg13g2_decap_8 FILLER_31_2751 ();
 sg13g2_decap_8 FILLER_31_2758 ();
 sg13g2_decap_8 FILLER_31_2765 ();
 sg13g2_decap_8 FILLER_31_2772 ();
 sg13g2_decap_8 FILLER_31_2779 ();
 sg13g2_decap_8 FILLER_31_2786 ();
 sg13g2_decap_8 FILLER_31_2793 ();
 sg13g2_decap_8 FILLER_31_2800 ();
 sg13g2_decap_8 FILLER_31_2807 ();
 sg13g2_decap_8 FILLER_31_2814 ();
 sg13g2_decap_8 FILLER_31_2821 ();
 sg13g2_decap_8 FILLER_31_2828 ();
 sg13g2_decap_8 FILLER_31_2835 ();
 sg13g2_decap_8 FILLER_31_2842 ();
 sg13g2_decap_8 FILLER_31_2849 ();
 sg13g2_decap_8 FILLER_31_2856 ();
 sg13g2_decap_8 FILLER_31_2863 ();
 sg13g2_decap_8 FILLER_31_2870 ();
 sg13g2_decap_8 FILLER_31_2877 ();
 sg13g2_decap_8 FILLER_31_2884 ();
 sg13g2_decap_8 FILLER_31_2891 ();
 sg13g2_decap_8 FILLER_31_2898 ();
 sg13g2_decap_8 FILLER_31_2905 ();
 sg13g2_decap_8 FILLER_31_2912 ();
 sg13g2_decap_8 FILLER_31_2919 ();
 sg13g2_decap_8 FILLER_31_2926 ();
 sg13g2_decap_8 FILLER_31_2933 ();
 sg13g2_decap_8 FILLER_31_2940 ();
 sg13g2_decap_8 FILLER_31_2947 ();
 sg13g2_decap_8 FILLER_31_2954 ();
 sg13g2_decap_8 FILLER_31_2961 ();
 sg13g2_decap_8 FILLER_31_2968 ();
 sg13g2_decap_8 FILLER_31_2975 ();
 sg13g2_decap_8 FILLER_31_2982 ();
 sg13g2_decap_8 FILLER_31_2989 ();
 sg13g2_decap_8 FILLER_31_2996 ();
 sg13g2_decap_8 FILLER_31_3003 ();
 sg13g2_decap_8 FILLER_31_3010 ();
 sg13g2_decap_8 FILLER_31_3017 ();
 sg13g2_decap_8 FILLER_31_3024 ();
 sg13g2_decap_8 FILLER_31_3031 ();
 sg13g2_decap_8 FILLER_31_3038 ();
 sg13g2_decap_8 FILLER_31_3045 ();
 sg13g2_decap_8 FILLER_31_3052 ();
 sg13g2_decap_8 FILLER_31_3059 ();
 sg13g2_decap_8 FILLER_31_3066 ();
 sg13g2_decap_8 FILLER_31_3073 ();
 sg13g2_decap_8 FILLER_31_3080 ();
 sg13g2_decap_8 FILLER_31_3087 ();
 sg13g2_decap_8 FILLER_31_3094 ();
 sg13g2_decap_8 FILLER_31_3101 ();
 sg13g2_decap_8 FILLER_31_3108 ();
 sg13g2_decap_8 FILLER_31_3115 ();
 sg13g2_decap_8 FILLER_31_3122 ();
 sg13g2_decap_8 FILLER_31_3129 ();
 sg13g2_decap_8 FILLER_31_3136 ();
 sg13g2_decap_8 FILLER_31_3143 ();
 sg13g2_decap_8 FILLER_31_3150 ();
 sg13g2_decap_8 FILLER_31_3157 ();
 sg13g2_decap_8 FILLER_31_3164 ();
 sg13g2_decap_8 FILLER_31_3171 ();
 sg13g2_decap_8 FILLER_31_3178 ();
 sg13g2_decap_8 FILLER_31_3185 ();
 sg13g2_decap_8 FILLER_31_3192 ();
 sg13g2_decap_8 FILLER_31_3199 ();
 sg13g2_decap_8 FILLER_31_3206 ();
 sg13g2_decap_8 FILLER_31_3213 ();
 sg13g2_decap_8 FILLER_31_3220 ();
 sg13g2_decap_8 FILLER_31_3227 ();
 sg13g2_decap_8 FILLER_31_3234 ();
 sg13g2_decap_8 FILLER_31_3241 ();
 sg13g2_decap_8 FILLER_31_3248 ();
 sg13g2_decap_8 FILLER_31_3255 ();
 sg13g2_decap_8 FILLER_31_3262 ();
 sg13g2_decap_8 FILLER_31_3269 ();
 sg13g2_decap_8 FILLER_31_3276 ();
 sg13g2_decap_8 FILLER_31_3283 ();
 sg13g2_decap_8 FILLER_31_3290 ();
 sg13g2_decap_8 FILLER_31_3297 ();
 sg13g2_decap_8 FILLER_31_3304 ();
 sg13g2_decap_8 FILLER_31_3311 ();
 sg13g2_decap_8 FILLER_31_3318 ();
 sg13g2_decap_8 FILLER_31_3325 ();
 sg13g2_decap_8 FILLER_31_3332 ();
 sg13g2_decap_8 FILLER_31_3339 ();
 sg13g2_decap_8 FILLER_31_3346 ();
 sg13g2_decap_8 FILLER_31_3353 ();
 sg13g2_decap_8 FILLER_31_3360 ();
 sg13g2_decap_8 FILLER_31_3367 ();
 sg13g2_decap_8 FILLER_31_3374 ();
 sg13g2_decap_8 FILLER_31_3381 ();
 sg13g2_decap_8 FILLER_31_3388 ();
 sg13g2_decap_8 FILLER_31_3395 ();
 sg13g2_decap_8 FILLER_31_3402 ();
 sg13g2_decap_8 FILLER_31_3409 ();
 sg13g2_decap_8 FILLER_31_3416 ();
 sg13g2_decap_8 FILLER_31_3423 ();
 sg13g2_decap_8 FILLER_31_3430 ();
 sg13g2_decap_8 FILLER_31_3437 ();
 sg13g2_decap_8 FILLER_31_3444 ();
 sg13g2_decap_8 FILLER_31_3451 ();
 sg13g2_decap_8 FILLER_31_3458 ();
 sg13g2_decap_8 FILLER_31_3465 ();
 sg13g2_decap_8 FILLER_31_3472 ();
 sg13g2_decap_8 FILLER_31_3479 ();
 sg13g2_decap_8 FILLER_31_3486 ();
 sg13g2_decap_8 FILLER_31_3493 ();
 sg13g2_decap_8 FILLER_31_3500 ();
 sg13g2_decap_8 FILLER_31_3507 ();
 sg13g2_decap_8 FILLER_31_3514 ();
 sg13g2_decap_8 FILLER_31_3521 ();
 sg13g2_decap_8 FILLER_31_3528 ();
 sg13g2_decap_8 FILLER_31_3535 ();
 sg13g2_decap_8 FILLER_31_3542 ();
 sg13g2_decap_8 FILLER_31_3549 ();
 sg13g2_decap_8 FILLER_31_3556 ();
 sg13g2_decap_8 FILLER_31_3563 ();
 sg13g2_decap_8 FILLER_31_3570 ();
 sg13g2_fill_2 FILLER_31_3577 ();
 sg13g2_fill_1 FILLER_31_3579 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_231 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_decap_8 FILLER_32_245 ();
 sg13g2_decap_8 FILLER_32_252 ();
 sg13g2_decap_8 FILLER_32_259 ();
 sg13g2_decap_8 FILLER_32_266 ();
 sg13g2_decap_8 FILLER_32_273 ();
 sg13g2_decap_8 FILLER_32_280 ();
 sg13g2_decap_8 FILLER_32_287 ();
 sg13g2_decap_8 FILLER_32_294 ();
 sg13g2_decap_8 FILLER_32_301 ();
 sg13g2_decap_8 FILLER_32_308 ();
 sg13g2_decap_8 FILLER_32_315 ();
 sg13g2_decap_8 FILLER_32_322 ();
 sg13g2_decap_8 FILLER_32_329 ();
 sg13g2_decap_8 FILLER_32_336 ();
 sg13g2_decap_8 FILLER_32_343 ();
 sg13g2_decap_8 FILLER_32_350 ();
 sg13g2_decap_8 FILLER_32_357 ();
 sg13g2_decap_8 FILLER_32_364 ();
 sg13g2_decap_8 FILLER_32_371 ();
 sg13g2_decap_8 FILLER_32_378 ();
 sg13g2_decap_8 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_decap_8 FILLER_32_406 ();
 sg13g2_decap_8 FILLER_32_413 ();
 sg13g2_decap_8 FILLER_32_420 ();
 sg13g2_decap_8 FILLER_32_427 ();
 sg13g2_decap_8 FILLER_32_434 ();
 sg13g2_decap_8 FILLER_32_441 ();
 sg13g2_decap_8 FILLER_32_448 ();
 sg13g2_decap_8 FILLER_32_455 ();
 sg13g2_decap_8 FILLER_32_462 ();
 sg13g2_decap_8 FILLER_32_469 ();
 sg13g2_decap_8 FILLER_32_476 ();
 sg13g2_decap_8 FILLER_32_483 ();
 sg13g2_decap_8 FILLER_32_490 ();
 sg13g2_decap_8 FILLER_32_497 ();
 sg13g2_decap_8 FILLER_32_504 ();
 sg13g2_decap_8 FILLER_32_511 ();
 sg13g2_decap_8 FILLER_32_518 ();
 sg13g2_decap_8 FILLER_32_525 ();
 sg13g2_decap_8 FILLER_32_532 ();
 sg13g2_decap_8 FILLER_32_539 ();
 sg13g2_decap_8 FILLER_32_546 ();
 sg13g2_decap_8 FILLER_32_553 ();
 sg13g2_decap_8 FILLER_32_560 ();
 sg13g2_decap_8 FILLER_32_567 ();
 sg13g2_decap_8 FILLER_32_574 ();
 sg13g2_decap_8 FILLER_32_581 ();
 sg13g2_decap_8 FILLER_32_588 ();
 sg13g2_decap_8 FILLER_32_595 ();
 sg13g2_decap_8 FILLER_32_602 ();
 sg13g2_decap_8 FILLER_32_609 ();
 sg13g2_decap_8 FILLER_32_616 ();
 sg13g2_decap_8 FILLER_32_623 ();
 sg13g2_decap_8 FILLER_32_630 ();
 sg13g2_decap_8 FILLER_32_637 ();
 sg13g2_decap_8 FILLER_32_644 ();
 sg13g2_decap_8 FILLER_32_651 ();
 sg13g2_decap_8 FILLER_32_658 ();
 sg13g2_decap_8 FILLER_32_665 ();
 sg13g2_decap_8 FILLER_32_672 ();
 sg13g2_decap_8 FILLER_32_679 ();
 sg13g2_decap_8 FILLER_32_686 ();
 sg13g2_decap_8 FILLER_32_693 ();
 sg13g2_decap_8 FILLER_32_700 ();
 sg13g2_decap_8 FILLER_32_707 ();
 sg13g2_decap_8 FILLER_32_714 ();
 sg13g2_decap_8 FILLER_32_721 ();
 sg13g2_decap_8 FILLER_32_728 ();
 sg13g2_decap_8 FILLER_32_735 ();
 sg13g2_decap_8 FILLER_32_742 ();
 sg13g2_decap_8 FILLER_32_749 ();
 sg13g2_decap_8 FILLER_32_756 ();
 sg13g2_decap_8 FILLER_32_763 ();
 sg13g2_decap_8 FILLER_32_770 ();
 sg13g2_decap_8 FILLER_32_777 ();
 sg13g2_decap_8 FILLER_32_784 ();
 sg13g2_decap_8 FILLER_32_791 ();
 sg13g2_decap_8 FILLER_32_798 ();
 sg13g2_decap_8 FILLER_32_805 ();
 sg13g2_decap_8 FILLER_32_812 ();
 sg13g2_decap_8 FILLER_32_819 ();
 sg13g2_decap_8 FILLER_32_826 ();
 sg13g2_decap_8 FILLER_32_833 ();
 sg13g2_decap_8 FILLER_32_840 ();
 sg13g2_decap_8 FILLER_32_847 ();
 sg13g2_decap_8 FILLER_32_854 ();
 sg13g2_decap_8 FILLER_32_861 ();
 sg13g2_decap_8 FILLER_32_868 ();
 sg13g2_decap_8 FILLER_32_875 ();
 sg13g2_decap_8 FILLER_32_882 ();
 sg13g2_decap_8 FILLER_32_889 ();
 sg13g2_decap_8 FILLER_32_896 ();
 sg13g2_decap_8 FILLER_32_903 ();
 sg13g2_decap_8 FILLER_32_910 ();
 sg13g2_decap_8 FILLER_32_917 ();
 sg13g2_decap_8 FILLER_32_924 ();
 sg13g2_decap_8 FILLER_32_931 ();
 sg13g2_decap_8 FILLER_32_938 ();
 sg13g2_decap_8 FILLER_32_945 ();
 sg13g2_decap_8 FILLER_32_952 ();
 sg13g2_decap_8 FILLER_32_959 ();
 sg13g2_decap_8 FILLER_32_966 ();
 sg13g2_decap_8 FILLER_32_973 ();
 sg13g2_decap_8 FILLER_32_980 ();
 sg13g2_decap_8 FILLER_32_987 ();
 sg13g2_decap_8 FILLER_32_994 ();
 sg13g2_decap_8 FILLER_32_1001 ();
 sg13g2_decap_8 FILLER_32_1008 ();
 sg13g2_decap_8 FILLER_32_1015 ();
 sg13g2_decap_8 FILLER_32_1022 ();
 sg13g2_decap_8 FILLER_32_1029 ();
 sg13g2_decap_8 FILLER_32_1036 ();
 sg13g2_decap_8 FILLER_32_1043 ();
 sg13g2_decap_8 FILLER_32_1050 ();
 sg13g2_decap_8 FILLER_32_1057 ();
 sg13g2_decap_8 FILLER_32_1064 ();
 sg13g2_decap_8 FILLER_32_1071 ();
 sg13g2_decap_8 FILLER_32_1078 ();
 sg13g2_decap_8 FILLER_32_1085 ();
 sg13g2_decap_8 FILLER_32_1092 ();
 sg13g2_decap_8 FILLER_32_1099 ();
 sg13g2_decap_8 FILLER_32_1106 ();
 sg13g2_decap_8 FILLER_32_1113 ();
 sg13g2_decap_8 FILLER_32_1120 ();
 sg13g2_decap_8 FILLER_32_1127 ();
 sg13g2_decap_8 FILLER_32_1134 ();
 sg13g2_decap_8 FILLER_32_1141 ();
 sg13g2_decap_8 FILLER_32_1148 ();
 sg13g2_decap_8 FILLER_32_1155 ();
 sg13g2_decap_8 FILLER_32_1162 ();
 sg13g2_decap_8 FILLER_32_1169 ();
 sg13g2_decap_8 FILLER_32_1176 ();
 sg13g2_decap_8 FILLER_32_1183 ();
 sg13g2_decap_8 FILLER_32_1190 ();
 sg13g2_decap_8 FILLER_32_1197 ();
 sg13g2_decap_8 FILLER_32_1204 ();
 sg13g2_decap_8 FILLER_32_1211 ();
 sg13g2_decap_8 FILLER_32_1218 ();
 sg13g2_decap_8 FILLER_32_1225 ();
 sg13g2_decap_8 FILLER_32_1232 ();
 sg13g2_decap_8 FILLER_32_1239 ();
 sg13g2_decap_8 FILLER_32_1246 ();
 sg13g2_decap_8 FILLER_32_1253 ();
 sg13g2_decap_8 FILLER_32_1260 ();
 sg13g2_decap_8 FILLER_32_1267 ();
 sg13g2_decap_8 FILLER_32_1274 ();
 sg13g2_decap_8 FILLER_32_1281 ();
 sg13g2_decap_8 FILLER_32_1288 ();
 sg13g2_decap_8 FILLER_32_1295 ();
 sg13g2_decap_8 FILLER_32_1302 ();
 sg13g2_decap_8 FILLER_32_1309 ();
 sg13g2_decap_8 FILLER_32_1316 ();
 sg13g2_decap_8 FILLER_32_1323 ();
 sg13g2_decap_8 FILLER_32_1330 ();
 sg13g2_decap_8 FILLER_32_1337 ();
 sg13g2_decap_8 FILLER_32_1344 ();
 sg13g2_decap_8 FILLER_32_1351 ();
 sg13g2_decap_8 FILLER_32_1358 ();
 sg13g2_decap_8 FILLER_32_1365 ();
 sg13g2_decap_8 FILLER_32_1372 ();
 sg13g2_decap_8 FILLER_32_1379 ();
 sg13g2_decap_8 FILLER_32_1386 ();
 sg13g2_decap_8 FILLER_32_1393 ();
 sg13g2_decap_8 FILLER_32_1400 ();
 sg13g2_decap_8 FILLER_32_1407 ();
 sg13g2_decap_8 FILLER_32_1414 ();
 sg13g2_decap_8 FILLER_32_1421 ();
 sg13g2_decap_8 FILLER_32_1428 ();
 sg13g2_decap_8 FILLER_32_1435 ();
 sg13g2_decap_8 FILLER_32_1442 ();
 sg13g2_decap_8 FILLER_32_1449 ();
 sg13g2_decap_8 FILLER_32_1456 ();
 sg13g2_decap_8 FILLER_32_1463 ();
 sg13g2_decap_8 FILLER_32_1470 ();
 sg13g2_decap_8 FILLER_32_1477 ();
 sg13g2_decap_8 FILLER_32_1484 ();
 sg13g2_decap_8 FILLER_32_1491 ();
 sg13g2_decap_8 FILLER_32_1498 ();
 sg13g2_decap_8 FILLER_32_1505 ();
 sg13g2_decap_8 FILLER_32_1512 ();
 sg13g2_decap_8 FILLER_32_1519 ();
 sg13g2_decap_8 FILLER_32_1526 ();
 sg13g2_decap_8 FILLER_32_1533 ();
 sg13g2_decap_8 FILLER_32_1540 ();
 sg13g2_decap_8 FILLER_32_1547 ();
 sg13g2_decap_8 FILLER_32_1554 ();
 sg13g2_decap_8 FILLER_32_1561 ();
 sg13g2_decap_8 FILLER_32_1568 ();
 sg13g2_decap_8 FILLER_32_1575 ();
 sg13g2_decap_8 FILLER_32_1582 ();
 sg13g2_decap_8 FILLER_32_1589 ();
 sg13g2_decap_8 FILLER_32_1596 ();
 sg13g2_decap_8 FILLER_32_1603 ();
 sg13g2_decap_8 FILLER_32_1610 ();
 sg13g2_decap_8 FILLER_32_1617 ();
 sg13g2_decap_8 FILLER_32_1624 ();
 sg13g2_decap_8 FILLER_32_1631 ();
 sg13g2_decap_8 FILLER_32_1638 ();
 sg13g2_decap_8 FILLER_32_1645 ();
 sg13g2_decap_8 FILLER_32_1652 ();
 sg13g2_decap_8 FILLER_32_1659 ();
 sg13g2_decap_8 FILLER_32_1666 ();
 sg13g2_decap_8 FILLER_32_1673 ();
 sg13g2_decap_8 FILLER_32_1680 ();
 sg13g2_decap_8 FILLER_32_1687 ();
 sg13g2_decap_8 FILLER_32_1694 ();
 sg13g2_decap_8 FILLER_32_1701 ();
 sg13g2_decap_8 FILLER_32_1708 ();
 sg13g2_decap_8 FILLER_32_1715 ();
 sg13g2_decap_8 FILLER_32_1722 ();
 sg13g2_decap_8 FILLER_32_1729 ();
 sg13g2_decap_8 FILLER_32_1736 ();
 sg13g2_decap_8 FILLER_32_1743 ();
 sg13g2_decap_8 FILLER_32_1750 ();
 sg13g2_decap_8 FILLER_32_1757 ();
 sg13g2_decap_8 FILLER_32_1764 ();
 sg13g2_decap_8 FILLER_32_1771 ();
 sg13g2_decap_8 FILLER_32_1778 ();
 sg13g2_decap_8 FILLER_32_1785 ();
 sg13g2_decap_8 FILLER_32_1792 ();
 sg13g2_decap_8 FILLER_32_1799 ();
 sg13g2_decap_8 FILLER_32_1806 ();
 sg13g2_decap_8 FILLER_32_1813 ();
 sg13g2_decap_8 FILLER_32_1820 ();
 sg13g2_decap_8 FILLER_32_1827 ();
 sg13g2_decap_8 FILLER_32_1834 ();
 sg13g2_decap_8 FILLER_32_1841 ();
 sg13g2_decap_8 FILLER_32_1848 ();
 sg13g2_decap_8 FILLER_32_1855 ();
 sg13g2_decap_8 FILLER_32_1862 ();
 sg13g2_decap_8 FILLER_32_1869 ();
 sg13g2_decap_8 FILLER_32_1876 ();
 sg13g2_decap_8 FILLER_32_1883 ();
 sg13g2_decap_8 FILLER_32_1890 ();
 sg13g2_decap_8 FILLER_32_1897 ();
 sg13g2_decap_8 FILLER_32_1904 ();
 sg13g2_decap_8 FILLER_32_1911 ();
 sg13g2_decap_8 FILLER_32_1918 ();
 sg13g2_decap_8 FILLER_32_1925 ();
 sg13g2_decap_8 FILLER_32_1932 ();
 sg13g2_decap_8 FILLER_32_1939 ();
 sg13g2_decap_8 FILLER_32_1946 ();
 sg13g2_decap_8 FILLER_32_1953 ();
 sg13g2_decap_8 FILLER_32_1960 ();
 sg13g2_decap_8 FILLER_32_1967 ();
 sg13g2_decap_8 FILLER_32_1974 ();
 sg13g2_decap_8 FILLER_32_1981 ();
 sg13g2_decap_8 FILLER_32_1988 ();
 sg13g2_decap_8 FILLER_32_1995 ();
 sg13g2_decap_8 FILLER_32_2002 ();
 sg13g2_decap_8 FILLER_32_2009 ();
 sg13g2_decap_8 FILLER_32_2016 ();
 sg13g2_decap_8 FILLER_32_2023 ();
 sg13g2_decap_8 FILLER_32_2030 ();
 sg13g2_decap_8 FILLER_32_2037 ();
 sg13g2_decap_8 FILLER_32_2044 ();
 sg13g2_decap_8 FILLER_32_2051 ();
 sg13g2_decap_8 FILLER_32_2058 ();
 sg13g2_decap_8 FILLER_32_2065 ();
 sg13g2_decap_8 FILLER_32_2072 ();
 sg13g2_decap_8 FILLER_32_2079 ();
 sg13g2_decap_8 FILLER_32_2086 ();
 sg13g2_decap_8 FILLER_32_2093 ();
 sg13g2_decap_8 FILLER_32_2100 ();
 sg13g2_decap_8 FILLER_32_2107 ();
 sg13g2_decap_8 FILLER_32_2114 ();
 sg13g2_decap_8 FILLER_32_2121 ();
 sg13g2_decap_8 FILLER_32_2128 ();
 sg13g2_decap_8 FILLER_32_2135 ();
 sg13g2_decap_8 FILLER_32_2142 ();
 sg13g2_decap_8 FILLER_32_2149 ();
 sg13g2_decap_8 FILLER_32_2156 ();
 sg13g2_decap_8 FILLER_32_2163 ();
 sg13g2_decap_8 FILLER_32_2170 ();
 sg13g2_decap_8 FILLER_32_2177 ();
 sg13g2_decap_8 FILLER_32_2184 ();
 sg13g2_decap_8 FILLER_32_2191 ();
 sg13g2_decap_8 FILLER_32_2198 ();
 sg13g2_decap_8 FILLER_32_2205 ();
 sg13g2_decap_8 FILLER_32_2212 ();
 sg13g2_decap_8 FILLER_32_2219 ();
 sg13g2_decap_8 FILLER_32_2226 ();
 sg13g2_decap_8 FILLER_32_2233 ();
 sg13g2_decap_8 FILLER_32_2240 ();
 sg13g2_decap_8 FILLER_32_2247 ();
 sg13g2_decap_8 FILLER_32_2254 ();
 sg13g2_decap_8 FILLER_32_2261 ();
 sg13g2_decap_8 FILLER_32_2268 ();
 sg13g2_decap_8 FILLER_32_2275 ();
 sg13g2_decap_8 FILLER_32_2282 ();
 sg13g2_decap_8 FILLER_32_2289 ();
 sg13g2_decap_8 FILLER_32_2296 ();
 sg13g2_decap_8 FILLER_32_2303 ();
 sg13g2_decap_8 FILLER_32_2310 ();
 sg13g2_decap_8 FILLER_32_2317 ();
 sg13g2_decap_8 FILLER_32_2324 ();
 sg13g2_decap_8 FILLER_32_2331 ();
 sg13g2_decap_8 FILLER_32_2338 ();
 sg13g2_decap_8 FILLER_32_2345 ();
 sg13g2_decap_8 FILLER_32_2352 ();
 sg13g2_decap_8 FILLER_32_2359 ();
 sg13g2_decap_8 FILLER_32_2366 ();
 sg13g2_decap_8 FILLER_32_2373 ();
 sg13g2_decap_8 FILLER_32_2380 ();
 sg13g2_decap_8 FILLER_32_2387 ();
 sg13g2_decap_8 FILLER_32_2394 ();
 sg13g2_decap_8 FILLER_32_2401 ();
 sg13g2_decap_8 FILLER_32_2408 ();
 sg13g2_decap_8 FILLER_32_2415 ();
 sg13g2_decap_8 FILLER_32_2422 ();
 sg13g2_decap_8 FILLER_32_2429 ();
 sg13g2_decap_8 FILLER_32_2436 ();
 sg13g2_decap_8 FILLER_32_2443 ();
 sg13g2_decap_8 FILLER_32_2450 ();
 sg13g2_decap_8 FILLER_32_2457 ();
 sg13g2_decap_8 FILLER_32_2464 ();
 sg13g2_decap_8 FILLER_32_2471 ();
 sg13g2_decap_8 FILLER_32_2478 ();
 sg13g2_decap_8 FILLER_32_2485 ();
 sg13g2_decap_8 FILLER_32_2492 ();
 sg13g2_decap_8 FILLER_32_2499 ();
 sg13g2_decap_8 FILLER_32_2506 ();
 sg13g2_decap_8 FILLER_32_2513 ();
 sg13g2_decap_8 FILLER_32_2520 ();
 sg13g2_decap_8 FILLER_32_2527 ();
 sg13g2_decap_8 FILLER_32_2534 ();
 sg13g2_decap_8 FILLER_32_2541 ();
 sg13g2_decap_8 FILLER_32_2548 ();
 sg13g2_decap_8 FILLER_32_2555 ();
 sg13g2_decap_8 FILLER_32_2562 ();
 sg13g2_decap_8 FILLER_32_2569 ();
 sg13g2_decap_8 FILLER_32_2576 ();
 sg13g2_decap_8 FILLER_32_2583 ();
 sg13g2_decap_8 FILLER_32_2590 ();
 sg13g2_decap_8 FILLER_32_2597 ();
 sg13g2_decap_8 FILLER_32_2604 ();
 sg13g2_decap_8 FILLER_32_2611 ();
 sg13g2_decap_8 FILLER_32_2618 ();
 sg13g2_decap_8 FILLER_32_2625 ();
 sg13g2_decap_8 FILLER_32_2632 ();
 sg13g2_decap_8 FILLER_32_2639 ();
 sg13g2_decap_8 FILLER_32_2646 ();
 sg13g2_decap_8 FILLER_32_2653 ();
 sg13g2_decap_8 FILLER_32_2660 ();
 sg13g2_decap_8 FILLER_32_2667 ();
 sg13g2_decap_8 FILLER_32_2674 ();
 sg13g2_decap_8 FILLER_32_2681 ();
 sg13g2_decap_8 FILLER_32_2688 ();
 sg13g2_decap_8 FILLER_32_2695 ();
 sg13g2_decap_8 FILLER_32_2702 ();
 sg13g2_decap_8 FILLER_32_2709 ();
 sg13g2_decap_8 FILLER_32_2716 ();
 sg13g2_decap_8 FILLER_32_2723 ();
 sg13g2_decap_8 FILLER_32_2730 ();
 sg13g2_decap_8 FILLER_32_2737 ();
 sg13g2_decap_8 FILLER_32_2744 ();
 sg13g2_decap_8 FILLER_32_2751 ();
 sg13g2_decap_8 FILLER_32_2758 ();
 sg13g2_decap_8 FILLER_32_2765 ();
 sg13g2_decap_8 FILLER_32_2772 ();
 sg13g2_decap_8 FILLER_32_2779 ();
 sg13g2_decap_8 FILLER_32_2786 ();
 sg13g2_decap_8 FILLER_32_2793 ();
 sg13g2_decap_8 FILLER_32_2800 ();
 sg13g2_decap_8 FILLER_32_2807 ();
 sg13g2_decap_8 FILLER_32_2814 ();
 sg13g2_decap_8 FILLER_32_2821 ();
 sg13g2_decap_8 FILLER_32_2828 ();
 sg13g2_decap_8 FILLER_32_2835 ();
 sg13g2_decap_8 FILLER_32_2842 ();
 sg13g2_decap_8 FILLER_32_2849 ();
 sg13g2_decap_8 FILLER_32_2856 ();
 sg13g2_decap_8 FILLER_32_2863 ();
 sg13g2_decap_8 FILLER_32_2870 ();
 sg13g2_decap_8 FILLER_32_2877 ();
 sg13g2_decap_8 FILLER_32_2884 ();
 sg13g2_decap_8 FILLER_32_2891 ();
 sg13g2_decap_8 FILLER_32_2898 ();
 sg13g2_decap_8 FILLER_32_2905 ();
 sg13g2_decap_8 FILLER_32_2912 ();
 sg13g2_decap_8 FILLER_32_2919 ();
 sg13g2_decap_8 FILLER_32_2926 ();
 sg13g2_decap_8 FILLER_32_2933 ();
 sg13g2_decap_8 FILLER_32_2940 ();
 sg13g2_decap_8 FILLER_32_2947 ();
 sg13g2_decap_8 FILLER_32_2954 ();
 sg13g2_decap_8 FILLER_32_2961 ();
 sg13g2_decap_8 FILLER_32_2968 ();
 sg13g2_decap_8 FILLER_32_2975 ();
 sg13g2_decap_8 FILLER_32_2982 ();
 sg13g2_decap_8 FILLER_32_2989 ();
 sg13g2_decap_8 FILLER_32_2996 ();
 sg13g2_decap_8 FILLER_32_3003 ();
 sg13g2_decap_8 FILLER_32_3010 ();
 sg13g2_decap_8 FILLER_32_3017 ();
 sg13g2_decap_8 FILLER_32_3024 ();
 sg13g2_decap_8 FILLER_32_3031 ();
 sg13g2_decap_8 FILLER_32_3038 ();
 sg13g2_decap_8 FILLER_32_3045 ();
 sg13g2_decap_8 FILLER_32_3052 ();
 sg13g2_decap_8 FILLER_32_3059 ();
 sg13g2_decap_8 FILLER_32_3066 ();
 sg13g2_decap_8 FILLER_32_3073 ();
 sg13g2_decap_8 FILLER_32_3080 ();
 sg13g2_decap_8 FILLER_32_3087 ();
 sg13g2_decap_8 FILLER_32_3094 ();
 sg13g2_decap_8 FILLER_32_3101 ();
 sg13g2_decap_8 FILLER_32_3108 ();
 sg13g2_decap_8 FILLER_32_3115 ();
 sg13g2_decap_8 FILLER_32_3122 ();
 sg13g2_decap_8 FILLER_32_3129 ();
 sg13g2_decap_8 FILLER_32_3136 ();
 sg13g2_decap_8 FILLER_32_3143 ();
 sg13g2_decap_8 FILLER_32_3150 ();
 sg13g2_decap_8 FILLER_32_3157 ();
 sg13g2_decap_8 FILLER_32_3164 ();
 sg13g2_decap_8 FILLER_32_3171 ();
 sg13g2_decap_8 FILLER_32_3178 ();
 sg13g2_decap_8 FILLER_32_3185 ();
 sg13g2_decap_8 FILLER_32_3192 ();
 sg13g2_decap_8 FILLER_32_3199 ();
 sg13g2_decap_8 FILLER_32_3206 ();
 sg13g2_decap_8 FILLER_32_3213 ();
 sg13g2_decap_8 FILLER_32_3220 ();
 sg13g2_decap_8 FILLER_32_3227 ();
 sg13g2_decap_8 FILLER_32_3234 ();
 sg13g2_decap_8 FILLER_32_3241 ();
 sg13g2_decap_8 FILLER_32_3248 ();
 sg13g2_decap_8 FILLER_32_3255 ();
 sg13g2_decap_8 FILLER_32_3262 ();
 sg13g2_decap_8 FILLER_32_3269 ();
 sg13g2_decap_8 FILLER_32_3276 ();
 sg13g2_decap_8 FILLER_32_3283 ();
 sg13g2_decap_8 FILLER_32_3290 ();
 sg13g2_decap_8 FILLER_32_3297 ();
 sg13g2_decap_8 FILLER_32_3304 ();
 sg13g2_decap_8 FILLER_32_3311 ();
 sg13g2_decap_8 FILLER_32_3318 ();
 sg13g2_decap_8 FILLER_32_3325 ();
 sg13g2_decap_8 FILLER_32_3332 ();
 sg13g2_decap_8 FILLER_32_3339 ();
 sg13g2_decap_8 FILLER_32_3346 ();
 sg13g2_decap_8 FILLER_32_3353 ();
 sg13g2_decap_8 FILLER_32_3360 ();
 sg13g2_decap_8 FILLER_32_3367 ();
 sg13g2_decap_8 FILLER_32_3374 ();
 sg13g2_decap_8 FILLER_32_3381 ();
 sg13g2_decap_8 FILLER_32_3388 ();
 sg13g2_decap_8 FILLER_32_3395 ();
 sg13g2_decap_8 FILLER_32_3402 ();
 sg13g2_decap_8 FILLER_32_3409 ();
 sg13g2_decap_8 FILLER_32_3416 ();
 sg13g2_decap_8 FILLER_32_3423 ();
 sg13g2_decap_8 FILLER_32_3430 ();
 sg13g2_decap_8 FILLER_32_3437 ();
 sg13g2_decap_8 FILLER_32_3444 ();
 sg13g2_decap_8 FILLER_32_3451 ();
 sg13g2_decap_8 FILLER_32_3458 ();
 sg13g2_decap_8 FILLER_32_3465 ();
 sg13g2_decap_8 FILLER_32_3472 ();
 sg13g2_decap_8 FILLER_32_3479 ();
 sg13g2_decap_8 FILLER_32_3486 ();
 sg13g2_decap_8 FILLER_32_3493 ();
 sg13g2_decap_8 FILLER_32_3500 ();
 sg13g2_decap_8 FILLER_32_3507 ();
 sg13g2_decap_8 FILLER_32_3514 ();
 sg13g2_decap_8 FILLER_32_3521 ();
 sg13g2_decap_8 FILLER_32_3528 ();
 sg13g2_decap_8 FILLER_32_3535 ();
 sg13g2_decap_8 FILLER_32_3542 ();
 sg13g2_decap_8 FILLER_32_3549 ();
 sg13g2_decap_8 FILLER_32_3556 ();
 sg13g2_decap_8 FILLER_32_3563 ();
 sg13g2_decap_8 FILLER_32_3570 ();
 sg13g2_fill_2 FILLER_32_3577 ();
 sg13g2_fill_1 FILLER_32_3579 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_259 ();
 sg13g2_decap_8 FILLER_33_266 ();
 sg13g2_decap_8 FILLER_33_273 ();
 sg13g2_decap_8 FILLER_33_280 ();
 sg13g2_decap_8 FILLER_33_287 ();
 sg13g2_decap_8 FILLER_33_294 ();
 sg13g2_decap_8 FILLER_33_301 ();
 sg13g2_decap_8 FILLER_33_308 ();
 sg13g2_decap_8 FILLER_33_315 ();
 sg13g2_decap_8 FILLER_33_322 ();
 sg13g2_decap_8 FILLER_33_329 ();
 sg13g2_decap_8 FILLER_33_336 ();
 sg13g2_decap_8 FILLER_33_343 ();
 sg13g2_decap_8 FILLER_33_350 ();
 sg13g2_decap_8 FILLER_33_357 ();
 sg13g2_decap_8 FILLER_33_364 ();
 sg13g2_decap_8 FILLER_33_371 ();
 sg13g2_decap_8 FILLER_33_378 ();
 sg13g2_decap_8 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_399 ();
 sg13g2_decap_8 FILLER_33_406 ();
 sg13g2_decap_8 FILLER_33_413 ();
 sg13g2_decap_8 FILLER_33_420 ();
 sg13g2_decap_8 FILLER_33_427 ();
 sg13g2_decap_8 FILLER_33_434 ();
 sg13g2_decap_8 FILLER_33_441 ();
 sg13g2_decap_8 FILLER_33_448 ();
 sg13g2_decap_8 FILLER_33_455 ();
 sg13g2_decap_8 FILLER_33_462 ();
 sg13g2_decap_8 FILLER_33_469 ();
 sg13g2_decap_8 FILLER_33_476 ();
 sg13g2_decap_8 FILLER_33_483 ();
 sg13g2_decap_8 FILLER_33_490 ();
 sg13g2_decap_8 FILLER_33_497 ();
 sg13g2_decap_8 FILLER_33_504 ();
 sg13g2_decap_8 FILLER_33_511 ();
 sg13g2_decap_8 FILLER_33_518 ();
 sg13g2_decap_8 FILLER_33_525 ();
 sg13g2_decap_8 FILLER_33_532 ();
 sg13g2_decap_8 FILLER_33_539 ();
 sg13g2_decap_8 FILLER_33_546 ();
 sg13g2_decap_8 FILLER_33_553 ();
 sg13g2_decap_8 FILLER_33_560 ();
 sg13g2_decap_8 FILLER_33_567 ();
 sg13g2_decap_8 FILLER_33_574 ();
 sg13g2_decap_8 FILLER_33_581 ();
 sg13g2_decap_8 FILLER_33_588 ();
 sg13g2_decap_8 FILLER_33_595 ();
 sg13g2_decap_8 FILLER_33_602 ();
 sg13g2_decap_8 FILLER_33_609 ();
 sg13g2_decap_8 FILLER_33_616 ();
 sg13g2_decap_8 FILLER_33_623 ();
 sg13g2_decap_8 FILLER_33_630 ();
 sg13g2_decap_8 FILLER_33_637 ();
 sg13g2_decap_8 FILLER_33_644 ();
 sg13g2_decap_8 FILLER_33_651 ();
 sg13g2_decap_8 FILLER_33_658 ();
 sg13g2_decap_8 FILLER_33_665 ();
 sg13g2_decap_8 FILLER_33_672 ();
 sg13g2_decap_8 FILLER_33_679 ();
 sg13g2_decap_8 FILLER_33_686 ();
 sg13g2_decap_8 FILLER_33_693 ();
 sg13g2_decap_8 FILLER_33_700 ();
 sg13g2_decap_8 FILLER_33_707 ();
 sg13g2_decap_8 FILLER_33_714 ();
 sg13g2_decap_8 FILLER_33_721 ();
 sg13g2_decap_8 FILLER_33_728 ();
 sg13g2_decap_8 FILLER_33_735 ();
 sg13g2_decap_8 FILLER_33_742 ();
 sg13g2_decap_8 FILLER_33_749 ();
 sg13g2_decap_8 FILLER_33_756 ();
 sg13g2_decap_8 FILLER_33_763 ();
 sg13g2_decap_8 FILLER_33_770 ();
 sg13g2_decap_8 FILLER_33_777 ();
 sg13g2_decap_8 FILLER_33_784 ();
 sg13g2_decap_8 FILLER_33_791 ();
 sg13g2_decap_8 FILLER_33_798 ();
 sg13g2_decap_8 FILLER_33_805 ();
 sg13g2_decap_8 FILLER_33_812 ();
 sg13g2_decap_8 FILLER_33_819 ();
 sg13g2_decap_8 FILLER_33_826 ();
 sg13g2_decap_8 FILLER_33_833 ();
 sg13g2_decap_8 FILLER_33_840 ();
 sg13g2_decap_8 FILLER_33_847 ();
 sg13g2_decap_8 FILLER_33_854 ();
 sg13g2_decap_8 FILLER_33_861 ();
 sg13g2_decap_8 FILLER_33_868 ();
 sg13g2_decap_8 FILLER_33_875 ();
 sg13g2_decap_8 FILLER_33_882 ();
 sg13g2_decap_8 FILLER_33_889 ();
 sg13g2_decap_8 FILLER_33_896 ();
 sg13g2_decap_8 FILLER_33_903 ();
 sg13g2_decap_8 FILLER_33_910 ();
 sg13g2_decap_8 FILLER_33_917 ();
 sg13g2_decap_8 FILLER_33_924 ();
 sg13g2_decap_8 FILLER_33_931 ();
 sg13g2_decap_8 FILLER_33_938 ();
 sg13g2_decap_8 FILLER_33_945 ();
 sg13g2_decap_8 FILLER_33_952 ();
 sg13g2_decap_8 FILLER_33_959 ();
 sg13g2_decap_8 FILLER_33_966 ();
 sg13g2_decap_8 FILLER_33_973 ();
 sg13g2_decap_8 FILLER_33_980 ();
 sg13g2_decap_8 FILLER_33_987 ();
 sg13g2_decap_8 FILLER_33_994 ();
 sg13g2_decap_8 FILLER_33_1001 ();
 sg13g2_decap_8 FILLER_33_1008 ();
 sg13g2_decap_8 FILLER_33_1015 ();
 sg13g2_decap_8 FILLER_33_1022 ();
 sg13g2_decap_8 FILLER_33_1029 ();
 sg13g2_decap_8 FILLER_33_1036 ();
 sg13g2_decap_8 FILLER_33_1043 ();
 sg13g2_decap_8 FILLER_33_1050 ();
 sg13g2_decap_8 FILLER_33_1057 ();
 sg13g2_decap_8 FILLER_33_1064 ();
 sg13g2_decap_8 FILLER_33_1071 ();
 sg13g2_decap_8 FILLER_33_1078 ();
 sg13g2_decap_8 FILLER_33_1085 ();
 sg13g2_decap_8 FILLER_33_1092 ();
 sg13g2_decap_8 FILLER_33_1099 ();
 sg13g2_decap_8 FILLER_33_1106 ();
 sg13g2_decap_8 FILLER_33_1113 ();
 sg13g2_decap_8 FILLER_33_1120 ();
 sg13g2_decap_8 FILLER_33_1127 ();
 sg13g2_decap_8 FILLER_33_1134 ();
 sg13g2_decap_8 FILLER_33_1141 ();
 sg13g2_decap_8 FILLER_33_1148 ();
 sg13g2_decap_8 FILLER_33_1155 ();
 sg13g2_decap_8 FILLER_33_1162 ();
 sg13g2_decap_8 FILLER_33_1169 ();
 sg13g2_decap_8 FILLER_33_1176 ();
 sg13g2_decap_8 FILLER_33_1183 ();
 sg13g2_decap_8 FILLER_33_1190 ();
 sg13g2_decap_8 FILLER_33_1197 ();
 sg13g2_decap_8 FILLER_33_1204 ();
 sg13g2_decap_8 FILLER_33_1211 ();
 sg13g2_decap_8 FILLER_33_1218 ();
 sg13g2_decap_8 FILLER_33_1225 ();
 sg13g2_decap_8 FILLER_33_1232 ();
 sg13g2_decap_8 FILLER_33_1239 ();
 sg13g2_decap_8 FILLER_33_1246 ();
 sg13g2_decap_8 FILLER_33_1253 ();
 sg13g2_decap_8 FILLER_33_1260 ();
 sg13g2_decap_8 FILLER_33_1267 ();
 sg13g2_decap_8 FILLER_33_1274 ();
 sg13g2_decap_8 FILLER_33_1281 ();
 sg13g2_decap_8 FILLER_33_1288 ();
 sg13g2_decap_8 FILLER_33_1295 ();
 sg13g2_decap_8 FILLER_33_1302 ();
 sg13g2_decap_8 FILLER_33_1309 ();
 sg13g2_decap_8 FILLER_33_1316 ();
 sg13g2_decap_8 FILLER_33_1323 ();
 sg13g2_decap_8 FILLER_33_1330 ();
 sg13g2_decap_8 FILLER_33_1337 ();
 sg13g2_decap_8 FILLER_33_1344 ();
 sg13g2_decap_8 FILLER_33_1351 ();
 sg13g2_decap_8 FILLER_33_1358 ();
 sg13g2_decap_8 FILLER_33_1365 ();
 sg13g2_decap_8 FILLER_33_1372 ();
 sg13g2_decap_8 FILLER_33_1379 ();
 sg13g2_decap_8 FILLER_33_1386 ();
 sg13g2_decap_8 FILLER_33_1393 ();
 sg13g2_decap_8 FILLER_33_1400 ();
 sg13g2_decap_8 FILLER_33_1407 ();
 sg13g2_decap_8 FILLER_33_1414 ();
 sg13g2_decap_8 FILLER_33_1421 ();
 sg13g2_decap_8 FILLER_33_1428 ();
 sg13g2_decap_8 FILLER_33_1435 ();
 sg13g2_decap_8 FILLER_33_1442 ();
 sg13g2_decap_8 FILLER_33_1449 ();
 sg13g2_decap_8 FILLER_33_1456 ();
 sg13g2_decap_8 FILLER_33_1463 ();
 sg13g2_decap_8 FILLER_33_1470 ();
 sg13g2_decap_8 FILLER_33_1477 ();
 sg13g2_decap_8 FILLER_33_1484 ();
 sg13g2_decap_8 FILLER_33_1491 ();
 sg13g2_decap_8 FILLER_33_1498 ();
 sg13g2_decap_8 FILLER_33_1505 ();
 sg13g2_decap_8 FILLER_33_1512 ();
 sg13g2_decap_8 FILLER_33_1519 ();
 sg13g2_decap_8 FILLER_33_1526 ();
 sg13g2_decap_8 FILLER_33_1533 ();
 sg13g2_decap_8 FILLER_33_1540 ();
 sg13g2_decap_8 FILLER_33_1547 ();
 sg13g2_decap_8 FILLER_33_1554 ();
 sg13g2_decap_8 FILLER_33_1561 ();
 sg13g2_decap_8 FILLER_33_1568 ();
 sg13g2_decap_8 FILLER_33_1575 ();
 sg13g2_decap_8 FILLER_33_1582 ();
 sg13g2_decap_8 FILLER_33_1589 ();
 sg13g2_decap_8 FILLER_33_1596 ();
 sg13g2_decap_8 FILLER_33_1603 ();
 sg13g2_decap_8 FILLER_33_1610 ();
 sg13g2_decap_8 FILLER_33_1617 ();
 sg13g2_decap_8 FILLER_33_1624 ();
 sg13g2_decap_8 FILLER_33_1631 ();
 sg13g2_decap_8 FILLER_33_1638 ();
 sg13g2_decap_8 FILLER_33_1645 ();
 sg13g2_decap_8 FILLER_33_1652 ();
 sg13g2_decap_8 FILLER_33_1659 ();
 sg13g2_decap_8 FILLER_33_1666 ();
 sg13g2_decap_8 FILLER_33_1673 ();
 sg13g2_decap_8 FILLER_33_1680 ();
 sg13g2_decap_8 FILLER_33_1687 ();
 sg13g2_decap_8 FILLER_33_1694 ();
 sg13g2_decap_8 FILLER_33_1701 ();
 sg13g2_decap_8 FILLER_33_1708 ();
 sg13g2_decap_8 FILLER_33_1715 ();
 sg13g2_decap_8 FILLER_33_1722 ();
 sg13g2_decap_8 FILLER_33_1729 ();
 sg13g2_decap_8 FILLER_33_1736 ();
 sg13g2_decap_8 FILLER_33_1743 ();
 sg13g2_decap_8 FILLER_33_1750 ();
 sg13g2_decap_8 FILLER_33_1757 ();
 sg13g2_decap_8 FILLER_33_1764 ();
 sg13g2_decap_8 FILLER_33_1771 ();
 sg13g2_decap_8 FILLER_33_1778 ();
 sg13g2_decap_8 FILLER_33_1785 ();
 sg13g2_decap_8 FILLER_33_1792 ();
 sg13g2_decap_8 FILLER_33_1799 ();
 sg13g2_decap_8 FILLER_33_1806 ();
 sg13g2_decap_8 FILLER_33_1813 ();
 sg13g2_decap_8 FILLER_33_1820 ();
 sg13g2_decap_8 FILLER_33_1827 ();
 sg13g2_decap_8 FILLER_33_1834 ();
 sg13g2_decap_8 FILLER_33_1841 ();
 sg13g2_decap_8 FILLER_33_1848 ();
 sg13g2_decap_8 FILLER_33_1855 ();
 sg13g2_decap_8 FILLER_33_1862 ();
 sg13g2_decap_8 FILLER_33_1869 ();
 sg13g2_decap_8 FILLER_33_1876 ();
 sg13g2_decap_8 FILLER_33_1883 ();
 sg13g2_decap_8 FILLER_33_1890 ();
 sg13g2_decap_8 FILLER_33_1897 ();
 sg13g2_decap_8 FILLER_33_1904 ();
 sg13g2_decap_8 FILLER_33_1911 ();
 sg13g2_decap_8 FILLER_33_1918 ();
 sg13g2_decap_8 FILLER_33_1925 ();
 sg13g2_decap_8 FILLER_33_1932 ();
 sg13g2_decap_8 FILLER_33_1939 ();
 sg13g2_decap_8 FILLER_33_1946 ();
 sg13g2_decap_8 FILLER_33_1953 ();
 sg13g2_decap_8 FILLER_33_1960 ();
 sg13g2_decap_8 FILLER_33_1967 ();
 sg13g2_decap_8 FILLER_33_1974 ();
 sg13g2_decap_8 FILLER_33_1981 ();
 sg13g2_decap_8 FILLER_33_1988 ();
 sg13g2_decap_8 FILLER_33_1995 ();
 sg13g2_decap_8 FILLER_33_2002 ();
 sg13g2_decap_8 FILLER_33_2009 ();
 sg13g2_decap_8 FILLER_33_2016 ();
 sg13g2_decap_8 FILLER_33_2023 ();
 sg13g2_decap_8 FILLER_33_2030 ();
 sg13g2_decap_8 FILLER_33_2037 ();
 sg13g2_decap_8 FILLER_33_2044 ();
 sg13g2_decap_8 FILLER_33_2051 ();
 sg13g2_decap_8 FILLER_33_2058 ();
 sg13g2_decap_8 FILLER_33_2065 ();
 sg13g2_decap_8 FILLER_33_2072 ();
 sg13g2_decap_8 FILLER_33_2079 ();
 sg13g2_decap_8 FILLER_33_2086 ();
 sg13g2_decap_8 FILLER_33_2093 ();
 sg13g2_decap_8 FILLER_33_2100 ();
 sg13g2_decap_8 FILLER_33_2107 ();
 sg13g2_decap_8 FILLER_33_2114 ();
 sg13g2_decap_8 FILLER_33_2121 ();
 sg13g2_decap_8 FILLER_33_2128 ();
 sg13g2_decap_8 FILLER_33_2135 ();
 sg13g2_decap_8 FILLER_33_2142 ();
 sg13g2_decap_8 FILLER_33_2149 ();
 sg13g2_decap_8 FILLER_33_2156 ();
 sg13g2_decap_8 FILLER_33_2163 ();
 sg13g2_decap_8 FILLER_33_2170 ();
 sg13g2_decap_8 FILLER_33_2177 ();
 sg13g2_decap_8 FILLER_33_2184 ();
 sg13g2_decap_8 FILLER_33_2191 ();
 sg13g2_decap_8 FILLER_33_2198 ();
 sg13g2_decap_8 FILLER_33_2205 ();
 sg13g2_decap_8 FILLER_33_2212 ();
 sg13g2_decap_8 FILLER_33_2219 ();
 sg13g2_decap_8 FILLER_33_2226 ();
 sg13g2_decap_8 FILLER_33_2233 ();
 sg13g2_decap_8 FILLER_33_2240 ();
 sg13g2_decap_8 FILLER_33_2247 ();
 sg13g2_decap_8 FILLER_33_2254 ();
 sg13g2_decap_8 FILLER_33_2261 ();
 sg13g2_decap_8 FILLER_33_2268 ();
 sg13g2_decap_8 FILLER_33_2275 ();
 sg13g2_decap_8 FILLER_33_2282 ();
 sg13g2_decap_8 FILLER_33_2289 ();
 sg13g2_decap_8 FILLER_33_2296 ();
 sg13g2_decap_8 FILLER_33_2303 ();
 sg13g2_decap_8 FILLER_33_2310 ();
 sg13g2_decap_8 FILLER_33_2317 ();
 sg13g2_decap_8 FILLER_33_2324 ();
 sg13g2_decap_8 FILLER_33_2331 ();
 sg13g2_decap_8 FILLER_33_2338 ();
 sg13g2_decap_8 FILLER_33_2345 ();
 sg13g2_decap_8 FILLER_33_2352 ();
 sg13g2_decap_8 FILLER_33_2359 ();
 sg13g2_decap_8 FILLER_33_2366 ();
 sg13g2_decap_8 FILLER_33_2373 ();
 sg13g2_decap_8 FILLER_33_2380 ();
 sg13g2_decap_8 FILLER_33_2387 ();
 sg13g2_decap_8 FILLER_33_2394 ();
 sg13g2_decap_8 FILLER_33_2401 ();
 sg13g2_decap_8 FILLER_33_2408 ();
 sg13g2_decap_8 FILLER_33_2415 ();
 sg13g2_decap_8 FILLER_33_2422 ();
 sg13g2_decap_8 FILLER_33_2429 ();
 sg13g2_decap_8 FILLER_33_2436 ();
 sg13g2_decap_8 FILLER_33_2443 ();
 sg13g2_decap_8 FILLER_33_2450 ();
 sg13g2_decap_8 FILLER_33_2457 ();
 sg13g2_decap_8 FILLER_33_2464 ();
 sg13g2_decap_8 FILLER_33_2471 ();
 sg13g2_decap_8 FILLER_33_2478 ();
 sg13g2_decap_8 FILLER_33_2485 ();
 sg13g2_decap_8 FILLER_33_2492 ();
 sg13g2_decap_8 FILLER_33_2499 ();
 sg13g2_decap_8 FILLER_33_2506 ();
 sg13g2_decap_8 FILLER_33_2513 ();
 sg13g2_decap_8 FILLER_33_2520 ();
 sg13g2_decap_8 FILLER_33_2527 ();
 sg13g2_decap_8 FILLER_33_2534 ();
 sg13g2_decap_8 FILLER_33_2541 ();
 sg13g2_decap_8 FILLER_33_2548 ();
 sg13g2_decap_8 FILLER_33_2555 ();
 sg13g2_decap_8 FILLER_33_2562 ();
 sg13g2_decap_8 FILLER_33_2569 ();
 sg13g2_decap_8 FILLER_33_2576 ();
 sg13g2_decap_8 FILLER_33_2583 ();
 sg13g2_decap_8 FILLER_33_2590 ();
 sg13g2_decap_8 FILLER_33_2597 ();
 sg13g2_decap_8 FILLER_33_2604 ();
 sg13g2_decap_8 FILLER_33_2611 ();
 sg13g2_decap_8 FILLER_33_2618 ();
 sg13g2_decap_8 FILLER_33_2625 ();
 sg13g2_decap_8 FILLER_33_2632 ();
 sg13g2_decap_8 FILLER_33_2639 ();
 sg13g2_decap_8 FILLER_33_2646 ();
 sg13g2_decap_8 FILLER_33_2653 ();
 sg13g2_decap_8 FILLER_33_2660 ();
 sg13g2_decap_8 FILLER_33_2667 ();
 sg13g2_decap_8 FILLER_33_2674 ();
 sg13g2_decap_8 FILLER_33_2681 ();
 sg13g2_decap_8 FILLER_33_2688 ();
 sg13g2_decap_8 FILLER_33_2695 ();
 sg13g2_decap_8 FILLER_33_2702 ();
 sg13g2_decap_8 FILLER_33_2709 ();
 sg13g2_decap_8 FILLER_33_2716 ();
 sg13g2_decap_8 FILLER_33_2723 ();
 sg13g2_decap_8 FILLER_33_2730 ();
 sg13g2_decap_8 FILLER_33_2737 ();
 sg13g2_decap_8 FILLER_33_2744 ();
 sg13g2_decap_8 FILLER_33_2751 ();
 sg13g2_decap_8 FILLER_33_2758 ();
 sg13g2_decap_8 FILLER_33_2765 ();
 sg13g2_decap_8 FILLER_33_2772 ();
 sg13g2_decap_8 FILLER_33_2779 ();
 sg13g2_decap_8 FILLER_33_2786 ();
 sg13g2_decap_8 FILLER_33_2793 ();
 sg13g2_decap_8 FILLER_33_2800 ();
 sg13g2_decap_8 FILLER_33_2807 ();
 sg13g2_decap_8 FILLER_33_2814 ();
 sg13g2_decap_8 FILLER_33_2821 ();
 sg13g2_decap_8 FILLER_33_2828 ();
 sg13g2_decap_8 FILLER_33_2835 ();
 sg13g2_decap_8 FILLER_33_2842 ();
 sg13g2_decap_8 FILLER_33_2849 ();
 sg13g2_decap_8 FILLER_33_2856 ();
 sg13g2_decap_8 FILLER_33_2863 ();
 sg13g2_decap_8 FILLER_33_2870 ();
 sg13g2_decap_8 FILLER_33_2877 ();
 sg13g2_decap_8 FILLER_33_2884 ();
 sg13g2_decap_8 FILLER_33_2891 ();
 sg13g2_decap_8 FILLER_33_2898 ();
 sg13g2_decap_8 FILLER_33_2905 ();
 sg13g2_decap_8 FILLER_33_2912 ();
 sg13g2_decap_8 FILLER_33_2919 ();
 sg13g2_decap_8 FILLER_33_2926 ();
 sg13g2_decap_8 FILLER_33_2933 ();
 sg13g2_decap_8 FILLER_33_2940 ();
 sg13g2_decap_8 FILLER_33_2947 ();
 sg13g2_decap_8 FILLER_33_2954 ();
 sg13g2_decap_8 FILLER_33_2961 ();
 sg13g2_decap_8 FILLER_33_2968 ();
 sg13g2_decap_8 FILLER_33_2975 ();
 sg13g2_decap_8 FILLER_33_2982 ();
 sg13g2_decap_8 FILLER_33_2989 ();
 sg13g2_decap_8 FILLER_33_2996 ();
 sg13g2_decap_8 FILLER_33_3003 ();
 sg13g2_decap_8 FILLER_33_3010 ();
 sg13g2_decap_8 FILLER_33_3017 ();
 sg13g2_decap_8 FILLER_33_3024 ();
 sg13g2_decap_8 FILLER_33_3031 ();
 sg13g2_decap_8 FILLER_33_3038 ();
 sg13g2_decap_8 FILLER_33_3045 ();
 sg13g2_decap_8 FILLER_33_3052 ();
 sg13g2_decap_8 FILLER_33_3059 ();
 sg13g2_decap_8 FILLER_33_3066 ();
 sg13g2_decap_8 FILLER_33_3073 ();
 sg13g2_decap_8 FILLER_33_3080 ();
 sg13g2_decap_8 FILLER_33_3087 ();
 sg13g2_decap_8 FILLER_33_3094 ();
 sg13g2_decap_8 FILLER_33_3101 ();
 sg13g2_decap_8 FILLER_33_3108 ();
 sg13g2_decap_8 FILLER_33_3115 ();
 sg13g2_decap_8 FILLER_33_3122 ();
 sg13g2_decap_8 FILLER_33_3129 ();
 sg13g2_decap_8 FILLER_33_3136 ();
 sg13g2_decap_8 FILLER_33_3143 ();
 sg13g2_decap_8 FILLER_33_3150 ();
 sg13g2_decap_8 FILLER_33_3157 ();
 sg13g2_decap_8 FILLER_33_3164 ();
 sg13g2_decap_8 FILLER_33_3171 ();
 sg13g2_decap_8 FILLER_33_3178 ();
 sg13g2_decap_8 FILLER_33_3185 ();
 sg13g2_decap_8 FILLER_33_3192 ();
 sg13g2_decap_8 FILLER_33_3199 ();
 sg13g2_decap_8 FILLER_33_3206 ();
 sg13g2_decap_8 FILLER_33_3213 ();
 sg13g2_decap_8 FILLER_33_3220 ();
 sg13g2_decap_8 FILLER_33_3227 ();
 sg13g2_decap_8 FILLER_33_3234 ();
 sg13g2_decap_8 FILLER_33_3241 ();
 sg13g2_decap_8 FILLER_33_3248 ();
 sg13g2_decap_8 FILLER_33_3255 ();
 sg13g2_decap_8 FILLER_33_3262 ();
 sg13g2_decap_8 FILLER_33_3269 ();
 sg13g2_decap_8 FILLER_33_3276 ();
 sg13g2_decap_8 FILLER_33_3283 ();
 sg13g2_decap_8 FILLER_33_3290 ();
 sg13g2_decap_8 FILLER_33_3297 ();
 sg13g2_decap_8 FILLER_33_3304 ();
 sg13g2_decap_8 FILLER_33_3311 ();
 sg13g2_decap_8 FILLER_33_3318 ();
 sg13g2_decap_8 FILLER_33_3325 ();
 sg13g2_decap_8 FILLER_33_3332 ();
 sg13g2_decap_8 FILLER_33_3339 ();
 sg13g2_decap_8 FILLER_33_3346 ();
 sg13g2_decap_8 FILLER_33_3353 ();
 sg13g2_decap_8 FILLER_33_3360 ();
 sg13g2_decap_8 FILLER_33_3367 ();
 sg13g2_decap_8 FILLER_33_3374 ();
 sg13g2_decap_8 FILLER_33_3381 ();
 sg13g2_decap_8 FILLER_33_3388 ();
 sg13g2_decap_8 FILLER_33_3395 ();
 sg13g2_decap_8 FILLER_33_3402 ();
 sg13g2_decap_8 FILLER_33_3409 ();
 sg13g2_decap_8 FILLER_33_3416 ();
 sg13g2_decap_8 FILLER_33_3423 ();
 sg13g2_decap_8 FILLER_33_3430 ();
 sg13g2_decap_8 FILLER_33_3437 ();
 sg13g2_decap_8 FILLER_33_3444 ();
 sg13g2_decap_8 FILLER_33_3451 ();
 sg13g2_decap_8 FILLER_33_3458 ();
 sg13g2_decap_8 FILLER_33_3465 ();
 sg13g2_decap_8 FILLER_33_3472 ();
 sg13g2_decap_8 FILLER_33_3479 ();
 sg13g2_decap_8 FILLER_33_3486 ();
 sg13g2_decap_8 FILLER_33_3493 ();
 sg13g2_decap_8 FILLER_33_3500 ();
 sg13g2_decap_8 FILLER_33_3507 ();
 sg13g2_decap_8 FILLER_33_3514 ();
 sg13g2_decap_8 FILLER_33_3521 ();
 sg13g2_decap_8 FILLER_33_3528 ();
 sg13g2_decap_8 FILLER_33_3535 ();
 sg13g2_decap_8 FILLER_33_3542 ();
 sg13g2_decap_8 FILLER_33_3549 ();
 sg13g2_decap_8 FILLER_33_3556 ();
 sg13g2_decap_8 FILLER_33_3563 ();
 sg13g2_decap_8 FILLER_33_3570 ();
 sg13g2_fill_2 FILLER_33_3577 ();
 sg13g2_fill_1 FILLER_33_3579 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_280 ();
 sg13g2_decap_8 FILLER_34_287 ();
 sg13g2_decap_8 FILLER_34_294 ();
 sg13g2_decap_8 FILLER_34_301 ();
 sg13g2_decap_8 FILLER_34_308 ();
 sg13g2_decap_8 FILLER_34_315 ();
 sg13g2_decap_8 FILLER_34_322 ();
 sg13g2_decap_8 FILLER_34_329 ();
 sg13g2_decap_8 FILLER_34_336 ();
 sg13g2_decap_8 FILLER_34_343 ();
 sg13g2_decap_8 FILLER_34_350 ();
 sg13g2_decap_8 FILLER_34_357 ();
 sg13g2_decap_8 FILLER_34_364 ();
 sg13g2_decap_8 FILLER_34_371 ();
 sg13g2_decap_8 FILLER_34_378 ();
 sg13g2_decap_8 FILLER_34_385 ();
 sg13g2_decap_8 FILLER_34_392 ();
 sg13g2_decap_8 FILLER_34_399 ();
 sg13g2_decap_8 FILLER_34_406 ();
 sg13g2_decap_8 FILLER_34_413 ();
 sg13g2_decap_8 FILLER_34_420 ();
 sg13g2_decap_8 FILLER_34_427 ();
 sg13g2_decap_8 FILLER_34_434 ();
 sg13g2_decap_8 FILLER_34_441 ();
 sg13g2_decap_8 FILLER_34_448 ();
 sg13g2_decap_8 FILLER_34_455 ();
 sg13g2_decap_8 FILLER_34_462 ();
 sg13g2_decap_8 FILLER_34_469 ();
 sg13g2_decap_8 FILLER_34_476 ();
 sg13g2_decap_8 FILLER_34_483 ();
 sg13g2_decap_8 FILLER_34_490 ();
 sg13g2_decap_8 FILLER_34_497 ();
 sg13g2_decap_8 FILLER_34_504 ();
 sg13g2_decap_8 FILLER_34_511 ();
 sg13g2_decap_8 FILLER_34_518 ();
 sg13g2_decap_8 FILLER_34_525 ();
 sg13g2_decap_8 FILLER_34_532 ();
 sg13g2_decap_8 FILLER_34_539 ();
 sg13g2_decap_8 FILLER_34_546 ();
 sg13g2_decap_8 FILLER_34_553 ();
 sg13g2_decap_8 FILLER_34_560 ();
 sg13g2_decap_8 FILLER_34_567 ();
 sg13g2_decap_8 FILLER_34_574 ();
 sg13g2_decap_8 FILLER_34_581 ();
 sg13g2_decap_8 FILLER_34_588 ();
 sg13g2_decap_8 FILLER_34_595 ();
 sg13g2_decap_8 FILLER_34_602 ();
 sg13g2_decap_8 FILLER_34_609 ();
 sg13g2_decap_8 FILLER_34_616 ();
 sg13g2_decap_8 FILLER_34_623 ();
 sg13g2_decap_8 FILLER_34_630 ();
 sg13g2_decap_8 FILLER_34_637 ();
 sg13g2_decap_8 FILLER_34_644 ();
 sg13g2_decap_8 FILLER_34_651 ();
 sg13g2_decap_8 FILLER_34_658 ();
 sg13g2_decap_8 FILLER_34_665 ();
 sg13g2_decap_8 FILLER_34_672 ();
 sg13g2_decap_8 FILLER_34_679 ();
 sg13g2_decap_8 FILLER_34_686 ();
 sg13g2_decap_8 FILLER_34_693 ();
 sg13g2_decap_8 FILLER_34_700 ();
 sg13g2_decap_8 FILLER_34_707 ();
 sg13g2_decap_8 FILLER_34_714 ();
 sg13g2_decap_8 FILLER_34_721 ();
 sg13g2_decap_8 FILLER_34_728 ();
 sg13g2_decap_8 FILLER_34_735 ();
 sg13g2_decap_8 FILLER_34_742 ();
 sg13g2_decap_8 FILLER_34_749 ();
 sg13g2_decap_8 FILLER_34_756 ();
 sg13g2_decap_8 FILLER_34_763 ();
 sg13g2_decap_8 FILLER_34_770 ();
 sg13g2_decap_8 FILLER_34_777 ();
 sg13g2_decap_8 FILLER_34_784 ();
 sg13g2_decap_8 FILLER_34_791 ();
 sg13g2_decap_8 FILLER_34_798 ();
 sg13g2_decap_8 FILLER_34_805 ();
 sg13g2_decap_8 FILLER_34_812 ();
 sg13g2_decap_8 FILLER_34_819 ();
 sg13g2_decap_8 FILLER_34_826 ();
 sg13g2_decap_8 FILLER_34_833 ();
 sg13g2_decap_8 FILLER_34_840 ();
 sg13g2_decap_8 FILLER_34_847 ();
 sg13g2_decap_8 FILLER_34_854 ();
 sg13g2_decap_8 FILLER_34_861 ();
 sg13g2_decap_8 FILLER_34_868 ();
 sg13g2_decap_8 FILLER_34_875 ();
 sg13g2_decap_8 FILLER_34_882 ();
 sg13g2_decap_8 FILLER_34_889 ();
 sg13g2_decap_8 FILLER_34_896 ();
 sg13g2_decap_8 FILLER_34_903 ();
 sg13g2_decap_8 FILLER_34_910 ();
 sg13g2_decap_8 FILLER_34_917 ();
 sg13g2_decap_8 FILLER_34_924 ();
 sg13g2_decap_8 FILLER_34_931 ();
 sg13g2_decap_8 FILLER_34_938 ();
 sg13g2_decap_8 FILLER_34_945 ();
 sg13g2_decap_8 FILLER_34_952 ();
 sg13g2_decap_8 FILLER_34_959 ();
 sg13g2_decap_8 FILLER_34_966 ();
 sg13g2_decap_8 FILLER_34_973 ();
 sg13g2_decap_8 FILLER_34_980 ();
 sg13g2_decap_8 FILLER_34_987 ();
 sg13g2_decap_8 FILLER_34_994 ();
 sg13g2_decap_8 FILLER_34_1001 ();
 sg13g2_decap_8 FILLER_34_1008 ();
 sg13g2_decap_8 FILLER_34_1015 ();
 sg13g2_decap_8 FILLER_34_1022 ();
 sg13g2_decap_8 FILLER_34_1029 ();
 sg13g2_decap_8 FILLER_34_1036 ();
 sg13g2_decap_8 FILLER_34_1043 ();
 sg13g2_decap_8 FILLER_34_1050 ();
 sg13g2_decap_8 FILLER_34_1057 ();
 sg13g2_decap_8 FILLER_34_1064 ();
 sg13g2_decap_8 FILLER_34_1071 ();
 sg13g2_decap_8 FILLER_34_1078 ();
 sg13g2_decap_8 FILLER_34_1085 ();
 sg13g2_decap_8 FILLER_34_1092 ();
 sg13g2_decap_8 FILLER_34_1099 ();
 sg13g2_decap_8 FILLER_34_1106 ();
 sg13g2_decap_8 FILLER_34_1113 ();
 sg13g2_decap_8 FILLER_34_1120 ();
 sg13g2_decap_8 FILLER_34_1127 ();
 sg13g2_decap_8 FILLER_34_1134 ();
 sg13g2_decap_8 FILLER_34_1141 ();
 sg13g2_decap_8 FILLER_34_1148 ();
 sg13g2_decap_8 FILLER_34_1155 ();
 sg13g2_decap_8 FILLER_34_1162 ();
 sg13g2_decap_8 FILLER_34_1169 ();
 sg13g2_decap_8 FILLER_34_1176 ();
 sg13g2_decap_8 FILLER_34_1183 ();
 sg13g2_decap_8 FILLER_34_1190 ();
 sg13g2_decap_8 FILLER_34_1197 ();
 sg13g2_decap_8 FILLER_34_1204 ();
 sg13g2_decap_8 FILLER_34_1211 ();
 sg13g2_decap_8 FILLER_34_1218 ();
 sg13g2_decap_8 FILLER_34_1225 ();
 sg13g2_decap_8 FILLER_34_1232 ();
 sg13g2_decap_8 FILLER_34_1239 ();
 sg13g2_decap_8 FILLER_34_1246 ();
 sg13g2_decap_8 FILLER_34_1253 ();
 sg13g2_decap_8 FILLER_34_1260 ();
 sg13g2_decap_8 FILLER_34_1267 ();
 sg13g2_decap_8 FILLER_34_1274 ();
 sg13g2_decap_8 FILLER_34_1281 ();
 sg13g2_decap_8 FILLER_34_1288 ();
 sg13g2_decap_8 FILLER_34_1295 ();
 sg13g2_decap_8 FILLER_34_1302 ();
 sg13g2_decap_8 FILLER_34_1309 ();
 sg13g2_decap_8 FILLER_34_1316 ();
 sg13g2_decap_8 FILLER_34_1323 ();
 sg13g2_decap_8 FILLER_34_1330 ();
 sg13g2_decap_8 FILLER_34_1337 ();
 sg13g2_decap_8 FILLER_34_1344 ();
 sg13g2_decap_8 FILLER_34_1351 ();
 sg13g2_decap_8 FILLER_34_1358 ();
 sg13g2_decap_8 FILLER_34_1365 ();
 sg13g2_decap_8 FILLER_34_1372 ();
 sg13g2_decap_8 FILLER_34_1379 ();
 sg13g2_decap_8 FILLER_34_1386 ();
 sg13g2_decap_8 FILLER_34_1393 ();
 sg13g2_decap_8 FILLER_34_1400 ();
 sg13g2_decap_8 FILLER_34_1407 ();
 sg13g2_decap_8 FILLER_34_1414 ();
 sg13g2_decap_8 FILLER_34_1421 ();
 sg13g2_decap_8 FILLER_34_1428 ();
 sg13g2_decap_8 FILLER_34_1435 ();
 sg13g2_decap_8 FILLER_34_1442 ();
 sg13g2_decap_8 FILLER_34_1449 ();
 sg13g2_decap_8 FILLER_34_1456 ();
 sg13g2_decap_8 FILLER_34_1463 ();
 sg13g2_decap_8 FILLER_34_1470 ();
 sg13g2_decap_8 FILLER_34_1477 ();
 sg13g2_decap_8 FILLER_34_1484 ();
 sg13g2_decap_8 FILLER_34_1491 ();
 sg13g2_decap_8 FILLER_34_1498 ();
 sg13g2_decap_8 FILLER_34_1505 ();
 sg13g2_decap_8 FILLER_34_1512 ();
 sg13g2_decap_8 FILLER_34_1519 ();
 sg13g2_decap_8 FILLER_34_1526 ();
 sg13g2_decap_8 FILLER_34_1533 ();
 sg13g2_decap_8 FILLER_34_1540 ();
 sg13g2_decap_8 FILLER_34_1547 ();
 sg13g2_decap_8 FILLER_34_1554 ();
 sg13g2_decap_8 FILLER_34_1561 ();
 sg13g2_decap_8 FILLER_34_1568 ();
 sg13g2_decap_8 FILLER_34_1575 ();
 sg13g2_decap_8 FILLER_34_1582 ();
 sg13g2_decap_8 FILLER_34_1589 ();
 sg13g2_decap_8 FILLER_34_1596 ();
 sg13g2_decap_8 FILLER_34_1603 ();
 sg13g2_decap_8 FILLER_34_1610 ();
 sg13g2_decap_8 FILLER_34_1617 ();
 sg13g2_decap_8 FILLER_34_1624 ();
 sg13g2_decap_8 FILLER_34_1631 ();
 sg13g2_decap_8 FILLER_34_1638 ();
 sg13g2_decap_8 FILLER_34_1645 ();
 sg13g2_decap_8 FILLER_34_1652 ();
 sg13g2_decap_8 FILLER_34_1659 ();
 sg13g2_decap_8 FILLER_34_1666 ();
 sg13g2_decap_8 FILLER_34_1673 ();
 sg13g2_decap_8 FILLER_34_1680 ();
 sg13g2_decap_8 FILLER_34_1687 ();
 sg13g2_decap_8 FILLER_34_1694 ();
 sg13g2_decap_8 FILLER_34_1701 ();
 sg13g2_decap_8 FILLER_34_1708 ();
 sg13g2_decap_8 FILLER_34_1715 ();
 sg13g2_decap_8 FILLER_34_1722 ();
 sg13g2_decap_8 FILLER_34_1729 ();
 sg13g2_decap_8 FILLER_34_1736 ();
 sg13g2_decap_8 FILLER_34_1743 ();
 sg13g2_decap_8 FILLER_34_1750 ();
 sg13g2_decap_8 FILLER_34_1757 ();
 sg13g2_decap_8 FILLER_34_1764 ();
 sg13g2_decap_8 FILLER_34_1771 ();
 sg13g2_decap_8 FILLER_34_1778 ();
 sg13g2_decap_8 FILLER_34_1785 ();
 sg13g2_decap_8 FILLER_34_1792 ();
 sg13g2_decap_8 FILLER_34_1799 ();
 sg13g2_decap_8 FILLER_34_1806 ();
 sg13g2_decap_8 FILLER_34_1813 ();
 sg13g2_decap_8 FILLER_34_1820 ();
 sg13g2_decap_8 FILLER_34_1827 ();
 sg13g2_decap_8 FILLER_34_1834 ();
 sg13g2_decap_8 FILLER_34_1841 ();
 sg13g2_decap_8 FILLER_34_1848 ();
 sg13g2_decap_8 FILLER_34_1855 ();
 sg13g2_decap_8 FILLER_34_1862 ();
 sg13g2_decap_8 FILLER_34_1869 ();
 sg13g2_decap_8 FILLER_34_1876 ();
 sg13g2_decap_8 FILLER_34_1883 ();
 sg13g2_decap_8 FILLER_34_1890 ();
 sg13g2_decap_8 FILLER_34_1897 ();
 sg13g2_decap_8 FILLER_34_1904 ();
 sg13g2_decap_8 FILLER_34_1911 ();
 sg13g2_decap_8 FILLER_34_1918 ();
 sg13g2_decap_8 FILLER_34_1925 ();
 sg13g2_decap_8 FILLER_34_1932 ();
 sg13g2_decap_8 FILLER_34_1939 ();
 sg13g2_decap_8 FILLER_34_1946 ();
 sg13g2_decap_8 FILLER_34_1953 ();
 sg13g2_decap_8 FILLER_34_1960 ();
 sg13g2_decap_8 FILLER_34_1967 ();
 sg13g2_decap_8 FILLER_34_1974 ();
 sg13g2_decap_8 FILLER_34_1981 ();
 sg13g2_decap_8 FILLER_34_1988 ();
 sg13g2_decap_8 FILLER_34_1995 ();
 sg13g2_decap_8 FILLER_34_2002 ();
 sg13g2_decap_8 FILLER_34_2009 ();
 sg13g2_decap_8 FILLER_34_2016 ();
 sg13g2_decap_8 FILLER_34_2023 ();
 sg13g2_decap_8 FILLER_34_2030 ();
 sg13g2_decap_8 FILLER_34_2037 ();
 sg13g2_decap_8 FILLER_34_2044 ();
 sg13g2_decap_8 FILLER_34_2051 ();
 sg13g2_decap_8 FILLER_34_2058 ();
 sg13g2_decap_8 FILLER_34_2065 ();
 sg13g2_decap_8 FILLER_34_2072 ();
 sg13g2_decap_8 FILLER_34_2079 ();
 sg13g2_decap_8 FILLER_34_2086 ();
 sg13g2_decap_8 FILLER_34_2093 ();
 sg13g2_decap_8 FILLER_34_2100 ();
 sg13g2_decap_8 FILLER_34_2107 ();
 sg13g2_decap_8 FILLER_34_2114 ();
 sg13g2_decap_8 FILLER_34_2121 ();
 sg13g2_decap_8 FILLER_34_2128 ();
 sg13g2_decap_8 FILLER_34_2135 ();
 sg13g2_decap_8 FILLER_34_2142 ();
 sg13g2_decap_8 FILLER_34_2149 ();
 sg13g2_decap_8 FILLER_34_2156 ();
 sg13g2_decap_8 FILLER_34_2163 ();
 sg13g2_decap_8 FILLER_34_2170 ();
 sg13g2_decap_8 FILLER_34_2177 ();
 sg13g2_decap_8 FILLER_34_2184 ();
 sg13g2_decap_8 FILLER_34_2191 ();
 sg13g2_decap_8 FILLER_34_2198 ();
 sg13g2_decap_8 FILLER_34_2205 ();
 sg13g2_decap_8 FILLER_34_2212 ();
 sg13g2_decap_8 FILLER_34_2219 ();
 sg13g2_decap_8 FILLER_34_2226 ();
 sg13g2_decap_8 FILLER_34_2233 ();
 sg13g2_decap_8 FILLER_34_2240 ();
 sg13g2_decap_8 FILLER_34_2247 ();
 sg13g2_decap_8 FILLER_34_2254 ();
 sg13g2_decap_8 FILLER_34_2261 ();
 sg13g2_decap_8 FILLER_34_2268 ();
 sg13g2_decap_8 FILLER_34_2275 ();
 sg13g2_decap_8 FILLER_34_2282 ();
 sg13g2_decap_8 FILLER_34_2289 ();
 sg13g2_decap_8 FILLER_34_2296 ();
 sg13g2_decap_8 FILLER_34_2303 ();
 sg13g2_decap_8 FILLER_34_2310 ();
 sg13g2_decap_8 FILLER_34_2317 ();
 sg13g2_decap_8 FILLER_34_2324 ();
 sg13g2_decap_8 FILLER_34_2331 ();
 sg13g2_decap_8 FILLER_34_2338 ();
 sg13g2_decap_8 FILLER_34_2345 ();
 sg13g2_decap_8 FILLER_34_2352 ();
 sg13g2_decap_8 FILLER_34_2359 ();
 sg13g2_decap_8 FILLER_34_2366 ();
 sg13g2_decap_8 FILLER_34_2373 ();
 sg13g2_decap_8 FILLER_34_2380 ();
 sg13g2_decap_8 FILLER_34_2387 ();
 sg13g2_decap_8 FILLER_34_2394 ();
 sg13g2_decap_8 FILLER_34_2401 ();
 sg13g2_decap_8 FILLER_34_2408 ();
 sg13g2_decap_8 FILLER_34_2415 ();
 sg13g2_decap_8 FILLER_34_2422 ();
 sg13g2_decap_8 FILLER_34_2429 ();
 sg13g2_decap_8 FILLER_34_2436 ();
 sg13g2_decap_8 FILLER_34_2443 ();
 sg13g2_decap_8 FILLER_34_2450 ();
 sg13g2_decap_8 FILLER_34_2457 ();
 sg13g2_decap_8 FILLER_34_2464 ();
 sg13g2_decap_8 FILLER_34_2471 ();
 sg13g2_decap_8 FILLER_34_2478 ();
 sg13g2_decap_8 FILLER_34_2485 ();
 sg13g2_decap_8 FILLER_34_2492 ();
 sg13g2_decap_8 FILLER_34_2499 ();
 sg13g2_decap_8 FILLER_34_2506 ();
 sg13g2_decap_8 FILLER_34_2513 ();
 sg13g2_decap_8 FILLER_34_2520 ();
 sg13g2_decap_8 FILLER_34_2527 ();
 sg13g2_decap_8 FILLER_34_2534 ();
 sg13g2_decap_8 FILLER_34_2541 ();
 sg13g2_decap_8 FILLER_34_2548 ();
 sg13g2_decap_8 FILLER_34_2555 ();
 sg13g2_decap_8 FILLER_34_2562 ();
 sg13g2_decap_8 FILLER_34_2569 ();
 sg13g2_decap_8 FILLER_34_2576 ();
 sg13g2_decap_8 FILLER_34_2583 ();
 sg13g2_decap_8 FILLER_34_2590 ();
 sg13g2_decap_8 FILLER_34_2597 ();
 sg13g2_decap_8 FILLER_34_2604 ();
 sg13g2_decap_8 FILLER_34_2611 ();
 sg13g2_decap_8 FILLER_34_2618 ();
 sg13g2_decap_8 FILLER_34_2625 ();
 sg13g2_decap_8 FILLER_34_2632 ();
 sg13g2_decap_8 FILLER_34_2639 ();
 sg13g2_decap_8 FILLER_34_2646 ();
 sg13g2_decap_8 FILLER_34_2653 ();
 sg13g2_decap_8 FILLER_34_2660 ();
 sg13g2_decap_8 FILLER_34_2667 ();
 sg13g2_decap_8 FILLER_34_2674 ();
 sg13g2_decap_8 FILLER_34_2681 ();
 sg13g2_decap_8 FILLER_34_2688 ();
 sg13g2_decap_8 FILLER_34_2695 ();
 sg13g2_decap_8 FILLER_34_2702 ();
 sg13g2_decap_8 FILLER_34_2709 ();
 sg13g2_decap_8 FILLER_34_2716 ();
 sg13g2_decap_8 FILLER_34_2723 ();
 sg13g2_decap_8 FILLER_34_2730 ();
 sg13g2_decap_8 FILLER_34_2737 ();
 sg13g2_decap_8 FILLER_34_2744 ();
 sg13g2_decap_8 FILLER_34_2751 ();
 sg13g2_decap_8 FILLER_34_2758 ();
 sg13g2_decap_8 FILLER_34_2765 ();
 sg13g2_decap_8 FILLER_34_2772 ();
 sg13g2_decap_8 FILLER_34_2779 ();
 sg13g2_decap_8 FILLER_34_2786 ();
 sg13g2_decap_8 FILLER_34_2793 ();
 sg13g2_decap_8 FILLER_34_2800 ();
 sg13g2_decap_8 FILLER_34_2807 ();
 sg13g2_decap_8 FILLER_34_2814 ();
 sg13g2_decap_8 FILLER_34_2821 ();
 sg13g2_decap_8 FILLER_34_2828 ();
 sg13g2_decap_8 FILLER_34_2835 ();
 sg13g2_decap_8 FILLER_34_2842 ();
 sg13g2_decap_8 FILLER_34_2849 ();
 sg13g2_decap_8 FILLER_34_2856 ();
 sg13g2_decap_8 FILLER_34_2863 ();
 sg13g2_decap_8 FILLER_34_2870 ();
 sg13g2_decap_8 FILLER_34_2877 ();
 sg13g2_decap_8 FILLER_34_2884 ();
 sg13g2_decap_8 FILLER_34_2891 ();
 sg13g2_decap_8 FILLER_34_2898 ();
 sg13g2_decap_8 FILLER_34_2905 ();
 sg13g2_decap_8 FILLER_34_2912 ();
 sg13g2_decap_8 FILLER_34_2919 ();
 sg13g2_decap_8 FILLER_34_2926 ();
 sg13g2_decap_8 FILLER_34_2933 ();
 sg13g2_decap_8 FILLER_34_2940 ();
 sg13g2_decap_8 FILLER_34_2947 ();
 sg13g2_decap_8 FILLER_34_2954 ();
 sg13g2_decap_8 FILLER_34_2961 ();
 sg13g2_decap_8 FILLER_34_2968 ();
 sg13g2_decap_8 FILLER_34_2975 ();
 sg13g2_decap_8 FILLER_34_2982 ();
 sg13g2_decap_8 FILLER_34_2989 ();
 sg13g2_decap_8 FILLER_34_2996 ();
 sg13g2_decap_8 FILLER_34_3003 ();
 sg13g2_decap_8 FILLER_34_3010 ();
 sg13g2_decap_8 FILLER_34_3017 ();
 sg13g2_decap_8 FILLER_34_3024 ();
 sg13g2_decap_8 FILLER_34_3031 ();
 sg13g2_decap_8 FILLER_34_3038 ();
 sg13g2_decap_8 FILLER_34_3045 ();
 sg13g2_decap_8 FILLER_34_3052 ();
 sg13g2_decap_8 FILLER_34_3059 ();
 sg13g2_decap_8 FILLER_34_3066 ();
 sg13g2_decap_8 FILLER_34_3073 ();
 sg13g2_decap_8 FILLER_34_3080 ();
 sg13g2_decap_8 FILLER_34_3087 ();
 sg13g2_decap_8 FILLER_34_3094 ();
 sg13g2_decap_8 FILLER_34_3101 ();
 sg13g2_decap_8 FILLER_34_3108 ();
 sg13g2_decap_8 FILLER_34_3115 ();
 sg13g2_decap_8 FILLER_34_3122 ();
 sg13g2_decap_8 FILLER_34_3129 ();
 sg13g2_decap_8 FILLER_34_3136 ();
 sg13g2_decap_8 FILLER_34_3143 ();
 sg13g2_decap_8 FILLER_34_3150 ();
 sg13g2_decap_8 FILLER_34_3157 ();
 sg13g2_decap_8 FILLER_34_3164 ();
 sg13g2_decap_8 FILLER_34_3171 ();
 sg13g2_decap_8 FILLER_34_3178 ();
 sg13g2_decap_8 FILLER_34_3185 ();
 sg13g2_decap_8 FILLER_34_3192 ();
 sg13g2_decap_8 FILLER_34_3199 ();
 sg13g2_decap_8 FILLER_34_3206 ();
 sg13g2_decap_8 FILLER_34_3213 ();
 sg13g2_decap_8 FILLER_34_3220 ();
 sg13g2_decap_8 FILLER_34_3227 ();
 sg13g2_decap_8 FILLER_34_3234 ();
 sg13g2_decap_8 FILLER_34_3241 ();
 sg13g2_decap_8 FILLER_34_3248 ();
 sg13g2_decap_8 FILLER_34_3255 ();
 sg13g2_decap_8 FILLER_34_3262 ();
 sg13g2_decap_8 FILLER_34_3269 ();
 sg13g2_decap_8 FILLER_34_3276 ();
 sg13g2_decap_8 FILLER_34_3283 ();
 sg13g2_decap_8 FILLER_34_3290 ();
 sg13g2_decap_8 FILLER_34_3297 ();
 sg13g2_decap_8 FILLER_34_3304 ();
 sg13g2_decap_8 FILLER_34_3311 ();
 sg13g2_decap_8 FILLER_34_3318 ();
 sg13g2_decap_8 FILLER_34_3325 ();
 sg13g2_decap_8 FILLER_34_3332 ();
 sg13g2_decap_8 FILLER_34_3339 ();
 sg13g2_decap_8 FILLER_34_3346 ();
 sg13g2_decap_8 FILLER_34_3353 ();
 sg13g2_decap_8 FILLER_34_3360 ();
 sg13g2_decap_8 FILLER_34_3367 ();
 sg13g2_decap_8 FILLER_34_3374 ();
 sg13g2_decap_8 FILLER_34_3381 ();
 sg13g2_decap_8 FILLER_34_3388 ();
 sg13g2_decap_8 FILLER_34_3395 ();
 sg13g2_decap_8 FILLER_34_3402 ();
 sg13g2_decap_8 FILLER_34_3409 ();
 sg13g2_decap_8 FILLER_34_3416 ();
 sg13g2_decap_8 FILLER_34_3423 ();
 sg13g2_decap_8 FILLER_34_3430 ();
 sg13g2_decap_8 FILLER_34_3437 ();
 sg13g2_decap_8 FILLER_34_3444 ();
 sg13g2_decap_8 FILLER_34_3451 ();
 sg13g2_decap_8 FILLER_34_3458 ();
 sg13g2_decap_8 FILLER_34_3465 ();
 sg13g2_decap_8 FILLER_34_3472 ();
 sg13g2_decap_8 FILLER_34_3479 ();
 sg13g2_decap_8 FILLER_34_3486 ();
 sg13g2_decap_8 FILLER_34_3493 ();
 sg13g2_decap_8 FILLER_34_3500 ();
 sg13g2_decap_8 FILLER_34_3507 ();
 sg13g2_decap_8 FILLER_34_3514 ();
 sg13g2_decap_8 FILLER_34_3521 ();
 sg13g2_decap_8 FILLER_34_3528 ();
 sg13g2_decap_8 FILLER_34_3535 ();
 sg13g2_decap_8 FILLER_34_3542 ();
 sg13g2_decap_8 FILLER_34_3549 ();
 sg13g2_decap_8 FILLER_34_3556 ();
 sg13g2_decap_8 FILLER_34_3563 ();
 sg13g2_decap_8 FILLER_34_3570 ();
 sg13g2_fill_2 FILLER_34_3577 ();
 sg13g2_fill_1 FILLER_34_3579 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_decap_8 FILLER_35_245 ();
 sg13g2_decap_8 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_decap_8 FILLER_35_266 ();
 sg13g2_decap_8 FILLER_35_273 ();
 sg13g2_decap_8 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_decap_8 FILLER_35_294 ();
 sg13g2_decap_8 FILLER_35_301 ();
 sg13g2_decap_8 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_315 ();
 sg13g2_decap_8 FILLER_35_322 ();
 sg13g2_decap_8 FILLER_35_329 ();
 sg13g2_decap_8 FILLER_35_336 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_decap_8 FILLER_35_350 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_decap_8 FILLER_35_406 ();
 sg13g2_decap_8 FILLER_35_413 ();
 sg13g2_decap_8 FILLER_35_420 ();
 sg13g2_decap_8 FILLER_35_427 ();
 sg13g2_decap_8 FILLER_35_434 ();
 sg13g2_decap_8 FILLER_35_441 ();
 sg13g2_decap_8 FILLER_35_448 ();
 sg13g2_decap_8 FILLER_35_455 ();
 sg13g2_decap_8 FILLER_35_462 ();
 sg13g2_decap_8 FILLER_35_469 ();
 sg13g2_decap_8 FILLER_35_476 ();
 sg13g2_decap_8 FILLER_35_483 ();
 sg13g2_decap_8 FILLER_35_490 ();
 sg13g2_decap_8 FILLER_35_497 ();
 sg13g2_decap_8 FILLER_35_504 ();
 sg13g2_decap_8 FILLER_35_511 ();
 sg13g2_decap_8 FILLER_35_518 ();
 sg13g2_decap_8 FILLER_35_525 ();
 sg13g2_decap_8 FILLER_35_532 ();
 sg13g2_decap_8 FILLER_35_539 ();
 sg13g2_decap_8 FILLER_35_546 ();
 sg13g2_decap_8 FILLER_35_553 ();
 sg13g2_decap_8 FILLER_35_560 ();
 sg13g2_decap_8 FILLER_35_567 ();
 sg13g2_decap_8 FILLER_35_574 ();
 sg13g2_decap_8 FILLER_35_581 ();
 sg13g2_decap_8 FILLER_35_588 ();
 sg13g2_decap_8 FILLER_35_595 ();
 sg13g2_decap_8 FILLER_35_602 ();
 sg13g2_decap_8 FILLER_35_609 ();
 sg13g2_decap_8 FILLER_35_616 ();
 sg13g2_decap_8 FILLER_35_623 ();
 sg13g2_decap_8 FILLER_35_630 ();
 sg13g2_decap_8 FILLER_35_637 ();
 sg13g2_decap_8 FILLER_35_644 ();
 sg13g2_decap_8 FILLER_35_651 ();
 sg13g2_decap_8 FILLER_35_658 ();
 sg13g2_decap_8 FILLER_35_665 ();
 sg13g2_decap_8 FILLER_35_672 ();
 sg13g2_decap_8 FILLER_35_679 ();
 sg13g2_decap_8 FILLER_35_686 ();
 sg13g2_decap_8 FILLER_35_693 ();
 sg13g2_decap_8 FILLER_35_700 ();
 sg13g2_decap_8 FILLER_35_707 ();
 sg13g2_decap_8 FILLER_35_714 ();
 sg13g2_decap_8 FILLER_35_721 ();
 sg13g2_decap_8 FILLER_35_728 ();
 sg13g2_decap_8 FILLER_35_735 ();
 sg13g2_decap_8 FILLER_35_742 ();
 sg13g2_decap_8 FILLER_35_749 ();
 sg13g2_decap_8 FILLER_35_756 ();
 sg13g2_decap_8 FILLER_35_763 ();
 sg13g2_decap_8 FILLER_35_770 ();
 sg13g2_decap_8 FILLER_35_777 ();
 sg13g2_decap_8 FILLER_35_784 ();
 sg13g2_decap_8 FILLER_35_791 ();
 sg13g2_decap_8 FILLER_35_798 ();
 sg13g2_decap_8 FILLER_35_805 ();
 sg13g2_decap_8 FILLER_35_812 ();
 sg13g2_decap_8 FILLER_35_819 ();
 sg13g2_decap_8 FILLER_35_826 ();
 sg13g2_decap_8 FILLER_35_833 ();
 sg13g2_decap_8 FILLER_35_840 ();
 sg13g2_decap_8 FILLER_35_847 ();
 sg13g2_decap_8 FILLER_35_854 ();
 sg13g2_decap_8 FILLER_35_861 ();
 sg13g2_decap_8 FILLER_35_868 ();
 sg13g2_decap_8 FILLER_35_875 ();
 sg13g2_decap_8 FILLER_35_882 ();
 sg13g2_decap_8 FILLER_35_889 ();
 sg13g2_decap_8 FILLER_35_896 ();
 sg13g2_decap_8 FILLER_35_903 ();
 sg13g2_decap_8 FILLER_35_910 ();
 sg13g2_decap_8 FILLER_35_917 ();
 sg13g2_decap_8 FILLER_35_924 ();
 sg13g2_decap_8 FILLER_35_931 ();
 sg13g2_decap_8 FILLER_35_938 ();
 sg13g2_decap_8 FILLER_35_945 ();
 sg13g2_decap_8 FILLER_35_952 ();
 sg13g2_decap_8 FILLER_35_959 ();
 sg13g2_decap_8 FILLER_35_966 ();
 sg13g2_decap_8 FILLER_35_973 ();
 sg13g2_decap_8 FILLER_35_980 ();
 sg13g2_decap_8 FILLER_35_987 ();
 sg13g2_decap_8 FILLER_35_994 ();
 sg13g2_decap_8 FILLER_35_1001 ();
 sg13g2_decap_8 FILLER_35_1008 ();
 sg13g2_decap_8 FILLER_35_1015 ();
 sg13g2_decap_8 FILLER_35_1022 ();
 sg13g2_decap_8 FILLER_35_1029 ();
 sg13g2_decap_8 FILLER_35_1036 ();
 sg13g2_decap_8 FILLER_35_1043 ();
 sg13g2_decap_8 FILLER_35_1050 ();
 sg13g2_decap_8 FILLER_35_1057 ();
 sg13g2_decap_8 FILLER_35_1064 ();
 sg13g2_decap_8 FILLER_35_1071 ();
 sg13g2_decap_8 FILLER_35_1078 ();
 sg13g2_decap_8 FILLER_35_1085 ();
 sg13g2_decap_8 FILLER_35_1092 ();
 sg13g2_decap_8 FILLER_35_1099 ();
 sg13g2_decap_8 FILLER_35_1106 ();
 sg13g2_decap_8 FILLER_35_1113 ();
 sg13g2_decap_8 FILLER_35_1120 ();
 sg13g2_decap_8 FILLER_35_1127 ();
 sg13g2_decap_8 FILLER_35_1134 ();
 sg13g2_decap_8 FILLER_35_1141 ();
 sg13g2_decap_8 FILLER_35_1148 ();
 sg13g2_decap_8 FILLER_35_1155 ();
 sg13g2_decap_8 FILLER_35_1162 ();
 sg13g2_decap_8 FILLER_35_1169 ();
 sg13g2_decap_8 FILLER_35_1176 ();
 sg13g2_decap_8 FILLER_35_1183 ();
 sg13g2_decap_8 FILLER_35_1190 ();
 sg13g2_decap_8 FILLER_35_1197 ();
 sg13g2_decap_8 FILLER_35_1204 ();
 sg13g2_decap_8 FILLER_35_1211 ();
 sg13g2_decap_8 FILLER_35_1218 ();
 sg13g2_decap_8 FILLER_35_1225 ();
 sg13g2_decap_8 FILLER_35_1232 ();
 sg13g2_decap_8 FILLER_35_1239 ();
 sg13g2_decap_8 FILLER_35_1246 ();
 sg13g2_decap_8 FILLER_35_1253 ();
 sg13g2_decap_8 FILLER_35_1260 ();
 sg13g2_decap_8 FILLER_35_1267 ();
 sg13g2_decap_8 FILLER_35_1274 ();
 sg13g2_decap_8 FILLER_35_1281 ();
 sg13g2_decap_8 FILLER_35_1288 ();
 sg13g2_decap_8 FILLER_35_1295 ();
 sg13g2_decap_8 FILLER_35_1302 ();
 sg13g2_decap_8 FILLER_35_1309 ();
 sg13g2_decap_8 FILLER_35_1316 ();
 sg13g2_decap_8 FILLER_35_1323 ();
 sg13g2_decap_8 FILLER_35_1330 ();
 sg13g2_decap_8 FILLER_35_1337 ();
 sg13g2_decap_8 FILLER_35_1344 ();
 sg13g2_decap_8 FILLER_35_1351 ();
 sg13g2_decap_8 FILLER_35_1358 ();
 sg13g2_decap_8 FILLER_35_1365 ();
 sg13g2_decap_8 FILLER_35_1372 ();
 sg13g2_decap_8 FILLER_35_1379 ();
 sg13g2_decap_8 FILLER_35_1386 ();
 sg13g2_decap_8 FILLER_35_1393 ();
 sg13g2_decap_8 FILLER_35_1400 ();
 sg13g2_decap_8 FILLER_35_1407 ();
 sg13g2_decap_8 FILLER_35_1414 ();
 sg13g2_decap_8 FILLER_35_1421 ();
 sg13g2_decap_8 FILLER_35_1428 ();
 sg13g2_decap_8 FILLER_35_1435 ();
 sg13g2_decap_8 FILLER_35_1442 ();
 sg13g2_decap_8 FILLER_35_1449 ();
 sg13g2_decap_8 FILLER_35_1456 ();
 sg13g2_decap_8 FILLER_35_1463 ();
 sg13g2_decap_8 FILLER_35_1470 ();
 sg13g2_decap_8 FILLER_35_1477 ();
 sg13g2_decap_8 FILLER_35_1484 ();
 sg13g2_decap_8 FILLER_35_1491 ();
 sg13g2_decap_8 FILLER_35_1498 ();
 sg13g2_decap_8 FILLER_35_1505 ();
 sg13g2_decap_8 FILLER_35_1512 ();
 sg13g2_decap_8 FILLER_35_1519 ();
 sg13g2_decap_8 FILLER_35_1526 ();
 sg13g2_decap_8 FILLER_35_1533 ();
 sg13g2_decap_8 FILLER_35_1540 ();
 sg13g2_decap_8 FILLER_35_1547 ();
 sg13g2_decap_8 FILLER_35_1554 ();
 sg13g2_decap_8 FILLER_35_1561 ();
 sg13g2_decap_8 FILLER_35_1568 ();
 sg13g2_decap_8 FILLER_35_1575 ();
 sg13g2_decap_8 FILLER_35_1582 ();
 sg13g2_decap_8 FILLER_35_1589 ();
 sg13g2_decap_8 FILLER_35_1596 ();
 sg13g2_decap_8 FILLER_35_1603 ();
 sg13g2_decap_8 FILLER_35_1610 ();
 sg13g2_decap_8 FILLER_35_1617 ();
 sg13g2_decap_8 FILLER_35_1624 ();
 sg13g2_decap_8 FILLER_35_1631 ();
 sg13g2_decap_8 FILLER_35_1638 ();
 sg13g2_decap_8 FILLER_35_1645 ();
 sg13g2_decap_8 FILLER_35_1652 ();
 sg13g2_decap_8 FILLER_35_1659 ();
 sg13g2_decap_8 FILLER_35_1666 ();
 sg13g2_decap_8 FILLER_35_1673 ();
 sg13g2_decap_8 FILLER_35_1680 ();
 sg13g2_decap_8 FILLER_35_1687 ();
 sg13g2_decap_8 FILLER_35_1694 ();
 sg13g2_decap_8 FILLER_35_1701 ();
 sg13g2_decap_8 FILLER_35_1708 ();
 sg13g2_decap_8 FILLER_35_1715 ();
 sg13g2_decap_8 FILLER_35_1722 ();
 sg13g2_decap_8 FILLER_35_1729 ();
 sg13g2_decap_8 FILLER_35_1736 ();
 sg13g2_decap_8 FILLER_35_1743 ();
 sg13g2_decap_8 FILLER_35_1750 ();
 sg13g2_decap_8 FILLER_35_1757 ();
 sg13g2_decap_8 FILLER_35_1764 ();
 sg13g2_decap_8 FILLER_35_1771 ();
 sg13g2_decap_8 FILLER_35_1778 ();
 sg13g2_decap_8 FILLER_35_1785 ();
 sg13g2_decap_8 FILLER_35_1792 ();
 sg13g2_decap_8 FILLER_35_1799 ();
 sg13g2_decap_8 FILLER_35_1806 ();
 sg13g2_decap_8 FILLER_35_1813 ();
 sg13g2_decap_8 FILLER_35_1820 ();
 sg13g2_decap_8 FILLER_35_1827 ();
 sg13g2_decap_8 FILLER_35_1834 ();
 sg13g2_decap_8 FILLER_35_1841 ();
 sg13g2_decap_8 FILLER_35_1848 ();
 sg13g2_decap_8 FILLER_35_1855 ();
 sg13g2_decap_8 FILLER_35_1862 ();
 sg13g2_decap_8 FILLER_35_1869 ();
 sg13g2_decap_8 FILLER_35_1876 ();
 sg13g2_decap_8 FILLER_35_1883 ();
 sg13g2_decap_8 FILLER_35_1890 ();
 sg13g2_decap_8 FILLER_35_1897 ();
 sg13g2_decap_8 FILLER_35_1904 ();
 sg13g2_decap_8 FILLER_35_1911 ();
 sg13g2_decap_8 FILLER_35_1918 ();
 sg13g2_decap_8 FILLER_35_1925 ();
 sg13g2_decap_8 FILLER_35_1932 ();
 sg13g2_decap_8 FILLER_35_1939 ();
 sg13g2_decap_8 FILLER_35_1946 ();
 sg13g2_decap_8 FILLER_35_1953 ();
 sg13g2_decap_8 FILLER_35_1960 ();
 sg13g2_decap_8 FILLER_35_1967 ();
 sg13g2_decap_8 FILLER_35_1974 ();
 sg13g2_decap_8 FILLER_35_1981 ();
 sg13g2_decap_8 FILLER_35_1988 ();
 sg13g2_decap_8 FILLER_35_1995 ();
 sg13g2_decap_8 FILLER_35_2002 ();
 sg13g2_decap_8 FILLER_35_2009 ();
 sg13g2_decap_8 FILLER_35_2016 ();
 sg13g2_decap_8 FILLER_35_2023 ();
 sg13g2_decap_8 FILLER_35_2030 ();
 sg13g2_decap_8 FILLER_35_2037 ();
 sg13g2_decap_8 FILLER_35_2044 ();
 sg13g2_decap_8 FILLER_35_2051 ();
 sg13g2_decap_8 FILLER_35_2058 ();
 sg13g2_decap_8 FILLER_35_2065 ();
 sg13g2_decap_8 FILLER_35_2072 ();
 sg13g2_decap_8 FILLER_35_2079 ();
 sg13g2_decap_8 FILLER_35_2086 ();
 sg13g2_decap_8 FILLER_35_2093 ();
 sg13g2_decap_8 FILLER_35_2100 ();
 sg13g2_decap_8 FILLER_35_2107 ();
 sg13g2_decap_8 FILLER_35_2114 ();
 sg13g2_decap_8 FILLER_35_2121 ();
 sg13g2_decap_8 FILLER_35_2128 ();
 sg13g2_decap_8 FILLER_35_2135 ();
 sg13g2_decap_8 FILLER_35_2142 ();
 sg13g2_decap_8 FILLER_35_2149 ();
 sg13g2_decap_8 FILLER_35_2156 ();
 sg13g2_decap_8 FILLER_35_2163 ();
 sg13g2_decap_8 FILLER_35_2170 ();
 sg13g2_decap_8 FILLER_35_2177 ();
 sg13g2_decap_8 FILLER_35_2184 ();
 sg13g2_decap_8 FILLER_35_2191 ();
 sg13g2_decap_8 FILLER_35_2198 ();
 sg13g2_decap_8 FILLER_35_2205 ();
 sg13g2_decap_8 FILLER_35_2212 ();
 sg13g2_decap_8 FILLER_35_2219 ();
 sg13g2_decap_8 FILLER_35_2226 ();
 sg13g2_decap_8 FILLER_35_2233 ();
 sg13g2_decap_8 FILLER_35_2240 ();
 sg13g2_decap_8 FILLER_35_2247 ();
 sg13g2_decap_8 FILLER_35_2254 ();
 sg13g2_decap_8 FILLER_35_2261 ();
 sg13g2_decap_8 FILLER_35_2268 ();
 sg13g2_decap_8 FILLER_35_2275 ();
 sg13g2_decap_8 FILLER_35_2282 ();
 sg13g2_decap_8 FILLER_35_2289 ();
 sg13g2_decap_8 FILLER_35_2296 ();
 sg13g2_decap_8 FILLER_35_2303 ();
 sg13g2_decap_8 FILLER_35_2310 ();
 sg13g2_decap_8 FILLER_35_2317 ();
 sg13g2_decap_8 FILLER_35_2324 ();
 sg13g2_decap_8 FILLER_35_2331 ();
 sg13g2_decap_8 FILLER_35_2338 ();
 sg13g2_decap_8 FILLER_35_2345 ();
 sg13g2_decap_8 FILLER_35_2352 ();
 sg13g2_decap_8 FILLER_35_2359 ();
 sg13g2_decap_8 FILLER_35_2366 ();
 sg13g2_decap_8 FILLER_35_2373 ();
 sg13g2_decap_8 FILLER_35_2380 ();
 sg13g2_decap_8 FILLER_35_2387 ();
 sg13g2_decap_8 FILLER_35_2394 ();
 sg13g2_decap_8 FILLER_35_2401 ();
 sg13g2_decap_8 FILLER_35_2408 ();
 sg13g2_decap_8 FILLER_35_2415 ();
 sg13g2_decap_8 FILLER_35_2422 ();
 sg13g2_decap_8 FILLER_35_2429 ();
 sg13g2_decap_8 FILLER_35_2436 ();
 sg13g2_decap_8 FILLER_35_2443 ();
 sg13g2_decap_8 FILLER_35_2450 ();
 sg13g2_decap_8 FILLER_35_2457 ();
 sg13g2_decap_8 FILLER_35_2464 ();
 sg13g2_decap_8 FILLER_35_2471 ();
 sg13g2_decap_8 FILLER_35_2478 ();
 sg13g2_decap_8 FILLER_35_2485 ();
 sg13g2_decap_8 FILLER_35_2492 ();
 sg13g2_decap_8 FILLER_35_2499 ();
 sg13g2_decap_8 FILLER_35_2506 ();
 sg13g2_decap_8 FILLER_35_2513 ();
 sg13g2_decap_8 FILLER_35_2520 ();
 sg13g2_decap_8 FILLER_35_2527 ();
 sg13g2_decap_8 FILLER_35_2534 ();
 sg13g2_decap_8 FILLER_35_2541 ();
 sg13g2_decap_8 FILLER_35_2548 ();
 sg13g2_decap_8 FILLER_35_2555 ();
 sg13g2_decap_8 FILLER_35_2562 ();
 sg13g2_decap_8 FILLER_35_2569 ();
 sg13g2_decap_8 FILLER_35_2576 ();
 sg13g2_decap_8 FILLER_35_2583 ();
 sg13g2_decap_8 FILLER_35_2590 ();
 sg13g2_decap_8 FILLER_35_2597 ();
 sg13g2_decap_8 FILLER_35_2604 ();
 sg13g2_decap_8 FILLER_35_2611 ();
 sg13g2_decap_8 FILLER_35_2618 ();
 sg13g2_decap_8 FILLER_35_2625 ();
 sg13g2_decap_8 FILLER_35_2632 ();
 sg13g2_decap_8 FILLER_35_2639 ();
 sg13g2_decap_8 FILLER_35_2646 ();
 sg13g2_decap_8 FILLER_35_2653 ();
 sg13g2_decap_8 FILLER_35_2660 ();
 sg13g2_decap_8 FILLER_35_2667 ();
 sg13g2_decap_8 FILLER_35_2674 ();
 sg13g2_decap_8 FILLER_35_2681 ();
 sg13g2_decap_8 FILLER_35_2688 ();
 sg13g2_decap_8 FILLER_35_2695 ();
 sg13g2_decap_8 FILLER_35_2702 ();
 sg13g2_decap_8 FILLER_35_2709 ();
 sg13g2_decap_8 FILLER_35_2716 ();
 sg13g2_decap_8 FILLER_35_2723 ();
 sg13g2_decap_8 FILLER_35_2730 ();
 sg13g2_decap_8 FILLER_35_2737 ();
 sg13g2_decap_8 FILLER_35_2744 ();
 sg13g2_decap_8 FILLER_35_2751 ();
 sg13g2_decap_8 FILLER_35_2758 ();
 sg13g2_decap_8 FILLER_35_2765 ();
 sg13g2_decap_8 FILLER_35_2772 ();
 sg13g2_decap_8 FILLER_35_2779 ();
 sg13g2_decap_8 FILLER_35_2786 ();
 sg13g2_decap_8 FILLER_35_2793 ();
 sg13g2_decap_8 FILLER_35_2800 ();
 sg13g2_decap_8 FILLER_35_2807 ();
 sg13g2_decap_8 FILLER_35_2814 ();
 sg13g2_decap_8 FILLER_35_2821 ();
 sg13g2_decap_8 FILLER_35_2828 ();
 sg13g2_decap_8 FILLER_35_2835 ();
 sg13g2_decap_8 FILLER_35_2842 ();
 sg13g2_decap_8 FILLER_35_2849 ();
 sg13g2_decap_8 FILLER_35_2856 ();
 sg13g2_decap_8 FILLER_35_2863 ();
 sg13g2_decap_8 FILLER_35_2870 ();
 sg13g2_decap_8 FILLER_35_2877 ();
 sg13g2_decap_8 FILLER_35_2884 ();
 sg13g2_decap_8 FILLER_35_2891 ();
 sg13g2_decap_8 FILLER_35_2898 ();
 sg13g2_decap_8 FILLER_35_2905 ();
 sg13g2_decap_8 FILLER_35_2912 ();
 sg13g2_decap_8 FILLER_35_2919 ();
 sg13g2_decap_8 FILLER_35_2926 ();
 sg13g2_decap_8 FILLER_35_2933 ();
 sg13g2_decap_8 FILLER_35_2940 ();
 sg13g2_decap_8 FILLER_35_2947 ();
 sg13g2_decap_8 FILLER_35_2954 ();
 sg13g2_decap_8 FILLER_35_2961 ();
 sg13g2_decap_8 FILLER_35_2968 ();
 sg13g2_decap_8 FILLER_35_2975 ();
 sg13g2_decap_8 FILLER_35_2982 ();
 sg13g2_decap_8 FILLER_35_2989 ();
 sg13g2_decap_8 FILLER_35_2996 ();
 sg13g2_decap_8 FILLER_35_3003 ();
 sg13g2_decap_8 FILLER_35_3010 ();
 sg13g2_decap_8 FILLER_35_3017 ();
 sg13g2_decap_8 FILLER_35_3024 ();
 sg13g2_decap_8 FILLER_35_3031 ();
 sg13g2_decap_8 FILLER_35_3038 ();
 sg13g2_decap_8 FILLER_35_3045 ();
 sg13g2_decap_8 FILLER_35_3052 ();
 sg13g2_decap_8 FILLER_35_3059 ();
 sg13g2_decap_8 FILLER_35_3066 ();
 sg13g2_decap_8 FILLER_35_3073 ();
 sg13g2_decap_8 FILLER_35_3080 ();
 sg13g2_decap_8 FILLER_35_3087 ();
 sg13g2_decap_8 FILLER_35_3094 ();
 sg13g2_decap_8 FILLER_35_3101 ();
 sg13g2_decap_8 FILLER_35_3108 ();
 sg13g2_decap_8 FILLER_35_3115 ();
 sg13g2_decap_8 FILLER_35_3122 ();
 sg13g2_decap_8 FILLER_35_3129 ();
 sg13g2_decap_8 FILLER_35_3136 ();
 sg13g2_decap_8 FILLER_35_3143 ();
 sg13g2_decap_8 FILLER_35_3150 ();
 sg13g2_decap_8 FILLER_35_3157 ();
 sg13g2_decap_8 FILLER_35_3164 ();
 sg13g2_decap_8 FILLER_35_3171 ();
 sg13g2_decap_8 FILLER_35_3178 ();
 sg13g2_decap_8 FILLER_35_3185 ();
 sg13g2_decap_8 FILLER_35_3192 ();
 sg13g2_decap_8 FILLER_35_3199 ();
 sg13g2_decap_8 FILLER_35_3206 ();
 sg13g2_decap_8 FILLER_35_3213 ();
 sg13g2_decap_8 FILLER_35_3220 ();
 sg13g2_decap_8 FILLER_35_3227 ();
 sg13g2_decap_8 FILLER_35_3234 ();
 sg13g2_decap_8 FILLER_35_3241 ();
 sg13g2_decap_8 FILLER_35_3248 ();
 sg13g2_decap_8 FILLER_35_3255 ();
 sg13g2_decap_8 FILLER_35_3262 ();
 sg13g2_decap_8 FILLER_35_3269 ();
 sg13g2_decap_8 FILLER_35_3276 ();
 sg13g2_decap_8 FILLER_35_3283 ();
 sg13g2_decap_8 FILLER_35_3290 ();
 sg13g2_decap_8 FILLER_35_3297 ();
 sg13g2_decap_8 FILLER_35_3304 ();
 sg13g2_decap_8 FILLER_35_3311 ();
 sg13g2_decap_8 FILLER_35_3318 ();
 sg13g2_decap_8 FILLER_35_3325 ();
 sg13g2_decap_8 FILLER_35_3332 ();
 sg13g2_decap_8 FILLER_35_3339 ();
 sg13g2_decap_8 FILLER_35_3346 ();
 sg13g2_decap_8 FILLER_35_3353 ();
 sg13g2_decap_8 FILLER_35_3360 ();
 sg13g2_decap_8 FILLER_35_3367 ();
 sg13g2_decap_8 FILLER_35_3374 ();
 sg13g2_decap_8 FILLER_35_3381 ();
 sg13g2_decap_8 FILLER_35_3388 ();
 sg13g2_decap_8 FILLER_35_3395 ();
 sg13g2_decap_8 FILLER_35_3402 ();
 sg13g2_decap_8 FILLER_35_3409 ();
 sg13g2_decap_8 FILLER_35_3416 ();
 sg13g2_decap_8 FILLER_35_3423 ();
 sg13g2_decap_8 FILLER_35_3430 ();
 sg13g2_decap_8 FILLER_35_3437 ();
 sg13g2_decap_8 FILLER_35_3444 ();
 sg13g2_decap_8 FILLER_35_3451 ();
 sg13g2_decap_8 FILLER_35_3458 ();
 sg13g2_decap_8 FILLER_35_3465 ();
 sg13g2_decap_8 FILLER_35_3472 ();
 sg13g2_decap_8 FILLER_35_3479 ();
 sg13g2_decap_8 FILLER_35_3486 ();
 sg13g2_decap_8 FILLER_35_3493 ();
 sg13g2_decap_8 FILLER_35_3500 ();
 sg13g2_decap_8 FILLER_35_3507 ();
 sg13g2_decap_8 FILLER_35_3514 ();
 sg13g2_decap_8 FILLER_35_3521 ();
 sg13g2_decap_8 FILLER_35_3528 ();
 sg13g2_decap_8 FILLER_35_3535 ();
 sg13g2_decap_8 FILLER_35_3542 ();
 sg13g2_decap_8 FILLER_35_3549 ();
 sg13g2_decap_8 FILLER_35_3556 ();
 sg13g2_decap_8 FILLER_35_3563 ();
 sg13g2_decap_8 FILLER_35_3570 ();
 sg13g2_fill_2 FILLER_35_3577 ();
 sg13g2_fill_1 FILLER_35_3579 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_decap_8 FILLER_36_231 ();
 sg13g2_decap_8 FILLER_36_238 ();
 sg13g2_decap_8 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_252 ();
 sg13g2_decap_8 FILLER_36_259 ();
 sg13g2_decap_8 FILLER_36_266 ();
 sg13g2_decap_8 FILLER_36_273 ();
 sg13g2_decap_8 FILLER_36_280 ();
 sg13g2_decap_8 FILLER_36_287 ();
 sg13g2_decap_8 FILLER_36_294 ();
 sg13g2_decap_8 FILLER_36_301 ();
 sg13g2_decap_8 FILLER_36_308 ();
 sg13g2_decap_8 FILLER_36_315 ();
 sg13g2_decap_8 FILLER_36_322 ();
 sg13g2_decap_8 FILLER_36_329 ();
 sg13g2_decap_8 FILLER_36_336 ();
 sg13g2_decap_8 FILLER_36_343 ();
 sg13g2_decap_8 FILLER_36_350 ();
 sg13g2_decap_8 FILLER_36_357 ();
 sg13g2_decap_8 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_385 ();
 sg13g2_decap_8 FILLER_36_392 ();
 sg13g2_decap_8 FILLER_36_399 ();
 sg13g2_decap_8 FILLER_36_406 ();
 sg13g2_decap_8 FILLER_36_413 ();
 sg13g2_decap_8 FILLER_36_420 ();
 sg13g2_decap_8 FILLER_36_427 ();
 sg13g2_decap_8 FILLER_36_434 ();
 sg13g2_decap_8 FILLER_36_441 ();
 sg13g2_decap_8 FILLER_36_448 ();
 sg13g2_decap_8 FILLER_36_455 ();
 sg13g2_decap_8 FILLER_36_462 ();
 sg13g2_decap_8 FILLER_36_469 ();
 sg13g2_decap_8 FILLER_36_476 ();
 sg13g2_decap_8 FILLER_36_483 ();
 sg13g2_decap_8 FILLER_36_490 ();
 sg13g2_decap_8 FILLER_36_497 ();
 sg13g2_decap_8 FILLER_36_504 ();
 sg13g2_decap_8 FILLER_36_511 ();
 sg13g2_decap_8 FILLER_36_518 ();
 sg13g2_decap_8 FILLER_36_525 ();
 sg13g2_decap_8 FILLER_36_532 ();
 sg13g2_decap_8 FILLER_36_539 ();
 sg13g2_decap_8 FILLER_36_546 ();
 sg13g2_decap_8 FILLER_36_553 ();
 sg13g2_decap_8 FILLER_36_560 ();
 sg13g2_decap_8 FILLER_36_567 ();
 sg13g2_decap_8 FILLER_36_574 ();
 sg13g2_decap_8 FILLER_36_581 ();
 sg13g2_decap_8 FILLER_36_588 ();
 sg13g2_decap_8 FILLER_36_595 ();
 sg13g2_decap_8 FILLER_36_602 ();
 sg13g2_decap_8 FILLER_36_609 ();
 sg13g2_decap_8 FILLER_36_616 ();
 sg13g2_decap_8 FILLER_36_623 ();
 sg13g2_decap_8 FILLER_36_630 ();
 sg13g2_decap_8 FILLER_36_637 ();
 sg13g2_decap_8 FILLER_36_644 ();
 sg13g2_decap_8 FILLER_36_651 ();
 sg13g2_decap_8 FILLER_36_658 ();
 sg13g2_decap_8 FILLER_36_665 ();
 sg13g2_decap_8 FILLER_36_672 ();
 sg13g2_decap_8 FILLER_36_679 ();
 sg13g2_decap_8 FILLER_36_686 ();
 sg13g2_decap_8 FILLER_36_693 ();
 sg13g2_decap_8 FILLER_36_700 ();
 sg13g2_decap_8 FILLER_36_707 ();
 sg13g2_decap_8 FILLER_36_714 ();
 sg13g2_decap_8 FILLER_36_721 ();
 sg13g2_decap_8 FILLER_36_728 ();
 sg13g2_decap_8 FILLER_36_735 ();
 sg13g2_decap_8 FILLER_36_742 ();
 sg13g2_decap_8 FILLER_36_749 ();
 sg13g2_decap_8 FILLER_36_756 ();
 sg13g2_decap_8 FILLER_36_763 ();
 sg13g2_decap_8 FILLER_36_770 ();
 sg13g2_decap_8 FILLER_36_777 ();
 sg13g2_decap_8 FILLER_36_784 ();
 sg13g2_decap_8 FILLER_36_791 ();
 sg13g2_decap_8 FILLER_36_798 ();
 sg13g2_decap_8 FILLER_36_805 ();
 sg13g2_decap_8 FILLER_36_812 ();
 sg13g2_decap_8 FILLER_36_819 ();
 sg13g2_decap_8 FILLER_36_826 ();
 sg13g2_decap_8 FILLER_36_833 ();
 sg13g2_decap_8 FILLER_36_840 ();
 sg13g2_decap_8 FILLER_36_847 ();
 sg13g2_decap_8 FILLER_36_854 ();
 sg13g2_decap_8 FILLER_36_861 ();
 sg13g2_decap_8 FILLER_36_868 ();
 sg13g2_decap_8 FILLER_36_875 ();
 sg13g2_decap_8 FILLER_36_882 ();
 sg13g2_decap_8 FILLER_36_889 ();
 sg13g2_decap_8 FILLER_36_896 ();
 sg13g2_decap_8 FILLER_36_903 ();
 sg13g2_decap_8 FILLER_36_910 ();
 sg13g2_decap_8 FILLER_36_917 ();
 sg13g2_decap_8 FILLER_36_924 ();
 sg13g2_decap_8 FILLER_36_931 ();
 sg13g2_decap_8 FILLER_36_938 ();
 sg13g2_decap_8 FILLER_36_945 ();
 sg13g2_decap_8 FILLER_36_952 ();
 sg13g2_decap_8 FILLER_36_959 ();
 sg13g2_decap_8 FILLER_36_966 ();
 sg13g2_decap_8 FILLER_36_973 ();
 sg13g2_decap_8 FILLER_36_980 ();
 sg13g2_decap_8 FILLER_36_987 ();
 sg13g2_decap_8 FILLER_36_994 ();
 sg13g2_decap_8 FILLER_36_1001 ();
 sg13g2_decap_8 FILLER_36_1008 ();
 sg13g2_decap_8 FILLER_36_1015 ();
 sg13g2_decap_8 FILLER_36_1022 ();
 sg13g2_decap_8 FILLER_36_1029 ();
 sg13g2_decap_8 FILLER_36_1036 ();
 sg13g2_decap_8 FILLER_36_1043 ();
 sg13g2_decap_8 FILLER_36_1050 ();
 sg13g2_decap_8 FILLER_36_1057 ();
 sg13g2_decap_8 FILLER_36_1064 ();
 sg13g2_decap_8 FILLER_36_1071 ();
 sg13g2_decap_8 FILLER_36_1078 ();
 sg13g2_decap_8 FILLER_36_1085 ();
 sg13g2_decap_8 FILLER_36_1092 ();
 sg13g2_decap_8 FILLER_36_1099 ();
 sg13g2_decap_8 FILLER_36_1106 ();
 sg13g2_decap_8 FILLER_36_1113 ();
 sg13g2_decap_8 FILLER_36_1120 ();
 sg13g2_decap_8 FILLER_36_1127 ();
 sg13g2_decap_8 FILLER_36_1134 ();
 sg13g2_decap_8 FILLER_36_1141 ();
 sg13g2_decap_8 FILLER_36_1148 ();
 sg13g2_decap_8 FILLER_36_1155 ();
 sg13g2_decap_8 FILLER_36_1162 ();
 sg13g2_decap_8 FILLER_36_1169 ();
 sg13g2_decap_8 FILLER_36_1176 ();
 sg13g2_decap_8 FILLER_36_1183 ();
 sg13g2_decap_8 FILLER_36_1190 ();
 sg13g2_decap_8 FILLER_36_1197 ();
 sg13g2_decap_8 FILLER_36_1204 ();
 sg13g2_decap_8 FILLER_36_1211 ();
 sg13g2_decap_8 FILLER_36_1218 ();
 sg13g2_decap_8 FILLER_36_1225 ();
 sg13g2_decap_8 FILLER_36_1232 ();
 sg13g2_decap_8 FILLER_36_1239 ();
 sg13g2_decap_8 FILLER_36_1246 ();
 sg13g2_decap_8 FILLER_36_1253 ();
 sg13g2_decap_8 FILLER_36_1260 ();
 sg13g2_decap_8 FILLER_36_1267 ();
 sg13g2_decap_8 FILLER_36_1274 ();
 sg13g2_decap_8 FILLER_36_1281 ();
 sg13g2_decap_8 FILLER_36_1288 ();
 sg13g2_decap_8 FILLER_36_1295 ();
 sg13g2_decap_8 FILLER_36_1302 ();
 sg13g2_decap_8 FILLER_36_1309 ();
 sg13g2_decap_8 FILLER_36_1316 ();
 sg13g2_decap_8 FILLER_36_1323 ();
 sg13g2_decap_8 FILLER_36_1330 ();
 sg13g2_decap_8 FILLER_36_1337 ();
 sg13g2_decap_8 FILLER_36_1344 ();
 sg13g2_decap_8 FILLER_36_1351 ();
 sg13g2_decap_8 FILLER_36_1358 ();
 sg13g2_decap_8 FILLER_36_1365 ();
 sg13g2_decap_8 FILLER_36_1372 ();
 sg13g2_decap_8 FILLER_36_1379 ();
 sg13g2_decap_8 FILLER_36_1386 ();
 sg13g2_decap_8 FILLER_36_1393 ();
 sg13g2_decap_8 FILLER_36_1400 ();
 sg13g2_decap_8 FILLER_36_1407 ();
 sg13g2_decap_8 FILLER_36_1414 ();
 sg13g2_decap_8 FILLER_36_1421 ();
 sg13g2_decap_8 FILLER_36_1428 ();
 sg13g2_decap_8 FILLER_36_1435 ();
 sg13g2_decap_8 FILLER_36_1442 ();
 sg13g2_decap_8 FILLER_36_1449 ();
 sg13g2_decap_8 FILLER_36_1456 ();
 sg13g2_decap_8 FILLER_36_1463 ();
 sg13g2_decap_8 FILLER_36_1470 ();
 sg13g2_decap_8 FILLER_36_1477 ();
 sg13g2_decap_8 FILLER_36_1484 ();
 sg13g2_decap_8 FILLER_36_1491 ();
 sg13g2_decap_8 FILLER_36_1498 ();
 sg13g2_decap_8 FILLER_36_1505 ();
 sg13g2_decap_8 FILLER_36_1512 ();
 sg13g2_decap_8 FILLER_36_1519 ();
 sg13g2_decap_8 FILLER_36_1526 ();
 sg13g2_decap_8 FILLER_36_1533 ();
 sg13g2_decap_8 FILLER_36_1540 ();
 sg13g2_decap_8 FILLER_36_1547 ();
 sg13g2_decap_8 FILLER_36_1554 ();
 sg13g2_decap_8 FILLER_36_1561 ();
 sg13g2_decap_8 FILLER_36_1568 ();
 sg13g2_decap_8 FILLER_36_1575 ();
 sg13g2_decap_8 FILLER_36_1582 ();
 sg13g2_decap_8 FILLER_36_1589 ();
 sg13g2_decap_8 FILLER_36_1596 ();
 sg13g2_decap_8 FILLER_36_1603 ();
 sg13g2_decap_8 FILLER_36_1610 ();
 sg13g2_decap_8 FILLER_36_1617 ();
 sg13g2_decap_8 FILLER_36_1624 ();
 sg13g2_decap_8 FILLER_36_1631 ();
 sg13g2_decap_8 FILLER_36_1638 ();
 sg13g2_decap_8 FILLER_36_1645 ();
 sg13g2_decap_8 FILLER_36_1652 ();
 sg13g2_decap_8 FILLER_36_1659 ();
 sg13g2_decap_8 FILLER_36_1666 ();
 sg13g2_decap_8 FILLER_36_1673 ();
 sg13g2_decap_8 FILLER_36_1680 ();
 sg13g2_decap_8 FILLER_36_1687 ();
 sg13g2_decap_8 FILLER_36_1694 ();
 sg13g2_decap_8 FILLER_36_1701 ();
 sg13g2_decap_8 FILLER_36_1708 ();
 sg13g2_decap_8 FILLER_36_1715 ();
 sg13g2_decap_8 FILLER_36_1722 ();
 sg13g2_decap_8 FILLER_36_1729 ();
 sg13g2_decap_8 FILLER_36_1736 ();
 sg13g2_decap_8 FILLER_36_1743 ();
 sg13g2_decap_8 FILLER_36_1750 ();
 sg13g2_decap_8 FILLER_36_1757 ();
 sg13g2_decap_8 FILLER_36_1764 ();
 sg13g2_decap_8 FILLER_36_1771 ();
 sg13g2_decap_8 FILLER_36_1778 ();
 sg13g2_decap_8 FILLER_36_1785 ();
 sg13g2_decap_8 FILLER_36_1792 ();
 sg13g2_decap_8 FILLER_36_1799 ();
 sg13g2_decap_8 FILLER_36_1806 ();
 sg13g2_decap_8 FILLER_36_1813 ();
 sg13g2_decap_8 FILLER_36_1820 ();
 sg13g2_decap_8 FILLER_36_1827 ();
 sg13g2_decap_8 FILLER_36_1834 ();
 sg13g2_decap_8 FILLER_36_1841 ();
 sg13g2_decap_8 FILLER_36_1848 ();
 sg13g2_decap_8 FILLER_36_1855 ();
 sg13g2_decap_8 FILLER_36_1862 ();
 sg13g2_decap_8 FILLER_36_1869 ();
 sg13g2_decap_8 FILLER_36_1876 ();
 sg13g2_decap_8 FILLER_36_1883 ();
 sg13g2_decap_8 FILLER_36_1890 ();
 sg13g2_decap_8 FILLER_36_1897 ();
 sg13g2_decap_8 FILLER_36_1904 ();
 sg13g2_decap_8 FILLER_36_1911 ();
 sg13g2_decap_8 FILLER_36_1918 ();
 sg13g2_decap_8 FILLER_36_1925 ();
 sg13g2_decap_8 FILLER_36_1932 ();
 sg13g2_decap_8 FILLER_36_1939 ();
 sg13g2_decap_8 FILLER_36_1946 ();
 sg13g2_decap_8 FILLER_36_1953 ();
 sg13g2_decap_8 FILLER_36_1960 ();
 sg13g2_decap_8 FILLER_36_1967 ();
 sg13g2_decap_8 FILLER_36_1974 ();
 sg13g2_decap_8 FILLER_36_1981 ();
 sg13g2_decap_8 FILLER_36_1988 ();
 sg13g2_decap_8 FILLER_36_1995 ();
 sg13g2_decap_8 FILLER_36_2002 ();
 sg13g2_decap_8 FILLER_36_2009 ();
 sg13g2_decap_8 FILLER_36_2016 ();
 sg13g2_decap_8 FILLER_36_2023 ();
 sg13g2_decap_8 FILLER_36_2030 ();
 sg13g2_decap_8 FILLER_36_2037 ();
 sg13g2_decap_8 FILLER_36_2044 ();
 sg13g2_decap_8 FILLER_36_2051 ();
 sg13g2_decap_8 FILLER_36_2058 ();
 sg13g2_decap_8 FILLER_36_2065 ();
 sg13g2_decap_8 FILLER_36_2072 ();
 sg13g2_decap_8 FILLER_36_2079 ();
 sg13g2_decap_8 FILLER_36_2086 ();
 sg13g2_decap_8 FILLER_36_2093 ();
 sg13g2_decap_8 FILLER_36_2100 ();
 sg13g2_decap_8 FILLER_36_2107 ();
 sg13g2_decap_8 FILLER_36_2114 ();
 sg13g2_decap_8 FILLER_36_2121 ();
 sg13g2_decap_8 FILLER_36_2128 ();
 sg13g2_decap_8 FILLER_36_2135 ();
 sg13g2_decap_8 FILLER_36_2142 ();
 sg13g2_decap_8 FILLER_36_2149 ();
 sg13g2_decap_8 FILLER_36_2156 ();
 sg13g2_decap_8 FILLER_36_2163 ();
 sg13g2_decap_8 FILLER_36_2170 ();
 sg13g2_decap_8 FILLER_36_2177 ();
 sg13g2_decap_8 FILLER_36_2184 ();
 sg13g2_decap_8 FILLER_36_2191 ();
 sg13g2_decap_8 FILLER_36_2198 ();
 sg13g2_decap_8 FILLER_36_2205 ();
 sg13g2_decap_8 FILLER_36_2212 ();
 sg13g2_decap_8 FILLER_36_2219 ();
 sg13g2_decap_8 FILLER_36_2226 ();
 sg13g2_decap_8 FILLER_36_2233 ();
 sg13g2_decap_8 FILLER_36_2240 ();
 sg13g2_decap_8 FILLER_36_2247 ();
 sg13g2_decap_8 FILLER_36_2254 ();
 sg13g2_decap_8 FILLER_36_2261 ();
 sg13g2_decap_8 FILLER_36_2268 ();
 sg13g2_decap_8 FILLER_36_2275 ();
 sg13g2_decap_8 FILLER_36_2282 ();
 sg13g2_decap_8 FILLER_36_2289 ();
 sg13g2_decap_8 FILLER_36_2296 ();
 sg13g2_decap_8 FILLER_36_2303 ();
 sg13g2_decap_8 FILLER_36_2310 ();
 sg13g2_decap_8 FILLER_36_2317 ();
 sg13g2_decap_8 FILLER_36_2324 ();
 sg13g2_decap_8 FILLER_36_2331 ();
 sg13g2_decap_8 FILLER_36_2338 ();
 sg13g2_decap_8 FILLER_36_2345 ();
 sg13g2_decap_8 FILLER_36_2352 ();
 sg13g2_decap_8 FILLER_36_2359 ();
 sg13g2_decap_8 FILLER_36_2366 ();
 sg13g2_decap_8 FILLER_36_2373 ();
 sg13g2_decap_8 FILLER_36_2380 ();
 sg13g2_decap_8 FILLER_36_2387 ();
 sg13g2_decap_8 FILLER_36_2394 ();
 sg13g2_decap_8 FILLER_36_2401 ();
 sg13g2_decap_8 FILLER_36_2408 ();
 sg13g2_decap_8 FILLER_36_2415 ();
 sg13g2_decap_8 FILLER_36_2422 ();
 sg13g2_decap_8 FILLER_36_2429 ();
 sg13g2_decap_8 FILLER_36_2436 ();
 sg13g2_decap_8 FILLER_36_2443 ();
 sg13g2_decap_8 FILLER_36_2450 ();
 sg13g2_decap_8 FILLER_36_2457 ();
 sg13g2_decap_8 FILLER_36_2464 ();
 sg13g2_decap_8 FILLER_36_2471 ();
 sg13g2_decap_8 FILLER_36_2478 ();
 sg13g2_decap_8 FILLER_36_2485 ();
 sg13g2_decap_8 FILLER_36_2492 ();
 sg13g2_decap_8 FILLER_36_2499 ();
 sg13g2_decap_8 FILLER_36_2506 ();
 sg13g2_decap_8 FILLER_36_2513 ();
 sg13g2_decap_8 FILLER_36_2520 ();
 sg13g2_decap_8 FILLER_36_2527 ();
 sg13g2_decap_8 FILLER_36_2534 ();
 sg13g2_decap_8 FILLER_36_2541 ();
 sg13g2_decap_8 FILLER_36_2548 ();
 sg13g2_decap_8 FILLER_36_2555 ();
 sg13g2_decap_8 FILLER_36_2562 ();
 sg13g2_decap_8 FILLER_36_2569 ();
 sg13g2_decap_8 FILLER_36_2576 ();
 sg13g2_decap_8 FILLER_36_2583 ();
 sg13g2_decap_8 FILLER_36_2590 ();
 sg13g2_decap_8 FILLER_36_2597 ();
 sg13g2_decap_8 FILLER_36_2604 ();
 sg13g2_decap_8 FILLER_36_2611 ();
 sg13g2_decap_8 FILLER_36_2618 ();
 sg13g2_decap_8 FILLER_36_2625 ();
 sg13g2_decap_8 FILLER_36_2632 ();
 sg13g2_decap_8 FILLER_36_2639 ();
 sg13g2_decap_8 FILLER_36_2646 ();
 sg13g2_decap_8 FILLER_36_2653 ();
 sg13g2_decap_8 FILLER_36_2660 ();
 sg13g2_decap_8 FILLER_36_2667 ();
 sg13g2_decap_8 FILLER_36_2674 ();
 sg13g2_decap_8 FILLER_36_2681 ();
 sg13g2_decap_8 FILLER_36_2688 ();
 sg13g2_decap_8 FILLER_36_2695 ();
 sg13g2_decap_8 FILLER_36_2702 ();
 sg13g2_decap_8 FILLER_36_2709 ();
 sg13g2_decap_8 FILLER_36_2716 ();
 sg13g2_decap_8 FILLER_36_2723 ();
 sg13g2_decap_8 FILLER_36_2730 ();
 sg13g2_decap_8 FILLER_36_2737 ();
 sg13g2_decap_8 FILLER_36_2744 ();
 sg13g2_decap_8 FILLER_36_2751 ();
 sg13g2_decap_8 FILLER_36_2758 ();
 sg13g2_decap_8 FILLER_36_2765 ();
 sg13g2_decap_8 FILLER_36_2772 ();
 sg13g2_decap_8 FILLER_36_2779 ();
 sg13g2_decap_8 FILLER_36_2786 ();
 sg13g2_decap_8 FILLER_36_2793 ();
 sg13g2_decap_8 FILLER_36_2800 ();
 sg13g2_decap_8 FILLER_36_2807 ();
 sg13g2_decap_8 FILLER_36_2814 ();
 sg13g2_decap_8 FILLER_36_2821 ();
 sg13g2_decap_8 FILLER_36_2828 ();
 sg13g2_decap_8 FILLER_36_2835 ();
 sg13g2_decap_8 FILLER_36_2842 ();
 sg13g2_decap_8 FILLER_36_2849 ();
 sg13g2_decap_8 FILLER_36_2856 ();
 sg13g2_decap_8 FILLER_36_2863 ();
 sg13g2_decap_8 FILLER_36_2870 ();
 sg13g2_decap_8 FILLER_36_2877 ();
 sg13g2_decap_8 FILLER_36_2884 ();
 sg13g2_decap_8 FILLER_36_2891 ();
 sg13g2_decap_8 FILLER_36_2898 ();
 sg13g2_decap_8 FILLER_36_2905 ();
 sg13g2_decap_8 FILLER_36_2912 ();
 sg13g2_decap_8 FILLER_36_2919 ();
 sg13g2_decap_8 FILLER_36_2926 ();
 sg13g2_decap_8 FILLER_36_2933 ();
 sg13g2_decap_8 FILLER_36_2940 ();
 sg13g2_decap_8 FILLER_36_2947 ();
 sg13g2_decap_8 FILLER_36_2954 ();
 sg13g2_decap_8 FILLER_36_2961 ();
 sg13g2_decap_8 FILLER_36_2968 ();
 sg13g2_decap_8 FILLER_36_2975 ();
 sg13g2_decap_8 FILLER_36_2982 ();
 sg13g2_decap_8 FILLER_36_2989 ();
 sg13g2_decap_8 FILLER_36_2996 ();
 sg13g2_decap_8 FILLER_36_3003 ();
 sg13g2_decap_8 FILLER_36_3010 ();
 sg13g2_decap_8 FILLER_36_3017 ();
 sg13g2_decap_8 FILLER_36_3024 ();
 sg13g2_decap_8 FILLER_36_3031 ();
 sg13g2_decap_8 FILLER_36_3038 ();
 sg13g2_decap_8 FILLER_36_3045 ();
 sg13g2_decap_8 FILLER_36_3052 ();
 sg13g2_decap_8 FILLER_36_3059 ();
 sg13g2_decap_8 FILLER_36_3066 ();
 sg13g2_decap_8 FILLER_36_3073 ();
 sg13g2_decap_8 FILLER_36_3080 ();
 sg13g2_decap_8 FILLER_36_3087 ();
 sg13g2_decap_8 FILLER_36_3094 ();
 sg13g2_decap_8 FILLER_36_3101 ();
 sg13g2_decap_8 FILLER_36_3108 ();
 sg13g2_decap_8 FILLER_36_3115 ();
 sg13g2_decap_8 FILLER_36_3122 ();
 sg13g2_decap_8 FILLER_36_3129 ();
 sg13g2_decap_8 FILLER_36_3136 ();
 sg13g2_decap_8 FILLER_36_3143 ();
 sg13g2_decap_8 FILLER_36_3150 ();
 sg13g2_decap_8 FILLER_36_3157 ();
 sg13g2_decap_8 FILLER_36_3164 ();
 sg13g2_decap_8 FILLER_36_3171 ();
 sg13g2_decap_8 FILLER_36_3178 ();
 sg13g2_decap_8 FILLER_36_3185 ();
 sg13g2_decap_8 FILLER_36_3192 ();
 sg13g2_decap_8 FILLER_36_3199 ();
 sg13g2_decap_8 FILLER_36_3206 ();
 sg13g2_decap_8 FILLER_36_3213 ();
 sg13g2_decap_8 FILLER_36_3220 ();
 sg13g2_decap_8 FILLER_36_3227 ();
 sg13g2_decap_8 FILLER_36_3234 ();
 sg13g2_decap_8 FILLER_36_3241 ();
 sg13g2_decap_8 FILLER_36_3248 ();
 sg13g2_decap_8 FILLER_36_3255 ();
 sg13g2_decap_8 FILLER_36_3262 ();
 sg13g2_decap_8 FILLER_36_3269 ();
 sg13g2_decap_8 FILLER_36_3276 ();
 sg13g2_decap_8 FILLER_36_3283 ();
 sg13g2_decap_8 FILLER_36_3290 ();
 sg13g2_decap_8 FILLER_36_3297 ();
 sg13g2_decap_8 FILLER_36_3304 ();
 sg13g2_decap_8 FILLER_36_3311 ();
 sg13g2_decap_8 FILLER_36_3318 ();
 sg13g2_decap_8 FILLER_36_3325 ();
 sg13g2_decap_8 FILLER_36_3332 ();
 sg13g2_decap_8 FILLER_36_3339 ();
 sg13g2_decap_8 FILLER_36_3346 ();
 sg13g2_decap_8 FILLER_36_3353 ();
 sg13g2_decap_8 FILLER_36_3360 ();
 sg13g2_decap_8 FILLER_36_3367 ();
 sg13g2_decap_8 FILLER_36_3374 ();
 sg13g2_decap_8 FILLER_36_3381 ();
 sg13g2_decap_8 FILLER_36_3388 ();
 sg13g2_decap_8 FILLER_36_3395 ();
 sg13g2_decap_8 FILLER_36_3402 ();
 sg13g2_decap_8 FILLER_36_3409 ();
 sg13g2_decap_8 FILLER_36_3416 ();
 sg13g2_decap_8 FILLER_36_3423 ();
 sg13g2_decap_8 FILLER_36_3430 ();
 sg13g2_decap_8 FILLER_36_3437 ();
 sg13g2_decap_8 FILLER_36_3444 ();
 sg13g2_decap_8 FILLER_36_3451 ();
 sg13g2_decap_8 FILLER_36_3458 ();
 sg13g2_decap_8 FILLER_36_3465 ();
 sg13g2_decap_8 FILLER_36_3472 ();
 sg13g2_decap_8 FILLER_36_3479 ();
 sg13g2_decap_8 FILLER_36_3486 ();
 sg13g2_decap_8 FILLER_36_3493 ();
 sg13g2_decap_8 FILLER_36_3500 ();
 sg13g2_decap_8 FILLER_36_3507 ();
 sg13g2_decap_8 FILLER_36_3514 ();
 sg13g2_decap_8 FILLER_36_3521 ();
 sg13g2_decap_8 FILLER_36_3528 ();
 sg13g2_decap_8 FILLER_36_3535 ();
 sg13g2_decap_8 FILLER_36_3542 ();
 sg13g2_decap_8 FILLER_36_3549 ();
 sg13g2_decap_8 FILLER_36_3556 ();
 sg13g2_decap_8 FILLER_36_3563 ();
 sg13g2_decap_8 FILLER_36_3570 ();
 sg13g2_fill_2 FILLER_36_3577 ();
 sg13g2_fill_1 FILLER_36_3579 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_245 ();
 sg13g2_decap_8 FILLER_37_252 ();
 sg13g2_decap_8 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_decap_8 FILLER_37_294 ();
 sg13g2_decap_8 FILLER_37_301 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_37_315 ();
 sg13g2_decap_8 FILLER_37_322 ();
 sg13g2_decap_8 FILLER_37_329 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_decap_8 FILLER_37_406 ();
 sg13g2_decap_8 FILLER_37_413 ();
 sg13g2_decap_8 FILLER_37_420 ();
 sg13g2_decap_8 FILLER_37_427 ();
 sg13g2_decap_8 FILLER_37_434 ();
 sg13g2_decap_8 FILLER_37_441 ();
 sg13g2_decap_8 FILLER_37_448 ();
 sg13g2_decap_8 FILLER_37_455 ();
 sg13g2_decap_8 FILLER_37_462 ();
 sg13g2_decap_8 FILLER_37_469 ();
 sg13g2_decap_8 FILLER_37_476 ();
 sg13g2_decap_8 FILLER_37_483 ();
 sg13g2_decap_8 FILLER_37_490 ();
 sg13g2_decap_8 FILLER_37_497 ();
 sg13g2_decap_8 FILLER_37_504 ();
 sg13g2_decap_8 FILLER_37_511 ();
 sg13g2_decap_8 FILLER_37_518 ();
 sg13g2_decap_8 FILLER_37_525 ();
 sg13g2_decap_8 FILLER_37_532 ();
 sg13g2_decap_8 FILLER_37_539 ();
 sg13g2_decap_8 FILLER_37_546 ();
 sg13g2_decap_8 FILLER_37_553 ();
 sg13g2_decap_8 FILLER_37_560 ();
 sg13g2_decap_8 FILLER_37_567 ();
 sg13g2_decap_8 FILLER_37_574 ();
 sg13g2_decap_8 FILLER_37_581 ();
 sg13g2_decap_8 FILLER_37_588 ();
 sg13g2_decap_8 FILLER_37_595 ();
 sg13g2_decap_8 FILLER_37_602 ();
 sg13g2_decap_8 FILLER_37_609 ();
 sg13g2_decap_8 FILLER_37_616 ();
 sg13g2_decap_8 FILLER_37_623 ();
 sg13g2_decap_8 FILLER_37_630 ();
 sg13g2_decap_8 FILLER_37_637 ();
 sg13g2_decap_8 FILLER_37_644 ();
 sg13g2_decap_8 FILLER_37_651 ();
 sg13g2_decap_8 FILLER_37_658 ();
 sg13g2_decap_8 FILLER_37_665 ();
 sg13g2_decap_8 FILLER_37_672 ();
 sg13g2_decap_8 FILLER_37_679 ();
 sg13g2_decap_8 FILLER_37_686 ();
 sg13g2_decap_8 FILLER_37_693 ();
 sg13g2_decap_8 FILLER_37_700 ();
 sg13g2_decap_8 FILLER_37_707 ();
 sg13g2_decap_8 FILLER_37_714 ();
 sg13g2_decap_8 FILLER_37_721 ();
 sg13g2_decap_8 FILLER_37_728 ();
 sg13g2_decap_8 FILLER_37_735 ();
 sg13g2_decap_8 FILLER_37_742 ();
 sg13g2_decap_8 FILLER_37_749 ();
 sg13g2_decap_8 FILLER_37_756 ();
 sg13g2_decap_8 FILLER_37_763 ();
 sg13g2_decap_8 FILLER_37_770 ();
 sg13g2_decap_8 FILLER_37_777 ();
 sg13g2_decap_8 FILLER_37_784 ();
 sg13g2_decap_8 FILLER_37_791 ();
 sg13g2_decap_8 FILLER_37_798 ();
 sg13g2_decap_8 FILLER_37_805 ();
 sg13g2_decap_8 FILLER_37_812 ();
 sg13g2_decap_8 FILLER_37_819 ();
 sg13g2_decap_8 FILLER_37_826 ();
 sg13g2_decap_8 FILLER_37_833 ();
 sg13g2_decap_8 FILLER_37_840 ();
 sg13g2_decap_8 FILLER_37_847 ();
 sg13g2_decap_8 FILLER_37_854 ();
 sg13g2_decap_8 FILLER_37_861 ();
 sg13g2_decap_8 FILLER_37_868 ();
 sg13g2_decap_8 FILLER_37_875 ();
 sg13g2_decap_8 FILLER_37_882 ();
 sg13g2_decap_8 FILLER_37_889 ();
 sg13g2_decap_8 FILLER_37_896 ();
 sg13g2_decap_8 FILLER_37_903 ();
 sg13g2_decap_8 FILLER_37_910 ();
 sg13g2_decap_8 FILLER_37_917 ();
 sg13g2_decap_8 FILLER_37_924 ();
 sg13g2_decap_8 FILLER_37_931 ();
 sg13g2_decap_8 FILLER_37_938 ();
 sg13g2_decap_8 FILLER_37_945 ();
 sg13g2_decap_8 FILLER_37_952 ();
 sg13g2_decap_8 FILLER_37_959 ();
 sg13g2_decap_8 FILLER_37_966 ();
 sg13g2_decap_8 FILLER_37_973 ();
 sg13g2_decap_8 FILLER_37_980 ();
 sg13g2_decap_8 FILLER_37_987 ();
 sg13g2_decap_8 FILLER_37_994 ();
 sg13g2_decap_8 FILLER_37_1001 ();
 sg13g2_decap_8 FILLER_37_1008 ();
 sg13g2_decap_8 FILLER_37_1015 ();
 sg13g2_decap_8 FILLER_37_1022 ();
 sg13g2_decap_8 FILLER_37_1029 ();
 sg13g2_decap_8 FILLER_37_1036 ();
 sg13g2_decap_8 FILLER_37_1043 ();
 sg13g2_decap_8 FILLER_37_1050 ();
 sg13g2_decap_8 FILLER_37_1057 ();
 sg13g2_decap_8 FILLER_37_1064 ();
 sg13g2_decap_8 FILLER_37_1071 ();
 sg13g2_decap_8 FILLER_37_1078 ();
 sg13g2_decap_8 FILLER_37_1085 ();
 sg13g2_decap_8 FILLER_37_1092 ();
 sg13g2_decap_8 FILLER_37_1099 ();
 sg13g2_decap_8 FILLER_37_1106 ();
 sg13g2_decap_8 FILLER_37_1113 ();
 sg13g2_decap_8 FILLER_37_1120 ();
 sg13g2_decap_8 FILLER_37_1127 ();
 sg13g2_decap_8 FILLER_37_1134 ();
 sg13g2_decap_8 FILLER_37_1141 ();
 sg13g2_decap_8 FILLER_37_1148 ();
 sg13g2_decap_8 FILLER_37_1155 ();
 sg13g2_decap_8 FILLER_37_1162 ();
 sg13g2_decap_8 FILLER_37_1169 ();
 sg13g2_decap_8 FILLER_37_1176 ();
 sg13g2_decap_8 FILLER_37_1183 ();
 sg13g2_decap_8 FILLER_37_1190 ();
 sg13g2_decap_8 FILLER_37_1197 ();
 sg13g2_decap_8 FILLER_37_1204 ();
 sg13g2_decap_8 FILLER_37_1211 ();
 sg13g2_decap_8 FILLER_37_1218 ();
 sg13g2_decap_8 FILLER_37_1225 ();
 sg13g2_decap_8 FILLER_37_1232 ();
 sg13g2_decap_8 FILLER_37_1239 ();
 sg13g2_decap_8 FILLER_37_1246 ();
 sg13g2_decap_8 FILLER_37_1253 ();
 sg13g2_decap_8 FILLER_37_1260 ();
 sg13g2_decap_8 FILLER_37_1267 ();
 sg13g2_decap_8 FILLER_37_1274 ();
 sg13g2_decap_8 FILLER_37_1281 ();
 sg13g2_decap_8 FILLER_37_1288 ();
 sg13g2_decap_8 FILLER_37_1295 ();
 sg13g2_decap_8 FILLER_37_1302 ();
 sg13g2_decap_8 FILLER_37_1309 ();
 sg13g2_decap_8 FILLER_37_1316 ();
 sg13g2_decap_8 FILLER_37_1323 ();
 sg13g2_decap_8 FILLER_37_1330 ();
 sg13g2_decap_8 FILLER_37_1337 ();
 sg13g2_decap_8 FILLER_37_1344 ();
 sg13g2_decap_8 FILLER_37_1351 ();
 sg13g2_decap_8 FILLER_37_1358 ();
 sg13g2_decap_8 FILLER_37_1365 ();
 sg13g2_decap_8 FILLER_37_1372 ();
 sg13g2_decap_8 FILLER_37_1379 ();
 sg13g2_decap_8 FILLER_37_1386 ();
 sg13g2_decap_8 FILLER_37_1393 ();
 sg13g2_decap_8 FILLER_37_1400 ();
 sg13g2_decap_8 FILLER_37_1407 ();
 sg13g2_decap_8 FILLER_37_1414 ();
 sg13g2_decap_8 FILLER_37_1421 ();
 sg13g2_decap_8 FILLER_37_1428 ();
 sg13g2_decap_8 FILLER_37_1435 ();
 sg13g2_decap_8 FILLER_37_1442 ();
 sg13g2_decap_8 FILLER_37_1449 ();
 sg13g2_decap_8 FILLER_37_1456 ();
 sg13g2_decap_8 FILLER_37_1463 ();
 sg13g2_decap_8 FILLER_37_1470 ();
 sg13g2_decap_8 FILLER_37_1477 ();
 sg13g2_decap_8 FILLER_37_1484 ();
 sg13g2_decap_8 FILLER_37_1491 ();
 sg13g2_decap_8 FILLER_37_1498 ();
 sg13g2_decap_8 FILLER_37_1505 ();
 sg13g2_decap_8 FILLER_37_1512 ();
 sg13g2_decap_8 FILLER_37_1519 ();
 sg13g2_decap_8 FILLER_37_1526 ();
 sg13g2_decap_8 FILLER_37_1533 ();
 sg13g2_decap_8 FILLER_37_1540 ();
 sg13g2_decap_8 FILLER_37_1547 ();
 sg13g2_decap_8 FILLER_37_1554 ();
 sg13g2_decap_8 FILLER_37_1561 ();
 sg13g2_decap_8 FILLER_37_1568 ();
 sg13g2_decap_8 FILLER_37_1575 ();
 sg13g2_decap_8 FILLER_37_1582 ();
 sg13g2_decap_8 FILLER_37_1589 ();
 sg13g2_decap_8 FILLER_37_1596 ();
 sg13g2_decap_8 FILLER_37_1603 ();
 sg13g2_decap_8 FILLER_37_1610 ();
 sg13g2_decap_8 FILLER_37_1617 ();
 sg13g2_decap_8 FILLER_37_1624 ();
 sg13g2_decap_8 FILLER_37_1631 ();
 sg13g2_decap_8 FILLER_37_1638 ();
 sg13g2_decap_8 FILLER_37_1645 ();
 sg13g2_decap_8 FILLER_37_1652 ();
 sg13g2_decap_8 FILLER_37_1659 ();
 sg13g2_decap_8 FILLER_37_1666 ();
 sg13g2_decap_8 FILLER_37_1673 ();
 sg13g2_decap_8 FILLER_37_1680 ();
 sg13g2_decap_8 FILLER_37_1687 ();
 sg13g2_decap_8 FILLER_37_1694 ();
 sg13g2_decap_8 FILLER_37_1701 ();
 sg13g2_decap_8 FILLER_37_1708 ();
 sg13g2_decap_8 FILLER_37_1715 ();
 sg13g2_decap_8 FILLER_37_1722 ();
 sg13g2_decap_8 FILLER_37_1729 ();
 sg13g2_decap_8 FILLER_37_1736 ();
 sg13g2_decap_8 FILLER_37_1743 ();
 sg13g2_decap_8 FILLER_37_1750 ();
 sg13g2_decap_8 FILLER_37_1757 ();
 sg13g2_decap_8 FILLER_37_1764 ();
 sg13g2_decap_8 FILLER_37_1771 ();
 sg13g2_decap_8 FILLER_37_1778 ();
 sg13g2_decap_8 FILLER_37_1785 ();
 sg13g2_decap_8 FILLER_37_1792 ();
 sg13g2_decap_8 FILLER_37_1799 ();
 sg13g2_decap_8 FILLER_37_1806 ();
 sg13g2_decap_8 FILLER_37_1813 ();
 sg13g2_decap_8 FILLER_37_1820 ();
 sg13g2_decap_8 FILLER_37_1827 ();
 sg13g2_decap_8 FILLER_37_1834 ();
 sg13g2_decap_8 FILLER_37_1841 ();
 sg13g2_decap_8 FILLER_37_1848 ();
 sg13g2_decap_8 FILLER_37_1855 ();
 sg13g2_decap_8 FILLER_37_1862 ();
 sg13g2_decap_8 FILLER_37_1869 ();
 sg13g2_decap_8 FILLER_37_1876 ();
 sg13g2_decap_8 FILLER_37_1883 ();
 sg13g2_decap_8 FILLER_37_1890 ();
 sg13g2_decap_8 FILLER_37_1897 ();
 sg13g2_decap_8 FILLER_37_1904 ();
 sg13g2_decap_8 FILLER_37_1911 ();
 sg13g2_decap_8 FILLER_37_1918 ();
 sg13g2_decap_8 FILLER_37_1925 ();
 sg13g2_decap_8 FILLER_37_1932 ();
 sg13g2_decap_8 FILLER_37_1939 ();
 sg13g2_decap_8 FILLER_37_1946 ();
 sg13g2_decap_8 FILLER_37_1953 ();
 sg13g2_decap_8 FILLER_37_1960 ();
 sg13g2_decap_8 FILLER_37_1967 ();
 sg13g2_decap_8 FILLER_37_1974 ();
 sg13g2_decap_8 FILLER_37_1981 ();
 sg13g2_decap_8 FILLER_37_1988 ();
 sg13g2_decap_8 FILLER_37_1995 ();
 sg13g2_decap_8 FILLER_37_2002 ();
 sg13g2_decap_8 FILLER_37_2009 ();
 sg13g2_decap_8 FILLER_37_2016 ();
 sg13g2_decap_8 FILLER_37_2023 ();
 sg13g2_decap_8 FILLER_37_2030 ();
 sg13g2_decap_8 FILLER_37_2037 ();
 sg13g2_decap_8 FILLER_37_2044 ();
 sg13g2_decap_8 FILLER_37_2051 ();
 sg13g2_decap_8 FILLER_37_2058 ();
 sg13g2_decap_8 FILLER_37_2065 ();
 sg13g2_decap_8 FILLER_37_2072 ();
 sg13g2_decap_8 FILLER_37_2079 ();
 sg13g2_decap_8 FILLER_37_2086 ();
 sg13g2_decap_8 FILLER_37_2093 ();
 sg13g2_decap_8 FILLER_37_2100 ();
 sg13g2_decap_8 FILLER_37_2107 ();
 sg13g2_decap_8 FILLER_37_2114 ();
 sg13g2_decap_8 FILLER_37_2121 ();
 sg13g2_decap_8 FILLER_37_2128 ();
 sg13g2_decap_8 FILLER_37_2135 ();
 sg13g2_decap_8 FILLER_37_2142 ();
 sg13g2_decap_8 FILLER_37_2149 ();
 sg13g2_decap_8 FILLER_37_2156 ();
 sg13g2_decap_8 FILLER_37_2163 ();
 sg13g2_decap_8 FILLER_37_2170 ();
 sg13g2_decap_8 FILLER_37_2177 ();
 sg13g2_decap_8 FILLER_37_2184 ();
 sg13g2_decap_8 FILLER_37_2191 ();
 sg13g2_decap_8 FILLER_37_2198 ();
 sg13g2_decap_8 FILLER_37_2205 ();
 sg13g2_decap_8 FILLER_37_2212 ();
 sg13g2_decap_8 FILLER_37_2219 ();
 sg13g2_decap_8 FILLER_37_2226 ();
 sg13g2_decap_8 FILLER_37_2233 ();
 sg13g2_decap_8 FILLER_37_2240 ();
 sg13g2_decap_8 FILLER_37_2247 ();
 sg13g2_decap_8 FILLER_37_2254 ();
 sg13g2_decap_8 FILLER_37_2261 ();
 sg13g2_decap_8 FILLER_37_2268 ();
 sg13g2_decap_8 FILLER_37_2275 ();
 sg13g2_decap_8 FILLER_37_2282 ();
 sg13g2_decap_8 FILLER_37_2289 ();
 sg13g2_decap_8 FILLER_37_2296 ();
 sg13g2_decap_8 FILLER_37_2303 ();
 sg13g2_decap_8 FILLER_37_2310 ();
 sg13g2_decap_8 FILLER_37_2317 ();
 sg13g2_decap_8 FILLER_37_2324 ();
 sg13g2_decap_8 FILLER_37_2331 ();
 sg13g2_decap_8 FILLER_37_2338 ();
 sg13g2_decap_8 FILLER_37_2345 ();
 sg13g2_decap_8 FILLER_37_2352 ();
 sg13g2_decap_8 FILLER_37_2359 ();
 sg13g2_decap_8 FILLER_37_2366 ();
 sg13g2_decap_8 FILLER_37_2373 ();
 sg13g2_decap_8 FILLER_37_2380 ();
 sg13g2_decap_8 FILLER_37_2387 ();
 sg13g2_decap_8 FILLER_37_2394 ();
 sg13g2_decap_8 FILLER_37_2401 ();
 sg13g2_decap_8 FILLER_37_2408 ();
 sg13g2_decap_8 FILLER_37_2415 ();
 sg13g2_decap_8 FILLER_37_2422 ();
 sg13g2_decap_8 FILLER_37_2429 ();
 sg13g2_decap_8 FILLER_37_2436 ();
 sg13g2_decap_8 FILLER_37_2443 ();
 sg13g2_decap_8 FILLER_37_2450 ();
 sg13g2_decap_8 FILLER_37_2457 ();
 sg13g2_decap_8 FILLER_37_2464 ();
 sg13g2_decap_8 FILLER_37_2471 ();
 sg13g2_decap_8 FILLER_37_2478 ();
 sg13g2_decap_8 FILLER_37_2485 ();
 sg13g2_decap_8 FILLER_37_2492 ();
 sg13g2_decap_8 FILLER_37_2499 ();
 sg13g2_decap_8 FILLER_37_2506 ();
 sg13g2_decap_8 FILLER_37_2513 ();
 sg13g2_decap_8 FILLER_37_2520 ();
 sg13g2_decap_8 FILLER_37_2527 ();
 sg13g2_decap_8 FILLER_37_2534 ();
 sg13g2_decap_8 FILLER_37_2541 ();
 sg13g2_decap_8 FILLER_37_2548 ();
 sg13g2_decap_8 FILLER_37_2555 ();
 sg13g2_decap_8 FILLER_37_2562 ();
 sg13g2_decap_8 FILLER_37_2569 ();
 sg13g2_decap_8 FILLER_37_2576 ();
 sg13g2_decap_8 FILLER_37_2583 ();
 sg13g2_decap_8 FILLER_37_2590 ();
 sg13g2_decap_8 FILLER_37_2597 ();
 sg13g2_decap_8 FILLER_37_2604 ();
 sg13g2_decap_8 FILLER_37_2611 ();
 sg13g2_decap_8 FILLER_37_2618 ();
 sg13g2_decap_8 FILLER_37_2625 ();
 sg13g2_decap_8 FILLER_37_2632 ();
 sg13g2_decap_8 FILLER_37_2639 ();
 sg13g2_decap_8 FILLER_37_2646 ();
 sg13g2_decap_8 FILLER_37_2653 ();
 sg13g2_decap_8 FILLER_37_2660 ();
 sg13g2_decap_8 FILLER_37_2667 ();
 sg13g2_decap_8 FILLER_37_2674 ();
 sg13g2_decap_8 FILLER_37_2681 ();
 sg13g2_decap_8 FILLER_37_2688 ();
 sg13g2_decap_8 FILLER_37_2695 ();
 sg13g2_decap_8 FILLER_37_2702 ();
 sg13g2_decap_8 FILLER_37_2709 ();
 sg13g2_decap_8 FILLER_37_2716 ();
 sg13g2_decap_8 FILLER_37_2723 ();
 sg13g2_decap_8 FILLER_37_2730 ();
 sg13g2_decap_8 FILLER_37_2737 ();
 sg13g2_decap_8 FILLER_37_2744 ();
 sg13g2_decap_8 FILLER_37_2751 ();
 sg13g2_decap_8 FILLER_37_2758 ();
 sg13g2_decap_8 FILLER_37_2765 ();
 sg13g2_decap_8 FILLER_37_2772 ();
 sg13g2_decap_8 FILLER_37_2779 ();
 sg13g2_decap_8 FILLER_37_2786 ();
 sg13g2_decap_8 FILLER_37_2793 ();
 sg13g2_decap_8 FILLER_37_2800 ();
 sg13g2_decap_8 FILLER_37_2807 ();
 sg13g2_decap_8 FILLER_37_2814 ();
 sg13g2_decap_8 FILLER_37_2821 ();
 sg13g2_decap_8 FILLER_37_2828 ();
 sg13g2_decap_8 FILLER_37_2835 ();
 sg13g2_decap_8 FILLER_37_2842 ();
 sg13g2_decap_8 FILLER_37_2849 ();
 sg13g2_decap_8 FILLER_37_2856 ();
 sg13g2_decap_8 FILLER_37_2863 ();
 sg13g2_decap_8 FILLER_37_2870 ();
 sg13g2_decap_8 FILLER_37_2877 ();
 sg13g2_decap_8 FILLER_37_2884 ();
 sg13g2_decap_8 FILLER_37_2891 ();
 sg13g2_decap_8 FILLER_37_2898 ();
 sg13g2_decap_8 FILLER_37_2905 ();
 sg13g2_decap_8 FILLER_37_2912 ();
 sg13g2_decap_8 FILLER_37_2919 ();
 sg13g2_decap_8 FILLER_37_2926 ();
 sg13g2_decap_8 FILLER_37_2933 ();
 sg13g2_decap_8 FILLER_37_2940 ();
 sg13g2_decap_8 FILLER_37_2947 ();
 sg13g2_decap_8 FILLER_37_2954 ();
 sg13g2_decap_8 FILLER_37_2961 ();
 sg13g2_decap_8 FILLER_37_2968 ();
 sg13g2_decap_8 FILLER_37_2975 ();
 sg13g2_decap_8 FILLER_37_2982 ();
 sg13g2_decap_8 FILLER_37_2989 ();
 sg13g2_decap_8 FILLER_37_2996 ();
 sg13g2_decap_8 FILLER_37_3003 ();
 sg13g2_decap_8 FILLER_37_3010 ();
 sg13g2_decap_8 FILLER_37_3017 ();
 sg13g2_decap_8 FILLER_37_3024 ();
 sg13g2_decap_8 FILLER_37_3031 ();
 sg13g2_decap_8 FILLER_37_3038 ();
 sg13g2_decap_8 FILLER_37_3045 ();
 sg13g2_decap_8 FILLER_37_3052 ();
 sg13g2_decap_8 FILLER_37_3059 ();
 sg13g2_decap_8 FILLER_37_3066 ();
 sg13g2_decap_8 FILLER_37_3073 ();
 sg13g2_decap_8 FILLER_37_3080 ();
 sg13g2_decap_8 FILLER_37_3087 ();
 sg13g2_decap_8 FILLER_37_3094 ();
 sg13g2_decap_8 FILLER_37_3101 ();
 sg13g2_decap_8 FILLER_37_3108 ();
 sg13g2_decap_8 FILLER_37_3115 ();
 sg13g2_decap_8 FILLER_37_3122 ();
 sg13g2_decap_8 FILLER_37_3129 ();
 sg13g2_decap_8 FILLER_37_3136 ();
 sg13g2_decap_8 FILLER_37_3143 ();
 sg13g2_decap_8 FILLER_37_3150 ();
 sg13g2_decap_8 FILLER_37_3157 ();
 sg13g2_decap_8 FILLER_37_3164 ();
 sg13g2_decap_8 FILLER_37_3171 ();
 sg13g2_decap_8 FILLER_37_3178 ();
 sg13g2_decap_8 FILLER_37_3185 ();
 sg13g2_decap_8 FILLER_37_3192 ();
 sg13g2_decap_8 FILLER_37_3199 ();
 sg13g2_decap_8 FILLER_37_3206 ();
 sg13g2_decap_8 FILLER_37_3213 ();
 sg13g2_decap_8 FILLER_37_3220 ();
 sg13g2_decap_8 FILLER_37_3227 ();
 sg13g2_decap_8 FILLER_37_3234 ();
 sg13g2_decap_8 FILLER_37_3241 ();
 sg13g2_decap_8 FILLER_37_3248 ();
 sg13g2_decap_8 FILLER_37_3255 ();
 sg13g2_decap_8 FILLER_37_3262 ();
 sg13g2_decap_8 FILLER_37_3269 ();
 sg13g2_decap_8 FILLER_37_3276 ();
 sg13g2_decap_8 FILLER_37_3283 ();
 sg13g2_decap_8 FILLER_37_3290 ();
 sg13g2_decap_8 FILLER_37_3297 ();
 sg13g2_decap_8 FILLER_37_3304 ();
 sg13g2_decap_8 FILLER_37_3311 ();
 sg13g2_decap_8 FILLER_37_3318 ();
 sg13g2_decap_8 FILLER_37_3325 ();
 sg13g2_decap_8 FILLER_37_3332 ();
 sg13g2_decap_8 FILLER_37_3339 ();
 sg13g2_decap_8 FILLER_37_3346 ();
 sg13g2_decap_8 FILLER_37_3353 ();
 sg13g2_decap_8 FILLER_37_3360 ();
 sg13g2_decap_8 FILLER_37_3367 ();
 sg13g2_decap_8 FILLER_37_3374 ();
 sg13g2_decap_8 FILLER_37_3381 ();
 sg13g2_decap_8 FILLER_37_3388 ();
 sg13g2_decap_8 FILLER_37_3395 ();
 sg13g2_decap_8 FILLER_37_3402 ();
 sg13g2_decap_8 FILLER_37_3409 ();
 sg13g2_decap_8 FILLER_37_3416 ();
 sg13g2_decap_8 FILLER_37_3423 ();
 sg13g2_decap_8 FILLER_37_3430 ();
 sg13g2_decap_8 FILLER_37_3437 ();
 sg13g2_decap_8 FILLER_37_3444 ();
 sg13g2_decap_8 FILLER_37_3451 ();
 sg13g2_decap_8 FILLER_37_3458 ();
 sg13g2_decap_8 FILLER_37_3465 ();
 sg13g2_decap_8 FILLER_37_3472 ();
 sg13g2_decap_8 FILLER_37_3479 ();
 sg13g2_decap_8 FILLER_37_3486 ();
 sg13g2_decap_8 FILLER_37_3493 ();
 sg13g2_decap_8 FILLER_37_3500 ();
 sg13g2_decap_8 FILLER_37_3507 ();
 sg13g2_decap_8 FILLER_37_3514 ();
 sg13g2_decap_8 FILLER_37_3521 ();
 sg13g2_decap_8 FILLER_37_3528 ();
 sg13g2_decap_8 FILLER_37_3535 ();
 sg13g2_decap_8 FILLER_37_3542 ();
 sg13g2_decap_8 FILLER_37_3549 ();
 sg13g2_decap_8 FILLER_37_3556 ();
 sg13g2_decap_8 FILLER_37_3563 ();
 sg13g2_decap_8 FILLER_37_3570 ();
 sg13g2_fill_2 FILLER_37_3577 ();
 sg13g2_fill_1 FILLER_37_3579 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_decap_8 FILLER_38_224 ();
 sg13g2_decap_8 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_decap_8 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_252 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_decap_8 FILLER_38_273 ();
 sg13g2_decap_8 FILLER_38_280 ();
 sg13g2_decap_8 FILLER_38_287 ();
 sg13g2_decap_8 FILLER_38_294 ();
 sg13g2_decap_8 FILLER_38_301 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_315 ();
 sg13g2_decap_8 FILLER_38_322 ();
 sg13g2_decap_8 FILLER_38_329 ();
 sg13g2_decap_8 FILLER_38_336 ();
 sg13g2_decap_8 FILLER_38_343 ();
 sg13g2_decap_8 FILLER_38_350 ();
 sg13g2_decap_8 FILLER_38_357 ();
 sg13g2_decap_8 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_371 ();
 sg13g2_decap_8 FILLER_38_378 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_decap_8 FILLER_38_406 ();
 sg13g2_decap_8 FILLER_38_413 ();
 sg13g2_decap_8 FILLER_38_420 ();
 sg13g2_decap_8 FILLER_38_427 ();
 sg13g2_decap_8 FILLER_38_434 ();
 sg13g2_decap_8 FILLER_38_441 ();
 sg13g2_decap_8 FILLER_38_448 ();
 sg13g2_decap_8 FILLER_38_455 ();
 sg13g2_decap_8 FILLER_38_462 ();
 sg13g2_decap_8 FILLER_38_469 ();
 sg13g2_decap_8 FILLER_38_476 ();
 sg13g2_decap_8 FILLER_38_483 ();
 sg13g2_decap_8 FILLER_38_490 ();
 sg13g2_decap_8 FILLER_38_497 ();
 sg13g2_decap_8 FILLER_38_504 ();
 sg13g2_decap_8 FILLER_38_511 ();
 sg13g2_decap_8 FILLER_38_518 ();
 sg13g2_decap_8 FILLER_38_525 ();
 sg13g2_decap_8 FILLER_38_532 ();
 sg13g2_decap_8 FILLER_38_539 ();
 sg13g2_decap_8 FILLER_38_546 ();
 sg13g2_decap_8 FILLER_38_553 ();
 sg13g2_decap_8 FILLER_38_560 ();
 sg13g2_decap_8 FILLER_38_567 ();
 sg13g2_decap_8 FILLER_38_574 ();
 sg13g2_decap_8 FILLER_38_581 ();
 sg13g2_decap_8 FILLER_38_588 ();
 sg13g2_decap_8 FILLER_38_595 ();
 sg13g2_decap_8 FILLER_38_602 ();
 sg13g2_decap_8 FILLER_38_609 ();
 sg13g2_decap_8 FILLER_38_616 ();
 sg13g2_decap_8 FILLER_38_623 ();
 sg13g2_decap_8 FILLER_38_630 ();
 sg13g2_decap_8 FILLER_38_637 ();
 sg13g2_decap_8 FILLER_38_644 ();
 sg13g2_decap_8 FILLER_38_651 ();
 sg13g2_decap_8 FILLER_38_658 ();
 sg13g2_decap_8 FILLER_38_665 ();
 sg13g2_decap_8 FILLER_38_672 ();
 sg13g2_decap_8 FILLER_38_679 ();
 sg13g2_decap_8 FILLER_38_686 ();
 sg13g2_decap_8 FILLER_38_693 ();
 sg13g2_decap_8 FILLER_38_700 ();
 sg13g2_decap_8 FILLER_38_707 ();
 sg13g2_decap_8 FILLER_38_714 ();
 sg13g2_decap_8 FILLER_38_721 ();
 sg13g2_decap_8 FILLER_38_728 ();
 sg13g2_decap_8 FILLER_38_735 ();
 sg13g2_decap_8 FILLER_38_742 ();
 sg13g2_decap_8 FILLER_38_749 ();
 sg13g2_decap_8 FILLER_38_756 ();
 sg13g2_decap_8 FILLER_38_763 ();
 sg13g2_decap_8 FILLER_38_770 ();
 sg13g2_decap_8 FILLER_38_777 ();
 sg13g2_decap_8 FILLER_38_784 ();
 sg13g2_decap_8 FILLER_38_791 ();
 sg13g2_decap_8 FILLER_38_798 ();
 sg13g2_decap_8 FILLER_38_805 ();
 sg13g2_decap_8 FILLER_38_812 ();
 sg13g2_decap_8 FILLER_38_819 ();
 sg13g2_decap_8 FILLER_38_826 ();
 sg13g2_decap_8 FILLER_38_833 ();
 sg13g2_decap_8 FILLER_38_840 ();
 sg13g2_decap_8 FILLER_38_847 ();
 sg13g2_decap_8 FILLER_38_854 ();
 sg13g2_decap_8 FILLER_38_861 ();
 sg13g2_decap_8 FILLER_38_868 ();
 sg13g2_decap_8 FILLER_38_875 ();
 sg13g2_decap_8 FILLER_38_882 ();
 sg13g2_decap_8 FILLER_38_889 ();
 sg13g2_decap_8 FILLER_38_896 ();
 sg13g2_decap_8 FILLER_38_903 ();
 sg13g2_decap_8 FILLER_38_910 ();
 sg13g2_decap_8 FILLER_38_917 ();
 sg13g2_decap_8 FILLER_38_924 ();
 sg13g2_decap_8 FILLER_38_931 ();
 sg13g2_decap_8 FILLER_38_938 ();
 sg13g2_decap_8 FILLER_38_945 ();
 sg13g2_decap_8 FILLER_38_952 ();
 sg13g2_decap_8 FILLER_38_959 ();
 sg13g2_decap_8 FILLER_38_966 ();
 sg13g2_decap_8 FILLER_38_973 ();
 sg13g2_decap_8 FILLER_38_980 ();
 sg13g2_decap_8 FILLER_38_987 ();
 sg13g2_decap_8 FILLER_38_994 ();
 sg13g2_decap_8 FILLER_38_1001 ();
 sg13g2_decap_8 FILLER_38_1008 ();
 sg13g2_decap_8 FILLER_38_1015 ();
 sg13g2_decap_8 FILLER_38_1022 ();
 sg13g2_decap_8 FILLER_38_1029 ();
 sg13g2_decap_8 FILLER_38_1036 ();
 sg13g2_decap_8 FILLER_38_1043 ();
 sg13g2_decap_8 FILLER_38_1050 ();
 sg13g2_decap_8 FILLER_38_1057 ();
 sg13g2_decap_8 FILLER_38_1064 ();
 sg13g2_decap_8 FILLER_38_1071 ();
 sg13g2_decap_8 FILLER_38_1078 ();
 sg13g2_decap_8 FILLER_38_1085 ();
 sg13g2_decap_8 FILLER_38_1092 ();
 sg13g2_decap_8 FILLER_38_1099 ();
 sg13g2_decap_8 FILLER_38_1106 ();
 sg13g2_decap_8 FILLER_38_1113 ();
 sg13g2_decap_8 FILLER_38_1120 ();
 sg13g2_decap_8 FILLER_38_1127 ();
 sg13g2_decap_8 FILLER_38_1134 ();
 sg13g2_decap_8 FILLER_38_1141 ();
 sg13g2_decap_8 FILLER_38_1148 ();
 sg13g2_decap_8 FILLER_38_1155 ();
 sg13g2_decap_8 FILLER_38_1162 ();
 sg13g2_decap_8 FILLER_38_1169 ();
 sg13g2_decap_8 FILLER_38_1176 ();
 sg13g2_decap_8 FILLER_38_1183 ();
 sg13g2_decap_8 FILLER_38_1190 ();
 sg13g2_decap_8 FILLER_38_1197 ();
 sg13g2_decap_8 FILLER_38_1204 ();
 sg13g2_decap_8 FILLER_38_1211 ();
 sg13g2_decap_8 FILLER_38_1218 ();
 sg13g2_decap_8 FILLER_38_1225 ();
 sg13g2_decap_8 FILLER_38_1232 ();
 sg13g2_decap_8 FILLER_38_1239 ();
 sg13g2_decap_8 FILLER_38_1246 ();
 sg13g2_decap_8 FILLER_38_1253 ();
 sg13g2_decap_8 FILLER_38_1260 ();
 sg13g2_decap_8 FILLER_38_1267 ();
 sg13g2_decap_8 FILLER_38_1274 ();
 sg13g2_decap_8 FILLER_38_1281 ();
 sg13g2_decap_8 FILLER_38_1288 ();
 sg13g2_decap_8 FILLER_38_1295 ();
 sg13g2_decap_8 FILLER_38_1302 ();
 sg13g2_decap_8 FILLER_38_1309 ();
 sg13g2_decap_8 FILLER_38_1316 ();
 sg13g2_decap_8 FILLER_38_1323 ();
 sg13g2_decap_8 FILLER_38_1330 ();
 sg13g2_decap_8 FILLER_38_1337 ();
 sg13g2_decap_8 FILLER_38_1344 ();
 sg13g2_decap_8 FILLER_38_1351 ();
 sg13g2_decap_8 FILLER_38_1358 ();
 sg13g2_decap_8 FILLER_38_1365 ();
 sg13g2_decap_8 FILLER_38_1372 ();
 sg13g2_decap_8 FILLER_38_1379 ();
 sg13g2_decap_8 FILLER_38_1386 ();
 sg13g2_decap_8 FILLER_38_1393 ();
 sg13g2_decap_8 FILLER_38_1400 ();
 sg13g2_decap_8 FILLER_38_1407 ();
 sg13g2_decap_8 FILLER_38_1414 ();
 sg13g2_decap_8 FILLER_38_1421 ();
 sg13g2_decap_8 FILLER_38_1428 ();
 sg13g2_decap_8 FILLER_38_1435 ();
 sg13g2_decap_8 FILLER_38_1442 ();
 sg13g2_decap_8 FILLER_38_1449 ();
 sg13g2_decap_8 FILLER_38_1456 ();
 sg13g2_decap_8 FILLER_38_1463 ();
 sg13g2_decap_8 FILLER_38_1470 ();
 sg13g2_decap_8 FILLER_38_1477 ();
 sg13g2_decap_8 FILLER_38_1484 ();
 sg13g2_decap_8 FILLER_38_1491 ();
 sg13g2_decap_8 FILLER_38_1498 ();
 sg13g2_decap_8 FILLER_38_1505 ();
 sg13g2_decap_8 FILLER_38_1512 ();
 sg13g2_decap_8 FILLER_38_1519 ();
 sg13g2_decap_8 FILLER_38_1526 ();
 sg13g2_decap_8 FILLER_38_1533 ();
 sg13g2_decap_8 FILLER_38_1540 ();
 sg13g2_decap_8 FILLER_38_1547 ();
 sg13g2_decap_8 FILLER_38_1554 ();
 sg13g2_decap_8 FILLER_38_1561 ();
 sg13g2_decap_8 FILLER_38_1568 ();
 sg13g2_decap_8 FILLER_38_1575 ();
 sg13g2_decap_8 FILLER_38_1582 ();
 sg13g2_decap_8 FILLER_38_1589 ();
 sg13g2_decap_8 FILLER_38_1596 ();
 sg13g2_decap_8 FILLER_38_1603 ();
 sg13g2_decap_8 FILLER_38_1610 ();
 sg13g2_decap_8 FILLER_38_1617 ();
 sg13g2_decap_8 FILLER_38_1624 ();
 sg13g2_decap_8 FILLER_38_1631 ();
 sg13g2_decap_8 FILLER_38_1638 ();
 sg13g2_decap_8 FILLER_38_1645 ();
 sg13g2_decap_8 FILLER_38_1652 ();
 sg13g2_decap_8 FILLER_38_1659 ();
 sg13g2_decap_8 FILLER_38_1666 ();
 sg13g2_decap_8 FILLER_38_1673 ();
 sg13g2_decap_8 FILLER_38_1680 ();
 sg13g2_decap_8 FILLER_38_1687 ();
 sg13g2_decap_8 FILLER_38_1694 ();
 sg13g2_decap_8 FILLER_38_1701 ();
 sg13g2_decap_8 FILLER_38_1708 ();
 sg13g2_decap_8 FILLER_38_1715 ();
 sg13g2_decap_8 FILLER_38_1722 ();
 sg13g2_decap_8 FILLER_38_1729 ();
 sg13g2_decap_8 FILLER_38_1736 ();
 sg13g2_decap_8 FILLER_38_1743 ();
 sg13g2_decap_8 FILLER_38_1750 ();
 sg13g2_decap_8 FILLER_38_1757 ();
 sg13g2_decap_8 FILLER_38_1764 ();
 sg13g2_decap_8 FILLER_38_1771 ();
 sg13g2_decap_8 FILLER_38_1778 ();
 sg13g2_decap_8 FILLER_38_1785 ();
 sg13g2_decap_8 FILLER_38_1792 ();
 sg13g2_decap_8 FILLER_38_1799 ();
 sg13g2_decap_8 FILLER_38_1806 ();
 sg13g2_decap_8 FILLER_38_1813 ();
 sg13g2_decap_8 FILLER_38_1820 ();
 sg13g2_decap_8 FILLER_38_1827 ();
 sg13g2_decap_8 FILLER_38_1834 ();
 sg13g2_decap_8 FILLER_38_1841 ();
 sg13g2_decap_8 FILLER_38_1848 ();
 sg13g2_decap_8 FILLER_38_1855 ();
 sg13g2_decap_8 FILLER_38_1862 ();
 sg13g2_decap_8 FILLER_38_1869 ();
 sg13g2_decap_8 FILLER_38_1876 ();
 sg13g2_decap_8 FILLER_38_1883 ();
 sg13g2_decap_8 FILLER_38_1890 ();
 sg13g2_decap_8 FILLER_38_1897 ();
 sg13g2_decap_8 FILLER_38_1904 ();
 sg13g2_decap_8 FILLER_38_1911 ();
 sg13g2_decap_8 FILLER_38_1918 ();
 sg13g2_decap_8 FILLER_38_1925 ();
 sg13g2_decap_8 FILLER_38_1932 ();
 sg13g2_decap_8 FILLER_38_1939 ();
 sg13g2_decap_8 FILLER_38_1946 ();
 sg13g2_decap_8 FILLER_38_1953 ();
 sg13g2_decap_8 FILLER_38_1960 ();
 sg13g2_decap_8 FILLER_38_1967 ();
 sg13g2_decap_8 FILLER_38_1974 ();
 sg13g2_decap_8 FILLER_38_1981 ();
 sg13g2_decap_8 FILLER_38_1988 ();
 sg13g2_decap_8 FILLER_38_1995 ();
 sg13g2_decap_8 FILLER_38_2002 ();
 sg13g2_decap_8 FILLER_38_2009 ();
 sg13g2_decap_8 FILLER_38_2016 ();
 sg13g2_decap_8 FILLER_38_2023 ();
 sg13g2_decap_8 FILLER_38_2030 ();
 sg13g2_decap_8 FILLER_38_2037 ();
 sg13g2_decap_8 FILLER_38_2044 ();
 sg13g2_decap_8 FILLER_38_2051 ();
 sg13g2_decap_8 FILLER_38_2058 ();
 sg13g2_decap_8 FILLER_38_2065 ();
 sg13g2_decap_8 FILLER_38_2072 ();
 sg13g2_decap_8 FILLER_38_2079 ();
 sg13g2_decap_8 FILLER_38_2086 ();
 sg13g2_decap_8 FILLER_38_2093 ();
 sg13g2_decap_8 FILLER_38_2100 ();
 sg13g2_decap_8 FILLER_38_2107 ();
 sg13g2_decap_8 FILLER_38_2114 ();
 sg13g2_decap_8 FILLER_38_2121 ();
 sg13g2_decap_8 FILLER_38_2128 ();
 sg13g2_decap_8 FILLER_38_2135 ();
 sg13g2_decap_8 FILLER_38_2142 ();
 sg13g2_decap_8 FILLER_38_2149 ();
 sg13g2_decap_8 FILLER_38_2156 ();
 sg13g2_decap_8 FILLER_38_2163 ();
 sg13g2_decap_8 FILLER_38_2170 ();
 sg13g2_decap_8 FILLER_38_2177 ();
 sg13g2_decap_8 FILLER_38_2184 ();
 sg13g2_decap_8 FILLER_38_2191 ();
 sg13g2_decap_8 FILLER_38_2198 ();
 sg13g2_decap_8 FILLER_38_2205 ();
 sg13g2_decap_8 FILLER_38_2212 ();
 sg13g2_decap_8 FILLER_38_2219 ();
 sg13g2_decap_8 FILLER_38_2226 ();
 sg13g2_decap_8 FILLER_38_2233 ();
 sg13g2_decap_8 FILLER_38_2240 ();
 sg13g2_decap_8 FILLER_38_2247 ();
 sg13g2_decap_8 FILLER_38_2254 ();
 sg13g2_decap_8 FILLER_38_2261 ();
 sg13g2_decap_8 FILLER_38_2268 ();
 sg13g2_decap_8 FILLER_38_2275 ();
 sg13g2_decap_8 FILLER_38_2282 ();
 sg13g2_decap_8 FILLER_38_2289 ();
 sg13g2_decap_8 FILLER_38_2296 ();
 sg13g2_decap_8 FILLER_38_2303 ();
 sg13g2_decap_8 FILLER_38_2310 ();
 sg13g2_decap_8 FILLER_38_2317 ();
 sg13g2_decap_8 FILLER_38_2324 ();
 sg13g2_decap_8 FILLER_38_2331 ();
 sg13g2_decap_8 FILLER_38_2338 ();
 sg13g2_decap_8 FILLER_38_2345 ();
 sg13g2_decap_8 FILLER_38_2352 ();
 sg13g2_decap_8 FILLER_38_2359 ();
 sg13g2_decap_8 FILLER_38_2366 ();
 sg13g2_decap_8 FILLER_38_2373 ();
 sg13g2_decap_8 FILLER_38_2380 ();
 sg13g2_decap_8 FILLER_38_2387 ();
 sg13g2_decap_8 FILLER_38_2394 ();
 sg13g2_decap_8 FILLER_38_2401 ();
 sg13g2_decap_8 FILLER_38_2408 ();
 sg13g2_decap_8 FILLER_38_2415 ();
 sg13g2_decap_8 FILLER_38_2422 ();
 sg13g2_decap_8 FILLER_38_2429 ();
 sg13g2_decap_8 FILLER_38_2436 ();
 sg13g2_decap_8 FILLER_38_2443 ();
 sg13g2_decap_8 FILLER_38_2450 ();
 sg13g2_decap_8 FILLER_38_2457 ();
 sg13g2_decap_8 FILLER_38_2464 ();
 sg13g2_decap_8 FILLER_38_2471 ();
 sg13g2_decap_8 FILLER_38_2478 ();
 sg13g2_decap_8 FILLER_38_2485 ();
 sg13g2_decap_8 FILLER_38_2492 ();
 sg13g2_decap_8 FILLER_38_2499 ();
 sg13g2_decap_8 FILLER_38_2506 ();
 sg13g2_decap_8 FILLER_38_2513 ();
 sg13g2_decap_8 FILLER_38_2520 ();
 sg13g2_decap_8 FILLER_38_2527 ();
 sg13g2_decap_8 FILLER_38_2534 ();
 sg13g2_decap_8 FILLER_38_2541 ();
 sg13g2_decap_8 FILLER_38_2548 ();
 sg13g2_decap_8 FILLER_38_2555 ();
 sg13g2_decap_8 FILLER_38_2562 ();
 sg13g2_decap_8 FILLER_38_2569 ();
 sg13g2_decap_8 FILLER_38_2576 ();
 sg13g2_decap_8 FILLER_38_2583 ();
 sg13g2_decap_8 FILLER_38_2590 ();
 sg13g2_decap_8 FILLER_38_2597 ();
 sg13g2_decap_8 FILLER_38_2604 ();
 sg13g2_decap_8 FILLER_38_2611 ();
 sg13g2_decap_8 FILLER_38_2618 ();
 sg13g2_decap_8 FILLER_38_2625 ();
 sg13g2_decap_8 FILLER_38_2632 ();
 sg13g2_decap_8 FILLER_38_2639 ();
 sg13g2_decap_8 FILLER_38_2646 ();
 sg13g2_decap_8 FILLER_38_2653 ();
 sg13g2_decap_8 FILLER_38_2660 ();
 sg13g2_decap_8 FILLER_38_2667 ();
 sg13g2_decap_8 FILLER_38_2674 ();
 sg13g2_decap_8 FILLER_38_2681 ();
 sg13g2_decap_8 FILLER_38_2688 ();
 sg13g2_decap_8 FILLER_38_2695 ();
 sg13g2_decap_8 FILLER_38_2702 ();
 sg13g2_decap_8 FILLER_38_2709 ();
 sg13g2_decap_8 FILLER_38_2716 ();
 sg13g2_decap_8 FILLER_38_2723 ();
 sg13g2_decap_8 FILLER_38_2730 ();
 sg13g2_decap_8 FILLER_38_2737 ();
 sg13g2_decap_8 FILLER_38_2744 ();
 sg13g2_decap_8 FILLER_38_2751 ();
 sg13g2_decap_8 FILLER_38_2758 ();
 sg13g2_decap_8 FILLER_38_2765 ();
 sg13g2_decap_8 FILLER_38_2772 ();
 sg13g2_decap_8 FILLER_38_2779 ();
 sg13g2_decap_8 FILLER_38_2786 ();
 sg13g2_decap_8 FILLER_38_2793 ();
 sg13g2_decap_8 FILLER_38_2800 ();
 sg13g2_decap_8 FILLER_38_2807 ();
 sg13g2_decap_8 FILLER_38_2814 ();
 sg13g2_decap_8 FILLER_38_2821 ();
 sg13g2_decap_8 FILLER_38_2828 ();
 sg13g2_decap_8 FILLER_38_2835 ();
 sg13g2_decap_8 FILLER_38_2842 ();
 sg13g2_decap_8 FILLER_38_2849 ();
 sg13g2_decap_8 FILLER_38_2856 ();
 sg13g2_decap_8 FILLER_38_2863 ();
 sg13g2_decap_8 FILLER_38_2870 ();
 sg13g2_decap_8 FILLER_38_2877 ();
 sg13g2_decap_8 FILLER_38_2884 ();
 sg13g2_decap_8 FILLER_38_2891 ();
 sg13g2_decap_8 FILLER_38_2898 ();
 sg13g2_decap_8 FILLER_38_2905 ();
 sg13g2_decap_8 FILLER_38_2912 ();
 sg13g2_decap_8 FILLER_38_2919 ();
 sg13g2_decap_8 FILLER_38_2926 ();
 sg13g2_decap_8 FILLER_38_2933 ();
 sg13g2_decap_8 FILLER_38_2940 ();
 sg13g2_decap_8 FILLER_38_2947 ();
 sg13g2_decap_8 FILLER_38_2954 ();
 sg13g2_decap_8 FILLER_38_2961 ();
 sg13g2_decap_8 FILLER_38_2968 ();
 sg13g2_decap_8 FILLER_38_2975 ();
 sg13g2_decap_8 FILLER_38_2982 ();
 sg13g2_decap_8 FILLER_38_2989 ();
 sg13g2_decap_8 FILLER_38_2996 ();
 sg13g2_decap_8 FILLER_38_3003 ();
 sg13g2_decap_8 FILLER_38_3010 ();
 sg13g2_decap_8 FILLER_38_3017 ();
 sg13g2_decap_8 FILLER_38_3024 ();
 sg13g2_decap_8 FILLER_38_3031 ();
 sg13g2_decap_8 FILLER_38_3038 ();
 sg13g2_decap_8 FILLER_38_3045 ();
 sg13g2_decap_8 FILLER_38_3052 ();
 sg13g2_decap_8 FILLER_38_3059 ();
 sg13g2_decap_8 FILLER_38_3066 ();
 sg13g2_decap_8 FILLER_38_3073 ();
 sg13g2_decap_8 FILLER_38_3080 ();
 sg13g2_decap_8 FILLER_38_3087 ();
 sg13g2_decap_8 FILLER_38_3094 ();
 sg13g2_decap_8 FILLER_38_3101 ();
 sg13g2_decap_8 FILLER_38_3108 ();
 sg13g2_decap_8 FILLER_38_3115 ();
 sg13g2_decap_8 FILLER_38_3122 ();
 sg13g2_decap_8 FILLER_38_3129 ();
 sg13g2_decap_8 FILLER_38_3136 ();
 sg13g2_decap_8 FILLER_38_3143 ();
 sg13g2_decap_8 FILLER_38_3150 ();
 sg13g2_decap_8 FILLER_38_3157 ();
 sg13g2_decap_8 FILLER_38_3164 ();
 sg13g2_decap_8 FILLER_38_3171 ();
 sg13g2_decap_8 FILLER_38_3178 ();
 sg13g2_decap_8 FILLER_38_3185 ();
 sg13g2_decap_8 FILLER_38_3192 ();
 sg13g2_decap_8 FILLER_38_3199 ();
 sg13g2_decap_8 FILLER_38_3206 ();
 sg13g2_decap_8 FILLER_38_3213 ();
 sg13g2_decap_8 FILLER_38_3220 ();
 sg13g2_decap_8 FILLER_38_3227 ();
 sg13g2_decap_8 FILLER_38_3234 ();
 sg13g2_decap_8 FILLER_38_3241 ();
 sg13g2_decap_8 FILLER_38_3248 ();
 sg13g2_decap_8 FILLER_38_3255 ();
 sg13g2_decap_8 FILLER_38_3262 ();
 sg13g2_decap_8 FILLER_38_3269 ();
 sg13g2_decap_8 FILLER_38_3276 ();
 sg13g2_decap_8 FILLER_38_3283 ();
 sg13g2_decap_8 FILLER_38_3290 ();
 sg13g2_decap_8 FILLER_38_3297 ();
 sg13g2_decap_8 FILLER_38_3304 ();
 sg13g2_decap_8 FILLER_38_3311 ();
 sg13g2_decap_8 FILLER_38_3318 ();
 sg13g2_decap_8 FILLER_38_3325 ();
 sg13g2_decap_8 FILLER_38_3332 ();
 sg13g2_decap_8 FILLER_38_3339 ();
 sg13g2_decap_8 FILLER_38_3346 ();
 sg13g2_decap_8 FILLER_38_3353 ();
 sg13g2_decap_8 FILLER_38_3360 ();
 sg13g2_decap_8 FILLER_38_3367 ();
 sg13g2_decap_8 FILLER_38_3374 ();
 sg13g2_decap_8 FILLER_38_3381 ();
 sg13g2_decap_8 FILLER_38_3388 ();
 sg13g2_decap_8 FILLER_38_3395 ();
 sg13g2_decap_8 FILLER_38_3402 ();
 sg13g2_decap_8 FILLER_38_3409 ();
 sg13g2_decap_8 FILLER_38_3416 ();
 sg13g2_decap_8 FILLER_38_3423 ();
 sg13g2_decap_8 FILLER_38_3430 ();
 sg13g2_decap_8 FILLER_38_3437 ();
 sg13g2_decap_8 FILLER_38_3444 ();
 sg13g2_decap_8 FILLER_38_3451 ();
 sg13g2_decap_8 FILLER_38_3458 ();
 sg13g2_decap_8 FILLER_38_3465 ();
 sg13g2_decap_8 FILLER_38_3472 ();
 sg13g2_decap_8 FILLER_38_3479 ();
 sg13g2_decap_8 FILLER_38_3486 ();
 sg13g2_decap_8 FILLER_38_3493 ();
 sg13g2_decap_8 FILLER_38_3500 ();
 sg13g2_decap_8 FILLER_38_3507 ();
 sg13g2_decap_8 FILLER_38_3514 ();
 sg13g2_decap_8 FILLER_38_3521 ();
 sg13g2_decap_8 FILLER_38_3528 ();
 sg13g2_decap_8 FILLER_38_3535 ();
 sg13g2_decap_8 FILLER_38_3542 ();
 sg13g2_decap_8 FILLER_38_3549 ();
 sg13g2_decap_8 FILLER_38_3556 ();
 sg13g2_decap_8 FILLER_38_3563 ();
 sg13g2_decap_8 FILLER_38_3570 ();
 sg13g2_fill_2 FILLER_38_3577 ();
 sg13g2_fill_1 FILLER_38_3579 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_decap_8 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_161 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_182 ();
 sg13g2_decap_8 FILLER_39_189 ();
 sg13g2_decap_8 FILLER_39_196 ();
 sg13g2_decap_8 FILLER_39_203 ();
 sg13g2_decap_8 FILLER_39_210 ();
 sg13g2_decap_8 FILLER_39_217 ();
 sg13g2_decap_8 FILLER_39_224 ();
 sg13g2_decap_8 FILLER_39_231 ();
 sg13g2_decap_8 FILLER_39_238 ();
 sg13g2_decap_8 FILLER_39_245 ();
 sg13g2_decap_8 FILLER_39_252 ();
 sg13g2_decap_8 FILLER_39_259 ();
 sg13g2_decap_8 FILLER_39_266 ();
 sg13g2_decap_8 FILLER_39_273 ();
 sg13g2_decap_8 FILLER_39_280 ();
 sg13g2_decap_8 FILLER_39_287 ();
 sg13g2_decap_8 FILLER_39_294 ();
 sg13g2_decap_8 FILLER_39_301 ();
 sg13g2_decap_8 FILLER_39_308 ();
 sg13g2_decap_8 FILLER_39_315 ();
 sg13g2_decap_8 FILLER_39_322 ();
 sg13g2_decap_8 FILLER_39_329 ();
 sg13g2_decap_8 FILLER_39_336 ();
 sg13g2_decap_8 FILLER_39_343 ();
 sg13g2_decap_8 FILLER_39_350 ();
 sg13g2_decap_8 FILLER_39_357 ();
 sg13g2_decap_8 FILLER_39_364 ();
 sg13g2_decap_8 FILLER_39_371 ();
 sg13g2_decap_8 FILLER_39_378 ();
 sg13g2_decap_8 FILLER_39_385 ();
 sg13g2_decap_8 FILLER_39_392 ();
 sg13g2_decap_8 FILLER_39_399 ();
 sg13g2_decap_8 FILLER_39_406 ();
 sg13g2_decap_8 FILLER_39_413 ();
 sg13g2_decap_8 FILLER_39_420 ();
 sg13g2_decap_8 FILLER_39_427 ();
 sg13g2_decap_8 FILLER_39_434 ();
 sg13g2_decap_8 FILLER_39_441 ();
 sg13g2_decap_8 FILLER_39_448 ();
 sg13g2_decap_8 FILLER_39_455 ();
 sg13g2_decap_8 FILLER_39_462 ();
 sg13g2_decap_8 FILLER_39_469 ();
 sg13g2_decap_8 FILLER_39_476 ();
 sg13g2_decap_8 FILLER_39_483 ();
 sg13g2_decap_8 FILLER_39_490 ();
 sg13g2_decap_8 FILLER_39_497 ();
 sg13g2_decap_8 FILLER_39_504 ();
 sg13g2_decap_8 FILLER_39_511 ();
 sg13g2_decap_8 FILLER_39_518 ();
 sg13g2_decap_8 FILLER_39_525 ();
 sg13g2_decap_8 FILLER_39_532 ();
 sg13g2_decap_8 FILLER_39_539 ();
 sg13g2_decap_8 FILLER_39_546 ();
 sg13g2_decap_8 FILLER_39_553 ();
 sg13g2_decap_8 FILLER_39_560 ();
 sg13g2_decap_8 FILLER_39_567 ();
 sg13g2_decap_8 FILLER_39_574 ();
 sg13g2_decap_8 FILLER_39_581 ();
 sg13g2_decap_8 FILLER_39_588 ();
 sg13g2_decap_8 FILLER_39_595 ();
 sg13g2_decap_8 FILLER_39_602 ();
 sg13g2_decap_8 FILLER_39_609 ();
 sg13g2_decap_8 FILLER_39_616 ();
 sg13g2_decap_8 FILLER_39_623 ();
 sg13g2_decap_8 FILLER_39_630 ();
 sg13g2_decap_8 FILLER_39_637 ();
 sg13g2_decap_8 FILLER_39_644 ();
 sg13g2_decap_8 FILLER_39_651 ();
 sg13g2_decap_8 FILLER_39_658 ();
 sg13g2_decap_8 FILLER_39_665 ();
 sg13g2_decap_8 FILLER_39_672 ();
 sg13g2_decap_8 FILLER_39_679 ();
 sg13g2_decap_8 FILLER_39_686 ();
 sg13g2_decap_8 FILLER_39_693 ();
 sg13g2_decap_8 FILLER_39_700 ();
 sg13g2_decap_8 FILLER_39_707 ();
 sg13g2_decap_8 FILLER_39_714 ();
 sg13g2_decap_8 FILLER_39_721 ();
 sg13g2_decap_8 FILLER_39_728 ();
 sg13g2_decap_8 FILLER_39_735 ();
 sg13g2_decap_8 FILLER_39_742 ();
 sg13g2_decap_8 FILLER_39_749 ();
 sg13g2_decap_8 FILLER_39_756 ();
 sg13g2_decap_8 FILLER_39_763 ();
 sg13g2_decap_8 FILLER_39_770 ();
 sg13g2_decap_8 FILLER_39_777 ();
 sg13g2_decap_8 FILLER_39_784 ();
 sg13g2_decap_8 FILLER_39_791 ();
 sg13g2_decap_8 FILLER_39_798 ();
 sg13g2_decap_8 FILLER_39_805 ();
 sg13g2_decap_8 FILLER_39_812 ();
 sg13g2_decap_8 FILLER_39_819 ();
 sg13g2_decap_8 FILLER_39_826 ();
 sg13g2_decap_8 FILLER_39_833 ();
 sg13g2_decap_8 FILLER_39_840 ();
 sg13g2_decap_8 FILLER_39_847 ();
 sg13g2_decap_8 FILLER_39_854 ();
 sg13g2_decap_8 FILLER_39_861 ();
 sg13g2_decap_8 FILLER_39_868 ();
 sg13g2_decap_8 FILLER_39_875 ();
 sg13g2_decap_8 FILLER_39_882 ();
 sg13g2_decap_8 FILLER_39_889 ();
 sg13g2_decap_8 FILLER_39_896 ();
 sg13g2_decap_8 FILLER_39_903 ();
 sg13g2_decap_8 FILLER_39_910 ();
 sg13g2_decap_8 FILLER_39_917 ();
 sg13g2_decap_8 FILLER_39_924 ();
 sg13g2_decap_8 FILLER_39_931 ();
 sg13g2_decap_8 FILLER_39_938 ();
 sg13g2_decap_8 FILLER_39_945 ();
 sg13g2_decap_8 FILLER_39_952 ();
 sg13g2_decap_8 FILLER_39_959 ();
 sg13g2_decap_8 FILLER_39_966 ();
 sg13g2_decap_8 FILLER_39_973 ();
 sg13g2_decap_8 FILLER_39_980 ();
 sg13g2_decap_8 FILLER_39_987 ();
 sg13g2_decap_8 FILLER_39_994 ();
 sg13g2_decap_8 FILLER_39_1001 ();
 sg13g2_decap_8 FILLER_39_1008 ();
 sg13g2_decap_8 FILLER_39_1015 ();
 sg13g2_decap_8 FILLER_39_1022 ();
 sg13g2_decap_8 FILLER_39_1029 ();
 sg13g2_decap_8 FILLER_39_1036 ();
 sg13g2_decap_8 FILLER_39_1043 ();
 sg13g2_decap_8 FILLER_39_1050 ();
 sg13g2_decap_8 FILLER_39_1057 ();
 sg13g2_decap_8 FILLER_39_1064 ();
 sg13g2_decap_8 FILLER_39_1071 ();
 sg13g2_decap_8 FILLER_39_1078 ();
 sg13g2_decap_8 FILLER_39_1085 ();
 sg13g2_decap_8 FILLER_39_1092 ();
 sg13g2_decap_8 FILLER_39_1099 ();
 sg13g2_decap_8 FILLER_39_1106 ();
 sg13g2_decap_8 FILLER_39_1113 ();
 sg13g2_decap_8 FILLER_39_1120 ();
 sg13g2_decap_8 FILLER_39_1127 ();
 sg13g2_decap_8 FILLER_39_1134 ();
 sg13g2_decap_8 FILLER_39_1141 ();
 sg13g2_decap_8 FILLER_39_1148 ();
 sg13g2_decap_8 FILLER_39_1155 ();
 sg13g2_decap_8 FILLER_39_1162 ();
 sg13g2_decap_8 FILLER_39_1169 ();
 sg13g2_decap_8 FILLER_39_1176 ();
 sg13g2_decap_8 FILLER_39_1183 ();
 sg13g2_decap_8 FILLER_39_1190 ();
 sg13g2_decap_8 FILLER_39_1197 ();
 sg13g2_decap_8 FILLER_39_1204 ();
 sg13g2_decap_8 FILLER_39_1211 ();
 sg13g2_decap_8 FILLER_39_1218 ();
 sg13g2_decap_8 FILLER_39_1225 ();
 sg13g2_decap_8 FILLER_39_1232 ();
 sg13g2_decap_8 FILLER_39_1239 ();
 sg13g2_decap_8 FILLER_39_1246 ();
 sg13g2_decap_8 FILLER_39_1253 ();
 sg13g2_decap_8 FILLER_39_1260 ();
 sg13g2_decap_8 FILLER_39_1267 ();
 sg13g2_decap_8 FILLER_39_1274 ();
 sg13g2_decap_8 FILLER_39_1281 ();
 sg13g2_decap_8 FILLER_39_1288 ();
 sg13g2_decap_8 FILLER_39_1295 ();
 sg13g2_decap_8 FILLER_39_1302 ();
 sg13g2_decap_8 FILLER_39_1309 ();
 sg13g2_decap_8 FILLER_39_1316 ();
 sg13g2_decap_8 FILLER_39_1323 ();
 sg13g2_decap_8 FILLER_39_1330 ();
 sg13g2_decap_8 FILLER_39_1337 ();
 sg13g2_decap_8 FILLER_39_1344 ();
 sg13g2_decap_8 FILLER_39_1351 ();
 sg13g2_decap_8 FILLER_39_1358 ();
 sg13g2_decap_8 FILLER_39_1365 ();
 sg13g2_decap_8 FILLER_39_1372 ();
 sg13g2_decap_8 FILLER_39_1379 ();
 sg13g2_decap_8 FILLER_39_1386 ();
 sg13g2_decap_8 FILLER_39_1393 ();
 sg13g2_decap_8 FILLER_39_1400 ();
 sg13g2_decap_8 FILLER_39_1407 ();
 sg13g2_decap_8 FILLER_39_1414 ();
 sg13g2_decap_8 FILLER_39_1421 ();
 sg13g2_decap_8 FILLER_39_1428 ();
 sg13g2_decap_8 FILLER_39_1435 ();
 sg13g2_decap_8 FILLER_39_1442 ();
 sg13g2_decap_8 FILLER_39_1449 ();
 sg13g2_decap_8 FILLER_39_1456 ();
 sg13g2_decap_8 FILLER_39_1463 ();
 sg13g2_decap_8 FILLER_39_1470 ();
 sg13g2_decap_8 FILLER_39_1477 ();
 sg13g2_decap_8 FILLER_39_1484 ();
 sg13g2_decap_8 FILLER_39_1491 ();
 sg13g2_decap_8 FILLER_39_1498 ();
 sg13g2_decap_8 FILLER_39_1505 ();
 sg13g2_decap_8 FILLER_39_1512 ();
 sg13g2_decap_8 FILLER_39_1519 ();
 sg13g2_decap_8 FILLER_39_1526 ();
 sg13g2_decap_8 FILLER_39_1533 ();
 sg13g2_decap_8 FILLER_39_1540 ();
 sg13g2_decap_8 FILLER_39_1547 ();
 sg13g2_decap_8 FILLER_39_1554 ();
 sg13g2_decap_8 FILLER_39_1561 ();
 sg13g2_decap_8 FILLER_39_1568 ();
 sg13g2_decap_8 FILLER_39_1575 ();
 sg13g2_decap_8 FILLER_39_1582 ();
 sg13g2_decap_8 FILLER_39_1589 ();
 sg13g2_decap_8 FILLER_39_1596 ();
 sg13g2_decap_8 FILLER_39_1603 ();
 sg13g2_decap_8 FILLER_39_1610 ();
 sg13g2_decap_8 FILLER_39_1617 ();
 sg13g2_decap_8 FILLER_39_1624 ();
 sg13g2_decap_8 FILLER_39_1631 ();
 sg13g2_decap_8 FILLER_39_1638 ();
 sg13g2_decap_8 FILLER_39_1645 ();
 sg13g2_decap_8 FILLER_39_1652 ();
 sg13g2_decap_8 FILLER_39_1659 ();
 sg13g2_decap_8 FILLER_39_1666 ();
 sg13g2_decap_8 FILLER_39_1673 ();
 sg13g2_decap_8 FILLER_39_1680 ();
 sg13g2_decap_8 FILLER_39_1687 ();
 sg13g2_decap_8 FILLER_39_1694 ();
 sg13g2_decap_8 FILLER_39_1701 ();
 sg13g2_decap_8 FILLER_39_1708 ();
 sg13g2_decap_8 FILLER_39_1715 ();
 sg13g2_decap_8 FILLER_39_1722 ();
 sg13g2_decap_8 FILLER_39_1729 ();
 sg13g2_decap_8 FILLER_39_1736 ();
 sg13g2_decap_8 FILLER_39_1743 ();
 sg13g2_decap_8 FILLER_39_1750 ();
 sg13g2_decap_8 FILLER_39_1757 ();
 sg13g2_decap_8 FILLER_39_1764 ();
 sg13g2_decap_8 FILLER_39_1771 ();
 sg13g2_decap_8 FILLER_39_1778 ();
 sg13g2_decap_8 FILLER_39_1785 ();
 sg13g2_decap_8 FILLER_39_1792 ();
 sg13g2_decap_8 FILLER_39_1799 ();
 sg13g2_decap_8 FILLER_39_1806 ();
 sg13g2_decap_8 FILLER_39_1813 ();
 sg13g2_decap_8 FILLER_39_1820 ();
 sg13g2_decap_8 FILLER_39_1827 ();
 sg13g2_decap_8 FILLER_39_1834 ();
 sg13g2_decap_8 FILLER_39_1841 ();
 sg13g2_decap_8 FILLER_39_1848 ();
 sg13g2_decap_8 FILLER_39_1855 ();
 sg13g2_decap_8 FILLER_39_1862 ();
 sg13g2_decap_8 FILLER_39_1869 ();
 sg13g2_decap_8 FILLER_39_1876 ();
 sg13g2_decap_8 FILLER_39_1883 ();
 sg13g2_decap_8 FILLER_39_1890 ();
 sg13g2_decap_8 FILLER_39_1897 ();
 sg13g2_decap_8 FILLER_39_1904 ();
 sg13g2_decap_8 FILLER_39_1911 ();
 sg13g2_decap_8 FILLER_39_1918 ();
 sg13g2_decap_8 FILLER_39_1925 ();
 sg13g2_decap_8 FILLER_39_1932 ();
 sg13g2_decap_8 FILLER_39_1939 ();
 sg13g2_decap_8 FILLER_39_1946 ();
 sg13g2_decap_8 FILLER_39_1953 ();
 sg13g2_decap_8 FILLER_39_1960 ();
 sg13g2_decap_8 FILLER_39_1967 ();
 sg13g2_decap_8 FILLER_39_1974 ();
 sg13g2_decap_8 FILLER_39_1981 ();
 sg13g2_decap_8 FILLER_39_1988 ();
 sg13g2_decap_8 FILLER_39_1995 ();
 sg13g2_decap_8 FILLER_39_2002 ();
 sg13g2_decap_8 FILLER_39_2009 ();
 sg13g2_decap_8 FILLER_39_2016 ();
 sg13g2_decap_8 FILLER_39_2023 ();
 sg13g2_decap_8 FILLER_39_2030 ();
 sg13g2_decap_8 FILLER_39_2037 ();
 sg13g2_decap_8 FILLER_39_2044 ();
 sg13g2_decap_8 FILLER_39_2051 ();
 sg13g2_decap_8 FILLER_39_2058 ();
 sg13g2_decap_8 FILLER_39_2065 ();
 sg13g2_decap_8 FILLER_39_2072 ();
 sg13g2_decap_8 FILLER_39_2079 ();
 sg13g2_decap_8 FILLER_39_2086 ();
 sg13g2_decap_8 FILLER_39_2093 ();
 sg13g2_decap_8 FILLER_39_2100 ();
 sg13g2_decap_8 FILLER_39_2107 ();
 sg13g2_decap_8 FILLER_39_2114 ();
 sg13g2_decap_8 FILLER_39_2121 ();
 sg13g2_decap_8 FILLER_39_2128 ();
 sg13g2_decap_8 FILLER_39_2135 ();
 sg13g2_decap_8 FILLER_39_2142 ();
 sg13g2_decap_8 FILLER_39_2149 ();
 sg13g2_decap_8 FILLER_39_2156 ();
 sg13g2_decap_8 FILLER_39_2163 ();
 sg13g2_decap_8 FILLER_39_2170 ();
 sg13g2_decap_8 FILLER_39_2177 ();
 sg13g2_decap_8 FILLER_39_2184 ();
 sg13g2_decap_8 FILLER_39_2191 ();
 sg13g2_decap_8 FILLER_39_2198 ();
 sg13g2_decap_8 FILLER_39_2205 ();
 sg13g2_decap_8 FILLER_39_2212 ();
 sg13g2_decap_8 FILLER_39_2219 ();
 sg13g2_decap_8 FILLER_39_2226 ();
 sg13g2_decap_8 FILLER_39_2233 ();
 sg13g2_decap_8 FILLER_39_2240 ();
 sg13g2_decap_8 FILLER_39_2247 ();
 sg13g2_decap_8 FILLER_39_2254 ();
 sg13g2_decap_8 FILLER_39_2261 ();
 sg13g2_decap_8 FILLER_39_2268 ();
 sg13g2_decap_8 FILLER_39_2275 ();
 sg13g2_decap_8 FILLER_39_2282 ();
 sg13g2_decap_8 FILLER_39_2289 ();
 sg13g2_decap_8 FILLER_39_2296 ();
 sg13g2_decap_8 FILLER_39_2303 ();
 sg13g2_decap_8 FILLER_39_2310 ();
 sg13g2_decap_8 FILLER_39_2317 ();
 sg13g2_decap_8 FILLER_39_2324 ();
 sg13g2_decap_8 FILLER_39_2331 ();
 sg13g2_decap_8 FILLER_39_2338 ();
 sg13g2_decap_8 FILLER_39_2345 ();
 sg13g2_decap_8 FILLER_39_2352 ();
 sg13g2_decap_8 FILLER_39_2359 ();
 sg13g2_decap_8 FILLER_39_2366 ();
 sg13g2_decap_8 FILLER_39_2373 ();
 sg13g2_decap_8 FILLER_39_2380 ();
 sg13g2_decap_8 FILLER_39_2387 ();
 sg13g2_decap_8 FILLER_39_2394 ();
 sg13g2_decap_8 FILLER_39_2401 ();
 sg13g2_decap_8 FILLER_39_2408 ();
 sg13g2_decap_8 FILLER_39_2415 ();
 sg13g2_decap_8 FILLER_39_2422 ();
 sg13g2_decap_8 FILLER_39_2429 ();
 sg13g2_decap_8 FILLER_39_2436 ();
 sg13g2_decap_8 FILLER_39_2443 ();
 sg13g2_decap_8 FILLER_39_2450 ();
 sg13g2_decap_8 FILLER_39_2457 ();
 sg13g2_decap_8 FILLER_39_2464 ();
 sg13g2_decap_8 FILLER_39_2471 ();
 sg13g2_decap_8 FILLER_39_2478 ();
 sg13g2_decap_8 FILLER_39_2485 ();
 sg13g2_decap_8 FILLER_39_2492 ();
 sg13g2_decap_8 FILLER_39_2499 ();
 sg13g2_decap_8 FILLER_39_2506 ();
 sg13g2_decap_8 FILLER_39_2513 ();
 sg13g2_decap_8 FILLER_39_2520 ();
 sg13g2_decap_8 FILLER_39_2527 ();
 sg13g2_decap_8 FILLER_39_2534 ();
 sg13g2_decap_8 FILLER_39_2541 ();
 sg13g2_decap_8 FILLER_39_2548 ();
 sg13g2_decap_8 FILLER_39_2555 ();
 sg13g2_decap_8 FILLER_39_2562 ();
 sg13g2_decap_8 FILLER_39_2569 ();
 sg13g2_decap_8 FILLER_39_2576 ();
 sg13g2_decap_8 FILLER_39_2583 ();
 sg13g2_decap_8 FILLER_39_2590 ();
 sg13g2_decap_8 FILLER_39_2597 ();
 sg13g2_decap_8 FILLER_39_2604 ();
 sg13g2_decap_8 FILLER_39_2611 ();
 sg13g2_decap_8 FILLER_39_2618 ();
 sg13g2_decap_8 FILLER_39_2625 ();
 sg13g2_decap_8 FILLER_39_2632 ();
 sg13g2_decap_8 FILLER_39_2639 ();
 sg13g2_decap_8 FILLER_39_2646 ();
 sg13g2_decap_8 FILLER_39_2653 ();
 sg13g2_decap_8 FILLER_39_2660 ();
 sg13g2_decap_8 FILLER_39_2667 ();
 sg13g2_decap_8 FILLER_39_2674 ();
 sg13g2_decap_8 FILLER_39_2681 ();
 sg13g2_decap_8 FILLER_39_2688 ();
 sg13g2_decap_8 FILLER_39_2695 ();
 sg13g2_decap_8 FILLER_39_2702 ();
 sg13g2_decap_8 FILLER_39_2709 ();
 sg13g2_decap_8 FILLER_39_2716 ();
 sg13g2_decap_8 FILLER_39_2723 ();
 sg13g2_decap_8 FILLER_39_2730 ();
 sg13g2_decap_8 FILLER_39_2737 ();
 sg13g2_decap_8 FILLER_39_2744 ();
 sg13g2_decap_8 FILLER_39_2751 ();
 sg13g2_decap_8 FILLER_39_2758 ();
 sg13g2_decap_8 FILLER_39_2765 ();
 sg13g2_decap_8 FILLER_39_2772 ();
 sg13g2_decap_8 FILLER_39_2779 ();
 sg13g2_decap_8 FILLER_39_2786 ();
 sg13g2_decap_8 FILLER_39_2793 ();
 sg13g2_decap_8 FILLER_39_2800 ();
 sg13g2_decap_8 FILLER_39_2807 ();
 sg13g2_decap_8 FILLER_39_2814 ();
 sg13g2_decap_8 FILLER_39_2821 ();
 sg13g2_decap_8 FILLER_39_2828 ();
 sg13g2_decap_8 FILLER_39_2835 ();
 sg13g2_decap_8 FILLER_39_2842 ();
 sg13g2_decap_8 FILLER_39_2849 ();
 sg13g2_decap_8 FILLER_39_2856 ();
 sg13g2_decap_8 FILLER_39_2863 ();
 sg13g2_decap_8 FILLER_39_2870 ();
 sg13g2_decap_8 FILLER_39_2877 ();
 sg13g2_decap_8 FILLER_39_2884 ();
 sg13g2_decap_8 FILLER_39_2891 ();
 sg13g2_decap_8 FILLER_39_2898 ();
 sg13g2_decap_8 FILLER_39_2905 ();
 sg13g2_decap_8 FILLER_39_2912 ();
 sg13g2_decap_8 FILLER_39_2919 ();
 sg13g2_decap_8 FILLER_39_2926 ();
 sg13g2_decap_8 FILLER_39_2933 ();
 sg13g2_decap_8 FILLER_39_2940 ();
 sg13g2_decap_8 FILLER_39_2947 ();
 sg13g2_decap_8 FILLER_39_2954 ();
 sg13g2_decap_8 FILLER_39_2961 ();
 sg13g2_decap_8 FILLER_39_2968 ();
 sg13g2_decap_8 FILLER_39_2975 ();
 sg13g2_decap_8 FILLER_39_2982 ();
 sg13g2_decap_8 FILLER_39_2989 ();
 sg13g2_decap_8 FILLER_39_2996 ();
 sg13g2_decap_8 FILLER_39_3003 ();
 sg13g2_decap_8 FILLER_39_3010 ();
 sg13g2_decap_8 FILLER_39_3017 ();
 sg13g2_decap_8 FILLER_39_3024 ();
 sg13g2_decap_8 FILLER_39_3031 ();
 sg13g2_decap_8 FILLER_39_3038 ();
 sg13g2_decap_8 FILLER_39_3045 ();
 sg13g2_decap_8 FILLER_39_3052 ();
 sg13g2_decap_8 FILLER_39_3059 ();
 sg13g2_decap_8 FILLER_39_3066 ();
 sg13g2_decap_8 FILLER_39_3073 ();
 sg13g2_decap_8 FILLER_39_3080 ();
 sg13g2_decap_8 FILLER_39_3087 ();
 sg13g2_decap_8 FILLER_39_3094 ();
 sg13g2_decap_8 FILLER_39_3101 ();
 sg13g2_decap_8 FILLER_39_3108 ();
 sg13g2_decap_8 FILLER_39_3115 ();
 sg13g2_decap_8 FILLER_39_3122 ();
 sg13g2_decap_8 FILLER_39_3129 ();
 sg13g2_decap_8 FILLER_39_3136 ();
 sg13g2_decap_8 FILLER_39_3143 ();
 sg13g2_decap_8 FILLER_39_3150 ();
 sg13g2_decap_8 FILLER_39_3157 ();
 sg13g2_decap_8 FILLER_39_3164 ();
 sg13g2_decap_8 FILLER_39_3171 ();
 sg13g2_decap_8 FILLER_39_3178 ();
 sg13g2_decap_8 FILLER_39_3185 ();
 sg13g2_decap_8 FILLER_39_3192 ();
 sg13g2_decap_8 FILLER_39_3199 ();
 sg13g2_decap_8 FILLER_39_3206 ();
 sg13g2_decap_8 FILLER_39_3213 ();
 sg13g2_decap_8 FILLER_39_3220 ();
 sg13g2_decap_8 FILLER_39_3227 ();
 sg13g2_decap_8 FILLER_39_3234 ();
 sg13g2_decap_8 FILLER_39_3241 ();
 sg13g2_decap_8 FILLER_39_3248 ();
 sg13g2_decap_8 FILLER_39_3255 ();
 sg13g2_decap_8 FILLER_39_3262 ();
 sg13g2_decap_8 FILLER_39_3269 ();
 sg13g2_decap_8 FILLER_39_3276 ();
 sg13g2_decap_8 FILLER_39_3283 ();
 sg13g2_decap_8 FILLER_39_3290 ();
 sg13g2_decap_8 FILLER_39_3297 ();
 sg13g2_decap_8 FILLER_39_3304 ();
 sg13g2_decap_8 FILLER_39_3311 ();
 sg13g2_decap_8 FILLER_39_3318 ();
 sg13g2_decap_8 FILLER_39_3325 ();
 sg13g2_decap_8 FILLER_39_3332 ();
 sg13g2_decap_8 FILLER_39_3339 ();
 sg13g2_decap_8 FILLER_39_3346 ();
 sg13g2_decap_8 FILLER_39_3353 ();
 sg13g2_decap_8 FILLER_39_3360 ();
 sg13g2_decap_8 FILLER_39_3367 ();
 sg13g2_decap_8 FILLER_39_3374 ();
 sg13g2_decap_8 FILLER_39_3381 ();
 sg13g2_decap_8 FILLER_39_3388 ();
 sg13g2_decap_8 FILLER_39_3395 ();
 sg13g2_decap_8 FILLER_39_3402 ();
 sg13g2_decap_8 FILLER_39_3409 ();
 sg13g2_decap_8 FILLER_39_3416 ();
 sg13g2_decap_8 FILLER_39_3423 ();
 sg13g2_decap_8 FILLER_39_3430 ();
 sg13g2_decap_8 FILLER_39_3437 ();
 sg13g2_decap_8 FILLER_39_3444 ();
 sg13g2_decap_8 FILLER_39_3451 ();
 sg13g2_decap_8 FILLER_39_3458 ();
 sg13g2_decap_8 FILLER_39_3465 ();
 sg13g2_decap_8 FILLER_39_3472 ();
 sg13g2_decap_8 FILLER_39_3479 ();
 sg13g2_decap_8 FILLER_39_3486 ();
 sg13g2_decap_8 FILLER_39_3493 ();
 sg13g2_decap_8 FILLER_39_3500 ();
 sg13g2_decap_8 FILLER_39_3507 ();
 sg13g2_decap_8 FILLER_39_3514 ();
 sg13g2_decap_8 FILLER_39_3521 ();
 sg13g2_decap_8 FILLER_39_3528 ();
 sg13g2_decap_8 FILLER_39_3535 ();
 sg13g2_decap_8 FILLER_39_3542 ();
 sg13g2_decap_8 FILLER_39_3549 ();
 sg13g2_decap_8 FILLER_39_3556 ();
 sg13g2_decap_8 FILLER_39_3563 ();
 sg13g2_decap_8 FILLER_39_3570 ();
 sg13g2_fill_2 FILLER_39_3577 ();
 sg13g2_fill_1 FILLER_39_3579 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_decap_8 FILLER_40_147 ();
 sg13g2_decap_8 FILLER_40_154 ();
 sg13g2_decap_8 FILLER_40_161 ();
 sg13g2_decap_8 FILLER_40_168 ();
 sg13g2_decap_8 FILLER_40_175 ();
 sg13g2_decap_8 FILLER_40_182 ();
 sg13g2_decap_8 FILLER_40_189 ();
 sg13g2_decap_8 FILLER_40_196 ();
 sg13g2_decap_8 FILLER_40_203 ();
 sg13g2_decap_8 FILLER_40_210 ();
 sg13g2_decap_8 FILLER_40_217 ();
 sg13g2_decap_8 FILLER_40_224 ();
 sg13g2_decap_8 FILLER_40_231 ();
 sg13g2_decap_8 FILLER_40_238 ();
 sg13g2_decap_8 FILLER_40_245 ();
 sg13g2_decap_8 FILLER_40_252 ();
 sg13g2_decap_8 FILLER_40_259 ();
 sg13g2_decap_8 FILLER_40_266 ();
 sg13g2_decap_8 FILLER_40_273 ();
 sg13g2_decap_8 FILLER_40_280 ();
 sg13g2_decap_8 FILLER_40_287 ();
 sg13g2_decap_8 FILLER_40_294 ();
 sg13g2_decap_8 FILLER_40_301 ();
 sg13g2_decap_8 FILLER_40_308 ();
 sg13g2_decap_8 FILLER_40_315 ();
 sg13g2_decap_8 FILLER_40_322 ();
 sg13g2_decap_8 FILLER_40_329 ();
 sg13g2_decap_8 FILLER_40_336 ();
 sg13g2_decap_8 FILLER_40_343 ();
 sg13g2_decap_8 FILLER_40_350 ();
 sg13g2_decap_8 FILLER_40_357 ();
 sg13g2_decap_8 FILLER_40_364 ();
 sg13g2_decap_8 FILLER_40_371 ();
 sg13g2_decap_8 FILLER_40_378 ();
 sg13g2_decap_8 FILLER_40_385 ();
 sg13g2_decap_8 FILLER_40_392 ();
 sg13g2_decap_8 FILLER_40_399 ();
 sg13g2_decap_8 FILLER_40_406 ();
 sg13g2_decap_8 FILLER_40_413 ();
 sg13g2_decap_8 FILLER_40_420 ();
 sg13g2_decap_8 FILLER_40_427 ();
 sg13g2_decap_8 FILLER_40_434 ();
 sg13g2_decap_8 FILLER_40_441 ();
 sg13g2_decap_8 FILLER_40_448 ();
 sg13g2_decap_8 FILLER_40_455 ();
 sg13g2_decap_8 FILLER_40_462 ();
 sg13g2_decap_8 FILLER_40_469 ();
 sg13g2_decap_8 FILLER_40_476 ();
 sg13g2_decap_8 FILLER_40_483 ();
 sg13g2_decap_8 FILLER_40_490 ();
 sg13g2_decap_8 FILLER_40_497 ();
 sg13g2_decap_8 FILLER_40_504 ();
 sg13g2_decap_8 FILLER_40_511 ();
 sg13g2_decap_8 FILLER_40_518 ();
 sg13g2_decap_8 FILLER_40_525 ();
 sg13g2_decap_8 FILLER_40_532 ();
 sg13g2_decap_8 FILLER_40_539 ();
 sg13g2_decap_8 FILLER_40_546 ();
 sg13g2_decap_8 FILLER_40_553 ();
 sg13g2_decap_8 FILLER_40_560 ();
 sg13g2_decap_8 FILLER_40_567 ();
 sg13g2_decap_8 FILLER_40_574 ();
 sg13g2_decap_8 FILLER_40_581 ();
 sg13g2_decap_8 FILLER_40_588 ();
 sg13g2_decap_8 FILLER_40_595 ();
 sg13g2_decap_8 FILLER_40_602 ();
 sg13g2_decap_8 FILLER_40_609 ();
 sg13g2_decap_8 FILLER_40_616 ();
 sg13g2_decap_8 FILLER_40_623 ();
 sg13g2_decap_8 FILLER_40_630 ();
 sg13g2_decap_8 FILLER_40_637 ();
 sg13g2_decap_8 FILLER_40_644 ();
 sg13g2_decap_8 FILLER_40_651 ();
 sg13g2_decap_8 FILLER_40_658 ();
 sg13g2_decap_8 FILLER_40_665 ();
 sg13g2_decap_8 FILLER_40_672 ();
 sg13g2_decap_8 FILLER_40_679 ();
 sg13g2_decap_8 FILLER_40_686 ();
 sg13g2_decap_8 FILLER_40_693 ();
 sg13g2_decap_8 FILLER_40_700 ();
 sg13g2_decap_8 FILLER_40_707 ();
 sg13g2_decap_8 FILLER_40_714 ();
 sg13g2_decap_8 FILLER_40_721 ();
 sg13g2_decap_8 FILLER_40_728 ();
 sg13g2_decap_8 FILLER_40_735 ();
 sg13g2_decap_8 FILLER_40_742 ();
 sg13g2_decap_8 FILLER_40_749 ();
 sg13g2_decap_8 FILLER_40_756 ();
 sg13g2_decap_8 FILLER_40_763 ();
 sg13g2_decap_8 FILLER_40_770 ();
 sg13g2_decap_8 FILLER_40_777 ();
 sg13g2_decap_8 FILLER_40_784 ();
 sg13g2_decap_8 FILLER_40_791 ();
 sg13g2_decap_8 FILLER_40_798 ();
 sg13g2_decap_8 FILLER_40_805 ();
 sg13g2_decap_8 FILLER_40_812 ();
 sg13g2_decap_8 FILLER_40_819 ();
 sg13g2_decap_8 FILLER_40_826 ();
 sg13g2_decap_8 FILLER_40_833 ();
 sg13g2_decap_8 FILLER_40_840 ();
 sg13g2_decap_8 FILLER_40_847 ();
 sg13g2_decap_8 FILLER_40_854 ();
 sg13g2_decap_8 FILLER_40_861 ();
 sg13g2_decap_8 FILLER_40_868 ();
 sg13g2_decap_8 FILLER_40_875 ();
 sg13g2_decap_8 FILLER_40_882 ();
 sg13g2_decap_8 FILLER_40_889 ();
 sg13g2_decap_8 FILLER_40_896 ();
 sg13g2_decap_8 FILLER_40_903 ();
 sg13g2_decap_8 FILLER_40_910 ();
 sg13g2_decap_8 FILLER_40_917 ();
 sg13g2_decap_8 FILLER_40_924 ();
 sg13g2_decap_8 FILLER_40_931 ();
 sg13g2_decap_8 FILLER_40_938 ();
 sg13g2_decap_8 FILLER_40_945 ();
 sg13g2_decap_8 FILLER_40_952 ();
 sg13g2_decap_8 FILLER_40_959 ();
 sg13g2_decap_8 FILLER_40_966 ();
 sg13g2_decap_8 FILLER_40_973 ();
 sg13g2_decap_8 FILLER_40_980 ();
 sg13g2_decap_8 FILLER_40_987 ();
 sg13g2_decap_8 FILLER_40_994 ();
 sg13g2_decap_8 FILLER_40_1001 ();
 sg13g2_decap_8 FILLER_40_1008 ();
 sg13g2_decap_8 FILLER_40_1015 ();
 sg13g2_decap_8 FILLER_40_1022 ();
 sg13g2_decap_8 FILLER_40_1029 ();
 sg13g2_decap_8 FILLER_40_1036 ();
 sg13g2_decap_8 FILLER_40_1043 ();
 sg13g2_decap_8 FILLER_40_1050 ();
 sg13g2_decap_8 FILLER_40_1057 ();
 sg13g2_decap_8 FILLER_40_1064 ();
 sg13g2_decap_8 FILLER_40_1071 ();
 sg13g2_decap_8 FILLER_40_1078 ();
 sg13g2_decap_8 FILLER_40_1085 ();
 sg13g2_decap_8 FILLER_40_1092 ();
 sg13g2_decap_8 FILLER_40_1099 ();
 sg13g2_decap_8 FILLER_40_1106 ();
 sg13g2_decap_8 FILLER_40_1113 ();
 sg13g2_decap_8 FILLER_40_1120 ();
 sg13g2_decap_8 FILLER_40_1127 ();
 sg13g2_decap_8 FILLER_40_1134 ();
 sg13g2_decap_8 FILLER_40_1141 ();
 sg13g2_decap_8 FILLER_40_1148 ();
 sg13g2_decap_8 FILLER_40_1155 ();
 sg13g2_decap_8 FILLER_40_1162 ();
 sg13g2_decap_8 FILLER_40_1169 ();
 sg13g2_decap_8 FILLER_40_1176 ();
 sg13g2_decap_8 FILLER_40_1183 ();
 sg13g2_decap_8 FILLER_40_1190 ();
 sg13g2_decap_8 FILLER_40_1197 ();
 sg13g2_decap_8 FILLER_40_1204 ();
 sg13g2_decap_8 FILLER_40_1211 ();
 sg13g2_decap_8 FILLER_40_1218 ();
 sg13g2_decap_8 FILLER_40_1225 ();
 sg13g2_decap_8 FILLER_40_1232 ();
 sg13g2_decap_8 FILLER_40_1239 ();
 sg13g2_decap_8 FILLER_40_1246 ();
 sg13g2_decap_8 FILLER_40_1253 ();
 sg13g2_decap_8 FILLER_40_1260 ();
 sg13g2_decap_8 FILLER_40_1267 ();
 sg13g2_decap_8 FILLER_40_1274 ();
 sg13g2_decap_8 FILLER_40_1281 ();
 sg13g2_decap_8 FILLER_40_1288 ();
 sg13g2_decap_8 FILLER_40_1295 ();
 sg13g2_decap_8 FILLER_40_1302 ();
 sg13g2_decap_8 FILLER_40_1309 ();
 sg13g2_decap_8 FILLER_40_1316 ();
 sg13g2_decap_8 FILLER_40_1323 ();
 sg13g2_decap_8 FILLER_40_1330 ();
 sg13g2_decap_8 FILLER_40_1337 ();
 sg13g2_decap_8 FILLER_40_1344 ();
 sg13g2_decap_8 FILLER_40_1351 ();
 sg13g2_decap_8 FILLER_40_1358 ();
 sg13g2_decap_8 FILLER_40_1365 ();
 sg13g2_decap_8 FILLER_40_1372 ();
 sg13g2_decap_8 FILLER_40_1379 ();
 sg13g2_decap_8 FILLER_40_1386 ();
 sg13g2_decap_8 FILLER_40_1393 ();
 sg13g2_decap_8 FILLER_40_1400 ();
 sg13g2_decap_8 FILLER_40_1407 ();
 sg13g2_decap_8 FILLER_40_1414 ();
 sg13g2_decap_8 FILLER_40_1421 ();
 sg13g2_decap_8 FILLER_40_1428 ();
 sg13g2_decap_8 FILLER_40_1435 ();
 sg13g2_decap_8 FILLER_40_1442 ();
 sg13g2_decap_8 FILLER_40_1449 ();
 sg13g2_decap_8 FILLER_40_1456 ();
 sg13g2_decap_8 FILLER_40_1463 ();
 sg13g2_decap_8 FILLER_40_1470 ();
 sg13g2_decap_8 FILLER_40_1477 ();
 sg13g2_decap_8 FILLER_40_1484 ();
 sg13g2_decap_8 FILLER_40_1491 ();
 sg13g2_decap_8 FILLER_40_1498 ();
 sg13g2_decap_8 FILLER_40_1505 ();
 sg13g2_decap_8 FILLER_40_1512 ();
 sg13g2_decap_8 FILLER_40_1519 ();
 sg13g2_decap_8 FILLER_40_1526 ();
 sg13g2_decap_8 FILLER_40_1533 ();
 sg13g2_decap_8 FILLER_40_1540 ();
 sg13g2_decap_8 FILLER_40_1547 ();
 sg13g2_decap_8 FILLER_40_1554 ();
 sg13g2_decap_8 FILLER_40_1561 ();
 sg13g2_decap_8 FILLER_40_1568 ();
 sg13g2_decap_8 FILLER_40_1575 ();
 sg13g2_decap_8 FILLER_40_1582 ();
 sg13g2_decap_8 FILLER_40_1589 ();
 sg13g2_decap_8 FILLER_40_1596 ();
 sg13g2_decap_8 FILLER_40_1603 ();
 sg13g2_decap_8 FILLER_40_1610 ();
 sg13g2_decap_8 FILLER_40_1617 ();
 sg13g2_decap_8 FILLER_40_1624 ();
 sg13g2_decap_8 FILLER_40_1631 ();
 sg13g2_decap_8 FILLER_40_1638 ();
 sg13g2_decap_8 FILLER_40_1645 ();
 sg13g2_decap_8 FILLER_40_1652 ();
 sg13g2_decap_8 FILLER_40_1659 ();
 sg13g2_decap_8 FILLER_40_1666 ();
 sg13g2_decap_8 FILLER_40_1673 ();
 sg13g2_decap_8 FILLER_40_1680 ();
 sg13g2_decap_8 FILLER_40_1687 ();
 sg13g2_decap_8 FILLER_40_1694 ();
 sg13g2_decap_8 FILLER_40_1701 ();
 sg13g2_decap_8 FILLER_40_1708 ();
 sg13g2_decap_8 FILLER_40_1715 ();
 sg13g2_decap_8 FILLER_40_1722 ();
 sg13g2_decap_8 FILLER_40_1729 ();
 sg13g2_decap_8 FILLER_40_1736 ();
 sg13g2_decap_8 FILLER_40_1743 ();
 sg13g2_decap_8 FILLER_40_1750 ();
 sg13g2_decap_8 FILLER_40_1757 ();
 sg13g2_decap_8 FILLER_40_1764 ();
 sg13g2_decap_8 FILLER_40_1771 ();
 sg13g2_decap_8 FILLER_40_1778 ();
 sg13g2_decap_8 FILLER_40_1785 ();
 sg13g2_decap_8 FILLER_40_1792 ();
 sg13g2_decap_8 FILLER_40_1799 ();
 sg13g2_decap_8 FILLER_40_1806 ();
 sg13g2_decap_8 FILLER_40_1813 ();
 sg13g2_decap_8 FILLER_40_1820 ();
 sg13g2_decap_8 FILLER_40_1827 ();
 sg13g2_decap_8 FILLER_40_1834 ();
 sg13g2_decap_8 FILLER_40_1841 ();
 sg13g2_decap_8 FILLER_40_1848 ();
 sg13g2_decap_8 FILLER_40_1855 ();
 sg13g2_decap_8 FILLER_40_1862 ();
 sg13g2_decap_8 FILLER_40_1869 ();
 sg13g2_decap_8 FILLER_40_1876 ();
 sg13g2_decap_8 FILLER_40_1883 ();
 sg13g2_decap_8 FILLER_40_1890 ();
 sg13g2_decap_8 FILLER_40_1897 ();
 sg13g2_decap_8 FILLER_40_1904 ();
 sg13g2_decap_8 FILLER_40_1911 ();
 sg13g2_decap_8 FILLER_40_1918 ();
 sg13g2_decap_8 FILLER_40_1925 ();
 sg13g2_decap_8 FILLER_40_1932 ();
 sg13g2_decap_8 FILLER_40_1939 ();
 sg13g2_decap_8 FILLER_40_1946 ();
 sg13g2_decap_8 FILLER_40_1953 ();
 sg13g2_decap_8 FILLER_40_1960 ();
 sg13g2_decap_8 FILLER_40_1967 ();
 sg13g2_decap_8 FILLER_40_1974 ();
 sg13g2_decap_8 FILLER_40_1981 ();
 sg13g2_decap_8 FILLER_40_1988 ();
 sg13g2_decap_8 FILLER_40_1995 ();
 sg13g2_decap_8 FILLER_40_2002 ();
 sg13g2_decap_8 FILLER_40_2009 ();
 sg13g2_decap_8 FILLER_40_2016 ();
 sg13g2_decap_8 FILLER_40_2023 ();
 sg13g2_decap_8 FILLER_40_2030 ();
 sg13g2_decap_8 FILLER_40_2037 ();
 sg13g2_decap_8 FILLER_40_2044 ();
 sg13g2_decap_8 FILLER_40_2051 ();
 sg13g2_decap_8 FILLER_40_2058 ();
 sg13g2_decap_8 FILLER_40_2065 ();
 sg13g2_decap_8 FILLER_40_2072 ();
 sg13g2_decap_8 FILLER_40_2079 ();
 sg13g2_decap_8 FILLER_40_2086 ();
 sg13g2_decap_8 FILLER_40_2093 ();
 sg13g2_decap_8 FILLER_40_2100 ();
 sg13g2_decap_8 FILLER_40_2107 ();
 sg13g2_decap_8 FILLER_40_2114 ();
 sg13g2_decap_8 FILLER_40_2121 ();
 sg13g2_decap_8 FILLER_40_2128 ();
 sg13g2_decap_8 FILLER_40_2135 ();
 sg13g2_decap_8 FILLER_40_2142 ();
 sg13g2_decap_8 FILLER_40_2149 ();
 sg13g2_decap_8 FILLER_40_2156 ();
 sg13g2_decap_8 FILLER_40_2163 ();
 sg13g2_decap_8 FILLER_40_2170 ();
 sg13g2_decap_8 FILLER_40_2177 ();
 sg13g2_decap_8 FILLER_40_2184 ();
 sg13g2_decap_8 FILLER_40_2191 ();
 sg13g2_decap_8 FILLER_40_2198 ();
 sg13g2_decap_8 FILLER_40_2205 ();
 sg13g2_decap_8 FILLER_40_2212 ();
 sg13g2_decap_8 FILLER_40_2219 ();
 sg13g2_decap_8 FILLER_40_2226 ();
 sg13g2_decap_8 FILLER_40_2233 ();
 sg13g2_decap_8 FILLER_40_2240 ();
 sg13g2_decap_8 FILLER_40_2247 ();
 sg13g2_decap_8 FILLER_40_2254 ();
 sg13g2_decap_8 FILLER_40_2261 ();
 sg13g2_decap_8 FILLER_40_2268 ();
 sg13g2_decap_8 FILLER_40_2275 ();
 sg13g2_decap_8 FILLER_40_2282 ();
 sg13g2_decap_8 FILLER_40_2289 ();
 sg13g2_decap_8 FILLER_40_2296 ();
 sg13g2_decap_8 FILLER_40_2303 ();
 sg13g2_decap_8 FILLER_40_2310 ();
 sg13g2_decap_8 FILLER_40_2317 ();
 sg13g2_decap_8 FILLER_40_2324 ();
 sg13g2_decap_8 FILLER_40_2331 ();
 sg13g2_decap_8 FILLER_40_2338 ();
 sg13g2_decap_8 FILLER_40_2345 ();
 sg13g2_decap_8 FILLER_40_2352 ();
 sg13g2_decap_8 FILLER_40_2359 ();
 sg13g2_decap_8 FILLER_40_2366 ();
 sg13g2_decap_8 FILLER_40_2373 ();
 sg13g2_decap_8 FILLER_40_2380 ();
 sg13g2_decap_8 FILLER_40_2387 ();
 sg13g2_decap_8 FILLER_40_2394 ();
 sg13g2_decap_8 FILLER_40_2401 ();
 sg13g2_decap_8 FILLER_40_2408 ();
 sg13g2_decap_8 FILLER_40_2415 ();
 sg13g2_decap_8 FILLER_40_2422 ();
 sg13g2_decap_8 FILLER_40_2429 ();
 sg13g2_decap_8 FILLER_40_2436 ();
 sg13g2_decap_8 FILLER_40_2443 ();
 sg13g2_decap_8 FILLER_40_2450 ();
 sg13g2_decap_8 FILLER_40_2457 ();
 sg13g2_decap_8 FILLER_40_2464 ();
 sg13g2_decap_8 FILLER_40_2471 ();
 sg13g2_decap_8 FILLER_40_2478 ();
 sg13g2_decap_8 FILLER_40_2485 ();
 sg13g2_decap_8 FILLER_40_2492 ();
 sg13g2_decap_8 FILLER_40_2499 ();
 sg13g2_decap_8 FILLER_40_2506 ();
 sg13g2_decap_8 FILLER_40_2513 ();
 sg13g2_decap_8 FILLER_40_2520 ();
 sg13g2_decap_8 FILLER_40_2527 ();
 sg13g2_decap_8 FILLER_40_2534 ();
 sg13g2_decap_8 FILLER_40_2541 ();
 sg13g2_decap_8 FILLER_40_2548 ();
 sg13g2_decap_8 FILLER_40_2555 ();
 sg13g2_decap_8 FILLER_40_2562 ();
 sg13g2_decap_8 FILLER_40_2569 ();
 sg13g2_decap_8 FILLER_40_2576 ();
 sg13g2_decap_8 FILLER_40_2583 ();
 sg13g2_decap_8 FILLER_40_2590 ();
 sg13g2_decap_8 FILLER_40_2597 ();
 sg13g2_decap_8 FILLER_40_2604 ();
 sg13g2_decap_8 FILLER_40_2611 ();
 sg13g2_decap_8 FILLER_40_2618 ();
 sg13g2_decap_8 FILLER_40_2625 ();
 sg13g2_decap_8 FILLER_40_2632 ();
 sg13g2_decap_8 FILLER_40_2639 ();
 sg13g2_decap_8 FILLER_40_2646 ();
 sg13g2_decap_8 FILLER_40_2653 ();
 sg13g2_decap_8 FILLER_40_2660 ();
 sg13g2_decap_8 FILLER_40_2667 ();
 sg13g2_decap_8 FILLER_40_2674 ();
 sg13g2_decap_8 FILLER_40_2681 ();
 sg13g2_decap_8 FILLER_40_2688 ();
 sg13g2_decap_8 FILLER_40_2695 ();
 sg13g2_decap_8 FILLER_40_2702 ();
 sg13g2_decap_8 FILLER_40_2709 ();
 sg13g2_decap_8 FILLER_40_2716 ();
 sg13g2_decap_8 FILLER_40_2723 ();
 sg13g2_decap_8 FILLER_40_2730 ();
 sg13g2_decap_8 FILLER_40_2737 ();
 sg13g2_decap_8 FILLER_40_2744 ();
 sg13g2_decap_8 FILLER_40_2751 ();
 sg13g2_decap_8 FILLER_40_2758 ();
 sg13g2_decap_8 FILLER_40_2765 ();
 sg13g2_decap_8 FILLER_40_2772 ();
 sg13g2_decap_8 FILLER_40_2779 ();
 sg13g2_decap_8 FILLER_40_2786 ();
 sg13g2_decap_8 FILLER_40_2793 ();
 sg13g2_decap_8 FILLER_40_2800 ();
 sg13g2_decap_8 FILLER_40_2807 ();
 sg13g2_decap_8 FILLER_40_2814 ();
 sg13g2_decap_8 FILLER_40_2821 ();
 sg13g2_decap_8 FILLER_40_2828 ();
 sg13g2_decap_8 FILLER_40_2835 ();
 sg13g2_decap_8 FILLER_40_2842 ();
 sg13g2_decap_8 FILLER_40_2849 ();
 sg13g2_decap_8 FILLER_40_2856 ();
 sg13g2_decap_8 FILLER_40_2863 ();
 sg13g2_decap_8 FILLER_40_2870 ();
 sg13g2_decap_8 FILLER_40_2877 ();
 sg13g2_decap_8 FILLER_40_2884 ();
 sg13g2_decap_8 FILLER_40_2891 ();
 sg13g2_decap_8 FILLER_40_2898 ();
 sg13g2_decap_8 FILLER_40_2905 ();
 sg13g2_decap_8 FILLER_40_2912 ();
 sg13g2_decap_8 FILLER_40_2919 ();
 sg13g2_decap_8 FILLER_40_2926 ();
 sg13g2_decap_8 FILLER_40_2933 ();
 sg13g2_decap_8 FILLER_40_2940 ();
 sg13g2_decap_8 FILLER_40_2947 ();
 sg13g2_decap_8 FILLER_40_2954 ();
 sg13g2_decap_8 FILLER_40_2961 ();
 sg13g2_decap_8 FILLER_40_2968 ();
 sg13g2_decap_8 FILLER_40_2975 ();
 sg13g2_decap_8 FILLER_40_2982 ();
 sg13g2_decap_8 FILLER_40_2989 ();
 sg13g2_decap_8 FILLER_40_2996 ();
 sg13g2_decap_8 FILLER_40_3003 ();
 sg13g2_decap_8 FILLER_40_3010 ();
 sg13g2_decap_8 FILLER_40_3017 ();
 sg13g2_decap_8 FILLER_40_3024 ();
 sg13g2_decap_8 FILLER_40_3031 ();
 sg13g2_decap_8 FILLER_40_3038 ();
 sg13g2_decap_8 FILLER_40_3045 ();
 sg13g2_decap_8 FILLER_40_3052 ();
 sg13g2_decap_8 FILLER_40_3059 ();
 sg13g2_decap_8 FILLER_40_3066 ();
 sg13g2_decap_8 FILLER_40_3073 ();
 sg13g2_decap_8 FILLER_40_3080 ();
 sg13g2_decap_8 FILLER_40_3087 ();
 sg13g2_decap_8 FILLER_40_3094 ();
 sg13g2_decap_8 FILLER_40_3101 ();
 sg13g2_decap_8 FILLER_40_3108 ();
 sg13g2_decap_8 FILLER_40_3115 ();
 sg13g2_decap_8 FILLER_40_3122 ();
 sg13g2_decap_8 FILLER_40_3129 ();
 sg13g2_decap_8 FILLER_40_3136 ();
 sg13g2_decap_8 FILLER_40_3143 ();
 sg13g2_decap_8 FILLER_40_3150 ();
 sg13g2_decap_8 FILLER_40_3157 ();
 sg13g2_decap_8 FILLER_40_3164 ();
 sg13g2_decap_8 FILLER_40_3171 ();
 sg13g2_decap_8 FILLER_40_3178 ();
 sg13g2_decap_8 FILLER_40_3185 ();
 sg13g2_decap_8 FILLER_40_3192 ();
 sg13g2_decap_8 FILLER_40_3199 ();
 sg13g2_decap_8 FILLER_40_3206 ();
 sg13g2_decap_8 FILLER_40_3213 ();
 sg13g2_decap_8 FILLER_40_3220 ();
 sg13g2_decap_8 FILLER_40_3227 ();
 sg13g2_decap_8 FILLER_40_3234 ();
 sg13g2_decap_8 FILLER_40_3241 ();
 sg13g2_decap_8 FILLER_40_3248 ();
 sg13g2_decap_8 FILLER_40_3255 ();
 sg13g2_decap_8 FILLER_40_3262 ();
 sg13g2_decap_8 FILLER_40_3269 ();
 sg13g2_decap_8 FILLER_40_3276 ();
 sg13g2_decap_8 FILLER_40_3283 ();
 sg13g2_decap_8 FILLER_40_3290 ();
 sg13g2_decap_8 FILLER_40_3297 ();
 sg13g2_decap_8 FILLER_40_3304 ();
 sg13g2_decap_8 FILLER_40_3311 ();
 sg13g2_decap_8 FILLER_40_3318 ();
 sg13g2_decap_8 FILLER_40_3325 ();
 sg13g2_decap_8 FILLER_40_3332 ();
 sg13g2_decap_8 FILLER_40_3339 ();
 sg13g2_decap_8 FILLER_40_3346 ();
 sg13g2_decap_8 FILLER_40_3353 ();
 sg13g2_decap_8 FILLER_40_3360 ();
 sg13g2_decap_8 FILLER_40_3367 ();
 sg13g2_decap_8 FILLER_40_3374 ();
 sg13g2_decap_8 FILLER_40_3381 ();
 sg13g2_decap_8 FILLER_40_3388 ();
 sg13g2_decap_8 FILLER_40_3395 ();
 sg13g2_decap_8 FILLER_40_3402 ();
 sg13g2_decap_8 FILLER_40_3409 ();
 sg13g2_decap_8 FILLER_40_3416 ();
 sg13g2_decap_8 FILLER_40_3423 ();
 sg13g2_decap_8 FILLER_40_3430 ();
 sg13g2_decap_8 FILLER_40_3437 ();
 sg13g2_decap_8 FILLER_40_3444 ();
 sg13g2_decap_8 FILLER_40_3451 ();
 sg13g2_decap_8 FILLER_40_3458 ();
 sg13g2_decap_8 FILLER_40_3465 ();
 sg13g2_decap_8 FILLER_40_3472 ();
 sg13g2_decap_8 FILLER_40_3479 ();
 sg13g2_decap_8 FILLER_40_3486 ();
 sg13g2_decap_8 FILLER_40_3493 ();
 sg13g2_decap_8 FILLER_40_3500 ();
 sg13g2_decap_8 FILLER_40_3507 ();
 sg13g2_decap_8 FILLER_40_3514 ();
 sg13g2_decap_8 FILLER_40_3521 ();
 sg13g2_decap_8 FILLER_40_3528 ();
 sg13g2_decap_8 FILLER_40_3535 ();
 sg13g2_decap_8 FILLER_40_3542 ();
 sg13g2_decap_8 FILLER_40_3549 ();
 sg13g2_decap_8 FILLER_40_3556 ();
 sg13g2_decap_8 FILLER_40_3563 ();
 sg13g2_decap_8 FILLER_40_3570 ();
 sg13g2_fill_2 FILLER_40_3577 ();
 sg13g2_fill_1 FILLER_40_3579 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_8 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_154 ();
 sg13g2_decap_8 FILLER_41_161 ();
 sg13g2_decap_8 FILLER_41_168 ();
 sg13g2_decap_8 FILLER_41_175 ();
 sg13g2_decap_8 FILLER_41_182 ();
 sg13g2_decap_8 FILLER_41_189 ();
 sg13g2_decap_8 FILLER_41_196 ();
 sg13g2_decap_8 FILLER_41_203 ();
 sg13g2_decap_8 FILLER_41_210 ();
 sg13g2_decap_8 FILLER_41_217 ();
 sg13g2_decap_8 FILLER_41_224 ();
 sg13g2_decap_8 FILLER_41_231 ();
 sg13g2_decap_8 FILLER_41_238 ();
 sg13g2_decap_8 FILLER_41_245 ();
 sg13g2_decap_8 FILLER_41_252 ();
 sg13g2_decap_8 FILLER_41_259 ();
 sg13g2_decap_8 FILLER_41_266 ();
 sg13g2_decap_8 FILLER_41_273 ();
 sg13g2_decap_8 FILLER_41_280 ();
 sg13g2_decap_8 FILLER_41_287 ();
 sg13g2_decap_8 FILLER_41_294 ();
 sg13g2_decap_8 FILLER_41_301 ();
 sg13g2_decap_8 FILLER_41_308 ();
 sg13g2_decap_8 FILLER_41_315 ();
 sg13g2_decap_8 FILLER_41_322 ();
 sg13g2_decap_8 FILLER_41_329 ();
 sg13g2_decap_8 FILLER_41_336 ();
 sg13g2_decap_8 FILLER_41_343 ();
 sg13g2_decap_8 FILLER_41_350 ();
 sg13g2_decap_8 FILLER_41_357 ();
 sg13g2_decap_8 FILLER_41_364 ();
 sg13g2_decap_8 FILLER_41_371 ();
 sg13g2_decap_8 FILLER_41_378 ();
 sg13g2_decap_8 FILLER_41_385 ();
 sg13g2_decap_8 FILLER_41_392 ();
 sg13g2_decap_8 FILLER_41_399 ();
 sg13g2_decap_8 FILLER_41_406 ();
 sg13g2_decap_8 FILLER_41_413 ();
 sg13g2_decap_8 FILLER_41_420 ();
 sg13g2_decap_8 FILLER_41_427 ();
 sg13g2_decap_8 FILLER_41_434 ();
 sg13g2_decap_8 FILLER_41_441 ();
 sg13g2_decap_8 FILLER_41_448 ();
 sg13g2_decap_8 FILLER_41_455 ();
 sg13g2_decap_8 FILLER_41_462 ();
 sg13g2_decap_8 FILLER_41_469 ();
 sg13g2_decap_8 FILLER_41_476 ();
 sg13g2_decap_8 FILLER_41_483 ();
 sg13g2_decap_8 FILLER_41_490 ();
 sg13g2_decap_8 FILLER_41_497 ();
 sg13g2_decap_8 FILLER_41_504 ();
 sg13g2_decap_8 FILLER_41_511 ();
 sg13g2_decap_8 FILLER_41_518 ();
 sg13g2_decap_8 FILLER_41_525 ();
 sg13g2_decap_8 FILLER_41_532 ();
 sg13g2_decap_8 FILLER_41_539 ();
 sg13g2_decap_8 FILLER_41_546 ();
 sg13g2_decap_8 FILLER_41_553 ();
 sg13g2_decap_8 FILLER_41_560 ();
 sg13g2_decap_8 FILLER_41_567 ();
 sg13g2_decap_8 FILLER_41_574 ();
 sg13g2_decap_8 FILLER_41_581 ();
 sg13g2_decap_8 FILLER_41_588 ();
 sg13g2_decap_8 FILLER_41_595 ();
 sg13g2_decap_8 FILLER_41_602 ();
 sg13g2_decap_8 FILLER_41_609 ();
 sg13g2_decap_8 FILLER_41_616 ();
 sg13g2_decap_8 FILLER_41_623 ();
 sg13g2_decap_8 FILLER_41_630 ();
 sg13g2_decap_8 FILLER_41_637 ();
 sg13g2_decap_8 FILLER_41_644 ();
 sg13g2_decap_8 FILLER_41_651 ();
 sg13g2_decap_8 FILLER_41_658 ();
 sg13g2_decap_8 FILLER_41_665 ();
 sg13g2_decap_8 FILLER_41_672 ();
 sg13g2_decap_8 FILLER_41_679 ();
 sg13g2_decap_8 FILLER_41_686 ();
 sg13g2_decap_8 FILLER_41_693 ();
 sg13g2_decap_8 FILLER_41_700 ();
 sg13g2_decap_8 FILLER_41_707 ();
 sg13g2_decap_8 FILLER_41_714 ();
 sg13g2_decap_8 FILLER_41_721 ();
 sg13g2_decap_8 FILLER_41_728 ();
 sg13g2_decap_8 FILLER_41_735 ();
 sg13g2_decap_8 FILLER_41_742 ();
 sg13g2_decap_8 FILLER_41_749 ();
 sg13g2_decap_8 FILLER_41_756 ();
 sg13g2_decap_8 FILLER_41_763 ();
 sg13g2_decap_8 FILLER_41_770 ();
 sg13g2_decap_8 FILLER_41_777 ();
 sg13g2_decap_8 FILLER_41_784 ();
 sg13g2_decap_8 FILLER_41_791 ();
 sg13g2_decap_8 FILLER_41_798 ();
 sg13g2_decap_8 FILLER_41_805 ();
 sg13g2_decap_8 FILLER_41_812 ();
 sg13g2_decap_8 FILLER_41_819 ();
 sg13g2_decap_8 FILLER_41_826 ();
 sg13g2_decap_8 FILLER_41_833 ();
 sg13g2_decap_8 FILLER_41_840 ();
 sg13g2_decap_8 FILLER_41_847 ();
 sg13g2_decap_8 FILLER_41_854 ();
 sg13g2_decap_8 FILLER_41_861 ();
 sg13g2_decap_8 FILLER_41_868 ();
 sg13g2_decap_8 FILLER_41_875 ();
 sg13g2_decap_8 FILLER_41_882 ();
 sg13g2_decap_8 FILLER_41_889 ();
 sg13g2_decap_8 FILLER_41_896 ();
 sg13g2_decap_8 FILLER_41_903 ();
 sg13g2_decap_8 FILLER_41_910 ();
 sg13g2_decap_8 FILLER_41_917 ();
 sg13g2_decap_8 FILLER_41_924 ();
 sg13g2_decap_8 FILLER_41_931 ();
 sg13g2_decap_8 FILLER_41_938 ();
 sg13g2_decap_8 FILLER_41_945 ();
 sg13g2_decap_8 FILLER_41_952 ();
 sg13g2_decap_8 FILLER_41_959 ();
 sg13g2_decap_8 FILLER_41_966 ();
 sg13g2_decap_8 FILLER_41_973 ();
 sg13g2_decap_8 FILLER_41_980 ();
 sg13g2_decap_8 FILLER_41_987 ();
 sg13g2_decap_8 FILLER_41_994 ();
 sg13g2_decap_8 FILLER_41_1001 ();
 sg13g2_decap_8 FILLER_41_1008 ();
 sg13g2_decap_8 FILLER_41_1015 ();
 sg13g2_decap_8 FILLER_41_1022 ();
 sg13g2_decap_8 FILLER_41_1029 ();
 sg13g2_decap_8 FILLER_41_1036 ();
 sg13g2_decap_8 FILLER_41_1043 ();
 sg13g2_decap_8 FILLER_41_1050 ();
 sg13g2_decap_8 FILLER_41_1057 ();
 sg13g2_decap_8 FILLER_41_1064 ();
 sg13g2_decap_8 FILLER_41_1071 ();
 sg13g2_decap_8 FILLER_41_1078 ();
 sg13g2_decap_8 FILLER_41_1085 ();
 sg13g2_decap_8 FILLER_41_1092 ();
 sg13g2_decap_8 FILLER_41_1099 ();
 sg13g2_decap_8 FILLER_41_1106 ();
 sg13g2_decap_8 FILLER_41_1113 ();
 sg13g2_decap_8 FILLER_41_1120 ();
 sg13g2_decap_8 FILLER_41_1127 ();
 sg13g2_decap_8 FILLER_41_1134 ();
 sg13g2_decap_8 FILLER_41_1141 ();
 sg13g2_decap_8 FILLER_41_1148 ();
 sg13g2_decap_8 FILLER_41_1155 ();
 sg13g2_decap_8 FILLER_41_1162 ();
 sg13g2_decap_8 FILLER_41_1169 ();
 sg13g2_decap_8 FILLER_41_1176 ();
 sg13g2_decap_8 FILLER_41_1183 ();
 sg13g2_decap_8 FILLER_41_1190 ();
 sg13g2_decap_8 FILLER_41_1197 ();
 sg13g2_decap_8 FILLER_41_1204 ();
 sg13g2_decap_8 FILLER_41_1211 ();
 sg13g2_decap_8 FILLER_41_1218 ();
 sg13g2_decap_8 FILLER_41_1225 ();
 sg13g2_decap_8 FILLER_41_1232 ();
 sg13g2_decap_8 FILLER_41_1239 ();
 sg13g2_decap_8 FILLER_41_1246 ();
 sg13g2_decap_8 FILLER_41_1253 ();
 sg13g2_decap_8 FILLER_41_1260 ();
 sg13g2_decap_8 FILLER_41_1267 ();
 sg13g2_decap_8 FILLER_41_1274 ();
 sg13g2_decap_8 FILLER_41_1281 ();
 sg13g2_decap_8 FILLER_41_1288 ();
 sg13g2_decap_8 FILLER_41_1295 ();
 sg13g2_decap_8 FILLER_41_1302 ();
 sg13g2_decap_8 FILLER_41_1309 ();
 sg13g2_decap_8 FILLER_41_1316 ();
 sg13g2_decap_8 FILLER_41_1323 ();
 sg13g2_decap_8 FILLER_41_1330 ();
 sg13g2_decap_8 FILLER_41_1337 ();
 sg13g2_decap_8 FILLER_41_1344 ();
 sg13g2_decap_8 FILLER_41_1351 ();
 sg13g2_decap_8 FILLER_41_1358 ();
 sg13g2_decap_8 FILLER_41_1365 ();
 sg13g2_decap_8 FILLER_41_1372 ();
 sg13g2_decap_8 FILLER_41_1379 ();
 sg13g2_decap_8 FILLER_41_1386 ();
 sg13g2_decap_8 FILLER_41_1393 ();
 sg13g2_decap_8 FILLER_41_1400 ();
 sg13g2_decap_8 FILLER_41_1407 ();
 sg13g2_decap_8 FILLER_41_1414 ();
 sg13g2_decap_8 FILLER_41_1421 ();
 sg13g2_decap_8 FILLER_41_1428 ();
 sg13g2_decap_8 FILLER_41_1435 ();
 sg13g2_decap_8 FILLER_41_1442 ();
 sg13g2_decap_8 FILLER_41_1449 ();
 sg13g2_decap_8 FILLER_41_1456 ();
 sg13g2_decap_8 FILLER_41_1463 ();
 sg13g2_decap_8 FILLER_41_1470 ();
 sg13g2_decap_8 FILLER_41_1477 ();
 sg13g2_decap_8 FILLER_41_1484 ();
 sg13g2_decap_8 FILLER_41_1491 ();
 sg13g2_decap_8 FILLER_41_1498 ();
 sg13g2_decap_8 FILLER_41_1505 ();
 sg13g2_decap_8 FILLER_41_1512 ();
 sg13g2_decap_8 FILLER_41_1519 ();
 sg13g2_decap_8 FILLER_41_1526 ();
 sg13g2_decap_8 FILLER_41_1533 ();
 sg13g2_decap_8 FILLER_41_1540 ();
 sg13g2_decap_8 FILLER_41_1547 ();
 sg13g2_decap_8 FILLER_41_1554 ();
 sg13g2_decap_8 FILLER_41_1561 ();
 sg13g2_decap_8 FILLER_41_1568 ();
 sg13g2_decap_8 FILLER_41_1575 ();
 sg13g2_decap_8 FILLER_41_1582 ();
 sg13g2_decap_8 FILLER_41_1589 ();
 sg13g2_decap_8 FILLER_41_1596 ();
 sg13g2_decap_8 FILLER_41_1603 ();
 sg13g2_decap_8 FILLER_41_1610 ();
 sg13g2_decap_8 FILLER_41_1617 ();
 sg13g2_decap_8 FILLER_41_1624 ();
 sg13g2_decap_8 FILLER_41_1631 ();
 sg13g2_decap_8 FILLER_41_1638 ();
 sg13g2_decap_8 FILLER_41_1645 ();
 sg13g2_decap_8 FILLER_41_1652 ();
 sg13g2_decap_8 FILLER_41_1659 ();
 sg13g2_decap_8 FILLER_41_1666 ();
 sg13g2_decap_8 FILLER_41_1673 ();
 sg13g2_decap_8 FILLER_41_1680 ();
 sg13g2_decap_8 FILLER_41_1687 ();
 sg13g2_decap_8 FILLER_41_1694 ();
 sg13g2_decap_8 FILLER_41_1701 ();
 sg13g2_decap_8 FILLER_41_1708 ();
 sg13g2_decap_8 FILLER_41_1715 ();
 sg13g2_decap_8 FILLER_41_1722 ();
 sg13g2_decap_8 FILLER_41_1729 ();
 sg13g2_decap_8 FILLER_41_1736 ();
 sg13g2_decap_8 FILLER_41_1743 ();
 sg13g2_decap_8 FILLER_41_1750 ();
 sg13g2_decap_8 FILLER_41_1757 ();
 sg13g2_decap_8 FILLER_41_1764 ();
 sg13g2_decap_8 FILLER_41_1771 ();
 sg13g2_decap_8 FILLER_41_1778 ();
 sg13g2_decap_8 FILLER_41_1785 ();
 sg13g2_decap_8 FILLER_41_1792 ();
 sg13g2_decap_8 FILLER_41_1799 ();
 sg13g2_decap_8 FILLER_41_1806 ();
 sg13g2_decap_8 FILLER_41_1813 ();
 sg13g2_decap_8 FILLER_41_1820 ();
 sg13g2_decap_8 FILLER_41_1827 ();
 sg13g2_decap_8 FILLER_41_1834 ();
 sg13g2_decap_8 FILLER_41_1841 ();
 sg13g2_decap_8 FILLER_41_1848 ();
 sg13g2_decap_8 FILLER_41_1855 ();
 sg13g2_decap_8 FILLER_41_1862 ();
 sg13g2_decap_8 FILLER_41_1869 ();
 sg13g2_decap_8 FILLER_41_1876 ();
 sg13g2_decap_8 FILLER_41_1883 ();
 sg13g2_decap_8 FILLER_41_1890 ();
 sg13g2_decap_8 FILLER_41_1897 ();
 sg13g2_decap_8 FILLER_41_1904 ();
 sg13g2_decap_8 FILLER_41_1911 ();
 sg13g2_decap_8 FILLER_41_1918 ();
 sg13g2_decap_8 FILLER_41_1925 ();
 sg13g2_decap_8 FILLER_41_1932 ();
 sg13g2_decap_8 FILLER_41_1939 ();
 sg13g2_decap_8 FILLER_41_1946 ();
 sg13g2_decap_8 FILLER_41_1953 ();
 sg13g2_decap_8 FILLER_41_1960 ();
 sg13g2_decap_8 FILLER_41_1967 ();
 sg13g2_decap_8 FILLER_41_1974 ();
 sg13g2_decap_8 FILLER_41_1981 ();
 sg13g2_decap_8 FILLER_41_1988 ();
 sg13g2_decap_8 FILLER_41_1995 ();
 sg13g2_decap_8 FILLER_41_2002 ();
 sg13g2_decap_8 FILLER_41_2009 ();
 sg13g2_decap_8 FILLER_41_2016 ();
 sg13g2_decap_8 FILLER_41_2023 ();
 sg13g2_decap_8 FILLER_41_2030 ();
 sg13g2_decap_8 FILLER_41_2037 ();
 sg13g2_decap_8 FILLER_41_2044 ();
 sg13g2_decap_8 FILLER_41_2051 ();
 sg13g2_decap_8 FILLER_41_2058 ();
 sg13g2_decap_8 FILLER_41_2065 ();
 sg13g2_decap_8 FILLER_41_2072 ();
 sg13g2_decap_8 FILLER_41_2079 ();
 sg13g2_decap_8 FILLER_41_2086 ();
 sg13g2_decap_8 FILLER_41_2093 ();
 sg13g2_decap_8 FILLER_41_2100 ();
 sg13g2_decap_8 FILLER_41_2107 ();
 sg13g2_decap_8 FILLER_41_2114 ();
 sg13g2_decap_8 FILLER_41_2121 ();
 sg13g2_decap_8 FILLER_41_2128 ();
 sg13g2_decap_8 FILLER_41_2135 ();
 sg13g2_decap_8 FILLER_41_2142 ();
 sg13g2_decap_8 FILLER_41_2149 ();
 sg13g2_decap_8 FILLER_41_2156 ();
 sg13g2_decap_8 FILLER_41_2163 ();
 sg13g2_decap_8 FILLER_41_2170 ();
 sg13g2_decap_8 FILLER_41_2177 ();
 sg13g2_decap_8 FILLER_41_2184 ();
 sg13g2_decap_8 FILLER_41_2191 ();
 sg13g2_decap_8 FILLER_41_2198 ();
 sg13g2_decap_8 FILLER_41_2205 ();
 sg13g2_decap_8 FILLER_41_2212 ();
 sg13g2_decap_8 FILLER_41_2219 ();
 sg13g2_decap_8 FILLER_41_2226 ();
 sg13g2_decap_8 FILLER_41_2233 ();
 sg13g2_decap_8 FILLER_41_2240 ();
 sg13g2_decap_8 FILLER_41_2247 ();
 sg13g2_decap_8 FILLER_41_2254 ();
 sg13g2_decap_8 FILLER_41_2261 ();
 sg13g2_decap_8 FILLER_41_2268 ();
 sg13g2_decap_8 FILLER_41_2275 ();
 sg13g2_decap_8 FILLER_41_2282 ();
 sg13g2_decap_8 FILLER_41_2289 ();
 sg13g2_decap_8 FILLER_41_2296 ();
 sg13g2_decap_8 FILLER_41_2303 ();
 sg13g2_decap_8 FILLER_41_2310 ();
 sg13g2_decap_8 FILLER_41_2317 ();
 sg13g2_decap_8 FILLER_41_2324 ();
 sg13g2_decap_8 FILLER_41_2331 ();
 sg13g2_decap_8 FILLER_41_2338 ();
 sg13g2_decap_8 FILLER_41_2345 ();
 sg13g2_decap_8 FILLER_41_2352 ();
 sg13g2_decap_8 FILLER_41_2359 ();
 sg13g2_decap_8 FILLER_41_2366 ();
 sg13g2_decap_8 FILLER_41_2373 ();
 sg13g2_decap_8 FILLER_41_2380 ();
 sg13g2_decap_8 FILLER_41_2387 ();
 sg13g2_decap_8 FILLER_41_2394 ();
 sg13g2_decap_8 FILLER_41_2401 ();
 sg13g2_decap_8 FILLER_41_2408 ();
 sg13g2_decap_8 FILLER_41_2415 ();
 sg13g2_decap_8 FILLER_41_2422 ();
 sg13g2_decap_8 FILLER_41_2429 ();
 sg13g2_decap_8 FILLER_41_2436 ();
 sg13g2_decap_8 FILLER_41_2443 ();
 sg13g2_decap_8 FILLER_41_2450 ();
 sg13g2_decap_8 FILLER_41_2457 ();
 sg13g2_decap_8 FILLER_41_2464 ();
 sg13g2_decap_8 FILLER_41_2471 ();
 sg13g2_decap_8 FILLER_41_2478 ();
 sg13g2_decap_8 FILLER_41_2485 ();
 sg13g2_decap_8 FILLER_41_2492 ();
 sg13g2_decap_8 FILLER_41_2499 ();
 sg13g2_decap_8 FILLER_41_2506 ();
 sg13g2_decap_8 FILLER_41_2513 ();
 sg13g2_decap_8 FILLER_41_2520 ();
 sg13g2_decap_8 FILLER_41_2527 ();
 sg13g2_decap_8 FILLER_41_2534 ();
 sg13g2_decap_8 FILLER_41_2541 ();
 sg13g2_decap_8 FILLER_41_2548 ();
 sg13g2_decap_8 FILLER_41_2555 ();
 sg13g2_decap_8 FILLER_41_2562 ();
 sg13g2_decap_8 FILLER_41_2569 ();
 sg13g2_decap_8 FILLER_41_2576 ();
 sg13g2_decap_8 FILLER_41_2583 ();
 sg13g2_decap_8 FILLER_41_2590 ();
 sg13g2_decap_8 FILLER_41_2597 ();
 sg13g2_decap_8 FILLER_41_2604 ();
 sg13g2_decap_8 FILLER_41_2611 ();
 sg13g2_decap_8 FILLER_41_2618 ();
 sg13g2_decap_8 FILLER_41_2625 ();
 sg13g2_decap_8 FILLER_41_2632 ();
 sg13g2_decap_8 FILLER_41_2639 ();
 sg13g2_decap_8 FILLER_41_2646 ();
 sg13g2_decap_8 FILLER_41_2653 ();
 sg13g2_decap_8 FILLER_41_2660 ();
 sg13g2_decap_8 FILLER_41_2667 ();
 sg13g2_decap_8 FILLER_41_2674 ();
 sg13g2_decap_8 FILLER_41_2681 ();
 sg13g2_decap_8 FILLER_41_2688 ();
 sg13g2_decap_8 FILLER_41_2695 ();
 sg13g2_decap_8 FILLER_41_2702 ();
 sg13g2_decap_8 FILLER_41_2709 ();
 sg13g2_decap_8 FILLER_41_2716 ();
 sg13g2_decap_8 FILLER_41_2723 ();
 sg13g2_decap_8 FILLER_41_2730 ();
 sg13g2_decap_8 FILLER_41_2737 ();
 sg13g2_decap_8 FILLER_41_2744 ();
 sg13g2_decap_8 FILLER_41_2751 ();
 sg13g2_decap_8 FILLER_41_2758 ();
 sg13g2_decap_8 FILLER_41_2765 ();
 sg13g2_decap_8 FILLER_41_2772 ();
 sg13g2_decap_8 FILLER_41_2779 ();
 sg13g2_decap_8 FILLER_41_2786 ();
 sg13g2_decap_8 FILLER_41_2793 ();
 sg13g2_decap_8 FILLER_41_2800 ();
 sg13g2_decap_8 FILLER_41_2807 ();
 sg13g2_decap_8 FILLER_41_2814 ();
 sg13g2_decap_8 FILLER_41_2821 ();
 sg13g2_decap_8 FILLER_41_2828 ();
 sg13g2_decap_8 FILLER_41_2835 ();
 sg13g2_decap_8 FILLER_41_2842 ();
 sg13g2_decap_8 FILLER_41_2849 ();
 sg13g2_decap_8 FILLER_41_2856 ();
 sg13g2_decap_8 FILLER_41_2863 ();
 sg13g2_decap_8 FILLER_41_2870 ();
 sg13g2_decap_8 FILLER_41_2877 ();
 sg13g2_decap_8 FILLER_41_2884 ();
 sg13g2_decap_8 FILLER_41_2891 ();
 sg13g2_decap_8 FILLER_41_2898 ();
 sg13g2_decap_8 FILLER_41_2905 ();
 sg13g2_decap_8 FILLER_41_2912 ();
 sg13g2_decap_8 FILLER_41_2919 ();
 sg13g2_decap_8 FILLER_41_2926 ();
 sg13g2_decap_8 FILLER_41_2933 ();
 sg13g2_decap_8 FILLER_41_2940 ();
 sg13g2_decap_8 FILLER_41_2947 ();
 sg13g2_decap_8 FILLER_41_2954 ();
 sg13g2_decap_8 FILLER_41_2961 ();
 sg13g2_decap_8 FILLER_41_2968 ();
 sg13g2_decap_8 FILLER_41_2975 ();
 sg13g2_decap_8 FILLER_41_2982 ();
 sg13g2_decap_8 FILLER_41_2989 ();
 sg13g2_decap_8 FILLER_41_2996 ();
 sg13g2_decap_8 FILLER_41_3003 ();
 sg13g2_decap_8 FILLER_41_3010 ();
 sg13g2_decap_8 FILLER_41_3017 ();
 sg13g2_decap_8 FILLER_41_3024 ();
 sg13g2_decap_8 FILLER_41_3031 ();
 sg13g2_decap_8 FILLER_41_3038 ();
 sg13g2_decap_8 FILLER_41_3045 ();
 sg13g2_decap_8 FILLER_41_3052 ();
 sg13g2_decap_8 FILLER_41_3059 ();
 sg13g2_decap_8 FILLER_41_3066 ();
 sg13g2_decap_8 FILLER_41_3073 ();
 sg13g2_decap_8 FILLER_41_3080 ();
 sg13g2_decap_8 FILLER_41_3087 ();
 sg13g2_decap_8 FILLER_41_3094 ();
 sg13g2_decap_8 FILLER_41_3101 ();
 sg13g2_decap_8 FILLER_41_3108 ();
 sg13g2_decap_8 FILLER_41_3115 ();
 sg13g2_decap_8 FILLER_41_3122 ();
 sg13g2_decap_8 FILLER_41_3129 ();
 sg13g2_decap_8 FILLER_41_3136 ();
 sg13g2_decap_8 FILLER_41_3143 ();
 sg13g2_decap_8 FILLER_41_3150 ();
 sg13g2_decap_8 FILLER_41_3157 ();
 sg13g2_decap_8 FILLER_41_3164 ();
 sg13g2_decap_8 FILLER_41_3171 ();
 sg13g2_decap_8 FILLER_41_3178 ();
 sg13g2_decap_8 FILLER_41_3185 ();
 sg13g2_decap_8 FILLER_41_3192 ();
 sg13g2_decap_8 FILLER_41_3199 ();
 sg13g2_decap_8 FILLER_41_3206 ();
 sg13g2_decap_8 FILLER_41_3213 ();
 sg13g2_decap_8 FILLER_41_3220 ();
 sg13g2_decap_8 FILLER_41_3227 ();
 sg13g2_decap_8 FILLER_41_3234 ();
 sg13g2_decap_8 FILLER_41_3241 ();
 sg13g2_decap_8 FILLER_41_3248 ();
 sg13g2_decap_8 FILLER_41_3255 ();
 sg13g2_decap_8 FILLER_41_3262 ();
 sg13g2_decap_8 FILLER_41_3269 ();
 sg13g2_decap_8 FILLER_41_3276 ();
 sg13g2_decap_8 FILLER_41_3283 ();
 sg13g2_decap_8 FILLER_41_3290 ();
 sg13g2_decap_8 FILLER_41_3297 ();
 sg13g2_decap_8 FILLER_41_3304 ();
 sg13g2_decap_8 FILLER_41_3311 ();
 sg13g2_decap_8 FILLER_41_3318 ();
 sg13g2_decap_8 FILLER_41_3325 ();
 sg13g2_decap_8 FILLER_41_3332 ();
 sg13g2_decap_8 FILLER_41_3339 ();
 sg13g2_decap_8 FILLER_41_3346 ();
 sg13g2_decap_8 FILLER_41_3353 ();
 sg13g2_decap_8 FILLER_41_3360 ();
 sg13g2_decap_8 FILLER_41_3367 ();
 sg13g2_decap_8 FILLER_41_3374 ();
 sg13g2_decap_8 FILLER_41_3381 ();
 sg13g2_decap_8 FILLER_41_3388 ();
 sg13g2_decap_8 FILLER_41_3395 ();
 sg13g2_decap_8 FILLER_41_3402 ();
 sg13g2_decap_8 FILLER_41_3409 ();
 sg13g2_decap_8 FILLER_41_3416 ();
 sg13g2_decap_8 FILLER_41_3423 ();
 sg13g2_decap_8 FILLER_41_3430 ();
 sg13g2_decap_8 FILLER_41_3437 ();
 sg13g2_decap_8 FILLER_41_3444 ();
 sg13g2_decap_8 FILLER_41_3451 ();
 sg13g2_decap_8 FILLER_41_3458 ();
 sg13g2_decap_8 FILLER_41_3465 ();
 sg13g2_decap_8 FILLER_41_3472 ();
 sg13g2_decap_8 FILLER_41_3479 ();
 sg13g2_decap_8 FILLER_41_3486 ();
 sg13g2_decap_8 FILLER_41_3493 ();
 sg13g2_decap_8 FILLER_41_3500 ();
 sg13g2_decap_8 FILLER_41_3507 ();
 sg13g2_decap_8 FILLER_41_3514 ();
 sg13g2_decap_8 FILLER_41_3521 ();
 sg13g2_decap_8 FILLER_41_3528 ();
 sg13g2_decap_8 FILLER_41_3535 ();
 sg13g2_decap_8 FILLER_41_3542 ();
 sg13g2_decap_8 FILLER_41_3549 ();
 sg13g2_decap_8 FILLER_41_3556 ();
 sg13g2_decap_8 FILLER_41_3563 ();
 sg13g2_decap_8 FILLER_41_3570 ();
 sg13g2_fill_2 FILLER_41_3577 ();
 sg13g2_fill_1 FILLER_41_3579 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_decap_8 FILLER_42_154 ();
 sg13g2_decap_8 FILLER_42_161 ();
 sg13g2_decap_8 FILLER_42_168 ();
 sg13g2_decap_8 FILLER_42_175 ();
 sg13g2_decap_8 FILLER_42_182 ();
 sg13g2_decap_8 FILLER_42_189 ();
 sg13g2_decap_8 FILLER_42_196 ();
 sg13g2_decap_8 FILLER_42_203 ();
 sg13g2_decap_8 FILLER_42_210 ();
 sg13g2_decap_8 FILLER_42_217 ();
 sg13g2_decap_8 FILLER_42_224 ();
 sg13g2_decap_8 FILLER_42_231 ();
 sg13g2_decap_8 FILLER_42_238 ();
 sg13g2_decap_8 FILLER_42_245 ();
 sg13g2_decap_8 FILLER_42_252 ();
 sg13g2_decap_8 FILLER_42_259 ();
 sg13g2_decap_8 FILLER_42_266 ();
 sg13g2_decap_8 FILLER_42_273 ();
 sg13g2_decap_8 FILLER_42_280 ();
 sg13g2_decap_8 FILLER_42_287 ();
 sg13g2_decap_8 FILLER_42_294 ();
 sg13g2_decap_8 FILLER_42_301 ();
 sg13g2_decap_8 FILLER_42_308 ();
 sg13g2_decap_8 FILLER_42_315 ();
 sg13g2_decap_8 FILLER_42_322 ();
 sg13g2_decap_8 FILLER_42_329 ();
 sg13g2_decap_8 FILLER_42_336 ();
 sg13g2_decap_8 FILLER_42_343 ();
 sg13g2_decap_8 FILLER_42_350 ();
 sg13g2_decap_8 FILLER_42_357 ();
 sg13g2_decap_8 FILLER_42_364 ();
 sg13g2_decap_8 FILLER_42_371 ();
 sg13g2_decap_8 FILLER_42_378 ();
 sg13g2_decap_8 FILLER_42_385 ();
 sg13g2_decap_8 FILLER_42_392 ();
 sg13g2_decap_8 FILLER_42_399 ();
 sg13g2_decap_8 FILLER_42_406 ();
 sg13g2_decap_8 FILLER_42_413 ();
 sg13g2_decap_8 FILLER_42_420 ();
 sg13g2_decap_8 FILLER_42_427 ();
 sg13g2_decap_8 FILLER_42_434 ();
 sg13g2_decap_8 FILLER_42_441 ();
 sg13g2_decap_8 FILLER_42_448 ();
 sg13g2_decap_8 FILLER_42_455 ();
 sg13g2_decap_8 FILLER_42_462 ();
 sg13g2_decap_8 FILLER_42_469 ();
 sg13g2_decap_8 FILLER_42_476 ();
 sg13g2_decap_8 FILLER_42_483 ();
 sg13g2_decap_8 FILLER_42_490 ();
 sg13g2_decap_8 FILLER_42_497 ();
 sg13g2_decap_8 FILLER_42_504 ();
 sg13g2_decap_8 FILLER_42_511 ();
 sg13g2_decap_8 FILLER_42_518 ();
 sg13g2_decap_8 FILLER_42_525 ();
 sg13g2_decap_8 FILLER_42_532 ();
 sg13g2_decap_8 FILLER_42_539 ();
 sg13g2_decap_8 FILLER_42_546 ();
 sg13g2_decap_8 FILLER_42_553 ();
 sg13g2_decap_8 FILLER_42_560 ();
 sg13g2_decap_8 FILLER_42_567 ();
 sg13g2_decap_8 FILLER_42_574 ();
 sg13g2_decap_8 FILLER_42_581 ();
 sg13g2_decap_8 FILLER_42_588 ();
 sg13g2_decap_8 FILLER_42_595 ();
 sg13g2_decap_8 FILLER_42_602 ();
 sg13g2_decap_8 FILLER_42_609 ();
 sg13g2_decap_8 FILLER_42_616 ();
 sg13g2_decap_8 FILLER_42_623 ();
 sg13g2_decap_8 FILLER_42_630 ();
 sg13g2_decap_8 FILLER_42_637 ();
 sg13g2_decap_8 FILLER_42_644 ();
 sg13g2_decap_8 FILLER_42_651 ();
 sg13g2_decap_8 FILLER_42_658 ();
 sg13g2_decap_8 FILLER_42_665 ();
 sg13g2_decap_8 FILLER_42_672 ();
 sg13g2_decap_8 FILLER_42_679 ();
 sg13g2_decap_8 FILLER_42_686 ();
 sg13g2_decap_8 FILLER_42_693 ();
 sg13g2_decap_8 FILLER_42_700 ();
 sg13g2_decap_8 FILLER_42_707 ();
 sg13g2_decap_8 FILLER_42_714 ();
 sg13g2_decap_8 FILLER_42_721 ();
 sg13g2_decap_8 FILLER_42_728 ();
 sg13g2_decap_8 FILLER_42_735 ();
 sg13g2_decap_8 FILLER_42_742 ();
 sg13g2_decap_8 FILLER_42_749 ();
 sg13g2_decap_8 FILLER_42_756 ();
 sg13g2_decap_8 FILLER_42_763 ();
 sg13g2_decap_8 FILLER_42_770 ();
 sg13g2_decap_8 FILLER_42_777 ();
 sg13g2_decap_8 FILLER_42_784 ();
 sg13g2_decap_8 FILLER_42_791 ();
 sg13g2_decap_8 FILLER_42_798 ();
 sg13g2_decap_8 FILLER_42_805 ();
 sg13g2_decap_8 FILLER_42_812 ();
 sg13g2_decap_8 FILLER_42_819 ();
 sg13g2_decap_8 FILLER_42_826 ();
 sg13g2_decap_8 FILLER_42_833 ();
 sg13g2_decap_8 FILLER_42_840 ();
 sg13g2_decap_8 FILLER_42_847 ();
 sg13g2_decap_8 FILLER_42_854 ();
 sg13g2_decap_8 FILLER_42_861 ();
 sg13g2_decap_8 FILLER_42_868 ();
 sg13g2_decap_8 FILLER_42_875 ();
 sg13g2_decap_8 FILLER_42_882 ();
 sg13g2_decap_8 FILLER_42_889 ();
 sg13g2_decap_8 FILLER_42_896 ();
 sg13g2_decap_8 FILLER_42_903 ();
 sg13g2_decap_8 FILLER_42_910 ();
 sg13g2_decap_8 FILLER_42_917 ();
 sg13g2_decap_8 FILLER_42_924 ();
 sg13g2_decap_8 FILLER_42_931 ();
 sg13g2_decap_8 FILLER_42_938 ();
 sg13g2_decap_8 FILLER_42_945 ();
 sg13g2_decap_8 FILLER_42_952 ();
 sg13g2_decap_8 FILLER_42_959 ();
 sg13g2_decap_8 FILLER_42_966 ();
 sg13g2_decap_8 FILLER_42_973 ();
 sg13g2_decap_8 FILLER_42_980 ();
 sg13g2_decap_8 FILLER_42_987 ();
 sg13g2_decap_8 FILLER_42_994 ();
 sg13g2_decap_8 FILLER_42_1001 ();
 sg13g2_decap_8 FILLER_42_1008 ();
 sg13g2_decap_8 FILLER_42_1015 ();
 sg13g2_decap_8 FILLER_42_1022 ();
 sg13g2_decap_8 FILLER_42_1029 ();
 sg13g2_decap_8 FILLER_42_1036 ();
 sg13g2_decap_8 FILLER_42_1043 ();
 sg13g2_decap_8 FILLER_42_1050 ();
 sg13g2_decap_8 FILLER_42_1057 ();
 sg13g2_decap_8 FILLER_42_1064 ();
 sg13g2_decap_8 FILLER_42_1071 ();
 sg13g2_decap_8 FILLER_42_1078 ();
 sg13g2_decap_8 FILLER_42_1085 ();
 sg13g2_decap_8 FILLER_42_1092 ();
 sg13g2_decap_8 FILLER_42_1099 ();
 sg13g2_decap_8 FILLER_42_1106 ();
 sg13g2_decap_8 FILLER_42_1113 ();
 sg13g2_decap_8 FILLER_42_1120 ();
 sg13g2_decap_8 FILLER_42_1127 ();
 sg13g2_decap_8 FILLER_42_1134 ();
 sg13g2_decap_8 FILLER_42_1141 ();
 sg13g2_decap_8 FILLER_42_1148 ();
 sg13g2_decap_8 FILLER_42_1155 ();
 sg13g2_decap_8 FILLER_42_1162 ();
 sg13g2_decap_8 FILLER_42_1169 ();
 sg13g2_decap_8 FILLER_42_1176 ();
 sg13g2_decap_8 FILLER_42_1183 ();
 sg13g2_decap_8 FILLER_42_1190 ();
 sg13g2_decap_8 FILLER_42_1197 ();
 sg13g2_decap_8 FILLER_42_1204 ();
 sg13g2_decap_8 FILLER_42_1211 ();
 sg13g2_decap_8 FILLER_42_1218 ();
 sg13g2_decap_8 FILLER_42_1225 ();
 sg13g2_decap_8 FILLER_42_1232 ();
 sg13g2_decap_8 FILLER_42_1239 ();
 sg13g2_decap_8 FILLER_42_1246 ();
 sg13g2_decap_8 FILLER_42_1253 ();
 sg13g2_decap_8 FILLER_42_1260 ();
 sg13g2_decap_8 FILLER_42_1267 ();
 sg13g2_decap_8 FILLER_42_1274 ();
 sg13g2_decap_8 FILLER_42_1281 ();
 sg13g2_decap_8 FILLER_42_1288 ();
 sg13g2_decap_8 FILLER_42_1295 ();
 sg13g2_decap_8 FILLER_42_1302 ();
 sg13g2_decap_8 FILLER_42_1309 ();
 sg13g2_decap_8 FILLER_42_1316 ();
 sg13g2_decap_8 FILLER_42_1323 ();
 sg13g2_decap_8 FILLER_42_1330 ();
 sg13g2_decap_8 FILLER_42_1337 ();
 sg13g2_decap_8 FILLER_42_1344 ();
 sg13g2_decap_8 FILLER_42_1351 ();
 sg13g2_decap_8 FILLER_42_1358 ();
 sg13g2_decap_8 FILLER_42_1365 ();
 sg13g2_decap_8 FILLER_42_1372 ();
 sg13g2_decap_8 FILLER_42_1379 ();
 sg13g2_decap_8 FILLER_42_1386 ();
 sg13g2_decap_8 FILLER_42_1393 ();
 sg13g2_decap_8 FILLER_42_1400 ();
 sg13g2_decap_8 FILLER_42_1407 ();
 sg13g2_decap_8 FILLER_42_1414 ();
 sg13g2_decap_8 FILLER_42_1421 ();
 sg13g2_decap_8 FILLER_42_1428 ();
 sg13g2_decap_8 FILLER_42_1435 ();
 sg13g2_decap_8 FILLER_42_1442 ();
 sg13g2_decap_8 FILLER_42_1449 ();
 sg13g2_decap_8 FILLER_42_1456 ();
 sg13g2_decap_8 FILLER_42_1463 ();
 sg13g2_decap_8 FILLER_42_1470 ();
 sg13g2_decap_8 FILLER_42_1477 ();
 sg13g2_decap_8 FILLER_42_1484 ();
 sg13g2_decap_8 FILLER_42_1491 ();
 sg13g2_decap_8 FILLER_42_1498 ();
 sg13g2_decap_8 FILLER_42_1505 ();
 sg13g2_decap_8 FILLER_42_1512 ();
 sg13g2_decap_8 FILLER_42_1519 ();
 sg13g2_decap_8 FILLER_42_1526 ();
 sg13g2_decap_8 FILLER_42_1533 ();
 sg13g2_decap_8 FILLER_42_1540 ();
 sg13g2_decap_8 FILLER_42_1547 ();
 sg13g2_decap_8 FILLER_42_1554 ();
 sg13g2_decap_8 FILLER_42_1561 ();
 sg13g2_decap_8 FILLER_42_1568 ();
 sg13g2_decap_8 FILLER_42_1575 ();
 sg13g2_decap_8 FILLER_42_1582 ();
 sg13g2_decap_8 FILLER_42_1589 ();
 sg13g2_decap_8 FILLER_42_1596 ();
 sg13g2_decap_8 FILLER_42_1603 ();
 sg13g2_decap_8 FILLER_42_1610 ();
 sg13g2_decap_8 FILLER_42_1617 ();
 sg13g2_decap_8 FILLER_42_1624 ();
 sg13g2_decap_8 FILLER_42_1631 ();
 sg13g2_decap_8 FILLER_42_1638 ();
 sg13g2_decap_8 FILLER_42_1645 ();
 sg13g2_decap_8 FILLER_42_1652 ();
 sg13g2_decap_8 FILLER_42_1659 ();
 sg13g2_decap_8 FILLER_42_1666 ();
 sg13g2_decap_8 FILLER_42_1673 ();
 sg13g2_decap_8 FILLER_42_1680 ();
 sg13g2_decap_8 FILLER_42_1687 ();
 sg13g2_decap_8 FILLER_42_1694 ();
 sg13g2_decap_8 FILLER_42_1701 ();
 sg13g2_decap_8 FILLER_42_1708 ();
 sg13g2_decap_8 FILLER_42_1715 ();
 sg13g2_decap_8 FILLER_42_1722 ();
 sg13g2_decap_8 FILLER_42_1729 ();
 sg13g2_decap_8 FILLER_42_1736 ();
 sg13g2_decap_8 FILLER_42_1743 ();
 sg13g2_decap_8 FILLER_42_1750 ();
 sg13g2_decap_8 FILLER_42_1757 ();
 sg13g2_decap_8 FILLER_42_1764 ();
 sg13g2_decap_8 FILLER_42_1771 ();
 sg13g2_decap_8 FILLER_42_1778 ();
 sg13g2_decap_8 FILLER_42_1785 ();
 sg13g2_decap_8 FILLER_42_1792 ();
 sg13g2_decap_8 FILLER_42_1799 ();
 sg13g2_decap_8 FILLER_42_1806 ();
 sg13g2_decap_8 FILLER_42_1813 ();
 sg13g2_decap_8 FILLER_42_1820 ();
 sg13g2_decap_8 FILLER_42_1827 ();
 sg13g2_decap_8 FILLER_42_1834 ();
 sg13g2_decap_8 FILLER_42_1841 ();
 sg13g2_decap_8 FILLER_42_1848 ();
 sg13g2_decap_8 FILLER_42_1855 ();
 sg13g2_decap_8 FILLER_42_1862 ();
 sg13g2_decap_8 FILLER_42_1869 ();
 sg13g2_decap_8 FILLER_42_1876 ();
 sg13g2_decap_8 FILLER_42_1883 ();
 sg13g2_decap_8 FILLER_42_1890 ();
 sg13g2_decap_8 FILLER_42_1897 ();
 sg13g2_decap_8 FILLER_42_1904 ();
 sg13g2_decap_8 FILLER_42_1911 ();
 sg13g2_decap_8 FILLER_42_1918 ();
 sg13g2_decap_8 FILLER_42_1925 ();
 sg13g2_decap_8 FILLER_42_1932 ();
 sg13g2_decap_8 FILLER_42_1939 ();
 sg13g2_decap_8 FILLER_42_1946 ();
 sg13g2_decap_8 FILLER_42_1953 ();
 sg13g2_decap_8 FILLER_42_1960 ();
 sg13g2_decap_8 FILLER_42_1967 ();
 sg13g2_decap_8 FILLER_42_1974 ();
 sg13g2_decap_8 FILLER_42_1981 ();
 sg13g2_decap_8 FILLER_42_1988 ();
 sg13g2_decap_8 FILLER_42_1995 ();
 sg13g2_decap_8 FILLER_42_2002 ();
 sg13g2_decap_8 FILLER_42_2009 ();
 sg13g2_decap_8 FILLER_42_2016 ();
 sg13g2_decap_8 FILLER_42_2023 ();
 sg13g2_decap_8 FILLER_42_2030 ();
 sg13g2_decap_8 FILLER_42_2037 ();
 sg13g2_decap_8 FILLER_42_2044 ();
 sg13g2_decap_8 FILLER_42_2051 ();
 sg13g2_decap_8 FILLER_42_2058 ();
 sg13g2_decap_8 FILLER_42_2065 ();
 sg13g2_decap_8 FILLER_42_2072 ();
 sg13g2_decap_8 FILLER_42_2079 ();
 sg13g2_decap_8 FILLER_42_2086 ();
 sg13g2_decap_8 FILLER_42_2093 ();
 sg13g2_decap_8 FILLER_42_2100 ();
 sg13g2_decap_8 FILLER_42_2107 ();
 sg13g2_decap_8 FILLER_42_2114 ();
 sg13g2_decap_8 FILLER_42_2121 ();
 sg13g2_decap_8 FILLER_42_2128 ();
 sg13g2_decap_8 FILLER_42_2135 ();
 sg13g2_decap_8 FILLER_42_2142 ();
 sg13g2_decap_8 FILLER_42_2149 ();
 sg13g2_decap_8 FILLER_42_2156 ();
 sg13g2_decap_8 FILLER_42_2163 ();
 sg13g2_decap_8 FILLER_42_2170 ();
 sg13g2_decap_8 FILLER_42_2177 ();
 sg13g2_decap_8 FILLER_42_2184 ();
 sg13g2_decap_8 FILLER_42_2191 ();
 sg13g2_decap_8 FILLER_42_2198 ();
 sg13g2_decap_8 FILLER_42_2205 ();
 sg13g2_decap_8 FILLER_42_2212 ();
 sg13g2_decap_8 FILLER_42_2219 ();
 sg13g2_decap_8 FILLER_42_2226 ();
 sg13g2_decap_8 FILLER_42_2233 ();
 sg13g2_decap_8 FILLER_42_2240 ();
 sg13g2_decap_8 FILLER_42_2247 ();
 sg13g2_decap_8 FILLER_42_2254 ();
 sg13g2_decap_8 FILLER_42_2261 ();
 sg13g2_decap_8 FILLER_42_2268 ();
 sg13g2_decap_8 FILLER_42_2275 ();
 sg13g2_decap_8 FILLER_42_2282 ();
 sg13g2_decap_8 FILLER_42_2289 ();
 sg13g2_decap_8 FILLER_42_2296 ();
 sg13g2_decap_8 FILLER_42_2303 ();
 sg13g2_decap_8 FILLER_42_2310 ();
 sg13g2_decap_8 FILLER_42_2317 ();
 sg13g2_decap_8 FILLER_42_2324 ();
 sg13g2_decap_8 FILLER_42_2331 ();
 sg13g2_decap_8 FILLER_42_2338 ();
 sg13g2_decap_8 FILLER_42_2345 ();
 sg13g2_decap_8 FILLER_42_2352 ();
 sg13g2_decap_8 FILLER_42_2359 ();
 sg13g2_decap_8 FILLER_42_2366 ();
 sg13g2_decap_8 FILLER_42_2373 ();
 sg13g2_decap_8 FILLER_42_2380 ();
 sg13g2_decap_8 FILLER_42_2387 ();
 sg13g2_decap_8 FILLER_42_2394 ();
 sg13g2_decap_8 FILLER_42_2401 ();
 sg13g2_decap_8 FILLER_42_2408 ();
 sg13g2_decap_8 FILLER_42_2415 ();
 sg13g2_decap_8 FILLER_42_2422 ();
 sg13g2_decap_8 FILLER_42_2429 ();
 sg13g2_decap_8 FILLER_42_2436 ();
 sg13g2_decap_8 FILLER_42_2443 ();
 sg13g2_decap_8 FILLER_42_2450 ();
 sg13g2_decap_8 FILLER_42_2457 ();
 sg13g2_decap_8 FILLER_42_2464 ();
 sg13g2_decap_8 FILLER_42_2471 ();
 sg13g2_decap_8 FILLER_42_2478 ();
 sg13g2_decap_8 FILLER_42_2485 ();
 sg13g2_decap_8 FILLER_42_2492 ();
 sg13g2_decap_8 FILLER_42_2499 ();
 sg13g2_decap_8 FILLER_42_2506 ();
 sg13g2_decap_8 FILLER_42_2513 ();
 sg13g2_decap_8 FILLER_42_2520 ();
 sg13g2_decap_8 FILLER_42_2527 ();
 sg13g2_decap_8 FILLER_42_2534 ();
 sg13g2_decap_8 FILLER_42_2541 ();
 sg13g2_decap_8 FILLER_42_2548 ();
 sg13g2_decap_8 FILLER_42_2555 ();
 sg13g2_decap_8 FILLER_42_2562 ();
 sg13g2_decap_8 FILLER_42_2569 ();
 sg13g2_decap_8 FILLER_42_2576 ();
 sg13g2_decap_8 FILLER_42_2583 ();
 sg13g2_decap_8 FILLER_42_2590 ();
 sg13g2_decap_8 FILLER_42_2597 ();
 sg13g2_decap_8 FILLER_42_2604 ();
 sg13g2_decap_8 FILLER_42_2611 ();
 sg13g2_decap_8 FILLER_42_2618 ();
 sg13g2_decap_8 FILLER_42_2625 ();
 sg13g2_decap_8 FILLER_42_2632 ();
 sg13g2_decap_8 FILLER_42_2639 ();
 sg13g2_decap_8 FILLER_42_2646 ();
 sg13g2_decap_8 FILLER_42_2653 ();
 sg13g2_decap_8 FILLER_42_2660 ();
 sg13g2_decap_8 FILLER_42_2667 ();
 sg13g2_decap_8 FILLER_42_2674 ();
 sg13g2_decap_8 FILLER_42_2681 ();
 sg13g2_decap_8 FILLER_42_2688 ();
 sg13g2_decap_8 FILLER_42_2695 ();
 sg13g2_decap_8 FILLER_42_2702 ();
 sg13g2_decap_8 FILLER_42_2709 ();
 sg13g2_decap_8 FILLER_42_2716 ();
 sg13g2_decap_8 FILLER_42_2723 ();
 sg13g2_decap_8 FILLER_42_2730 ();
 sg13g2_decap_8 FILLER_42_2737 ();
 sg13g2_decap_8 FILLER_42_2744 ();
 sg13g2_decap_8 FILLER_42_2751 ();
 sg13g2_decap_8 FILLER_42_2758 ();
 sg13g2_decap_8 FILLER_42_2765 ();
 sg13g2_decap_8 FILLER_42_2772 ();
 sg13g2_decap_8 FILLER_42_2779 ();
 sg13g2_decap_8 FILLER_42_2786 ();
 sg13g2_decap_8 FILLER_42_2793 ();
 sg13g2_decap_8 FILLER_42_2800 ();
 sg13g2_decap_8 FILLER_42_2807 ();
 sg13g2_decap_8 FILLER_42_2814 ();
 sg13g2_decap_8 FILLER_42_2821 ();
 sg13g2_decap_8 FILLER_42_2828 ();
 sg13g2_decap_8 FILLER_42_2835 ();
 sg13g2_decap_8 FILLER_42_2842 ();
 sg13g2_decap_8 FILLER_42_2849 ();
 sg13g2_decap_8 FILLER_42_2856 ();
 sg13g2_decap_8 FILLER_42_2863 ();
 sg13g2_decap_8 FILLER_42_2870 ();
 sg13g2_decap_8 FILLER_42_2877 ();
 sg13g2_decap_8 FILLER_42_2884 ();
 sg13g2_decap_8 FILLER_42_2891 ();
 sg13g2_decap_8 FILLER_42_2898 ();
 sg13g2_decap_8 FILLER_42_2905 ();
 sg13g2_decap_8 FILLER_42_2912 ();
 sg13g2_decap_8 FILLER_42_2919 ();
 sg13g2_decap_8 FILLER_42_2926 ();
 sg13g2_decap_8 FILLER_42_2933 ();
 sg13g2_decap_8 FILLER_42_2940 ();
 sg13g2_decap_8 FILLER_42_2947 ();
 sg13g2_decap_8 FILLER_42_2954 ();
 sg13g2_decap_8 FILLER_42_2961 ();
 sg13g2_decap_8 FILLER_42_2968 ();
 sg13g2_decap_8 FILLER_42_2975 ();
 sg13g2_decap_8 FILLER_42_2982 ();
 sg13g2_decap_8 FILLER_42_2989 ();
 sg13g2_decap_8 FILLER_42_2996 ();
 sg13g2_decap_8 FILLER_42_3003 ();
 sg13g2_decap_8 FILLER_42_3010 ();
 sg13g2_decap_8 FILLER_42_3017 ();
 sg13g2_decap_8 FILLER_42_3024 ();
 sg13g2_decap_8 FILLER_42_3031 ();
 sg13g2_decap_8 FILLER_42_3038 ();
 sg13g2_decap_8 FILLER_42_3045 ();
 sg13g2_decap_8 FILLER_42_3052 ();
 sg13g2_decap_8 FILLER_42_3059 ();
 sg13g2_decap_8 FILLER_42_3066 ();
 sg13g2_decap_8 FILLER_42_3073 ();
 sg13g2_decap_8 FILLER_42_3080 ();
 sg13g2_decap_8 FILLER_42_3087 ();
 sg13g2_decap_8 FILLER_42_3094 ();
 sg13g2_decap_8 FILLER_42_3101 ();
 sg13g2_decap_8 FILLER_42_3108 ();
 sg13g2_decap_8 FILLER_42_3115 ();
 sg13g2_decap_8 FILLER_42_3122 ();
 sg13g2_decap_8 FILLER_42_3129 ();
 sg13g2_decap_8 FILLER_42_3136 ();
 sg13g2_decap_8 FILLER_42_3143 ();
 sg13g2_decap_8 FILLER_42_3150 ();
 sg13g2_decap_8 FILLER_42_3157 ();
 sg13g2_decap_8 FILLER_42_3164 ();
 sg13g2_decap_8 FILLER_42_3171 ();
 sg13g2_decap_8 FILLER_42_3178 ();
 sg13g2_decap_8 FILLER_42_3185 ();
 sg13g2_decap_8 FILLER_42_3192 ();
 sg13g2_decap_8 FILLER_42_3199 ();
 sg13g2_decap_8 FILLER_42_3206 ();
 sg13g2_decap_8 FILLER_42_3213 ();
 sg13g2_decap_8 FILLER_42_3220 ();
 sg13g2_decap_8 FILLER_42_3227 ();
 sg13g2_decap_8 FILLER_42_3234 ();
 sg13g2_decap_8 FILLER_42_3241 ();
 sg13g2_decap_8 FILLER_42_3248 ();
 sg13g2_decap_8 FILLER_42_3255 ();
 sg13g2_decap_8 FILLER_42_3262 ();
 sg13g2_decap_8 FILLER_42_3269 ();
 sg13g2_decap_8 FILLER_42_3276 ();
 sg13g2_decap_8 FILLER_42_3283 ();
 sg13g2_decap_8 FILLER_42_3290 ();
 sg13g2_decap_8 FILLER_42_3297 ();
 sg13g2_decap_8 FILLER_42_3304 ();
 sg13g2_decap_8 FILLER_42_3311 ();
 sg13g2_decap_8 FILLER_42_3318 ();
 sg13g2_decap_8 FILLER_42_3325 ();
 sg13g2_decap_8 FILLER_42_3332 ();
 sg13g2_decap_8 FILLER_42_3339 ();
 sg13g2_decap_8 FILLER_42_3346 ();
 sg13g2_decap_8 FILLER_42_3353 ();
 sg13g2_decap_8 FILLER_42_3360 ();
 sg13g2_decap_8 FILLER_42_3367 ();
 sg13g2_decap_8 FILLER_42_3374 ();
 sg13g2_decap_8 FILLER_42_3381 ();
 sg13g2_decap_8 FILLER_42_3388 ();
 sg13g2_decap_8 FILLER_42_3395 ();
 sg13g2_decap_8 FILLER_42_3402 ();
 sg13g2_decap_8 FILLER_42_3409 ();
 sg13g2_decap_8 FILLER_42_3416 ();
 sg13g2_decap_8 FILLER_42_3423 ();
 sg13g2_decap_8 FILLER_42_3430 ();
 sg13g2_decap_8 FILLER_42_3437 ();
 sg13g2_decap_8 FILLER_42_3444 ();
 sg13g2_decap_8 FILLER_42_3451 ();
 sg13g2_decap_8 FILLER_42_3458 ();
 sg13g2_decap_8 FILLER_42_3465 ();
 sg13g2_decap_8 FILLER_42_3472 ();
 sg13g2_decap_8 FILLER_42_3479 ();
 sg13g2_decap_8 FILLER_42_3486 ();
 sg13g2_decap_8 FILLER_42_3493 ();
 sg13g2_decap_8 FILLER_42_3500 ();
 sg13g2_decap_8 FILLER_42_3507 ();
 sg13g2_decap_8 FILLER_42_3514 ();
 sg13g2_decap_8 FILLER_42_3521 ();
 sg13g2_decap_8 FILLER_42_3528 ();
 sg13g2_decap_8 FILLER_42_3535 ();
 sg13g2_decap_8 FILLER_42_3542 ();
 sg13g2_decap_8 FILLER_42_3549 ();
 sg13g2_decap_8 FILLER_42_3556 ();
 sg13g2_decap_8 FILLER_42_3563 ();
 sg13g2_decap_8 FILLER_42_3570 ();
 sg13g2_fill_2 FILLER_42_3577 ();
 sg13g2_fill_1 FILLER_42_3579 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_decap_8 FILLER_43_133 ();
 sg13g2_decap_8 FILLER_43_140 ();
 sg13g2_decap_8 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_154 ();
 sg13g2_decap_8 FILLER_43_161 ();
 sg13g2_decap_8 FILLER_43_168 ();
 sg13g2_decap_8 FILLER_43_175 ();
 sg13g2_decap_8 FILLER_43_182 ();
 sg13g2_decap_8 FILLER_43_189 ();
 sg13g2_decap_8 FILLER_43_196 ();
 sg13g2_decap_8 FILLER_43_203 ();
 sg13g2_decap_8 FILLER_43_210 ();
 sg13g2_decap_8 FILLER_43_217 ();
 sg13g2_decap_8 FILLER_43_224 ();
 sg13g2_decap_8 FILLER_43_231 ();
 sg13g2_decap_8 FILLER_43_238 ();
 sg13g2_decap_8 FILLER_43_245 ();
 sg13g2_decap_8 FILLER_43_252 ();
 sg13g2_decap_8 FILLER_43_259 ();
 sg13g2_decap_8 FILLER_43_266 ();
 sg13g2_decap_8 FILLER_43_273 ();
 sg13g2_decap_8 FILLER_43_280 ();
 sg13g2_decap_8 FILLER_43_287 ();
 sg13g2_decap_8 FILLER_43_294 ();
 sg13g2_decap_8 FILLER_43_301 ();
 sg13g2_decap_8 FILLER_43_308 ();
 sg13g2_decap_8 FILLER_43_315 ();
 sg13g2_decap_8 FILLER_43_322 ();
 sg13g2_decap_8 FILLER_43_329 ();
 sg13g2_decap_8 FILLER_43_336 ();
 sg13g2_decap_8 FILLER_43_343 ();
 sg13g2_decap_8 FILLER_43_350 ();
 sg13g2_decap_8 FILLER_43_357 ();
 sg13g2_decap_8 FILLER_43_364 ();
 sg13g2_decap_8 FILLER_43_371 ();
 sg13g2_decap_8 FILLER_43_378 ();
 sg13g2_decap_8 FILLER_43_385 ();
 sg13g2_decap_8 FILLER_43_392 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_decap_8 FILLER_43_406 ();
 sg13g2_decap_8 FILLER_43_413 ();
 sg13g2_decap_8 FILLER_43_420 ();
 sg13g2_decap_8 FILLER_43_427 ();
 sg13g2_decap_8 FILLER_43_434 ();
 sg13g2_decap_8 FILLER_43_441 ();
 sg13g2_decap_8 FILLER_43_448 ();
 sg13g2_decap_8 FILLER_43_455 ();
 sg13g2_decap_8 FILLER_43_462 ();
 sg13g2_decap_8 FILLER_43_469 ();
 sg13g2_decap_8 FILLER_43_476 ();
 sg13g2_decap_8 FILLER_43_483 ();
 sg13g2_decap_8 FILLER_43_490 ();
 sg13g2_decap_8 FILLER_43_497 ();
 sg13g2_decap_8 FILLER_43_504 ();
 sg13g2_decap_8 FILLER_43_511 ();
 sg13g2_decap_8 FILLER_43_518 ();
 sg13g2_decap_8 FILLER_43_525 ();
 sg13g2_decap_8 FILLER_43_532 ();
 sg13g2_decap_8 FILLER_43_539 ();
 sg13g2_decap_8 FILLER_43_546 ();
 sg13g2_decap_8 FILLER_43_553 ();
 sg13g2_decap_8 FILLER_43_560 ();
 sg13g2_decap_8 FILLER_43_567 ();
 sg13g2_decap_8 FILLER_43_574 ();
 sg13g2_decap_8 FILLER_43_581 ();
 sg13g2_decap_8 FILLER_43_588 ();
 sg13g2_decap_8 FILLER_43_595 ();
 sg13g2_decap_8 FILLER_43_602 ();
 sg13g2_decap_8 FILLER_43_609 ();
 sg13g2_decap_8 FILLER_43_616 ();
 sg13g2_decap_8 FILLER_43_623 ();
 sg13g2_decap_8 FILLER_43_630 ();
 sg13g2_decap_8 FILLER_43_637 ();
 sg13g2_decap_8 FILLER_43_644 ();
 sg13g2_decap_8 FILLER_43_651 ();
 sg13g2_decap_8 FILLER_43_658 ();
 sg13g2_decap_8 FILLER_43_665 ();
 sg13g2_decap_8 FILLER_43_672 ();
 sg13g2_decap_8 FILLER_43_679 ();
 sg13g2_decap_8 FILLER_43_686 ();
 sg13g2_decap_8 FILLER_43_693 ();
 sg13g2_decap_8 FILLER_43_700 ();
 sg13g2_decap_8 FILLER_43_707 ();
 sg13g2_decap_8 FILLER_43_714 ();
 sg13g2_decap_8 FILLER_43_721 ();
 sg13g2_decap_8 FILLER_43_728 ();
 sg13g2_decap_8 FILLER_43_735 ();
 sg13g2_decap_8 FILLER_43_742 ();
 sg13g2_decap_8 FILLER_43_749 ();
 sg13g2_decap_8 FILLER_43_756 ();
 sg13g2_decap_8 FILLER_43_763 ();
 sg13g2_decap_8 FILLER_43_770 ();
 sg13g2_decap_8 FILLER_43_777 ();
 sg13g2_decap_8 FILLER_43_784 ();
 sg13g2_decap_8 FILLER_43_791 ();
 sg13g2_decap_8 FILLER_43_798 ();
 sg13g2_decap_8 FILLER_43_805 ();
 sg13g2_decap_8 FILLER_43_812 ();
 sg13g2_decap_8 FILLER_43_819 ();
 sg13g2_decap_8 FILLER_43_826 ();
 sg13g2_decap_8 FILLER_43_833 ();
 sg13g2_decap_8 FILLER_43_840 ();
 sg13g2_decap_8 FILLER_43_847 ();
 sg13g2_decap_8 FILLER_43_854 ();
 sg13g2_decap_8 FILLER_43_861 ();
 sg13g2_decap_8 FILLER_43_868 ();
 sg13g2_decap_8 FILLER_43_875 ();
 sg13g2_decap_8 FILLER_43_882 ();
 sg13g2_decap_8 FILLER_43_889 ();
 sg13g2_decap_8 FILLER_43_896 ();
 sg13g2_decap_8 FILLER_43_903 ();
 sg13g2_decap_8 FILLER_43_910 ();
 sg13g2_decap_8 FILLER_43_917 ();
 sg13g2_decap_8 FILLER_43_924 ();
 sg13g2_decap_8 FILLER_43_931 ();
 sg13g2_decap_8 FILLER_43_938 ();
 sg13g2_decap_8 FILLER_43_945 ();
 sg13g2_decap_8 FILLER_43_952 ();
 sg13g2_decap_8 FILLER_43_959 ();
 sg13g2_decap_8 FILLER_43_966 ();
 sg13g2_decap_8 FILLER_43_973 ();
 sg13g2_decap_8 FILLER_43_980 ();
 sg13g2_decap_8 FILLER_43_987 ();
 sg13g2_decap_8 FILLER_43_994 ();
 sg13g2_decap_8 FILLER_43_1001 ();
 sg13g2_decap_8 FILLER_43_1008 ();
 sg13g2_decap_8 FILLER_43_1015 ();
 sg13g2_decap_8 FILLER_43_1022 ();
 sg13g2_decap_8 FILLER_43_1029 ();
 sg13g2_decap_8 FILLER_43_1036 ();
 sg13g2_decap_8 FILLER_43_1043 ();
 sg13g2_decap_8 FILLER_43_1050 ();
 sg13g2_decap_8 FILLER_43_1057 ();
 sg13g2_decap_8 FILLER_43_1064 ();
 sg13g2_decap_8 FILLER_43_1071 ();
 sg13g2_decap_8 FILLER_43_1078 ();
 sg13g2_decap_8 FILLER_43_1085 ();
 sg13g2_decap_8 FILLER_43_1092 ();
 sg13g2_decap_8 FILLER_43_1099 ();
 sg13g2_decap_8 FILLER_43_1106 ();
 sg13g2_decap_8 FILLER_43_1113 ();
 sg13g2_decap_8 FILLER_43_1120 ();
 sg13g2_decap_8 FILLER_43_1127 ();
 sg13g2_decap_8 FILLER_43_1134 ();
 sg13g2_decap_8 FILLER_43_1141 ();
 sg13g2_decap_8 FILLER_43_1148 ();
 sg13g2_decap_8 FILLER_43_1155 ();
 sg13g2_decap_8 FILLER_43_1162 ();
 sg13g2_decap_8 FILLER_43_1169 ();
 sg13g2_decap_8 FILLER_43_1176 ();
 sg13g2_decap_8 FILLER_43_1183 ();
 sg13g2_decap_8 FILLER_43_1190 ();
 sg13g2_decap_8 FILLER_43_1197 ();
 sg13g2_decap_8 FILLER_43_1204 ();
 sg13g2_decap_8 FILLER_43_1211 ();
 sg13g2_decap_8 FILLER_43_1218 ();
 sg13g2_decap_8 FILLER_43_1225 ();
 sg13g2_decap_8 FILLER_43_1232 ();
 sg13g2_decap_8 FILLER_43_1239 ();
 sg13g2_decap_8 FILLER_43_1246 ();
 sg13g2_decap_8 FILLER_43_1253 ();
 sg13g2_decap_8 FILLER_43_1260 ();
 sg13g2_decap_8 FILLER_43_1267 ();
 sg13g2_decap_8 FILLER_43_1274 ();
 sg13g2_decap_8 FILLER_43_1281 ();
 sg13g2_decap_8 FILLER_43_1288 ();
 sg13g2_decap_8 FILLER_43_1295 ();
 sg13g2_decap_8 FILLER_43_1302 ();
 sg13g2_decap_8 FILLER_43_1309 ();
 sg13g2_decap_8 FILLER_43_1316 ();
 sg13g2_decap_8 FILLER_43_1323 ();
 sg13g2_decap_8 FILLER_43_1330 ();
 sg13g2_decap_8 FILLER_43_1337 ();
 sg13g2_decap_8 FILLER_43_1344 ();
 sg13g2_decap_8 FILLER_43_1351 ();
 sg13g2_decap_8 FILLER_43_1358 ();
 sg13g2_decap_8 FILLER_43_1365 ();
 sg13g2_decap_8 FILLER_43_1372 ();
 sg13g2_decap_8 FILLER_43_1379 ();
 sg13g2_decap_8 FILLER_43_1386 ();
 sg13g2_decap_8 FILLER_43_1393 ();
 sg13g2_decap_8 FILLER_43_1400 ();
 sg13g2_decap_8 FILLER_43_1407 ();
 sg13g2_decap_8 FILLER_43_1414 ();
 sg13g2_decap_8 FILLER_43_1421 ();
 sg13g2_decap_8 FILLER_43_1428 ();
 sg13g2_decap_8 FILLER_43_1435 ();
 sg13g2_decap_8 FILLER_43_1442 ();
 sg13g2_decap_8 FILLER_43_1449 ();
 sg13g2_decap_8 FILLER_43_1456 ();
 sg13g2_decap_8 FILLER_43_1463 ();
 sg13g2_decap_8 FILLER_43_1470 ();
 sg13g2_decap_8 FILLER_43_1477 ();
 sg13g2_decap_8 FILLER_43_1484 ();
 sg13g2_decap_8 FILLER_43_1491 ();
 sg13g2_decap_8 FILLER_43_1498 ();
 sg13g2_decap_8 FILLER_43_1505 ();
 sg13g2_decap_8 FILLER_43_1512 ();
 sg13g2_decap_8 FILLER_43_1519 ();
 sg13g2_decap_8 FILLER_43_1526 ();
 sg13g2_decap_8 FILLER_43_1533 ();
 sg13g2_decap_8 FILLER_43_1540 ();
 sg13g2_decap_8 FILLER_43_1547 ();
 sg13g2_decap_8 FILLER_43_1554 ();
 sg13g2_decap_8 FILLER_43_1561 ();
 sg13g2_decap_8 FILLER_43_1568 ();
 sg13g2_decap_8 FILLER_43_1575 ();
 sg13g2_decap_8 FILLER_43_1582 ();
 sg13g2_decap_8 FILLER_43_1589 ();
 sg13g2_decap_8 FILLER_43_1596 ();
 sg13g2_decap_8 FILLER_43_1603 ();
 sg13g2_decap_8 FILLER_43_1610 ();
 sg13g2_decap_8 FILLER_43_1617 ();
 sg13g2_decap_8 FILLER_43_1624 ();
 sg13g2_decap_8 FILLER_43_1631 ();
 sg13g2_decap_8 FILLER_43_1638 ();
 sg13g2_decap_8 FILLER_43_1645 ();
 sg13g2_decap_8 FILLER_43_1652 ();
 sg13g2_decap_8 FILLER_43_1659 ();
 sg13g2_decap_8 FILLER_43_1666 ();
 sg13g2_decap_8 FILLER_43_1673 ();
 sg13g2_decap_8 FILLER_43_1680 ();
 sg13g2_decap_8 FILLER_43_1687 ();
 sg13g2_decap_8 FILLER_43_1694 ();
 sg13g2_decap_8 FILLER_43_1701 ();
 sg13g2_decap_8 FILLER_43_1708 ();
 sg13g2_decap_8 FILLER_43_1715 ();
 sg13g2_decap_8 FILLER_43_1722 ();
 sg13g2_decap_8 FILLER_43_1729 ();
 sg13g2_decap_8 FILLER_43_1736 ();
 sg13g2_decap_8 FILLER_43_1743 ();
 sg13g2_decap_8 FILLER_43_1750 ();
 sg13g2_decap_8 FILLER_43_1757 ();
 sg13g2_decap_8 FILLER_43_1764 ();
 sg13g2_decap_8 FILLER_43_1771 ();
 sg13g2_decap_8 FILLER_43_1778 ();
 sg13g2_decap_8 FILLER_43_1785 ();
 sg13g2_decap_8 FILLER_43_1792 ();
 sg13g2_decap_8 FILLER_43_1799 ();
 sg13g2_decap_8 FILLER_43_1806 ();
 sg13g2_decap_8 FILLER_43_1813 ();
 sg13g2_decap_8 FILLER_43_1820 ();
 sg13g2_decap_8 FILLER_43_1827 ();
 sg13g2_decap_8 FILLER_43_1834 ();
 sg13g2_decap_8 FILLER_43_1841 ();
 sg13g2_decap_8 FILLER_43_1848 ();
 sg13g2_decap_8 FILLER_43_1855 ();
 sg13g2_decap_8 FILLER_43_1862 ();
 sg13g2_decap_8 FILLER_43_1869 ();
 sg13g2_decap_8 FILLER_43_1876 ();
 sg13g2_decap_8 FILLER_43_1883 ();
 sg13g2_decap_8 FILLER_43_1890 ();
 sg13g2_decap_8 FILLER_43_1897 ();
 sg13g2_decap_8 FILLER_43_1904 ();
 sg13g2_decap_8 FILLER_43_1911 ();
 sg13g2_decap_8 FILLER_43_1918 ();
 sg13g2_decap_8 FILLER_43_1925 ();
 sg13g2_decap_8 FILLER_43_1932 ();
 sg13g2_decap_8 FILLER_43_1939 ();
 sg13g2_decap_8 FILLER_43_1946 ();
 sg13g2_decap_8 FILLER_43_1953 ();
 sg13g2_decap_8 FILLER_43_1960 ();
 sg13g2_decap_8 FILLER_43_1967 ();
 sg13g2_decap_8 FILLER_43_1974 ();
 sg13g2_decap_8 FILLER_43_1981 ();
 sg13g2_decap_8 FILLER_43_1988 ();
 sg13g2_decap_8 FILLER_43_1995 ();
 sg13g2_decap_8 FILLER_43_2002 ();
 sg13g2_decap_8 FILLER_43_2009 ();
 sg13g2_decap_8 FILLER_43_2016 ();
 sg13g2_decap_8 FILLER_43_2023 ();
 sg13g2_decap_8 FILLER_43_2030 ();
 sg13g2_decap_8 FILLER_43_2037 ();
 sg13g2_decap_8 FILLER_43_2044 ();
 sg13g2_decap_8 FILLER_43_2051 ();
 sg13g2_decap_8 FILLER_43_2058 ();
 sg13g2_decap_8 FILLER_43_2065 ();
 sg13g2_decap_8 FILLER_43_2072 ();
 sg13g2_decap_8 FILLER_43_2079 ();
 sg13g2_decap_8 FILLER_43_2086 ();
 sg13g2_decap_8 FILLER_43_2093 ();
 sg13g2_decap_8 FILLER_43_2100 ();
 sg13g2_decap_8 FILLER_43_2107 ();
 sg13g2_decap_8 FILLER_43_2114 ();
 sg13g2_decap_8 FILLER_43_2121 ();
 sg13g2_decap_8 FILLER_43_2128 ();
 sg13g2_decap_8 FILLER_43_2135 ();
 sg13g2_decap_8 FILLER_43_2142 ();
 sg13g2_decap_8 FILLER_43_2149 ();
 sg13g2_decap_8 FILLER_43_2156 ();
 sg13g2_decap_8 FILLER_43_2163 ();
 sg13g2_decap_8 FILLER_43_2170 ();
 sg13g2_decap_8 FILLER_43_2177 ();
 sg13g2_decap_8 FILLER_43_2184 ();
 sg13g2_decap_8 FILLER_43_2191 ();
 sg13g2_decap_8 FILLER_43_2198 ();
 sg13g2_decap_8 FILLER_43_2205 ();
 sg13g2_decap_8 FILLER_43_2212 ();
 sg13g2_decap_8 FILLER_43_2219 ();
 sg13g2_decap_8 FILLER_43_2226 ();
 sg13g2_decap_8 FILLER_43_2233 ();
 sg13g2_decap_8 FILLER_43_2240 ();
 sg13g2_decap_8 FILLER_43_2247 ();
 sg13g2_decap_8 FILLER_43_2254 ();
 sg13g2_decap_8 FILLER_43_2261 ();
 sg13g2_decap_8 FILLER_43_2268 ();
 sg13g2_decap_8 FILLER_43_2275 ();
 sg13g2_decap_8 FILLER_43_2282 ();
 sg13g2_decap_8 FILLER_43_2289 ();
 sg13g2_decap_8 FILLER_43_2296 ();
 sg13g2_decap_8 FILLER_43_2303 ();
 sg13g2_decap_8 FILLER_43_2310 ();
 sg13g2_decap_8 FILLER_43_2317 ();
 sg13g2_decap_8 FILLER_43_2324 ();
 sg13g2_decap_8 FILLER_43_2331 ();
 sg13g2_decap_8 FILLER_43_2338 ();
 sg13g2_decap_8 FILLER_43_2345 ();
 sg13g2_decap_8 FILLER_43_2352 ();
 sg13g2_decap_8 FILLER_43_2359 ();
 sg13g2_decap_8 FILLER_43_2366 ();
 sg13g2_decap_8 FILLER_43_2373 ();
 sg13g2_decap_8 FILLER_43_2380 ();
 sg13g2_decap_8 FILLER_43_2387 ();
 sg13g2_decap_8 FILLER_43_2394 ();
 sg13g2_decap_8 FILLER_43_2401 ();
 sg13g2_decap_8 FILLER_43_2408 ();
 sg13g2_decap_8 FILLER_43_2415 ();
 sg13g2_decap_8 FILLER_43_2422 ();
 sg13g2_decap_8 FILLER_43_2429 ();
 sg13g2_decap_8 FILLER_43_2436 ();
 sg13g2_decap_8 FILLER_43_2443 ();
 sg13g2_decap_8 FILLER_43_2450 ();
 sg13g2_decap_8 FILLER_43_2457 ();
 sg13g2_decap_8 FILLER_43_2464 ();
 sg13g2_decap_8 FILLER_43_2471 ();
 sg13g2_decap_8 FILLER_43_2478 ();
 sg13g2_decap_8 FILLER_43_2485 ();
 sg13g2_decap_8 FILLER_43_2492 ();
 sg13g2_decap_8 FILLER_43_2499 ();
 sg13g2_decap_8 FILLER_43_2506 ();
 sg13g2_decap_8 FILLER_43_2513 ();
 sg13g2_decap_8 FILLER_43_2520 ();
 sg13g2_decap_8 FILLER_43_2527 ();
 sg13g2_decap_8 FILLER_43_2534 ();
 sg13g2_decap_8 FILLER_43_2541 ();
 sg13g2_decap_8 FILLER_43_2548 ();
 sg13g2_decap_8 FILLER_43_2555 ();
 sg13g2_decap_8 FILLER_43_2562 ();
 sg13g2_decap_8 FILLER_43_2569 ();
 sg13g2_decap_8 FILLER_43_2576 ();
 sg13g2_decap_8 FILLER_43_2583 ();
 sg13g2_decap_8 FILLER_43_2590 ();
 sg13g2_decap_8 FILLER_43_2597 ();
 sg13g2_decap_8 FILLER_43_2604 ();
 sg13g2_decap_8 FILLER_43_2611 ();
 sg13g2_decap_8 FILLER_43_2618 ();
 sg13g2_decap_8 FILLER_43_2625 ();
 sg13g2_decap_8 FILLER_43_2632 ();
 sg13g2_decap_8 FILLER_43_2639 ();
 sg13g2_decap_8 FILLER_43_2646 ();
 sg13g2_decap_8 FILLER_43_2653 ();
 sg13g2_decap_8 FILLER_43_2660 ();
 sg13g2_decap_8 FILLER_43_2667 ();
 sg13g2_decap_8 FILLER_43_2674 ();
 sg13g2_decap_8 FILLER_43_2681 ();
 sg13g2_decap_8 FILLER_43_2688 ();
 sg13g2_decap_8 FILLER_43_2695 ();
 sg13g2_decap_8 FILLER_43_2702 ();
 sg13g2_decap_8 FILLER_43_2709 ();
 sg13g2_decap_8 FILLER_43_2716 ();
 sg13g2_decap_8 FILLER_43_2723 ();
 sg13g2_decap_8 FILLER_43_2730 ();
 sg13g2_decap_8 FILLER_43_2737 ();
 sg13g2_decap_8 FILLER_43_2744 ();
 sg13g2_decap_8 FILLER_43_2751 ();
 sg13g2_decap_8 FILLER_43_2758 ();
 sg13g2_decap_8 FILLER_43_2765 ();
 sg13g2_decap_8 FILLER_43_2772 ();
 sg13g2_decap_8 FILLER_43_2779 ();
 sg13g2_decap_8 FILLER_43_2786 ();
 sg13g2_decap_8 FILLER_43_2793 ();
 sg13g2_decap_8 FILLER_43_2800 ();
 sg13g2_decap_8 FILLER_43_2807 ();
 sg13g2_decap_8 FILLER_43_2814 ();
 sg13g2_decap_8 FILLER_43_2821 ();
 sg13g2_decap_8 FILLER_43_2828 ();
 sg13g2_decap_8 FILLER_43_2835 ();
 sg13g2_decap_8 FILLER_43_2842 ();
 sg13g2_decap_8 FILLER_43_2849 ();
 sg13g2_decap_8 FILLER_43_2856 ();
 sg13g2_decap_8 FILLER_43_2863 ();
 sg13g2_decap_8 FILLER_43_2870 ();
 sg13g2_decap_8 FILLER_43_2877 ();
 sg13g2_decap_8 FILLER_43_2884 ();
 sg13g2_decap_8 FILLER_43_2891 ();
 sg13g2_decap_8 FILLER_43_2898 ();
 sg13g2_decap_8 FILLER_43_2905 ();
 sg13g2_decap_8 FILLER_43_2912 ();
 sg13g2_decap_8 FILLER_43_2919 ();
 sg13g2_decap_8 FILLER_43_2926 ();
 sg13g2_decap_8 FILLER_43_2933 ();
 sg13g2_decap_8 FILLER_43_2940 ();
 sg13g2_decap_8 FILLER_43_2947 ();
 sg13g2_decap_8 FILLER_43_2954 ();
 sg13g2_decap_8 FILLER_43_2961 ();
 sg13g2_decap_8 FILLER_43_2968 ();
 sg13g2_decap_8 FILLER_43_2975 ();
 sg13g2_decap_8 FILLER_43_2982 ();
 sg13g2_decap_8 FILLER_43_2989 ();
 sg13g2_decap_8 FILLER_43_2996 ();
 sg13g2_decap_8 FILLER_43_3003 ();
 sg13g2_decap_8 FILLER_43_3010 ();
 sg13g2_decap_8 FILLER_43_3017 ();
 sg13g2_decap_8 FILLER_43_3024 ();
 sg13g2_decap_8 FILLER_43_3031 ();
 sg13g2_decap_8 FILLER_43_3038 ();
 sg13g2_decap_8 FILLER_43_3045 ();
 sg13g2_decap_8 FILLER_43_3052 ();
 sg13g2_decap_8 FILLER_43_3059 ();
 sg13g2_decap_8 FILLER_43_3066 ();
 sg13g2_decap_8 FILLER_43_3073 ();
 sg13g2_decap_8 FILLER_43_3080 ();
 sg13g2_decap_8 FILLER_43_3087 ();
 sg13g2_decap_8 FILLER_43_3094 ();
 sg13g2_decap_8 FILLER_43_3101 ();
 sg13g2_decap_8 FILLER_43_3108 ();
 sg13g2_decap_8 FILLER_43_3115 ();
 sg13g2_decap_8 FILLER_43_3122 ();
 sg13g2_decap_8 FILLER_43_3129 ();
 sg13g2_decap_8 FILLER_43_3136 ();
 sg13g2_decap_8 FILLER_43_3143 ();
 sg13g2_decap_8 FILLER_43_3150 ();
 sg13g2_decap_8 FILLER_43_3157 ();
 sg13g2_decap_8 FILLER_43_3164 ();
 sg13g2_decap_8 FILLER_43_3171 ();
 sg13g2_decap_8 FILLER_43_3178 ();
 sg13g2_decap_8 FILLER_43_3185 ();
 sg13g2_decap_8 FILLER_43_3192 ();
 sg13g2_decap_8 FILLER_43_3199 ();
 sg13g2_decap_8 FILLER_43_3206 ();
 sg13g2_decap_8 FILLER_43_3213 ();
 sg13g2_decap_8 FILLER_43_3220 ();
 sg13g2_decap_8 FILLER_43_3227 ();
 sg13g2_decap_8 FILLER_43_3234 ();
 sg13g2_decap_8 FILLER_43_3241 ();
 sg13g2_decap_8 FILLER_43_3248 ();
 sg13g2_decap_8 FILLER_43_3255 ();
 sg13g2_decap_8 FILLER_43_3262 ();
 sg13g2_decap_8 FILLER_43_3269 ();
 sg13g2_decap_8 FILLER_43_3276 ();
 sg13g2_decap_8 FILLER_43_3283 ();
 sg13g2_decap_8 FILLER_43_3290 ();
 sg13g2_decap_8 FILLER_43_3297 ();
 sg13g2_decap_8 FILLER_43_3304 ();
 sg13g2_decap_8 FILLER_43_3311 ();
 sg13g2_decap_8 FILLER_43_3318 ();
 sg13g2_decap_8 FILLER_43_3325 ();
 sg13g2_decap_8 FILLER_43_3332 ();
 sg13g2_decap_8 FILLER_43_3339 ();
 sg13g2_decap_8 FILLER_43_3346 ();
 sg13g2_decap_8 FILLER_43_3353 ();
 sg13g2_decap_8 FILLER_43_3360 ();
 sg13g2_decap_8 FILLER_43_3367 ();
 sg13g2_decap_8 FILLER_43_3374 ();
 sg13g2_decap_8 FILLER_43_3381 ();
 sg13g2_decap_8 FILLER_43_3388 ();
 sg13g2_decap_8 FILLER_43_3395 ();
 sg13g2_decap_8 FILLER_43_3402 ();
 sg13g2_decap_8 FILLER_43_3409 ();
 sg13g2_decap_8 FILLER_43_3416 ();
 sg13g2_decap_8 FILLER_43_3423 ();
 sg13g2_decap_8 FILLER_43_3430 ();
 sg13g2_decap_8 FILLER_43_3437 ();
 sg13g2_decap_8 FILLER_43_3444 ();
 sg13g2_decap_8 FILLER_43_3451 ();
 sg13g2_decap_8 FILLER_43_3458 ();
 sg13g2_decap_8 FILLER_43_3465 ();
 sg13g2_decap_8 FILLER_43_3472 ();
 sg13g2_decap_8 FILLER_43_3479 ();
 sg13g2_decap_8 FILLER_43_3486 ();
 sg13g2_decap_8 FILLER_43_3493 ();
 sg13g2_decap_8 FILLER_43_3500 ();
 sg13g2_decap_8 FILLER_43_3507 ();
 sg13g2_decap_8 FILLER_43_3514 ();
 sg13g2_decap_8 FILLER_43_3521 ();
 sg13g2_decap_8 FILLER_43_3528 ();
 sg13g2_decap_8 FILLER_43_3535 ();
 sg13g2_decap_8 FILLER_43_3542 ();
 sg13g2_decap_8 FILLER_43_3549 ();
 sg13g2_decap_8 FILLER_43_3556 ();
 sg13g2_decap_8 FILLER_43_3563 ();
 sg13g2_decap_8 FILLER_43_3570 ();
 sg13g2_fill_2 FILLER_43_3577 ();
 sg13g2_fill_1 FILLER_43_3579 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_decap_8 FILLER_44_133 ();
 sg13g2_decap_8 FILLER_44_140 ();
 sg13g2_decap_8 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_154 ();
 sg13g2_decap_8 FILLER_44_161 ();
 sg13g2_decap_8 FILLER_44_168 ();
 sg13g2_decap_8 FILLER_44_175 ();
 sg13g2_decap_8 FILLER_44_182 ();
 sg13g2_decap_8 FILLER_44_189 ();
 sg13g2_decap_8 FILLER_44_196 ();
 sg13g2_decap_8 FILLER_44_203 ();
 sg13g2_decap_8 FILLER_44_210 ();
 sg13g2_decap_8 FILLER_44_217 ();
 sg13g2_decap_8 FILLER_44_224 ();
 sg13g2_decap_8 FILLER_44_231 ();
 sg13g2_decap_8 FILLER_44_238 ();
 sg13g2_decap_8 FILLER_44_245 ();
 sg13g2_decap_8 FILLER_44_252 ();
 sg13g2_decap_8 FILLER_44_259 ();
 sg13g2_decap_8 FILLER_44_266 ();
 sg13g2_decap_8 FILLER_44_273 ();
 sg13g2_decap_8 FILLER_44_280 ();
 sg13g2_decap_8 FILLER_44_287 ();
 sg13g2_decap_8 FILLER_44_294 ();
 sg13g2_decap_8 FILLER_44_301 ();
 sg13g2_decap_8 FILLER_44_308 ();
 sg13g2_decap_8 FILLER_44_315 ();
 sg13g2_decap_8 FILLER_44_322 ();
 sg13g2_decap_8 FILLER_44_329 ();
 sg13g2_decap_8 FILLER_44_336 ();
 sg13g2_decap_8 FILLER_44_343 ();
 sg13g2_decap_8 FILLER_44_350 ();
 sg13g2_decap_8 FILLER_44_357 ();
 sg13g2_decap_8 FILLER_44_364 ();
 sg13g2_decap_8 FILLER_44_371 ();
 sg13g2_decap_8 FILLER_44_378 ();
 sg13g2_decap_8 FILLER_44_385 ();
 sg13g2_decap_8 FILLER_44_392 ();
 sg13g2_decap_8 FILLER_44_399 ();
 sg13g2_decap_8 FILLER_44_406 ();
 sg13g2_decap_8 FILLER_44_413 ();
 sg13g2_decap_8 FILLER_44_420 ();
 sg13g2_decap_8 FILLER_44_427 ();
 sg13g2_decap_8 FILLER_44_434 ();
 sg13g2_decap_8 FILLER_44_441 ();
 sg13g2_decap_8 FILLER_44_448 ();
 sg13g2_decap_8 FILLER_44_455 ();
 sg13g2_decap_8 FILLER_44_462 ();
 sg13g2_decap_8 FILLER_44_469 ();
 sg13g2_decap_8 FILLER_44_476 ();
 sg13g2_decap_8 FILLER_44_483 ();
 sg13g2_decap_8 FILLER_44_490 ();
 sg13g2_decap_8 FILLER_44_497 ();
 sg13g2_decap_8 FILLER_44_504 ();
 sg13g2_decap_8 FILLER_44_511 ();
 sg13g2_decap_8 FILLER_44_518 ();
 sg13g2_decap_8 FILLER_44_525 ();
 sg13g2_decap_8 FILLER_44_532 ();
 sg13g2_decap_8 FILLER_44_539 ();
 sg13g2_decap_8 FILLER_44_546 ();
 sg13g2_decap_8 FILLER_44_553 ();
 sg13g2_decap_8 FILLER_44_560 ();
 sg13g2_decap_8 FILLER_44_567 ();
 sg13g2_decap_8 FILLER_44_574 ();
 sg13g2_decap_8 FILLER_44_581 ();
 sg13g2_decap_8 FILLER_44_588 ();
 sg13g2_decap_8 FILLER_44_595 ();
 sg13g2_decap_8 FILLER_44_602 ();
 sg13g2_decap_8 FILLER_44_609 ();
 sg13g2_decap_8 FILLER_44_616 ();
 sg13g2_decap_8 FILLER_44_623 ();
 sg13g2_decap_8 FILLER_44_630 ();
 sg13g2_decap_8 FILLER_44_637 ();
 sg13g2_decap_8 FILLER_44_644 ();
 sg13g2_decap_8 FILLER_44_651 ();
 sg13g2_decap_8 FILLER_44_658 ();
 sg13g2_decap_8 FILLER_44_665 ();
 sg13g2_decap_8 FILLER_44_672 ();
 sg13g2_decap_8 FILLER_44_679 ();
 sg13g2_decap_8 FILLER_44_686 ();
 sg13g2_decap_8 FILLER_44_693 ();
 sg13g2_decap_8 FILLER_44_700 ();
 sg13g2_decap_8 FILLER_44_707 ();
 sg13g2_decap_8 FILLER_44_714 ();
 sg13g2_decap_8 FILLER_44_721 ();
 sg13g2_decap_8 FILLER_44_728 ();
 sg13g2_decap_8 FILLER_44_735 ();
 sg13g2_decap_8 FILLER_44_742 ();
 sg13g2_decap_8 FILLER_44_749 ();
 sg13g2_decap_8 FILLER_44_756 ();
 sg13g2_decap_8 FILLER_44_763 ();
 sg13g2_decap_8 FILLER_44_770 ();
 sg13g2_decap_8 FILLER_44_777 ();
 sg13g2_decap_8 FILLER_44_784 ();
 sg13g2_decap_8 FILLER_44_791 ();
 sg13g2_decap_8 FILLER_44_798 ();
 sg13g2_decap_8 FILLER_44_805 ();
 sg13g2_decap_8 FILLER_44_812 ();
 sg13g2_decap_8 FILLER_44_819 ();
 sg13g2_decap_8 FILLER_44_826 ();
 sg13g2_decap_8 FILLER_44_833 ();
 sg13g2_decap_8 FILLER_44_840 ();
 sg13g2_decap_8 FILLER_44_847 ();
 sg13g2_decap_8 FILLER_44_854 ();
 sg13g2_decap_8 FILLER_44_861 ();
 sg13g2_decap_8 FILLER_44_868 ();
 sg13g2_decap_8 FILLER_44_875 ();
 sg13g2_decap_8 FILLER_44_882 ();
 sg13g2_decap_8 FILLER_44_889 ();
 sg13g2_decap_8 FILLER_44_896 ();
 sg13g2_decap_8 FILLER_44_903 ();
 sg13g2_decap_8 FILLER_44_910 ();
 sg13g2_decap_8 FILLER_44_917 ();
 sg13g2_decap_8 FILLER_44_924 ();
 sg13g2_decap_8 FILLER_44_931 ();
 sg13g2_decap_8 FILLER_44_938 ();
 sg13g2_decap_8 FILLER_44_945 ();
 sg13g2_decap_8 FILLER_44_952 ();
 sg13g2_decap_8 FILLER_44_959 ();
 sg13g2_decap_8 FILLER_44_966 ();
 sg13g2_decap_8 FILLER_44_973 ();
 sg13g2_decap_8 FILLER_44_980 ();
 sg13g2_decap_8 FILLER_44_987 ();
 sg13g2_decap_8 FILLER_44_994 ();
 sg13g2_decap_8 FILLER_44_1001 ();
 sg13g2_decap_8 FILLER_44_1008 ();
 sg13g2_decap_8 FILLER_44_1015 ();
 sg13g2_decap_8 FILLER_44_1022 ();
 sg13g2_decap_8 FILLER_44_1029 ();
 sg13g2_decap_8 FILLER_44_1036 ();
 sg13g2_decap_8 FILLER_44_1043 ();
 sg13g2_decap_8 FILLER_44_1050 ();
 sg13g2_decap_8 FILLER_44_1057 ();
 sg13g2_decap_8 FILLER_44_1064 ();
 sg13g2_decap_8 FILLER_44_1071 ();
 sg13g2_decap_8 FILLER_44_1078 ();
 sg13g2_decap_8 FILLER_44_1085 ();
 sg13g2_decap_8 FILLER_44_1092 ();
 sg13g2_decap_8 FILLER_44_1099 ();
 sg13g2_decap_8 FILLER_44_1106 ();
 sg13g2_decap_8 FILLER_44_1113 ();
 sg13g2_decap_8 FILLER_44_1120 ();
 sg13g2_decap_8 FILLER_44_1127 ();
 sg13g2_decap_8 FILLER_44_1134 ();
 sg13g2_decap_8 FILLER_44_1141 ();
 sg13g2_decap_8 FILLER_44_1148 ();
 sg13g2_decap_8 FILLER_44_1155 ();
 sg13g2_decap_8 FILLER_44_1162 ();
 sg13g2_decap_8 FILLER_44_1169 ();
 sg13g2_decap_8 FILLER_44_1176 ();
 sg13g2_decap_8 FILLER_44_1183 ();
 sg13g2_decap_8 FILLER_44_1190 ();
 sg13g2_decap_8 FILLER_44_1197 ();
 sg13g2_decap_8 FILLER_44_1204 ();
 sg13g2_decap_8 FILLER_44_1211 ();
 sg13g2_decap_8 FILLER_44_1218 ();
 sg13g2_decap_8 FILLER_44_1225 ();
 sg13g2_decap_8 FILLER_44_1232 ();
 sg13g2_decap_8 FILLER_44_1239 ();
 sg13g2_decap_8 FILLER_44_1246 ();
 sg13g2_decap_8 FILLER_44_1253 ();
 sg13g2_decap_8 FILLER_44_1260 ();
 sg13g2_decap_8 FILLER_44_1267 ();
 sg13g2_decap_8 FILLER_44_1274 ();
 sg13g2_decap_8 FILLER_44_1281 ();
 sg13g2_decap_8 FILLER_44_1288 ();
 sg13g2_decap_8 FILLER_44_1295 ();
 sg13g2_decap_8 FILLER_44_1302 ();
 sg13g2_decap_8 FILLER_44_1309 ();
 sg13g2_decap_8 FILLER_44_1316 ();
 sg13g2_decap_8 FILLER_44_1323 ();
 sg13g2_decap_8 FILLER_44_1330 ();
 sg13g2_decap_8 FILLER_44_1337 ();
 sg13g2_decap_8 FILLER_44_1344 ();
 sg13g2_decap_8 FILLER_44_1351 ();
 sg13g2_decap_8 FILLER_44_1358 ();
 sg13g2_decap_8 FILLER_44_1365 ();
 sg13g2_decap_8 FILLER_44_1372 ();
 sg13g2_decap_8 FILLER_44_1379 ();
 sg13g2_decap_8 FILLER_44_1386 ();
 sg13g2_decap_8 FILLER_44_1393 ();
 sg13g2_decap_8 FILLER_44_1400 ();
 sg13g2_decap_8 FILLER_44_1407 ();
 sg13g2_decap_8 FILLER_44_1414 ();
 sg13g2_decap_8 FILLER_44_1421 ();
 sg13g2_decap_8 FILLER_44_1428 ();
 sg13g2_decap_8 FILLER_44_1435 ();
 sg13g2_decap_8 FILLER_44_1442 ();
 sg13g2_decap_8 FILLER_44_1449 ();
 sg13g2_decap_8 FILLER_44_1456 ();
 sg13g2_decap_8 FILLER_44_1463 ();
 sg13g2_decap_8 FILLER_44_1470 ();
 sg13g2_decap_8 FILLER_44_1477 ();
 sg13g2_decap_8 FILLER_44_1484 ();
 sg13g2_decap_8 FILLER_44_1491 ();
 sg13g2_decap_8 FILLER_44_1498 ();
 sg13g2_decap_8 FILLER_44_1505 ();
 sg13g2_decap_8 FILLER_44_1512 ();
 sg13g2_decap_8 FILLER_44_1519 ();
 sg13g2_decap_8 FILLER_44_1526 ();
 sg13g2_decap_8 FILLER_44_1533 ();
 sg13g2_decap_8 FILLER_44_1540 ();
 sg13g2_decap_8 FILLER_44_1547 ();
 sg13g2_decap_8 FILLER_44_1554 ();
 sg13g2_decap_8 FILLER_44_1561 ();
 sg13g2_decap_8 FILLER_44_1568 ();
 sg13g2_decap_8 FILLER_44_1575 ();
 sg13g2_decap_8 FILLER_44_1582 ();
 sg13g2_decap_8 FILLER_44_1589 ();
 sg13g2_decap_8 FILLER_44_1596 ();
 sg13g2_decap_8 FILLER_44_1603 ();
 sg13g2_decap_8 FILLER_44_1610 ();
 sg13g2_decap_8 FILLER_44_1617 ();
 sg13g2_decap_8 FILLER_44_1624 ();
 sg13g2_decap_8 FILLER_44_1631 ();
 sg13g2_decap_8 FILLER_44_1638 ();
 sg13g2_decap_8 FILLER_44_1645 ();
 sg13g2_decap_8 FILLER_44_1652 ();
 sg13g2_decap_8 FILLER_44_1659 ();
 sg13g2_decap_8 FILLER_44_1666 ();
 sg13g2_decap_8 FILLER_44_1673 ();
 sg13g2_decap_8 FILLER_44_1680 ();
 sg13g2_decap_8 FILLER_44_1687 ();
 sg13g2_decap_8 FILLER_44_1694 ();
 sg13g2_decap_8 FILLER_44_1701 ();
 sg13g2_decap_8 FILLER_44_1708 ();
 sg13g2_decap_8 FILLER_44_1715 ();
 sg13g2_decap_8 FILLER_44_1722 ();
 sg13g2_decap_8 FILLER_44_1729 ();
 sg13g2_decap_8 FILLER_44_1736 ();
 sg13g2_decap_8 FILLER_44_1743 ();
 sg13g2_decap_8 FILLER_44_1750 ();
 sg13g2_decap_8 FILLER_44_1757 ();
 sg13g2_decap_8 FILLER_44_1764 ();
 sg13g2_decap_8 FILLER_44_1771 ();
 sg13g2_decap_8 FILLER_44_1778 ();
 sg13g2_decap_8 FILLER_44_1785 ();
 sg13g2_decap_8 FILLER_44_1792 ();
 sg13g2_decap_8 FILLER_44_1799 ();
 sg13g2_decap_8 FILLER_44_1806 ();
 sg13g2_decap_8 FILLER_44_1813 ();
 sg13g2_decap_8 FILLER_44_1820 ();
 sg13g2_decap_8 FILLER_44_1827 ();
 sg13g2_decap_8 FILLER_44_1834 ();
 sg13g2_decap_8 FILLER_44_1841 ();
 sg13g2_decap_8 FILLER_44_1848 ();
 sg13g2_decap_8 FILLER_44_1855 ();
 sg13g2_decap_8 FILLER_44_1862 ();
 sg13g2_decap_8 FILLER_44_1869 ();
 sg13g2_decap_8 FILLER_44_1876 ();
 sg13g2_decap_8 FILLER_44_1883 ();
 sg13g2_decap_8 FILLER_44_1890 ();
 sg13g2_decap_8 FILLER_44_1897 ();
 sg13g2_decap_8 FILLER_44_1904 ();
 sg13g2_decap_8 FILLER_44_1911 ();
 sg13g2_decap_8 FILLER_44_1918 ();
 sg13g2_decap_8 FILLER_44_1925 ();
 sg13g2_decap_8 FILLER_44_1932 ();
 sg13g2_decap_8 FILLER_44_1939 ();
 sg13g2_decap_8 FILLER_44_1946 ();
 sg13g2_decap_8 FILLER_44_1953 ();
 sg13g2_decap_8 FILLER_44_1960 ();
 sg13g2_decap_8 FILLER_44_1967 ();
 sg13g2_decap_8 FILLER_44_1974 ();
 sg13g2_decap_8 FILLER_44_1981 ();
 sg13g2_decap_8 FILLER_44_1988 ();
 sg13g2_decap_8 FILLER_44_1995 ();
 sg13g2_decap_8 FILLER_44_2002 ();
 sg13g2_decap_8 FILLER_44_2009 ();
 sg13g2_decap_8 FILLER_44_2016 ();
 sg13g2_decap_8 FILLER_44_2023 ();
 sg13g2_decap_8 FILLER_44_2030 ();
 sg13g2_decap_8 FILLER_44_2037 ();
 sg13g2_decap_8 FILLER_44_2044 ();
 sg13g2_decap_8 FILLER_44_2051 ();
 sg13g2_decap_8 FILLER_44_2058 ();
 sg13g2_decap_8 FILLER_44_2065 ();
 sg13g2_decap_8 FILLER_44_2072 ();
 sg13g2_decap_8 FILLER_44_2079 ();
 sg13g2_decap_8 FILLER_44_2086 ();
 sg13g2_decap_8 FILLER_44_2093 ();
 sg13g2_decap_8 FILLER_44_2100 ();
 sg13g2_decap_8 FILLER_44_2107 ();
 sg13g2_decap_8 FILLER_44_2114 ();
 sg13g2_decap_8 FILLER_44_2121 ();
 sg13g2_decap_8 FILLER_44_2128 ();
 sg13g2_decap_8 FILLER_44_2135 ();
 sg13g2_decap_8 FILLER_44_2142 ();
 sg13g2_decap_8 FILLER_44_2149 ();
 sg13g2_decap_8 FILLER_44_2156 ();
 sg13g2_decap_8 FILLER_44_2163 ();
 sg13g2_decap_8 FILLER_44_2170 ();
 sg13g2_decap_8 FILLER_44_2177 ();
 sg13g2_decap_8 FILLER_44_2184 ();
 sg13g2_decap_8 FILLER_44_2191 ();
 sg13g2_decap_8 FILLER_44_2198 ();
 sg13g2_decap_8 FILLER_44_2205 ();
 sg13g2_decap_8 FILLER_44_2212 ();
 sg13g2_decap_8 FILLER_44_2219 ();
 sg13g2_decap_8 FILLER_44_2226 ();
 sg13g2_decap_8 FILLER_44_2233 ();
 sg13g2_decap_8 FILLER_44_2240 ();
 sg13g2_decap_8 FILLER_44_2247 ();
 sg13g2_decap_8 FILLER_44_2254 ();
 sg13g2_decap_8 FILLER_44_2261 ();
 sg13g2_decap_8 FILLER_44_2268 ();
 sg13g2_decap_8 FILLER_44_2275 ();
 sg13g2_decap_8 FILLER_44_2282 ();
 sg13g2_decap_8 FILLER_44_2289 ();
 sg13g2_decap_8 FILLER_44_2296 ();
 sg13g2_decap_8 FILLER_44_2303 ();
 sg13g2_decap_8 FILLER_44_2310 ();
 sg13g2_decap_8 FILLER_44_2317 ();
 sg13g2_decap_8 FILLER_44_2324 ();
 sg13g2_decap_8 FILLER_44_2331 ();
 sg13g2_decap_8 FILLER_44_2338 ();
 sg13g2_decap_8 FILLER_44_2345 ();
 sg13g2_decap_8 FILLER_44_2352 ();
 sg13g2_decap_8 FILLER_44_2359 ();
 sg13g2_decap_8 FILLER_44_2366 ();
 sg13g2_decap_8 FILLER_44_2373 ();
 sg13g2_decap_8 FILLER_44_2380 ();
 sg13g2_decap_8 FILLER_44_2387 ();
 sg13g2_decap_8 FILLER_44_2394 ();
 sg13g2_decap_8 FILLER_44_2401 ();
 sg13g2_decap_8 FILLER_44_2408 ();
 sg13g2_decap_8 FILLER_44_2415 ();
 sg13g2_decap_8 FILLER_44_2422 ();
 sg13g2_decap_8 FILLER_44_2429 ();
 sg13g2_decap_8 FILLER_44_2436 ();
 sg13g2_decap_8 FILLER_44_2443 ();
 sg13g2_decap_8 FILLER_44_2450 ();
 sg13g2_decap_8 FILLER_44_2457 ();
 sg13g2_decap_8 FILLER_44_2464 ();
 sg13g2_decap_8 FILLER_44_2471 ();
 sg13g2_decap_8 FILLER_44_2478 ();
 sg13g2_decap_8 FILLER_44_2485 ();
 sg13g2_decap_8 FILLER_44_2492 ();
 sg13g2_decap_8 FILLER_44_2499 ();
 sg13g2_decap_8 FILLER_44_2506 ();
 sg13g2_decap_8 FILLER_44_2513 ();
 sg13g2_decap_8 FILLER_44_2520 ();
 sg13g2_decap_8 FILLER_44_2527 ();
 sg13g2_decap_8 FILLER_44_2534 ();
 sg13g2_decap_8 FILLER_44_2541 ();
 sg13g2_decap_8 FILLER_44_2548 ();
 sg13g2_decap_8 FILLER_44_2555 ();
 sg13g2_decap_8 FILLER_44_2562 ();
 sg13g2_decap_8 FILLER_44_2569 ();
 sg13g2_decap_8 FILLER_44_2576 ();
 sg13g2_decap_8 FILLER_44_2583 ();
 sg13g2_decap_8 FILLER_44_2590 ();
 sg13g2_decap_8 FILLER_44_2597 ();
 sg13g2_decap_8 FILLER_44_2604 ();
 sg13g2_decap_8 FILLER_44_2611 ();
 sg13g2_decap_8 FILLER_44_2618 ();
 sg13g2_decap_8 FILLER_44_2625 ();
 sg13g2_decap_8 FILLER_44_2632 ();
 sg13g2_decap_8 FILLER_44_2639 ();
 sg13g2_decap_8 FILLER_44_2646 ();
 sg13g2_decap_8 FILLER_44_2653 ();
 sg13g2_decap_8 FILLER_44_2660 ();
 sg13g2_decap_8 FILLER_44_2667 ();
 sg13g2_decap_8 FILLER_44_2674 ();
 sg13g2_decap_8 FILLER_44_2681 ();
 sg13g2_decap_8 FILLER_44_2688 ();
 sg13g2_decap_8 FILLER_44_2695 ();
 sg13g2_decap_8 FILLER_44_2702 ();
 sg13g2_decap_8 FILLER_44_2709 ();
 sg13g2_decap_8 FILLER_44_2716 ();
 sg13g2_decap_8 FILLER_44_2723 ();
 sg13g2_decap_8 FILLER_44_2730 ();
 sg13g2_decap_8 FILLER_44_2737 ();
 sg13g2_decap_8 FILLER_44_2744 ();
 sg13g2_decap_8 FILLER_44_2751 ();
 sg13g2_decap_8 FILLER_44_2758 ();
 sg13g2_decap_8 FILLER_44_2765 ();
 sg13g2_decap_8 FILLER_44_2772 ();
 sg13g2_decap_8 FILLER_44_2779 ();
 sg13g2_decap_8 FILLER_44_2786 ();
 sg13g2_decap_8 FILLER_44_2793 ();
 sg13g2_decap_8 FILLER_44_2800 ();
 sg13g2_decap_8 FILLER_44_2807 ();
 sg13g2_decap_8 FILLER_44_2814 ();
 sg13g2_decap_8 FILLER_44_2821 ();
 sg13g2_decap_8 FILLER_44_2828 ();
 sg13g2_decap_8 FILLER_44_2835 ();
 sg13g2_decap_8 FILLER_44_2842 ();
 sg13g2_decap_8 FILLER_44_2849 ();
 sg13g2_decap_8 FILLER_44_2856 ();
 sg13g2_decap_8 FILLER_44_2863 ();
 sg13g2_decap_8 FILLER_44_2870 ();
 sg13g2_decap_8 FILLER_44_2877 ();
 sg13g2_decap_8 FILLER_44_2884 ();
 sg13g2_decap_8 FILLER_44_2891 ();
 sg13g2_decap_8 FILLER_44_2898 ();
 sg13g2_decap_8 FILLER_44_2905 ();
 sg13g2_decap_8 FILLER_44_2912 ();
 sg13g2_decap_8 FILLER_44_2919 ();
 sg13g2_decap_8 FILLER_44_2926 ();
 sg13g2_decap_8 FILLER_44_2933 ();
 sg13g2_decap_8 FILLER_44_2940 ();
 sg13g2_decap_8 FILLER_44_2947 ();
 sg13g2_decap_8 FILLER_44_2954 ();
 sg13g2_decap_8 FILLER_44_2961 ();
 sg13g2_decap_8 FILLER_44_2968 ();
 sg13g2_decap_8 FILLER_44_2975 ();
 sg13g2_decap_8 FILLER_44_2982 ();
 sg13g2_decap_8 FILLER_44_2989 ();
 sg13g2_decap_8 FILLER_44_2996 ();
 sg13g2_decap_8 FILLER_44_3003 ();
 sg13g2_decap_8 FILLER_44_3010 ();
 sg13g2_decap_8 FILLER_44_3017 ();
 sg13g2_decap_8 FILLER_44_3024 ();
 sg13g2_decap_8 FILLER_44_3031 ();
 sg13g2_decap_8 FILLER_44_3038 ();
 sg13g2_decap_8 FILLER_44_3045 ();
 sg13g2_decap_8 FILLER_44_3052 ();
 sg13g2_decap_8 FILLER_44_3059 ();
 sg13g2_decap_8 FILLER_44_3066 ();
 sg13g2_decap_8 FILLER_44_3073 ();
 sg13g2_decap_8 FILLER_44_3080 ();
 sg13g2_decap_8 FILLER_44_3087 ();
 sg13g2_decap_8 FILLER_44_3094 ();
 sg13g2_decap_8 FILLER_44_3101 ();
 sg13g2_decap_8 FILLER_44_3108 ();
 sg13g2_decap_8 FILLER_44_3115 ();
 sg13g2_decap_8 FILLER_44_3122 ();
 sg13g2_decap_8 FILLER_44_3129 ();
 sg13g2_decap_8 FILLER_44_3136 ();
 sg13g2_decap_8 FILLER_44_3143 ();
 sg13g2_decap_8 FILLER_44_3150 ();
 sg13g2_decap_8 FILLER_44_3157 ();
 sg13g2_decap_8 FILLER_44_3164 ();
 sg13g2_decap_8 FILLER_44_3171 ();
 sg13g2_decap_8 FILLER_44_3178 ();
 sg13g2_decap_8 FILLER_44_3185 ();
 sg13g2_decap_8 FILLER_44_3192 ();
 sg13g2_decap_8 FILLER_44_3199 ();
 sg13g2_decap_8 FILLER_44_3206 ();
 sg13g2_decap_8 FILLER_44_3213 ();
 sg13g2_decap_8 FILLER_44_3220 ();
 sg13g2_decap_8 FILLER_44_3227 ();
 sg13g2_decap_8 FILLER_44_3234 ();
 sg13g2_decap_8 FILLER_44_3241 ();
 sg13g2_decap_8 FILLER_44_3248 ();
 sg13g2_decap_8 FILLER_44_3255 ();
 sg13g2_decap_8 FILLER_44_3262 ();
 sg13g2_decap_8 FILLER_44_3269 ();
 sg13g2_decap_8 FILLER_44_3276 ();
 sg13g2_decap_8 FILLER_44_3283 ();
 sg13g2_decap_8 FILLER_44_3290 ();
 sg13g2_decap_8 FILLER_44_3297 ();
 sg13g2_decap_8 FILLER_44_3304 ();
 sg13g2_decap_8 FILLER_44_3311 ();
 sg13g2_decap_8 FILLER_44_3318 ();
 sg13g2_decap_8 FILLER_44_3325 ();
 sg13g2_decap_8 FILLER_44_3332 ();
 sg13g2_decap_8 FILLER_44_3339 ();
 sg13g2_decap_8 FILLER_44_3346 ();
 sg13g2_decap_8 FILLER_44_3353 ();
 sg13g2_decap_8 FILLER_44_3360 ();
 sg13g2_decap_8 FILLER_44_3367 ();
 sg13g2_decap_8 FILLER_44_3374 ();
 sg13g2_decap_8 FILLER_44_3381 ();
 sg13g2_decap_8 FILLER_44_3388 ();
 sg13g2_decap_8 FILLER_44_3395 ();
 sg13g2_decap_8 FILLER_44_3402 ();
 sg13g2_decap_8 FILLER_44_3409 ();
 sg13g2_decap_8 FILLER_44_3416 ();
 sg13g2_decap_8 FILLER_44_3423 ();
 sg13g2_decap_8 FILLER_44_3430 ();
 sg13g2_decap_8 FILLER_44_3437 ();
 sg13g2_decap_8 FILLER_44_3444 ();
 sg13g2_decap_8 FILLER_44_3451 ();
 sg13g2_decap_8 FILLER_44_3458 ();
 sg13g2_decap_8 FILLER_44_3465 ();
 sg13g2_decap_8 FILLER_44_3472 ();
 sg13g2_decap_8 FILLER_44_3479 ();
 sg13g2_decap_8 FILLER_44_3486 ();
 sg13g2_decap_8 FILLER_44_3493 ();
 sg13g2_decap_8 FILLER_44_3500 ();
 sg13g2_decap_8 FILLER_44_3507 ();
 sg13g2_decap_8 FILLER_44_3514 ();
 sg13g2_decap_8 FILLER_44_3521 ();
 sg13g2_decap_8 FILLER_44_3528 ();
 sg13g2_decap_8 FILLER_44_3535 ();
 sg13g2_decap_8 FILLER_44_3542 ();
 sg13g2_decap_8 FILLER_44_3549 ();
 sg13g2_decap_8 FILLER_44_3556 ();
 sg13g2_decap_8 FILLER_44_3563 ();
 sg13g2_decap_8 FILLER_44_3570 ();
 sg13g2_fill_2 FILLER_44_3577 ();
 sg13g2_fill_1 FILLER_44_3579 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_decap_8 FILLER_45_133 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_decap_8 FILLER_45_147 ();
 sg13g2_decap_8 FILLER_45_154 ();
 sg13g2_decap_8 FILLER_45_161 ();
 sg13g2_decap_8 FILLER_45_168 ();
 sg13g2_decap_8 FILLER_45_175 ();
 sg13g2_decap_8 FILLER_45_182 ();
 sg13g2_decap_8 FILLER_45_189 ();
 sg13g2_decap_8 FILLER_45_196 ();
 sg13g2_decap_8 FILLER_45_203 ();
 sg13g2_decap_8 FILLER_45_210 ();
 sg13g2_decap_8 FILLER_45_217 ();
 sg13g2_decap_8 FILLER_45_224 ();
 sg13g2_decap_8 FILLER_45_231 ();
 sg13g2_decap_8 FILLER_45_238 ();
 sg13g2_decap_8 FILLER_45_245 ();
 sg13g2_decap_8 FILLER_45_252 ();
 sg13g2_decap_8 FILLER_45_259 ();
 sg13g2_decap_8 FILLER_45_266 ();
 sg13g2_decap_8 FILLER_45_273 ();
 sg13g2_decap_8 FILLER_45_280 ();
 sg13g2_decap_8 FILLER_45_287 ();
 sg13g2_decap_8 FILLER_45_294 ();
 sg13g2_decap_8 FILLER_45_301 ();
 sg13g2_decap_8 FILLER_45_308 ();
 sg13g2_decap_8 FILLER_45_315 ();
 sg13g2_decap_8 FILLER_45_322 ();
 sg13g2_decap_8 FILLER_45_329 ();
 sg13g2_decap_8 FILLER_45_336 ();
 sg13g2_decap_8 FILLER_45_343 ();
 sg13g2_decap_8 FILLER_45_350 ();
 sg13g2_decap_8 FILLER_45_357 ();
 sg13g2_decap_8 FILLER_45_364 ();
 sg13g2_decap_8 FILLER_45_371 ();
 sg13g2_decap_8 FILLER_45_378 ();
 sg13g2_decap_8 FILLER_45_385 ();
 sg13g2_decap_8 FILLER_45_392 ();
 sg13g2_decap_8 FILLER_45_399 ();
 sg13g2_decap_8 FILLER_45_406 ();
 sg13g2_decap_8 FILLER_45_413 ();
 sg13g2_decap_8 FILLER_45_420 ();
 sg13g2_decap_8 FILLER_45_427 ();
 sg13g2_decap_8 FILLER_45_434 ();
 sg13g2_decap_8 FILLER_45_441 ();
 sg13g2_decap_8 FILLER_45_448 ();
 sg13g2_decap_8 FILLER_45_455 ();
 sg13g2_decap_8 FILLER_45_462 ();
 sg13g2_decap_8 FILLER_45_469 ();
 sg13g2_decap_8 FILLER_45_476 ();
 sg13g2_decap_8 FILLER_45_483 ();
 sg13g2_decap_8 FILLER_45_490 ();
 sg13g2_decap_8 FILLER_45_497 ();
 sg13g2_decap_8 FILLER_45_504 ();
 sg13g2_decap_8 FILLER_45_511 ();
 sg13g2_decap_8 FILLER_45_518 ();
 sg13g2_decap_8 FILLER_45_525 ();
 sg13g2_decap_8 FILLER_45_532 ();
 sg13g2_decap_8 FILLER_45_539 ();
 sg13g2_decap_8 FILLER_45_546 ();
 sg13g2_decap_8 FILLER_45_553 ();
 sg13g2_decap_8 FILLER_45_560 ();
 sg13g2_decap_8 FILLER_45_567 ();
 sg13g2_decap_8 FILLER_45_574 ();
 sg13g2_decap_8 FILLER_45_581 ();
 sg13g2_decap_8 FILLER_45_588 ();
 sg13g2_decap_8 FILLER_45_595 ();
 sg13g2_decap_8 FILLER_45_602 ();
 sg13g2_decap_8 FILLER_45_609 ();
 sg13g2_decap_8 FILLER_45_616 ();
 sg13g2_decap_8 FILLER_45_623 ();
 sg13g2_decap_8 FILLER_45_630 ();
 sg13g2_decap_8 FILLER_45_637 ();
 sg13g2_decap_8 FILLER_45_644 ();
 sg13g2_decap_8 FILLER_45_651 ();
 sg13g2_decap_8 FILLER_45_658 ();
 sg13g2_decap_8 FILLER_45_665 ();
 sg13g2_decap_8 FILLER_45_672 ();
 sg13g2_decap_8 FILLER_45_679 ();
 sg13g2_decap_8 FILLER_45_686 ();
 sg13g2_decap_8 FILLER_45_693 ();
 sg13g2_decap_8 FILLER_45_700 ();
 sg13g2_decap_8 FILLER_45_707 ();
 sg13g2_decap_8 FILLER_45_714 ();
 sg13g2_decap_8 FILLER_45_721 ();
 sg13g2_decap_8 FILLER_45_728 ();
 sg13g2_decap_8 FILLER_45_735 ();
 sg13g2_decap_8 FILLER_45_742 ();
 sg13g2_decap_8 FILLER_45_749 ();
 sg13g2_decap_8 FILLER_45_756 ();
 sg13g2_decap_8 FILLER_45_763 ();
 sg13g2_decap_8 FILLER_45_770 ();
 sg13g2_decap_8 FILLER_45_777 ();
 sg13g2_decap_8 FILLER_45_784 ();
 sg13g2_decap_8 FILLER_45_791 ();
 sg13g2_decap_8 FILLER_45_798 ();
 sg13g2_decap_8 FILLER_45_805 ();
 sg13g2_decap_8 FILLER_45_812 ();
 sg13g2_decap_8 FILLER_45_819 ();
 sg13g2_decap_8 FILLER_45_826 ();
 sg13g2_decap_8 FILLER_45_833 ();
 sg13g2_decap_8 FILLER_45_840 ();
 sg13g2_decap_8 FILLER_45_847 ();
 sg13g2_decap_8 FILLER_45_854 ();
 sg13g2_decap_8 FILLER_45_861 ();
 sg13g2_decap_8 FILLER_45_868 ();
 sg13g2_decap_8 FILLER_45_875 ();
 sg13g2_decap_8 FILLER_45_882 ();
 sg13g2_decap_8 FILLER_45_889 ();
 sg13g2_decap_8 FILLER_45_896 ();
 sg13g2_decap_8 FILLER_45_903 ();
 sg13g2_decap_8 FILLER_45_910 ();
 sg13g2_decap_8 FILLER_45_917 ();
 sg13g2_decap_8 FILLER_45_924 ();
 sg13g2_decap_8 FILLER_45_931 ();
 sg13g2_decap_8 FILLER_45_938 ();
 sg13g2_decap_8 FILLER_45_945 ();
 sg13g2_decap_8 FILLER_45_952 ();
 sg13g2_decap_8 FILLER_45_959 ();
 sg13g2_decap_8 FILLER_45_966 ();
 sg13g2_decap_8 FILLER_45_973 ();
 sg13g2_decap_8 FILLER_45_980 ();
 sg13g2_decap_8 FILLER_45_987 ();
 sg13g2_decap_8 FILLER_45_994 ();
 sg13g2_decap_8 FILLER_45_1001 ();
 sg13g2_decap_8 FILLER_45_1008 ();
 sg13g2_decap_8 FILLER_45_1015 ();
 sg13g2_decap_8 FILLER_45_1022 ();
 sg13g2_decap_8 FILLER_45_1029 ();
 sg13g2_decap_8 FILLER_45_1036 ();
 sg13g2_decap_8 FILLER_45_1043 ();
 sg13g2_decap_8 FILLER_45_1050 ();
 sg13g2_decap_8 FILLER_45_1057 ();
 sg13g2_decap_8 FILLER_45_1064 ();
 sg13g2_decap_8 FILLER_45_1071 ();
 sg13g2_decap_8 FILLER_45_1078 ();
 sg13g2_decap_8 FILLER_45_1085 ();
 sg13g2_decap_8 FILLER_45_1092 ();
 sg13g2_decap_8 FILLER_45_1099 ();
 sg13g2_decap_8 FILLER_45_1106 ();
 sg13g2_decap_8 FILLER_45_1113 ();
 sg13g2_decap_8 FILLER_45_1120 ();
 sg13g2_decap_8 FILLER_45_1127 ();
 sg13g2_decap_8 FILLER_45_1134 ();
 sg13g2_decap_8 FILLER_45_1141 ();
 sg13g2_decap_8 FILLER_45_1148 ();
 sg13g2_decap_8 FILLER_45_1155 ();
 sg13g2_decap_8 FILLER_45_1162 ();
 sg13g2_decap_8 FILLER_45_1169 ();
 sg13g2_decap_8 FILLER_45_1176 ();
 sg13g2_decap_8 FILLER_45_1183 ();
 sg13g2_decap_8 FILLER_45_1190 ();
 sg13g2_decap_8 FILLER_45_1197 ();
 sg13g2_decap_8 FILLER_45_1204 ();
 sg13g2_decap_8 FILLER_45_1211 ();
 sg13g2_decap_8 FILLER_45_1218 ();
 sg13g2_decap_8 FILLER_45_1225 ();
 sg13g2_decap_8 FILLER_45_1232 ();
 sg13g2_decap_8 FILLER_45_1239 ();
 sg13g2_decap_8 FILLER_45_1246 ();
 sg13g2_decap_8 FILLER_45_1253 ();
 sg13g2_decap_8 FILLER_45_1260 ();
 sg13g2_decap_8 FILLER_45_1267 ();
 sg13g2_decap_8 FILLER_45_1274 ();
 sg13g2_decap_8 FILLER_45_1281 ();
 sg13g2_decap_8 FILLER_45_1288 ();
 sg13g2_decap_8 FILLER_45_1295 ();
 sg13g2_decap_8 FILLER_45_1302 ();
 sg13g2_decap_8 FILLER_45_1309 ();
 sg13g2_decap_8 FILLER_45_1316 ();
 sg13g2_decap_8 FILLER_45_1323 ();
 sg13g2_decap_8 FILLER_45_1330 ();
 sg13g2_decap_8 FILLER_45_1337 ();
 sg13g2_decap_8 FILLER_45_1344 ();
 sg13g2_decap_8 FILLER_45_1351 ();
 sg13g2_decap_8 FILLER_45_1358 ();
 sg13g2_decap_8 FILLER_45_1365 ();
 sg13g2_decap_8 FILLER_45_1372 ();
 sg13g2_decap_8 FILLER_45_1379 ();
 sg13g2_decap_8 FILLER_45_1386 ();
 sg13g2_decap_8 FILLER_45_1393 ();
 sg13g2_decap_8 FILLER_45_1400 ();
 sg13g2_decap_8 FILLER_45_1407 ();
 sg13g2_decap_8 FILLER_45_1414 ();
 sg13g2_decap_8 FILLER_45_1421 ();
 sg13g2_decap_8 FILLER_45_1428 ();
 sg13g2_decap_8 FILLER_45_1435 ();
 sg13g2_decap_8 FILLER_45_1442 ();
 sg13g2_decap_8 FILLER_45_1449 ();
 sg13g2_decap_8 FILLER_45_1456 ();
 sg13g2_decap_8 FILLER_45_1463 ();
 sg13g2_decap_8 FILLER_45_1470 ();
 sg13g2_decap_8 FILLER_45_1477 ();
 sg13g2_decap_8 FILLER_45_1484 ();
 sg13g2_decap_8 FILLER_45_1491 ();
 sg13g2_decap_8 FILLER_45_1498 ();
 sg13g2_decap_8 FILLER_45_1505 ();
 sg13g2_decap_8 FILLER_45_1512 ();
 sg13g2_decap_8 FILLER_45_1519 ();
 sg13g2_decap_8 FILLER_45_1526 ();
 sg13g2_decap_8 FILLER_45_1533 ();
 sg13g2_decap_8 FILLER_45_1540 ();
 sg13g2_decap_8 FILLER_45_1547 ();
 sg13g2_decap_8 FILLER_45_1554 ();
 sg13g2_decap_8 FILLER_45_1561 ();
 sg13g2_decap_8 FILLER_45_1568 ();
 sg13g2_decap_8 FILLER_45_1575 ();
 sg13g2_decap_8 FILLER_45_1582 ();
 sg13g2_decap_8 FILLER_45_1589 ();
 sg13g2_decap_8 FILLER_45_1596 ();
 sg13g2_decap_8 FILLER_45_1603 ();
 sg13g2_decap_8 FILLER_45_1610 ();
 sg13g2_decap_8 FILLER_45_1617 ();
 sg13g2_decap_8 FILLER_45_1624 ();
 sg13g2_decap_8 FILLER_45_1631 ();
 sg13g2_decap_8 FILLER_45_1638 ();
 sg13g2_decap_8 FILLER_45_1645 ();
 sg13g2_decap_8 FILLER_45_1652 ();
 sg13g2_decap_8 FILLER_45_1659 ();
 sg13g2_decap_8 FILLER_45_1666 ();
 sg13g2_decap_8 FILLER_45_1673 ();
 sg13g2_decap_8 FILLER_45_1680 ();
 sg13g2_decap_8 FILLER_45_1687 ();
 sg13g2_decap_8 FILLER_45_1694 ();
 sg13g2_decap_8 FILLER_45_1701 ();
 sg13g2_decap_8 FILLER_45_1708 ();
 sg13g2_decap_8 FILLER_45_1715 ();
 sg13g2_decap_8 FILLER_45_1722 ();
 sg13g2_decap_8 FILLER_45_1729 ();
 sg13g2_decap_8 FILLER_45_1736 ();
 sg13g2_decap_8 FILLER_45_1743 ();
 sg13g2_decap_8 FILLER_45_1750 ();
 sg13g2_decap_8 FILLER_45_1757 ();
 sg13g2_decap_8 FILLER_45_1764 ();
 sg13g2_decap_8 FILLER_45_1771 ();
 sg13g2_decap_8 FILLER_45_1778 ();
 sg13g2_decap_8 FILLER_45_1785 ();
 sg13g2_decap_8 FILLER_45_1792 ();
 sg13g2_decap_8 FILLER_45_1799 ();
 sg13g2_decap_8 FILLER_45_1806 ();
 sg13g2_decap_8 FILLER_45_1813 ();
 sg13g2_decap_8 FILLER_45_1820 ();
 sg13g2_decap_8 FILLER_45_1827 ();
 sg13g2_decap_8 FILLER_45_1834 ();
 sg13g2_decap_8 FILLER_45_1841 ();
 sg13g2_decap_8 FILLER_45_1848 ();
 sg13g2_decap_8 FILLER_45_1855 ();
 sg13g2_decap_8 FILLER_45_1862 ();
 sg13g2_decap_8 FILLER_45_1869 ();
 sg13g2_decap_8 FILLER_45_1876 ();
 sg13g2_decap_8 FILLER_45_1883 ();
 sg13g2_decap_8 FILLER_45_1890 ();
 sg13g2_decap_8 FILLER_45_1897 ();
 sg13g2_decap_8 FILLER_45_1904 ();
 sg13g2_decap_8 FILLER_45_1911 ();
 sg13g2_decap_8 FILLER_45_1918 ();
 sg13g2_decap_8 FILLER_45_1925 ();
 sg13g2_decap_8 FILLER_45_1932 ();
 sg13g2_decap_8 FILLER_45_1939 ();
 sg13g2_decap_8 FILLER_45_1946 ();
 sg13g2_decap_8 FILLER_45_1953 ();
 sg13g2_decap_8 FILLER_45_1960 ();
 sg13g2_decap_8 FILLER_45_1967 ();
 sg13g2_decap_8 FILLER_45_1974 ();
 sg13g2_decap_8 FILLER_45_1981 ();
 sg13g2_decap_8 FILLER_45_1988 ();
 sg13g2_decap_8 FILLER_45_1995 ();
 sg13g2_decap_8 FILLER_45_2002 ();
 sg13g2_decap_8 FILLER_45_2009 ();
 sg13g2_decap_8 FILLER_45_2016 ();
 sg13g2_decap_8 FILLER_45_2023 ();
 sg13g2_decap_8 FILLER_45_2030 ();
 sg13g2_decap_8 FILLER_45_2037 ();
 sg13g2_decap_8 FILLER_45_2044 ();
 sg13g2_decap_8 FILLER_45_2051 ();
 sg13g2_decap_8 FILLER_45_2058 ();
 sg13g2_decap_8 FILLER_45_2065 ();
 sg13g2_decap_8 FILLER_45_2072 ();
 sg13g2_decap_8 FILLER_45_2079 ();
 sg13g2_decap_8 FILLER_45_2086 ();
 sg13g2_decap_8 FILLER_45_2093 ();
 sg13g2_decap_8 FILLER_45_2100 ();
 sg13g2_decap_8 FILLER_45_2107 ();
 sg13g2_decap_8 FILLER_45_2114 ();
 sg13g2_decap_8 FILLER_45_2121 ();
 sg13g2_decap_8 FILLER_45_2128 ();
 sg13g2_decap_8 FILLER_45_2135 ();
 sg13g2_decap_8 FILLER_45_2142 ();
 sg13g2_decap_8 FILLER_45_2149 ();
 sg13g2_decap_8 FILLER_45_2156 ();
 sg13g2_decap_8 FILLER_45_2163 ();
 sg13g2_decap_8 FILLER_45_2170 ();
 sg13g2_decap_8 FILLER_45_2177 ();
 sg13g2_decap_8 FILLER_45_2184 ();
 sg13g2_decap_8 FILLER_45_2191 ();
 sg13g2_decap_8 FILLER_45_2198 ();
 sg13g2_decap_8 FILLER_45_2205 ();
 sg13g2_decap_8 FILLER_45_2212 ();
 sg13g2_decap_8 FILLER_45_2219 ();
 sg13g2_decap_8 FILLER_45_2226 ();
 sg13g2_decap_8 FILLER_45_2233 ();
 sg13g2_decap_8 FILLER_45_2240 ();
 sg13g2_decap_8 FILLER_45_2247 ();
 sg13g2_decap_8 FILLER_45_2254 ();
 sg13g2_decap_8 FILLER_45_2261 ();
 sg13g2_decap_8 FILLER_45_2268 ();
 sg13g2_decap_8 FILLER_45_2275 ();
 sg13g2_decap_8 FILLER_45_2282 ();
 sg13g2_decap_8 FILLER_45_2289 ();
 sg13g2_decap_8 FILLER_45_2296 ();
 sg13g2_decap_8 FILLER_45_2303 ();
 sg13g2_decap_8 FILLER_45_2310 ();
 sg13g2_decap_8 FILLER_45_2317 ();
 sg13g2_decap_8 FILLER_45_2324 ();
 sg13g2_decap_8 FILLER_45_2331 ();
 sg13g2_decap_8 FILLER_45_2338 ();
 sg13g2_decap_8 FILLER_45_2345 ();
 sg13g2_decap_8 FILLER_45_2352 ();
 sg13g2_decap_8 FILLER_45_2359 ();
 sg13g2_decap_8 FILLER_45_2366 ();
 sg13g2_decap_8 FILLER_45_2373 ();
 sg13g2_decap_8 FILLER_45_2380 ();
 sg13g2_decap_8 FILLER_45_2387 ();
 sg13g2_decap_8 FILLER_45_2394 ();
 sg13g2_decap_8 FILLER_45_2401 ();
 sg13g2_decap_8 FILLER_45_2408 ();
 sg13g2_decap_8 FILLER_45_2415 ();
 sg13g2_decap_8 FILLER_45_2422 ();
 sg13g2_decap_8 FILLER_45_2429 ();
 sg13g2_decap_8 FILLER_45_2436 ();
 sg13g2_decap_8 FILLER_45_2443 ();
 sg13g2_decap_8 FILLER_45_2450 ();
 sg13g2_decap_8 FILLER_45_2457 ();
 sg13g2_decap_8 FILLER_45_2464 ();
 sg13g2_decap_8 FILLER_45_2471 ();
 sg13g2_decap_8 FILLER_45_2478 ();
 sg13g2_decap_8 FILLER_45_2485 ();
 sg13g2_decap_8 FILLER_45_2492 ();
 sg13g2_decap_8 FILLER_45_2499 ();
 sg13g2_decap_8 FILLER_45_2506 ();
 sg13g2_decap_8 FILLER_45_2513 ();
 sg13g2_decap_8 FILLER_45_2520 ();
 sg13g2_decap_8 FILLER_45_2527 ();
 sg13g2_decap_8 FILLER_45_2534 ();
 sg13g2_decap_8 FILLER_45_2541 ();
 sg13g2_decap_8 FILLER_45_2548 ();
 sg13g2_decap_8 FILLER_45_2555 ();
 sg13g2_decap_8 FILLER_45_2562 ();
 sg13g2_decap_8 FILLER_45_2569 ();
 sg13g2_decap_8 FILLER_45_2576 ();
 sg13g2_decap_8 FILLER_45_2583 ();
 sg13g2_decap_8 FILLER_45_2590 ();
 sg13g2_decap_8 FILLER_45_2597 ();
 sg13g2_decap_8 FILLER_45_2604 ();
 sg13g2_decap_8 FILLER_45_2611 ();
 sg13g2_decap_8 FILLER_45_2618 ();
 sg13g2_decap_8 FILLER_45_2625 ();
 sg13g2_decap_8 FILLER_45_2632 ();
 sg13g2_decap_8 FILLER_45_2639 ();
 sg13g2_decap_8 FILLER_45_2646 ();
 sg13g2_decap_8 FILLER_45_2653 ();
 sg13g2_decap_8 FILLER_45_2660 ();
 sg13g2_decap_8 FILLER_45_2667 ();
 sg13g2_decap_8 FILLER_45_2674 ();
 sg13g2_decap_8 FILLER_45_2681 ();
 sg13g2_decap_8 FILLER_45_2688 ();
 sg13g2_decap_8 FILLER_45_2695 ();
 sg13g2_decap_8 FILLER_45_2702 ();
 sg13g2_decap_8 FILLER_45_2709 ();
 sg13g2_decap_8 FILLER_45_2716 ();
 sg13g2_decap_8 FILLER_45_2723 ();
 sg13g2_decap_8 FILLER_45_2730 ();
 sg13g2_decap_8 FILLER_45_2737 ();
 sg13g2_decap_8 FILLER_45_2744 ();
 sg13g2_decap_8 FILLER_45_2751 ();
 sg13g2_decap_8 FILLER_45_2758 ();
 sg13g2_decap_8 FILLER_45_2765 ();
 sg13g2_decap_8 FILLER_45_2772 ();
 sg13g2_decap_8 FILLER_45_2779 ();
 sg13g2_decap_8 FILLER_45_2786 ();
 sg13g2_decap_8 FILLER_45_2793 ();
 sg13g2_decap_8 FILLER_45_2800 ();
 sg13g2_decap_8 FILLER_45_2807 ();
 sg13g2_decap_8 FILLER_45_2814 ();
 sg13g2_decap_8 FILLER_45_2821 ();
 sg13g2_decap_8 FILLER_45_2828 ();
 sg13g2_decap_8 FILLER_45_2835 ();
 sg13g2_decap_8 FILLER_45_2842 ();
 sg13g2_decap_8 FILLER_45_2849 ();
 sg13g2_decap_8 FILLER_45_2856 ();
 sg13g2_decap_8 FILLER_45_2863 ();
 sg13g2_decap_8 FILLER_45_2870 ();
 sg13g2_decap_8 FILLER_45_2877 ();
 sg13g2_decap_8 FILLER_45_2884 ();
 sg13g2_decap_8 FILLER_45_2891 ();
 sg13g2_decap_8 FILLER_45_2898 ();
 sg13g2_decap_8 FILLER_45_2905 ();
 sg13g2_decap_8 FILLER_45_2912 ();
 sg13g2_decap_8 FILLER_45_2919 ();
 sg13g2_decap_8 FILLER_45_2926 ();
 sg13g2_decap_8 FILLER_45_2933 ();
 sg13g2_decap_8 FILLER_45_2940 ();
 sg13g2_decap_8 FILLER_45_2947 ();
 sg13g2_decap_8 FILLER_45_2954 ();
 sg13g2_decap_8 FILLER_45_2961 ();
 sg13g2_decap_8 FILLER_45_2968 ();
 sg13g2_decap_8 FILLER_45_2975 ();
 sg13g2_decap_8 FILLER_45_2982 ();
 sg13g2_decap_8 FILLER_45_2989 ();
 sg13g2_decap_8 FILLER_45_2996 ();
 sg13g2_decap_8 FILLER_45_3003 ();
 sg13g2_decap_8 FILLER_45_3010 ();
 sg13g2_decap_8 FILLER_45_3017 ();
 sg13g2_decap_8 FILLER_45_3024 ();
 sg13g2_decap_8 FILLER_45_3031 ();
 sg13g2_decap_8 FILLER_45_3038 ();
 sg13g2_decap_8 FILLER_45_3045 ();
 sg13g2_decap_8 FILLER_45_3052 ();
 sg13g2_decap_8 FILLER_45_3059 ();
 sg13g2_decap_8 FILLER_45_3066 ();
 sg13g2_decap_8 FILLER_45_3073 ();
 sg13g2_decap_8 FILLER_45_3080 ();
 sg13g2_decap_8 FILLER_45_3087 ();
 sg13g2_decap_8 FILLER_45_3094 ();
 sg13g2_decap_8 FILLER_45_3101 ();
 sg13g2_decap_8 FILLER_45_3108 ();
 sg13g2_decap_8 FILLER_45_3115 ();
 sg13g2_decap_8 FILLER_45_3122 ();
 sg13g2_decap_8 FILLER_45_3129 ();
 sg13g2_decap_8 FILLER_45_3136 ();
 sg13g2_decap_8 FILLER_45_3143 ();
 sg13g2_decap_8 FILLER_45_3150 ();
 sg13g2_decap_8 FILLER_45_3157 ();
 sg13g2_decap_8 FILLER_45_3164 ();
 sg13g2_decap_8 FILLER_45_3171 ();
 sg13g2_decap_8 FILLER_45_3178 ();
 sg13g2_decap_8 FILLER_45_3185 ();
 sg13g2_decap_8 FILLER_45_3192 ();
 sg13g2_decap_8 FILLER_45_3199 ();
 sg13g2_decap_8 FILLER_45_3206 ();
 sg13g2_decap_8 FILLER_45_3213 ();
 sg13g2_decap_8 FILLER_45_3220 ();
 sg13g2_decap_8 FILLER_45_3227 ();
 sg13g2_decap_8 FILLER_45_3234 ();
 sg13g2_decap_8 FILLER_45_3241 ();
 sg13g2_decap_8 FILLER_45_3248 ();
 sg13g2_decap_8 FILLER_45_3255 ();
 sg13g2_decap_8 FILLER_45_3262 ();
 sg13g2_decap_8 FILLER_45_3269 ();
 sg13g2_decap_8 FILLER_45_3276 ();
 sg13g2_decap_8 FILLER_45_3283 ();
 sg13g2_decap_8 FILLER_45_3290 ();
 sg13g2_decap_8 FILLER_45_3297 ();
 sg13g2_decap_8 FILLER_45_3304 ();
 sg13g2_decap_8 FILLER_45_3311 ();
 sg13g2_decap_8 FILLER_45_3318 ();
 sg13g2_decap_8 FILLER_45_3325 ();
 sg13g2_decap_8 FILLER_45_3332 ();
 sg13g2_decap_8 FILLER_45_3339 ();
 sg13g2_decap_8 FILLER_45_3346 ();
 sg13g2_decap_8 FILLER_45_3353 ();
 sg13g2_decap_8 FILLER_45_3360 ();
 sg13g2_decap_8 FILLER_45_3367 ();
 sg13g2_decap_8 FILLER_45_3374 ();
 sg13g2_decap_8 FILLER_45_3381 ();
 sg13g2_decap_8 FILLER_45_3388 ();
 sg13g2_decap_8 FILLER_45_3395 ();
 sg13g2_decap_8 FILLER_45_3402 ();
 sg13g2_decap_8 FILLER_45_3409 ();
 sg13g2_decap_8 FILLER_45_3416 ();
 sg13g2_decap_8 FILLER_45_3423 ();
 sg13g2_decap_8 FILLER_45_3430 ();
 sg13g2_decap_8 FILLER_45_3437 ();
 sg13g2_decap_8 FILLER_45_3444 ();
 sg13g2_decap_8 FILLER_45_3451 ();
 sg13g2_decap_8 FILLER_45_3458 ();
 sg13g2_decap_8 FILLER_45_3465 ();
 sg13g2_decap_8 FILLER_45_3472 ();
 sg13g2_decap_8 FILLER_45_3479 ();
 sg13g2_decap_8 FILLER_45_3486 ();
 sg13g2_decap_8 FILLER_45_3493 ();
 sg13g2_decap_8 FILLER_45_3500 ();
 sg13g2_decap_8 FILLER_45_3507 ();
 sg13g2_decap_8 FILLER_45_3514 ();
 sg13g2_decap_8 FILLER_45_3521 ();
 sg13g2_decap_8 FILLER_45_3528 ();
 sg13g2_decap_8 FILLER_45_3535 ();
 sg13g2_decap_8 FILLER_45_3542 ();
 sg13g2_decap_8 FILLER_45_3549 ();
 sg13g2_decap_8 FILLER_45_3556 ();
 sg13g2_decap_8 FILLER_45_3563 ();
 sg13g2_decap_8 FILLER_45_3570 ();
 sg13g2_fill_2 FILLER_45_3577 ();
 sg13g2_fill_1 FILLER_45_3579 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_8 FILLER_46_133 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_decap_8 FILLER_46_147 ();
 sg13g2_decap_8 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_161 ();
 sg13g2_decap_8 FILLER_46_168 ();
 sg13g2_decap_8 FILLER_46_175 ();
 sg13g2_decap_8 FILLER_46_182 ();
 sg13g2_decap_8 FILLER_46_189 ();
 sg13g2_decap_8 FILLER_46_196 ();
 sg13g2_decap_8 FILLER_46_203 ();
 sg13g2_decap_8 FILLER_46_210 ();
 sg13g2_decap_8 FILLER_46_217 ();
 sg13g2_decap_8 FILLER_46_224 ();
 sg13g2_decap_8 FILLER_46_231 ();
 sg13g2_decap_8 FILLER_46_238 ();
 sg13g2_decap_8 FILLER_46_245 ();
 sg13g2_decap_8 FILLER_46_252 ();
 sg13g2_decap_8 FILLER_46_259 ();
 sg13g2_decap_8 FILLER_46_266 ();
 sg13g2_decap_8 FILLER_46_273 ();
 sg13g2_decap_8 FILLER_46_280 ();
 sg13g2_decap_8 FILLER_46_287 ();
 sg13g2_decap_8 FILLER_46_294 ();
 sg13g2_decap_8 FILLER_46_301 ();
 sg13g2_decap_8 FILLER_46_308 ();
 sg13g2_decap_8 FILLER_46_315 ();
 sg13g2_decap_8 FILLER_46_322 ();
 sg13g2_decap_8 FILLER_46_329 ();
 sg13g2_decap_8 FILLER_46_336 ();
 sg13g2_decap_8 FILLER_46_343 ();
 sg13g2_decap_8 FILLER_46_350 ();
 sg13g2_decap_8 FILLER_46_357 ();
 sg13g2_decap_8 FILLER_46_364 ();
 sg13g2_decap_8 FILLER_46_371 ();
 sg13g2_decap_8 FILLER_46_378 ();
 sg13g2_decap_8 FILLER_46_385 ();
 sg13g2_decap_8 FILLER_46_392 ();
 sg13g2_decap_8 FILLER_46_399 ();
 sg13g2_decap_8 FILLER_46_406 ();
 sg13g2_decap_8 FILLER_46_413 ();
 sg13g2_decap_8 FILLER_46_420 ();
 sg13g2_decap_8 FILLER_46_427 ();
 sg13g2_decap_8 FILLER_46_434 ();
 sg13g2_decap_8 FILLER_46_441 ();
 sg13g2_decap_8 FILLER_46_448 ();
 sg13g2_decap_8 FILLER_46_455 ();
 sg13g2_decap_8 FILLER_46_462 ();
 sg13g2_decap_8 FILLER_46_469 ();
 sg13g2_decap_8 FILLER_46_476 ();
 sg13g2_decap_8 FILLER_46_483 ();
 sg13g2_decap_8 FILLER_46_490 ();
 sg13g2_decap_8 FILLER_46_497 ();
 sg13g2_decap_8 FILLER_46_504 ();
 sg13g2_decap_8 FILLER_46_511 ();
 sg13g2_decap_8 FILLER_46_518 ();
 sg13g2_decap_8 FILLER_46_525 ();
 sg13g2_decap_8 FILLER_46_532 ();
 sg13g2_decap_8 FILLER_46_539 ();
 sg13g2_decap_8 FILLER_46_546 ();
 sg13g2_decap_8 FILLER_46_553 ();
 sg13g2_decap_8 FILLER_46_560 ();
 sg13g2_decap_8 FILLER_46_567 ();
 sg13g2_decap_8 FILLER_46_574 ();
 sg13g2_decap_8 FILLER_46_581 ();
 sg13g2_decap_8 FILLER_46_588 ();
 sg13g2_decap_8 FILLER_46_595 ();
 sg13g2_decap_8 FILLER_46_602 ();
 sg13g2_decap_8 FILLER_46_609 ();
 sg13g2_decap_8 FILLER_46_616 ();
 sg13g2_decap_8 FILLER_46_623 ();
 sg13g2_decap_8 FILLER_46_630 ();
 sg13g2_decap_8 FILLER_46_637 ();
 sg13g2_decap_8 FILLER_46_644 ();
 sg13g2_decap_8 FILLER_46_651 ();
 sg13g2_decap_8 FILLER_46_658 ();
 sg13g2_decap_8 FILLER_46_665 ();
 sg13g2_decap_8 FILLER_46_672 ();
 sg13g2_decap_8 FILLER_46_679 ();
 sg13g2_decap_8 FILLER_46_686 ();
 sg13g2_decap_8 FILLER_46_693 ();
 sg13g2_decap_8 FILLER_46_700 ();
 sg13g2_decap_8 FILLER_46_707 ();
 sg13g2_decap_8 FILLER_46_714 ();
 sg13g2_decap_8 FILLER_46_721 ();
 sg13g2_decap_8 FILLER_46_728 ();
 sg13g2_decap_8 FILLER_46_735 ();
 sg13g2_decap_8 FILLER_46_742 ();
 sg13g2_decap_8 FILLER_46_749 ();
 sg13g2_decap_8 FILLER_46_756 ();
 sg13g2_decap_8 FILLER_46_763 ();
 sg13g2_decap_8 FILLER_46_770 ();
 sg13g2_decap_8 FILLER_46_777 ();
 sg13g2_decap_8 FILLER_46_784 ();
 sg13g2_decap_8 FILLER_46_791 ();
 sg13g2_decap_8 FILLER_46_798 ();
 sg13g2_decap_8 FILLER_46_805 ();
 sg13g2_decap_8 FILLER_46_812 ();
 sg13g2_decap_8 FILLER_46_819 ();
 sg13g2_decap_8 FILLER_46_826 ();
 sg13g2_decap_8 FILLER_46_833 ();
 sg13g2_decap_8 FILLER_46_840 ();
 sg13g2_decap_8 FILLER_46_847 ();
 sg13g2_decap_8 FILLER_46_854 ();
 sg13g2_decap_8 FILLER_46_861 ();
 sg13g2_decap_8 FILLER_46_868 ();
 sg13g2_decap_8 FILLER_46_875 ();
 sg13g2_decap_8 FILLER_46_882 ();
 sg13g2_decap_8 FILLER_46_889 ();
 sg13g2_decap_8 FILLER_46_896 ();
 sg13g2_decap_8 FILLER_46_903 ();
 sg13g2_decap_8 FILLER_46_910 ();
 sg13g2_decap_8 FILLER_46_917 ();
 sg13g2_decap_8 FILLER_46_924 ();
 sg13g2_decap_8 FILLER_46_931 ();
 sg13g2_decap_8 FILLER_46_938 ();
 sg13g2_decap_8 FILLER_46_945 ();
 sg13g2_decap_8 FILLER_46_952 ();
 sg13g2_decap_8 FILLER_46_959 ();
 sg13g2_decap_8 FILLER_46_966 ();
 sg13g2_decap_8 FILLER_46_973 ();
 sg13g2_decap_8 FILLER_46_980 ();
 sg13g2_decap_8 FILLER_46_987 ();
 sg13g2_decap_8 FILLER_46_994 ();
 sg13g2_decap_8 FILLER_46_1001 ();
 sg13g2_decap_8 FILLER_46_1008 ();
 sg13g2_decap_8 FILLER_46_1015 ();
 sg13g2_decap_8 FILLER_46_1022 ();
 sg13g2_decap_8 FILLER_46_1029 ();
 sg13g2_decap_8 FILLER_46_1036 ();
 sg13g2_decap_8 FILLER_46_1043 ();
 sg13g2_decap_8 FILLER_46_1050 ();
 sg13g2_decap_8 FILLER_46_1057 ();
 sg13g2_decap_8 FILLER_46_1064 ();
 sg13g2_decap_8 FILLER_46_1071 ();
 sg13g2_decap_8 FILLER_46_1078 ();
 sg13g2_decap_8 FILLER_46_1085 ();
 sg13g2_decap_8 FILLER_46_1092 ();
 sg13g2_decap_8 FILLER_46_1099 ();
 sg13g2_decap_8 FILLER_46_1106 ();
 sg13g2_decap_8 FILLER_46_1113 ();
 sg13g2_decap_8 FILLER_46_1120 ();
 sg13g2_decap_8 FILLER_46_1127 ();
 sg13g2_decap_8 FILLER_46_1134 ();
 sg13g2_decap_8 FILLER_46_1141 ();
 sg13g2_decap_8 FILLER_46_1148 ();
 sg13g2_decap_8 FILLER_46_1155 ();
 sg13g2_decap_8 FILLER_46_1162 ();
 sg13g2_decap_8 FILLER_46_1169 ();
 sg13g2_decap_8 FILLER_46_1176 ();
 sg13g2_decap_8 FILLER_46_1183 ();
 sg13g2_decap_8 FILLER_46_1190 ();
 sg13g2_decap_8 FILLER_46_1197 ();
 sg13g2_decap_8 FILLER_46_1204 ();
 sg13g2_decap_8 FILLER_46_1211 ();
 sg13g2_decap_8 FILLER_46_1218 ();
 sg13g2_decap_8 FILLER_46_1225 ();
 sg13g2_decap_8 FILLER_46_1232 ();
 sg13g2_decap_8 FILLER_46_1239 ();
 sg13g2_decap_8 FILLER_46_1246 ();
 sg13g2_decap_8 FILLER_46_1253 ();
 sg13g2_decap_8 FILLER_46_1260 ();
 sg13g2_decap_8 FILLER_46_1267 ();
 sg13g2_decap_8 FILLER_46_1274 ();
 sg13g2_decap_8 FILLER_46_1281 ();
 sg13g2_decap_8 FILLER_46_1288 ();
 sg13g2_decap_8 FILLER_46_1295 ();
 sg13g2_decap_8 FILLER_46_1302 ();
 sg13g2_decap_8 FILLER_46_1309 ();
 sg13g2_decap_8 FILLER_46_1316 ();
 sg13g2_decap_8 FILLER_46_1323 ();
 sg13g2_decap_8 FILLER_46_1330 ();
 sg13g2_decap_8 FILLER_46_1337 ();
 sg13g2_decap_8 FILLER_46_1344 ();
 sg13g2_decap_8 FILLER_46_1351 ();
 sg13g2_decap_8 FILLER_46_1358 ();
 sg13g2_decap_8 FILLER_46_1365 ();
 sg13g2_decap_8 FILLER_46_1372 ();
 sg13g2_decap_8 FILLER_46_1379 ();
 sg13g2_decap_8 FILLER_46_1386 ();
 sg13g2_decap_8 FILLER_46_1393 ();
 sg13g2_decap_8 FILLER_46_1400 ();
 sg13g2_decap_8 FILLER_46_1407 ();
 sg13g2_decap_8 FILLER_46_1414 ();
 sg13g2_decap_8 FILLER_46_1421 ();
 sg13g2_decap_8 FILLER_46_1428 ();
 sg13g2_decap_8 FILLER_46_1435 ();
 sg13g2_decap_8 FILLER_46_1442 ();
 sg13g2_decap_8 FILLER_46_1449 ();
 sg13g2_decap_8 FILLER_46_1456 ();
 sg13g2_decap_8 FILLER_46_1463 ();
 sg13g2_decap_8 FILLER_46_1470 ();
 sg13g2_decap_8 FILLER_46_1477 ();
 sg13g2_decap_8 FILLER_46_1484 ();
 sg13g2_decap_8 FILLER_46_1491 ();
 sg13g2_decap_8 FILLER_46_1498 ();
 sg13g2_decap_8 FILLER_46_1505 ();
 sg13g2_decap_8 FILLER_46_1512 ();
 sg13g2_decap_8 FILLER_46_1519 ();
 sg13g2_decap_8 FILLER_46_1526 ();
 sg13g2_decap_8 FILLER_46_1533 ();
 sg13g2_decap_8 FILLER_46_1540 ();
 sg13g2_decap_8 FILLER_46_1547 ();
 sg13g2_decap_8 FILLER_46_1554 ();
 sg13g2_decap_8 FILLER_46_1561 ();
 sg13g2_decap_8 FILLER_46_1568 ();
 sg13g2_decap_8 FILLER_46_1575 ();
 sg13g2_decap_8 FILLER_46_1582 ();
 sg13g2_decap_8 FILLER_46_1589 ();
 sg13g2_decap_8 FILLER_46_1596 ();
 sg13g2_decap_8 FILLER_46_1603 ();
 sg13g2_decap_8 FILLER_46_1610 ();
 sg13g2_decap_8 FILLER_46_1617 ();
 sg13g2_decap_8 FILLER_46_1624 ();
 sg13g2_decap_8 FILLER_46_1631 ();
 sg13g2_decap_8 FILLER_46_1638 ();
 sg13g2_decap_8 FILLER_46_1645 ();
 sg13g2_decap_8 FILLER_46_1652 ();
 sg13g2_decap_8 FILLER_46_1659 ();
 sg13g2_decap_8 FILLER_46_1666 ();
 sg13g2_decap_8 FILLER_46_1673 ();
 sg13g2_decap_8 FILLER_46_1680 ();
 sg13g2_decap_8 FILLER_46_1687 ();
 sg13g2_decap_8 FILLER_46_1694 ();
 sg13g2_decap_8 FILLER_46_1701 ();
 sg13g2_decap_8 FILLER_46_1708 ();
 sg13g2_decap_8 FILLER_46_1715 ();
 sg13g2_decap_8 FILLER_46_1722 ();
 sg13g2_decap_8 FILLER_46_1729 ();
 sg13g2_decap_8 FILLER_46_1736 ();
 sg13g2_decap_8 FILLER_46_1743 ();
 sg13g2_decap_8 FILLER_46_1750 ();
 sg13g2_decap_8 FILLER_46_1757 ();
 sg13g2_decap_8 FILLER_46_1764 ();
 sg13g2_decap_8 FILLER_46_1771 ();
 sg13g2_decap_8 FILLER_46_1778 ();
 sg13g2_decap_8 FILLER_46_1785 ();
 sg13g2_decap_8 FILLER_46_1792 ();
 sg13g2_decap_8 FILLER_46_1799 ();
 sg13g2_decap_8 FILLER_46_1806 ();
 sg13g2_decap_8 FILLER_46_1813 ();
 sg13g2_decap_8 FILLER_46_1820 ();
 sg13g2_decap_8 FILLER_46_1827 ();
 sg13g2_decap_8 FILLER_46_1834 ();
 sg13g2_decap_8 FILLER_46_1841 ();
 sg13g2_decap_8 FILLER_46_1848 ();
 sg13g2_decap_8 FILLER_46_1855 ();
 sg13g2_decap_8 FILLER_46_1862 ();
 sg13g2_decap_8 FILLER_46_1869 ();
 sg13g2_decap_8 FILLER_46_1876 ();
 sg13g2_decap_8 FILLER_46_1883 ();
 sg13g2_decap_8 FILLER_46_1890 ();
 sg13g2_decap_8 FILLER_46_1897 ();
 sg13g2_decap_8 FILLER_46_1904 ();
 sg13g2_decap_8 FILLER_46_1911 ();
 sg13g2_decap_8 FILLER_46_1918 ();
 sg13g2_decap_8 FILLER_46_1925 ();
 sg13g2_decap_8 FILLER_46_1932 ();
 sg13g2_decap_8 FILLER_46_1939 ();
 sg13g2_decap_8 FILLER_46_1946 ();
 sg13g2_decap_8 FILLER_46_1953 ();
 sg13g2_decap_8 FILLER_46_1960 ();
 sg13g2_decap_8 FILLER_46_1967 ();
 sg13g2_decap_8 FILLER_46_1974 ();
 sg13g2_decap_8 FILLER_46_1981 ();
 sg13g2_decap_8 FILLER_46_1988 ();
 sg13g2_decap_8 FILLER_46_1995 ();
 sg13g2_decap_8 FILLER_46_2002 ();
 sg13g2_decap_8 FILLER_46_2009 ();
 sg13g2_decap_8 FILLER_46_2016 ();
 sg13g2_decap_8 FILLER_46_2023 ();
 sg13g2_decap_8 FILLER_46_2030 ();
 sg13g2_decap_8 FILLER_46_2037 ();
 sg13g2_decap_8 FILLER_46_2044 ();
 sg13g2_decap_8 FILLER_46_2051 ();
 sg13g2_decap_8 FILLER_46_2058 ();
 sg13g2_decap_8 FILLER_46_2065 ();
 sg13g2_decap_8 FILLER_46_2072 ();
 sg13g2_decap_8 FILLER_46_2079 ();
 sg13g2_decap_8 FILLER_46_2086 ();
 sg13g2_decap_8 FILLER_46_2093 ();
 sg13g2_decap_8 FILLER_46_2100 ();
 sg13g2_decap_8 FILLER_46_2107 ();
 sg13g2_decap_8 FILLER_46_2114 ();
 sg13g2_decap_8 FILLER_46_2121 ();
 sg13g2_decap_8 FILLER_46_2128 ();
 sg13g2_decap_8 FILLER_46_2135 ();
 sg13g2_decap_8 FILLER_46_2142 ();
 sg13g2_decap_8 FILLER_46_2149 ();
 sg13g2_decap_8 FILLER_46_2156 ();
 sg13g2_decap_8 FILLER_46_2163 ();
 sg13g2_decap_8 FILLER_46_2170 ();
 sg13g2_decap_8 FILLER_46_2177 ();
 sg13g2_decap_8 FILLER_46_2184 ();
 sg13g2_decap_8 FILLER_46_2191 ();
 sg13g2_decap_8 FILLER_46_2198 ();
 sg13g2_decap_8 FILLER_46_2205 ();
 sg13g2_decap_8 FILLER_46_2212 ();
 sg13g2_decap_8 FILLER_46_2219 ();
 sg13g2_decap_8 FILLER_46_2226 ();
 sg13g2_decap_8 FILLER_46_2233 ();
 sg13g2_decap_8 FILLER_46_2240 ();
 sg13g2_decap_8 FILLER_46_2247 ();
 sg13g2_decap_8 FILLER_46_2254 ();
 sg13g2_decap_8 FILLER_46_2261 ();
 sg13g2_decap_8 FILLER_46_2268 ();
 sg13g2_decap_8 FILLER_46_2275 ();
 sg13g2_decap_8 FILLER_46_2282 ();
 sg13g2_decap_8 FILLER_46_2289 ();
 sg13g2_decap_8 FILLER_46_2296 ();
 sg13g2_decap_8 FILLER_46_2303 ();
 sg13g2_decap_8 FILLER_46_2310 ();
 sg13g2_decap_8 FILLER_46_2317 ();
 sg13g2_decap_8 FILLER_46_2324 ();
 sg13g2_decap_8 FILLER_46_2331 ();
 sg13g2_decap_8 FILLER_46_2338 ();
 sg13g2_decap_8 FILLER_46_2345 ();
 sg13g2_decap_8 FILLER_46_2352 ();
 sg13g2_decap_8 FILLER_46_2359 ();
 sg13g2_decap_8 FILLER_46_2366 ();
 sg13g2_decap_8 FILLER_46_2373 ();
 sg13g2_decap_8 FILLER_46_2380 ();
 sg13g2_decap_8 FILLER_46_2387 ();
 sg13g2_decap_8 FILLER_46_2394 ();
 sg13g2_decap_8 FILLER_46_2401 ();
 sg13g2_decap_8 FILLER_46_2408 ();
 sg13g2_decap_8 FILLER_46_2415 ();
 sg13g2_decap_8 FILLER_46_2422 ();
 sg13g2_decap_8 FILLER_46_2429 ();
 sg13g2_decap_8 FILLER_46_2436 ();
 sg13g2_decap_8 FILLER_46_2443 ();
 sg13g2_decap_8 FILLER_46_2450 ();
 sg13g2_decap_8 FILLER_46_2457 ();
 sg13g2_decap_8 FILLER_46_2464 ();
 sg13g2_decap_8 FILLER_46_2471 ();
 sg13g2_decap_8 FILLER_46_2478 ();
 sg13g2_decap_8 FILLER_46_2485 ();
 sg13g2_decap_8 FILLER_46_2492 ();
 sg13g2_decap_8 FILLER_46_2499 ();
 sg13g2_decap_8 FILLER_46_2506 ();
 sg13g2_decap_8 FILLER_46_2513 ();
 sg13g2_decap_8 FILLER_46_2520 ();
 sg13g2_decap_8 FILLER_46_2527 ();
 sg13g2_decap_8 FILLER_46_2534 ();
 sg13g2_decap_8 FILLER_46_2541 ();
 sg13g2_decap_8 FILLER_46_2548 ();
 sg13g2_decap_8 FILLER_46_2555 ();
 sg13g2_decap_8 FILLER_46_2562 ();
 sg13g2_decap_8 FILLER_46_2569 ();
 sg13g2_decap_8 FILLER_46_2576 ();
 sg13g2_decap_8 FILLER_46_2583 ();
 sg13g2_decap_8 FILLER_46_2590 ();
 sg13g2_decap_8 FILLER_46_2597 ();
 sg13g2_decap_8 FILLER_46_2604 ();
 sg13g2_decap_8 FILLER_46_2611 ();
 sg13g2_decap_8 FILLER_46_2618 ();
 sg13g2_decap_8 FILLER_46_2625 ();
 sg13g2_decap_8 FILLER_46_2632 ();
 sg13g2_decap_8 FILLER_46_2639 ();
 sg13g2_decap_8 FILLER_46_2646 ();
 sg13g2_decap_8 FILLER_46_2653 ();
 sg13g2_decap_8 FILLER_46_2660 ();
 sg13g2_decap_8 FILLER_46_2667 ();
 sg13g2_decap_8 FILLER_46_2674 ();
 sg13g2_decap_8 FILLER_46_2681 ();
 sg13g2_decap_8 FILLER_46_2688 ();
 sg13g2_decap_8 FILLER_46_2695 ();
 sg13g2_decap_8 FILLER_46_2702 ();
 sg13g2_decap_8 FILLER_46_2709 ();
 sg13g2_decap_8 FILLER_46_2716 ();
 sg13g2_decap_8 FILLER_46_2723 ();
 sg13g2_decap_8 FILLER_46_2730 ();
 sg13g2_decap_8 FILLER_46_2737 ();
 sg13g2_decap_8 FILLER_46_2744 ();
 sg13g2_decap_8 FILLER_46_2751 ();
 sg13g2_decap_8 FILLER_46_2758 ();
 sg13g2_decap_8 FILLER_46_2765 ();
 sg13g2_decap_8 FILLER_46_2772 ();
 sg13g2_decap_8 FILLER_46_2779 ();
 sg13g2_decap_8 FILLER_46_2786 ();
 sg13g2_decap_8 FILLER_46_2793 ();
 sg13g2_decap_8 FILLER_46_2800 ();
 sg13g2_decap_8 FILLER_46_2807 ();
 sg13g2_decap_8 FILLER_46_2814 ();
 sg13g2_decap_8 FILLER_46_2821 ();
 sg13g2_decap_8 FILLER_46_2828 ();
 sg13g2_decap_8 FILLER_46_2835 ();
 sg13g2_decap_8 FILLER_46_2842 ();
 sg13g2_decap_8 FILLER_46_2849 ();
 sg13g2_decap_8 FILLER_46_2856 ();
 sg13g2_decap_8 FILLER_46_2863 ();
 sg13g2_decap_8 FILLER_46_2870 ();
 sg13g2_decap_8 FILLER_46_2877 ();
 sg13g2_decap_8 FILLER_46_2884 ();
 sg13g2_decap_8 FILLER_46_2891 ();
 sg13g2_decap_8 FILLER_46_2898 ();
 sg13g2_decap_8 FILLER_46_2905 ();
 sg13g2_decap_8 FILLER_46_2912 ();
 sg13g2_decap_8 FILLER_46_2919 ();
 sg13g2_decap_8 FILLER_46_2926 ();
 sg13g2_decap_8 FILLER_46_2933 ();
 sg13g2_decap_8 FILLER_46_2940 ();
 sg13g2_decap_8 FILLER_46_2947 ();
 sg13g2_decap_8 FILLER_46_2954 ();
 sg13g2_decap_8 FILLER_46_2961 ();
 sg13g2_decap_8 FILLER_46_2968 ();
 sg13g2_decap_8 FILLER_46_2975 ();
 sg13g2_decap_8 FILLER_46_2982 ();
 sg13g2_decap_8 FILLER_46_2989 ();
 sg13g2_decap_8 FILLER_46_2996 ();
 sg13g2_decap_8 FILLER_46_3003 ();
 sg13g2_decap_8 FILLER_46_3010 ();
 sg13g2_decap_8 FILLER_46_3017 ();
 sg13g2_decap_8 FILLER_46_3024 ();
 sg13g2_decap_8 FILLER_46_3031 ();
 sg13g2_decap_8 FILLER_46_3038 ();
 sg13g2_decap_8 FILLER_46_3045 ();
 sg13g2_decap_8 FILLER_46_3052 ();
 sg13g2_decap_8 FILLER_46_3059 ();
 sg13g2_decap_8 FILLER_46_3066 ();
 sg13g2_decap_8 FILLER_46_3073 ();
 sg13g2_decap_8 FILLER_46_3080 ();
 sg13g2_decap_8 FILLER_46_3087 ();
 sg13g2_decap_8 FILLER_46_3094 ();
 sg13g2_decap_8 FILLER_46_3101 ();
 sg13g2_decap_8 FILLER_46_3108 ();
 sg13g2_decap_8 FILLER_46_3115 ();
 sg13g2_decap_8 FILLER_46_3122 ();
 sg13g2_decap_8 FILLER_46_3129 ();
 sg13g2_decap_8 FILLER_46_3136 ();
 sg13g2_decap_8 FILLER_46_3143 ();
 sg13g2_decap_8 FILLER_46_3150 ();
 sg13g2_decap_8 FILLER_46_3157 ();
 sg13g2_decap_8 FILLER_46_3164 ();
 sg13g2_decap_8 FILLER_46_3171 ();
 sg13g2_decap_8 FILLER_46_3178 ();
 sg13g2_decap_8 FILLER_46_3185 ();
 sg13g2_decap_8 FILLER_46_3192 ();
 sg13g2_decap_8 FILLER_46_3199 ();
 sg13g2_decap_8 FILLER_46_3206 ();
 sg13g2_decap_8 FILLER_46_3213 ();
 sg13g2_decap_8 FILLER_46_3220 ();
 sg13g2_decap_8 FILLER_46_3227 ();
 sg13g2_decap_8 FILLER_46_3234 ();
 sg13g2_decap_8 FILLER_46_3241 ();
 sg13g2_decap_8 FILLER_46_3248 ();
 sg13g2_decap_8 FILLER_46_3255 ();
 sg13g2_decap_8 FILLER_46_3262 ();
 sg13g2_decap_8 FILLER_46_3269 ();
 sg13g2_decap_8 FILLER_46_3276 ();
 sg13g2_decap_8 FILLER_46_3283 ();
 sg13g2_decap_8 FILLER_46_3290 ();
 sg13g2_decap_8 FILLER_46_3297 ();
 sg13g2_decap_8 FILLER_46_3304 ();
 sg13g2_decap_8 FILLER_46_3311 ();
 sg13g2_decap_8 FILLER_46_3318 ();
 sg13g2_decap_8 FILLER_46_3325 ();
 sg13g2_decap_8 FILLER_46_3332 ();
 sg13g2_decap_8 FILLER_46_3339 ();
 sg13g2_decap_8 FILLER_46_3346 ();
 sg13g2_decap_8 FILLER_46_3353 ();
 sg13g2_decap_8 FILLER_46_3360 ();
 sg13g2_decap_8 FILLER_46_3367 ();
 sg13g2_decap_8 FILLER_46_3374 ();
 sg13g2_decap_8 FILLER_46_3381 ();
 sg13g2_decap_8 FILLER_46_3388 ();
 sg13g2_decap_8 FILLER_46_3395 ();
 sg13g2_decap_8 FILLER_46_3402 ();
 sg13g2_decap_8 FILLER_46_3409 ();
 sg13g2_decap_8 FILLER_46_3416 ();
 sg13g2_decap_8 FILLER_46_3423 ();
 sg13g2_decap_8 FILLER_46_3430 ();
 sg13g2_decap_8 FILLER_46_3437 ();
 sg13g2_decap_8 FILLER_46_3444 ();
 sg13g2_decap_8 FILLER_46_3451 ();
 sg13g2_decap_8 FILLER_46_3458 ();
 sg13g2_decap_8 FILLER_46_3465 ();
 sg13g2_decap_8 FILLER_46_3472 ();
 sg13g2_decap_8 FILLER_46_3479 ();
 sg13g2_decap_8 FILLER_46_3486 ();
 sg13g2_decap_8 FILLER_46_3493 ();
 sg13g2_decap_8 FILLER_46_3500 ();
 sg13g2_decap_8 FILLER_46_3507 ();
 sg13g2_decap_8 FILLER_46_3514 ();
 sg13g2_decap_8 FILLER_46_3521 ();
 sg13g2_decap_8 FILLER_46_3528 ();
 sg13g2_decap_8 FILLER_46_3535 ();
 sg13g2_decap_8 FILLER_46_3542 ();
 sg13g2_decap_8 FILLER_46_3549 ();
 sg13g2_decap_8 FILLER_46_3556 ();
 sg13g2_decap_8 FILLER_46_3563 ();
 sg13g2_decap_8 FILLER_46_3570 ();
 sg13g2_fill_2 FILLER_46_3577 ();
 sg13g2_fill_1 FILLER_46_3579 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_decap_8 FILLER_47_175 ();
 sg13g2_decap_8 FILLER_47_182 ();
 sg13g2_decap_8 FILLER_47_189 ();
 sg13g2_decap_8 FILLER_47_196 ();
 sg13g2_decap_8 FILLER_47_203 ();
 sg13g2_decap_8 FILLER_47_210 ();
 sg13g2_decap_8 FILLER_47_217 ();
 sg13g2_decap_8 FILLER_47_224 ();
 sg13g2_decap_8 FILLER_47_231 ();
 sg13g2_decap_8 FILLER_47_238 ();
 sg13g2_decap_8 FILLER_47_245 ();
 sg13g2_decap_8 FILLER_47_252 ();
 sg13g2_decap_8 FILLER_47_259 ();
 sg13g2_decap_8 FILLER_47_266 ();
 sg13g2_decap_8 FILLER_47_273 ();
 sg13g2_decap_8 FILLER_47_280 ();
 sg13g2_decap_8 FILLER_47_287 ();
 sg13g2_decap_8 FILLER_47_294 ();
 sg13g2_decap_8 FILLER_47_301 ();
 sg13g2_decap_8 FILLER_47_308 ();
 sg13g2_decap_8 FILLER_47_315 ();
 sg13g2_decap_8 FILLER_47_322 ();
 sg13g2_decap_8 FILLER_47_329 ();
 sg13g2_decap_8 FILLER_47_336 ();
 sg13g2_decap_8 FILLER_47_343 ();
 sg13g2_decap_8 FILLER_47_350 ();
 sg13g2_decap_8 FILLER_47_357 ();
 sg13g2_decap_8 FILLER_47_364 ();
 sg13g2_decap_8 FILLER_47_371 ();
 sg13g2_decap_8 FILLER_47_378 ();
 sg13g2_decap_8 FILLER_47_385 ();
 sg13g2_decap_8 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_399 ();
 sg13g2_decap_8 FILLER_47_406 ();
 sg13g2_decap_8 FILLER_47_413 ();
 sg13g2_decap_8 FILLER_47_420 ();
 sg13g2_decap_8 FILLER_47_427 ();
 sg13g2_decap_8 FILLER_47_434 ();
 sg13g2_decap_8 FILLER_47_441 ();
 sg13g2_decap_8 FILLER_47_448 ();
 sg13g2_decap_8 FILLER_47_455 ();
 sg13g2_decap_8 FILLER_47_462 ();
 sg13g2_decap_8 FILLER_47_469 ();
 sg13g2_decap_8 FILLER_47_476 ();
 sg13g2_decap_8 FILLER_47_483 ();
 sg13g2_decap_8 FILLER_47_490 ();
 sg13g2_decap_8 FILLER_47_497 ();
 sg13g2_decap_8 FILLER_47_504 ();
 sg13g2_decap_8 FILLER_47_511 ();
 sg13g2_decap_8 FILLER_47_518 ();
 sg13g2_decap_8 FILLER_47_525 ();
 sg13g2_decap_8 FILLER_47_532 ();
 sg13g2_decap_8 FILLER_47_539 ();
 sg13g2_decap_8 FILLER_47_546 ();
 sg13g2_decap_8 FILLER_47_553 ();
 sg13g2_decap_8 FILLER_47_560 ();
 sg13g2_decap_8 FILLER_47_567 ();
 sg13g2_decap_8 FILLER_47_574 ();
 sg13g2_decap_8 FILLER_47_581 ();
 sg13g2_decap_8 FILLER_47_588 ();
 sg13g2_decap_8 FILLER_47_595 ();
 sg13g2_decap_8 FILLER_47_602 ();
 sg13g2_decap_8 FILLER_47_609 ();
 sg13g2_decap_8 FILLER_47_616 ();
 sg13g2_decap_8 FILLER_47_623 ();
 sg13g2_decap_8 FILLER_47_630 ();
 sg13g2_decap_8 FILLER_47_637 ();
 sg13g2_decap_8 FILLER_47_644 ();
 sg13g2_decap_8 FILLER_47_651 ();
 sg13g2_decap_8 FILLER_47_658 ();
 sg13g2_decap_8 FILLER_47_665 ();
 sg13g2_decap_8 FILLER_47_672 ();
 sg13g2_decap_8 FILLER_47_679 ();
 sg13g2_decap_8 FILLER_47_686 ();
 sg13g2_decap_8 FILLER_47_693 ();
 sg13g2_decap_8 FILLER_47_700 ();
 sg13g2_decap_8 FILLER_47_707 ();
 sg13g2_decap_8 FILLER_47_714 ();
 sg13g2_decap_8 FILLER_47_721 ();
 sg13g2_decap_8 FILLER_47_728 ();
 sg13g2_decap_8 FILLER_47_735 ();
 sg13g2_decap_8 FILLER_47_742 ();
 sg13g2_decap_8 FILLER_47_749 ();
 sg13g2_decap_8 FILLER_47_756 ();
 sg13g2_decap_8 FILLER_47_763 ();
 sg13g2_decap_8 FILLER_47_770 ();
 sg13g2_decap_8 FILLER_47_777 ();
 sg13g2_decap_8 FILLER_47_784 ();
 sg13g2_decap_8 FILLER_47_791 ();
 sg13g2_decap_8 FILLER_47_798 ();
 sg13g2_decap_8 FILLER_47_805 ();
 sg13g2_decap_8 FILLER_47_812 ();
 sg13g2_decap_8 FILLER_47_819 ();
 sg13g2_decap_8 FILLER_47_826 ();
 sg13g2_decap_8 FILLER_47_833 ();
 sg13g2_decap_8 FILLER_47_840 ();
 sg13g2_decap_8 FILLER_47_847 ();
 sg13g2_decap_8 FILLER_47_854 ();
 sg13g2_decap_8 FILLER_47_861 ();
 sg13g2_decap_8 FILLER_47_868 ();
 sg13g2_decap_8 FILLER_47_875 ();
 sg13g2_decap_8 FILLER_47_882 ();
 sg13g2_decap_8 FILLER_47_889 ();
 sg13g2_decap_8 FILLER_47_896 ();
 sg13g2_decap_8 FILLER_47_903 ();
 sg13g2_decap_8 FILLER_47_910 ();
 sg13g2_decap_8 FILLER_47_917 ();
 sg13g2_decap_8 FILLER_47_924 ();
 sg13g2_decap_8 FILLER_47_931 ();
 sg13g2_decap_8 FILLER_47_938 ();
 sg13g2_decap_8 FILLER_47_945 ();
 sg13g2_decap_8 FILLER_47_952 ();
 sg13g2_decap_8 FILLER_47_959 ();
 sg13g2_decap_8 FILLER_47_966 ();
 sg13g2_decap_8 FILLER_47_973 ();
 sg13g2_decap_8 FILLER_47_980 ();
 sg13g2_decap_8 FILLER_47_987 ();
 sg13g2_decap_8 FILLER_47_994 ();
 sg13g2_decap_8 FILLER_47_1001 ();
 sg13g2_decap_8 FILLER_47_1008 ();
 sg13g2_decap_8 FILLER_47_1015 ();
 sg13g2_decap_8 FILLER_47_1022 ();
 sg13g2_decap_8 FILLER_47_1029 ();
 sg13g2_decap_8 FILLER_47_1036 ();
 sg13g2_decap_8 FILLER_47_1043 ();
 sg13g2_decap_8 FILLER_47_1050 ();
 sg13g2_decap_8 FILLER_47_1057 ();
 sg13g2_decap_8 FILLER_47_1064 ();
 sg13g2_decap_8 FILLER_47_1071 ();
 sg13g2_decap_8 FILLER_47_1078 ();
 sg13g2_decap_8 FILLER_47_1085 ();
 sg13g2_decap_8 FILLER_47_1092 ();
 sg13g2_decap_8 FILLER_47_1099 ();
 sg13g2_decap_8 FILLER_47_1106 ();
 sg13g2_decap_8 FILLER_47_1113 ();
 sg13g2_decap_8 FILLER_47_1120 ();
 sg13g2_decap_8 FILLER_47_1127 ();
 sg13g2_decap_8 FILLER_47_1134 ();
 sg13g2_decap_8 FILLER_47_1141 ();
 sg13g2_decap_8 FILLER_47_1148 ();
 sg13g2_decap_8 FILLER_47_1155 ();
 sg13g2_decap_8 FILLER_47_1162 ();
 sg13g2_decap_8 FILLER_47_1169 ();
 sg13g2_decap_8 FILLER_47_1176 ();
 sg13g2_decap_8 FILLER_47_1183 ();
 sg13g2_decap_8 FILLER_47_1190 ();
 sg13g2_decap_8 FILLER_47_1197 ();
 sg13g2_decap_8 FILLER_47_1204 ();
 sg13g2_decap_8 FILLER_47_1211 ();
 sg13g2_decap_8 FILLER_47_1218 ();
 sg13g2_decap_8 FILLER_47_1225 ();
 sg13g2_decap_8 FILLER_47_1232 ();
 sg13g2_decap_8 FILLER_47_1239 ();
 sg13g2_decap_8 FILLER_47_1246 ();
 sg13g2_decap_8 FILLER_47_1253 ();
 sg13g2_decap_8 FILLER_47_1260 ();
 sg13g2_decap_8 FILLER_47_1267 ();
 sg13g2_decap_8 FILLER_47_1274 ();
 sg13g2_decap_8 FILLER_47_1281 ();
 sg13g2_decap_8 FILLER_47_1288 ();
 sg13g2_decap_8 FILLER_47_1295 ();
 sg13g2_decap_8 FILLER_47_1302 ();
 sg13g2_decap_8 FILLER_47_1309 ();
 sg13g2_decap_8 FILLER_47_1316 ();
 sg13g2_decap_8 FILLER_47_1323 ();
 sg13g2_decap_8 FILLER_47_1330 ();
 sg13g2_decap_8 FILLER_47_1337 ();
 sg13g2_decap_8 FILLER_47_1344 ();
 sg13g2_decap_8 FILLER_47_1351 ();
 sg13g2_decap_8 FILLER_47_1358 ();
 sg13g2_decap_8 FILLER_47_1365 ();
 sg13g2_decap_8 FILLER_47_1372 ();
 sg13g2_decap_8 FILLER_47_1379 ();
 sg13g2_decap_8 FILLER_47_1386 ();
 sg13g2_decap_8 FILLER_47_1393 ();
 sg13g2_decap_8 FILLER_47_1400 ();
 sg13g2_decap_8 FILLER_47_1407 ();
 sg13g2_decap_8 FILLER_47_1414 ();
 sg13g2_decap_8 FILLER_47_1421 ();
 sg13g2_decap_8 FILLER_47_1428 ();
 sg13g2_decap_8 FILLER_47_1435 ();
 sg13g2_decap_8 FILLER_47_1442 ();
 sg13g2_decap_8 FILLER_47_1449 ();
 sg13g2_decap_8 FILLER_47_1456 ();
 sg13g2_decap_8 FILLER_47_1463 ();
 sg13g2_decap_8 FILLER_47_1470 ();
 sg13g2_decap_8 FILLER_47_1477 ();
 sg13g2_decap_8 FILLER_47_1484 ();
 sg13g2_decap_8 FILLER_47_1491 ();
 sg13g2_decap_8 FILLER_47_1498 ();
 sg13g2_decap_8 FILLER_47_1505 ();
 sg13g2_decap_8 FILLER_47_1512 ();
 sg13g2_decap_8 FILLER_47_1519 ();
 sg13g2_decap_8 FILLER_47_1526 ();
 sg13g2_decap_8 FILLER_47_1533 ();
 sg13g2_decap_8 FILLER_47_1540 ();
 sg13g2_decap_8 FILLER_47_1547 ();
 sg13g2_decap_8 FILLER_47_1554 ();
 sg13g2_decap_8 FILLER_47_1561 ();
 sg13g2_decap_8 FILLER_47_1568 ();
 sg13g2_decap_8 FILLER_47_1575 ();
 sg13g2_decap_8 FILLER_47_1582 ();
 sg13g2_decap_8 FILLER_47_1589 ();
 sg13g2_decap_8 FILLER_47_1596 ();
 sg13g2_decap_8 FILLER_47_1603 ();
 sg13g2_decap_8 FILLER_47_1610 ();
 sg13g2_decap_8 FILLER_47_1617 ();
 sg13g2_decap_8 FILLER_47_1624 ();
 sg13g2_decap_8 FILLER_47_1631 ();
 sg13g2_decap_8 FILLER_47_1638 ();
 sg13g2_decap_8 FILLER_47_1645 ();
 sg13g2_decap_8 FILLER_47_1652 ();
 sg13g2_decap_8 FILLER_47_1659 ();
 sg13g2_decap_8 FILLER_47_1666 ();
 sg13g2_decap_8 FILLER_47_1673 ();
 sg13g2_decap_8 FILLER_47_1680 ();
 sg13g2_decap_8 FILLER_47_1687 ();
 sg13g2_decap_8 FILLER_47_1694 ();
 sg13g2_decap_8 FILLER_47_1701 ();
 sg13g2_decap_8 FILLER_47_1708 ();
 sg13g2_decap_8 FILLER_47_1715 ();
 sg13g2_decap_8 FILLER_47_1722 ();
 sg13g2_decap_8 FILLER_47_1729 ();
 sg13g2_decap_8 FILLER_47_1736 ();
 sg13g2_decap_8 FILLER_47_1743 ();
 sg13g2_decap_8 FILLER_47_1750 ();
 sg13g2_decap_8 FILLER_47_1757 ();
 sg13g2_decap_8 FILLER_47_1764 ();
 sg13g2_decap_8 FILLER_47_1771 ();
 sg13g2_decap_8 FILLER_47_1778 ();
 sg13g2_decap_8 FILLER_47_1785 ();
 sg13g2_decap_8 FILLER_47_1792 ();
 sg13g2_decap_8 FILLER_47_1799 ();
 sg13g2_decap_8 FILLER_47_1806 ();
 sg13g2_decap_8 FILLER_47_1813 ();
 sg13g2_decap_8 FILLER_47_1820 ();
 sg13g2_decap_8 FILLER_47_1827 ();
 sg13g2_decap_8 FILLER_47_1834 ();
 sg13g2_decap_8 FILLER_47_1841 ();
 sg13g2_decap_8 FILLER_47_1848 ();
 sg13g2_decap_8 FILLER_47_1855 ();
 sg13g2_decap_8 FILLER_47_1862 ();
 sg13g2_decap_8 FILLER_47_1869 ();
 sg13g2_decap_8 FILLER_47_1876 ();
 sg13g2_decap_8 FILLER_47_1883 ();
 sg13g2_decap_8 FILLER_47_1890 ();
 sg13g2_decap_8 FILLER_47_1897 ();
 sg13g2_decap_8 FILLER_47_1904 ();
 sg13g2_decap_8 FILLER_47_1911 ();
 sg13g2_decap_8 FILLER_47_1918 ();
 sg13g2_decap_8 FILLER_47_1925 ();
 sg13g2_decap_8 FILLER_47_1932 ();
 sg13g2_decap_8 FILLER_47_1939 ();
 sg13g2_decap_8 FILLER_47_1946 ();
 sg13g2_decap_8 FILLER_47_1953 ();
 sg13g2_decap_8 FILLER_47_1960 ();
 sg13g2_decap_8 FILLER_47_1967 ();
 sg13g2_decap_8 FILLER_47_1974 ();
 sg13g2_decap_8 FILLER_47_1981 ();
 sg13g2_decap_8 FILLER_47_1988 ();
 sg13g2_decap_8 FILLER_47_1995 ();
 sg13g2_decap_8 FILLER_47_2002 ();
 sg13g2_decap_8 FILLER_47_2009 ();
 sg13g2_decap_8 FILLER_47_2016 ();
 sg13g2_decap_8 FILLER_47_2023 ();
 sg13g2_decap_8 FILLER_47_2030 ();
 sg13g2_decap_8 FILLER_47_2037 ();
 sg13g2_decap_8 FILLER_47_2044 ();
 sg13g2_decap_8 FILLER_47_2051 ();
 sg13g2_decap_8 FILLER_47_2058 ();
 sg13g2_decap_8 FILLER_47_2065 ();
 sg13g2_decap_8 FILLER_47_2072 ();
 sg13g2_decap_8 FILLER_47_2079 ();
 sg13g2_decap_8 FILLER_47_2086 ();
 sg13g2_decap_8 FILLER_47_2093 ();
 sg13g2_decap_8 FILLER_47_2100 ();
 sg13g2_decap_8 FILLER_47_2107 ();
 sg13g2_decap_8 FILLER_47_2114 ();
 sg13g2_decap_8 FILLER_47_2121 ();
 sg13g2_decap_8 FILLER_47_2128 ();
 sg13g2_decap_8 FILLER_47_2135 ();
 sg13g2_decap_8 FILLER_47_2142 ();
 sg13g2_decap_8 FILLER_47_2149 ();
 sg13g2_decap_8 FILLER_47_2156 ();
 sg13g2_decap_8 FILLER_47_2163 ();
 sg13g2_decap_8 FILLER_47_2170 ();
 sg13g2_decap_8 FILLER_47_2177 ();
 sg13g2_decap_8 FILLER_47_2184 ();
 sg13g2_decap_8 FILLER_47_2191 ();
 sg13g2_decap_8 FILLER_47_2198 ();
 sg13g2_decap_8 FILLER_47_2205 ();
 sg13g2_decap_8 FILLER_47_2212 ();
 sg13g2_decap_8 FILLER_47_2219 ();
 sg13g2_decap_8 FILLER_47_2226 ();
 sg13g2_decap_8 FILLER_47_2233 ();
 sg13g2_decap_8 FILLER_47_2240 ();
 sg13g2_decap_8 FILLER_47_2247 ();
 sg13g2_decap_8 FILLER_47_2254 ();
 sg13g2_decap_8 FILLER_47_2261 ();
 sg13g2_decap_8 FILLER_47_2268 ();
 sg13g2_decap_8 FILLER_47_2275 ();
 sg13g2_decap_8 FILLER_47_2282 ();
 sg13g2_decap_8 FILLER_47_2289 ();
 sg13g2_decap_8 FILLER_47_2296 ();
 sg13g2_decap_8 FILLER_47_2303 ();
 sg13g2_decap_8 FILLER_47_2310 ();
 sg13g2_decap_8 FILLER_47_2317 ();
 sg13g2_decap_8 FILLER_47_2324 ();
 sg13g2_decap_8 FILLER_47_2331 ();
 sg13g2_decap_8 FILLER_47_2338 ();
 sg13g2_decap_8 FILLER_47_2345 ();
 sg13g2_decap_8 FILLER_47_2352 ();
 sg13g2_decap_8 FILLER_47_2359 ();
 sg13g2_decap_8 FILLER_47_2366 ();
 sg13g2_decap_8 FILLER_47_2373 ();
 sg13g2_decap_8 FILLER_47_2380 ();
 sg13g2_decap_8 FILLER_47_2387 ();
 sg13g2_decap_8 FILLER_47_2394 ();
 sg13g2_decap_8 FILLER_47_2401 ();
 sg13g2_decap_8 FILLER_47_2408 ();
 sg13g2_decap_8 FILLER_47_2415 ();
 sg13g2_decap_8 FILLER_47_2422 ();
 sg13g2_decap_8 FILLER_47_2429 ();
 sg13g2_decap_8 FILLER_47_2436 ();
 sg13g2_decap_8 FILLER_47_2443 ();
 sg13g2_decap_8 FILLER_47_2450 ();
 sg13g2_decap_8 FILLER_47_2457 ();
 sg13g2_decap_8 FILLER_47_2464 ();
 sg13g2_decap_8 FILLER_47_2471 ();
 sg13g2_decap_8 FILLER_47_2478 ();
 sg13g2_decap_8 FILLER_47_2485 ();
 sg13g2_decap_8 FILLER_47_2492 ();
 sg13g2_decap_8 FILLER_47_2499 ();
 sg13g2_decap_8 FILLER_47_2506 ();
 sg13g2_decap_8 FILLER_47_2513 ();
 sg13g2_decap_8 FILLER_47_2520 ();
 sg13g2_decap_8 FILLER_47_2527 ();
 sg13g2_decap_8 FILLER_47_2534 ();
 sg13g2_decap_8 FILLER_47_2541 ();
 sg13g2_decap_8 FILLER_47_2548 ();
 sg13g2_decap_8 FILLER_47_2555 ();
 sg13g2_decap_8 FILLER_47_2562 ();
 sg13g2_decap_8 FILLER_47_2569 ();
 sg13g2_decap_8 FILLER_47_2576 ();
 sg13g2_decap_8 FILLER_47_2583 ();
 sg13g2_decap_8 FILLER_47_2590 ();
 sg13g2_decap_8 FILLER_47_2597 ();
 sg13g2_decap_8 FILLER_47_2604 ();
 sg13g2_decap_8 FILLER_47_2611 ();
 sg13g2_decap_8 FILLER_47_2618 ();
 sg13g2_decap_8 FILLER_47_2625 ();
 sg13g2_decap_8 FILLER_47_2632 ();
 sg13g2_decap_8 FILLER_47_2639 ();
 sg13g2_decap_8 FILLER_47_2646 ();
 sg13g2_decap_8 FILLER_47_2653 ();
 sg13g2_decap_8 FILLER_47_2660 ();
 sg13g2_decap_8 FILLER_47_2667 ();
 sg13g2_decap_8 FILLER_47_2674 ();
 sg13g2_decap_8 FILLER_47_2681 ();
 sg13g2_decap_8 FILLER_47_2688 ();
 sg13g2_decap_8 FILLER_47_2695 ();
 sg13g2_decap_8 FILLER_47_2702 ();
 sg13g2_decap_8 FILLER_47_2709 ();
 sg13g2_decap_8 FILLER_47_2716 ();
 sg13g2_decap_8 FILLER_47_2723 ();
 sg13g2_decap_8 FILLER_47_2730 ();
 sg13g2_decap_8 FILLER_47_2737 ();
 sg13g2_decap_8 FILLER_47_2744 ();
 sg13g2_decap_8 FILLER_47_2751 ();
 sg13g2_decap_8 FILLER_47_2758 ();
 sg13g2_decap_8 FILLER_47_2765 ();
 sg13g2_decap_8 FILLER_47_2772 ();
 sg13g2_decap_8 FILLER_47_2779 ();
 sg13g2_decap_8 FILLER_47_2786 ();
 sg13g2_decap_8 FILLER_47_2793 ();
 sg13g2_decap_8 FILLER_47_2800 ();
 sg13g2_decap_8 FILLER_47_2807 ();
 sg13g2_decap_8 FILLER_47_2814 ();
 sg13g2_decap_8 FILLER_47_2821 ();
 sg13g2_decap_8 FILLER_47_2828 ();
 sg13g2_decap_8 FILLER_47_2835 ();
 sg13g2_decap_8 FILLER_47_2842 ();
 sg13g2_decap_8 FILLER_47_2849 ();
 sg13g2_decap_8 FILLER_47_2856 ();
 sg13g2_decap_8 FILLER_47_2863 ();
 sg13g2_decap_8 FILLER_47_2870 ();
 sg13g2_decap_8 FILLER_47_2877 ();
 sg13g2_decap_8 FILLER_47_2884 ();
 sg13g2_decap_8 FILLER_47_2891 ();
 sg13g2_decap_8 FILLER_47_2898 ();
 sg13g2_decap_8 FILLER_47_2905 ();
 sg13g2_decap_8 FILLER_47_2912 ();
 sg13g2_decap_8 FILLER_47_2919 ();
 sg13g2_decap_8 FILLER_47_2926 ();
 sg13g2_decap_8 FILLER_47_2933 ();
 sg13g2_decap_8 FILLER_47_2940 ();
 sg13g2_decap_8 FILLER_47_2947 ();
 sg13g2_decap_8 FILLER_47_2954 ();
 sg13g2_decap_8 FILLER_47_2961 ();
 sg13g2_decap_8 FILLER_47_2968 ();
 sg13g2_decap_8 FILLER_47_2975 ();
 sg13g2_decap_8 FILLER_47_2982 ();
 sg13g2_decap_8 FILLER_47_2989 ();
 sg13g2_decap_8 FILLER_47_2996 ();
 sg13g2_decap_8 FILLER_47_3003 ();
 sg13g2_decap_8 FILLER_47_3010 ();
 sg13g2_decap_8 FILLER_47_3017 ();
 sg13g2_decap_8 FILLER_47_3024 ();
 sg13g2_decap_8 FILLER_47_3031 ();
 sg13g2_decap_8 FILLER_47_3038 ();
 sg13g2_decap_8 FILLER_47_3045 ();
 sg13g2_decap_8 FILLER_47_3052 ();
 sg13g2_decap_8 FILLER_47_3059 ();
 sg13g2_decap_8 FILLER_47_3066 ();
 sg13g2_decap_8 FILLER_47_3073 ();
 sg13g2_decap_8 FILLER_47_3080 ();
 sg13g2_decap_8 FILLER_47_3087 ();
 sg13g2_decap_8 FILLER_47_3094 ();
 sg13g2_decap_8 FILLER_47_3101 ();
 sg13g2_decap_8 FILLER_47_3108 ();
 sg13g2_decap_8 FILLER_47_3115 ();
 sg13g2_decap_8 FILLER_47_3122 ();
 sg13g2_decap_8 FILLER_47_3129 ();
 sg13g2_decap_8 FILLER_47_3136 ();
 sg13g2_decap_8 FILLER_47_3143 ();
 sg13g2_decap_8 FILLER_47_3150 ();
 sg13g2_decap_8 FILLER_47_3157 ();
 sg13g2_decap_8 FILLER_47_3164 ();
 sg13g2_decap_8 FILLER_47_3171 ();
 sg13g2_decap_8 FILLER_47_3178 ();
 sg13g2_decap_8 FILLER_47_3185 ();
 sg13g2_decap_8 FILLER_47_3192 ();
 sg13g2_decap_8 FILLER_47_3199 ();
 sg13g2_decap_8 FILLER_47_3206 ();
 sg13g2_decap_8 FILLER_47_3213 ();
 sg13g2_decap_8 FILLER_47_3220 ();
 sg13g2_decap_8 FILLER_47_3227 ();
 sg13g2_decap_8 FILLER_47_3234 ();
 sg13g2_decap_8 FILLER_47_3241 ();
 sg13g2_decap_8 FILLER_47_3248 ();
 sg13g2_decap_8 FILLER_47_3255 ();
 sg13g2_decap_8 FILLER_47_3262 ();
 sg13g2_decap_8 FILLER_47_3269 ();
 sg13g2_decap_8 FILLER_47_3276 ();
 sg13g2_decap_8 FILLER_47_3283 ();
 sg13g2_decap_8 FILLER_47_3290 ();
 sg13g2_decap_8 FILLER_47_3297 ();
 sg13g2_decap_8 FILLER_47_3304 ();
 sg13g2_decap_8 FILLER_47_3311 ();
 sg13g2_decap_8 FILLER_47_3318 ();
 sg13g2_decap_8 FILLER_47_3325 ();
 sg13g2_decap_8 FILLER_47_3332 ();
 sg13g2_decap_8 FILLER_47_3339 ();
 sg13g2_decap_8 FILLER_47_3346 ();
 sg13g2_decap_8 FILLER_47_3353 ();
 sg13g2_decap_8 FILLER_47_3360 ();
 sg13g2_decap_8 FILLER_47_3367 ();
 sg13g2_decap_8 FILLER_47_3374 ();
 sg13g2_decap_8 FILLER_47_3381 ();
 sg13g2_decap_8 FILLER_47_3388 ();
 sg13g2_decap_8 FILLER_47_3395 ();
 sg13g2_decap_8 FILLER_47_3402 ();
 sg13g2_decap_8 FILLER_47_3409 ();
 sg13g2_decap_8 FILLER_47_3416 ();
 sg13g2_decap_8 FILLER_47_3423 ();
 sg13g2_decap_8 FILLER_47_3430 ();
 sg13g2_decap_8 FILLER_47_3437 ();
 sg13g2_decap_8 FILLER_47_3444 ();
 sg13g2_decap_8 FILLER_47_3451 ();
 sg13g2_decap_8 FILLER_47_3458 ();
 sg13g2_decap_8 FILLER_47_3465 ();
 sg13g2_decap_8 FILLER_47_3472 ();
 sg13g2_decap_8 FILLER_47_3479 ();
 sg13g2_decap_8 FILLER_47_3486 ();
 sg13g2_decap_8 FILLER_47_3493 ();
 sg13g2_decap_8 FILLER_47_3500 ();
 sg13g2_decap_8 FILLER_47_3507 ();
 sg13g2_decap_8 FILLER_47_3514 ();
 sg13g2_decap_8 FILLER_47_3521 ();
 sg13g2_decap_8 FILLER_47_3528 ();
 sg13g2_decap_8 FILLER_47_3535 ();
 sg13g2_decap_8 FILLER_47_3542 ();
 sg13g2_decap_8 FILLER_47_3549 ();
 sg13g2_decap_8 FILLER_47_3556 ();
 sg13g2_decap_8 FILLER_47_3563 ();
 sg13g2_decap_8 FILLER_47_3570 ();
 sg13g2_fill_2 FILLER_47_3577 ();
 sg13g2_fill_1 FILLER_47_3579 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_147 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_168 ();
 sg13g2_decap_8 FILLER_48_175 ();
 sg13g2_decap_8 FILLER_48_182 ();
 sg13g2_decap_8 FILLER_48_189 ();
 sg13g2_decap_8 FILLER_48_196 ();
 sg13g2_decap_8 FILLER_48_203 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_decap_8 FILLER_48_217 ();
 sg13g2_decap_8 FILLER_48_224 ();
 sg13g2_decap_8 FILLER_48_231 ();
 sg13g2_decap_8 FILLER_48_238 ();
 sg13g2_decap_8 FILLER_48_245 ();
 sg13g2_decap_8 FILLER_48_252 ();
 sg13g2_decap_8 FILLER_48_259 ();
 sg13g2_decap_8 FILLER_48_266 ();
 sg13g2_decap_8 FILLER_48_273 ();
 sg13g2_decap_8 FILLER_48_280 ();
 sg13g2_decap_8 FILLER_48_287 ();
 sg13g2_decap_8 FILLER_48_294 ();
 sg13g2_decap_8 FILLER_48_301 ();
 sg13g2_decap_8 FILLER_48_308 ();
 sg13g2_decap_8 FILLER_48_315 ();
 sg13g2_decap_8 FILLER_48_322 ();
 sg13g2_decap_8 FILLER_48_329 ();
 sg13g2_decap_8 FILLER_48_336 ();
 sg13g2_decap_8 FILLER_48_343 ();
 sg13g2_decap_8 FILLER_48_350 ();
 sg13g2_decap_8 FILLER_48_357 ();
 sg13g2_decap_8 FILLER_48_364 ();
 sg13g2_decap_8 FILLER_48_371 ();
 sg13g2_decap_8 FILLER_48_378 ();
 sg13g2_decap_8 FILLER_48_385 ();
 sg13g2_decap_8 FILLER_48_392 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_decap_8 FILLER_48_406 ();
 sg13g2_decap_8 FILLER_48_413 ();
 sg13g2_decap_8 FILLER_48_420 ();
 sg13g2_decap_8 FILLER_48_427 ();
 sg13g2_decap_8 FILLER_48_434 ();
 sg13g2_decap_8 FILLER_48_441 ();
 sg13g2_decap_8 FILLER_48_448 ();
 sg13g2_decap_8 FILLER_48_455 ();
 sg13g2_decap_8 FILLER_48_462 ();
 sg13g2_decap_8 FILLER_48_469 ();
 sg13g2_decap_8 FILLER_48_476 ();
 sg13g2_decap_8 FILLER_48_483 ();
 sg13g2_decap_8 FILLER_48_490 ();
 sg13g2_decap_8 FILLER_48_497 ();
 sg13g2_decap_8 FILLER_48_504 ();
 sg13g2_decap_8 FILLER_48_511 ();
 sg13g2_decap_8 FILLER_48_518 ();
 sg13g2_decap_8 FILLER_48_525 ();
 sg13g2_decap_8 FILLER_48_532 ();
 sg13g2_decap_8 FILLER_48_539 ();
 sg13g2_decap_8 FILLER_48_546 ();
 sg13g2_decap_8 FILLER_48_553 ();
 sg13g2_decap_8 FILLER_48_560 ();
 sg13g2_decap_8 FILLER_48_567 ();
 sg13g2_decap_8 FILLER_48_574 ();
 sg13g2_decap_8 FILLER_48_581 ();
 sg13g2_decap_8 FILLER_48_588 ();
 sg13g2_decap_8 FILLER_48_595 ();
 sg13g2_decap_8 FILLER_48_602 ();
 sg13g2_decap_8 FILLER_48_609 ();
 sg13g2_decap_8 FILLER_48_616 ();
 sg13g2_decap_8 FILLER_48_623 ();
 sg13g2_decap_8 FILLER_48_630 ();
 sg13g2_decap_8 FILLER_48_637 ();
 sg13g2_decap_8 FILLER_48_644 ();
 sg13g2_decap_8 FILLER_48_651 ();
 sg13g2_decap_8 FILLER_48_658 ();
 sg13g2_decap_8 FILLER_48_665 ();
 sg13g2_decap_8 FILLER_48_672 ();
 sg13g2_decap_8 FILLER_48_679 ();
 sg13g2_decap_8 FILLER_48_686 ();
 sg13g2_decap_8 FILLER_48_693 ();
 sg13g2_decap_8 FILLER_48_700 ();
 sg13g2_decap_8 FILLER_48_707 ();
 sg13g2_decap_8 FILLER_48_714 ();
 sg13g2_decap_8 FILLER_48_721 ();
 sg13g2_decap_8 FILLER_48_728 ();
 sg13g2_decap_8 FILLER_48_735 ();
 sg13g2_decap_8 FILLER_48_742 ();
 sg13g2_decap_8 FILLER_48_749 ();
 sg13g2_decap_8 FILLER_48_756 ();
 sg13g2_decap_8 FILLER_48_763 ();
 sg13g2_decap_8 FILLER_48_770 ();
 sg13g2_decap_8 FILLER_48_777 ();
 sg13g2_decap_8 FILLER_48_784 ();
 sg13g2_decap_8 FILLER_48_791 ();
 sg13g2_decap_8 FILLER_48_798 ();
 sg13g2_decap_8 FILLER_48_805 ();
 sg13g2_decap_8 FILLER_48_812 ();
 sg13g2_decap_8 FILLER_48_819 ();
 sg13g2_decap_8 FILLER_48_826 ();
 sg13g2_decap_8 FILLER_48_833 ();
 sg13g2_decap_8 FILLER_48_840 ();
 sg13g2_decap_8 FILLER_48_847 ();
 sg13g2_decap_8 FILLER_48_854 ();
 sg13g2_decap_8 FILLER_48_861 ();
 sg13g2_decap_8 FILLER_48_868 ();
 sg13g2_decap_8 FILLER_48_875 ();
 sg13g2_decap_8 FILLER_48_882 ();
 sg13g2_decap_8 FILLER_48_889 ();
 sg13g2_decap_8 FILLER_48_896 ();
 sg13g2_decap_8 FILLER_48_903 ();
 sg13g2_decap_8 FILLER_48_910 ();
 sg13g2_decap_8 FILLER_48_917 ();
 sg13g2_decap_8 FILLER_48_924 ();
 sg13g2_decap_8 FILLER_48_931 ();
 sg13g2_decap_8 FILLER_48_938 ();
 sg13g2_decap_8 FILLER_48_945 ();
 sg13g2_decap_8 FILLER_48_952 ();
 sg13g2_decap_8 FILLER_48_959 ();
 sg13g2_decap_8 FILLER_48_966 ();
 sg13g2_decap_8 FILLER_48_973 ();
 sg13g2_decap_8 FILLER_48_980 ();
 sg13g2_decap_8 FILLER_48_987 ();
 sg13g2_decap_8 FILLER_48_994 ();
 sg13g2_decap_8 FILLER_48_1001 ();
 sg13g2_decap_8 FILLER_48_1008 ();
 sg13g2_decap_8 FILLER_48_1015 ();
 sg13g2_decap_8 FILLER_48_1022 ();
 sg13g2_decap_8 FILLER_48_1029 ();
 sg13g2_decap_8 FILLER_48_1036 ();
 sg13g2_decap_8 FILLER_48_1043 ();
 sg13g2_decap_8 FILLER_48_1050 ();
 sg13g2_decap_8 FILLER_48_1057 ();
 sg13g2_decap_8 FILLER_48_1064 ();
 sg13g2_decap_8 FILLER_48_1071 ();
 sg13g2_decap_8 FILLER_48_1078 ();
 sg13g2_decap_8 FILLER_48_1085 ();
 sg13g2_decap_8 FILLER_48_1092 ();
 sg13g2_decap_8 FILLER_48_1099 ();
 sg13g2_decap_8 FILLER_48_1106 ();
 sg13g2_decap_8 FILLER_48_1113 ();
 sg13g2_decap_8 FILLER_48_1120 ();
 sg13g2_decap_8 FILLER_48_1127 ();
 sg13g2_decap_8 FILLER_48_1134 ();
 sg13g2_decap_8 FILLER_48_1141 ();
 sg13g2_decap_8 FILLER_48_1148 ();
 sg13g2_decap_8 FILLER_48_1155 ();
 sg13g2_decap_8 FILLER_48_1162 ();
 sg13g2_decap_8 FILLER_48_1169 ();
 sg13g2_decap_8 FILLER_48_1176 ();
 sg13g2_decap_8 FILLER_48_1183 ();
 sg13g2_decap_8 FILLER_48_1190 ();
 sg13g2_decap_8 FILLER_48_1197 ();
 sg13g2_decap_8 FILLER_48_1204 ();
 sg13g2_decap_8 FILLER_48_1211 ();
 sg13g2_decap_8 FILLER_48_1218 ();
 sg13g2_decap_8 FILLER_48_1225 ();
 sg13g2_decap_8 FILLER_48_1232 ();
 sg13g2_decap_8 FILLER_48_1239 ();
 sg13g2_decap_8 FILLER_48_1246 ();
 sg13g2_decap_8 FILLER_48_1253 ();
 sg13g2_decap_8 FILLER_48_1260 ();
 sg13g2_decap_8 FILLER_48_1267 ();
 sg13g2_decap_8 FILLER_48_1274 ();
 sg13g2_decap_8 FILLER_48_1281 ();
 sg13g2_decap_8 FILLER_48_1288 ();
 sg13g2_decap_8 FILLER_48_1295 ();
 sg13g2_decap_8 FILLER_48_1302 ();
 sg13g2_decap_8 FILLER_48_1309 ();
 sg13g2_decap_8 FILLER_48_1316 ();
 sg13g2_decap_8 FILLER_48_1323 ();
 sg13g2_decap_8 FILLER_48_1330 ();
 sg13g2_decap_8 FILLER_48_1337 ();
 sg13g2_decap_8 FILLER_48_1344 ();
 sg13g2_decap_8 FILLER_48_1351 ();
 sg13g2_decap_8 FILLER_48_1358 ();
 sg13g2_decap_8 FILLER_48_1365 ();
 sg13g2_decap_8 FILLER_48_1372 ();
 sg13g2_decap_8 FILLER_48_1379 ();
 sg13g2_decap_8 FILLER_48_1386 ();
 sg13g2_decap_8 FILLER_48_1393 ();
 sg13g2_decap_8 FILLER_48_1400 ();
 sg13g2_decap_8 FILLER_48_1407 ();
 sg13g2_decap_8 FILLER_48_1414 ();
 sg13g2_decap_8 FILLER_48_1421 ();
 sg13g2_decap_8 FILLER_48_1428 ();
 sg13g2_decap_8 FILLER_48_1435 ();
 sg13g2_decap_8 FILLER_48_1442 ();
 sg13g2_decap_8 FILLER_48_1449 ();
 sg13g2_decap_8 FILLER_48_1456 ();
 sg13g2_decap_8 FILLER_48_1463 ();
 sg13g2_decap_8 FILLER_48_1470 ();
 sg13g2_decap_8 FILLER_48_1477 ();
 sg13g2_decap_8 FILLER_48_1484 ();
 sg13g2_decap_8 FILLER_48_1491 ();
 sg13g2_decap_8 FILLER_48_1498 ();
 sg13g2_decap_8 FILLER_48_1505 ();
 sg13g2_decap_8 FILLER_48_1512 ();
 sg13g2_decap_8 FILLER_48_1519 ();
 sg13g2_decap_8 FILLER_48_1526 ();
 sg13g2_decap_8 FILLER_48_1533 ();
 sg13g2_decap_8 FILLER_48_1540 ();
 sg13g2_decap_8 FILLER_48_1547 ();
 sg13g2_decap_8 FILLER_48_1554 ();
 sg13g2_decap_8 FILLER_48_1561 ();
 sg13g2_decap_8 FILLER_48_1568 ();
 sg13g2_decap_8 FILLER_48_1575 ();
 sg13g2_decap_8 FILLER_48_1582 ();
 sg13g2_decap_8 FILLER_48_1589 ();
 sg13g2_decap_8 FILLER_48_1596 ();
 sg13g2_decap_8 FILLER_48_1603 ();
 sg13g2_decap_8 FILLER_48_1610 ();
 sg13g2_decap_8 FILLER_48_1617 ();
 sg13g2_decap_8 FILLER_48_1624 ();
 sg13g2_decap_8 FILLER_48_1631 ();
 sg13g2_decap_8 FILLER_48_1638 ();
 sg13g2_decap_8 FILLER_48_1645 ();
 sg13g2_decap_8 FILLER_48_1652 ();
 sg13g2_decap_8 FILLER_48_1659 ();
 sg13g2_decap_8 FILLER_48_1666 ();
 sg13g2_decap_8 FILLER_48_1673 ();
 sg13g2_decap_8 FILLER_48_1680 ();
 sg13g2_decap_8 FILLER_48_1687 ();
 sg13g2_decap_8 FILLER_48_1694 ();
 sg13g2_decap_8 FILLER_48_1701 ();
 sg13g2_decap_8 FILLER_48_1708 ();
 sg13g2_decap_8 FILLER_48_1715 ();
 sg13g2_decap_8 FILLER_48_1722 ();
 sg13g2_decap_8 FILLER_48_1729 ();
 sg13g2_decap_8 FILLER_48_1736 ();
 sg13g2_decap_8 FILLER_48_1743 ();
 sg13g2_decap_8 FILLER_48_1750 ();
 sg13g2_decap_8 FILLER_48_1757 ();
 sg13g2_decap_8 FILLER_48_1764 ();
 sg13g2_decap_8 FILLER_48_1771 ();
 sg13g2_decap_8 FILLER_48_1778 ();
 sg13g2_decap_8 FILLER_48_1785 ();
 sg13g2_decap_8 FILLER_48_1792 ();
 sg13g2_decap_8 FILLER_48_1799 ();
 sg13g2_decap_8 FILLER_48_1806 ();
 sg13g2_decap_8 FILLER_48_1813 ();
 sg13g2_decap_8 FILLER_48_1820 ();
 sg13g2_decap_8 FILLER_48_1827 ();
 sg13g2_decap_8 FILLER_48_1834 ();
 sg13g2_decap_8 FILLER_48_1841 ();
 sg13g2_decap_8 FILLER_48_1848 ();
 sg13g2_decap_8 FILLER_48_1855 ();
 sg13g2_decap_8 FILLER_48_1862 ();
 sg13g2_decap_8 FILLER_48_1869 ();
 sg13g2_decap_8 FILLER_48_1876 ();
 sg13g2_decap_8 FILLER_48_1883 ();
 sg13g2_decap_8 FILLER_48_1890 ();
 sg13g2_decap_8 FILLER_48_1897 ();
 sg13g2_decap_8 FILLER_48_1904 ();
 sg13g2_decap_8 FILLER_48_1911 ();
 sg13g2_decap_8 FILLER_48_1918 ();
 sg13g2_decap_8 FILLER_48_1925 ();
 sg13g2_decap_8 FILLER_48_1932 ();
 sg13g2_decap_8 FILLER_48_1939 ();
 sg13g2_decap_8 FILLER_48_1946 ();
 sg13g2_decap_8 FILLER_48_1953 ();
 sg13g2_decap_8 FILLER_48_1960 ();
 sg13g2_decap_8 FILLER_48_1967 ();
 sg13g2_decap_8 FILLER_48_1974 ();
 sg13g2_decap_8 FILLER_48_1981 ();
 sg13g2_decap_8 FILLER_48_1988 ();
 sg13g2_decap_8 FILLER_48_1995 ();
 sg13g2_decap_8 FILLER_48_2002 ();
 sg13g2_decap_8 FILLER_48_2009 ();
 sg13g2_decap_8 FILLER_48_2016 ();
 sg13g2_decap_8 FILLER_48_2023 ();
 sg13g2_decap_8 FILLER_48_2030 ();
 sg13g2_decap_8 FILLER_48_2037 ();
 sg13g2_decap_8 FILLER_48_2044 ();
 sg13g2_decap_8 FILLER_48_2051 ();
 sg13g2_decap_8 FILLER_48_2058 ();
 sg13g2_decap_8 FILLER_48_2065 ();
 sg13g2_decap_8 FILLER_48_2072 ();
 sg13g2_decap_8 FILLER_48_2079 ();
 sg13g2_decap_8 FILLER_48_2086 ();
 sg13g2_decap_8 FILLER_48_2093 ();
 sg13g2_decap_8 FILLER_48_2100 ();
 sg13g2_decap_8 FILLER_48_2107 ();
 sg13g2_decap_8 FILLER_48_2114 ();
 sg13g2_decap_8 FILLER_48_2121 ();
 sg13g2_decap_8 FILLER_48_2128 ();
 sg13g2_decap_8 FILLER_48_2135 ();
 sg13g2_decap_8 FILLER_48_2142 ();
 sg13g2_decap_8 FILLER_48_2149 ();
 sg13g2_decap_8 FILLER_48_2156 ();
 sg13g2_decap_8 FILLER_48_2163 ();
 sg13g2_decap_8 FILLER_48_2170 ();
 sg13g2_decap_8 FILLER_48_2177 ();
 sg13g2_decap_8 FILLER_48_2184 ();
 sg13g2_decap_8 FILLER_48_2191 ();
 sg13g2_decap_8 FILLER_48_2198 ();
 sg13g2_decap_8 FILLER_48_2205 ();
 sg13g2_decap_8 FILLER_48_2212 ();
 sg13g2_decap_8 FILLER_48_2219 ();
 sg13g2_decap_8 FILLER_48_2226 ();
 sg13g2_decap_8 FILLER_48_2233 ();
 sg13g2_decap_8 FILLER_48_2240 ();
 sg13g2_decap_8 FILLER_48_2247 ();
 sg13g2_decap_8 FILLER_48_2254 ();
 sg13g2_decap_8 FILLER_48_2261 ();
 sg13g2_decap_8 FILLER_48_2268 ();
 sg13g2_decap_8 FILLER_48_2275 ();
 sg13g2_decap_8 FILLER_48_2282 ();
 sg13g2_decap_8 FILLER_48_2289 ();
 sg13g2_decap_8 FILLER_48_2296 ();
 sg13g2_decap_8 FILLER_48_2303 ();
 sg13g2_decap_8 FILLER_48_2310 ();
 sg13g2_decap_8 FILLER_48_2317 ();
 sg13g2_decap_8 FILLER_48_2324 ();
 sg13g2_decap_8 FILLER_48_2331 ();
 sg13g2_decap_8 FILLER_48_2338 ();
 sg13g2_decap_8 FILLER_48_2345 ();
 sg13g2_decap_8 FILLER_48_2352 ();
 sg13g2_decap_8 FILLER_48_2359 ();
 sg13g2_decap_8 FILLER_48_2366 ();
 sg13g2_decap_8 FILLER_48_2373 ();
 sg13g2_decap_8 FILLER_48_2380 ();
 sg13g2_decap_8 FILLER_48_2387 ();
 sg13g2_decap_8 FILLER_48_2394 ();
 sg13g2_decap_8 FILLER_48_2401 ();
 sg13g2_decap_8 FILLER_48_2408 ();
 sg13g2_decap_8 FILLER_48_2415 ();
 sg13g2_decap_8 FILLER_48_2422 ();
 sg13g2_decap_8 FILLER_48_2429 ();
 sg13g2_decap_8 FILLER_48_2436 ();
 sg13g2_decap_8 FILLER_48_2443 ();
 sg13g2_decap_8 FILLER_48_2450 ();
 sg13g2_decap_8 FILLER_48_2457 ();
 sg13g2_decap_8 FILLER_48_2464 ();
 sg13g2_decap_8 FILLER_48_2471 ();
 sg13g2_decap_8 FILLER_48_2478 ();
 sg13g2_decap_8 FILLER_48_2485 ();
 sg13g2_decap_8 FILLER_48_2492 ();
 sg13g2_decap_8 FILLER_48_2499 ();
 sg13g2_decap_8 FILLER_48_2506 ();
 sg13g2_decap_8 FILLER_48_2513 ();
 sg13g2_decap_8 FILLER_48_2520 ();
 sg13g2_decap_8 FILLER_48_2527 ();
 sg13g2_decap_8 FILLER_48_2534 ();
 sg13g2_decap_8 FILLER_48_2541 ();
 sg13g2_decap_8 FILLER_48_2548 ();
 sg13g2_decap_8 FILLER_48_2555 ();
 sg13g2_decap_8 FILLER_48_2562 ();
 sg13g2_decap_8 FILLER_48_2569 ();
 sg13g2_decap_8 FILLER_48_2576 ();
 sg13g2_decap_8 FILLER_48_2583 ();
 sg13g2_decap_8 FILLER_48_2590 ();
 sg13g2_decap_8 FILLER_48_2597 ();
 sg13g2_decap_8 FILLER_48_2604 ();
 sg13g2_decap_8 FILLER_48_2611 ();
 sg13g2_decap_8 FILLER_48_2618 ();
 sg13g2_decap_8 FILLER_48_2625 ();
 sg13g2_decap_8 FILLER_48_2632 ();
 sg13g2_decap_8 FILLER_48_2639 ();
 sg13g2_decap_8 FILLER_48_2646 ();
 sg13g2_decap_8 FILLER_48_2653 ();
 sg13g2_decap_8 FILLER_48_2660 ();
 sg13g2_decap_8 FILLER_48_2667 ();
 sg13g2_decap_8 FILLER_48_2674 ();
 sg13g2_decap_8 FILLER_48_2681 ();
 sg13g2_decap_8 FILLER_48_2688 ();
 sg13g2_decap_8 FILLER_48_2695 ();
 sg13g2_decap_8 FILLER_48_2702 ();
 sg13g2_decap_8 FILLER_48_2709 ();
 sg13g2_decap_8 FILLER_48_2716 ();
 sg13g2_decap_8 FILLER_48_2723 ();
 sg13g2_decap_8 FILLER_48_2730 ();
 sg13g2_decap_8 FILLER_48_2737 ();
 sg13g2_decap_8 FILLER_48_2744 ();
 sg13g2_decap_8 FILLER_48_2751 ();
 sg13g2_decap_8 FILLER_48_2758 ();
 sg13g2_decap_8 FILLER_48_2765 ();
 sg13g2_decap_8 FILLER_48_2772 ();
 sg13g2_decap_8 FILLER_48_2779 ();
 sg13g2_decap_8 FILLER_48_2786 ();
 sg13g2_decap_8 FILLER_48_2793 ();
 sg13g2_decap_8 FILLER_48_2800 ();
 sg13g2_decap_8 FILLER_48_2807 ();
 sg13g2_decap_8 FILLER_48_2814 ();
 sg13g2_decap_8 FILLER_48_2821 ();
 sg13g2_decap_8 FILLER_48_2828 ();
 sg13g2_decap_8 FILLER_48_2835 ();
 sg13g2_decap_8 FILLER_48_2842 ();
 sg13g2_decap_8 FILLER_48_2849 ();
 sg13g2_decap_8 FILLER_48_2856 ();
 sg13g2_decap_8 FILLER_48_2863 ();
 sg13g2_decap_8 FILLER_48_2870 ();
 sg13g2_decap_8 FILLER_48_2877 ();
 sg13g2_decap_8 FILLER_48_2884 ();
 sg13g2_decap_8 FILLER_48_2891 ();
 sg13g2_decap_8 FILLER_48_2898 ();
 sg13g2_decap_8 FILLER_48_2905 ();
 sg13g2_decap_8 FILLER_48_2912 ();
 sg13g2_decap_8 FILLER_48_2919 ();
 sg13g2_decap_8 FILLER_48_2926 ();
 sg13g2_decap_8 FILLER_48_2933 ();
 sg13g2_decap_8 FILLER_48_2940 ();
 sg13g2_decap_8 FILLER_48_2947 ();
 sg13g2_decap_8 FILLER_48_2954 ();
 sg13g2_decap_8 FILLER_48_2961 ();
 sg13g2_decap_8 FILLER_48_2968 ();
 sg13g2_decap_8 FILLER_48_2975 ();
 sg13g2_decap_8 FILLER_48_2982 ();
 sg13g2_decap_8 FILLER_48_2989 ();
 sg13g2_decap_8 FILLER_48_2996 ();
 sg13g2_decap_8 FILLER_48_3003 ();
 sg13g2_decap_8 FILLER_48_3010 ();
 sg13g2_decap_8 FILLER_48_3017 ();
 sg13g2_decap_8 FILLER_48_3024 ();
 sg13g2_decap_8 FILLER_48_3031 ();
 sg13g2_decap_8 FILLER_48_3038 ();
 sg13g2_decap_8 FILLER_48_3045 ();
 sg13g2_decap_8 FILLER_48_3052 ();
 sg13g2_decap_8 FILLER_48_3059 ();
 sg13g2_decap_8 FILLER_48_3066 ();
 sg13g2_decap_8 FILLER_48_3073 ();
 sg13g2_decap_8 FILLER_48_3080 ();
 sg13g2_decap_8 FILLER_48_3087 ();
 sg13g2_decap_8 FILLER_48_3094 ();
 sg13g2_decap_8 FILLER_48_3101 ();
 sg13g2_decap_8 FILLER_48_3108 ();
 sg13g2_decap_8 FILLER_48_3115 ();
 sg13g2_decap_8 FILLER_48_3122 ();
 sg13g2_decap_8 FILLER_48_3129 ();
 sg13g2_decap_8 FILLER_48_3136 ();
 sg13g2_decap_8 FILLER_48_3143 ();
 sg13g2_decap_8 FILLER_48_3150 ();
 sg13g2_decap_8 FILLER_48_3157 ();
 sg13g2_decap_8 FILLER_48_3164 ();
 sg13g2_decap_8 FILLER_48_3171 ();
 sg13g2_decap_8 FILLER_48_3178 ();
 sg13g2_decap_8 FILLER_48_3185 ();
 sg13g2_decap_8 FILLER_48_3192 ();
 sg13g2_decap_8 FILLER_48_3199 ();
 sg13g2_decap_8 FILLER_48_3206 ();
 sg13g2_decap_8 FILLER_48_3213 ();
 sg13g2_decap_8 FILLER_48_3220 ();
 sg13g2_decap_8 FILLER_48_3227 ();
 sg13g2_decap_8 FILLER_48_3234 ();
 sg13g2_decap_8 FILLER_48_3241 ();
 sg13g2_decap_8 FILLER_48_3248 ();
 sg13g2_decap_8 FILLER_48_3255 ();
 sg13g2_decap_8 FILLER_48_3262 ();
 sg13g2_decap_8 FILLER_48_3269 ();
 sg13g2_decap_8 FILLER_48_3276 ();
 sg13g2_decap_8 FILLER_48_3283 ();
 sg13g2_decap_8 FILLER_48_3290 ();
 sg13g2_decap_8 FILLER_48_3297 ();
 sg13g2_decap_8 FILLER_48_3304 ();
 sg13g2_decap_8 FILLER_48_3311 ();
 sg13g2_decap_8 FILLER_48_3318 ();
 sg13g2_decap_8 FILLER_48_3325 ();
 sg13g2_decap_8 FILLER_48_3332 ();
 sg13g2_decap_8 FILLER_48_3339 ();
 sg13g2_decap_8 FILLER_48_3346 ();
 sg13g2_decap_8 FILLER_48_3353 ();
 sg13g2_decap_8 FILLER_48_3360 ();
 sg13g2_decap_8 FILLER_48_3367 ();
 sg13g2_decap_8 FILLER_48_3374 ();
 sg13g2_decap_8 FILLER_48_3381 ();
 sg13g2_decap_8 FILLER_48_3388 ();
 sg13g2_decap_8 FILLER_48_3395 ();
 sg13g2_decap_8 FILLER_48_3402 ();
 sg13g2_decap_8 FILLER_48_3409 ();
 sg13g2_decap_8 FILLER_48_3416 ();
 sg13g2_decap_8 FILLER_48_3423 ();
 sg13g2_decap_8 FILLER_48_3430 ();
 sg13g2_decap_8 FILLER_48_3437 ();
 sg13g2_decap_8 FILLER_48_3444 ();
 sg13g2_decap_8 FILLER_48_3451 ();
 sg13g2_decap_8 FILLER_48_3458 ();
 sg13g2_decap_8 FILLER_48_3465 ();
 sg13g2_decap_8 FILLER_48_3472 ();
 sg13g2_decap_8 FILLER_48_3479 ();
 sg13g2_decap_8 FILLER_48_3486 ();
 sg13g2_decap_8 FILLER_48_3493 ();
 sg13g2_decap_8 FILLER_48_3500 ();
 sg13g2_decap_8 FILLER_48_3507 ();
 sg13g2_decap_8 FILLER_48_3514 ();
 sg13g2_decap_8 FILLER_48_3521 ();
 sg13g2_decap_8 FILLER_48_3528 ();
 sg13g2_decap_8 FILLER_48_3535 ();
 sg13g2_decap_8 FILLER_48_3542 ();
 sg13g2_decap_8 FILLER_48_3549 ();
 sg13g2_decap_8 FILLER_48_3556 ();
 sg13g2_decap_8 FILLER_48_3563 ();
 sg13g2_decap_8 FILLER_48_3570 ();
 sg13g2_fill_2 FILLER_48_3577 ();
 sg13g2_fill_1 FILLER_48_3579 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_decap_8 FILLER_49_133 ();
 sg13g2_decap_8 FILLER_49_140 ();
 sg13g2_decap_8 FILLER_49_147 ();
 sg13g2_decap_8 FILLER_49_154 ();
 sg13g2_decap_8 FILLER_49_161 ();
 sg13g2_decap_8 FILLER_49_168 ();
 sg13g2_decap_8 FILLER_49_175 ();
 sg13g2_decap_8 FILLER_49_182 ();
 sg13g2_decap_8 FILLER_49_189 ();
 sg13g2_decap_8 FILLER_49_196 ();
 sg13g2_decap_8 FILLER_49_203 ();
 sg13g2_decap_8 FILLER_49_210 ();
 sg13g2_decap_8 FILLER_49_217 ();
 sg13g2_decap_8 FILLER_49_224 ();
 sg13g2_decap_8 FILLER_49_231 ();
 sg13g2_decap_8 FILLER_49_238 ();
 sg13g2_decap_8 FILLER_49_245 ();
 sg13g2_decap_8 FILLER_49_252 ();
 sg13g2_decap_8 FILLER_49_259 ();
 sg13g2_decap_8 FILLER_49_266 ();
 sg13g2_decap_8 FILLER_49_273 ();
 sg13g2_decap_8 FILLER_49_280 ();
 sg13g2_decap_8 FILLER_49_287 ();
 sg13g2_decap_8 FILLER_49_294 ();
 sg13g2_decap_8 FILLER_49_301 ();
 sg13g2_decap_8 FILLER_49_308 ();
 sg13g2_decap_8 FILLER_49_315 ();
 sg13g2_decap_8 FILLER_49_322 ();
 sg13g2_decap_8 FILLER_49_329 ();
 sg13g2_decap_8 FILLER_49_336 ();
 sg13g2_decap_8 FILLER_49_343 ();
 sg13g2_decap_8 FILLER_49_350 ();
 sg13g2_decap_8 FILLER_49_357 ();
 sg13g2_decap_8 FILLER_49_364 ();
 sg13g2_decap_8 FILLER_49_371 ();
 sg13g2_decap_8 FILLER_49_378 ();
 sg13g2_decap_8 FILLER_49_385 ();
 sg13g2_decap_8 FILLER_49_392 ();
 sg13g2_decap_8 FILLER_49_399 ();
 sg13g2_decap_8 FILLER_49_406 ();
 sg13g2_decap_8 FILLER_49_413 ();
 sg13g2_decap_8 FILLER_49_420 ();
 sg13g2_decap_8 FILLER_49_427 ();
 sg13g2_decap_8 FILLER_49_434 ();
 sg13g2_decap_8 FILLER_49_441 ();
 sg13g2_decap_8 FILLER_49_448 ();
 sg13g2_decap_8 FILLER_49_455 ();
 sg13g2_decap_8 FILLER_49_462 ();
 sg13g2_decap_8 FILLER_49_469 ();
 sg13g2_decap_8 FILLER_49_476 ();
 sg13g2_decap_8 FILLER_49_483 ();
 sg13g2_decap_8 FILLER_49_490 ();
 sg13g2_decap_8 FILLER_49_497 ();
 sg13g2_decap_8 FILLER_49_504 ();
 sg13g2_decap_8 FILLER_49_511 ();
 sg13g2_decap_8 FILLER_49_518 ();
 sg13g2_decap_8 FILLER_49_525 ();
 sg13g2_decap_8 FILLER_49_532 ();
 sg13g2_decap_8 FILLER_49_539 ();
 sg13g2_decap_8 FILLER_49_546 ();
 sg13g2_decap_8 FILLER_49_553 ();
 sg13g2_decap_8 FILLER_49_560 ();
 sg13g2_decap_8 FILLER_49_567 ();
 sg13g2_decap_8 FILLER_49_574 ();
 sg13g2_decap_8 FILLER_49_581 ();
 sg13g2_decap_8 FILLER_49_588 ();
 sg13g2_decap_8 FILLER_49_595 ();
 sg13g2_decap_8 FILLER_49_602 ();
 sg13g2_decap_8 FILLER_49_609 ();
 sg13g2_decap_8 FILLER_49_616 ();
 sg13g2_decap_8 FILLER_49_623 ();
 sg13g2_decap_8 FILLER_49_630 ();
 sg13g2_decap_8 FILLER_49_637 ();
 sg13g2_decap_8 FILLER_49_644 ();
 sg13g2_decap_8 FILLER_49_651 ();
 sg13g2_decap_8 FILLER_49_658 ();
 sg13g2_decap_8 FILLER_49_665 ();
 sg13g2_decap_8 FILLER_49_672 ();
 sg13g2_decap_8 FILLER_49_679 ();
 sg13g2_decap_8 FILLER_49_686 ();
 sg13g2_decap_8 FILLER_49_693 ();
 sg13g2_decap_8 FILLER_49_700 ();
 sg13g2_decap_8 FILLER_49_707 ();
 sg13g2_decap_8 FILLER_49_714 ();
 sg13g2_decap_8 FILLER_49_721 ();
 sg13g2_decap_8 FILLER_49_728 ();
 sg13g2_decap_8 FILLER_49_735 ();
 sg13g2_decap_8 FILLER_49_742 ();
 sg13g2_decap_8 FILLER_49_749 ();
 sg13g2_decap_8 FILLER_49_756 ();
 sg13g2_decap_8 FILLER_49_763 ();
 sg13g2_decap_8 FILLER_49_770 ();
 sg13g2_decap_8 FILLER_49_777 ();
 sg13g2_decap_8 FILLER_49_784 ();
 sg13g2_decap_8 FILLER_49_791 ();
 sg13g2_decap_8 FILLER_49_798 ();
 sg13g2_decap_8 FILLER_49_805 ();
 sg13g2_decap_8 FILLER_49_812 ();
 sg13g2_decap_8 FILLER_49_819 ();
 sg13g2_decap_8 FILLER_49_826 ();
 sg13g2_decap_8 FILLER_49_833 ();
 sg13g2_decap_8 FILLER_49_840 ();
 sg13g2_decap_8 FILLER_49_847 ();
 sg13g2_decap_8 FILLER_49_854 ();
 sg13g2_decap_8 FILLER_49_861 ();
 sg13g2_decap_8 FILLER_49_868 ();
 sg13g2_decap_8 FILLER_49_875 ();
 sg13g2_decap_8 FILLER_49_882 ();
 sg13g2_decap_8 FILLER_49_889 ();
 sg13g2_decap_8 FILLER_49_896 ();
 sg13g2_decap_8 FILLER_49_903 ();
 sg13g2_decap_8 FILLER_49_910 ();
 sg13g2_decap_8 FILLER_49_917 ();
 sg13g2_decap_8 FILLER_49_924 ();
 sg13g2_decap_8 FILLER_49_931 ();
 sg13g2_decap_8 FILLER_49_938 ();
 sg13g2_decap_8 FILLER_49_945 ();
 sg13g2_decap_8 FILLER_49_952 ();
 sg13g2_decap_8 FILLER_49_959 ();
 sg13g2_decap_8 FILLER_49_966 ();
 sg13g2_decap_8 FILLER_49_973 ();
 sg13g2_decap_8 FILLER_49_980 ();
 sg13g2_decap_8 FILLER_49_987 ();
 sg13g2_decap_8 FILLER_49_994 ();
 sg13g2_decap_8 FILLER_49_1001 ();
 sg13g2_decap_8 FILLER_49_1008 ();
 sg13g2_decap_8 FILLER_49_1015 ();
 sg13g2_decap_8 FILLER_49_1022 ();
 sg13g2_decap_8 FILLER_49_1029 ();
 sg13g2_decap_8 FILLER_49_1036 ();
 sg13g2_decap_8 FILLER_49_1043 ();
 sg13g2_decap_8 FILLER_49_1050 ();
 sg13g2_decap_8 FILLER_49_1057 ();
 sg13g2_decap_8 FILLER_49_1064 ();
 sg13g2_decap_8 FILLER_49_1071 ();
 sg13g2_decap_8 FILLER_49_1078 ();
 sg13g2_decap_8 FILLER_49_1085 ();
 sg13g2_decap_8 FILLER_49_1092 ();
 sg13g2_decap_8 FILLER_49_1099 ();
 sg13g2_decap_8 FILLER_49_1106 ();
 sg13g2_decap_8 FILLER_49_1113 ();
 sg13g2_decap_8 FILLER_49_1120 ();
 sg13g2_decap_8 FILLER_49_1127 ();
 sg13g2_decap_8 FILLER_49_1134 ();
 sg13g2_decap_8 FILLER_49_1141 ();
 sg13g2_decap_8 FILLER_49_1148 ();
 sg13g2_decap_8 FILLER_49_1155 ();
 sg13g2_decap_8 FILLER_49_1162 ();
 sg13g2_decap_8 FILLER_49_1169 ();
 sg13g2_decap_8 FILLER_49_1176 ();
 sg13g2_decap_8 FILLER_49_1183 ();
 sg13g2_decap_8 FILLER_49_1190 ();
 sg13g2_decap_8 FILLER_49_1197 ();
 sg13g2_decap_8 FILLER_49_1204 ();
 sg13g2_decap_8 FILLER_49_1211 ();
 sg13g2_decap_8 FILLER_49_1218 ();
 sg13g2_decap_8 FILLER_49_1225 ();
 sg13g2_decap_8 FILLER_49_1232 ();
 sg13g2_decap_8 FILLER_49_1239 ();
 sg13g2_decap_8 FILLER_49_1246 ();
 sg13g2_decap_8 FILLER_49_1253 ();
 sg13g2_decap_8 FILLER_49_1260 ();
 sg13g2_decap_8 FILLER_49_1267 ();
 sg13g2_decap_8 FILLER_49_1274 ();
 sg13g2_decap_8 FILLER_49_1281 ();
 sg13g2_decap_8 FILLER_49_1288 ();
 sg13g2_decap_8 FILLER_49_1295 ();
 sg13g2_decap_8 FILLER_49_1302 ();
 sg13g2_decap_8 FILLER_49_1309 ();
 sg13g2_decap_8 FILLER_49_1316 ();
 sg13g2_decap_8 FILLER_49_1323 ();
 sg13g2_decap_8 FILLER_49_1330 ();
 sg13g2_decap_8 FILLER_49_1337 ();
 sg13g2_decap_8 FILLER_49_1344 ();
 sg13g2_decap_8 FILLER_49_1351 ();
 sg13g2_decap_8 FILLER_49_1358 ();
 sg13g2_decap_8 FILLER_49_1365 ();
 sg13g2_decap_8 FILLER_49_1372 ();
 sg13g2_decap_8 FILLER_49_1379 ();
 sg13g2_decap_8 FILLER_49_1386 ();
 sg13g2_decap_8 FILLER_49_1393 ();
 sg13g2_decap_8 FILLER_49_1400 ();
 sg13g2_decap_8 FILLER_49_1407 ();
 sg13g2_decap_8 FILLER_49_1414 ();
 sg13g2_decap_8 FILLER_49_1421 ();
 sg13g2_decap_8 FILLER_49_1428 ();
 sg13g2_decap_8 FILLER_49_1435 ();
 sg13g2_decap_8 FILLER_49_1442 ();
 sg13g2_decap_8 FILLER_49_1449 ();
 sg13g2_decap_8 FILLER_49_1456 ();
 sg13g2_decap_8 FILLER_49_1463 ();
 sg13g2_decap_8 FILLER_49_1470 ();
 sg13g2_decap_8 FILLER_49_1477 ();
 sg13g2_decap_8 FILLER_49_1484 ();
 sg13g2_decap_8 FILLER_49_1491 ();
 sg13g2_decap_8 FILLER_49_1498 ();
 sg13g2_decap_8 FILLER_49_1505 ();
 sg13g2_decap_8 FILLER_49_1512 ();
 sg13g2_decap_8 FILLER_49_1519 ();
 sg13g2_decap_8 FILLER_49_1526 ();
 sg13g2_decap_8 FILLER_49_1533 ();
 sg13g2_decap_8 FILLER_49_1540 ();
 sg13g2_decap_8 FILLER_49_1547 ();
 sg13g2_decap_8 FILLER_49_1554 ();
 sg13g2_decap_8 FILLER_49_1561 ();
 sg13g2_decap_8 FILLER_49_1568 ();
 sg13g2_decap_8 FILLER_49_1575 ();
 sg13g2_decap_8 FILLER_49_1582 ();
 sg13g2_decap_8 FILLER_49_1589 ();
 sg13g2_decap_8 FILLER_49_1596 ();
 sg13g2_decap_8 FILLER_49_1603 ();
 sg13g2_decap_8 FILLER_49_1610 ();
 sg13g2_decap_8 FILLER_49_1617 ();
 sg13g2_decap_8 FILLER_49_1624 ();
 sg13g2_decap_8 FILLER_49_1631 ();
 sg13g2_decap_8 FILLER_49_1638 ();
 sg13g2_decap_8 FILLER_49_1645 ();
 sg13g2_decap_8 FILLER_49_1652 ();
 sg13g2_decap_8 FILLER_49_1659 ();
 sg13g2_decap_8 FILLER_49_1666 ();
 sg13g2_decap_8 FILLER_49_1673 ();
 sg13g2_decap_8 FILLER_49_1680 ();
 sg13g2_decap_8 FILLER_49_1687 ();
 sg13g2_decap_8 FILLER_49_1694 ();
 sg13g2_decap_8 FILLER_49_1701 ();
 sg13g2_decap_8 FILLER_49_1708 ();
 sg13g2_decap_8 FILLER_49_1715 ();
 sg13g2_decap_8 FILLER_49_1722 ();
 sg13g2_decap_8 FILLER_49_1729 ();
 sg13g2_decap_8 FILLER_49_1736 ();
 sg13g2_decap_8 FILLER_49_1743 ();
 sg13g2_decap_8 FILLER_49_1750 ();
 sg13g2_decap_8 FILLER_49_1757 ();
 sg13g2_decap_8 FILLER_49_1764 ();
 sg13g2_decap_8 FILLER_49_1771 ();
 sg13g2_decap_8 FILLER_49_1778 ();
 sg13g2_decap_8 FILLER_49_1785 ();
 sg13g2_decap_8 FILLER_49_1792 ();
 sg13g2_decap_8 FILLER_49_1799 ();
 sg13g2_decap_8 FILLER_49_1806 ();
 sg13g2_decap_8 FILLER_49_1813 ();
 sg13g2_decap_8 FILLER_49_1820 ();
 sg13g2_decap_8 FILLER_49_1827 ();
 sg13g2_decap_8 FILLER_49_1834 ();
 sg13g2_decap_8 FILLER_49_1841 ();
 sg13g2_decap_8 FILLER_49_1848 ();
 sg13g2_decap_8 FILLER_49_1855 ();
 sg13g2_decap_8 FILLER_49_1862 ();
 sg13g2_decap_8 FILLER_49_1869 ();
 sg13g2_decap_8 FILLER_49_1876 ();
 sg13g2_decap_8 FILLER_49_1883 ();
 sg13g2_decap_8 FILLER_49_1890 ();
 sg13g2_decap_8 FILLER_49_1897 ();
 sg13g2_decap_8 FILLER_49_1904 ();
 sg13g2_decap_8 FILLER_49_1911 ();
 sg13g2_decap_8 FILLER_49_1918 ();
 sg13g2_decap_8 FILLER_49_1925 ();
 sg13g2_decap_8 FILLER_49_1932 ();
 sg13g2_decap_8 FILLER_49_1939 ();
 sg13g2_decap_8 FILLER_49_1946 ();
 sg13g2_decap_8 FILLER_49_1953 ();
 sg13g2_decap_8 FILLER_49_1960 ();
 sg13g2_decap_8 FILLER_49_1967 ();
 sg13g2_decap_8 FILLER_49_1974 ();
 sg13g2_decap_8 FILLER_49_1981 ();
 sg13g2_decap_8 FILLER_49_1988 ();
 sg13g2_decap_8 FILLER_49_1995 ();
 sg13g2_decap_8 FILLER_49_2002 ();
 sg13g2_decap_8 FILLER_49_2009 ();
 sg13g2_decap_8 FILLER_49_2016 ();
 sg13g2_decap_8 FILLER_49_2023 ();
 sg13g2_decap_8 FILLER_49_2030 ();
 sg13g2_decap_8 FILLER_49_2037 ();
 sg13g2_decap_8 FILLER_49_2044 ();
 sg13g2_decap_8 FILLER_49_2051 ();
 sg13g2_decap_8 FILLER_49_2058 ();
 sg13g2_decap_8 FILLER_49_2065 ();
 sg13g2_decap_8 FILLER_49_2072 ();
 sg13g2_decap_8 FILLER_49_2079 ();
 sg13g2_decap_8 FILLER_49_2086 ();
 sg13g2_decap_8 FILLER_49_2093 ();
 sg13g2_decap_8 FILLER_49_2100 ();
 sg13g2_decap_8 FILLER_49_2107 ();
 sg13g2_decap_8 FILLER_49_2114 ();
 sg13g2_decap_8 FILLER_49_2121 ();
 sg13g2_decap_8 FILLER_49_2128 ();
 sg13g2_decap_8 FILLER_49_2135 ();
 sg13g2_decap_8 FILLER_49_2142 ();
 sg13g2_decap_8 FILLER_49_2149 ();
 sg13g2_decap_8 FILLER_49_2156 ();
 sg13g2_decap_8 FILLER_49_2163 ();
 sg13g2_decap_8 FILLER_49_2170 ();
 sg13g2_decap_8 FILLER_49_2177 ();
 sg13g2_decap_8 FILLER_49_2184 ();
 sg13g2_decap_8 FILLER_49_2191 ();
 sg13g2_decap_8 FILLER_49_2198 ();
 sg13g2_decap_8 FILLER_49_2205 ();
 sg13g2_decap_8 FILLER_49_2212 ();
 sg13g2_decap_8 FILLER_49_2219 ();
 sg13g2_decap_8 FILLER_49_2226 ();
 sg13g2_decap_8 FILLER_49_2233 ();
 sg13g2_decap_8 FILLER_49_2240 ();
 sg13g2_decap_8 FILLER_49_2247 ();
 sg13g2_decap_8 FILLER_49_2254 ();
 sg13g2_decap_8 FILLER_49_2261 ();
 sg13g2_decap_8 FILLER_49_2268 ();
 sg13g2_decap_8 FILLER_49_2275 ();
 sg13g2_decap_8 FILLER_49_2282 ();
 sg13g2_decap_8 FILLER_49_2289 ();
 sg13g2_decap_8 FILLER_49_2296 ();
 sg13g2_decap_8 FILLER_49_2303 ();
 sg13g2_decap_8 FILLER_49_2310 ();
 sg13g2_decap_8 FILLER_49_2317 ();
 sg13g2_decap_8 FILLER_49_2324 ();
 sg13g2_decap_8 FILLER_49_2331 ();
 sg13g2_decap_8 FILLER_49_2338 ();
 sg13g2_decap_8 FILLER_49_2345 ();
 sg13g2_decap_8 FILLER_49_2352 ();
 sg13g2_decap_8 FILLER_49_2359 ();
 sg13g2_decap_8 FILLER_49_2366 ();
 sg13g2_decap_8 FILLER_49_2373 ();
 sg13g2_decap_8 FILLER_49_2380 ();
 sg13g2_decap_8 FILLER_49_2387 ();
 sg13g2_decap_8 FILLER_49_2394 ();
 sg13g2_decap_8 FILLER_49_2401 ();
 sg13g2_decap_8 FILLER_49_2408 ();
 sg13g2_decap_8 FILLER_49_2415 ();
 sg13g2_decap_8 FILLER_49_2422 ();
 sg13g2_decap_8 FILLER_49_2429 ();
 sg13g2_decap_8 FILLER_49_2436 ();
 sg13g2_decap_8 FILLER_49_2443 ();
 sg13g2_decap_8 FILLER_49_2450 ();
 sg13g2_decap_8 FILLER_49_2457 ();
 sg13g2_decap_8 FILLER_49_2464 ();
 sg13g2_decap_8 FILLER_49_2471 ();
 sg13g2_decap_8 FILLER_49_2478 ();
 sg13g2_decap_8 FILLER_49_2485 ();
 sg13g2_decap_8 FILLER_49_2492 ();
 sg13g2_decap_8 FILLER_49_2499 ();
 sg13g2_decap_8 FILLER_49_2506 ();
 sg13g2_decap_8 FILLER_49_2513 ();
 sg13g2_decap_8 FILLER_49_2520 ();
 sg13g2_decap_8 FILLER_49_2527 ();
 sg13g2_decap_8 FILLER_49_2534 ();
 sg13g2_decap_8 FILLER_49_2541 ();
 sg13g2_decap_8 FILLER_49_2548 ();
 sg13g2_decap_8 FILLER_49_2555 ();
 sg13g2_decap_8 FILLER_49_2562 ();
 sg13g2_decap_8 FILLER_49_2569 ();
 sg13g2_decap_8 FILLER_49_2576 ();
 sg13g2_decap_8 FILLER_49_2583 ();
 sg13g2_decap_8 FILLER_49_2590 ();
 sg13g2_decap_8 FILLER_49_2597 ();
 sg13g2_decap_8 FILLER_49_2604 ();
 sg13g2_decap_8 FILLER_49_2611 ();
 sg13g2_decap_8 FILLER_49_2618 ();
 sg13g2_decap_8 FILLER_49_2625 ();
 sg13g2_decap_8 FILLER_49_2632 ();
 sg13g2_decap_8 FILLER_49_2639 ();
 sg13g2_decap_8 FILLER_49_2646 ();
 sg13g2_decap_8 FILLER_49_2653 ();
 sg13g2_decap_8 FILLER_49_2660 ();
 sg13g2_decap_8 FILLER_49_2667 ();
 sg13g2_decap_8 FILLER_49_2674 ();
 sg13g2_decap_8 FILLER_49_2681 ();
 sg13g2_decap_8 FILLER_49_2688 ();
 sg13g2_decap_8 FILLER_49_2695 ();
 sg13g2_decap_8 FILLER_49_2702 ();
 sg13g2_decap_8 FILLER_49_2709 ();
 sg13g2_decap_8 FILLER_49_2716 ();
 sg13g2_decap_8 FILLER_49_2723 ();
 sg13g2_decap_8 FILLER_49_2730 ();
 sg13g2_decap_8 FILLER_49_2737 ();
 sg13g2_decap_8 FILLER_49_2744 ();
 sg13g2_decap_8 FILLER_49_2751 ();
 sg13g2_decap_8 FILLER_49_2758 ();
 sg13g2_decap_8 FILLER_49_2765 ();
 sg13g2_decap_8 FILLER_49_2772 ();
 sg13g2_decap_8 FILLER_49_2779 ();
 sg13g2_decap_8 FILLER_49_2786 ();
 sg13g2_decap_8 FILLER_49_2793 ();
 sg13g2_decap_8 FILLER_49_2800 ();
 sg13g2_decap_8 FILLER_49_2807 ();
 sg13g2_decap_8 FILLER_49_2814 ();
 sg13g2_decap_8 FILLER_49_2821 ();
 sg13g2_decap_8 FILLER_49_2828 ();
 sg13g2_decap_8 FILLER_49_2835 ();
 sg13g2_decap_8 FILLER_49_2842 ();
 sg13g2_decap_8 FILLER_49_2849 ();
 sg13g2_decap_8 FILLER_49_2856 ();
 sg13g2_decap_8 FILLER_49_2863 ();
 sg13g2_decap_8 FILLER_49_2870 ();
 sg13g2_decap_8 FILLER_49_2877 ();
 sg13g2_decap_8 FILLER_49_2884 ();
 sg13g2_decap_8 FILLER_49_2891 ();
 sg13g2_decap_8 FILLER_49_2898 ();
 sg13g2_decap_8 FILLER_49_2905 ();
 sg13g2_decap_8 FILLER_49_2912 ();
 sg13g2_decap_8 FILLER_49_2919 ();
 sg13g2_decap_8 FILLER_49_2926 ();
 sg13g2_decap_8 FILLER_49_2933 ();
 sg13g2_decap_8 FILLER_49_2940 ();
 sg13g2_decap_8 FILLER_49_2947 ();
 sg13g2_decap_8 FILLER_49_2954 ();
 sg13g2_decap_8 FILLER_49_2961 ();
 sg13g2_decap_8 FILLER_49_2968 ();
 sg13g2_decap_8 FILLER_49_2975 ();
 sg13g2_decap_8 FILLER_49_2982 ();
 sg13g2_decap_8 FILLER_49_2989 ();
 sg13g2_decap_8 FILLER_49_2996 ();
 sg13g2_decap_8 FILLER_49_3003 ();
 sg13g2_decap_8 FILLER_49_3010 ();
 sg13g2_decap_8 FILLER_49_3017 ();
 sg13g2_decap_8 FILLER_49_3024 ();
 sg13g2_decap_8 FILLER_49_3031 ();
 sg13g2_decap_8 FILLER_49_3038 ();
 sg13g2_decap_8 FILLER_49_3045 ();
 sg13g2_decap_8 FILLER_49_3052 ();
 sg13g2_decap_8 FILLER_49_3059 ();
 sg13g2_decap_8 FILLER_49_3066 ();
 sg13g2_decap_8 FILLER_49_3073 ();
 sg13g2_decap_8 FILLER_49_3080 ();
 sg13g2_decap_8 FILLER_49_3087 ();
 sg13g2_decap_8 FILLER_49_3094 ();
 sg13g2_decap_8 FILLER_49_3101 ();
 sg13g2_decap_8 FILLER_49_3108 ();
 sg13g2_decap_8 FILLER_49_3115 ();
 sg13g2_decap_8 FILLER_49_3122 ();
 sg13g2_decap_8 FILLER_49_3129 ();
 sg13g2_decap_8 FILLER_49_3136 ();
 sg13g2_decap_8 FILLER_49_3143 ();
 sg13g2_decap_8 FILLER_49_3150 ();
 sg13g2_decap_8 FILLER_49_3157 ();
 sg13g2_decap_8 FILLER_49_3164 ();
 sg13g2_decap_8 FILLER_49_3171 ();
 sg13g2_decap_8 FILLER_49_3178 ();
 sg13g2_decap_8 FILLER_49_3185 ();
 sg13g2_decap_8 FILLER_49_3192 ();
 sg13g2_decap_8 FILLER_49_3199 ();
 sg13g2_decap_8 FILLER_49_3206 ();
 sg13g2_decap_8 FILLER_49_3213 ();
 sg13g2_decap_8 FILLER_49_3220 ();
 sg13g2_decap_8 FILLER_49_3227 ();
 sg13g2_decap_8 FILLER_49_3234 ();
 sg13g2_decap_8 FILLER_49_3241 ();
 sg13g2_decap_8 FILLER_49_3248 ();
 sg13g2_decap_8 FILLER_49_3255 ();
 sg13g2_decap_8 FILLER_49_3262 ();
 sg13g2_decap_8 FILLER_49_3269 ();
 sg13g2_decap_8 FILLER_49_3276 ();
 sg13g2_decap_8 FILLER_49_3283 ();
 sg13g2_decap_8 FILLER_49_3290 ();
 sg13g2_decap_8 FILLER_49_3297 ();
 sg13g2_decap_8 FILLER_49_3304 ();
 sg13g2_decap_8 FILLER_49_3311 ();
 sg13g2_decap_8 FILLER_49_3318 ();
 sg13g2_decap_8 FILLER_49_3325 ();
 sg13g2_decap_8 FILLER_49_3332 ();
 sg13g2_decap_8 FILLER_49_3339 ();
 sg13g2_decap_8 FILLER_49_3346 ();
 sg13g2_decap_8 FILLER_49_3353 ();
 sg13g2_decap_8 FILLER_49_3360 ();
 sg13g2_decap_8 FILLER_49_3367 ();
 sg13g2_decap_8 FILLER_49_3374 ();
 sg13g2_decap_8 FILLER_49_3381 ();
 sg13g2_decap_8 FILLER_49_3388 ();
 sg13g2_decap_8 FILLER_49_3395 ();
 sg13g2_decap_8 FILLER_49_3402 ();
 sg13g2_decap_8 FILLER_49_3409 ();
 sg13g2_decap_8 FILLER_49_3416 ();
 sg13g2_decap_8 FILLER_49_3423 ();
 sg13g2_decap_8 FILLER_49_3430 ();
 sg13g2_decap_8 FILLER_49_3437 ();
 sg13g2_decap_8 FILLER_49_3444 ();
 sg13g2_decap_8 FILLER_49_3451 ();
 sg13g2_decap_8 FILLER_49_3458 ();
 sg13g2_decap_8 FILLER_49_3465 ();
 sg13g2_decap_8 FILLER_49_3472 ();
 sg13g2_decap_8 FILLER_49_3479 ();
 sg13g2_decap_8 FILLER_49_3486 ();
 sg13g2_decap_8 FILLER_49_3493 ();
 sg13g2_decap_8 FILLER_49_3500 ();
 sg13g2_decap_8 FILLER_49_3507 ();
 sg13g2_decap_8 FILLER_49_3514 ();
 sg13g2_decap_8 FILLER_49_3521 ();
 sg13g2_decap_8 FILLER_49_3528 ();
 sg13g2_decap_8 FILLER_49_3535 ();
 sg13g2_decap_8 FILLER_49_3542 ();
 sg13g2_decap_8 FILLER_49_3549 ();
 sg13g2_decap_8 FILLER_49_3556 ();
 sg13g2_decap_8 FILLER_49_3563 ();
 sg13g2_decap_8 FILLER_49_3570 ();
 sg13g2_fill_2 FILLER_49_3577 ();
 sg13g2_fill_1 FILLER_49_3579 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_98 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_decap_8 FILLER_50_112 ();
 sg13g2_decap_8 FILLER_50_119 ();
 sg13g2_decap_8 FILLER_50_126 ();
 sg13g2_decap_8 FILLER_50_133 ();
 sg13g2_decap_8 FILLER_50_140 ();
 sg13g2_decap_8 FILLER_50_147 ();
 sg13g2_decap_8 FILLER_50_154 ();
 sg13g2_decap_8 FILLER_50_161 ();
 sg13g2_decap_8 FILLER_50_168 ();
 sg13g2_decap_8 FILLER_50_175 ();
 sg13g2_decap_8 FILLER_50_182 ();
 sg13g2_decap_8 FILLER_50_189 ();
 sg13g2_decap_8 FILLER_50_196 ();
 sg13g2_decap_8 FILLER_50_203 ();
 sg13g2_decap_8 FILLER_50_210 ();
 sg13g2_decap_8 FILLER_50_217 ();
 sg13g2_decap_8 FILLER_50_224 ();
 sg13g2_decap_8 FILLER_50_231 ();
 sg13g2_decap_8 FILLER_50_238 ();
 sg13g2_decap_8 FILLER_50_245 ();
 sg13g2_decap_8 FILLER_50_252 ();
 sg13g2_decap_8 FILLER_50_259 ();
 sg13g2_decap_8 FILLER_50_266 ();
 sg13g2_decap_8 FILLER_50_273 ();
 sg13g2_decap_8 FILLER_50_280 ();
 sg13g2_decap_8 FILLER_50_287 ();
 sg13g2_decap_8 FILLER_50_294 ();
 sg13g2_decap_8 FILLER_50_301 ();
 sg13g2_decap_8 FILLER_50_308 ();
 sg13g2_decap_8 FILLER_50_315 ();
 sg13g2_decap_8 FILLER_50_322 ();
 sg13g2_decap_8 FILLER_50_329 ();
 sg13g2_decap_8 FILLER_50_336 ();
 sg13g2_decap_8 FILLER_50_343 ();
 sg13g2_decap_8 FILLER_50_350 ();
 sg13g2_decap_8 FILLER_50_357 ();
 sg13g2_decap_8 FILLER_50_364 ();
 sg13g2_decap_8 FILLER_50_371 ();
 sg13g2_decap_8 FILLER_50_378 ();
 sg13g2_decap_8 FILLER_50_385 ();
 sg13g2_decap_8 FILLER_50_392 ();
 sg13g2_decap_8 FILLER_50_399 ();
 sg13g2_decap_8 FILLER_50_406 ();
 sg13g2_decap_8 FILLER_50_413 ();
 sg13g2_decap_8 FILLER_50_420 ();
 sg13g2_decap_8 FILLER_50_427 ();
 sg13g2_decap_8 FILLER_50_434 ();
 sg13g2_decap_8 FILLER_50_441 ();
 sg13g2_decap_8 FILLER_50_448 ();
 sg13g2_decap_8 FILLER_50_455 ();
 sg13g2_decap_8 FILLER_50_462 ();
 sg13g2_decap_8 FILLER_50_469 ();
 sg13g2_decap_8 FILLER_50_476 ();
 sg13g2_decap_8 FILLER_50_483 ();
 sg13g2_decap_8 FILLER_50_490 ();
 sg13g2_decap_8 FILLER_50_497 ();
 sg13g2_decap_8 FILLER_50_504 ();
 sg13g2_decap_8 FILLER_50_511 ();
 sg13g2_decap_8 FILLER_50_518 ();
 sg13g2_decap_8 FILLER_50_525 ();
 sg13g2_decap_8 FILLER_50_532 ();
 sg13g2_decap_8 FILLER_50_539 ();
 sg13g2_decap_8 FILLER_50_546 ();
 sg13g2_decap_8 FILLER_50_553 ();
 sg13g2_decap_8 FILLER_50_560 ();
 sg13g2_decap_8 FILLER_50_567 ();
 sg13g2_decap_8 FILLER_50_574 ();
 sg13g2_decap_8 FILLER_50_581 ();
 sg13g2_decap_8 FILLER_50_588 ();
 sg13g2_decap_8 FILLER_50_595 ();
 sg13g2_decap_8 FILLER_50_602 ();
 sg13g2_decap_8 FILLER_50_609 ();
 sg13g2_decap_8 FILLER_50_616 ();
 sg13g2_decap_8 FILLER_50_623 ();
 sg13g2_decap_8 FILLER_50_630 ();
 sg13g2_decap_8 FILLER_50_637 ();
 sg13g2_decap_8 FILLER_50_644 ();
 sg13g2_decap_8 FILLER_50_651 ();
 sg13g2_decap_8 FILLER_50_658 ();
 sg13g2_decap_8 FILLER_50_665 ();
 sg13g2_decap_8 FILLER_50_672 ();
 sg13g2_decap_8 FILLER_50_679 ();
 sg13g2_decap_8 FILLER_50_686 ();
 sg13g2_decap_8 FILLER_50_693 ();
 sg13g2_decap_8 FILLER_50_700 ();
 sg13g2_decap_8 FILLER_50_707 ();
 sg13g2_decap_8 FILLER_50_714 ();
 sg13g2_decap_8 FILLER_50_721 ();
 sg13g2_decap_8 FILLER_50_728 ();
 sg13g2_decap_8 FILLER_50_735 ();
 sg13g2_decap_8 FILLER_50_742 ();
 sg13g2_decap_8 FILLER_50_749 ();
 sg13g2_decap_8 FILLER_50_756 ();
 sg13g2_decap_8 FILLER_50_763 ();
 sg13g2_decap_8 FILLER_50_770 ();
 sg13g2_decap_8 FILLER_50_777 ();
 sg13g2_decap_8 FILLER_50_784 ();
 sg13g2_decap_8 FILLER_50_791 ();
 sg13g2_decap_8 FILLER_50_798 ();
 sg13g2_decap_8 FILLER_50_805 ();
 sg13g2_decap_8 FILLER_50_812 ();
 sg13g2_decap_8 FILLER_50_819 ();
 sg13g2_decap_8 FILLER_50_826 ();
 sg13g2_decap_8 FILLER_50_833 ();
 sg13g2_decap_8 FILLER_50_840 ();
 sg13g2_decap_8 FILLER_50_847 ();
 sg13g2_decap_8 FILLER_50_854 ();
 sg13g2_decap_8 FILLER_50_861 ();
 sg13g2_decap_8 FILLER_50_868 ();
 sg13g2_decap_8 FILLER_50_875 ();
 sg13g2_decap_8 FILLER_50_882 ();
 sg13g2_decap_8 FILLER_50_889 ();
 sg13g2_decap_8 FILLER_50_896 ();
 sg13g2_decap_8 FILLER_50_903 ();
 sg13g2_decap_8 FILLER_50_910 ();
 sg13g2_decap_8 FILLER_50_917 ();
 sg13g2_decap_8 FILLER_50_924 ();
 sg13g2_decap_8 FILLER_50_931 ();
 sg13g2_decap_8 FILLER_50_938 ();
 sg13g2_decap_8 FILLER_50_945 ();
 sg13g2_decap_8 FILLER_50_952 ();
 sg13g2_decap_8 FILLER_50_959 ();
 sg13g2_decap_8 FILLER_50_966 ();
 sg13g2_decap_8 FILLER_50_973 ();
 sg13g2_decap_8 FILLER_50_980 ();
 sg13g2_decap_8 FILLER_50_987 ();
 sg13g2_decap_8 FILLER_50_994 ();
 sg13g2_decap_8 FILLER_50_1001 ();
 sg13g2_decap_8 FILLER_50_1008 ();
 sg13g2_decap_8 FILLER_50_1015 ();
 sg13g2_decap_8 FILLER_50_1022 ();
 sg13g2_decap_8 FILLER_50_1029 ();
 sg13g2_decap_8 FILLER_50_1036 ();
 sg13g2_decap_8 FILLER_50_1043 ();
 sg13g2_decap_8 FILLER_50_1050 ();
 sg13g2_decap_8 FILLER_50_1057 ();
 sg13g2_decap_8 FILLER_50_1064 ();
 sg13g2_decap_8 FILLER_50_1071 ();
 sg13g2_decap_8 FILLER_50_1078 ();
 sg13g2_decap_8 FILLER_50_1085 ();
 sg13g2_decap_8 FILLER_50_1092 ();
 sg13g2_decap_8 FILLER_50_1099 ();
 sg13g2_decap_8 FILLER_50_1106 ();
 sg13g2_decap_8 FILLER_50_1113 ();
 sg13g2_decap_8 FILLER_50_1120 ();
 sg13g2_decap_8 FILLER_50_1127 ();
 sg13g2_decap_8 FILLER_50_1134 ();
 sg13g2_decap_8 FILLER_50_1141 ();
 sg13g2_decap_8 FILLER_50_1148 ();
 sg13g2_decap_8 FILLER_50_1155 ();
 sg13g2_decap_8 FILLER_50_1162 ();
 sg13g2_decap_8 FILLER_50_1169 ();
 sg13g2_decap_8 FILLER_50_1176 ();
 sg13g2_decap_8 FILLER_50_1183 ();
 sg13g2_decap_8 FILLER_50_1190 ();
 sg13g2_decap_8 FILLER_50_1197 ();
 sg13g2_decap_8 FILLER_50_1204 ();
 sg13g2_decap_8 FILLER_50_1211 ();
 sg13g2_decap_8 FILLER_50_1218 ();
 sg13g2_decap_8 FILLER_50_1225 ();
 sg13g2_decap_8 FILLER_50_1232 ();
 sg13g2_decap_8 FILLER_50_1239 ();
 sg13g2_decap_8 FILLER_50_1246 ();
 sg13g2_decap_8 FILLER_50_1253 ();
 sg13g2_decap_8 FILLER_50_1260 ();
 sg13g2_decap_8 FILLER_50_1267 ();
 sg13g2_decap_8 FILLER_50_1274 ();
 sg13g2_decap_8 FILLER_50_1281 ();
 sg13g2_decap_8 FILLER_50_1288 ();
 sg13g2_decap_8 FILLER_50_1295 ();
 sg13g2_decap_8 FILLER_50_1302 ();
 sg13g2_decap_8 FILLER_50_1309 ();
 sg13g2_decap_8 FILLER_50_1316 ();
 sg13g2_decap_8 FILLER_50_1323 ();
 sg13g2_decap_8 FILLER_50_1330 ();
 sg13g2_decap_8 FILLER_50_1337 ();
 sg13g2_decap_8 FILLER_50_1344 ();
 sg13g2_decap_8 FILLER_50_1351 ();
 sg13g2_decap_8 FILLER_50_1358 ();
 sg13g2_decap_8 FILLER_50_1365 ();
 sg13g2_decap_8 FILLER_50_1372 ();
 sg13g2_decap_8 FILLER_50_1379 ();
 sg13g2_decap_8 FILLER_50_1386 ();
 sg13g2_decap_8 FILLER_50_1393 ();
 sg13g2_decap_8 FILLER_50_1400 ();
 sg13g2_decap_8 FILLER_50_1407 ();
 sg13g2_decap_8 FILLER_50_1414 ();
 sg13g2_decap_8 FILLER_50_1421 ();
 sg13g2_decap_8 FILLER_50_1428 ();
 sg13g2_decap_8 FILLER_50_1435 ();
 sg13g2_decap_8 FILLER_50_1442 ();
 sg13g2_decap_8 FILLER_50_1449 ();
 sg13g2_decap_8 FILLER_50_1456 ();
 sg13g2_decap_8 FILLER_50_1463 ();
 sg13g2_decap_8 FILLER_50_1470 ();
 sg13g2_decap_8 FILLER_50_1477 ();
 sg13g2_decap_8 FILLER_50_1484 ();
 sg13g2_decap_8 FILLER_50_1491 ();
 sg13g2_decap_8 FILLER_50_1498 ();
 sg13g2_decap_8 FILLER_50_1505 ();
 sg13g2_decap_8 FILLER_50_1512 ();
 sg13g2_decap_8 FILLER_50_1519 ();
 sg13g2_decap_8 FILLER_50_1526 ();
 sg13g2_decap_8 FILLER_50_1533 ();
 sg13g2_decap_8 FILLER_50_1540 ();
 sg13g2_decap_8 FILLER_50_1547 ();
 sg13g2_decap_8 FILLER_50_1554 ();
 sg13g2_decap_8 FILLER_50_1561 ();
 sg13g2_decap_8 FILLER_50_1568 ();
 sg13g2_decap_8 FILLER_50_1575 ();
 sg13g2_decap_8 FILLER_50_1582 ();
 sg13g2_decap_8 FILLER_50_1589 ();
 sg13g2_decap_8 FILLER_50_1596 ();
 sg13g2_decap_8 FILLER_50_1603 ();
 sg13g2_decap_8 FILLER_50_1610 ();
 sg13g2_decap_8 FILLER_50_1617 ();
 sg13g2_decap_8 FILLER_50_1624 ();
 sg13g2_decap_8 FILLER_50_1631 ();
 sg13g2_decap_8 FILLER_50_1638 ();
 sg13g2_decap_8 FILLER_50_1645 ();
 sg13g2_decap_8 FILLER_50_1652 ();
 sg13g2_decap_8 FILLER_50_1659 ();
 sg13g2_decap_8 FILLER_50_1666 ();
 sg13g2_decap_8 FILLER_50_1673 ();
 sg13g2_decap_8 FILLER_50_1680 ();
 sg13g2_decap_8 FILLER_50_1687 ();
 sg13g2_decap_8 FILLER_50_1694 ();
 sg13g2_decap_8 FILLER_50_1701 ();
 sg13g2_decap_8 FILLER_50_1708 ();
 sg13g2_decap_8 FILLER_50_1715 ();
 sg13g2_decap_8 FILLER_50_1722 ();
 sg13g2_decap_8 FILLER_50_1729 ();
 sg13g2_decap_8 FILLER_50_1736 ();
 sg13g2_decap_8 FILLER_50_1743 ();
 sg13g2_decap_8 FILLER_50_1750 ();
 sg13g2_decap_8 FILLER_50_1757 ();
 sg13g2_decap_8 FILLER_50_1764 ();
 sg13g2_decap_8 FILLER_50_1771 ();
 sg13g2_decap_8 FILLER_50_1778 ();
 sg13g2_decap_8 FILLER_50_1785 ();
 sg13g2_decap_8 FILLER_50_1792 ();
 sg13g2_decap_8 FILLER_50_1799 ();
 sg13g2_decap_8 FILLER_50_1806 ();
 sg13g2_decap_8 FILLER_50_1813 ();
 sg13g2_decap_8 FILLER_50_1820 ();
 sg13g2_decap_8 FILLER_50_1827 ();
 sg13g2_decap_8 FILLER_50_1834 ();
 sg13g2_decap_8 FILLER_50_1841 ();
 sg13g2_decap_8 FILLER_50_1848 ();
 sg13g2_decap_8 FILLER_50_1855 ();
 sg13g2_decap_8 FILLER_50_1862 ();
 sg13g2_decap_8 FILLER_50_1869 ();
 sg13g2_decap_8 FILLER_50_1876 ();
 sg13g2_decap_8 FILLER_50_1883 ();
 sg13g2_decap_8 FILLER_50_1890 ();
 sg13g2_decap_8 FILLER_50_1897 ();
 sg13g2_decap_8 FILLER_50_1904 ();
 sg13g2_decap_8 FILLER_50_1911 ();
 sg13g2_decap_8 FILLER_50_1918 ();
 sg13g2_decap_8 FILLER_50_1925 ();
 sg13g2_decap_8 FILLER_50_1932 ();
 sg13g2_decap_8 FILLER_50_1939 ();
 sg13g2_decap_8 FILLER_50_1946 ();
 sg13g2_decap_8 FILLER_50_1953 ();
 sg13g2_decap_8 FILLER_50_1960 ();
 sg13g2_decap_8 FILLER_50_1967 ();
 sg13g2_decap_8 FILLER_50_1974 ();
 sg13g2_decap_8 FILLER_50_1981 ();
 sg13g2_decap_8 FILLER_50_1988 ();
 sg13g2_decap_8 FILLER_50_1995 ();
 sg13g2_decap_8 FILLER_50_2002 ();
 sg13g2_decap_8 FILLER_50_2009 ();
 sg13g2_decap_8 FILLER_50_2016 ();
 sg13g2_decap_8 FILLER_50_2023 ();
 sg13g2_decap_8 FILLER_50_2030 ();
 sg13g2_decap_8 FILLER_50_2037 ();
 sg13g2_decap_8 FILLER_50_2044 ();
 sg13g2_decap_8 FILLER_50_2051 ();
 sg13g2_decap_8 FILLER_50_2058 ();
 sg13g2_decap_8 FILLER_50_2065 ();
 sg13g2_decap_8 FILLER_50_2072 ();
 sg13g2_decap_8 FILLER_50_2079 ();
 sg13g2_decap_8 FILLER_50_2086 ();
 sg13g2_decap_8 FILLER_50_2093 ();
 sg13g2_decap_8 FILLER_50_2100 ();
 sg13g2_decap_8 FILLER_50_2107 ();
 sg13g2_decap_8 FILLER_50_2114 ();
 sg13g2_decap_8 FILLER_50_2121 ();
 sg13g2_decap_8 FILLER_50_2128 ();
 sg13g2_decap_8 FILLER_50_2135 ();
 sg13g2_decap_8 FILLER_50_2142 ();
 sg13g2_decap_8 FILLER_50_2149 ();
 sg13g2_decap_8 FILLER_50_2156 ();
 sg13g2_decap_8 FILLER_50_2163 ();
 sg13g2_decap_8 FILLER_50_2170 ();
 sg13g2_decap_8 FILLER_50_2177 ();
 sg13g2_decap_8 FILLER_50_2184 ();
 sg13g2_decap_8 FILLER_50_2191 ();
 sg13g2_decap_8 FILLER_50_2198 ();
 sg13g2_decap_8 FILLER_50_2205 ();
 sg13g2_decap_8 FILLER_50_2212 ();
 sg13g2_decap_8 FILLER_50_2219 ();
 sg13g2_decap_8 FILLER_50_2226 ();
 sg13g2_decap_8 FILLER_50_2233 ();
 sg13g2_decap_8 FILLER_50_2240 ();
 sg13g2_decap_8 FILLER_50_2247 ();
 sg13g2_decap_8 FILLER_50_2254 ();
 sg13g2_decap_8 FILLER_50_2261 ();
 sg13g2_decap_8 FILLER_50_2268 ();
 sg13g2_decap_8 FILLER_50_2275 ();
 sg13g2_decap_8 FILLER_50_2282 ();
 sg13g2_decap_8 FILLER_50_2289 ();
 sg13g2_decap_8 FILLER_50_2296 ();
 sg13g2_decap_8 FILLER_50_2303 ();
 sg13g2_decap_8 FILLER_50_2310 ();
 sg13g2_decap_8 FILLER_50_2317 ();
 sg13g2_decap_8 FILLER_50_2324 ();
 sg13g2_decap_8 FILLER_50_2331 ();
 sg13g2_decap_8 FILLER_50_2338 ();
 sg13g2_decap_8 FILLER_50_2345 ();
 sg13g2_decap_8 FILLER_50_2352 ();
 sg13g2_decap_8 FILLER_50_2359 ();
 sg13g2_decap_8 FILLER_50_2366 ();
 sg13g2_decap_8 FILLER_50_2373 ();
 sg13g2_decap_8 FILLER_50_2380 ();
 sg13g2_decap_8 FILLER_50_2387 ();
 sg13g2_decap_8 FILLER_50_2394 ();
 sg13g2_decap_8 FILLER_50_2401 ();
 sg13g2_decap_8 FILLER_50_2408 ();
 sg13g2_decap_8 FILLER_50_2415 ();
 sg13g2_decap_8 FILLER_50_2422 ();
 sg13g2_decap_8 FILLER_50_2429 ();
 sg13g2_decap_8 FILLER_50_2436 ();
 sg13g2_decap_8 FILLER_50_2443 ();
 sg13g2_decap_8 FILLER_50_2450 ();
 sg13g2_decap_8 FILLER_50_2457 ();
 sg13g2_decap_8 FILLER_50_2464 ();
 sg13g2_decap_8 FILLER_50_2471 ();
 sg13g2_decap_8 FILLER_50_2478 ();
 sg13g2_decap_8 FILLER_50_2485 ();
 sg13g2_decap_8 FILLER_50_2492 ();
 sg13g2_decap_8 FILLER_50_2499 ();
 sg13g2_decap_8 FILLER_50_2506 ();
 sg13g2_decap_8 FILLER_50_2513 ();
 sg13g2_decap_8 FILLER_50_2520 ();
 sg13g2_decap_8 FILLER_50_2527 ();
 sg13g2_decap_8 FILLER_50_2534 ();
 sg13g2_decap_8 FILLER_50_2541 ();
 sg13g2_decap_8 FILLER_50_2548 ();
 sg13g2_decap_8 FILLER_50_2555 ();
 sg13g2_decap_8 FILLER_50_2562 ();
 sg13g2_decap_8 FILLER_50_2569 ();
 sg13g2_decap_8 FILLER_50_2576 ();
 sg13g2_decap_8 FILLER_50_2583 ();
 sg13g2_decap_8 FILLER_50_2590 ();
 sg13g2_decap_8 FILLER_50_2597 ();
 sg13g2_decap_8 FILLER_50_2604 ();
 sg13g2_decap_8 FILLER_50_2611 ();
 sg13g2_decap_8 FILLER_50_2618 ();
 sg13g2_decap_8 FILLER_50_2625 ();
 sg13g2_decap_8 FILLER_50_2632 ();
 sg13g2_decap_8 FILLER_50_2639 ();
 sg13g2_decap_8 FILLER_50_2646 ();
 sg13g2_decap_8 FILLER_50_2653 ();
 sg13g2_decap_8 FILLER_50_2660 ();
 sg13g2_decap_8 FILLER_50_2667 ();
 sg13g2_decap_8 FILLER_50_2674 ();
 sg13g2_decap_8 FILLER_50_2681 ();
 sg13g2_decap_8 FILLER_50_2688 ();
 sg13g2_decap_8 FILLER_50_2695 ();
 sg13g2_decap_8 FILLER_50_2702 ();
 sg13g2_decap_8 FILLER_50_2709 ();
 sg13g2_decap_8 FILLER_50_2716 ();
 sg13g2_decap_8 FILLER_50_2723 ();
 sg13g2_decap_8 FILLER_50_2730 ();
 sg13g2_decap_8 FILLER_50_2737 ();
 sg13g2_decap_8 FILLER_50_2744 ();
 sg13g2_decap_8 FILLER_50_2751 ();
 sg13g2_decap_8 FILLER_50_2758 ();
 sg13g2_decap_8 FILLER_50_2765 ();
 sg13g2_decap_8 FILLER_50_2772 ();
 sg13g2_decap_8 FILLER_50_2779 ();
 sg13g2_decap_8 FILLER_50_2786 ();
 sg13g2_decap_8 FILLER_50_2793 ();
 sg13g2_decap_8 FILLER_50_2800 ();
 sg13g2_decap_8 FILLER_50_2807 ();
 sg13g2_decap_8 FILLER_50_2814 ();
 sg13g2_decap_8 FILLER_50_2821 ();
 sg13g2_decap_8 FILLER_50_2828 ();
 sg13g2_decap_8 FILLER_50_2835 ();
 sg13g2_decap_8 FILLER_50_2842 ();
 sg13g2_decap_8 FILLER_50_2849 ();
 sg13g2_decap_8 FILLER_50_2856 ();
 sg13g2_decap_8 FILLER_50_2863 ();
 sg13g2_decap_8 FILLER_50_2870 ();
 sg13g2_decap_8 FILLER_50_2877 ();
 sg13g2_decap_8 FILLER_50_2884 ();
 sg13g2_decap_8 FILLER_50_2891 ();
 sg13g2_decap_8 FILLER_50_2898 ();
 sg13g2_decap_8 FILLER_50_2905 ();
 sg13g2_decap_8 FILLER_50_2912 ();
 sg13g2_decap_8 FILLER_50_2919 ();
 sg13g2_decap_8 FILLER_50_2926 ();
 sg13g2_decap_8 FILLER_50_2933 ();
 sg13g2_decap_8 FILLER_50_2940 ();
 sg13g2_decap_8 FILLER_50_2947 ();
 sg13g2_decap_8 FILLER_50_2954 ();
 sg13g2_decap_8 FILLER_50_2961 ();
 sg13g2_decap_8 FILLER_50_2968 ();
 sg13g2_decap_8 FILLER_50_2975 ();
 sg13g2_decap_8 FILLER_50_2982 ();
 sg13g2_decap_8 FILLER_50_2989 ();
 sg13g2_decap_8 FILLER_50_2996 ();
 sg13g2_decap_8 FILLER_50_3003 ();
 sg13g2_decap_8 FILLER_50_3010 ();
 sg13g2_decap_8 FILLER_50_3017 ();
 sg13g2_decap_8 FILLER_50_3024 ();
 sg13g2_decap_8 FILLER_50_3031 ();
 sg13g2_decap_8 FILLER_50_3038 ();
 sg13g2_decap_8 FILLER_50_3045 ();
 sg13g2_decap_8 FILLER_50_3052 ();
 sg13g2_decap_8 FILLER_50_3059 ();
 sg13g2_decap_8 FILLER_50_3066 ();
 sg13g2_decap_8 FILLER_50_3073 ();
 sg13g2_decap_8 FILLER_50_3080 ();
 sg13g2_decap_8 FILLER_50_3087 ();
 sg13g2_decap_8 FILLER_50_3094 ();
 sg13g2_decap_8 FILLER_50_3101 ();
 sg13g2_decap_8 FILLER_50_3108 ();
 sg13g2_decap_8 FILLER_50_3115 ();
 sg13g2_decap_8 FILLER_50_3122 ();
 sg13g2_decap_8 FILLER_50_3129 ();
 sg13g2_decap_8 FILLER_50_3136 ();
 sg13g2_decap_8 FILLER_50_3143 ();
 sg13g2_decap_8 FILLER_50_3150 ();
 sg13g2_decap_8 FILLER_50_3157 ();
 sg13g2_decap_8 FILLER_50_3164 ();
 sg13g2_decap_8 FILLER_50_3171 ();
 sg13g2_decap_8 FILLER_50_3178 ();
 sg13g2_decap_8 FILLER_50_3185 ();
 sg13g2_decap_8 FILLER_50_3192 ();
 sg13g2_decap_8 FILLER_50_3199 ();
 sg13g2_decap_8 FILLER_50_3206 ();
 sg13g2_decap_8 FILLER_50_3213 ();
 sg13g2_decap_8 FILLER_50_3220 ();
 sg13g2_decap_8 FILLER_50_3227 ();
 sg13g2_decap_8 FILLER_50_3234 ();
 sg13g2_decap_8 FILLER_50_3241 ();
 sg13g2_decap_8 FILLER_50_3248 ();
 sg13g2_decap_8 FILLER_50_3255 ();
 sg13g2_decap_8 FILLER_50_3262 ();
 sg13g2_decap_8 FILLER_50_3269 ();
 sg13g2_decap_8 FILLER_50_3276 ();
 sg13g2_decap_8 FILLER_50_3283 ();
 sg13g2_decap_8 FILLER_50_3290 ();
 sg13g2_decap_8 FILLER_50_3297 ();
 sg13g2_decap_8 FILLER_50_3304 ();
 sg13g2_decap_8 FILLER_50_3311 ();
 sg13g2_decap_8 FILLER_50_3318 ();
 sg13g2_decap_8 FILLER_50_3325 ();
 sg13g2_decap_8 FILLER_50_3332 ();
 sg13g2_decap_8 FILLER_50_3339 ();
 sg13g2_decap_8 FILLER_50_3346 ();
 sg13g2_decap_8 FILLER_50_3353 ();
 sg13g2_decap_8 FILLER_50_3360 ();
 sg13g2_decap_8 FILLER_50_3367 ();
 sg13g2_decap_8 FILLER_50_3374 ();
 sg13g2_decap_8 FILLER_50_3381 ();
 sg13g2_decap_8 FILLER_50_3388 ();
 sg13g2_decap_8 FILLER_50_3395 ();
 sg13g2_decap_8 FILLER_50_3402 ();
 sg13g2_decap_8 FILLER_50_3409 ();
 sg13g2_decap_8 FILLER_50_3416 ();
 sg13g2_decap_8 FILLER_50_3423 ();
 sg13g2_decap_8 FILLER_50_3430 ();
 sg13g2_decap_8 FILLER_50_3437 ();
 sg13g2_decap_8 FILLER_50_3444 ();
 sg13g2_decap_8 FILLER_50_3451 ();
 sg13g2_decap_8 FILLER_50_3458 ();
 sg13g2_decap_8 FILLER_50_3465 ();
 sg13g2_decap_8 FILLER_50_3472 ();
 sg13g2_decap_8 FILLER_50_3479 ();
 sg13g2_decap_8 FILLER_50_3486 ();
 sg13g2_decap_8 FILLER_50_3493 ();
 sg13g2_decap_8 FILLER_50_3500 ();
 sg13g2_decap_8 FILLER_50_3507 ();
 sg13g2_decap_8 FILLER_50_3514 ();
 sg13g2_decap_8 FILLER_50_3521 ();
 sg13g2_decap_8 FILLER_50_3528 ();
 sg13g2_decap_8 FILLER_50_3535 ();
 sg13g2_decap_8 FILLER_50_3542 ();
 sg13g2_decap_8 FILLER_50_3549 ();
 sg13g2_decap_8 FILLER_50_3556 ();
 sg13g2_decap_8 FILLER_50_3563 ();
 sg13g2_decap_8 FILLER_50_3570 ();
 sg13g2_fill_2 FILLER_50_3577 ();
 sg13g2_fill_1 FILLER_50_3579 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_98 ();
 sg13g2_decap_8 FILLER_51_105 ();
 sg13g2_decap_8 FILLER_51_112 ();
 sg13g2_decap_8 FILLER_51_119 ();
 sg13g2_decap_8 FILLER_51_126 ();
 sg13g2_decap_8 FILLER_51_133 ();
 sg13g2_decap_8 FILLER_51_140 ();
 sg13g2_decap_8 FILLER_51_147 ();
 sg13g2_decap_8 FILLER_51_154 ();
 sg13g2_decap_8 FILLER_51_161 ();
 sg13g2_decap_8 FILLER_51_168 ();
 sg13g2_decap_8 FILLER_51_175 ();
 sg13g2_decap_8 FILLER_51_182 ();
 sg13g2_decap_8 FILLER_51_189 ();
 sg13g2_decap_8 FILLER_51_196 ();
 sg13g2_decap_8 FILLER_51_203 ();
 sg13g2_decap_8 FILLER_51_210 ();
 sg13g2_decap_8 FILLER_51_217 ();
 sg13g2_decap_8 FILLER_51_224 ();
 sg13g2_decap_8 FILLER_51_231 ();
 sg13g2_decap_8 FILLER_51_238 ();
 sg13g2_decap_8 FILLER_51_245 ();
 sg13g2_decap_8 FILLER_51_252 ();
 sg13g2_decap_8 FILLER_51_259 ();
 sg13g2_decap_8 FILLER_51_266 ();
 sg13g2_decap_8 FILLER_51_273 ();
 sg13g2_decap_8 FILLER_51_280 ();
 sg13g2_decap_8 FILLER_51_287 ();
 sg13g2_decap_8 FILLER_51_294 ();
 sg13g2_decap_8 FILLER_51_301 ();
 sg13g2_decap_8 FILLER_51_308 ();
 sg13g2_decap_8 FILLER_51_315 ();
 sg13g2_decap_8 FILLER_51_322 ();
 sg13g2_decap_8 FILLER_51_329 ();
 sg13g2_decap_8 FILLER_51_336 ();
 sg13g2_decap_8 FILLER_51_343 ();
 sg13g2_decap_8 FILLER_51_350 ();
 sg13g2_decap_8 FILLER_51_357 ();
 sg13g2_decap_8 FILLER_51_364 ();
 sg13g2_decap_8 FILLER_51_371 ();
 sg13g2_decap_8 FILLER_51_378 ();
 sg13g2_decap_8 FILLER_51_385 ();
 sg13g2_decap_8 FILLER_51_392 ();
 sg13g2_decap_8 FILLER_51_399 ();
 sg13g2_decap_8 FILLER_51_406 ();
 sg13g2_decap_8 FILLER_51_413 ();
 sg13g2_decap_8 FILLER_51_420 ();
 sg13g2_decap_8 FILLER_51_427 ();
 sg13g2_decap_8 FILLER_51_434 ();
 sg13g2_decap_8 FILLER_51_441 ();
 sg13g2_decap_8 FILLER_51_448 ();
 sg13g2_decap_8 FILLER_51_455 ();
 sg13g2_decap_8 FILLER_51_462 ();
 sg13g2_decap_8 FILLER_51_469 ();
 sg13g2_decap_8 FILLER_51_476 ();
 sg13g2_decap_8 FILLER_51_483 ();
 sg13g2_decap_8 FILLER_51_490 ();
 sg13g2_decap_8 FILLER_51_497 ();
 sg13g2_decap_8 FILLER_51_504 ();
 sg13g2_decap_8 FILLER_51_511 ();
 sg13g2_decap_8 FILLER_51_518 ();
 sg13g2_decap_8 FILLER_51_525 ();
 sg13g2_decap_8 FILLER_51_532 ();
 sg13g2_decap_8 FILLER_51_539 ();
 sg13g2_decap_8 FILLER_51_546 ();
 sg13g2_decap_8 FILLER_51_553 ();
 sg13g2_decap_8 FILLER_51_560 ();
 sg13g2_decap_8 FILLER_51_567 ();
 sg13g2_decap_8 FILLER_51_574 ();
 sg13g2_decap_8 FILLER_51_581 ();
 sg13g2_decap_8 FILLER_51_588 ();
 sg13g2_decap_8 FILLER_51_595 ();
 sg13g2_decap_8 FILLER_51_602 ();
 sg13g2_decap_8 FILLER_51_609 ();
 sg13g2_decap_8 FILLER_51_616 ();
 sg13g2_decap_8 FILLER_51_623 ();
 sg13g2_decap_8 FILLER_51_630 ();
 sg13g2_decap_8 FILLER_51_637 ();
 sg13g2_decap_8 FILLER_51_644 ();
 sg13g2_decap_8 FILLER_51_651 ();
 sg13g2_decap_8 FILLER_51_658 ();
 sg13g2_decap_8 FILLER_51_665 ();
 sg13g2_decap_8 FILLER_51_672 ();
 sg13g2_decap_8 FILLER_51_679 ();
 sg13g2_decap_8 FILLER_51_686 ();
 sg13g2_decap_8 FILLER_51_693 ();
 sg13g2_decap_8 FILLER_51_700 ();
 sg13g2_decap_8 FILLER_51_707 ();
 sg13g2_decap_8 FILLER_51_714 ();
 sg13g2_decap_8 FILLER_51_721 ();
 sg13g2_decap_8 FILLER_51_728 ();
 sg13g2_decap_8 FILLER_51_735 ();
 sg13g2_decap_8 FILLER_51_742 ();
 sg13g2_decap_8 FILLER_51_749 ();
 sg13g2_decap_8 FILLER_51_756 ();
 sg13g2_decap_8 FILLER_51_763 ();
 sg13g2_decap_8 FILLER_51_770 ();
 sg13g2_decap_8 FILLER_51_777 ();
 sg13g2_decap_8 FILLER_51_784 ();
 sg13g2_decap_8 FILLER_51_791 ();
 sg13g2_decap_8 FILLER_51_798 ();
 sg13g2_decap_8 FILLER_51_805 ();
 sg13g2_decap_8 FILLER_51_812 ();
 sg13g2_decap_8 FILLER_51_819 ();
 sg13g2_decap_8 FILLER_51_826 ();
 sg13g2_decap_8 FILLER_51_833 ();
 sg13g2_decap_8 FILLER_51_840 ();
 sg13g2_decap_8 FILLER_51_847 ();
 sg13g2_decap_8 FILLER_51_854 ();
 sg13g2_decap_8 FILLER_51_861 ();
 sg13g2_decap_8 FILLER_51_868 ();
 sg13g2_decap_8 FILLER_51_875 ();
 sg13g2_decap_8 FILLER_51_882 ();
 sg13g2_decap_8 FILLER_51_889 ();
 sg13g2_decap_8 FILLER_51_896 ();
 sg13g2_decap_8 FILLER_51_903 ();
 sg13g2_decap_8 FILLER_51_910 ();
 sg13g2_decap_8 FILLER_51_917 ();
 sg13g2_decap_8 FILLER_51_924 ();
 sg13g2_decap_8 FILLER_51_931 ();
 sg13g2_decap_8 FILLER_51_938 ();
 sg13g2_decap_8 FILLER_51_945 ();
 sg13g2_decap_8 FILLER_51_952 ();
 sg13g2_decap_8 FILLER_51_959 ();
 sg13g2_decap_8 FILLER_51_966 ();
 sg13g2_decap_8 FILLER_51_973 ();
 sg13g2_decap_8 FILLER_51_980 ();
 sg13g2_decap_8 FILLER_51_987 ();
 sg13g2_decap_8 FILLER_51_994 ();
 sg13g2_decap_8 FILLER_51_1001 ();
 sg13g2_decap_8 FILLER_51_1008 ();
 sg13g2_decap_8 FILLER_51_1015 ();
 sg13g2_decap_8 FILLER_51_1022 ();
 sg13g2_decap_8 FILLER_51_1029 ();
 sg13g2_decap_8 FILLER_51_1036 ();
 sg13g2_decap_8 FILLER_51_1043 ();
 sg13g2_decap_8 FILLER_51_1050 ();
 sg13g2_decap_8 FILLER_51_1057 ();
 sg13g2_decap_8 FILLER_51_1064 ();
 sg13g2_decap_8 FILLER_51_1071 ();
 sg13g2_decap_8 FILLER_51_1078 ();
 sg13g2_decap_8 FILLER_51_1085 ();
 sg13g2_decap_8 FILLER_51_1092 ();
 sg13g2_decap_8 FILLER_51_1099 ();
 sg13g2_decap_8 FILLER_51_1106 ();
 sg13g2_decap_8 FILLER_51_1113 ();
 sg13g2_decap_8 FILLER_51_1120 ();
 sg13g2_decap_8 FILLER_51_1127 ();
 sg13g2_decap_8 FILLER_51_1134 ();
 sg13g2_decap_8 FILLER_51_1141 ();
 sg13g2_decap_8 FILLER_51_1148 ();
 sg13g2_decap_8 FILLER_51_1155 ();
 sg13g2_decap_8 FILLER_51_1162 ();
 sg13g2_decap_8 FILLER_51_1169 ();
 sg13g2_decap_8 FILLER_51_1176 ();
 sg13g2_decap_8 FILLER_51_1183 ();
 sg13g2_decap_8 FILLER_51_1190 ();
 sg13g2_decap_8 FILLER_51_1197 ();
 sg13g2_decap_8 FILLER_51_1204 ();
 sg13g2_decap_8 FILLER_51_1211 ();
 sg13g2_decap_8 FILLER_51_1218 ();
 sg13g2_decap_8 FILLER_51_1225 ();
 sg13g2_decap_8 FILLER_51_1232 ();
 sg13g2_decap_8 FILLER_51_1239 ();
 sg13g2_decap_8 FILLER_51_1246 ();
 sg13g2_decap_8 FILLER_51_1253 ();
 sg13g2_decap_8 FILLER_51_1260 ();
 sg13g2_decap_8 FILLER_51_1267 ();
 sg13g2_decap_8 FILLER_51_1274 ();
 sg13g2_decap_8 FILLER_51_1281 ();
 sg13g2_decap_8 FILLER_51_1288 ();
 sg13g2_decap_8 FILLER_51_1295 ();
 sg13g2_decap_8 FILLER_51_1302 ();
 sg13g2_decap_8 FILLER_51_1309 ();
 sg13g2_decap_8 FILLER_51_1316 ();
 sg13g2_decap_8 FILLER_51_1323 ();
 sg13g2_decap_8 FILLER_51_1330 ();
 sg13g2_decap_8 FILLER_51_1337 ();
 sg13g2_decap_8 FILLER_51_1344 ();
 sg13g2_decap_8 FILLER_51_1351 ();
 sg13g2_decap_8 FILLER_51_1358 ();
 sg13g2_decap_8 FILLER_51_1365 ();
 sg13g2_decap_8 FILLER_51_1372 ();
 sg13g2_decap_8 FILLER_51_1379 ();
 sg13g2_decap_8 FILLER_51_1386 ();
 sg13g2_decap_8 FILLER_51_1393 ();
 sg13g2_decap_8 FILLER_51_1400 ();
 sg13g2_decap_8 FILLER_51_1407 ();
 sg13g2_decap_8 FILLER_51_1414 ();
 sg13g2_decap_8 FILLER_51_1421 ();
 sg13g2_decap_8 FILLER_51_1428 ();
 sg13g2_decap_8 FILLER_51_1435 ();
 sg13g2_decap_8 FILLER_51_1442 ();
 sg13g2_decap_8 FILLER_51_1449 ();
 sg13g2_decap_8 FILLER_51_1456 ();
 sg13g2_decap_8 FILLER_51_1463 ();
 sg13g2_decap_8 FILLER_51_1470 ();
 sg13g2_decap_8 FILLER_51_1477 ();
 sg13g2_decap_8 FILLER_51_1484 ();
 sg13g2_decap_8 FILLER_51_1491 ();
 sg13g2_decap_8 FILLER_51_1498 ();
 sg13g2_decap_8 FILLER_51_1505 ();
 sg13g2_decap_8 FILLER_51_1512 ();
 sg13g2_decap_8 FILLER_51_1519 ();
 sg13g2_decap_8 FILLER_51_1526 ();
 sg13g2_decap_8 FILLER_51_1533 ();
 sg13g2_decap_8 FILLER_51_1540 ();
 sg13g2_decap_8 FILLER_51_1547 ();
 sg13g2_decap_8 FILLER_51_1554 ();
 sg13g2_decap_8 FILLER_51_1561 ();
 sg13g2_decap_8 FILLER_51_1568 ();
 sg13g2_decap_8 FILLER_51_1575 ();
 sg13g2_decap_8 FILLER_51_1582 ();
 sg13g2_decap_8 FILLER_51_1589 ();
 sg13g2_decap_8 FILLER_51_1596 ();
 sg13g2_decap_8 FILLER_51_1603 ();
 sg13g2_decap_8 FILLER_51_1610 ();
 sg13g2_decap_8 FILLER_51_1617 ();
 sg13g2_decap_8 FILLER_51_1624 ();
 sg13g2_decap_8 FILLER_51_1631 ();
 sg13g2_decap_8 FILLER_51_1638 ();
 sg13g2_decap_8 FILLER_51_1645 ();
 sg13g2_decap_8 FILLER_51_1652 ();
 sg13g2_decap_8 FILLER_51_1659 ();
 sg13g2_decap_8 FILLER_51_1666 ();
 sg13g2_decap_8 FILLER_51_1673 ();
 sg13g2_decap_8 FILLER_51_1680 ();
 sg13g2_decap_8 FILLER_51_1687 ();
 sg13g2_decap_8 FILLER_51_1694 ();
 sg13g2_decap_8 FILLER_51_1701 ();
 sg13g2_decap_8 FILLER_51_1708 ();
 sg13g2_decap_8 FILLER_51_1715 ();
 sg13g2_decap_8 FILLER_51_1722 ();
 sg13g2_decap_8 FILLER_51_1729 ();
 sg13g2_decap_8 FILLER_51_1736 ();
 sg13g2_decap_8 FILLER_51_1743 ();
 sg13g2_decap_8 FILLER_51_1750 ();
 sg13g2_decap_8 FILLER_51_1757 ();
 sg13g2_decap_8 FILLER_51_1764 ();
 sg13g2_decap_8 FILLER_51_1771 ();
 sg13g2_decap_8 FILLER_51_1778 ();
 sg13g2_decap_8 FILLER_51_1785 ();
 sg13g2_decap_8 FILLER_51_1792 ();
 sg13g2_decap_8 FILLER_51_1799 ();
 sg13g2_decap_8 FILLER_51_1806 ();
 sg13g2_decap_8 FILLER_51_1813 ();
 sg13g2_decap_8 FILLER_51_1820 ();
 sg13g2_decap_8 FILLER_51_1827 ();
 sg13g2_decap_8 FILLER_51_1834 ();
 sg13g2_decap_8 FILLER_51_1841 ();
 sg13g2_decap_8 FILLER_51_1848 ();
 sg13g2_decap_8 FILLER_51_1855 ();
 sg13g2_decap_8 FILLER_51_1862 ();
 sg13g2_decap_8 FILLER_51_1869 ();
 sg13g2_decap_8 FILLER_51_1876 ();
 sg13g2_decap_8 FILLER_51_1883 ();
 sg13g2_decap_8 FILLER_51_1890 ();
 sg13g2_decap_8 FILLER_51_1897 ();
 sg13g2_decap_8 FILLER_51_1904 ();
 sg13g2_decap_8 FILLER_51_1911 ();
 sg13g2_decap_8 FILLER_51_1918 ();
 sg13g2_decap_8 FILLER_51_1925 ();
 sg13g2_decap_8 FILLER_51_1932 ();
 sg13g2_decap_8 FILLER_51_1939 ();
 sg13g2_decap_8 FILLER_51_1946 ();
 sg13g2_decap_8 FILLER_51_1953 ();
 sg13g2_decap_8 FILLER_51_1960 ();
 sg13g2_decap_8 FILLER_51_1967 ();
 sg13g2_decap_8 FILLER_51_1974 ();
 sg13g2_decap_8 FILLER_51_1981 ();
 sg13g2_decap_8 FILLER_51_1988 ();
 sg13g2_decap_8 FILLER_51_1995 ();
 sg13g2_decap_8 FILLER_51_2002 ();
 sg13g2_decap_8 FILLER_51_2009 ();
 sg13g2_decap_8 FILLER_51_2016 ();
 sg13g2_decap_8 FILLER_51_2023 ();
 sg13g2_decap_8 FILLER_51_2030 ();
 sg13g2_decap_8 FILLER_51_2037 ();
 sg13g2_decap_8 FILLER_51_2044 ();
 sg13g2_decap_8 FILLER_51_2051 ();
 sg13g2_decap_8 FILLER_51_2058 ();
 sg13g2_decap_8 FILLER_51_2065 ();
 sg13g2_decap_8 FILLER_51_2072 ();
 sg13g2_decap_8 FILLER_51_2079 ();
 sg13g2_decap_8 FILLER_51_2086 ();
 sg13g2_decap_8 FILLER_51_2093 ();
 sg13g2_decap_8 FILLER_51_2100 ();
 sg13g2_decap_8 FILLER_51_2107 ();
 sg13g2_decap_8 FILLER_51_2114 ();
 sg13g2_decap_8 FILLER_51_2121 ();
 sg13g2_decap_8 FILLER_51_2128 ();
 sg13g2_decap_8 FILLER_51_2135 ();
 sg13g2_decap_8 FILLER_51_2142 ();
 sg13g2_decap_8 FILLER_51_2149 ();
 sg13g2_decap_8 FILLER_51_2156 ();
 sg13g2_decap_8 FILLER_51_2163 ();
 sg13g2_decap_8 FILLER_51_2170 ();
 sg13g2_decap_8 FILLER_51_2177 ();
 sg13g2_decap_8 FILLER_51_2184 ();
 sg13g2_decap_8 FILLER_51_2191 ();
 sg13g2_decap_8 FILLER_51_2198 ();
 sg13g2_decap_8 FILLER_51_2205 ();
 sg13g2_decap_8 FILLER_51_2212 ();
 sg13g2_decap_8 FILLER_51_2219 ();
 sg13g2_decap_8 FILLER_51_2226 ();
 sg13g2_decap_8 FILLER_51_2233 ();
 sg13g2_decap_8 FILLER_51_2240 ();
 sg13g2_decap_8 FILLER_51_2247 ();
 sg13g2_decap_8 FILLER_51_2254 ();
 sg13g2_decap_8 FILLER_51_2261 ();
 sg13g2_decap_8 FILLER_51_2268 ();
 sg13g2_decap_8 FILLER_51_2275 ();
 sg13g2_decap_8 FILLER_51_2282 ();
 sg13g2_decap_8 FILLER_51_2289 ();
 sg13g2_decap_8 FILLER_51_2296 ();
 sg13g2_decap_8 FILLER_51_2303 ();
 sg13g2_decap_8 FILLER_51_2310 ();
 sg13g2_decap_8 FILLER_51_2317 ();
 sg13g2_decap_8 FILLER_51_2324 ();
 sg13g2_decap_8 FILLER_51_2331 ();
 sg13g2_decap_8 FILLER_51_2338 ();
 sg13g2_decap_8 FILLER_51_2345 ();
 sg13g2_decap_8 FILLER_51_2352 ();
 sg13g2_decap_8 FILLER_51_2359 ();
 sg13g2_decap_8 FILLER_51_2366 ();
 sg13g2_decap_8 FILLER_51_2373 ();
 sg13g2_decap_8 FILLER_51_2380 ();
 sg13g2_decap_8 FILLER_51_2387 ();
 sg13g2_decap_8 FILLER_51_2394 ();
 sg13g2_decap_8 FILLER_51_2401 ();
 sg13g2_decap_8 FILLER_51_2408 ();
 sg13g2_decap_8 FILLER_51_2415 ();
 sg13g2_decap_8 FILLER_51_2422 ();
 sg13g2_decap_8 FILLER_51_2429 ();
 sg13g2_decap_8 FILLER_51_2436 ();
 sg13g2_decap_8 FILLER_51_2443 ();
 sg13g2_decap_8 FILLER_51_2450 ();
 sg13g2_decap_8 FILLER_51_2457 ();
 sg13g2_decap_8 FILLER_51_2464 ();
 sg13g2_decap_8 FILLER_51_2471 ();
 sg13g2_decap_8 FILLER_51_2478 ();
 sg13g2_decap_8 FILLER_51_2485 ();
 sg13g2_decap_8 FILLER_51_2492 ();
 sg13g2_decap_8 FILLER_51_2499 ();
 sg13g2_decap_8 FILLER_51_2506 ();
 sg13g2_decap_8 FILLER_51_2513 ();
 sg13g2_decap_8 FILLER_51_2520 ();
 sg13g2_decap_8 FILLER_51_2527 ();
 sg13g2_decap_8 FILLER_51_2534 ();
 sg13g2_decap_8 FILLER_51_2541 ();
 sg13g2_decap_8 FILLER_51_2548 ();
 sg13g2_decap_8 FILLER_51_2555 ();
 sg13g2_decap_8 FILLER_51_2562 ();
 sg13g2_decap_8 FILLER_51_2569 ();
 sg13g2_decap_8 FILLER_51_2576 ();
 sg13g2_decap_8 FILLER_51_2583 ();
 sg13g2_decap_8 FILLER_51_2590 ();
 sg13g2_decap_8 FILLER_51_2597 ();
 sg13g2_decap_8 FILLER_51_2604 ();
 sg13g2_decap_8 FILLER_51_2611 ();
 sg13g2_decap_8 FILLER_51_2618 ();
 sg13g2_decap_8 FILLER_51_2625 ();
 sg13g2_decap_8 FILLER_51_2632 ();
 sg13g2_decap_8 FILLER_51_2639 ();
 sg13g2_decap_8 FILLER_51_2646 ();
 sg13g2_decap_8 FILLER_51_2653 ();
 sg13g2_decap_8 FILLER_51_2660 ();
 sg13g2_decap_8 FILLER_51_2667 ();
 sg13g2_decap_8 FILLER_51_2674 ();
 sg13g2_decap_8 FILLER_51_2681 ();
 sg13g2_decap_8 FILLER_51_2688 ();
 sg13g2_decap_8 FILLER_51_2695 ();
 sg13g2_decap_8 FILLER_51_2702 ();
 sg13g2_decap_8 FILLER_51_2709 ();
 sg13g2_decap_8 FILLER_51_2716 ();
 sg13g2_decap_8 FILLER_51_2723 ();
 sg13g2_decap_8 FILLER_51_2730 ();
 sg13g2_decap_8 FILLER_51_2737 ();
 sg13g2_decap_8 FILLER_51_2744 ();
 sg13g2_decap_8 FILLER_51_2751 ();
 sg13g2_decap_8 FILLER_51_2758 ();
 sg13g2_decap_8 FILLER_51_2765 ();
 sg13g2_decap_8 FILLER_51_2772 ();
 sg13g2_decap_8 FILLER_51_2779 ();
 sg13g2_decap_8 FILLER_51_2786 ();
 sg13g2_decap_8 FILLER_51_2793 ();
 sg13g2_decap_8 FILLER_51_2800 ();
 sg13g2_decap_8 FILLER_51_2807 ();
 sg13g2_decap_8 FILLER_51_2814 ();
 sg13g2_decap_8 FILLER_51_2821 ();
 sg13g2_decap_8 FILLER_51_2828 ();
 sg13g2_decap_8 FILLER_51_2835 ();
 sg13g2_decap_8 FILLER_51_2842 ();
 sg13g2_decap_8 FILLER_51_2849 ();
 sg13g2_decap_8 FILLER_51_2856 ();
 sg13g2_decap_8 FILLER_51_2863 ();
 sg13g2_decap_8 FILLER_51_2870 ();
 sg13g2_decap_8 FILLER_51_2877 ();
 sg13g2_decap_8 FILLER_51_2884 ();
 sg13g2_decap_8 FILLER_51_2891 ();
 sg13g2_decap_8 FILLER_51_2898 ();
 sg13g2_decap_8 FILLER_51_2905 ();
 sg13g2_decap_8 FILLER_51_2912 ();
 sg13g2_decap_8 FILLER_51_2919 ();
 sg13g2_decap_8 FILLER_51_2926 ();
 sg13g2_decap_8 FILLER_51_2933 ();
 sg13g2_decap_8 FILLER_51_2940 ();
 sg13g2_decap_8 FILLER_51_2947 ();
 sg13g2_decap_8 FILLER_51_2954 ();
 sg13g2_decap_8 FILLER_51_2961 ();
 sg13g2_decap_8 FILLER_51_2968 ();
 sg13g2_decap_8 FILLER_51_2975 ();
 sg13g2_decap_8 FILLER_51_2982 ();
 sg13g2_decap_8 FILLER_51_2989 ();
 sg13g2_decap_8 FILLER_51_2996 ();
 sg13g2_decap_8 FILLER_51_3003 ();
 sg13g2_decap_8 FILLER_51_3010 ();
 sg13g2_decap_8 FILLER_51_3017 ();
 sg13g2_decap_8 FILLER_51_3024 ();
 sg13g2_decap_8 FILLER_51_3031 ();
 sg13g2_decap_8 FILLER_51_3038 ();
 sg13g2_decap_8 FILLER_51_3045 ();
 sg13g2_decap_8 FILLER_51_3052 ();
 sg13g2_decap_8 FILLER_51_3059 ();
 sg13g2_decap_8 FILLER_51_3066 ();
 sg13g2_decap_8 FILLER_51_3073 ();
 sg13g2_decap_8 FILLER_51_3080 ();
 sg13g2_decap_8 FILLER_51_3087 ();
 sg13g2_decap_8 FILLER_51_3094 ();
 sg13g2_decap_8 FILLER_51_3101 ();
 sg13g2_decap_8 FILLER_51_3108 ();
 sg13g2_decap_8 FILLER_51_3115 ();
 sg13g2_decap_8 FILLER_51_3122 ();
 sg13g2_decap_8 FILLER_51_3129 ();
 sg13g2_decap_8 FILLER_51_3136 ();
 sg13g2_decap_8 FILLER_51_3143 ();
 sg13g2_decap_8 FILLER_51_3150 ();
 sg13g2_decap_8 FILLER_51_3157 ();
 sg13g2_decap_8 FILLER_51_3164 ();
 sg13g2_decap_8 FILLER_51_3171 ();
 sg13g2_decap_8 FILLER_51_3178 ();
 sg13g2_decap_8 FILLER_51_3185 ();
 sg13g2_decap_8 FILLER_51_3192 ();
 sg13g2_decap_8 FILLER_51_3199 ();
 sg13g2_decap_8 FILLER_51_3206 ();
 sg13g2_decap_8 FILLER_51_3213 ();
 sg13g2_decap_8 FILLER_51_3220 ();
 sg13g2_decap_8 FILLER_51_3227 ();
 sg13g2_decap_8 FILLER_51_3234 ();
 sg13g2_decap_8 FILLER_51_3241 ();
 sg13g2_decap_8 FILLER_51_3248 ();
 sg13g2_decap_8 FILLER_51_3255 ();
 sg13g2_decap_8 FILLER_51_3262 ();
 sg13g2_decap_8 FILLER_51_3269 ();
 sg13g2_decap_8 FILLER_51_3276 ();
 sg13g2_decap_8 FILLER_51_3283 ();
 sg13g2_decap_8 FILLER_51_3290 ();
 sg13g2_decap_8 FILLER_51_3297 ();
 sg13g2_decap_8 FILLER_51_3304 ();
 sg13g2_decap_8 FILLER_51_3311 ();
 sg13g2_decap_8 FILLER_51_3318 ();
 sg13g2_decap_8 FILLER_51_3325 ();
 sg13g2_decap_8 FILLER_51_3332 ();
 sg13g2_decap_8 FILLER_51_3339 ();
 sg13g2_decap_8 FILLER_51_3346 ();
 sg13g2_decap_8 FILLER_51_3353 ();
 sg13g2_decap_8 FILLER_51_3360 ();
 sg13g2_decap_8 FILLER_51_3367 ();
 sg13g2_decap_8 FILLER_51_3374 ();
 sg13g2_decap_8 FILLER_51_3381 ();
 sg13g2_decap_8 FILLER_51_3388 ();
 sg13g2_decap_8 FILLER_51_3395 ();
 sg13g2_decap_8 FILLER_51_3402 ();
 sg13g2_decap_8 FILLER_51_3409 ();
 sg13g2_decap_8 FILLER_51_3416 ();
 sg13g2_decap_8 FILLER_51_3423 ();
 sg13g2_decap_8 FILLER_51_3430 ();
 sg13g2_decap_8 FILLER_51_3437 ();
 sg13g2_decap_8 FILLER_51_3444 ();
 sg13g2_decap_8 FILLER_51_3451 ();
 sg13g2_decap_8 FILLER_51_3458 ();
 sg13g2_decap_8 FILLER_51_3465 ();
 sg13g2_decap_8 FILLER_51_3472 ();
 sg13g2_decap_8 FILLER_51_3479 ();
 sg13g2_decap_8 FILLER_51_3486 ();
 sg13g2_decap_8 FILLER_51_3493 ();
 sg13g2_decap_8 FILLER_51_3500 ();
 sg13g2_decap_8 FILLER_51_3507 ();
 sg13g2_decap_8 FILLER_51_3514 ();
 sg13g2_decap_8 FILLER_51_3521 ();
 sg13g2_decap_8 FILLER_51_3528 ();
 sg13g2_decap_8 FILLER_51_3535 ();
 sg13g2_decap_8 FILLER_51_3542 ();
 sg13g2_decap_8 FILLER_51_3549 ();
 sg13g2_decap_8 FILLER_51_3556 ();
 sg13g2_decap_8 FILLER_51_3563 ();
 sg13g2_decap_8 FILLER_51_3570 ();
 sg13g2_fill_2 FILLER_51_3577 ();
 sg13g2_fill_1 FILLER_51_3579 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_decap_8 FILLER_52_112 ();
 sg13g2_decap_8 FILLER_52_119 ();
 sg13g2_decap_8 FILLER_52_126 ();
 sg13g2_decap_8 FILLER_52_133 ();
 sg13g2_decap_8 FILLER_52_140 ();
 sg13g2_decap_8 FILLER_52_147 ();
 sg13g2_decap_8 FILLER_52_154 ();
 sg13g2_decap_8 FILLER_52_161 ();
 sg13g2_decap_8 FILLER_52_168 ();
 sg13g2_decap_8 FILLER_52_175 ();
 sg13g2_decap_8 FILLER_52_182 ();
 sg13g2_decap_8 FILLER_52_189 ();
 sg13g2_decap_8 FILLER_52_196 ();
 sg13g2_decap_8 FILLER_52_203 ();
 sg13g2_decap_8 FILLER_52_210 ();
 sg13g2_decap_8 FILLER_52_217 ();
 sg13g2_decap_8 FILLER_52_224 ();
 sg13g2_decap_8 FILLER_52_231 ();
 sg13g2_decap_8 FILLER_52_238 ();
 sg13g2_decap_8 FILLER_52_245 ();
 sg13g2_decap_8 FILLER_52_252 ();
 sg13g2_decap_8 FILLER_52_259 ();
 sg13g2_decap_8 FILLER_52_266 ();
 sg13g2_decap_8 FILLER_52_273 ();
 sg13g2_decap_8 FILLER_52_280 ();
 sg13g2_decap_8 FILLER_52_287 ();
 sg13g2_decap_8 FILLER_52_294 ();
 sg13g2_decap_8 FILLER_52_301 ();
 sg13g2_decap_8 FILLER_52_308 ();
 sg13g2_decap_8 FILLER_52_315 ();
 sg13g2_decap_8 FILLER_52_322 ();
 sg13g2_decap_8 FILLER_52_329 ();
 sg13g2_decap_8 FILLER_52_336 ();
 sg13g2_decap_8 FILLER_52_343 ();
 sg13g2_decap_8 FILLER_52_350 ();
 sg13g2_decap_8 FILLER_52_357 ();
 sg13g2_decap_8 FILLER_52_364 ();
 sg13g2_decap_8 FILLER_52_371 ();
 sg13g2_decap_8 FILLER_52_378 ();
 sg13g2_decap_8 FILLER_52_385 ();
 sg13g2_decap_8 FILLER_52_392 ();
 sg13g2_decap_8 FILLER_52_399 ();
 sg13g2_decap_8 FILLER_52_406 ();
 sg13g2_decap_8 FILLER_52_413 ();
 sg13g2_decap_8 FILLER_52_420 ();
 sg13g2_decap_8 FILLER_52_427 ();
 sg13g2_decap_8 FILLER_52_434 ();
 sg13g2_decap_8 FILLER_52_441 ();
 sg13g2_decap_8 FILLER_52_448 ();
 sg13g2_decap_8 FILLER_52_455 ();
 sg13g2_decap_8 FILLER_52_462 ();
 sg13g2_decap_8 FILLER_52_469 ();
 sg13g2_decap_8 FILLER_52_476 ();
 sg13g2_decap_8 FILLER_52_483 ();
 sg13g2_decap_8 FILLER_52_490 ();
 sg13g2_decap_8 FILLER_52_497 ();
 sg13g2_decap_8 FILLER_52_504 ();
 sg13g2_decap_8 FILLER_52_511 ();
 sg13g2_decap_8 FILLER_52_518 ();
 sg13g2_decap_8 FILLER_52_525 ();
 sg13g2_decap_8 FILLER_52_532 ();
 sg13g2_decap_8 FILLER_52_539 ();
 sg13g2_decap_8 FILLER_52_546 ();
 sg13g2_decap_8 FILLER_52_553 ();
 sg13g2_decap_8 FILLER_52_560 ();
 sg13g2_decap_8 FILLER_52_567 ();
 sg13g2_decap_8 FILLER_52_574 ();
 sg13g2_decap_8 FILLER_52_581 ();
 sg13g2_decap_8 FILLER_52_588 ();
 sg13g2_decap_8 FILLER_52_595 ();
 sg13g2_decap_8 FILLER_52_602 ();
 sg13g2_decap_8 FILLER_52_609 ();
 sg13g2_decap_8 FILLER_52_616 ();
 sg13g2_decap_8 FILLER_52_623 ();
 sg13g2_decap_8 FILLER_52_630 ();
 sg13g2_decap_8 FILLER_52_637 ();
 sg13g2_decap_8 FILLER_52_644 ();
 sg13g2_decap_8 FILLER_52_651 ();
 sg13g2_decap_8 FILLER_52_658 ();
 sg13g2_decap_8 FILLER_52_665 ();
 sg13g2_decap_8 FILLER_52_672 ();
 sg13g2_decap_8 FILLER_52_679 ();
 sg13g2_decap_8 FILLER_52_686 ();
 sg13g2_decap_8 FILLER_52_693 ();
 sg13g2_decap_8 FILLER_52_700 ();
 sg13g2_decap_8 FILLER_52_707 ();
 sg13g2_decap_8 FILLER_52_714 ();
 sg13g2_decap_8 FILLER_52_721 ();
 sg13g2_decap_8 FILLER_52_728 ();
 sg13g2_decap_8 FILLER_52_735 ();
 sg13g2_decap_8 FILLER_52_742 ();
 sg13g2_decap_8 FILLER_52_749 ();
 sg13g2_decap_8 FILLER_52_756 ();
 sg13g2_decap_8 FILLER_52_763 ();
 sg13g2_decap_8 FILLER_52_770 ();
 sg13g2_decap_8 FILLER_52_777 ();
 sg13g2_decap_8 FILLER_52_784 ();
 sg13g2_decap_8 FILLER_52_791 ();
 sg13g2_decap_8 FILLER_52_798 ();
 sg13g2_decap_8 FILLER_52_805 ();
 sg13g2_decap_8 FILLER_52_812 ();
 sg13g2_decap_8 FILLER_52_819 ();
 sg13g2_decap_8 FILLER_52_826 ();
 sg13g2_decap_8 FILLER_52_833 ();
 sg13g2_decap_8 FILLER_52_840 ();
 sg13g2_decap_8 FILLER_52_847 ();
 sg13g2_decap_8 FILLER_52_854 ();
 sg13g2_decap_8 FILLER_52_861 ();
 sg13g2_decap_8 FILLER_52_868 ();
 sg13g2_decap_8 FILLER_52_875 ();
 sg13g2_decap_8 FILLER_52_882 ();
 sg13g2_decap_8 FILLER_52_889 ();
 sg13g2_decap_8 FILLER_52_896 ();
 sg13g2_decap_8 FILLER_52_903 ();
 sg13g2_decap_8 FILLER_52_910 ();
 sg13g2_decap_8 FILLER_52_917 ();
 sg13g2_decap_8 FILLER_52_924 ();
 sg13g2_decap_8 FILLER_52_931 ();
 sg13g2_decap_8 FILLER_52_938 ();
 sg13g2_decap_8 FILLER_52_945 ();
 sg13g2_decap_8 FILLER_52_952 ();
 sg13g2_decap_8 FILLER_52_959 ();
 sg13g2_decap_8 FILLER_52_966 ();
 sg13g2_decap_8 FILLER_52_973 ();
 sg13g2_decap_8 FILLER_52_980 ();
 sg13g2_decap_8 FILLER_52_987 ();
 sg13g2_decap_8 FILLER_52_994 ();
 sg13g2_decap_8 FILLER_52_1001 ();
 sg13g2_decap_8 FILLER_52_1008 ();
 sg13g2_decap_8 FILLER_52_1015 ();
 sg13g2_decap_8 FILLER_52_1022 ();
 sg13g2_decap_8 FILLER_52_1029 ();
 sg13g2_decap_8 FILLER_52_1036 ();
 sg13g2_decap_8 FILLER_52_1043 ();
 sg13g2_decap_8 FILLER_52_1050 ();
 sg13g2_decap_8 FILLER_52_1057 ();
 sg13g2_decap_8 FILLER_52_1064 ();
 sg13g2_decap_8 FILLER_52_1071 ();
 sg13g2_decap_8 FILLER_52_1078 ();
 sg13g2_decap_8 FILLER_52_1085 ();
 sg13g2_decap_8 FILLER_52_1092 ();
 sg13g2_decap_8 FILLER_52_1099 ();
 sg13g2_decap_8 FILLER_52_1106 ();
 sg13g2_decap_8 FILLER_52_1113 ();
 sg13g2_decap_8 FILLER_52_1120 ();
 sg13g2_decap_8 FILLER_52_1127 ();
 sg13g2_decap_8 FILLER_52_1134 ();
 sg13g2_decap_8 FILLER_52_1141 ();
 sg13g2_decap_8 FILLER_52_1148 ();
 sg13g2_decap_8 FILLER_52_1155 ();
 sg13g2_decap_8 FILLER_52_1162 ();
 sg13g2_decap_8 FILLER_52_1169 ();
 sg13g2_decap_8 FILLER_52_1176 ();
 sg13g2_decap_8 FILLER_52_1183 ();
 sg13g2_decap_8 FILLER_52_1190 ();
 sg13g2_decap_8 FILLER_52_1197 ();
 sg13g2_decap_8 FILLER_52_1204 ();
 sg13g2_decap_8 FILLER_52_1211 ();
 sg13g2_decap_8 FILLER_52_1218 ();
 sg13g2_decap_8 FILLER_52_1225 ();
 sg13g2_decap_8 FILLER_52_1232 ();
 sg13g2_decap_8 FILLER_52_1239 ();
 sg13g2_decap_8 FILLER_52_1246 ();
 sg13g2_decap_8 FILLER_52_1253 ();
 sg13g2_decap_8 FILLER_52_1260 ();
 sg13g2_decap_8 FILLER_52_1267 ();
 sg13g2_decap_8 FILLER_52_1274 ();
 sg13g2_decap_8 FILLER_52_1281 ();
 sg13g2_decap_8 FILLER_52_1288 ();
 sg13g2_decap_8 FILLER_52_1295 ();
 sg13g2_decap_8 FILLER_52_1302 ();
 sg13g2_decap_8 FILLER_52_1309 ();
 sg13g2_decap_8 FILLER_52_1316 ();
 sg13g2_decap_8 FILLER_52_1323 ();
 sg13g2_decap_8 FILLER_52_1330 ();
 sg13g2_decap_8 FILLER_52_1337 ();
 sg13g2_decap_8 FILLER_52_1344 ();
 sg13g2_decap_8 FILLER_52_1351 ();
 sg13g2_decap_8 FILLER_52_1358 ();
 sg13g2_decap_8 FILLER_52_1365 ();
 sg13g2_decap_8 FILLER_52_1372 ();
 sg13g2_decap_8 FILLER_52_1379 ();
 sg13g2_decap_8 FILLER_52_1386 ();
 sg13g2_decap_8 FILLER_52_1393 ();
 sg13g2_decap_8 FILLER_52_1400 ();
 sg13g2_decap_8 FILLER_52_1407 ();
 sg13g2_decap_8 FILLER_52_1414 ();
 sg13g2_decap_8 FILLER_52_1421 ();
 sg13g2_decap_8 FILLER_52_1428 ();
 sg13g2_decap_8 FILLER_52_1435 ();
 sg13g2_decap_8 FILLER_52_1442 ();
 sg13g2_decap_8 FILLER_52_1449 ();
 sg13g2_decap_8 FILLER_52_1456 ();
 sg13g2_decap_8 FILLER_52_1463 ();
 sg13g2_decap_8 FILLER_52_1470 ();
 sg13g2_decap_8 FILLER_52_1477 ();
 sg13g2_decap_8 FILLER_52_1484 ();
 sg13g2_decap_8 FILLER_52_1491 ();
 sg13g2_decap_8 FILLER_52_1498 ();
 sg13g2_decap_8 FILLER_52_1505 ();
 sg13g2_decap_8 FILLER_52_1512 ();
 sg13g2_decap_8 FILLER_52_1519 ();
 sg13g2_decap_8 FILLER_52_1526 ();
 sg13g2_decap_8 FILLER_52_1533 ();
 sg13g2_decap_8 FILLER_52_1540 ();
 sg13g2_decap_8 FILLER_52_1547 ();
 sg13g2_decap_8 FILLER_52_1554 ();
 sg13g2_decap_8 FILLER_52_1561 ();
 sg13g2_decap_8 FILLER_52_1568 ();
 sg13g2_decap_8 FILLER_52_1575 ();
 sg13g2_decap_8 FILLER_52_1582 ();
 sg13g2_decap_8 FILLER_52_1589 ();
 sg13g2_decap_8 FILLER_52_1596 ();
 sg13g2_decap_8 FILLER_52_1603 ();
 sg13g2_decap_8 FILLER_52_1610 ();
 sg13g2_decap_8 FILLER_52_1617 ();
 sg13g2_decap_8 FILLER_52_1624 ();
 sg13g2_decap_8 FILLER_52_1631 ();
 sg13g2_decap_8 FILLER_52_1638 ();
 sg13g2_decap_8 FILLER_52_1645 ();
 sg13g2_decap_8 FILLER_52_1652 ();
 sg13g2_decap_8 FILLER_52_1659 ();
 sg13g2_decap_8 FILLER_52_1666 ();
 sg13g2_decap_8 FILLER_52_1673 ();
 sg13g2_decap_8 FILLER_52_1680 ();
 sg13g2_decap_8 FILLER_52_1687 ();
 sg13g2_decap_8 FILLER_52_1694 ();
 sg13g2_decap_8 FILLER_52_1701 ();
 sg13g2_decap_8 FILLER_52_1708 ();
 sg13g2_decap_8 FILLER_52_1715 ();
 sg13g2_decap_8 FILLER_52_1722 ();
 sg13g2_decap_8 FILLER_52_1729 ();
 sg13g2_decap_8 FILLER_52_1736 ();
 sg13g2_decap_8 FILLER_52_1743 ();
 sg13g2_decap_8 FILLER_52_1750 ();
 sg13g2_decap_8 FILLER_52_1757 ();
 sg13g2_decap_8 FILLER_52_1764 ();
 sg13g2_decap_8 FILLER_52_1771 ();
 sg13g2_decap_8 FILLER_52_1778 ();
 sg13g2_decap_8 FILLER_52_1785 ();
 sg13g2_decap_8 FILLER_52_1792 ();
 sg13g2_decap_8 FILLER_52_1799 ();
 sg13g2_decap_8 FILLER_52_1806 ();
 sg13g2_decap_8 FILLER_52_1813 ();
 sg13g2_decap_8 FILLER_52_1820 ();
 sg13g2_decap_8 FILLER_52_1827 ();
 sg13g2_decap_8 FILLER_52_1834 ();
 sg13g2_decap_8 FILLER_52_1841 ();
 sg13g2_decap_8 FILLER_52_1848 ();
 sg13g2_decap_8 FILLER_52_1855 ();
 sg13g2_decap_8 FILLER_52_1862 ();
 sg13g2_decap_8 FILLER_52_1869 ();
 sg13g2_decap_8 FILLER_52_1876 ();
 sg13g2_decap_8 FILLER_52_1883 ();
 sg13g2_decap_8 FILLER_52_1890 ();
 sg13g2_decap_8 FILLER_52_1897 ();
 sg13g2_decap_8 FILLER_52_1904 ();
 sg13g2_decap_8 FILLER_52_1911 ();
 sg13g2_decap_8 FILLER_52_1918 ();
 sg13g2_decap_8 FILLER_52_1925 ();
 sg13g2_decap_8 FILLER_52_1932 ();
 sg13g2_decap_8 FILLER_52_1939 ();
 sg13g2_decap_8 FILLER_52_1946 ();
 sg13g2_decap_8 FILLER_52_1953 ();
 sg13g2_decap_8 FILLER_52_1960 ();
 sg13g2_decap_8 FILLER_52_1967 ();
 sg13g2_decap_8 FILLER_52_1974 ();
 sg13g2_decap_8 FILLER_52_1981 ();
 sg13g2_decap_8 FILLER_52_1988 ();
 sg13g2_decap_8 FILLER_52_1995 ();
 sg13g2_decap_8 FILLER_52_2002 ();
 sg13g2_decap_8 FILLER_52_2009 ();
 sg13g2_decap_8 FILLER_52_2016 ();
 sg13g2_decap_8 FILLER_52_2023 ();
 sg13g2_decap_8 FILLER_52_2030 ();
 sg13g2_decap_8 FILLER_52_2037 ();
 sg13g2_decap_8 FILLER_52_2044 ();
 sg13g2_decap_8 FILLER_52_2051 ();
 sg13g2_decap_8 FILLER_52_2058 ();
 sg13g2_decap_8 FILLER_52_2065 ();
 sg13g2_decap_8 FILLER_52_2072 ();
 sg13g2_decap_8 FILLER_52_2079 ();
 sg13g2_decap_8 FILLER_52_2086 ();
 sg13g2_decap_8 FILLER_52_2093 ();
 sg13g2_decap_8 FILLER_52_2100 ();
 sg13g2_decap_8 FILLER_52_2107 ();
 sg13g2_decap_8 FILLER_52_2114 ();
 sg13g2_decap_8 FILLER_52_2121 ();
 sg13g2_decap_8 FILLER_52_2128 ();
 sg13g2_decap_8 FILLER_52_2135 ();
 sg13g2_decap_8 FILLER_52_2142 ();
 sg13g2_decap_8 FILLER_52_2149 ();
 sg13g2_decap_8 FILLER_52_2156 ();
 sg13g2_decap_8 FILLER_52_2163 ();
 sg13g2_decap_8 FILLER_52_2170 ();
 sg13g2_decap_8 FILLER_52_2177 ();
 sg13g2_decap_8 FILLER_52_2184 ();
 sg13g2_decap_8 FILLER_52_2191 ();
 sg13g2_decap_8 FILLER_52_2198 ();
 sg13g2_decap_8 FILLER_52_2205 ();
 sg13g2_decap_8 FILLER_52_2212 ();
 sg13g2_decap_8 FILLER_52_2219 ();
 sg13g2_decap_8 FILLER_52_2226 ();
 sg13g2_decap_8 FILLER_52_2233 ();
 sg13g2_decap_8 FILLER_52_2240 ();
 sg13g2_decap_8 FILLER_52_2247 ();
 sg13g2_decap_8 FILLER_52_2254 ();
 sg13g2_decap_8 FILLER_52_2261 ();
 sg13g2_decap_8 FILLER_52_2268 ();
 sg13g2_decap_8 FILLER_52_2275 ();
 sg13g2_decap_8 FILLER_52_2282 ();
 sg13g2_decap_8 FILLER_52_2289 ();
 sg13g2_decap_8 FILLER_52_2296 ();
 sg13g2_decap_8 FILLER_52_2303 ();
 sg13g2_decap_8 FILLER_52_2310 ();
 sg13g2_decap_8 FILLER_52_2317 ();
 sg13g2_decap_8 FILLER_52_2324 ();
 sg13g2_decap_8 FILLER_52_2331 ();
 sg13g2_decap_8 FILLER_52_2338 ();
 sg13g2_decap_8 FILLER_52_2345 ();
 sg13g2_decap_8 FILLER_52_2352 ();
 sg13g2_decap_8 FILLER_52_2359 ();
 sg13g2_decap_8 FILLER_52_2366 ();
 sg13g2_decap_8 FILLER_52_2373 ();
 sg13g2_decap_8 FILLER_52_2380 ();
 sg13g2_decap_8 FILLER_52_2387 ();
 sg13g2_decap_8 FILLER_52_2394 ();
 sg13g2_decap_8 FILLER_52_2401 ();
 sg13g2_decap_8 FILLER_52_2408 ();
 sg13g2_decap_8 FILLER_52_2415 ();
 sg13g2_decap_8 FILLER_52_2422 ();
 sg13g2_decap_8 FILLER_52_2429 ();
 sg13g2_decap_8 FILLER_52_2436 ();
 sg13g2_decap_8 FILLER_52_2443 ();
 sg13g2_decap_8 FILLER_52_2450 ();
 sg13g2_decap_8 FILLER_52_2457 ();
 sg13g2_decap_8 FILLER_52_2464 ();
 sg13g2_decap_8 FILLER_52_2471 ();
 sg13g2_decap_8 FILLER_52_2478 ();
 sg13g2_decap_8 FILLER_52_2485 ();
 sg13g2_decap_8 FILLER_52_2492 ();
 sg13g2_decap_8 FILLER_52_2499 ();
 sg13g2_decap_8 FILLER_52_2506 ();
 sg13g2_decap_8 FILLER_52_2513 ();
 sg13g2_decap_8 FILLER_52_2520 ();
 sg13g2_decap_8 FILLER_52_2527 ();
 sg13g2_decap_8 FILLER_52_2534 ();
 sg13g2_decap_8 FILLER_52_2541 ();
 sg13g2_decap_8 FILLER_52_2548 ();
 sg13g2_decap_8 FILLER_52_2555 ();
 sg13g2_decap_8 FILLER_52_2562 ();
 sg13g2_decap_8 FILLER_52_2569 ();
 sg13g2_decap_8 FILLER_52_2576 ();
 sg13g2_decap_8 FILLER_52_2583 ();
 sg13g2_decap_8 FILLER_52_2590 ();
 sg13g2_decap_8 FILLER_52_2597 ();
 sg13g2_decap_8 FILLER_52_2604 ();
 sg13g2_decap_8 FILLER_52_2611 ();
 sg13g2_decap_8 FILLER_52_2618 ();
 sg13g2_decap_8 FILLER_52_2625 ();
 sg13g2_decap_8 FILLER_52_2632 ();
 sg13g2_decap_8 FILLER_52_2639 ();
 sg13g2_decap_8 FILLER_52_2646 ();
 sg13g2_decap_8 FILLER_52_2653 ();
 sg13g2_decap_8 FILLER_52_2660 ();
 sg13g2_decap_8 FILLER_52_2667 ();
 sg13g2_decap_8 FILLER_52_2674 ();
 sg13g2_decap_8 FILLER_52_2681 ();
 sg13g2_decap_8 FILLER_52_2688 ();
 sg13g2_decap_8 FILLER_52_2695 ();
 sg13g2_decap_8 FILLER_52_2702 ();
 sg13g2_decap_8 FILLER_52_2709 ();
 sg13g2_decap_8 FILLER_52_2716 ();
 sg13g2_decap_8 FILLER_52_2723 ();
 sg13g2_decap_8 FILLER_52_2730 ();
 sg13g2_decap_8 FILLER_52_2737 ();
 sg13g2_decap_8 FILLER_52_2744 ();
 sg13g2_decap_8 FILLER_52_2751 ();
 sg13g2_decap_8 FILLER_52_2758 ();
 sg13g2_decap_8 FILLER_52_2765 ();
 sg13g2_decap_8 FILLER_52_2772 ();
 sg13g2_decap_8 FILLER_52_2779 ();
 sg13g2_decap_8 FILLER_52_2786 ();
 sg13g2_decap_8 FILLER_52_2793 ();
 sg13g2_decap_8 FILLER_52_2800 ();
 sg13g2_decap_8 FILLER_52_2807 ();
 sg13g2_decap_8 FILLER_52_2814 ();
 sg13g2_decap_8 FILLER_52_2821 ();
 sg13g2_decap_8 FILLER_52_2828 ();
 sg13g2_decap_8 FILLER_52_2835 ();
 sg13g2_decap_8 FILLER_52_2842 ();
 sg13g2_decap_8 FILLER_52_2849 ();
 sg13g2_decap_8 FILLER_52_2856 ();
 sg13g2_decap_8 FILLER_52_2863 ();
 sg13g2_decap_8 FILLER_52_2870 ();
 sg13g2_decap_8 FILLER_52_2877 ();
 sg13g2_decap_8 FILLER_52_2884 ();
 sg13g2_decap_8 FILLER_52_2891 ();
 sg13g2_decap_8 FILLER_52_2898 ();
 sg13g2_decap_8 FILLER_52_2905 ();
 sg13g2_decap_8 FILLER_52_2912 ();
 sg13g2_decap_8 FILLER_52_2919 ();
 sg13g2_decap_8 FILLER_52_2926 ();
 sg13g2_decap_8 FILLER_52_2933 ();
 sg13g2_decap_8 FILLER_52_2940 ();
 sg13g2_decap_8 FILLER_52_2947 ();
 sg13g2_decap_8 FILLER_52_2954 ();
 sg13g2_decap_8 FILLER_52_2961 ();
 sg13g2_decap_8 FILLER_52_2968 ();
 sg13g2_decap_8 FILLER_52_2975 ();
 sg13g2_decap_8 FILLER_52_2982 ();
 sg13g2_decap_8 FILLER_52_2989 ();
 sg13g2_decap_8 FILLER_52_2996 ();
 sg13g2_decap_8 FILLER_52_3003 ();
 sg13g2_decap_8 FILLER_52_3010 ();
 sg13g2_decap_8 FILLER_52_3017 ();
 sg13g2_decap_8 FILLER_52_3024 ();
 sg13g2_decap_8 FILLER_52_3031 ();
 sg13g2_decap_8 FILLER_52_3038 ();
 sg13g2_decap_8 FILLER_52_3045 ();
 sg13g2_decap_8 FILLER_52_3052 ();
 sg13g2_decap_8 FILLER_52_3059 ();
 sg13g2_decap_8 FILLER_52_3066 ();
 sg13g2_decap_8 FILLER_52_3073 ();
 sg13g2_decap_8 FILLER_52_3080 ();
 sg13g2_decap_8 FILLER_52_3087 ();
 sg13g2_decap_8 FILLER_52_3094 ();
 sg13g2_decap_8 FILLER_52_3101 ();
 sg13g2_decap_8 FILLER_52_3108 ();
 sg13g2_decap_8 FILLER_52_3115 ();
 sg13g2_decap_8 FILLER_52_3122 ();
 sg13g2_decap_8 FILLER_52_3129 ();
 sg13g2_decap_8 FILLER_52_3136 ();
 sg13g2_decap_8 FILLER_52_3143 ();
 sg13g2_decap_8 FILLER_52_3150 ();
 sg13g2_decap_8 FILLER_52_3157 ();
 sg13g2_decap_8 FILLER_52_3164 ();
 sg13g2_decap_8 FILLER_52_3171 ();
 sg13g2_decap_8 FILLER_52_3178 ();
 sg13g2_decap_8 FILLER_52_3185 ();
 sg13g2_decap_8 FILLER_52_3192 ();
 sg13g2_decap_8 FILLER_52_3199 ();
 sg13g2_decap_8 FILLER_52_3206 ();
 sg13g2_decap_8 FILLER_52_3213 ();
 sg13g2_decap_8 FILLER_52_3220 ();
 sg13g2_decap_8 FILLER_52_3227 ();
 sg13g2_decap_8 FILLER_52_3234 ();
 sg13g2_decap_8 FILLER_52_3241 ();
 sg13g2_decap_8 FILLER_52_3248 ();
 sg13g2_decap_8 FILLER_52_3255 ();
 sg13g2_decap_8 FILLER_52_3262 ();
 sg13g2_decap_8 FILLER_52_3269 ();
 sg13g2_decap_8 FILLER_52_3276 ();
 sg13g2_decap_8 FILLER_52_3283 ();
 sg13g2_decap_8 FILLER_52_3290 ();
 sg13g2_decap_8 FILLER_52_3297 ();
 sg13g2_decap_8 FILLER_52_3304 ();
 sg13g2_decap_8 FILLER_52_3311 ();
 sg13g2_decap_8 FILLER_52_3318 ();
 sg13g2_decap_8 FILLER_52_3325 ();
 sg13g2_decap_8 FILLER_52_3332 ();
 sg13g2_decap_8 FILLER_52_3339 ();
 sg13g2_decap_8 FILLER_52_3346 ();
 sg13g2_decap_8 FILLER_52_3353 ();
 sg13g2_decap_8 FILLER_52_3360 ();
 sg13g2_decap_8 FILLER_52_3367 ();
 sg13g2_decap_8 FILLER_52_3374 ();
 sg13g2_decap_8 FILLER_52_3381 ();
 sg13g2_decap_8 FILLER_52_3388 ();
 sg13g2_decap_8 FILLER_52_3395 ();
 sg13g2_decap_8 FILLER_52_3402 ();
 sg13g2_decap_8 FILLER_52_3409 ();
 sg13g2_decap_8 FILLER_52_3416 ();
 sg13g2_decap_8 FILLER_52_3423 ();
 sg13g2_decap_8 FILLER_52_3430 ();
 sg13g2_decap_8 FILLER_52_3437 ();
 sg13g2_decap_8 FILLER_52_3444 ();
 sg13g2_decap_8 FILLER_52_3451 ();
 sg13g2_decap_8 FILLER_52_3458 ();
 sg13g2_decap_8 FILLER_52_3465 ();
 sg13g2_decap_8 FILLER_52_3472 ();
 sg13g2_decap_8 FILLER_52_3479 ();
 sg13g2_decap_8 FILLER_52_3486 ();
 sg13g2_decap_8 FILLER_52_3493 ();
 sg13g2_decap_8 FILLER_52_3500 ();
 sg13g2_decap_8 FILLER_52_3507 ();
 sg13g2_decap_8 FILLER_52_3514 ();
 sg13g2_decap_8 FILLER_52_3521 ();
 sg13g2_decap_8 FILLER_52_3528 ();
 sg13g2_decap_8 FILLER_52_3535 ();
 sg13g2_decap_8 FILLER_52_3542 ();
 sg13g2_decap_8 FILLER_52_3549 ();
 sg13g2_decap_8 FILLER_52_3556 ();
 sg13g2_decap_8 FILLER_52_3563 ();
 sg13g2_decap_8 FILLER_52_3570 ();
 sg13g2_fill_2 FILLER_52_3577 ();
 sg13g2_fill_1 FILLER_52_3579 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_8 FILLER_53_105 ();
 sg13g2_decap_8 FILLER_53_112 ();
 sg13g2_decap_8 FILLER_53_119 ();
 sg13g2_decap_8 FILLER_53_126 ();
 sg13g2_decap_8 FILLER_53_133 ();
 sg13g2_decap_8 FILLER_53_140 ();
 sg13g2_decap_8 FILLER_53_147 ();
 sg13g2_decap_8 FILLER_53_154 ();
 sg13g2_decap_8 FILLER_53_161 ();
 sg13g2_decap_8 FILLER_53_168 ();
 sg13g2_decap_8 FILLER_53_175 ();
 sg13g2_decap_8 FILLER_53_182 ();
 sg13g2_decap_8 FILLER_53_189 ();
 sg13g2_decap_8 FILLER_53_196 ();
 sg13g2_decap_8 FILLER_53_203 ();
 sg13g2_decap_8 FILLER_53_210 ();
 sg13g2_decap_8 FILLER_53_217 ();
 sg13g2_decap_8 FILLER_53_224 ();
 sg13g2_decap_8 FILLER_53_231 ();
 sg13g2_decap_8 FILLER_53_238 ();
 sg13g2_decap_8 FILLER_53_245 ();
 sg13g2_decap_8 FILLER_53_252 ();
 sg13g2_decap_8 FILLER_53_259 ();
 sg13g2_decap_8 FILLER_53_266 ();
 sg13g2_decap_8 FILLER_53_273 ();
 sg13g2_decap_8 FILLER_53_280 ();
 sg13g2_decap_8 FILLER_53_287 ();
 sg13g2_decap_8 FILLER_53_294 ();
 sg13g2_decap_8 FILLER_53_301 ();
 sg13g2_decap_8 FILLER_53_308 ();
 sg13g2_decap_8 FILLER_53_315 ();
 sg13g2_decap_8 FILLER_53_322 ();
 sg13g2_decap_8 FILLER_53_329 ();
 sg13g2_decap_8 FILLER_53_336 ();
 sg13g2_decap_8 FILLER_53_343 ();
 sg13g2_decap_8 FILLER_53_350 ();
 sg13g2_decap_8 FILLER_53_357 ();
 sg13g2_decap_8 FILLER_53_364 ();
 sg13g2_decap_8 FILLER_53_371 ();
 sg13g2_decap_8 FILLER_53_378 ();
 sg13g2_decap_8 FILLER_53_385 ();
 sg13g2_decap_8 FILLER_53_392 ();
 sg13g2_decap_8 FILLER_53_399 ();
 sg13g2_decap_8 FILLER_53_406 ();
 sg13g2_decap_8 FILLER_53_413 ();
 sg13g2_decap_8 FILLER_53_420 ();
 sg13g2_decap_8 FILLER_53_427 ();
 sg13g2_decap_8 FILLER_53_434 ();
 sg13g2_decap_8 FILLER_53_441 ();
 sg13g2_decap_8 FILLER_53_448 ();
 sg13g2_decap_8 FILLER_53_455 ();
 sg13g2_decap_8 FILLER_53_462 ();
 sg13g2_decap_8 FILLER_53_469 ();
 sg13g2_decap_8 FILLER_53_476 ();
 sg13g2_decap_8 FILLER_53_483 ();
 sg13g2_decap_8 FILLER_53_490 ();
 sg13g2_decap_8 FILLER_53_497 ();
 sg13g2_decap_8 FILLER_53_504 ();
 sg13g2_decap_8 FILLER_53_511 ();
 sg13g2_decap_8 FILLER_53_518 ();
 sg13g2_decap_8 FILLER_53_525 ();
 sg13g2_decap_8 FILLER_53_532 ();
 sg13g2_decap_8 FILLER_53_539 ();
 sg13g2_decap_8 FILLER_53_546 ();
 sg13g2_decap_8 FILLER_53_553 ();
 sg13g2_decap_8 FILLER_53_560 ();
 sg13g2_decap_8 FILLER_53_567 ();
 sg13g2_decap_8 FILLER_53_574 ();
 sg13g2_decap_8 FILLER_53_581 ();
 sg13g2_decap_8 FILLER_53_588 ();
 sg13g2_decap_8 FILLER_53_595 ();
 sg13g2_decap_8 FILLER_53_602 ();
 sg13g2_decap_8 FILLER_53_609 ();
 sg13g2_decap_8 FILLER_53_616 ();
 sg13g2_decap_8 FILLER_53_623 ();
 sg13g2_decap_8 FILLER_53_630 ();
 sg13g2_decap_8 FILLER_53_637 ();
 sg13g2_decap_8 FILLER_53_644 ();
 sg13g2_decap_8 FILLER_53_651 ();
 sg13g2_decap_8 FILLER_53_658 ();
 sg13g2_decap_8 FILLER_53_665 ();
 sg13g2_decap_8 FILLER_53_672 ();
 sg13g2_decap_8 FILLER_53_679 ();
 sg13g2_decap_8 FILLER_53_686 ();
 sg13g2_decap_8 FILLER_53_693 ();
 sg13g2_decap_8 FILLER_53_700 ();
 sg13g2_decap_8 FILLER_53_707 ();
 sg13g2_decap_8 FILLER_53_714 ();
 sg13g2_decap_8 FILLER_53_721 ();
 sg13g2_decap_8 FILLER_53_728 ();
 sg13g2_decap_8 FILLER_53_735 ();
 sg13g2_decap_8 FILLER_53_742 ();
 sg13g2_decap_8 FILLER_53_749 ();
 sg13g2_decap_8 FILLER_53_756 ();
 sg13g2_decap_8 FILLER_53_763 ();
 sg13g2_decap_8 FILLER_53_770 ();
 sg13g2_decap_8 FILLER_53_777 ();
 sg13g2_decap_8 FILLER_53_784 ();
 sg13g2_decap_8 FILLER_53_791 ();
 sg13g2_decap_8 FILLER_53_798 ();
 sg13g2_decap_8 FILLER_53_805 ();
 sg13g2_decap_8 FILLER_53_812 ();
 sg13g2_decap_8 FILLER_53_819 ();
 sg13g2_decap_8 FILLER_53_826 ();
 sg13g2_decap_8 FILLER_53_833 ();
 sg13g2_decap_8 FILLER_53_840 ();
 sg13g2_decap_8 FILLER_53_847 ();
 sg13g2_decap_8 FILLER_53_854 ();
 sg13g2_decap_8 FILLER_53_861 ();
 sg13g2_decap_8 FILLER_53_868 ();
 sg13g2_decap_8 FILLER_53_875 ();
 sg13g2_decap_8 FILLER_53_882 ();
 sg13g2_decap_8 FILLER_53_889 ();
 sg13g2_decap_8 FILLER_53_896 ();
 sg13g2_decap_8 FILLER_53_903 ();
 sg13g2_decap_8 FILLER_53_910 ();
 sg13g2_decap_8 FILLER_53_917 ();
 sg13g2_decap_8 FILLER_53_924 ();
 sg13g2_decap_8 FILLER_53_931 ();
 sg13g2_decap_8 FILLER_53_938 ();
 sg13g2_decap_8 FILLER_53_945 ();
 sg13g2_decap_8 FILLER_53_952 ();
 sg13g2_decap_8 FILLER_53_959 ();
 sg13g2_decap_8 FILLER_53_966 ();
 sg13g2_decap_8 FILLER_53_973 ();
 sg13g2_decap_8 FILLER_53_980 ();
 sg13g2_decap_8 FILLER_53_987 ();
 sg13g2_decap_8 FILLER_53_994 ();
 sg13g2_decap_8 FILLER_53_1001 ();
 sg13g2_decap_8 FILLER_53_1008 ();
 sg13g2_decap_8 FILLER_53_1015 ();
 sg13g2_decap_8 FILLER_53_1022 ();
 sg13g2_decap_8 FILLER_53_1029 ();
 sg13g2_decap_8 FILLER_53_1036 ();
 sg13g2_decap_8 FILLER_53_1043 ();
 sg13g2_decap_8 FILLER_53_1050 ();
 sg13g2_decap_8 FILLER_53_1057 ();
 sg13g2_decap_8 FILLER_53_1064 ();
 sg13g2_decap_8 FILLER_53_1071 ();
 sg13g2_decap_8 FILLER_53_1078 ();
 sg13g2_decap_8 FILLER_53_1085 ();
 sg13g2_decap_8 FILLER_53_1092 ();
 sg13g2_decap_8 FILLER_53_1099 ();
 sg13g2_decap_8 FILLER_53_1106 ();
 sg13g2_decap_8 FILLER_53_1113 ();
 sg13g2_decap_8 FILLER_53_1120 ();
 sg13g2_decap_8 FILLER_53_1127 ();
 sg13g2_decap_8 FILLER_53_1134 ();
 sg13g2_decap_8 FILLER_53_1141 ();
 sg13g2_decap_8 FILLER_53_1148 ();
 sg13g2_decap_8 FILLER_53_1155 ();
 sg13g2_decap_8 FILLER_53_1162 ();
 sg13g2_decap_8 FILLER_53_1169 ();
 sg13g2_decap_8 FILLER_53_1176 ();
 sg13g2_decap_8 FILLER_53_1183 ();
 sg13g2_decap_8 FILLER_53_1190 ();
 sg13g2_decap_8 FILLER_53_1197 ();
 sg13g2_decap_8 FILLER_53_1204 ();
 sg13g2_decap_8 FILLER_53_1211 ();
 sg13g2_decap_8 FILLER_53_1218 ();
 sg13g2_decap_8 FILLER_53_1225 ();
 sg13g2_decap_8 FILLER_53_1232 ();
 sg13g2_decap_8 FILLER_53_1239 ();
 sg13g2_decap_8 FILLER_53_1246 ();
 sg13g2_decap_8 FILLER_53_1253 ();
 sg13g2_decap_8 FILLER_53_1260 ();
 sg13g2_decap_8 FILLER_53_1267 ();
 sg13g2_decap_8 FILLER_53_1274 ();
 sg13g2_decap_8 FILLER_53_1281 ();
 sg13g2_decap_8 FILLER_53_1288 ();
 sg13g2_decap_8 FILLER_53_1295 ();
 sg13g2_decap_8 FILLER_53_1302 ();
 sg13g2_decap_8 FILLER_53_1309 ();
 sg13g2_decap_8 FILLER_53_1316 ();
 sg13g2_decap_8 FILLER_53_1323 ();
 sg13g2_decap_8 FILLER_53_1330 ();
 sg13g2_decap_8 FILLER_53_1337 ();
 sg13g2_decap_8 FILLER_53_1344 ();
 sg13g2_decap_8 FILLER_53_1351 ();
 sg13g2_decap_8 FILLER_53_1358 ();
 sg13g2_decap_8 FILLER_53_1365 ();
 sg13g2_decap_8 FILLER_53_1372 ();
 sg13g2_decap_8 FILLER_53_1379 ();
 sg13g2_decap_8 FILLER_53_1386 ();
 sg13g2_decap_8 FILLER_53_1393 ();
 sg13g2_decap_8 FILLER_53_1400 ();
 sg13g2_decap_8 FILLER_53_1407 ();
 sg13g2_decap_8 FILLER_53_1414 ();
 sg13g2_decap_8 FILLER_53_1421 ();
 sg13g2_decap_8 FILLER_53_1428 ();
 sg13g2_decap_8 FILLER_53_1435 ();
 sg13g2_decap_8 FILLER_53_1442 ();
 sg13g2_decap_8 FILLER_53_1449 ();
 sg13g2_decap_8 FILLER_53_1456 ();
 sg13g2_decap_8 FILLER_53_1463 ();
 sg13g2_decap_8 FILLER_53_1470 ();
 sg13g2_decap_8 FILLER_53_1477 ();
 sg13g2_decap_8 FILLER_53_1484 ();
 sg13g2_decap_8 FILLER_53_1491 ();
 sg13g2_decap_8 FILLER_53_1498 ();
 sg13g2_decap_8 FILLER_53_1505 ();
 sg13g2_decap_8 FILLER_53_1512 ();
 sg13g2_decap_8 FILLER_53_1519 ();
 sg13g2_decap_8 FILLER_53_1526 ();
 sg13g2_decap_8 FILLER_53_1533 ();
 sg13g2_decap_8 FILLER_53_1540 ();
 sg13g2_decap_8 FILLER_53_1547 ();
 sg13g2_decap_8 FILLER_53_1554 ();
 sg13g2_decap_8 FILLER_53_1561 ();
 sg13g2_decap_8 FILLER_53_1568 ();
 sg13g2_decap_8 FILLER_53_1575 ();
 sg13g2_decap_8 FILLER_53_1582 ();
 sg13g2_decap_8 FILLER_53_1589 ();
 sg13g2_decap_8 FILLER_53_1596 ();
 sg13g2_decap_8 FILLER_53_1603 ();
 sg13g2_decap_8 FILLER_53_1610 ();
 sg13g2_decap_8 FILLER_53_1617 ();
 sg13g2_decap_8 FILLER_53_1624 ();
 sg13g2_decap_8 FILLER_53_1631 ();
 sg13g2_decap_8 FILLER_53_1638 ();
 sg13g2_decap_8 FILLER_53_1645 ();
 sg13g2_decap_8 FILLER_53_1652 ();
 sg13g2_decap_8 FILLER_53_1659 ();
 sg13g2_decap_8 FILLER_53_1666 ();
 sg13g2_decap_8 FILLER_53_1673 ();
 sg13g2_decap_8 FILLER_53_1680 ();
 sg13g2_decap_8 FILLER_53_1687 ();
 sg13g2_decap_8 FILLER_53_1694 ();
 sg13g2_decap_8 FILLER_53_1701 ();
 sg13g2_decap_8 FILLER_53_1708 ();
 sg13g2_decap_8 FILLER_53_1715 ();
 sg13g2_decap_8 FILLER_53_1722 ();
 sg13g2_decap_8 FILLER_53_1729 ();
 sg13g2_decap_8 FILLER_53_1736 ();
 sg13g2_decap_8 FILLER_53_1743 ();
 sg13g2_decap_8 FILLER_53_1750 ();
 sg13g2_decap_8 FILLER_53_1757 ();
 sg13g2_decap_8 FILLER_53_1764 ();
 sg13g2_decap_8 FILLER_53_1771 ();
 sg13g2_decap_8 FILLER_53_1778 ();
 sg13g2_decap_8 FILLER_53_1785 ();
 sg13g2_decap_8 FILLER_53_1792 ();
 sg13g2_decap_8 FILLER_53_1799 ();
 sg13g2_decap_8 FILLER_53_1806 ();
 sg13g2_decap_8 FILLER_53_1813 ();
 sg13g2_decap_8 FILLER_53_1820 ();
 sg13g2_decap_8 FILLER_53_1827 ();
 sg13g2_decap_8 FILLER_53_1834 ();
 sg13g2_decap_8 FILLER_53_1841 ();
 sg13g2_decap_8 FILLER_53_1848 ();
 sg13g2_decap_8 FILLER_53_1855 ();
 sg13g2_decap_8 FILLER_53_1862 ();
 sg13g2_decap_8 FILLER_53_1869 ();
 sg13g2_decap_8 FILLER_53_1876 ();
 sg13g2_decap_8 FILLER_53_1883 ();
 sg13g2_decap_8 FILLER_53_1890 ();
 sg13g2_decap_8 FILLER_53_1897 ();
 sg13g2_decap_8 FILLER_53_1904 ();
 sg13g2_decap_8 FILLER_53_1911 ();
 sg13g2_decap_8 FILLER_53_1918 ();
 sg13g2_decap_8 FILLER_53_1925 ();
 sg13g2_decap_8 FILLER_53_1932 ();
 sg13g2_decap_8 FILLER_53_1939 ();
 sg13g2_decap_8 FILLER_53_1946 ();
 sg13g2_decap_8 FILLER_53_1953 ();
 sg13g2_decap_8 FILLER_53_1960 ();
 sg13g2_decap_8 FILLER_53_1967 ();
 sg13g2_decap_8 FILLER_53_1974 ();
 sg13g2_decap_8 FILLER_53_1981 ();
 sg13g2_decap_8 FILLER_53_1988 ();
 sg13g2_decap_8 FILLER_53_1995 ();
 sg13g2_decap_8 FILLER_53_2002 ();
 sg13g2_decap_8 FILLER_53_2009 ();
 sg13g2_decap_8 FILLER_53_2016 ();
 sg13g2_decap_8 FILLER_53_2023 ();
 sg13g2_decap_8 FILLER_53_2030 ();
 sg13g2_decap_8 FILLER_53_2037 ();
 sg13g2_decap_8 FILLER_53_2044 ();
 sg13g2_decap_8 FILLER_53_2051 ();
 sg13g2_decap_8 FILLER_53_2058 ();
 sg13g2_decap_8 FILLER_53_2065 ();
 sg13g2_decap_8 FILLER_53_2072 ();
 sg13g2_decap_8 FILLER_53_2079 ();
 sg13g2_decap_8 FILLER_53_2086 ();
 sg13g2_decap_8 FILLER_53_2093 ();
 sg13g2_decap_8 FILLER_53_2100 ();
 sg13g2_decap_8 FILLER_53_2107 ();
 sg13g2_decap_8 FILLER_53_2114 ();
 sg13g2_decap_8 FILLER_53_2121 ();
 sg13g2_decap_8 FILLER_53_2128 ();
 sg13g2_decap_8 FILLER_53_2135 ();
 sg13g2_decap_8 FILLER_53_2142 ();
 sg13g2_decap_8 FILLER_53_2149 ();
 sg13g2_decap_8 FILLER_53_2156 ();
 sg13g2_decap_8 FILLER_53_2163 ();
 sg13g2_decap_8 FILLER_53_2170 ();
 sg13g2_decap_8 FILLER_53_2177 ();
 sg13g2_decap_8 FILLER_53_2184 ();
 sg13g2_decap_8 FILLER_53_2191 ();
 sg13g2_decap_8 FILLER_53_2198 ();
 sg13g2_decap_8 FILLER_53_2205 ();
 sg13g2_decap_8 FILLER_53_2212 ();
 sg13g2_decap_8 FILLER_53_2219 ();
 sg13g2_decap_8 FILLER_53_2226 ();
 sg13g2_decap_8 FILLER_53_2233 ();
 sg13g2_decap_8 FILLER_53_2240 ();
 sg13g2_decap_8 FILLER_53_2247 ();
 sg13g2_decap_8 FILLER_53_2254 ();
 sg13g2_decap_8 FILLER_53_2261 ();
 sg13g2_decap_8 FILLER_53_2268 ();
 sg13g2_decap_8 FILLER_53_2275 ();
 sg13g2_decap_8 FILLER_53_2282 ();
 sg13g2_decap_8 FILLER_53_2289 ();
 sg13g2_decap_8 FILLER_53_2296 ();
 sg13g2_decap_8 FILLER_53_2303 ();
 sg13g2_decap_8 FILLER_53_2310 ();
 sg13g2_decap_8 FILLER_53_2317 ();
 sg13g2_decap_8 FILLER_53_2324 ();
 sg13g2_decap_8 FILLER_53_2331 ();
 sg13g2_decap_8 FILLER_53_2338 ();
 sg13g2_decap_8 FILLER_53_2345 ();
 sg13g2_decap_8 FILLER_53_2352 ();
 sg13g2_decap_8 FILLER_53_2359 ();
 sg13g2_decap_8 FILLER_53_2366 ();
 sg13g2_decap_8 FILLER_53_2373 ();
 sg13g2_decap_8 FILLER_53_2380 ();
 sg13g2_decap_8 FILLER_53_2387 ();
 sg13g2_decap_8 FILLER_53_2394 ();
 sg13g2_decap_8 FILLER_53_2401 ();
 sg13g2_decap_8 FILLER_53_2408 ();
 sg13g2_decap_8 FILLER_53_2415 ();
 sg13g2_decap_8 FILLER_53_2422 ();
 sg13g2_decap_8 FILLER_53_2429 ();
 sg13g2_decap_8 FILLER_53_2436 ();
 sg13g2_decap_8 FILLER_53_2443 ();
 sg13g2_decap_8 FILLER_53_2450 ();
 sg13g2_decap_8 FILLER_53_2457 ();
 sg13g2_decap_8 FILLER_53_2464 ();
 sg13g2_decap_8 FILLER_53_2471 ();
 sg13g2_decap_8 FILLER_53_2478 ();
 sg13g2_decap_8 FILLER_53_2485 ();
 sg13g2_decap_8 FILLER_53_2492 ();
 sg13g2_decap_8 FILLER_53_2499 ();
 sg13g2_decap_8 FILLER_53_2506 ();
 sg13g2_decap_8 FILLER_53_2513 ();
 sg13g2_decap_8 FILLER_53_2520 ();
 sg13g2_decap_8 FILLER_53_2527 ();
 sg13g2_decap_8 FILLER_53_2534 ();
 sg13g2_decap_8 FILLER_53_2541 ();
 sg13g2_decap_8 FILLER_53_2548 ();
 sg13g2_decap_8 FILLER_53_2555 ();
 sg13g2_decap_8 FILLER_53_2562 ();
 sg13g2_decap_8 FILLER_53_2569 ();
 sg13g2_decap_8 FILLER_53_2576 ();
 sg13g2_decap_8 FILLER_53_2583 ();
 sg13g2_decap_8 FILLER_53_2590 ();
 sg13g2_decap_8 FILLER_53_2597 ();
 sg13g2_decap_8 FILLER_53_2604 ();
 sg13g2_decap_8 FILLER_53_2611 ();
 sg13g2_decap_8 FILLER_53_2618 ();
 sg13g2_decap_8 FILLER_53_2625 ();
 sg13g2_decap_8 FILLER_53_2632 ();
 sg13g2_decap_8 FILLER_53_2639 ();
 sg13g2_decap_8 FILLER_53_2646 ();
 sg13g2_decap_8 FILLER_53_2653 ();
 sg13g2_decap_8 FILLER_53_2660 ();
 sg13g2_decap_8 FILLER_53_2667 ();
 sg13g2_decap_8 FILLER_53_2674 ();
 sg13g2_decap_8 FILLER_53_2681 ();
 sg13g2_decap_8 FILLER_53_2688 ();
 sg13g2_decap_8 FILLER_53_2695 ();
 sg13g2_decap_8 FILLER_53_2702 ();
 sg13g2_decap_8 FILLER_53_2709 ();
 sg13g2_decap_8 FILLER_53_2716 ();
 sg13g2_decap_8 FILLER_53_2723 ();
 sg13g2_decap_8 FILLER_53_2730 ();
 sg13g2_decap_8 FILLER_53_2737 ();
 sg13g2_decap_8 FILLER_53_2744 ();
 sg13g2_decap_8 FILLER_53_2751 ();
 sg13g2_decap_8 FILLER_53_2758 ();
 sg13g2_decap_8 FILLER_53_2765 ();
 sg13g2_decap_8 FILLER_53_2772 ();
 sg13g2_decap_8 FILLER_53_2779 ();
 sg13g2_decap_8 FILLER_53_2786 ();
 sg13g2_decap_8 FILLER_53_2793 ();
 sg13g2_decap_8 FILLER_53_2800 ();
 sg13g2_decap_8 FILLER_53_2807 ();
 sg13g2_decap_8 FILLER_53_2814 ();
 sg13g2_decap_8 FILLER_53_2821 ();
 sg13g2_decap_8 FILLER_53_2828 ();
 sg13g2_decap_8 FILLER_53_2835 ();
 sg13g2_decap_8 FILLER_53_2842 ();
 sg13g2_decap_8 FILLER_53_2849 ();
 sg13g2_decap_8 FILLER_53_2856 ();
 sg13g2_decap_8 FILLER_53_2863 ();
 sg13g2_decap_8 FILLER_53_2870 ();
 sg13g2_decap_8 FILLER_53_2877 ();
 sg13g2_decap_8 FILLER_53_2884 ();
 sg13g2_decap_8 FILLER_53_2891 ();
 sg13g2_decap_8 FILLER_53_2898 ();
 sg13g2_decap_8 FILLER_53_2905 ();
 sg13g2_decap_8 FILLER_53_2912 ();
 sg13g2_decap_8 FILLER_53_2919 ();
 sg13g2_decap_8 FILLER_53_2926 ();
 sg13g2_decap_8 FILLER_53_2933 ();
 sg13g2_decap_8 FILLER_53_2940 ();
 sg13g2_decap_8 FILLER_53_2947 ();
 sg13g2_decap_8 FILLER_53_2954 ();
 sg13g2_decap_8 FILLER_53_2961 ();
 sg13g2_decap_8 FILLER_53_2968 ();
 sg13g2_decap_8 FILLER_53_2975 ();
 sg13g2_decap_8 FILLER_53_2982 ();
 sg13g2_decap_8 FILLER_53_2989 ();
 sg13g2_decap_8 FILLER_53_2996 ();
 sg13g2_decap_8 FILLER_53_3003 ();
 sg13g2_decap_8 FILLER_53_3010 ();
 sg13g2_decap_8 FILLER_53_3017 ();
 sg13g2_decap_8 FILLER_53_3024 ();
 sg13g2_decap_8 FILLER_53_3031 ();
 sg13g2_decap_8 FILLER_53_3038 ();
 sg13g2_decap_8 FILLER_53_3045 ();
 sg13g2_decap_8 FILLER_53_3052 ();
 sg13g2_decap_8 FILLER_53_3059 ();
 sg13g2_decap_8 FILLER_53_3066 ();
 sg13g2_decap_8 FILLER_53_3073 ();
 sg13g2_decap_8 FILLER_53_3080 ();
 sg13g2_decap_8 FILLER_53_3087 ();
 sg13g2_decap_8 FILLER_53_3094 ();
 sg13g2_decap_8 FILLER_53_3101 ();
 sg13g2_decap_8 FILLER_53_3108 ();
 sg13g2_decap_8 FILLER_53_3115 ();
 sg13g2_decap_8 FILLER_53_3122 ();
 sg13g2_decap_8 FILLER_53_3129 ();
 sg13g2_decap_8 FILLER_53_3136 ();
 sg13g2_decap_8 FILLER_53_3143 ();
 sg13g2_decap_8 FILLER_53_3150 ();
 sg13g2_decap_8 FILLER_53_3157 ();
 sg13g2_decap_8 FILLER_53_3164 ();
 sg13g2_decap_8 FILLER_53_3171 ();
 sg13g2_decap_8 FILLER_53_3178 ();
 sg13g2_decap_8 FILLER_53_3185 ();
 sg13g2_decap_8 FILLER_53_3192 ();
 sg13g2_decap_8 FILLER_53_3199 ();
 sg13g2_decap_8 FILLER_53_3206 ();
 sg13g2_decap_8 FILLER_53_3213 ();
 sg13g2_decap_8 FILLER_53_3220 ();
 sg13g2_decap_8 FILLER_53_3227 ();
 sg13g2_decap_8 FILLER_53_3234 ();
 sg13g2_decap_8 FILLER_53_3241 ();
 sg13g2_decap_8 FILLER_53_3248 ();
 sg13g2_decap_8 FILLER_53_3255 ();
 sg13g2_decap_8 FILLER_53_3262 ();
 sg13g2_decap_8 FILLER_53_3269 ();
 sg13g2_decap_8 FILLER_53_3276 ();
 sg13g2_decap_8 FILLER_53_3283 ();
 sg13g2_decap_8 FILLER_53_3290 ();
 sg13g2_decap_8 FILLER_53_3297 ();
 sg13g2_decap_8 FILLER_53_3304 ();
 sg13g2_decap_8 FILLER_53_3311 ();
 sg13g2_decap_8 FILLER_53_3318 ();
 sg13g2_decap_8 FILLER_53_3325 ();
 sg13g2_decap_8 FILLER_53_3332 ();
 sg13g2_decap_8 FILLER_53_3339 ();
 sg13g2_decap_8 FILLER_53_3346 ();
 sg13g2_decap_8 FILLER_53_3353 ();
 sg13g2_decap_8 FILLER_53_3360 ();
 sg13g2_decap_8 FILLER_53_3367 ();
 sg13g2_decap_8 FILLER_53_3374 ();
 sg13g2_decap_8 FILLER_53_3381 ();
 sg13g2_decap_8 FILLER_53_3388 ();
 sg13g2_decap_8 FILLER_53_3395 ();
 sg13g2_decap_8 FILLER_53_3402 ();
 sg13g2_decap_8 FILLER_53_3409 ();
 sg13g2_decap_8 FILLER_53_3416 ();
 sg13g2_decap_8 FILLER_53_3423 ();
 sg13g2_decap_8 FILLER_53_3430 ();
 sg13g2_decap_8 FILLER_53_3437 ();
 sg13g2_decap_8 FILLER_53_3444 ();
 sg13g2_decap_8 FILLER_53_3451 ();
 sg13g2_decap_8 FILLER_53_3458 ();
 sg13g2_decap_8 FILLER_53_3465 ();
 sg13g2_decap_8 FILLER_53_3472 ();
 sg13g2_decap_8 FILLER_53_3479 ();
 sg13g2_decap_8 FILLER_53_3486 ();
 sg13g2_decap_8 FILLER_53_3493 ();
 sg13g2_decap_8 FILLER_53_3500 ();
 sg13g2_decap_8 FILLER_53_3507 ();
 sg13g2_decap_8 FILLER_53_3514 ();
 sg13g2_decap_8 FILLER_53_3521 ();
 sg13g2_decap_8 FILLER_53_3528 ();
 sg13g2_decap_8 FILLER_53_3535 ();
 sg13g2_decap_8 FILLER_53_3542 ();
 sg13g2_decap_8 FILLER_53_3549 ();
 sg13g2_decap_8 FILLER_53_3556 ();
 sg13g2_decap_8 FILLER_53_3563 ();
 sg13g2_decap_8 FILLER_53_3570 ();
 sg13g2_fill_2 FILLER_53_3577 ();
 sg13g2_fill_1 FILLER_53_3579 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_decap_8 FILLER_54_105 ();
 sg13g2_decap_8 FILLER_54_112 ();
 sg13g2_decap_8 FILLER_54_119 ();
 sg13g2_decap_8 FILLER_54_126 ();
 sg13g2_decap_8 FILLER_54_133 ();
 sg13g2_decap_8 FILLER_54_140 ();
 sg13g2_decap_8 FILLER_54_147 ();
 sg13g2_decap_8 FILLER_54_154 ();
 sg13g2_decap_8 FILLER_54_161 ();
 sg13g2_decap_8 FILLER_54_168 ();
 sg13g2_decap_8 FILLER_54_175 ();
 sg13g2_decap_8 FILLER_54_182 ();
 sg13g2_decap_8 FILLER_54_189 ();
 sg13g2_decap_8 FILLER_54_196 ();
 sg13g2_decap_8 FILLER_54_203 ();
 sg13g2_decap_8 FILLER_54_210 ();
 sg13g2_decap_8 FILLER_54_217 ();
 sg13g2_decap_8 FILLER_54_224 ();
 sg13g2_decap_8 FILLER_54_231 ();
 sg13g2_decap_8 FILLER_54_238 ();
 sg13g2_decap_8 FILLER_54_245 ();
 sg13g2_decap_8 FILLER_54_252 ();
 sg13g2_decap_8 FILLER_54_259 ();
 sg13g2_decap_8 FILLER_54_266 ();
 sg13g2_decap_8 FILLER_54_273 ();
 sg13g2_decap_8 FILLER_54_280 ();
 sg13g2_decap_8 FILLER_54_287 ();
 sg13g2_decap_8 FILLER_54_294 ();
 sg13g2_decap_8 FILLER_54_301 ();
 sg13g2_decap_8 FILLER_54_308 ();
 sg13g2_decap_8 FILLER_54_315 ();
 sg13g2_decap_8 FILLER_54_322 ();
 sg13g2_decap_8 FILLER_54_329 ();
 sg13g2_decap_8 FILLER_54_336 ();
 sg13g2_decap_8 FILLER_54_343 ();
 sg13g2_decap_8 FILLER_54_350 ();
 sg13g2_decap_8 FILLER_54_357 ();
 sg13g2_decap_8 FILLER_54_364 ();
 sg13g2_decap_8 FILLER_54_371 ();
 sg13g2_decap_8 FILLER_54_378 ();
 sg13g2_decap_8 FILLER_54_385 ();
 sg13g2_decap_8 FILLER_54_392 ();
 sg13g2_decap_8 FILLER_54_399 ();
 sg13g2_decap_8 FILLER_54_406 ();
 sg13g2_decap_8 FILLER_54_413 ();
 sg13g2_decap_8 FILLER_54_420 ();
 sg13g2_decap_8 FILLER_54_427 ();
 sg13g2_decap_8 FILLER_54_434 ();
 sg13g2_decap_8 FILLER_54_441 ();
 sg13g2_decap_8 FILLER_54_448 ();
 sg13g2_decap_8 FILLER_54_455 ();
 sg13g2_decap_8 FILLER_54_462 ();
 sg13g2_decap_8 FILLER_54_469 ();
 sg13g2_decap_8 FILLER_54_476 ();
 sg13g2_decap_8 FILLER_54_483 ();
 sg13g2_decap_8 FILLER_54_490 ();
 sg13g2_decap_8 FILLER_54_497 ();
 sg13g2_decap_8 FILLER_54_504 ();
 sg13g2_decap_8 FILLER_54_511 ();
 sg13g2_decap_8 FILLER_54_518 ();
 sg13g2_decap_8 FILLER_54_525 ();
 sg13g2_decap_8 FILLER_54_532 ();
 sg13g2_decap_8 FILLER_54_539 ();
 sg13g2_decap_8 FILLER_54_546 ();
 sg13g2_decap_8 FILLER_54_553 ();
 sg13g2_decap_8 FILLER_54_560 ();
 sg13g2_decap_8 FILLER_54_567 ();
 sg13g2_decap_8 FILLER_54_574 ();
 sg13g2_decap_8 FILLER_54_581 ();
 sg13g2_decap_8 FILLER_54_588 ();
 sg13g2_decap_8 FILLER_54_595 ();
 sg13g2_decap_8 FILLER_54_602 ();
 sg13g2_decap_8 FILLER_54_609 ();
 sg13g2_decap_8 FILLER_54_616 ();
 sg13g2_decap_8 FILLER_54_623 ();
 sg13g2_decap_8 FILLER_54_630 ();
 sg13g2_decap_8 FILLER_54_637 ();
 sg13g2_decap_8 FILLER_54_644 ();
 sg13g2_decap_8 FILLER_54_651 ();
 sg13g2_decap_8 FILLER_54_658 ();
 sg13g2_decap_8 FILLER_54_665 ();
 sg13g2_decap_8 FILLER_54_672 ();
 sg13g2_decap_8 FILLER_54_679 ();
 sg13g2_decap_8 FILLER_54_686 ();
 sg13g2_decap_8 FILLER_54_693 ();
 sg13g2_decap_8 FILLER_54_700 ();
 sg13g2_decap_8 FILLER_54_707 ();
 sg13g2_decap_8 FILLER_54_714 ();
 sg13g2_decap_8 FILLER_54_721 ();
 sg13g2_decap_8 FILLER_54_728 ();
 sg13g2_decap_8 FILLER_54_735 ();
 sg13g2_decap_8 FILLER_54_742 ();
 sg13g2_decap_8 FILLER_54_749 ();
 sg13g2_decap_8 FILLER_54_756 ();
 sg13g2_decap_8 FILLER_54_763 ();
 sg13g2_decap_8 FILLER_54_770 ();
 sg13g2_decap_8 FILLER_54_777 ();
 sg13g2_decap_8 FILLER_54_784 ();
 sg13g2_decap_8 FILLER_54_791 ();
 sg13g2_decap_8 FILLER_54_798 ();
 sg13g2_decap_8 FILLER_54_805 ();
 sg13g2_decap_8 FILLER_54_812 ();
 sg13g2_decap_8 FILLER_54_819 ();
 sg13g2_decap_8 FILLER_54_826 ();
 sg13g2_decap_8 FILLER_54_833 ();
 sg13g2_decap_8 FILLER_54_840 ();
 sg13g2_decap_8 FILLER_54_847 ();
 sg13g2_decap_8 FILLER_54_854 ();
 sg13g2_decap_8 FILLER_54_861 ();
 sg13g2_decap_8 FILLER_54_868 ();
 sg13g2_decap_8 FILLER_54_875 ();
 sg13g2_decap_8 FILLER_54_882 ();
 sg13g2_decap_8 FILLER_54_889 ();
 sg13g2_decap_8 FILLER_54_896 ();
 sg13g2_decap_8 FILLER_54_903 ();
 sg13g2_decap_8 FILLER_54_910 ();
 sg13g2_decap_8 FILLER_54_917 ();
 sg13g2_decap_8 FILLER_54_924 ();
 sg13g2_decap_8 FILLER_54_931 ();
 sg13g2_decap_8 FILLER_54_938 ();
 sg13g2_decap_8 FILLER_54_945 ();
 sg13g2_decap_8 FILLER_54_952 ();
 sg13g2_decap_8 FILLER_54_959 ();
 sg13g2_decap_8 FILLER_54_966 ();
 sg13g2_decap_8 FILLER_54_973 ();
 sg13g2_decap_8 FILLER_54_980 ();
 sg13g2_decap_8 FILLER_54_987 ();
 sg13g2_decap_8 FILLER_54_994 ();
 sg13g2_decap_8 FILLER_54_1001 ();
 sg13g2_decap_8 FILLER_54_1008 ();
 sg13g2_decap_8 FILLER_54_1015 ();
 sg13g2_decap_8 FILLER_54_1022 ();
 sg13g2_decap_8 FILLER_54_1029 ();
 sg13g2_decap_8 FILLER_54_1036 ();
 sg13g2_decap_8 FILLER_54_1043 ();
 sg13g2_decap_8 FILLER_54_1050 ();
 sg13g2_decap_8 FILLER_54_1057 ();
 sg13g2_decap_8 FILLER_54_1064 ();
 sg13g2_decap_8 FILLER_54_1071 ();
 sg13g2_decap_8 FILLER_54_1078 ();
 sg13g2_decap_8 FILLER_54_1085 ();
 sg13g2_decap_8 FILLER_54_1092 ();
 sg13g2_decap_8 FILLER_54_1099 ();
 sg13g2_decap_8 FILLER_54_1106 ();
 sg13g2_decap_8 FILLER_54_1113 ();
 sg13g2_decap_8 FILLER_54_1120 ();
 sg13g2_decap_8 FILLER_54_1127 ();
 sg13g2_decap_8 FILLER_54_1134 ();
 sg13g2_decap_8 FILLER_54_1141 ();
 sg13g2_decap_8 FILLER_54_1148 ();
 sg13g2_decap_8 FILLER_54_1155 ();
 sg13g2_decap_8 FILLER_54_1162 ();
 sg13g2_decap_8 FILLER_54_1169 ();
 sg13g2_decap_8 FILLER_54_1176 ();
 sg13g2_decap_8 FILLER_54_1183 ();
 sg13g2_decap_8 FILLER_54_1190 ();
 sg13g2_decap_8 FILLER_54_1197 ();
 sg13g2_decap_8 FILLER_54_1204 ();
 sg13g2_decap_8 FILLER_54_1211 ();
 sg13g2_decap_8 FILLER_54_1218 ();
 sg13g2_decap_8 FILLER_54_1225 ();
 sg13g2_decap_8 FILLER_54_1232 ();
 sg13g2_decap_8 FILLER_54_1239 ();
 sg13g2_decap_8 FILLER_54_1246 ();
 sg13g2_decap_8 FILLER_54_1253 ();
 sg13g2_decap_8 FILLER_54_1260 ();
 sg13g2_decap_8 FILLER_54_1267 ();
 sg13g2_decap_8 FILLER_54_1274 ();
 sg13g2_decap_8 FILLER_54_1281 ();
 sg13g2_decap_8 FILLER_54_1288 ();
 sg13g2_decap_8 FILLER_54_1295 ();
 sg13g2_decap_8 FILLER_54_1302 ();
 sg13g2_decap_8 FILLER_54_1309 ();
 sg13g2_decap_8 FILLER_54_1316 ();
 sg13g2_decap_8 FILLER_54_1323 ();
 sg13g2_decap_8 FILLER_54_1330 ();
 sg13g2_decap_8 FILLER_54_1337 ();
 sg13g2_decap_8 FILLER_54_1344 ();
 sg13g2_decap_8 FILLER_54_1351 ();
 sg13g2_decap_8 FILLER_54_1358 ();
 sg13g2_decap_8 FILLER_54_1365 ();
 sg13g2_decap_8 FILLER_54_1372 ();
 sg13g2_decap_8 FILLER_54_1379 ();
 sg13g2_decap_8 FILLER_54_1386 ();
 sg13g2_decap_8 FILLER_54_1393 ();
 sg13g2_decap_8 FILLER_54_1400 ();
 sg13g2_decap_8 FILLER_54_1407 ();
 sg13g2_decap_8 FILLER_54_1414 ();
 sg13g2_decap_8 FILLER_54_1421 ();
 sg13g2_decap_8 FILLER_54_1428 ();
 sg13g2_decap_8 FILLER_54_1435 ();
 sg13g2_decap_8 FILLER_54_1442 ();
 sg13g2_decap_8 FILLER_54_1449 ();
 sg13g2_decap_8 FILLER_54_1456 ();
 sg13g2_decap_8 FILLER_54_1463 ();
 sg13g2_decap_8 FILLER_54_1470 ();
 sg13g2_decap_8 FILLER_54_1477 ();
 sg13g2_decap_8 FILLER_54_1484 ();
 sg13g2_decap_8 FILLER_54_1491 ();
 sg13g2_decap_8 FILLER_54_1498 ();
 sg13g2_decap_8 FILLER_54_1505 ();
 sg13g2_decap_8 FILLER_54_1512 ();
 sg13g2_decap_8 FILLER_54_1519 ();
 sg13g2_decap_8 FILLER_54_1526 ();
 sg13g2_decap_8 FILLER_54_1533 ();
 sg13g2_decap_8 FILLER_54_1540 ();
 sg13g2_decap_8 FILLER_54_1547 ();
 sg13g2_decap_8 FILLER_54_1554 ();
 sg13g2_decap_8 FILLER_54_1561 ();
 sg13g2_decap_8 FILLER_54_1568 ();
 sg13g2_decap_8 FILLER_54_1575 ();
 sg13g2_decap_8 FILLER_54_1582 ();
 sg13g2_decap_8 FILLER_54_1589 ();
 sg13g2_decap_8 FILLER_54_1596 ();
 sg13g2_decap_8 FILLER_54_1603 ();
 sg13g2_decap_8 FILLER_54_1610 ();
 sg13g2_decap_8 FILLER_54_1617 ();
 sg13g2_decap_8 FILLER_54_1624 ();
 sg13g2_decap_8 FILLER_54_1631 ();
 sg13g2_decap_8 FILLER_54_1638 ();
 sg13g2_decap_8 FILLER_54_1645 ();
 sg13g2_decap_8 FILLER_54_1652 ();
 sg13g2_decap_8 FILLER_54_1659 ();
 sg13g2_decap_8 FILLER_54_1666 ();
 sg13g2_decap_8 FILLER_54_1673 ();
 sg13g2_decap_8 FILLER_54_1680 ();
 sg13g2_decap_8 FILLER_54_1687 ();
 sg13g2_decap_8 FILLER_54_1694 ();
 sg13g2_decap_8 FILLER_54_1701 ();
 sg13g2_decap_8 FILLER_54_1708 ();
 sg13g2_decap_8 FILLER_54_1715 ();
 sg13g2_decap_8 FILLER_54_1722 ();
 sg13g2_decap_8 FILLER_54_1729 ();
 sg13g2_decap_8 FILLER_54_1736 ();
 sg13g2_decap_8 FILLER_54_1743 ();
 sg13g2_decap_8 FILLER_54_1750 ();
 sg13g2_decap_8 FILLER_54_1757 ();
 sg13g2_decap_8 FILLER_54_1764 ();
 sg13g2_decap_8 FILLER_54_1771 ();
 sg13g2_decap_8 FILLER_54_1778 ();
 sg13g2_decap_8 FILLER_54_1785 ();
 sg13g2_decap_8 FILLER_54_1792 ();
 sg13g2_decap_8 FILLER_54_1799 ();
 sg13g2_decap_8 FILLER_54_1806 ();
 sg13g2_decap_8 FILLER_54_1813 ();
 sg13g2_decap_8 FILLER_54_1820 ();
 sg13g2_decap_8 FILLER_54_1827 ();
 sg13g2_decap_8 FILLER_54_1834 ();
 sg13g2_decap_8 FILLER_54_1841 ();
 sg13g2_decap_8 FILLER_54_1848 ();
 sg13g2_decap_8 FILLER_54_1855 ();
 sg13g2_decap_8 FILLER_54_1862 ();
 sg13g2_decap_8 FILLER_54_1869 ();
 sg13g2_decap_8 FILLER_54_1876 ();
 sg13g2_decap_8 FILLER_54_1883 ();
 sg13g2_decap_8 FILLER_54_1890 ();
 sg13g2_decap_8 FILLER_54_1897 ();
 sg13g2_decap_8 FILLER_54_1904 ();
 sg13g2_decap_8 FILLER_54_1911 ();
 sg13g2_decap_8 FILLER_54_1918 ();
 sg13g2_decap_8 FILLER_54_1925 ();
 sg13g2_decap_8 FILLER_54_1932 ();
 sg13g2_decap_8 FILLER_54_1939 ();
 sg13g2_decap_8 FILLER_54_1946 ();
 sg13g2_decap_8 FILLER_54_1953 ();
 sg13g2_decap_8 FILLER_54_1960 ();
 sg13g2_decap_8 FILLER_54_1967 ();
 sg13g2_decap_8 FILLER_54_1974 ();
 sg13g2_decap_8 FILLER_54_1981 ();
 sg13g2_decap_8 FILLER_54_1988 ();
 sg13g2_decap_8 FILLER_54_1995 ();
 sg13g2_decap_8 FILLER_54_2002 ();
 sg13g2_decap_8 FILLER_54_2009 ();
 sg13g2_decap_8 FILLER_54_2016 ();
 sg13g2_decap_8 FILLER_54_2023 ();
 sg13g2_decap_8 FILLER_54_2030 ();
 sg13g2_decap_8 FILLER_54_2037 ();
 sg13g2_decap_8 FILLER_54_2044 ();
 sg13g2_decap_8 FILLER_54_2051 ();
 sg13g2_decap_8 FILLER_54_2058 ();
 sg13g2_decap_8 FILLER_54_2065 ();
 sg13g2_decap_8 FILLER_54_2072 ();
 sg13g2_decap_8 FILLER_54_2079 ();
 sg13g2_decap_8 FILLER_54_2086 ();
 sg13g2_decap_8 FILLER_54_2093 ();
 sg13g2_decap_8 FILLER_54_2100 ();
 sg13g2_decap_8 FILLER_54_2107 ();
 sg13g2_decap_8 FILLER_54_2114 ();
 sg13g2_decap_8 FILLER_54_2121 ();
 sg13g2_decap_8 FILLER_54_2128 ();
 sg13g2_decap_8 FILLER_54_2135 ();
 sg13g2_decap_8 FILLER_54_2142 ();
 sg13g2_decap_8 FILLER_54_2149 ();
 sg13g2_decap_8 FILLER_54_2156 ();
 sg13g2_decap_8 FILLER_54_2163 ();
 sg13g2_decap_8 FILLER_54_2170 ();
 sg13g2_decap_8 FILLER_54_2177 ();
 sg13g2_decap_8 FILLER_54_2184 ();
 sg13g2_decap_8 FILLER_54_2191 ();
 sg13g2_decap_8 FILLER_54_2198 ();
 sg13g2_decap_8 FILLER_54_2205 ();
 sg13g2_decap_8 FILLER_54_2212 ();
 sg13g2_decap_8 FILLER_54_2219 ();
 sg13g2_decap_8 FILLER_54_2226 ();
 sg13g2_decap_8 FILLER_54_2233 ();
 sg13g2_decap_8 FILLER_54_2240 ();
 sg13g2_decap_8 FILLER_54_2247 ();
 sg13g2_decap_8 FILLER_54_2254 ();
 sg13g2_decap_8 FILLER_54_2261 ();
 sg13g2_decap_8 FILLER_54_2268 ();
 sg13g2_decap_8 FILLER_54_2275 ();
 sg13g2_decap_8 FILLER_54_2282 ();
 sg13g2_decap_8 FILLER_54_2289 ();
 sg13g2_decap_8 FILLER_54_2296 ();
 sg13g2_decap_8 FILLER_54_2303 ();
 sg13g2_decap_8 FILLER_54_2310 ();
 sg13g2_decap_8 FILLER_54_2317 ();
 sg13g2_decap_8 FILLER_54_2324 ();
 sg13g2_decap_8 FILLER_54_2331 ();
 sg13g2_decap_8 FILLER_54_2338 ();
 sg13g2_decap_8 FILLER_54_2345 ();
 sg13g2_decap_8 FILLER_54_2352 ();
 sg13g2_decap_8 FILLER_54_2359 ();
 sg13g2_decap_8 FILLER_54_2366 ();
 sg13g2_decap_8 FILLER_54_2373 ();
 sg13g2_decap_8 FILLER_54_2380 ();
 sg13g2_decap_8 FILLER_54_2387 ();
 sg13g2_decap_8 FILLER_54_2394 ();
 sg13g2_decap_8 FILLER_54_2401 ();
 sg13g2_decap_8 FILLER_54_2408 ();
 sg13g2_decap_8 FILLER_54_2415 ();
 sg13g2_decap_8 FILLER_54_2422 ();
 sg13g2_decap_8 FILLER_54_2429 ();
 sg13g2_decap_8 FILLER_54_2436 ();
 sg13g2_decap_8 FILLER_54_2443 ();
 sg13g2_decap_8 FILLER_54_2450 ();
 sg13g2_decap_8 FILLER_54_2457 ();
 sg13g2_decap_8 FILLER_54_2464 ();
 sg13g2_decap_8 FILLER_54_2471 ();
 sg13g2_decap_8 FILLER_54_2478 ();
 sg13g2_decap_8 FILLER_54_2485 ();
 sg13g2_decap_8 FILLER_54_2492 ();
 sg13g2_decap_8 FILLER_54_2499 ();
 sg13g2_decap_8 FILLER_54_2506 ();
 sg13g2_decap_8 FILLER_54_2513 ();
 sg13g2_decap_8 FILLER_54_2520 ();
 sg13g2_decap_8 FILLER_54_2527 ();
 sg13g2_decap_8 FILLER_54_2534 ();
 sg13g2_decap_8 FILLER_54_2541 ();
 sg13g2_decap_8 FILLER_54_2548 ();
 sg13g2_decap_8 FILLER_54_2555 ();
 sg13g2_decap_8 FILLER_54_2562 ();
 sg13g2_decap_8 FILLER_54_2569 ();
 sg13g2_decap_8 FILLER_54_2576 ();
 sg13g2_decap_8 FILLER_54_2583 ();
 sg13g2_decap_8 FILLER_54_2590 ();
 sg13g2_decap_8 FILLER_54_2597 ();
 sg13g2_decap_8 FILLER_54_2604 ();
 sg13g2_decap_8 FILLER_54_2611 ();
 sg13g2_decap_8 FILLER_54_2618 ();
 sg13g2_decap_8 FILLER_54_2625 ();
 sg13g2_decap_8 FILLER_54_2632 ();
 sg13g2_decap_8 FILLER_54_2639 ();
 sg13g2_decap_8 FILLER_54_2646 ();
 sg13g2_decap_8 FILLER_54_2653 ();
 sg13g2_decap_8 FILLER_54_2660 ();
 sg13g2_decap_8 FILLER_54_2667 ();
 sg13g2_decap_8 FILLER_54_2674 ();
 sg13g2_decap_8 FILLER_54_2681 ();
 sg13g2_decap_8 FILLER_54_2688 ();
 sg13g2_decap_8 FILLER_54_2695 ();
 sg13g2_decap_8 FILLER_54_2702 ();
 sg13g2_decap_8 FILLER_54_2709 ();
 sg13g2_decap_8 FILLER_54_2716 ();
 sg13g2_decap_8 FILLER_54_2723 ();
 sg13g2_decap_8 FILLER_54_2730 ();
 sg13g2_decap_8 FILLER_54_2737 ();
 sg13g2_decap_8 FILLER_54_2744 ();
 sg13g2_decap_8 FILLER_54_2751 ();
 sg13g2_decap_8 FILLER_54_2758 ();
 sg13g2_decap_8 FILLER_54_2765 ();
 sg13g2_decap_8 FILLER_54_2772 ();
 sg13g2_decap_8 FILLER_54_2779 ();
 sg13g2_decap_8 FILLER_54_2786 ();
 sg13g2_decap_8 FILLER_54_2793 ();
 sg13g2_decap_8 FILLER_54_2800 ();
 sg13g2_decap_8 FILLER_54_2807 ();
 sg13g2_decap_8 FILLER_54_2814 ();
 sg13g2_decap_8 FILLER_54_2821 ();
 sg13g2_decap_8 FILLER_54_2828 ();
 sg13g2_decap_8 FILLER_54_2835 ();
 sg13g2_decap_8 FILLER_54_2842 ();
 sg13g2_decap_8 FILLER_54_2849 ();
 sg13g2_decap_8 FILLER_54_2856 ();
 sg13g2_decap_8 FILLER_54_2863 ();
 sg13g2_decap_8 FILLER_54_2870 ();
 sg13g2_decap_8 FILLER_54_2877 ();
 sg13g2_decap_8 FILLER_54_2884 ();
 sg13g2_decap_8 FILLER_54_2891 ();
 sg13g2_decap_8 FILLER_54_2898 ();
 sg13g2_decap_8 FILLER_54_2905 ();
 sg13g2_decap_8 FILLER_54_2912 ();
 sg13g2_decap_8 FILLER_54_2919 ();
 sg13g2_decap_8 FILLER_54_2926 ();
 sg13g2_decap_8 FILLER_54_2933 ();
 sg13g2_decap_8 FILLER_54_2940 ();
 sg13g2_decap_8 FILLER_54_2947 ();
 sg13g2_decap_8 FILLER_54_2954 ();
 sg13g2_decap_8 FILLER_54_2961 ();
 sg13g2_decap_8 FILLER_54_2968 ();
 sg13g2_decap_8 FILLER_54_2975 ();
 sg13g2_decap_8 FILLER_54_2982 ();
 sg13g2_decap_8 FILLER_54_2989 ();
 sg13g2_decap_8 FILLER_54_2996 ();
 sg13g2_decap_8 FILLER_54_3003 ();
 sg13g2_decap_8 FILLER_54_3010 ();
 sg13g2_decap_8 FILLER_54_3017 ();
 sg13g2_decap_8 FILLER_54_3024 ();
 sg13g2_decap_8 FILLER_54_3031 ();
 sg13g2_decap_8 FILLER_54_3038 ();
 sg13g2_decap_8 FILLER_54_3045 ();
 sg13g2_decap_8 FILLER_54_3052 ();
 sg13g2_decap_8 FILLER_54_3059 ();
 sg13g2_decap_8 FILLER_54_3066 ();
 sg13g2_decap_8 FILLER_54_3073 ();
 sg13g2_decap_8 FILLER_54_3080 ();
 sg13g2_decap_8 FILLER_54_3087 ();
 sg13g2_decap_8 FILLER_54_3094 ();
 sg13g2_decap_8 FILLER_54_3101 ();
 sg13g2_decap_8 FILLER_54_3108 ();
 sg13g2_decap_8 FILLER_54_3115 ();
 sg13g2_decap_8 FILLER_54_3122 ();
 sg13g2_decap_8 FILLER_54_3129 ();
 sg13g2_decap_8 FILLER_54_3136 ();
 sg13g2_decap_8 FILLER_54_3143 ();
 sg13g2_decap_8 FILLER_54_3150 ();
 sg13g2_decap_8 FILLER_54_3157 ();
 sg13g2_decap_8 FILLER_54_3164 ();
 sg13g2_decap_8 FILLER_54_3171 ();
 sg13g2_decap_8 FILLER_54_3178 ();
 sg13g2_decap_8 FILLER_54_3185 ();
 sg13g2_decap_8 FILLER_54_3192 ();
 sg13g2_decap_8 FILLER_54_3199 ();
 sg13g2_decap_8 FILLER_54_3206 ();
 sg13g2_decap_8 FILLER_54_3213 ();
 sg13g2_decap_8 FILLER_54_3220 ();
 sg13g2_decap_8 FILLER_54_3227 ();
 sg13g2_decap_8 FILLER_54_3234 ();
 sg13g2_decap_8 FILLER_54_3241 ();
 sg13g2_decap_8 FILLER_54_3248 ();
 sg13g2_decap_8 FILLER_54_3255 ();
 sg13g2_decap_8 FILLER_54_3262 ();
 sg13g2_decap_8 FILLER_54_3269 ();
 sg13g2_decap_8 FILLER_54_3276 ();
 sg13g2_decap_8 FILLER_54_3283 ();
 sg13g2_decap_8 FILLER_54_3290 ();
 sg13g2_decap_8 FILLER_54_3297 ();
 sg13g2_decap_8 FILLER_54_3304 ();
 sg13g2_decap_8 FILLER_54_3311 ();
 sg13g2_decap_8 FILLER_54_3318 ();
 sg13g2_decap_8 FILLER_54_3325 ();
 sg13g2_decap_8 FILLER_54_3332 ();
 sg13g2_decap_8 FILLER_54_3339 ();
 sg13g2_decap_8 FILLER_54_3346 ();
 sg13g2_decap_8 FILLER_54_3353 ();
 sg13g2_decap_8 FILLER_54_3360 ();
 sg13g2_decap_8 FILLER_54_3367 ();
 sg13g2_decap_8 FILLER_54_3374 ();
 sg13g2_decap_8 FILLER_54_3381 ();
 sg13g2_decap_8 FILLER_54_3388 ();
 sg13g2_decap_8 FILLER_54_3395 ();
 sg13g2_decap_8 FILLER_54_3402 ();
 sg13g2_decap_8 FILLER_54_3409 ();
 sg13g2_decap_8 FILLER_54_3416 ();
 sg13g2_decap_8 FILLER_54_3423 ();
 sg13g2_decap_8 FILLER_54_3430 ();
 sg13g2_decap_8 FILLER_54_3437 ();
 sg13g2_decap_8 FILLER_54_3444 ();
 sg13g2_decap_8 FILLER_54_3451 ();
 sg13g2_decap_8 FILLER_54_3458 ();
 sg13g2_decap_8 FILLER_54_3465 ();
 sg13g2_decap_8 FILLER_54_3472 ();
 sg13g2_decap_8 FILLER_54_3479 ();
 sg13g2_decap_8 FILLER_54_3486 ();
 sg13g2_decap_8 FILLER_54_3493 ();
 sg13g2_decap_8 FILLER_54_3500 ();
 sg13g2_decap_8 FILLER_54_3507 ();
 sg13g2_decap_8 FILLER_54_3514 ();
 sg13g2_decap_8 FILLER_54_3521 ();
 sg13g2_decap_8 FILLER_54_3528 ();
 sg13g2_decap_8 FILLER_54_3535 ();
 sg13g2_decap_8 FILLER_54_3542 ();
 sg13g2_decap_8 FILLER_54_3549 ();
 sg13g2_decap_8 FILLER_54_3556 ();
 sg13g2_decap_8 FILLER_54_3563 ();
 sg13g2_decap_8 FILLER_54_3570 ();
 sg13g2_fill_2 FILLER_54_3577 ();
 sg13g2_fill_1 FILLER_54_3579 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_98 ();
 sg13g2_decap_8 FILLER_55_105 ();
 sg13g2_decap_8 FILLER_55_112 ();
 sg13g2_decap_8 FILLER_55_119 ();
 sg13g2_decap_8 FILLER_55_126 ();
 sg13g2_decap_8 FILLER_55_133 ();
 sg13g2_decap_8 FILLER_55_140 ();
 sg13g2_decap_8 FILLER_55_147 ();
 sg13g2_decap_8 FILLER_55_154 ();
 sg13g2_decap_8 FILLER_55_161 ();
 sg13g2_decap_8 FILLER_55_168 ();
 sg13g2_decap_8 FILLER_55_175 ();
 sg13g2_decap_8 FILLER_55_182 ();
 sg13g2_decap_8 FILLER_55_189 ();
 sg13g2_decap_8 FILLER_55_196 ();
 sg13g2_decap_8 FILLER_55_203 ();
 sg13g2_decap_8 FILLER_55_210 ();
 sg13g2_decap_8 FILLER_55_217 ();
 sg13g2_decap_8 FILLER_55_224 ();
 sg13g2_decap_8 FILLER_55_231 ();
 sg13g2_decap_8 FILLER_55_238 ();
 sg13g2_decap_8 FILLER_55_245 ();
 sg13g2_decap_8 FILLER_55_252 ();
 sg13g2_decap_8 FILLER_55_259 ();
 sg13g2_decap_8 FILLER_55_266 ();
 sg13g2_decap_8 FILLER_55_273 ();
 sg13g2_decap_8 FILLER_55_280 ();
 sg13g2_decap_8 FILLER_55_287 ();
 sg13g2_decap_8 FILLER_55_294 ();
 sg13g2_decap_8 FILLER_55_301 ();
 sg13g2_decap_8 FILLER_55_308 ();
 sg13g2_decap_8 FILLER_55_315 ();
 sg13g2_decap_8 FILLER_55_322 ();
 sg13g2_decap_8 FILLER_55_329 ();
 sg13g2_decap_8 FILLER_55_336 ();
 sg13g2_decap_8 FILLER_55_343 ();
 sg13g2_decap_8 FILLER_55_350 ();
 sg13g2_decap_8 FILLER_55_357 ();
 sg13g2_decap_8 FILLER_55_364 ();
 sg13g2_decap_8 FILLER_55_371 ();
 sg13g2_decap_8 FILLER_55_378 ();
 sg13g2_decap_8 FILLER_55_385 ();
 sg13g2_decap_8 FILLER_55_392 ();
 sg13g2_decap_8 FILLER_55_399 ();
 sg13g2_decap_8 FILLER_55_406 ();
 sg13g2_decap_8 FILLER_55_413 ();
 sg13g2_decap_8 FILLER_55_420 ();
 sg13g2_decap_8 FILLER_55_427 ();
 sg13g2_decap_8 FILLER_55_434 ();
 sg13g2_decap_8 FILLER_55_441 ();
 sg13g2_decap_8 FILLER_55_448 ();
 sg13g2_decap_8 FILLER_55_455 ();
 sg13g2_decap_8 FILLER_55_462 ();
 sg13g2_decap_8 FILLER_55_469 ();
 sg13g2_decap_8 FILLER_55_476 ();
 sg13g2_decap_8 FILLER_55_483 ();
 sg13g2_decap_8 FILLER_55_490 ();
 sg13g2_decap_8 FILLER_55_497 ();
 sg13g2_decap_8 FILLER_55_504 ();
 sg13g2_decap_8 FILLER_55_511 ();
 sg13g2_decap_8 FILLER_55_518 ();
 sg13g2_decap_8 FILLER_55_525 ();
 sg13g2_decap_8 FILLER_55_532 ();
 sg13g2_decap_8 FILLER_55_539 ();
 sg13g2_decap_8 FILLER_55_546 ();
 sg13g2_decap_8 FILLER_55_553 ();
 sg13g2_decap_8 FILLER_55_560 ();
 sg13g2_decap_8 FILLER_55_567 ();
 sg13g2_decap_8 FILLER_55_574 ();
 sg13g2_decap_8 FILLER_55_581 ();
 sg13g2_decap_8 FILLER_55_588 ();
 sg13g2_decap_8 FILLER_55_595 ();
 sg13g2_decap_8 FILLER_55_602 ();
 sg13g2_decap_8 FILLER_55_609 ();
 sg13g2_decap_8 FILLER_55_616 ();
 sg13g2_decap_8 FILLER_55_623 ();
 sg13g2_decap_8 FILLER_55_630 ();
 sg13g2_decap_8 FILLER_55_637 ();
 sg13g2_decap_8 FILLER_55_644 ();
 sg13g2_decap_8 FILLER_55_651 ();
 sg13g2_decap_8 FILLER_55_658 ();
 sg13g2_decap_8 FILLER_55_665 ();
 sg13g2_decap_8 FILLER_55_672 ();
 sg13g2_decap_8 FILLER_55_679 ();
 sg13g2_decap_8 FILLER_55_686 ();
 sg13g2_decap_8 FILLER_55_693 ();
 sg13g2_decap_8 FILLER_55_700 ();
 sg13g2_decap_8 FILLER_55_707 ();
 sg13g2_decap_8 FILLER_55_714 ();
 sg13g2_decap_8 FILLER_55_721 ();
 sg13g2_decap_8 FILLER_55_728 ();
 sg13g2_decap_8 FILLER_55_735 ();
 sg13g2_decap_8 FILLER_55_742 ();
 sg13g2_decap_8 FILLER_55_749 ();
 sg13g2_decap_8 FILLER_55_756 ();
 sg13g2_decap_8 FILLER_55_763 ();
 sg13g2_decap_8 FILLER_55_770 ();
 sg13g2_decap_8 FILLER_55_777 ();
 sg13g2_decap_8 FILLER_55_784 ();
 sg13g2_decap_8 FILLER_55_791 ();
 sg13g2_decap_8 FILLER_55_798 ();
 sg13g2_decap_8 FILLER_55_805 ();
 sg13g2_decap_8 FILLER_55_812 ();
 sg13g2_decap_8 FILLER_55_819 ();
 sg13g2_decap_8 FILLER_55_826 ();
 sg13g2_decap_8 FILLER_55_833 ();
 sg13g2_decap_8 FILLER_55_840 ();
 sg13g2_decap_8 FILLER_55_847 ();
 sg13g2_decap_8 FILLER_55_854 ();
 sg13g2_decap_8 FILLER_55_861 ();
 sg13g2_decap_8 FILLER_55_868 ();
 sg13g2_decap_8 FILLER_55_875 ();
 sg13g2_decap_8 FILLER_55_882 ();
 sg13g2_decap_8 FILLER_55_889 ();
 sg13g2_decap_8 FILLER_55_896 ();
 sg13g2_decap_8 FILLER_55_903 ();
 sg13g2_decap_8 FILLER_55_910 ();
 sg13g2_decap_8 FILLER_55_917 ();
 sg13g2_decap_8 FILLER_55_924 ();
 sg13g2_decap_8 FILLER_55_931 ();
 sg13g2_decap_8 FILLER_55_938 ();
 sg13g2_decap_8 FILLER_55_945 ();
 sg13g2_decap_8 FILLER_55_952 ();
 sg13g2_decap_8 FILLER_55_959 ();
 sg13g2_decap_8 FILLER_55_966 ();
 sg13g2_decap_8 FILLER_55_973 ();
 sg13g2_decap_8 FILLER_55_980 ();
 sg13g2_decap_8 FILLER_55_987 ();
 sg13g2_decap_8 FILLER_55_994 ();
 sg13g2_decap_8 FILLER_55_1001 ();
 sg13g2_decap_8 FILLER_55_1008 ();
 sg13g2_decap_8 FILLER_55_1015 ();
 sg13g2_decap_8 FILLER_55_1022 ();
 sg13g2_decap_8 FILLER_55_1029 ();
 sg13g2_decap_8 FILLER_55_1036 ();
 sg13g2_decap_8 FILLER_55_1043 ();
 sg13g2_decap_8 FILLER_55_1050 ();
 sg13g2_decap_8 FILLER_55_1057 ();
 sg13g2_decap_8 FILLER_55_1064 ();
 sg13g2_decap_8 FILLER_55_1071 ();
 sg13g2_decap_8 FILLER_55_1078 ();
 sg13g2_decap_8 FILLER_55_1085 ();
 sg13g2_decap_8 FILLER_55_1092 ();
 sg13g2_decap_8 FILLER_55_1099 ();
 sg13g2_decap_8 FILLER_55_1106 ();
 sg13g2_decap_8 FILLER_55_1113 ();
 sg13g2_decap_8 FILLER_55_1120 ();
 sg13g2_decap_8 FILLER_55_1127 ();
 sg13g2_decap_8 FILLER_55_1134 ();
 sg13g2_decap_8 FILLER_55_1141 ();
 sg13g2_decap_8 FILLER_55_1148 ();
 sg13g2_decap_8 FILLER_55_1155 ();
 sg13g2_decap_8 FILLER_55_1162 ();
 sg13g2_decap_8 FILLER_55_1169 ();
 sg13g2_decap_8 FILLER_55_1176 ();
 sg13g2_decap_8 FILLER_55_1183 ();
 sg13g2_decap_8 FILLER_55_1190 ();
 sg13g2_decap_8 FILLER_55_1197 ();
 sg13g2_decap_8 FILLER_55_1204 ();
 sg13g2_decap_8 FILLER_55_1211 ();
 sg13g2_decap_8 FILLER_55_1218 ();
 sg13g2_decap_8 FILLER_55_1225 ();
 sg13g2_decap_8 FILLER_55_1232 ();
 sg13g2_decap_8 FILLER_55_1239 ();
 sg13g2_decap_8 FILLER_55_1246 ();
 sg13g2_decap_8 FILLER_55_1253 ();
 sg13g2_decap_8 FILLER_55_1260 ();
 sg13g2_decap_8 FILLER_55_1267 ();
 sg13g2_decap_8 FILLER_55_1274 ();
 sg13g2_decap_8 FILLER_55_1281 ();
 sg13g2_decap_8 FILLER_55_1288 ();
 sg13g2_decap_8 FILLER_55_1295 ();
 sg13g2_decap_8 FILLER_55_1302 ();
 sg13g2_decap_8 FILLER_55_1309 ();
 sg13g2_decap_8 FILLER_55_1316 ();
 sg13g2_decap_8 FILLER_55_1323 ();
 sg13g2_decap_8 FILLER_55_1330 ();
 sg13g2_decap_8 FILLER_55_1337 ();
 sg13g2_decap_8 FILLER_55_1344 ();
 sg13g2_decap_8 FILLER_55_1351 ();
 sg13g2_decap_8 FILLER_55_1358 ();
 sg13g2_decap_8 FILLER_55_1365 ();
 sg13g2_decap_8 FILLER_55_1372 ();
 sg13g2_decap_8 FILLER_55_1379 ();
 sg13g2_decap_8 FILLER_55_1386 ();
 sg13g2_decap_8 FILLER_55_1393 ();
 sg13g2_decap_8 FILLER_55_1400 ();
 sg13g2_decap_8 FILLER_55_1407 ();
 sg13g2_decap_8 FILLER_55_1414 ();
 sg13g2_decap_8 FILLER_55_1421 ();
 sg13g2_decap_8 FILLER_55_1428 ();
 sg13g2_decap_8 FILLER_55_1435 ();
 sg13g2_decap_8 FILLER_55_1442 ();
 sg13g2_decap_8 FILLER_55_1449 ();
 sg13g2_decap_8 FILLER_55_1456 ();
 sg13g2_decap_8 FILLER_55_1463 ();
 sg13g2_decap_8 FILLER_55_1470 ();
 sg13g2_decap_8 FILLER_55_1477 ();
 sg13g2_decap_8 FILLER_55_1484 ();
 sg13g2_decap_8 FILLER_55_1491 ();
 sg13g2_decap_8 FILLER_55_1498 ();
 sg13g2_decap_8 FILLER_55_1505 ();
 sg13g2_decap_8 FILLER_55_1512 ();
 sg13g2_decap_8 FILLER_55_1519 ();
 sg13g2_decap_8 FILLER_55_1526 ();
 sg13g2_decap_8 FILLER_55_1533 ();
 sg13g2_decap_8 FILLER_55_1540 ();
 sg13g2_decap_8 FILLER_55_1547 ();
 sg13g2_decap_8 FILLER_55_1554 ();
 sg13g2_decap_8 FILLER_55_1561 ();
 sg13g2_decap_8 FILLER_55_1568 ();
 sg13g2_decap_8 FILLER_55_1575 ();
 sg13g2_decap_8 FILLER_55_1582 ();
 sg13g2_decap_8 FILLER_55_1589 ();
 sg13g2_decap_8 FILLER_55_1596 ();
 sg13g2_decap_8 FILLER_55_1603 ();
 sg13g2_decap_8 FILLER_55_1610 ();
 sg13g2_decap_8 FILLER_55_1617 ();
 sg13g2_decap_8 FILLER_55_1624 ();
 sg13g2_decap_8 FILLER_55_1631 ();
 sg13g2_decap_8 FILLER_55_1638 ();
 sg13g2_decap_8 FILLER_55_1645 ();
 sg13g2_decap_8 FILLER_55_1652 ();
 sg13g2_decap_8 FILLER_55_1659 ();
 sg13g2_decap_8 FILLER_55_1666 ();
 sg13g2_decap_8 FILLER_55_1673 ();
 sg13g2_decap_8 FILLER_55_1680 ();
 sg13g2_decap_8 FILLER_55_1687 ();
 sg13g2_decap_8 FILLER_55_1694 ();
 sg13g2_decap_8 FILLER_55_1701 ();
 sg13g2_decap_8 FILLER_55_1708 ();
 sg13g2_decap_8 FILLER_55_1715 ();
 sg13g2_decap_8 FILLER_55_1722 ();
 sg13g2_decap_8 FILLER_55_1729 ();
 sg13g2_decap_8 FILLER_55_1736 ();
 sg13g2_decap_8 FILLER_55_1743 ();
 sg13g2_decap_8 FILLER_55_1750 ();
 sg13g2_decap_8 FILLER_55_1757 ();
 sg13g2_decap_8 FILLER_55_1764 ();
 sg13g2_decap_8 FILLER_55_1771 ();
 sg13g2_decap_8 FILLER_55_1778 ();
 sg13g2_decap_8 FILLER_55_1785 ();
 sg13g2_decap_8 FILLER_55_1792 ();
 sg13g2_decap_8 FILLER_55_1799 ();
 sg13g2_decap_8 FILLER_55_1806 ();
 sg13g2_decap_8 FILLER_55_1813 ();
 sg13g2_decap_8 FILLER_55_1820 ();
 sg13g2_decap_8 FILLER_55_1827 ();
 sg13g2_decap_8 FILLER_55_1834 ();
 sg13g2_decap_8 FILLER_55_1841 ();
 sg13g2_decap_8 FILLER_55_1848 ();
 sg13g2_decap_8 FILLER_55_1855 ();
 sg13g2_decap_8 FILLER_55_1862 ();
 sg13g2_decap_8 FILLER_55_1869 ();
 sg13g2_decap_8 FILLER_55_1876 ();
 sg13g2_decap_8 FILLER_55_1883 ();
 sg13g2_decap_8 FILLER_55_1890 ();
 sg13g2_decap_8 FILLER_55_1897 ();
 sg13g2_decap_8 FILLER_55_1904 ();
 sg13g2_decap_8 FILLER_55_1911 ();
 sg13g2_decap_8 FILLER_55_1918 ();
 sg13g2_decap_8 FILLER_55_1925 ();
 sg13g2_decap_8 FILLER_55_1932 ();
 sg13g2_decap_8 FILLER_55_1939 ();
 sg13g2_decap_8 FILLER_55_1946 ();
 sg13g2_decap_8 FILLER_55_1953 ();
 sg13g2_decap_8 FILLER_55_1960 ();
 sg13g2_decap_8 FILLER_55_1967 ();
 sg13g2_decap_8 FILLER_55_1974 ();
 sg13g2_decap_8 FILLER_55_1981 ();
 sg13g2_decap_8 FILLER_55_1988 ();
 sg13g2_decap_8 FILLER_55_1995 ();
 sg13g2_decap_8 FILLER_55_2002 ();
 sg13g2_decap_8 FILLER_55_2009 ();
 sg13g2_decap_8 FILLER_55_2016 ();
 sg13g2_decap_8 FILLER_55_2023 ();
 sg13g2_decap_8 FILLER_55_2030 ();
 sg13g2_decap_8 FILLER_55_2037 ();
 sg13g2_decap_8 FILLER_55_2044 ();
 sg13g2_decap_8 FILLER_55_2051 ();
 sg13g2_decap_8 FILLER_55_2058 ();
 sg13g2_decap_8 FILLER_55_2065 ();
 sg13g2_decap_8 FILLER_55_2072 ();
 sg13g2_decap_8 FILLER_55_2079 ();
 sg13g2_decap_8 FILLER_55_2086 ();
 sg13g2_decap_8 FILLER_55_2093 ();
 sg13g2_decap_8 FILLER_55_2100 ();
 sg13g2_decap_8 FILLER_55_2107 ();
 sg13g2_decap_8 FILLER_55_2114 ();
 sg13g2_decap_8 FILLER_55_2121 ();
 sg13g2_decap_8 FILLER_55_2128 ();
 sg13g2_decap_8 FILLER_55_2135 ();
 sg13g2_decap_8 FILLER_55_2142 ();
 sg13g2_decap_8 FILLER_55_2149 ();
 sg13g2_decap_8 FILLER_55_2156 ();
 sg13g2_decap_8 FILLER_55_2163 ();
 sg13g2_decap_8 FILLER_55_2170 ();
 sg13g2_decap_8 FILLER_55_2177 ();
 sg13g2_decap_8 FILLER_55_2184 ();
 sg13g2_decap_8 FILLER_55_2191 ();
 sg13g2_decap_8 FILLER_55_2198 ();
 sg13g2_decap_8 FILLER_55_2205 ();
 sg13g2_decap_8 FILLER_55_2212 ();
 sg13g2_decap_8 FILLER_55_2219 ();
 sg13g2_decap_8 FILLER_55_2226 ();
 sg13g2_decap_8 FILLER_55_2233 ();
 sg13g2_decap_8 FILLER_55_2240 ();
 sg13g2_decap_8 FILLER_55_2247 ();
 sg13g2_decap_8 FILLER_55_2254 ();
 sg13g2_decap_8 FILLER_55_2261 ();
 sg13g2_decap_8 FILLER_55_2268 ();
 sg13g2_decap_8 FILLER_55_2275 ();
 sg13g2_decap_8 FILLER_55_2282 ();
 sg13g2_decap_8 FILLER_55_2289 ();
 sg13g2_decap_8 FILLER_55_2296 ();
 sg13g2_decap_8 FILLER_55_2303 ();
 sg13g2_decap_8 FILLER_55_2310 ();
 sg13g2_decap_8 FILLER_55_2317 ();
 sg13g2_decap_8 FILLER_55_2324 ();
 sg13g2_decap_8 FILLER_55_2331 ();
 sg13g2_decap_8 FILLER_55_2338 ();
 sg13g2_decap_8 FILLER_55_2345 ();
 sg13g2_decap_8 FILLER_55_2352 ();
 sg13g2_decap_8 FILLER_55_2359 ();
 sg13g2_decap_8 FILLER_55_2366 ();
 sg13g2_decap_8 FILLER_55_2373 ();
 sg13g2_decap_8 FILLER_55_2380 ();
 sg13g2_decap_8 FILLER_55_2387 ();
 sg13g2_decap_8 FILLER_55_2394 ();
 sg13g2_decap_8 FILLER_55_2401 ();
 sg13g2_decap_8 FILLER_55_2408 ();
 sg13g2_decap_8 FILLER_55_2415 ();
 sg13g2_decap_8 FILLER_55_2422 ();
 sg13g2_decap_8 FILLER_55_2429 ();
 sg13g2_decap_8 FILLER_55_2436 ();
 sg13g2_decap_8 FILLER_55_2443 ();
 sg13g2_decap_8 FILLER_55_2450 ();
 sg13g2_decap_8 FILLER_55_2457 ();
 sg13g2_decap_8 FILLER_55_2464 ();
 sg13g2_decap_8 FILLER_55_2471 ();
 sg13g2_decap_8 FILLER_55_2478 ();
 sg13g2_decap_8 FILLER_55_2485 ();
 sg13g2_decap_8 FILLER_55_2492 ();
 sg13g2_decap_8 FILLER_55_2499 ();
 sg13g2_decap_8 FILLER_55_2506 ();
 sg13g2_decap_8 FILLER_55_2513 ();
 sg13g2_decap_8 FILLER_55_2520 ();
 sg13g2_decap_8 FILLER_55_2527 ();
 sg13g2_decap_8 FILLER_55_2534 ();
 sg13g2_decap_8 FILLER_55_2541 ();
 sg13g2_decap_8 FILLER_55_2548 ();
 sg13g2_decap_8 FILLER_55_2555 ();
 sg13g2_decap_8 FILLER_55_2562 ();
 sg13g2_decap_8 FILLER_55_2569 ();
 sg13g2_decap_8 FILLER_55_2576 ();
 sg13g2_decap_8 FILLER_55_2583 ();
 sg13g2_decap_8 FILLER_55_2590 ();
 sg13g2_decap_8 FILLER_55_2597 ();
 sg13g2_decap_8 FILLER_55_2604 ();
 sg13g2_decap_8 FILLER_55_2611 ();
 sg13g2_decap_8 FILLER_55_2618 ();
 sg13g2_decap_8 FILLER_55_2625 ();
 sg13g2_decap_8 FILLER_55_2632 ();
 sg13g2_decap_8 FILLER_55_2639 ();
 sg13g2_decap_8 FILLER_55_2646 ();
 sg13g2_decap_8 FILLER_55_2653 ();
 sg13g2_decap_8 FILLER_55_2660 ();
 sg13g2_decap_8 FILLER_55_2667 ();
 sg13g2_decap_8 FILLER_55_2674 ();
 sg13g2_decap_8 FILLER_55_2681 ();
 sg13g2_decap_8 FILLER_55_2688 ();
 sg13g2_decap_8 FILLER_55_2695 ();
 sg13g2_decap_8 FILLER_55_2702 ();
 sg13g2_decap_8 FILLER_55_2709 ();
 sg13g2_decap_8 FILLER_55_2716 ();
 sg13g2_decap_8 FILLER_55_2723 ();
 sg13g2_decap_8 FILLER_55_2730 ();
 sg13g2_decap_8 FILLER_55_2737 ();
 sg13g2_decap_8 FILLER_55_2744 ();
 sg13g2_decap_8 FILLER_55_2751 ();
 sg13g2_decap_8 FILLER_55_2758 ();
 sg13g2_decap_8 FILLER_55_2765 ();
 sg13g2_decap_8 FILLER_55_2772 ();
 sg13g2_decap_8 FILLER_55_2779 ();
 sg13g2_decap_8 FILLER_55_2786 ();
 sg13g2_decap_8 FILLER_55_2793 ();
 sg13g2_decap_8 FILLER_55_2800 ();
 sg13g2_decap_8 FILLER_55_2807 ();
 sg13g2_decap_8 FILLER_55_2814 ();
 sg13g2_decap_8 FILLER_55_2821 ();
 sg13g2_decap_8 FILLER_55_2828 ();
 sg13g2_decap_8 FILLER_55_2835 ();
 sg13g2_decap_8 FILLER_55_2842 ();
 sg13g2_decap_8 FILLER_55_2849 ();
 sg13g2_decap_8 FILLER_55_2856 ();
 sg13g2_decap_8 FILLER_55_2863 ();
 sg13g2_decap_8 FILLER_55_2870 ();
 sg13g2_decap_8 FILLER_55_2877 ();
 sg13g2_decap_8 FILLER_55_2884 ();
 sg13g2_decap_8 FILLER_55_2891 ();
 sg13g2_decap_8 FILLER_55_2898 ();
 sg13g2_decap_8 FILLER_55_2905 ();
 sg13g2_decap_8 FILLER_55_2912 ();
 sg13g2_decap_8 FILLER_55_2919 ();
 sg13g2_decap_8 FILLER_55_2926 ();
 sg13g2_decap_8 FILLER_55_2933 ();
 sg13g2_decap_8 FILLER_55_2940 ();
 sg13g2_decap_8 FILLER_55_2947 ();
 sg13g2_decap_8 FILLER_55_2954 ();
 sg13g2_decap_8 FILLER_55_2961 ();
 sg13g2_decap_8 FILLER_55_2968 ();
 sg13g2_decap_8 FILLER_55_2975 ();
 sg13g2_decap_8 FILLER_55_2982 ();
 sg13g2_decap_8 FILLER_55_2989 ();
 sg13g2_decap_8 FILLER_55_2996 ();
 sg13g2_decap_8 FILLER_55_3003 ();
 sg13g2_decap_8 FILLER_55_3010 ();
 sg13g2_decap_8 FILLER_55_3017 ();
 sg13g2_decap_8 FILLER_55_3024 ();
 sg13g2_decap_8 FILLER_55_3031 ();
 sg13g2_decap_8 FILLER_55_3038 ();
 sg13g2_decap_8 FILLER_55_3045 ();
 sg13g2_decap_8 FILLER_55_3052 ();
 sg13g2_decap_8 FILLER_55_3059 ();
 sg13g2_decap_8 FILLER_55_3066 ();
 sg13g2_decap_8 FILLER_55_3073 ();
 sg13g2_decap_8 FILLER_55_3080 ();
 sg13g2_decap_8 FILLER_55_3087 ();
 sg13g2_decap_8 FILLER_55_3094 ();
 sg13g2_decap_8 FILLER_55_3101 ();
 sg13g2_decap_8 FILLER_55_3108 ();
 sg13g2_decap_8 FILLER_55_3115 ();
 sg13g2_decap_8 FILLER_55_3122 ();
 sg13g2_decap_8 FILLER_55_3129 ();
 sg13g2_decap_8 FILLER_55_3136 ();
 sg13g2_decap_8 FILLER_55_3143 ();
 sg13g2_decap_8 FILLER_55_3150 ();
 sg13g2_decap_8 FILLER_55_3157 ();
 sg13g2_decap_8 FILLER_55_3164 ();
 sg13g2_decap_8 FILLER_55_3171 ();
 sg13g2_decap_8 FILLER_55_3178 ();
 sg13g2_decap_8 FILLER_55_3185 ();
 sg13g2_decap_8 FILLER_55_3192 ();
 sg13g2_decap_8 FILLER_55_3199 ();
 sg13g2_decap_8 FILLER_55_3206 ();
 sg13g2_decap_8 FILLER_55_3213 ();
 sg13g2_decap_8 FILLER_55_3220 ();
 sg13g2_decap_8 FILLER_55_3227 ();
 sg13g2_decap_8 FILLER_55_3234 ();
 sg13g2_decap_8 FILLER_55_3241 ();
 sg13g2_decap_8 FILLER_55_3248 ();
 sg13g2_decap_8 FILLER_55_3255 ();
 sg13g2_decap_8 FILLER_55_3262 ();
 sg13g2_decap_8 FILLER_55_3269 ();
 sg13g2_decap_8 FILLER_55_3276 ();
 sg13g2_decap_8 FILLER_55_3283 ();
 sg13g2_decap_8 FILLER_55_3290 ();
 sg13g2_decap_8 FILLER_55_3297 ();
 sg13g2_decap_8 FILLER_55_3304 ();
 sg13g2_decap_8 FILLER_55_3311 ();
 sg13g2_decap_8 FILLER_55_3318 ();
 sg13g2_decap_8 FILLER_55_3325 ();
 sg13g2_decap_8 FILLER_55_3332 ();
 sg13g2_decap_8 FILLER_55_3339 ();
 sg13g2_decap_8 FILLER_55_3346 ();
 sg13g2_decap_8 FILLER_55_3353 ();
 sg13g2_decap_8 FILLER_55_3360 ();
 sg13g2_decap_8 FILLER_55_3367 ();
 sg13g2_decap_8 FILLER_55_3374 ();
 sg13g2_decap_8 FILLER_55_3381 ();
 sg13g2_decap_8 FILLER_55_3388 ();
 sg13g2_decap_8 FILLER_55_3395 ();
 sg13g2_decap_8 FILLER_55_3402 ();
 sg13g2_decap_8 FILLER_55_3409 ();
 sg13g2_decap_8 FILLER_55_3416 ();
 sg13g2_decap_8 FILLER_55_3423 ();
 sg13g2_decap_8 FILLER_55_3430 ();
 sg13g2_decap_8 FILLER_55_3437 ();
 sg13g2_decap_8 FILLER_55_3444 ();
 sg13g2_decap_8 FILLER_55_3451 ();
 sg13g2_decap_8 FILLER_55_3458 ();
 sg13g2_decap_8 FILLER_55_3465 ();
 sg13g2_decap_8 FILLER_55_3472 ();
 sg13g2_decap_8 FILLER_55_3479 ();
 sg13g2_decap_8 FILLER_55_3486 ();
 sg13g2_decap_8 FILLER_55_3493 ();
 sg13g2_decap_8 FILLER_55_3500 ();
 sg13g2_decap_8 FILLER_55_3507 ();
 sg13g2_decap_8 FILLER_55_3514 ();
 sg13g2_decap_8 FILLER_55_3521 ();
 sg13g2_decap_8 FILLER_55_3528 ();
 sg13g2_decap_8 FILLER_55_3535 ();
 sg13g2_decap_8 FILLER_55_3542 ();
 sg13g2_decap_8 FILLER_55_3549 ();
 sg13g2_decap_8 FILLER_55_3556 ();
 sg13g2_decap_8 FILLER_55_3563 ();
 sg13g2_decap_8 FILLER_55_3570 ();
 sg13g2_fill_2 FILLER_55_3577 ();
 sg13g2_fill_1 FILLER_55_3579 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_decap_8 FILLER_56_105 ();
 sg13g2_decap_8 FILLER_56_112 ();
 sg13g2_decap_8 FILLER_56_119 ();
 sg13g2_decap_8 FILLER_56_126 ();
 sg13g2_decap_8 FILLER_56_133 ();
 sg13g2_decap_8 FILLER_56_140 ();
 sg13g2_decap_8 FILLER_56_147 ();
 sg13g2_decap_8 FILLER_56_154 ();
 sg13g2_decap_8 FILLER_56_161 ();
 sg13g2_decap_8 FILLER_56_168 ();
 sg13g2_decap_8 FILLER_56_175 ();
 sg13g2_decap_8 FILLER_56_182 ();
 sg13g2_decap_8 FILLER_56_189 ();
 sg13g2_decap_8 FILLER_56_196 ();
 sg13g2_decap_8 FILLER_56_203 ();
 sg13g2_decap_8 FILLER_56_210 ();
 sg13g2_decap_8 FILLER_56_217 ();
 sg13g2_decap_8 FILLER_56_224 ();
 sg13g2_decap_8 FILLER_56_231 ();
 sg13g2_decap_8 FILLER_56_238 ();
 sg13g2_decap_8 FILLER_56_245 ();
 sg13g2_decap_8 FILLER_56_252 ();
 sg13g2_decap_8 FILLER_56_259 ();
 sg13g2_decap_8 FILLER_56_266 ();
 sg13g2_decap_8 FILLER_56_273 ();
 sg13g2_decap_8 FILLER_56_280 ();
 sg13g2_decap_8 FILLER_56_287 ();
 sg13g2_decap_8 FILLER_56_294 ();
 sg13g2_decap_8 FILLER_56_301 ();
 sg13g2_decap_8 FILLER_56_308 ();
 sg13g2_decap_8 FILLER_56_315 ();
 sg13g2_decap_8 FILLER_56_322 ();
 sg13g2_decap_8 FILLER_56_329 ();
 sg13g2_decap_8 FILLER_56_336 ();
 sg13g2_decap_8 FILLER_56_343 ();
 sg13g2_decap_8 FILLER_56_350 ();
 sg13g2_decap_8 FILLER_56_357 ();
 sg13g2_decap_8 FILLER_56_364 ();
 sg13g2_decap_8 FILLER_56_371 ();
 sg13g2_decap_8 FILLER_56_378 ();
 sg13g2_decap_8 FILLER_56_385 ();
 sg13g2_decap_8 FILLER_56_392 ();
 sg13g2_decap_8 FILLER_56_399 ();
 sg13g2_decap_8 FILLER_56_406 ();
 sg13g2_decap_8 FILLER_56_413 ();
 sg13g2_decap_8 FILLER_56_420 ();
 sg13g2_decap_8 FILLER_56_427 ();
 sg13g2_decap_8 FILLER_56_434 ();
 sg13g2_decap_8 FILLER_56_441 ();
 sg13g2_decap_8 FILLER_56_448 ();
 sg13g2_decap_8 FILLER_56_455 ();
 sg13g2_decap_8 FILLER_56_462 ();
 sg13g2_decap_8 FILLER_56_469 ();
 sg13g2_decap_8 FILLER_56_476 ();
 sg13g2_decap_8 FILLER_56_483 ();
 sg13g2_decap_8 FILLER_56_490 ();
 sg13g2_decap_8 FILLER_56_497 ();
 sg13g2_decap_8 FILLER_56_504 ();
 sg13g2_decap_8 FILLER_56_511 ();
 sg13g2_decap_8 FILLER_56_518 ();
 sg13g2_decap_8 FILLER_56_525 ();
 sg13g2_decap_8 FILLER_56_532 ();
 sg13g2_decap_8 FILLER_56_539 ();
 sg13g2_decap_8 FILLER_56_546 ();
 sg13g2_decap_8 FILLER_56_553 ();
 sg13g2_decap_8 FILLER_56_560 ();
 sg13g2_decap_8 FILLER_56_567 ();
 sg13g2_decap_8 FILLER_56_574 ();
 sg13g2_decap_8 FILLER_56_581 ();
 sg13g2_decap_8 FILLER_56_588 ();
 sg13g2_decap_8 FILLER_56_595 ();
 sg13g2_decap_8 FILLER_56_602 ();
 sg13g2_decap_8 FILLER_56_609 ();
 sg13g2_decap_8 FILLER_56_616 ();
 sg13g2_decap_8 FILLER_56_623 ();
 sg13g2_decap_8 FILLER_56_630 ();
 sg13g2_decap_8 FILLER_56_637 ();
 sg13g2_decap_8 FILLER_56_644 ();
 sg13g2_decap_8 FILLER_56_651 ();
 sg13g2_decap_8 FILLER_56_658 ();
 sg13g2_decap_8 FILLER_56_665 ();
 sg13g2_decap_8 FILLER_56_672 ();
 sg13g2_decap_8 FILLER_56_679 ();
 sg13g2_decap_8 FILLER_56_686 ();
 sg13g2_decap_8 FILLER_56_693 ();
 sg13g2_decap_8 FILLER_56_700 ();
 sg13g2_decap_8 FILLER_56_707 ();
 sg13g2_decap_8 FILLER_56_714 ();
 sg13g2_decap_8 FILLER_56_721 ();
 sg13g2_decap_8 FILLER_56_728 ();
 sg13g2_decap_8 FILLER_56_735 ();
 sg13g2_decap_8 FILLER_56_742 ();
 sg13g2_decap_8 FILLER_56_749 ();
 sg13g2_decap_8 FILLER_56_756 ();
 sg13g2_decap_8 FILLER_56_763 ();
 sg13g2_decap_8 FILLER_56_770 ();
 sg13g2_decap_8 FILLER_56_777 ();
 sg13g2_decap_8 FILLER_56_784 ();
 sg13g2_decap_8 FILLER_56_791 ();
 sg13g2_decap_8 FILLER_56_798 ();
 sg13g2_decap_8 FILLER_56_805 ();
 sg13g2_decap_8 FILLER_56_812 ();
 sg13g2_decap_8 FILLER_56_819 ();
 sg13g2_decap_8 FILLER_56_826 ();
 sg13g2_decap_8 FILLER_56_833 ();
 sg13g2_decap_8 FILLER_56_840 ();
 sg13g2_decap_8 FILLER_56_847 ();
 sg13g2_decap_8 FILLER_56_854 ();
 sg13g2_decap_8 FILLER_56_861 ();
 sg13g2_decap_8 FILLER_56_868 ();
 sg13g2_decap_8 FILLER_56_875 ();
 sg13g2_decap_8 FILLER_56_882 ();
 sg13g2_decap_8 FILLER_56_889 ();
 sg13g2_decap_8 FILLER_56_896 ();
 sg13g2_decap_8 FILLER_56_903 ();
 sg13g2_decap_8 FILLER_56_910 ();
 sg13g2_decap_8 FILLER_56_917 ();
 sg13g2_decap_8 FILLER_56_924 ();
 sg13g2_decap_8 FILLER_56_931 ();
 sg13g2_decap_8 FILLER_56_938 ();
 sg13g2_decap_8 FILLER_56_945 ();
 sg13g2_decap_8 FILLER_56_952 ();
 sg13g2_decap_8 FILLER_56_959 ();
 sg13g2_decap_8 FILLER_56_966 ();
 sg13g2_decap_8 FILLER_56_973 ();
 sg13g2_decap_8 FILLER_56_980 ();
 sg13g2_decap_8 FILLER_56_987 ();
 sg13g2_decap_8 FILLER_56_994 ();
 sg13g2_decap_8 FILLER_56_1001 ();
 sg13g2_decap_8 FILLER_56_1008 ();
 sg13g2_decap_8 FILLER_56_1015 ();
 sg13g2_decap_8 FILLER_56_1022 ();
 sg13g2_decap_8 FILLER_56_1029 ();
 sg13g2_decap_8 FILLER_56_1036 ();
 sg13g2_decap_8 FILLER_56_1043 ();
 sg13g2_decap_8 FILLER_56_1050 ();
 sg13g2_decap_8 FILLER_56_1057 ();
 sg13g2_decap_8 FILLER_56_1064 ();
 sg13g2_decap_8 FILLER_56_1071 ();
 sg13g2_decap_8 FILLER_56_1078 ();
 sg13g2_decap_8 FILLER_56_1085 ();
 sg13g2_decap_8 FILLER_56_1092 ();
 sg13g2_decap_8 FILLER_56_1099 ();
 sg13g2_decap_8 FILLER_56_1106 ();
 sg13g2_decap_8 FILLER_56_1113 ();
 sg13g2_decap_8 FILLER_56_1120 ();
 sg13g2_decap_8 FILLER_56_1127 ();
 sg13g2_decap_8 FILLER_56_1134 ();
 sg13g2_decap_8 FILLER_56_1141 ();
 sg13g2_decap_8 FILLER_56_1148 ();
 sg13g2_decap_8 FILLER_56_1155 ();
 sg13g2_decap_8 FILLER_56_1162 ();
 sg13g2_decap_8 FILLER_56_1169 ();
 sg13g2_decap_8 FILLER_56_1176 ();
 sg13g2_decap_8 FILLER_56_1183 ();
 sg13g2_decap_8 FILLER_56_1190 ();
 sg13g2_decap_8 FILLER_56_1197 ();
 sg13g2_decap_8 FILLER_56_1204 ();
 sg13g2_decap_8 FILLER_56_1211 ();
 sg13g2_decap_8 FILLER_56_1218 ();
 sg13g2_decap_8 FILLER_56_1225 ();
 sg13g2_decap_8 FILLER_56_1232 ();
 sg13g2_decap_8 FILLER_56_1239 ();
 sg13g2_decap_8 FILLER_56_1246 ();
 sg13g2_decap_8 FILLER_56_1253 ();
 sg13g2_decap_8 FILLER_56_1260 ();
 sg13g2_decap_8 FILLER_56_1267 ();
 sg13g2_decap_8 FILLER_56_1274 ();
 sg13g2_decap_8 FILLER_56_1281 ();
 sg13g2_decap_8 FILLER_56_1288 ();
 sg13g2_decap_8 FILLER_56_1295 ();
 sg13g2_decap_8 FILLER_56_1302 ();
 sg13g2_decap_8 FILLER_56_1309 ();
 sg13g2_decap_8 FILLER_56_1316 ();
 sg13g2_decap_8 FILLER_56_1323 ();
 sg13g2_decap_8 FILLER_56_1330 ();
 sg13g2_decap_8 FILLER_56_1337 ();
 sg13g2_decap_8 FILLER_56_1344 ();
 sg13g2_decap_8 FILLER_56_1351 ();
 sg13g2_decap_8 FILLER_56_1358 ();
 sg13g2_decap_8 FILLER_56_1365 ();
 sg13g2_decap_8 FILLER_56_1372 ();
 sg13g2_decap_8 FILLER_56_1379 ();
 sg13g2_decap_8 FILLER_56_1386 ();
 sg13g2_decap_8 FILLER_56_1393 ();
 sg13g2_decap_8 FILLER_56_1400 ();
 sg13g2_decap_8 FILLER_56_1407 ();
 sg13g2_decap_8 FILLER_56_1414 ();
 sg13g2_decap_8 FILLER_56_1421 ();
 sg13g2_decap_8 FILLER_56_1428 ();
 sg13g2_decap_8 FILLER_56_1435 ();
 sg13g2_decap_8 FILLER_56_1442 ();
 sg13g2_decap_8 FILLER_56_1449 ();
 sg13g2_decap_8 FILLER_56_1456 ();
 sg13g2_decap_8 FILLER_56_1463 ();
 sg13g2_decap_8 FILLER_56_1470 ();
 sg13g2_decap_8 FILLER_56_1477 ();
 sg13g2_decap_8 FILLER_56_1484 ();
 sg13g2_decap_8 FILLER_56_1491 ();
 sg13g2_decap_8 FILLER_56_1498 ();
 sg13g2_decap_8 FILLER_56_1505 ();
 sg13g2_decap_8 FILLER_56_1512 ();
 sg13g2_decap_8 FILLER_56_1519 ();
 sg13g2_decap_8 FILLER_56_1526 ();
 sg13g2_decap_8 FILLER_56_1533 ();
 sg13g2_decap_8 FILLER_56_1540 ();
 sg13g2_decap_8 FILLER_56_1547 ();
 sg13g2_decap_8 FILLER_56_1554 ();
 sg13g2_decap_8 FILLER_56_1561 ();
 sg13g2_decap_8 FILLER_56_1568 ();
 sg13g2_decap_8 FILLER_56_1575 ();
 sg13g2_decap_8 FILLER_56_1582 ();
 sg13g2_decap_8 FILLER_56_1589 ();
 sg13g2_decap_8 FILLER_56_1596 ();
 sg13g2_decap_8 FILLER_56_1603 ();
 sg13g2_decap_8 FILLER_56_1610 ();
 sg13g2_decap_8 FILLER_56_1617 ();
 sg13g2_decap_8 FILLER_56_1624 ();
 sg13g2_decap_8 FILLER_56_1631 ();
 sg13g2_decap_8 FILLER_56_1638 ();
 sg13g2_decap_8 FILLER_56_1645 ();
 sg13g2_decap_8 FILLER_56_1652 ();
 sg13g2_decap_8 FILLER_56_1659 ();
 sg13g2_decap_8 FILLER_56_1666 ();
 sg13g2_decap_8 FILLER_56_1673 ();
 sg13g2_decap_8 FILLER_56_1680 ();
 sg13g2_decap_8 FILLER_56_1687 ();
 sg13g2_decap_8 FILLER_56_1694 ();
 sg13g2_decap_8 FILLER_56_1701 ();
 sg13g2_decap_8 FILLER_56_1708 ();
 sg13g2_decap_8 FILLER_56_1715 ();
 sg13g2_decap_8 FILLER_56_1722 ();
 sg13g2_decap_8 FILLER_56_1729 ();
 sg13g2_decap_8 FILLER_56_1736 ();
 sg13g2_decap_8 FILLER_56_1743 ();
 sg13g2_decap_8 FILLER_56_1750 ();
 sg13g2_decap_8 FILLER_56_1757 ();
 sg13g2_decap_8 FILLER_56_1764 ();
 sg13g2_decap_8 FILLER_56_1771 ();
 sg13g2_decap_8 FILLER_56_1778 ();
 sg13g2_decap_8 FILLER_56_1785 ();
 sg13g2_decap_8 FILLER_56_1792 ();
 sg13g2_decap_8 FILLER_56_1799 ();
 sg13g2_decap_8 FILLER_56_1806 ();
 sg13g2_decap_8 FILLER_56_1813 ();
 sg13g2_decap_8 FILLER_56_1820 ();
 sg13g2_decap_8 FILLER_56_1827 ();
 sg13g2_decap_8 FILLER_56_1834 ();
 sg13g2_decap_8 FILLER_56_1841 ();
 sg13g2_decap_8 FILLER_56_1848 ();
 sg13g2_decap_8 FILLER_56_1855 ();
 sg13g2_decap_8 FILLER_56_1862 ();
 sg13g2_decap_8 FILLER_56_1869 ();
 sg13g2_decap_8 FILLER_56_1876 ();
 sg13g2_decap_8 FILLER_56_1883 ();
 sg13g2_decap_8 FILLER_56_1890 ();
 sg13g2_decap_8 FILLER_56_1897 ();
 sg13g2_decap_8 FILLER_56_1904 ();
 sg13g2_decap_8 FILLER_56_1911 ();
 sg13g2_decap_8 FILLER_56_1918 ();
 sg13g2_decap_8 FILLER_56_1925 ();
 sg13g2_decap_8 FILLER_56_1932 ();
 sg13g2_decap_8 FILLER_56_1939 ();
 sg13g2_decap_8 FILLER_56_1946 ();
 sg13g2_decap_8 FILLER_56_1953 ();
 sg13g2_decap_8 FILLER_56_1960 ();
 sg13g2_decap_8 FILLER_56_1967 ();
 sg13g2_decap_8 FILLER_56_1974 ();
 sg13g2_decap_8 FILLER_56_1981 ();
 sg13g2_decap_8 FILLER_56_1988 ();
 sg13g2_decap_8 FILLER_56_1995 ();
 sg13g2_decap_8 FILLER_56_2002 ();
 sg13g2_decap_8 FILLER_56_2009 ();
 sg13g2_decap_8 FILLER_56_2016 ();
 sg13g2_decap_8 FILLER_56_2023 ();
 sg13g2_decap_8 FILLER_56_2030 ();
 sg13g2_decap_8 FILLER_56_2037 ();
 sg13g2_decap_8 FILLER_56_2044 ();
 sg13g2_decap_8 FILLER_56_2051 ();
 sg13g2_decap_8 FILLER_56_2058 ();
 sg13g2_decap_8 FILLER_56_2065 ();
 sg13g2_decap_8 FILLER_56_2072 ();
 sg13g2_decap_8 FILLER_56_2079 ();
 sg13g2_decap_8 FILLER_56_2086 ();
 sg13g2_decap_8 FILLER_56_2093 ();
 sg13g2_decap_8 FILLER_56_2100 ();
 sg13g2_decap_8 FILLER_56_2107 ();
 sg13g2_decap_8 FILLER_56_2114 ();
 sg13g2_decap_8 FILLER_56_2121 ();
 sg13g2_decap_8 FILLER_56_2128 ();
 sg13g2_decap_8 FILLER_56_2135 ();
 sg13g2_decap_8 FILLER_56_2142 ();
 sg13g2_decap_8 FILLER_56_2149 ();
 sg13g2_decap_8 FILLER_56_2156 ();
 sg13g2_decap_8 FILLER_56_2163 ();
 sg13g2_decap_8 FILLER_56_2170 ();
 sg13g2_decap_8 FILLER_56_2177 ();
 sg13g2_decap_8 FILLER_56_2184 ();
 sg13g2_decap_8 FILLER_56_2191 ();
 sg13g2_decap_8 FILLER_56_2198 ();
 sg13g2_decap_8 FILLER_56_2205 ();
 sg13g2_decap_8 FILLER_56_2212 ();
 sg13g2_decap_8 FILLER_56_2219 ();
 sg13g2_decap_8 FILLER_56_2226 ();
 sg13g2_decap_8 FILLER_56_2233 ();
 sg13g2_decap_8 FILLER_56_2240 ();
 sg13g2_decap_8 FILLER_56_2247 ();
 sg13g2_decap_8 FILLER_56_2254 ();
 sg13g2_decap_8 FILLER_56_2261 ();
 sg13g2_decap_8 FILLER_56_2268 ();
 sg13g2_decap_8 FILLER_56_2275 ();
 sg13g2_decap_8 FILLER_56_2282 ();
 sg13g2_decap_8 FILLER_56_2289 ();
 sg13g2_decap_8 FILLER_56_2296 ();
 sg13g2_decap_8 FILLER_56_2303 ();
 sg13g2_decap_8 FILLER_56_2310 ();
 sg13g2_decap_8 FILLER_56_2317 ();
 sg13g2_decap_8 FILLER_56_2324 ();
 sg13g2_decap_8 FILLER_56_2331 ();
 sg13g2_decap_8 FILLER_56_2338 ();
 sg13g2_decap_8 FILLER_56_2345 ();
 sg13g2_decap_8 FILLER_56_2352 ();
 sg13g2_decap_8 FILLER_56_2359 ();
 sg13g2_decap_8 FILLER_56_2366 ();
 sg13g2_decap_8 FILLER_56_2373 ();
 sg13g2_decap_8 FILLER_56_2380 ();
 sg13g2_decap_8 FILLER_56_2387 ();
 sg13g2_decap_8 FILLER_56_2394 ();
 sg13g2_decap_8 FILLER_56_2401 ();
 sg13g2_decap_8 FILLER_56_2408 ();
 sg13g2_decap_8 FILLER_56_2415 ();
 sg13g2_decap_8 FILLER_56_2422 ();
 sg13g2_decap_8 FILLER_56_2429 ();
 sg13g2_decap_8 FILLER_56_2436 ();
 sg13g2_decap_8 FILLER_56_2443 ();
 sg13g2_decap_8 FILLER_56_2450 ();
 sg13g2_decap_8 FILLER_56_2457 ();
 sg13g2_decap_8 FILLER_56_2464 ();
 sg13g2_decap_8 FILLER_56_2471 ();
 sg13g2_decap_8 FILLER_56_2478 ();
 sg13g2_decap_8 FILLER_56_2485 ();
 sg13g2_decap_8 FILLER_56_2492 ();
 sg13g2_decap_8 FILLER_56_2499 ();
 sg13g2_decap_8 FILLER_56_2506 ();
 sg13g2_decap_8 FILLER_56_2513 ();
 sg13g2_decap_8 FILLER_56_2520 ();
 sg13g2_decap_8 FILLER_56_2527 ();
 sg13g2_decap_8 FILLER_56_2534 ();
 sg13g2_decap_8 FILLER_56_2541 ();
 sg13g2_decap_8 FILLER_56_2548 ();
 sg13g2_decap_8 FILLER_56_2555 ();
 sg13g2_decap_8 FILLER_56_2562 ();
 sg13g2_decap_8 FILLER_56_2569 ();
 sg13g2_decap_8 FILLER_56_2576 ();
 sg13g2_decap_8 FILLER_56_2583 ();
 sg13g2_decap_8 FILLER_56_2590 ();
 sg13g2_decap_8 FILLER_56_2597 ();
 sg13g2_decap_8 FILLER_56_2604 ();
 sg13g2_decap_8 FILLER_56_2611 ();
 sg13g2_decap_8 FILLER_56_2618 ();
 sg13g2_decap_8 FILLER_56_2625 ();
 sg13g2_decap_8 FILLER_56_2632 ();
 sg13g2_decap_8 FILLER_56_2639 ();
 sg13g2_decap_8 FILLER_56_2646 ();
 sg13g2_decap_8 FILLER_56_2653 ();
 sg13g2_decap_8 FILLER_56_2660 ();
 sg13g2_decap_8 FILLER_56_2667 ();
 sg13g2_decap_8 FILLER_56_2674 ();
 sg13g2_decap_8 FILLER_56_2681 ();
 sg13g2_decap_8 FILLER_56_2688 ();
 sg13g2_decap_8 FILLER_56_2695 ();
 sg13g2_decap_8 FILLER_56_2702 ();
 sg13g2_decap_8 FILLER_56_2709 ();
 sg13g2_decap_8 FILLER_56_2716 ();
 sg13g2_decap_8 FILLER_56_2723 ();
 sg13g2_decap_8 FILLER_56_2730 ();
 sg13g2_decap_8 FILLER_56_2737 ();
 sg13g2_decap_8 FILLER_56_2744 ();
 sg13g2_decap_8 FILLER_56_2751 ();
 sg13g2_decap_8 FILLER_56_2758 ();
 sg13g2_decap_8 FILLER_56_2765 ();
 sg13g2_decap_8 FILLER_56_2772 ();
 sg13g2_decap_8 FILLER_56_2779 ();
 sg13g2_decap_8 FILLER_56_2786 ();
 sg13g2_decap_8 FILLER_56_2793 ();
 sg13g2_decap_8 FILLER_56_2800 ();
 sg13g2_decap_8 FILLER_56_2807 ();
 sg13g2_decap_8 FILLER_56_2814 ();
 sg13g2_decap_8 FILLER_56_2821 ();
 sg13g2_decap_8 FILLER_56_2828 ();
 sg13g2_decap_8 FILLER_56_2835 ();
 sg13g2_decap_8 FILLER_56_2842 ();
 sg13g2_decap_8 FILLER_56_2849 ();
 sg13g2_decap_8 FILLER_56_2856 ();
 sg13g2_decap_8 FILLER_56_2863 ();
 sg13g2_decap_8 FILLER_56_2870 ();
 sg13g2_decap_8 FILLER_56_2877 ();
 sg13g2_decap_8 FILLER_56_2884 ();
 sg13g2_decap_8 FILLER_56_2891 ();
 sg13g2_decap_8 FILLER_56_2898 ();
 sg13g2_decap_8 FILLER_56_2905 ();
 sg13g2_decap_8 FILLER_56_2912 ();
 sg13g2_decap_8 FILLER_56_2919 ();
 sg13g2_decap_8 FILLER_56_2926 ();
 sg13g2_decap_8 FILLER_56_2933 ();
 sg13g2_decap_8 FILLER_56_2940 ();
 sg13g2_decap_8 FILLER_56_2947 ();
 sg13g2_decap_8 FILLER_56_2954 ();
 sg13g2_decap_8 FILLER_56_2961 ();
 sg13g2_decap_8 FILLER_56_2968 ();
 sg13g2_decap_8 FILLER_56_2975 ();
 sg13g2_decap_8 FILLER_56_2982 ();
 sg13g2_decap_8 FILLER_56_2989 ();
 sg13g2_decap_8 FILLER_56_2996 ();
 sg13g2_decap_8 FILLER_56_3003 ();
 sg13g2_decap_8 FILLER_56_3010 ();
 sg13g2_decap_8 FILLER_56_3017 ();
 sg13g2_decap_8 FILLER_56_3024 ();
 sg13g2_decap_8 FILLER_56_3031 ();
 sg13g2_decap_8 FILLER_56_3038 ();
 sg13g2_decap_8 FILLER_56_3045 ();
 sg13g2_decap_8 FILLER_56_3052 ();
 sg13g2_decap_8 FILLER_56_3059 ();
 sg13g2_decap_8 FILLER_56_3066 ();
 sg13g2_decap_8 FILLER_56_3073 ();
 sg13g2_decap_8 FILLER_56_3080 ();
 sg13g2_decap_8 FILLER_56_3087 ();
 sg13g2_decap_8 FILLER_56_3094 ();
 sg13g2_decap_8 FILLER_56_3101 ();
 sg13g2_decap_8 FILLER_56_3108 ();
 sg13g2_decap_8 FILLER_56_3115 ();
 sg13g2_decap_8 FILLER_56_3122 ();
 sg13g2_decap_8 FILLER_56_3129 ();
 sg13g2_decap_8 FILLER_56_3136 ();
 sg13g2_decap_8 FILLER_56_3143 ();
 sg13g2_decap_8 FILLER_56_3150 ();
 sg13g2_decap_8 FILLER_56_3157 ();
 sg13g2_decap_8 FILLER_56_3164 ();
 sg13g2_decap_8 FILLER_56_3171 ();
 sg13g2_decap_8 FILLER_56_3178 ();
 sg13g2_decap_8 FILLER_56_3185 ();
 sg13g2_decap_8 FILLER_56_3192 ();
 sg13g2_decap_8 FILLER_56_3199 ();
 sg13g2_decap_8 FILLER_56_3206 ();
 sg13g2_decap_8 FILLER_56_3213 ();
 sg13g2_decap_8 FILLER_56_3220 ();
 sg13g2_decap_8 FILLER_56_3227 ();
 sg13g2_decap_8 FILLER_56_3234 ();
 sg13g2_decap_8 FILLER_56_3241 ();
 sg13g2_decap_8 FILLER_56_3248 ();
 sg13g2_decap_8 FILLER_56_3255 ();
 sg13g2_decap_8 FILLER_56_3262 ();
 sg13g2_decap_8 FILLER_56_3269 ();
 sg13g2_decap_8 FILLER_56_3276 ();
 sg13g2_decap_8 FILLER_56_3283 ();
 sg13g2_decap_8 FILLER_56_3290 ();
 sg13g2_decap_8 FILLER_56_3297 ();
 sg13g2_decap_8 FILLER_56_3304 ();
 sg13g2_decap_8 FILLER_56_3311 ();
 sg13g2_decap_8 FILLER_56_3318 ();
 sg13g2_decap_8 FILLER_56_3325 ();
 sg13g2_decap_8 FILLER_56_3332 ();
 sg13g2_decap_8 FILLER_56_3339 ();
 sg13g2_decap_8 FILLER_56_3346 ();
 sg13g2_decap_8 FILLER_56_3353 ();
 sg13g2_decap_8 FILLER_56_3360 ();
 sg13g2_decap_8 FILLER_56_3367 ();
 sg13g2_decap_8 FILLER_56_3374 ();
 sg13g2_decap_8 FILLER_56_3381 ();
 sg13g2_decap_8 FILLER_56_3388 ();
 sg13g2_decap_8 FILLER_56_3395 ();
 sg13g2_decap_8 FILLER_56_3402 ();
 sg13g2_decap_8 FILLER_56_3409 ();
 sg13g2_decap_8 FILLER_56_3416 ();
 sg13g2_decap_8 FILLER_56_3423 ();
 sg13g2_decap_8 FILLER_56_3430 ();
 sg13g2_decap_8 FILLER_56_3437 ();
 sg13g2_decap_8 FILLER_56_3444 ();
 sg13g2_decap_8 FILLER_56_3451 ();
 sg13g2_decap_8 FILLER_56_3458 ();
 sg13g2_decap_8 FILLER_56_3465 ();
 sg13g2_decap_8 FILLER_56_3472 ();
 sg13g2_decap_8 FILLER_56_3479 ();
 sg13g2_decap_8 FILLER_56_3486 ();
 sg13g2_decap_8 FILLER_56_3493 ();
 sg13g2_decap_8 FILLER_56_3500 ();
 sg13g2_decap_8 FILLER_56_3507 ();
 sg13g2_decap_8 FILLER_56_3514 ();
 sg13g2_decap_8 FILLER_56_3521 ();
 sg13g2_decap_8 FILLER_56_3528 ();
 sg13g2_decap_8 FILLER_56_3535 ();
 sg13g2_decap_8 FILLER_56_3542 ();
 sg13g2_decap_8 FILLER_56_3549 ();
 sg13g2_decap_8 FILLER_56_3556 ();
 sg13g2_decap_8 FILLER_56_3563 ();
 sg13g2_decap_8 FILLER_56_3570 ();
 sg13g2_fill_2 FILLER_56_3577 ();
 sg13g2_fill_1 FILLER_56_3579 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_98 ();
 sg13g2_decap_8 FILLER_57_105 ();
 sg13g2_decap_8 FILLER_57_112 ();
 sg13g2_decap_8 FILLER_57_119 ();
 sg13g2_decap_8 FILLER_57_126 ();
 sg13g2_decap_8 FILLER_57_133 ();
 sg13g2_decap_8 FILLER_57_140 ();
 sg13g2_decap_8 FILLER_57_147 ();
 sg13g2_decap_8 FILLER_57_154 ();
 sg13g2_decap_8 FILLER_57_161 ();
 sg13g2_decap_8 FILLER_57_168 ();
 sg13g2_decap_8 FILLER_57_175 ();
 sg13g2_decap_8 FILLER_57_182 ();
 sg13g2_decap_8 FILLER_57_189 ();
 sg13g2_decap_8 FILLER_57_196 ();
 sg13g2_decap_8 FILLER_57_203 ();
 sg13g2_decap_8 FILLER_57_210 ();
 sg13g2_decap_8 FILLER_57_217 ();
 sg13g2_decap_8 FILLER_57_224 ();
 sg13g2_decap_8 FILLER_57_231 ();
 sg13g2_decap_8 FILLER_57_238 ();
 sg13g2_decap_8 FILLER_57_245 ();
 sg13g2_decap_8 FILLER_57_252 ();
 sg13g2_decap_8 FILLER_57_259 ();
 sg13g2_decap_8 FILLER_57_266 ();
 sg13g2_decap_8 FILLER_57_273 ();
 sg13g2_decap_8 FILLER_57_280 ();
 sg13g2_decap_8 FILLER_57_287 ();
 sg13g2_decap_8 FILLER_57_294 ();
 sg13g2_decap_8 FILLER_57_301 ();
 sg13g2_decap_8 FILLER_57_308 ();
 sg13g2_decap_8 FILLER_57_315 ();
 sg13g2_decap_8 FILLER_57_322 ();
 sg13g2_decap_8 FILLER_57_329 ();
 sg13g2_decap_8 FILLER_57_336 ();
 sg13g2_decap_8 FILLER_57_343 ();
 sg13g2_decap_8 FILLER_57_350 ();
 sg13g2_decap_8 FILLER_57_357 ();
 sg13g2_decap_8 FILLER_57_364 ();
 sg13g2_decap_8 FILLER_57_371 ();
 sg13g2_decap_8 FILLER_57_378 ();
 sg13g2_decap_8 FILLER_57_385 ();
 sg13g2_decap_8 FILLER_57_392 ();
 sg13g2_decap_8 FILLER_57_399 ();
 sg13g2_decap_8 FILLER_57_406 ();
 sg13g2_decap_8 FILLER_57_413 ();
 sg13g2_decap_8 FILLER_57_420 ();
 sg13g2_decap_8 FILLER_57_427 ();
 sg13g2_decap_8 FILLER_57_434 ();
 sg13g2_decap_8 FILLER_57_441 ();
 sg13g2_decap_8 FILLER_57_448 ();
 sg13g2_decap_8 FILLER_57_455 ();
 sg13g2_decap_8 FILLER_57_462 ();
 sg13g2_decap_8 FILLER_57_469 ();
 sg13g2_decap_8 FILLER_57_476 ();
 sg13g2_decap_8 FILLER_57_483 ();
 sg13g2_decap_8 FILLER_57_490 ();
 sg13g2_decap_8 FILLER_57_497 ();
 sg13g2_decap_8 FILLER_57_504 ();
 sg13g2_decap_8 FILLER_57_511 ();
 sg13g2_decap_8 FILLER_57_518 ();
 sg13g2_decap_8 FILLER_57_525 ();
 sg13g2_decap_8 FILLER_57_532 ();
 sg13g2_decap_8 FILLER_57_539 ();
 sg13g2_decap_8 FILLER_57_546 ();
 sg13g2_decap_8 FILLER_57_553 ();
 sg13g2_decap_8 FILLER_57_560 ();
 sg13g2_decap_8 FILLER_57_567 ();
 sg13g2_decap_8 FILLER_57_574 ();
 sg13g2_decap_8 FILLER_57_581 ();
 sg13g2_decap_8 FILLER_57_588 ();
 sg13g2_decap_8 FILLER_57_595 ();
 sg13g2_decap_8 FILLER_57_602 ();
 sg13g2_decap_8 FILLER_57_609 ();
 sg13g2_decap_8 FILLER_57_616 ();
 sg13g2_decap_8 FILLER_57_623 ();
 sg13g2_decap_8 FILLER_57_630 ();
 sg13g2_decap_8 FILLER_57_637 ();
 sg13g2_decap_8 FILLER_57_644 ();
 sg13g2_decap_8 FILLER_57_651 ();
 sg13g2_decap_8 FILLER_57_658 ();
 sg13g2_decap_8 FILLER_57_665 ();
 sg13g2_decap_8 FILLER_57_672 ();
 sg13g2_decap_8 FILLER_57_679 ();
 sg13g2_decap_8 FILLER_57_686 ();
 sg13g2_decap_8 FILLER_57_693 ();
 sg13g2_decap_8 FILLER_57_700 ();
 sg13g2_decap_8 FILLER_57_707 ();
 sg13g2_decap_8 FILLER_57_714 ();
 sg13g2_decap_8 FILLER_57_721 ();
 sg13g2_decap_8 FILLER_57_728 ();
 sg13g2_decap_8 FILLER_57_735 ();
 sg13g2_decap_8 FILLER_57_742 ();
 sg13g2_decap_8 FILLER_57_749 ();
 sg13g2_decap_8 FILLER_57_756 ();
 sg13g2_decap_8 FILLER_57_763 ();
 sg13g2_decap_8 FILLER_57_770 ();
 sg13g2_decap_8 FILLER_57_777 ();
 sg13g2_decap_8 FILLER_57_784 ();
 sg13g2_decap_8 FILLER_57_791 ();
 sg13g2_decap_8 FILLER_57_798 ();
 sg13g2_decap_8 FILLER_57_805 ();
 sg13g2_decap_8 FILLER_57_812 ();
 sg13g2_decap_8 FILLER_57_819 ();
 sg13g2_decap_8 FILLER_57_826 ();
 sg13g2_decap_8 FILLER_57_833 ();
 sg13g2_decap_8 FILLER_57_840 ();
 sg13g2_decap_8 FILLER_57_847 ();
 sg13g2_decap_8 FILLER_57_854 ();
 sg13g2_decap_8 FILLER_57_861 ();
 sg13g2_decap_8 FILLER_57_868 ();
 sg13g2_decap_8 FILLER_57_875 ();
 sg13g2_decap_8 FILLER_57_882 ();
 sg13g2_decap_8 FILLER_57_889 ();
 sg13g2_decap_8 FILLER_57_896 ();
 sg13g2_decap_8 FILLER_57_903 ();
 sg13g2_decap_8 FILLER_57_910 ();
 sg13g2_decap_8 FILLER_57_917 ();
 sg13g2_decap_8 FILLER_57_924 ();
 sg13g2_decap_8 FILLER_57_931 ();
 sg13g2_decap_8 FILLER_57_938 ();
 sg13g2_decap_8 FILLER_57_945 ();
 sg13g2_decap_8 FILLER_57_952 ();
 sg13g2_decap_8 FILLER_57_959 ();
 sg13g2_decap_8 FILLER_57_966 ();
 sg13g2_decap_8 FILLER_57_973 ();
 sg13g2_decap_8 FILLER_57_980 ();
 sg13g2_decap_8 FILLER_57_987 ();
 sg13g2_decap_8 FILLER_57_994 ();
 sg13g2_decap_8 FILLER_57_1001 ();
 sg13g2_decap_8 FILLER_57_1008 ();
 sg13g2_decap_8 FILLER_57_1015 ();
 sg13g2_decap_8 FILLER_57_1022 ();
 sg13g2_decap_8 FILLER_57_1029 ();
 sg13g2_decap_8 FILLER_57_1036 ();
 sg13g2_decap_8 FILLER_57_1043 ();
 sg13g2_decap_8 FILLER_57_1050 ();
 sg13g2_decap_8 FILLER_57_1057 ();
 sg13g2_decap_8 FILLER_57_1064 ();
 sg13g2_decap_8 FILLER_57_1071 ();
 sg13g2_decap_8 FILLER_57_1078 ();
 sg13g2_decap_8 FILLER_57_1085 ();
 sg13g2_decap_8 FILLER_57_1092 ();
 sg13g2_decap_8 FILLER_57_1099 ();
 sg13g2_decap_8 FILLER_57_1106 ();
 sg13g2_decap_8 FILLER_57_1113 ();
 sg13g2_decap_8 FILLER_57_1120 ();
 sg13g2_decap_8 FILLER_57_1127 ();
 sg13g2_decap_8 FILLER_57_1134 ();
 sg13g2_decap_8 FILLER_57_1141 ();
 sg13g2_decap_8 FILLER_57_1148 ();
 sg13g2_decap_8 FILLER_57_1155 ();
 sg13g2_decap_8 FILLER_57_1162 ();
 sg13g2_decap_8 FILLER_57_1169 ();
 sg13g2_decap_8 FILLER_57_1176 ();
 sg13g2_decap_8 FILLER_57_1183 ();
 sg13g2_decap_8 FILLER_57_1190 ();
 sg13g2_decap_8 FILLER_57_1197 ();
 sg13g2_decap_8 FILLER_57_1204 ();
 sg13g2_decap_8 FILLER_57_1211 ();
 sg13g2_decap_8 FILLER_57_1218 ();
 sg13g2_decap_8 FILLER_57_1225 ();
 sg13g2_decap_8 FILLER_57_1232 ();
 sg13g2_decap_8 FILLER_57_1239 ();
 sg13g2_decap_8 FILLER_57_1246 ();
 sg13g2_decap_8 FILLER_57_1253 ();
 sg13g2_decap_8 FILLER_57_1260 ();
 sg13g2_decap_8 FILLER_57_1267 ();
 sg13g2_decap_8 FILLER_57_1274 ();
 sg13g2_decap_8 FILLER_57_1281 ();
 sg13g2_decap_8 FILLER_57_1288 ();
 sg13g2_decap_8 FILLER_57_1295 ();
 sg13g2_decap_8 FILLER_57_1302 ();
 sg13g2_decap_8 FILLER_57_1309 ();
 sg13g2_decap_8 FILLER_57_1316 ();
 sg13g2_decap_8 FILLER_57_1323 ();
 sg13g2_decap_8 FILLER_57_1330 ();
 sg13g2_decap_8 FILLER_57_1337 ();
 sg13g2_decap_8 FILLER_57_1344 ();
 sg13g2_decap_8 FILLER_57_1351 ();
 sg13g2_decap_8 FILLER_57_1358 ();
 sg13g2_decap_8 FILLER_57_1365 ();
 sg13g2_decap_8 FILLER_57_1372 ();
 sg13g2_decap_8 FILLER_57_1379 ();
 sg13g2_decap_8 FILLER_57_1386 ();
 sg13g2_decap_8 FILLER_57_1393 ();
 sg13g2_decap_8 FILLER_57_1400 ();
 sg13g2_decap_8 FILLER_57_1407 ();
 sg13g2_decap_8 FILLER_57_1414 ();
 sg13g2_decap_8 FILLER_57_1421 ();
 sg13g2_decap_8 FILLER_57_1428 ();
 sg13g2_decap_8 FILLER_57_1435 ();
 sg13g2_decap_8 FILLER_57_1442 ();
 sg13g2_decap_8 FILLER_57_1449 ();
 sg13g2_decap_8 FILLER_57_1456 ();
 sg13g2_decap_8 FILLER_57_1463 ();
 sg13g2_decap_8 FILLER_57_1470 ();
 sg13g2_decap_8 FILLER_57_1477 ();
 sg13g2_decap_8 FILLER_57_1484 ();
 sg13g2_decap_8 FILLER_57_1491 ();
 sg13g2_decap_8 FILLER_57_1498 ();
 sg13g2_decap_8 FILLER_57_1505 ();
 sg13g2_decap_8 FILLER_57_1512 ();
 sg13g2_decap_8 FILLER_57_1519 ();
 sg13g2_decap_8 FILLER_57_1526 ();
 sg13g2_decap_8 FILLER_57_1533 ();
 sg13g2_decap_8 FILLER_57_1540 ();
 sg13g2_decap_8 FILLER_57_1547 ();
 sg13g2_decap_8 FILLER_57_1554 ();
 sg13g2_decap_8 FILLER_57_1561 ();
 sg13g2_decap_8 FILLER_57_1568 ();
 sg13g2_decap_8 FILLER_57_1575 ();
 sg13g2_decap_8 FILLER_57_1582 ();
 sg13g2_decap_8 FILLER_57_1589 ();
 sg13g2_decap_8 FILLER_57_1596 ();
 sg13g2_decap_8 FILLER_57_1603 ();
 sg13g2_decap_8 FILLER_57_1610 ();
 sg13g2_decap_8 FILLER_57_1617 ();
 sg13g2_decap_8 FILLER_57_1624 ();
 sg13g2_decap_8 FILLER_57_1631 ();
 sg13g2_decap_8 FILLER_57_1638 ();
 sg13g2_decap_8 FILLER_57_1645 ();
 sg13g2_decap_8 FILLER_57_1652 ();
 sg13g2_decap_8 FILLER_57_1659 ();
 sg13g2_decap_8 FILLER_57_1666 ();
 sg13g2_decap_8 FILLER_57_1673 ();
 sg13g2_decap_8 FILLER_57_1680 ();
 sg13g2_decap_8 FILLER_57_1687 ();
 sg13g2_decap_8 FILLER_57_1694 ();
 sg13g2_decap_8 FILLER_57_1701 ();
 sg13g2_decap_8 FILLER_57_1708 ();
 sg13g2_decap_8 FILLER_57_1715 ();
 sg13g2_decap_8 FILLER_57_1722 ();
 sg13g2_decap_8 FILLER_57_1729 ();
 sg13g2_decap_8 FILLER_57_1736 ();
 sg13g2_decap_8 FILLER_57_1743 ();
 sg13g2_decap_8 FILLER_57_1750 ();
 sg13g2_decap_8 FILLER_57_1757 ();
 sg13g2_decap_8 FILLER_57_1764 ();
 sg13g2_decap_8 FILLER_57_1771 ();
 sg13g2_decap_8 FILLER_57_1778 ();
 sg13g2_decap_8 FILLER_57_1785 ();
 sg13g2_decap_8 FILLER_57_1792 ();
 sg13g2_decap_8 FILLER_57_1799 ();
 sg13g2_decap_8 FILLER_57_1806 ();
 sg13g2_decap_8 FILLER_57_1813 ();
 sg13g2_decap_8 FILLER_57_1820 ();
 sg13g2_decap_8 FILLER_57_1827 ();
 sg13g2_decap_8 FILLER_57_1834 ();
 sg13g2_decap_8 FILLER_57_1841 ();
 sg13g2_decap_8 FILLER_57_1848 ();
 sg13g2_decap_8 FILLER_57_1855 ();
 sg13g2_decap_8 FILLER_57_1862 ();
 sg13g2_decap_8 FILLER_57_1869 ();
 sg13g2_decap_8 FILLER_57_1876 ();
 sg13g2_decap_8 FILLER_57_1883 ();
 sg13g2_decap_8 FILLER_57_1890 ();
 sg13g2_decap_8 FILLER_57_1897 ();
 sg13g2_decap_8 FILLER_57_1904 ();
 sg13g2_decap_8 FILLER_57_1911 ();
 sg13g2_decap_8 FILLER_57_1918 ();
 sg13g2_decap_8 FILLER_57_1925 ();
 sg13g2_decap_8 FILLER_57_1932 ();
 sg13g2_decap_8 FILLER_57_1939 ();
 sg13g2_decap_8 FILLER_57_1946 ();
 sg13g2_decap_8 FILLER_57_1953 ();
 sg13g2_decap_8 FILLER_57_1960 ();
 sg13g2_decap_8 FILLER_57_1967 ();
 sg13g2_decap_8 FILLER_57_1974 ();
 sg13g2_decap_8 FILLER_57_1981 ();
 sg13g2_decap_8 FILLER_57_1988 ();
 sg13g2_decap_8 FILLER_57_1995 ();
 sg13g2_decap_8 FILLER_57_2002 ();
 sg13g2_decap_8 FILLER_57_2009 ();
 sg13g2_decap_8 FILLER_57_2016 ();
 sg13g2_decap_8 FILLER_57_2023 ();
 sg13g2_decap_8 FILLER_57_2030 ();
 sg13g2_decap_8 FILLER_57_2037 ();
 sg13g2_decap_8 FILLER_57_2044 ();
 sg13g2_decap_8 FILLER_57_2051 ();
 sg13g2_decap_8 FILLER_57_2058 ();
 sg13g2_decap_8 FILLER_57_2065 ();
 sg13g2_decap_8 FILLER_57_2072 ();
 sg13g2_decap_8 FILLER_57_2079 ();
 sg13g2_decap_8 FILLER_57_2086 ();
 sg13g2_decap_8 FILLER_57_2093 ();
 sg13g2_decap_8 FILLER_57_2100 ();
 sg13g2_decap_8 FILLER_57_2107 ();
 sg13g2_decap_8 FILLER_57_2114 ();
 sg13g2_decap_8 FILLER_57_2121 ();
 sg13g2_decap_8 FILLER_57_2128 ();
 sg13g2_decap_8 FILLER_57_2135 ();
 sg13g2_decap_8 FILLER_57_2142 ();
 sg13g2_decap_8 FILLER_57_2149 ();
 sg13g2_decap_8 FILLER_57_2156 ();
 sg13g2_decap_8 FILLER_57_2163 ();
 sg13g2_decap_8 FILLER_57_2170 ();
 sg13g2_decap_8 FILLER_57_2177 ();
 sg13g2_decap_8 FILLER_57_2184 ();
 sg13g2_decap_8 FILLER_57_2191 ();
 sg13g2_decap_8 FILLER_57_2198 ();
 sg13g2_decap_8 FILLER_57_2205 ();
 sg13g2_decap_8 FILLER_57_2212 ();
 sg13g2_decap_8 FILLER_57_2219 ();
 sg13g2_decap_8 FILLER_57_2226 ();
 sg13g2_decap_8 FILLER_57_2233 ();
 sg13g2_decap_8 FILLER_57_2240 ();
 sg13g2_decap_8 FILLER_57_2247 ();
 sg13g2_decap_8 FILLER_57_2254 ();
 sg13g2_decap_8 FILLER_57_2261 ();
 sg13g2_decap_8 FILLER_57_2268 ();
 sg13g2_decap_8 FILLER_57_2275 ();
 sg13g2_decap_8 FILLER_57_2282 ();
 sg13g2_decap_8 FILLER_57_2289 ();
 sg13g2_decap_8 FILLER_57_2296 ();
 sg13g2_decap_8 FILLER_57_2303 ();
 sg13g2_decap_8 FILLER_57_2310 ();
 sg13g2_decap_8 FILLER_57_2317 ();
 sg13g2_decap_8 FILLER_57_2324 ();
 sg13g2_decap_8 FILLER_57_2331 ();
 sg13g2_decap_8 FILLER_57_2338 ();
 sg13g2_decap_8 FILLER_57_2345 ();
 sg13g2_decap_8 FILLER_57_2352 ();
 sg13g2_decap_8 FILLER_57_2359 ();
 sg13g2_decap_8 FILLER_57_2366 ();
 sg13g2_decap_8 FILLER_57_2373 ();
 sg13g2_decap_8 FILLER_57_2380 ();
 sg13g2_decap_8 FILLER_57_2387 ();
 sg13g2_decap_8 FILLER_57_2394 ();
 sg13g2_decap_8 FILLER_57_2401 ();
 sg13g2_decap_8 FILLER_57_2408 ();
 sg13g2_decap_8 FILLER_57_2415 ();
 sg13g2_decap_8 FILLER_57_2422 ();
 sg13g2_decap_8 FILLER_57_2429 ();
 sg13g2_decap_8 FILLER_57_2436 ();
 sg13g2_decap_8 FILLER_57_2443 ();
 sg13g2_decap_8 FILLER_57_2450 ();
 sg13g2_decap_8 FILLER_57_2457 ();
 sg13g2_decap_8 FILLER_57_2464 ();
 sg13g2_decap_8 FILLER_57_2471 ();
 sg13g2_decap_8 FILLER_57_2478 ();
 sg13g2_decap_8 FILLER_57_2485 ();
 sg13g2_decap_8 FILLER_57_2492 ();
 sg13g2_decap_8 FILLER_57_2499 ();
 sg13g2_decap_8 FILLER_57_2506 ();
 sg13g2_decap_8 FILLER_57_2513 ();
 sg13g2_decap_8 FILLER_57_2520 ();
 sg13g2_decap_8 FILLER_57_2527 ();
 sg13g2_decap_8 FILLER_57_2534 ();
 sg13g2_decap_8 FILLER_57_2541 ();
 sg13g2_decap_8 FILLER_57_2548 ();
 sg13g2_decap_8 FILLER_57_2555 ();
 sg13g2_decap_8 FILLER_57_2562 ();
 sg13g2_decap_8 FILLER_57_2569 ();
 sg13g2_decap_8 FILLER_57_2576 ();
 sg13g2_decap_8 FILLER_57_2583 ();
 sg13g2_decap_8 FILLER_57_2590 ();
 sg13g2_decap_8 FILLER_57_2597 ();
 sg13g2_decap_8 FILLER_57_2604 ();
 sg13g2_decap_8 FILLER_57_2611 ();
 sg13g2_decap_8 FILLER_57_2618 ();
 sg13g2_decap_8 FILLER_57_2625 ();
 sg13g2_decap_8 FILLER_57_2632 ();
 sg13g2_decap_8 FILLER_57_2639 ();
 sg13g2_decap_8 FILLER_57_2646 ();
 sg13g2_decap_8 FILLER_57_2653 ();
 sg13g2_decap_8 FILLER_57_2660 ();
 sg13g2_decap_8 FILLER_57_2667 ();
 sg13g2_decap_8 FILLER_57_2674 ();
 sg13g2_decap_8 FILLER_57_2681 ();
 sg13g2_decap_8 FILLER_57_2688 ();
 sg13g2_decap_8 FILLER_57_2695 ();
 sg13g2_decap_8 FILLER_57_2702 ();
 sg13g2_decap_8 FILLER_57_2709 ();
 sg13g2_decap_8 FILLER_57_2716 ();
 sg13g2_decap_8 FILLER_57_2723 ();
 sg13g2_decap_8 FILLER_57_2730 ();
 sg13g2_decap_8 FILLER_57_2737 ();
 sg13g2_decap_8 FILLER_57_2744 ();
 sg13g2_decap_8 FILLER_57_2751 ();
 sg13g2_decap_8 FILLER_57_2758 ();
 sg13g2_decap_8 FILLER_57_2765 ();
 sg13g2_decap_8 FILLER_57_2772 ();
 sg13g2_decap_8 FILLER_57_2779 ();
 sg13g2_decap_8 FILLER_57_2786 ();
 sg13g2_decap_8 FILLER_57_2793 ();
 sg13g2_decap_8 FILLER_57_2800 ();
 sg13g2_decap_8 FILLER_57_2807 ();
 sg13g2_decap_8 FILLER_57_2814 ();
 sg13g2_decap_8 FILLER_57_2821 ();
 sg13g2_decap_8 FILLER_57_2828 ();
 sg13g2_decap_8 FILLER_57_2835 ();
 sg13g2_decap_8 FILLER_57_2842 ();
 sg13g2_decap_8 FILLER_57_2849 ();
 sg13g2_decap_8 FILLER_57_2856 ();
 sg13g2_decap_8 FILLER_57_2863 ();
 sg13g2_decap_8 FILLER_57_2870 ();
 sg13g2_decap_8 FILLER_57_2877 ();
 sg13g2_decap_8 FILLER_57_2884 ();
 sg13g2_decap_8 FILLER_57_2891 ();
 sg13g2_decap_8 FILLER_57_2898 ();
 sg13g2_decap_8 FILLER_57_2905 ();
 sg13g2_decap_8 FILLER_57_2912 ();
 sg13g2_decap_8 FILLER_57_2919 ();
 sg13g2_decap_8 FILLER_57_2926 ();
 sg13g2_decap_8 FILLER_57_2933 ();
 sg13g2_decap_8 FILLER_57_2940 ();
 sg13g2_decap_8 FILLER_57_2947 ();
 sg13g2_decap_8 FILLER_57_2954 ();
 sg13g2_decap_8 FILLER_57_2961 ();
 sg13g2_decap_8 FILLER_57_2968 ();
 sg13g2_decap_8 FILLER_57_2975 ();
 sg13g2_decap_8 FILLER_57_2982 ();
 sg13g2_decap_8 FILLER_57_2989 ();
 sg13g2_decap_8 FILLER_57_2996 ();
 sg13g2_decap_8 FILLER_57_3003 ();
 sg13g2_decap_8 FILLER_57_3010 ();
 sg13g2_decap_8 FILLER_57_3017 ();
 sg13g2_decap_8 FILLER_57_3024 ();
 sg13g2_decap_8 FILLER_57_3031 ();
 sg13g2_decap_8 FILLER_57_3038 ();
 sg13g2_decap_8 FILLER_57_3045 ();
 sg13g2_decap_8 FILLER_57_3052 ();
 sg13g2_decap_8 FILLER_57_3059 ();
 sg13g2_decap_8 FILLER_57_3066 ();
 sg13g2_decap_8 FILLER_57_3073 ();
 sg13g2_decap_8 FILLER_57_3080 ();
 sg13g2_decap_8 FILLER_57_3087 ();
 sg13g2_decap_8 FILLER_57_3094 ();
 sg13g2_decap_8 FILLER_57_3101 ();
 sg13g2_decap_8 FILLER_57_3108 ();
 sg13g2_decap_8 FILLER_57_3115 ();
 sg13g2_decap_8 FILLER_57_3122 ();
 sg13g2_decap_8 FILLER_57_3129 ();
 sg13g2_decap_8 FILLER_57_3136 ();
 sg13g2_decap_8 FILLER_57_3143 ();
 sg13g2_decap_8 FILLER_57_3150 ();
 sg13g2_decap_8 FILLER_57_3157 ();
 sg13g2_decap_8 FILLER_57_3164 ();
 sg13g2_decap_8 FILLER_57_3171 ();
 sg13g2_decap_8 FILLER_57_3178 ();
 sg13g2_decap_8 FILLER_57_3185 ();
 sg13g2_decap_8 FILLER_57_3192 ();
 sg13g2_decap_8 FILLER_57_3199 ();
 sg13g2_decap_8 FILLER_57_3206 ();
 sg13g2_decap_8 FILLER_57_3213 ();
 sg13g2_decap_8 FILLER_57_3220 ();
 sg13g2_decap_8 FILLER_57_3227 ();
 sg13g2_decap_8 FILLER_57_3234 ();
 sg13g2_decap_8 FILLER_57_3241 ();
 sg13g2_decap_8 FILLER_57_3248 ();
 sg13g2_decap_8 FILLER_57_3255 ();
 sg13g2_decap_8 FILLER_57_3262 ();
 sg13g2_decap_8 FILLER_57_3269 ();
 sg13g2_decap_8 FILLER_57_3276 ();
 sg13g2_decap_8 FILLER_57_3283 ();
 sg13g2_decap_8 FILLER_57_3290 ();
 sg13g2_decap_8 FILLER_57_3297 ();
 sg13g2_decap_8 FILLER_57_3304 ();
 sg13g2_decap_8 FILLER_57_3311 ();
 sg13g2_decap_8 FILLER_57_3318 ();
 sg13g2_decap_8 FILLER_57_3325 ();
 sg13g2_decap_8 FILLER_57_3332 ();
 sg13g2_decap_8 FILLER_57_3339 ();
 sg13g2_decap_8 FILLER_57_3346 ();
 sg13g2_decap_8 FILLER_57_3353 ();
 sg13g2_decap_8 FILLER_57_3360 ();
 sg13g2_decap_8 FILLER_57_3367 ();
 sg13g2_decap_8 FILLER_57_3374 ();
 sg13g2_decap_8 FILLER_57_3381 ();
 sg13g2_decap_8 FILLER_57_3388 ();
 sg13g2_decap_8 FILLER_57_3395 ();
 sg13g2_decap_8 FILLER_57_3402 ();
 sg13g2_decap_8 FILLER_57_3409 ();
 sg13g2_decap_8 FILLER_57_3416 ();
 sg13g2_decap_8 FILLER_57_3423 ();
 sg13g2_decap_8 FILLER_57_3430 ();
 sg13g2_decap_8 FILLER_57_3437 ();
 sg13g2_decap_8 FILLER_57_3444 ();
 sg13g2_decap_8 FILLER_57_3451 ();
 sg13g2_decap_8 FILLER_57_3458 ();
 sg13g2_decap_8 FILLER_57_3465 ();
 sg13g2_decap_8 FILLER_57_3472 ();
 sg13g2_decap_8 FILLER_57_3479 ();
 sg13g2_decap_8 FILLER_57_3486 ();
 sg13g2_decap_8 FILLER_57_3493 ();
 sg13g2_decap_8 FILLER_57_3500 ();
 sg13g2_decap_8 FILLER_57_3507 ();
 sg13g2_decap_8 FILLER_57_3514 ();
 sg13g2_decap_8 FILLER_57_3521 ();
 sg13g2_decap_8 FILLER_57_3528 ();
 sg13g2_decap_8 FILLER_57_3535 ();
 sg13g2_decap_8 FILLER_57_3542 ();
 sg13g2_decap_8 FILLER_57_3549 ();
 sg13g2_decap_8 FILLER_57_3556 ();
 sg13g2_decap_8 FILLER_57_3563 ();
 sg13g2_decap_8 FILLER_57_3570 ();
 sg13g2_fill_2 FILLER_57_3577 ();
 sg13g2_fill_1 FILLER_57_3579 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_decap_8 FILLER_58_112 ();
 sg13g2_decap_8 FILLER_58_119 ();
 sg13g2_decap_8 FILLER_58_126 ();
 sg13g2_decap_8 FILLER_58_133 ();
 sg13g2_decap_8 FILLER_58_140 ();
 sg13g2_decap_8 FILLER_58_147 ();
 sg13g2_decap_8 FILLER_58_154 ();
 sg13g2_decap_8 FILLER_58_161 ();
 sg13g2_decap_8 FILLER_58_168 ();
 sg13g2_decap_8 FILLER_58_175 ();
 sg13g2_decap_8 FILLER_58_182 ();
 sg13g2_decap_8 FILLER_58_189 ();
 sg13g2_decap_8 FILLER_58_196 ();
 sg13g2_decap_8 FILLER_58_203 ();
 sg13g2_decap_8 FILLER_58_210 ();
 sg13g2_decap_8 FILLER_58_217 ();
 sg13g2_decap_8 FILLER_58_224 ();
 sg13g2_decap_8 FILLER_58_231 ();
 sg13g2_decap_8 FILLER_58_238 ();
 sg13g2_decap_8 FILLER_58_245 ();
 sg13g2_decap_8 FILLER_58_252 ();
 sg13g2_decap_8 FILLER_58_259 ();
 sg13g2_decap_8 FILLER_58_266 ();
 sg13g2_decap_8 FILLER_58_273 ();
 sg13g2_decap_8 FILLER_58_280 ();
 sg13g2_decap_8 FILLER_58_287 ();
 sg13g2_decap_8 FILLER_58_294 ();
 sg13g2_decap_8 FILLER_58_301 ();
 sg13g2_decap_8 FILLER_58_308 ();
 sg13g2_decap_8 FILLER_58_315 ();
 sg13g2_decap_8 FILLER_58_322 ();
 sg13g2_decap_8 FILLER_58_329 ();
 sg13g2_decap_8 FILLER_58_336 ();
 sg13g2_decap_8 FILLER_58_343 ();
 sg13g2_decap_8 FILLER_58_350 ();
 sg13g2_decap_8 FILLER_58_357 ();
 sg13g2_decap_8 FILLER_58_364 ();
 sg13g2_decap_8 FILLER_58_371 ();
 sg13g2_decap_8 FILLER_58_378 ();
 sg13g2_decap_8 FILLER_58_385 ();
 sg13g2_decap_8 FILLER_58_392 ();
 sg13g2_decap_8 FILLER_58_399 ();
 sg13g2_decap_8 FILLER_58_406 ();
 sg13g2_decap_8 FILLER_58_413 ();
 sg13g2_decap_8 FILLER_58_420 ();
 sg13g2_decap_8 FILLER_58_427 ();
 sg13g2_decap_8 FILLER_58_434 ();
 sg13g2_decap_8 FILLER_58_441 ();
 sg13g2_decap_8 FILLER_58_448 ();
 sg13g2_decap_8 FILLER_58_455 ();
 sg13g2_decap_8 FILLER_58_462 ();
 sg13g2_decap_8 FILLER_58_469 ();
 sg13g2_decap_8 FILLER_58_476 ();
 sg13g2_decap_8 FILLER_58_483 ();
 sg13g2_decap_8 FILLER_58_490 ();
 sg13g2_decap_8 FILLER_58_497 ();
 sg13g2_decap_8 FILLER_58_504 ();
 sg13g2_decap_8 FILLER_58_511 ();
 sg13g2_decap_8 FILLER_58_518 ();
 sg13g2_decap_8 FILLER_58_525 ();
 sg13g2_decap_8 FILLER_58_532 ();
 sg13g2_decap_8 FILLER_58_539 ();
 sg13g2_decap_8 FILLER_58_546 ();
 sg13g2_decap_8 FILLER_58_553 ();
 sg13g2_decap_8 FILLER_58_560 ();
 sg13g2_decap_8 FILLER_58_567 ();
 sg13g2_decap_8 FILLER_58_574 ();
 sg13g2_decap_8 FILLER_58_581 ();
 sg13g2_decap_8 FILLER_58_588 ();
 sg13g2_decap_8 FILLER_58_595 ();
 sg13g2_decap_8 FILLER_58_602 ();
 sg13g2_decap_8 FILLER_58_609 ();
 sg13g2_decap_8 FILLER_58_616 ();
 sg13g2_decap_8 FILLER_58_623 ();
 sg13g2_decap_8 FILLER_58_630 ();
 sg13g2_decap_8 FILLER_58_637 ();
 sg13g2_decap_8 FILLER_58_644 ();
 sg13g2_decap_8 FILLER_58_651 ();
 sg13g2_decap_8 FILLER_58_658 ();
 sg13g2_decap_8 FILLER_58_665 ();
 sg13g2_decap_8 FILLER_58_672 ();
 sg13g2_decap_8 FILLER_58_679 ();
 sg13g2_decap_8 FILLER_58_686 ();
 sg13g2_decap_8 FILLER_58_693 ();
 sg13g2_decap_8 FILLER_58_700 ();
 sg13g2_decap_8 FILLER_58_707 ();
 sg13g2_decap_8 FILLER_58_714 ();
 sg13g2_decap_8 FILLER_58_721 ();
 sg13g2_decap_8 FILLER_58_728 ();
 sg13g2_decap_8 FILLER_58_735 ();
 sg13g2_decap_8 FILLER_58_742 ();
 sg13g2_decap_8 FILLER_58_749 ();
 sg13g2_decap_8 FILLER_58_756 ();
 sg13g2_decap_8 FILLER_58_763 ();
 sg13g2_decap_8 FILLER_58_770 ();
 sg13g2_decap_8 FILLER_58_777 ();
 sg13g2_decap_8 FILLER_58_784 ();
 sg13g2_decap_8 FILLER_58_791 ();
 sg13g2_decap_8 FILLER_58_798 ();
 sg13g2_decap_8 FILLER_58_805 ();
 sg13g2_decap_8 FILLER_58_812 ();
 sg13g2_decap_8 FILLER_58_819 ();
 sg13g2_decap_8 FILLER_58_826 ();
 sg13g2_decap_8 FILLER_58_833 ();
 sg13g2_decap_8 FILLER_58_840 ();
 sg13g2_decap_8 FILLER_58_847 ();
 sg13g2_decap_8 FILLER_58_854 ();
 sg13g2_decap_8 FILLER_58_861 ();
 sg13g2_decap_8 FILLER_58_868 ();
 sg13g2_decap_8 FILLER_58_875 ();
 sg13g2_decap_8 FILLER_58_882 ();
 sg13g2_decap_8 FILLER_58_889 ();
 sg13g2_decap_8 FILLER_58_896 ();
 sg13g2_decap_8 FILLER_58_903 ();
 sg13g2_decap_8 FILLER_58_910 ();
 sg13g2_decap_8 FILLER_58_917 ();
 sg13g2_decap_8 FILLER_58_924 ();
 sg13g2_decap_8 FILLER_58_931 ();
 sg13g2_decap_8 FILLER_58_938 ();
 sg13g2_decap_8 FILLER_58_945 ();
 sg13g2_decap_8 FILLER_58_952 ();
 sg13g2_decap_8 FILLER_58_959 ();
 sg13g2_decap_8 FILLER_58_966 ();
 sg13g2_decap_8 FILLER_58_973 ();
 sg13g2_decap_8 FILLER_58_980 ();
 sg13g2_decap_8 FILLER_58_987 ();
 sg13g2_decap_8 FILLER_58_994 ();
 sg13g2_decap_8 FILLER_58_1001 ();
 sg13g2_decap_8 FILLER_58_1008 ();
 sg13g2_decap_8 FILLER_58_1015 ();
 sg13g2_decap_8 FILLER_58_1022 ();
 sg13g2_decap_8 FILLER_58_1029 ();
 sg13g2_decap_8 FILLER_58_1036 ();
 sg13g2_decap_8 FILLER_58_1043 ();
 sg13g2_decap_8 FILLER_58_1050 ();
 sg13g2_decap_8 FILLER_58_1057 ();
 sg13g2_decap_8 FILLER_58_1064 ();
 sg13g2_decap_8 FILLER_58_1071 ();
 sg13g2_decap_8 FILLER_58_1078 ();
 sg13g2_decap_8 FILLER_58_1085 ();
 sg13g2_decap_8 FILLER_58_1092 ();
 sg13g2_decap_8 FILLER_58_1099 ();
 sg13g2_decap_8 FILLER_58_1106 ();
 sg13g2_decap_8 FILLER_58_1113 ();
 sg13g2_decap_8 FILLER_58_1120 ();
 sg13g2_decap_8 FILLER_58_1127 ();
 sg13g2_decap_8 FILLER_58_1134 ();
 sg13g2_decap_8 FILLER_58_1141 ();
 sg13g2_decap_8 FILLER_58_1148 ();
 sg13g2_decap_8 FILLER_58_1155 ();
 sg13g2_decap_8 FILLER_58_1162 ();
 sg13g2_decap_8 FILLER_58_1169 ();
 sg13g2_decap_8 FILLER_58_1176 ();
 sg13g2_decap_8 FILLER_58_1183 ();
 sg13g2_decap_8 FILLER_58_1190 ();
 sg13g2_decap_8 FILLER_58_1197 ();
 sg13g2_decap_8 FILLER_58_1204 ();
 sg13g2_decap_8 FILLER_58_1211 ();
 sg13g2_decap_8 FILLER_58_1218 ();
 sg13g2_decap_8 FILLER_58_1225 ();
 sg13g2_decap_8 FILLER_58_1232 ();
 sg13g2_decap_8 FILLER_58_1239 ();
 sg13g2_decap_8 FILLER_58_1246 ();
 sg13g2_decap_8 FILLER_58_1253 ();
 sg13g2_decap_8 FILLER_58_1260 ();
 sg13g2_decap_8 FILLER_58_1267 ();
 sg13g2_decap_8 FILLER_58_1274 ();
 sg13g2_decap_8 FILLER_58_1281 ();
 sg13g2_decap_8 FILLER_58_1288 ();
 sg13g2_decap_8 FILLER_58_1295 ();
 sg13g2_decap_8 FILLER_58_1302 ();
 sg13g2_decap_8 FILLER_58_1309 ();
 sg13g2_decap_8 FILLER_58_1316 ();
 sg13g2_decap_8 FILLER_58_1323 ();
 sg13g2_decap_8 FILLER_58_1330 ();
 sg13g2_decap_8 FILLER_58_1337 ();
 sg13g2_decap_8 FILLER_58_1344 ();
 sg13g2_decap_8 FILLER_58_1351 ();
 sg13g2_decap_8 FILLER_58_1358 ();
 sg13g2_decap_8 FILLER_58_1365 ();
 sg13g2_decap_8 FILLER_58_1372 ();
 sg13g2_decap_8 FILLER_58_1379 ();
 sg13g2_decap_8 FILLER_58_1386 ();
 sg13g2_decap_8 FILLER_58_1393 ();
 sg13g2_decap_8 FILLER_58_1400 ();
 sg13g2_decap_8 FILLER_58_1407 ();
 sg13g2_decap_8 FILLER_58_1414 ();
 sg13g2_decap_8 FILLER_58_1421 ();
 sg13g2_decap_8 FILLER_58_1428 ();
 sg13g2_decap_8 FILLER_58_1435 ();
 sg13g2_decap_8 FILLER_58_1442 ();
 sg13g2_decap_8 FILLER_58_1449 ();
 sg13g2_decap_8 FILLER_58_1456 ();
 sg13g2_decap_8 FILLER_58_1463 ();
 sg13g2_decap_8 FILLER_58_1470 ();
 sg13g2_decap_8 FILLER_58_1477 ();
 sg13g2_decap_8 FILLER_58_1484 ();
 sg13g2_decap_8 FILLER_58_1491 ();
 sg13g2_decap_8 FILLER_58_1498 ();
 sg13g2_decap_8 FILLER_58_1505 ();
 sg13g2_decap_8 FILLER_58_1512 ();
 sg13g2_decap_8 FILLER_58_1519 ();
 sg13g2_decap_8 FILLER_58_1526 ();
 sg13g2_decap_8 FILLER_58_1533 ();
 sg13g2_decap_8 FILLER_58_1540 ();
 sg13g2_decap_8 FILLER_58_1547 ();
 sg13g2_decap_8 FILLER_58_1554 ();
 sg13g2_decap_8 FILLER_58_1561 ();
 sg13g2_decap_8 FILLER_58_1568 ();
 sg13g2_decap_8 FILLER_58_1575 ();
 sg13g2_decap_8 FILLER_58_1582 ();
 sg13g2_decap_8 FILLER_58_1589 ();
 sg13g2_decap_8 FILLER_58_1596 ();
 sg13g2_decap_8 FILLER_58_1603 ();
 sg13g2_decap_8 FILLER_58_1610 ();
 sg13g2_decap_8 FILLER_58_1617 ();
 sg13g2_decap_8 FILLER_58_1624 ();
 sg13g2_decap_8 FILLER_58_1631 ();
 sg13g2_decap_8 FILLER_58_1638 ();
 sg13g2_decap_8 FILLER_58_1645 ();
 sg13g2_decap_8 FILLER_58_1652 ();
 sg13g2_decap_8 FILLER_58_1659 ();
 sg13g2_decap_8 FILLER_58_1666 ();
 sg13g2_decap_8 FILLER_58_1673 ();
 sg13g2_decap_8 FILLER_58_1680 ();
 sg13g2_decap_8 FILLER_58_1687 ();
 sg13g2_decap_8 FILLER_58_1694 ();
 sg13g2_decap_8 FILLER_58_1701 ();
 sg13g2_decap_8 FILLER_58_1708 ();
 sg13g2_decap_8 FILLER_58_1715 ();
 sg13g2_decap_8 FILLER_58_1722 ();
 sg13g2_decap_8 FILLER_58_1729 ();
 sg13g2_decap_8 FILLER_58_1736 ();
 sg13g2_decap_8 FILLER_58_1743 ();
 sg13g2_decap_8 FILLER_58_1750 ();
 sg13g2_decap_8 FILLER_58_1757 ();
 sg13g2_decap_8 FILLER_58_1764 ();
 sg13g2_decap_8 FILLER_58_1771 ();
 sg13g2_decap_8 FILLER_58_1778 ();
 sg13g2_decap_8 FILLER_58_1785 ();
 sg13g2_decap_8 FILLER_58_1792 ();
 sg13g2_decap_8 FILLER_58_1799 ();
 sg13g2_decap_8 FILLER_58_1806 ();
 sg13g2_decap_8 FILLER_58_1813 ();
 sg13g2_decap_8 FILLER_58_1820 ();
 sg13g2_decap_8 FILLER_58_1827 ();
 sg13g2_decap_8 FILLER_58_1834 ();
 sg13g2_decap_8 FILLER_58_1841 ();
 sg13g2_decap_8 FILLER_58_1848 ();
 sg13g2_decap_8 FILLER_58_1855 ();
 sg13g2_decap_8 FILLER_58_1862 ();
 sg13g2_decap_8 FILLER_58_1869 ();
 sg13g2_decap_8 FILLER_58_1876 ();
 sg13g2_decap_8 FILLER_58_1883 ();
 sg13g2_decap_8 FILLER_58_1890 ();
 sg13g2_decap_8 FILLER_58_1897 ();
 sg13g2_decap_8 FILLER_58_1904 ();
 sg13g2_decap_8 FILLER_58_1911 ();
 sg13g2_decap_8 FILLER_58_1918 ();
 sg13g2_decap_8 FILLER_58_1925 ();
 sg13g2_decap_8 FILLER_58_1932 ();
 sg13g2_decap_8 FILLER_58_1939 ();
 sg13g2_decap_8 FILLER_58_1946 ();
 sg13g2_decap_8 FILLER_58_1953 ();
 sg13g2_decap_8 FILLER_58_1960 ();
 sg13g2_decap_8 FILLER_58_1967 ();
 sg13g2_decap_8 FILLER_58_1974 ();
 sg13g2_decap_8 FILLER_58_1981 ();
 sg13g2_decap_8 FILLER_58_1988 ();
 sg13g2_decap_8 FILLER_58_1995 ();
 sg13g2_decap_8 FILLER_58_2002 ();
 sg13g2_decap_8 FILLER_58_2009 ();
 sg13g2_decap_8 FILLER_58_2016 ();
 sg13g2_decap_8 FILLER_58_2023 ();
 sg13g2_decap_8 FILLER_58_2030 ();
 sg13g2_decap_8 FILLER_58_2037 ();
 sg13g2_decap_8 FILLER_58_2044 ();
 sg13g2_decap_8 FILLER_58_2051 ();
 sg13g2_decap_8 FILLER_58_2058 ();
 sg13g2_decap_8 FILLER_58_2065 ();
 sg13g2_decap_8 FILLER_58_2072 ();
 sg13g2_decap_8 FILLER_58_2079 ();
 sg13g2_decap_8 FILLER_58_2086 ();
 sg13g2_decap_8 FILLER_58_2093 ();
 sg13g2_decap_8 FILLER_58_2100 ();
 sg13g2_decap_8 FILLER_58_2107 ();
 sg13g2_decap_8 FILLER_58_2114 ();
 sg13g2_decap_8 FILLER_58_2121 ();
 sg13g2_decap_8 FILLER_58_2128 ();
 sg13g2_decap_8 FILLER_58_2135 ();
 sg13g2_decap_8 FILLER_58_2142 ();
 sg13g2_decap_8 FILLER_58_2149 ();
 sg13g2_decap_8 FILLER_58_2156 ();
 sg13g2_decap_8 FILLER_58_2163 ();
 sg13g2_decap_8 FILLER_58_2170 ();
 sg13g2_decap_8 FILLER_58_2177 ();
 sg13g2_decap_8 FILLER_58_2184 ();
 sg13g2_decap_8 FILLER_58_2191 ();
 sg13g2_decap_8 FILLER_58_2198 ();
 sg13g2_decap_8 FILLER_58_2205 ();
 sg13g2_decap_8 FILLER_58_2212 ();
 sg13g2_decap_8 FILLER_58_2219 ();
 sg13g2_decap_8 FILLER_58_2226 ();
 sg13g2_decap_8 FILLER_58_2233 ();
 sg13g2_decap_8 FILLER_58_2240 ();
 sg13g2_decap_8 FILLER_58_2247 ();
 sg13g2_decap_8 FILLER_58_2254 ();
 sg13g2_decap_8 FILLER_58_2261 ();
 sg13g2_decap_8 FILLER_58_2268 ();
 sg13g2_decap_8 FILLER_58_2275 ();
 sg13g2_decap_8 FILLER_58_2282 ();
 sg13g2_decap_8 FILLER_58_2289 ();
 sg13g2_decap_8 FILLER_58_2296 ();
 sg13g2_decap_8 FILLER_58_2303 ();
 sg13g2_decap_8 FILLER_58_2310 ();
 sg13g2_decap_8 FILLER_58_2317 ();
 sg13g2_decap_8 FILLER_58_2324 ();
 sg13g2_decap_8 FILLER_58_2331 ();
 sg13g2_decap_8 FILLER_58_2338 ();
 sg13g2_decap_8 FILLER_58_2345 ();
 sg13g2_decap_8 FILLER_58_2352 ();
 sg13g2_decap_8 FILLER_58_2359 ();
 sg13g2_decap_8 FILLER_58_2366 ();
 sg13g2_decap_8 FILLER_58_2373 ();
 sg13g2_decap_8 FILLER_58_2380 ();
 sg13g2_decap_8 FILLER_58_2387 ();
 sg13g2_decap_8 FILLER_58_2394 ();
 sg13g2_decap_8 FILLER_58_2401 ();
 sg13g2_decap_8 FILLER_58_2408 ();
 sg13g2_decap_8 FILLER_58_2415 ();
 sg13g2_decap_8 FILLER_58_2422 ();
 sg13g2_decap_8 FILLER_58_2429 ();
 sg13g2_decap_8 FILLER_58_2436 ();
 sg13g2_decap_8 FILLER_58_2443 ();
 sg13g2_decap_8 FILLER_58_2450 ();
 sg13g2_decap_8 FILLER_58_2457 ();
 sg13g2_decap_8 FILLER_58_2464 ();
 sg13g2_decap_8 FILLER_58_2471 ();
 sg13g2_decap_8 FILLER_58_2478 ();
 sg13g2_decap_8 FILLER_58_2485 ();
 sg13g2_decap_8 FILLER_58_2492 ();
 sg13g2_decap_8 FILLER_58_2499 ();
 sg13g2_decap_8 FILLER_58_2506 ();
 sg13g2_decap_8 FILLER_58_2513 ();
 sg13g2_decap_8 FILLER_58_2520 ();
 sg13g2_decap_8 FILLER_58_2527 ();
 sg13g2_decap_8 FILLER_58_2534 ();
 sg13g2_decap_8 FILLER_58_2541 ();
 sg13g2_decap_8 FILLER_58_2548 ();
 sg13g2_decap_8 FILLER_58_2555 ();
 sg13g2_decap_8 FILLER_58_2562 ();
 sg13g2_decap_8 FILLER_58_2569 ();
 sg13g2_decap_8 FILLER_58_2576 ();
 sg13g2_decap_8 FILLER_58_2583 ();
 sg13g2_decap_8 FILLER_58_2590 ();
 sg13g2_decap_8 FILLER_58_2597 ();
 sg13g2_decap_8 FILLER_58_2604 ();
 sg13g2_decap_8 FILLER_58_2611 ();
 sg13g2_decap_8 FILLER_58_2618 ();
 sg13g2_decap_8 FILLER_58_2625 ();
 sg13g2_decap_8 FILLER_58_2632 ();
 sg13g2_decap_8 FILLER_58_2639 ();
 sg13g2_decap_8 FILLER_58_2646 ();
 sg13g2_decap_8 FILLER_58_2653 ();
 sg13g2_decap_8 FILLER_58_2660 ();
 sg13g2_decap_8 FILLER_58_2667 ();
 sg13g2_decap_8 FILLER_58_2674 ();
 sg13g2_decap_8 FILLER_58_2681 ();
 sg13g2_decap_8 FILLER_58_2688 ();
 sg13g2_decap_8 FILLER_58_2695 ();
 sg13g2_decap_8 FILLER_58_2702 ();
 sg13g2_decap_8 FILLER_58_2709 ();
 sg13g2_decap_8 FILLER_58_2716 ();
 sg13g2_decap_8 FILLER_58_2723 ();
 sg13g2_decap_8 FILLER_58_2730 ();
 sg13g2_decap_8 FILLER_58_2737 ();
 sg13g2_decap_8 FILLER_58_2744 ();
 sg13g2_decap_8 FILLER_58_2751 ();
 sg13g2_decap_8 FILLER_58_2758 ();
 sg13g2_decap_8 FILLER_58_2765 ();
 sg13g2_decap_8 FILLER_58_2772 ();
 sg13g2_decap_8 FILLER_58_2779 ();
 sg13g2_decap_8 FILLER_58_2786 ();
 sg13g2_decap_8 FILLER_58_2793 ();
 sg13g2_decap_8 FILLER_58_2800 ();
 sg13g2_decap_8 FILLER_58_2807 ();
 sg13g2_decap_8 FILLER_58_2814 ();
 sg13g2_decap_8 FILLER_58_2821 ();
 sg13g2_decap_8 FILLER_58_2828 ();
 sg13g2_decap_8 FILLER_58_2835 ();
 sg13g2_decap_8 FILLER_58_2842 ();
 sg13g2_decap_8 FILLER_58_2849 ();
 sg13g2_decap_8 FILLER_58_2856 ();
 sg13g2_decap_8 FILLER_58_2863 ();
 sg13g2_decap_8 FILLER_58_2870 ();
 sg13g2_decap_8 FILLER_58_2877 ();
 sg13g2_decap_8 FILLER_58_2884 ();
 sg13g2_decap_8 FILLER_58_2891 ();
 sg13g2_decap_8 FILLER_58_2898 ();
 sg13g2_decap_8 FILLER_58_2905 ();
 sg13g2_decap_8 FILLER_58_2912 ();
 sg13g2_decap_8 FILLER_58_2919 ();
 sg13g2_decap_8 FILLER_58_2926 ();
 sg13g2_decap_8 FILLER_58_2933 ();
 sg13g2_decap_8 FILLER_58_2940 ();
 sg13g2_decap_8 FILLER_58_2947 ();
 sg13g2_decap_8 FILLER_58_2954 ();
 sg13g2_decap_8 FILLER_58_2961 ();
 sg13g2_decap_8 FILLER_58_2968 ();
 sg13g2_decap_8 FILLER_58_2975 ();
 sg13g2_decap_8 FILLER_58_2982 ();
 sg13g2_decap_8 FILLER_58_2989 ();
 sg13g2_decap_8 FILLER_58_2996 ();
 sg13g2_decap_8 FILLER_58_3003 ();
 sg13g2_decap_8 FILLER_58_3010 ();
 sg13g2_decap_8 FILLER_58_3017 ();
 sg13g2_decap_8 FILLER_58_3024 ();
 sg13g2_decap_8 FILLER_58_3031 ();
 sg13g2_decap_8 FILLER_58_3038 ();
 sg13g2_decap_8 FILLER_58_3045 ();
 sg13g2_decap_8 FILLER_58_3052 ();
 sg13g2_decap_8 FILLER_58_3059 ();
 sg13g2_decap_8 FILLER_58_3066 ();
 sg13g2_decap_8 FILLER_58_3073 ();
 sg13g2_decap_8 FILLER_58_3080 ();
 sg13g2_decap_8 FILLER_58_3087 ();
 sg13g2_decap_8 FILLER_58_3094 ();
 sg13g2_decap_8 FILLER_58_3101 ();
 sg13g2_decap_8 FILLER_58_3108 ();
 sg13g2_decap_8 FILLER_58_3115 ();
 sg13g2_decap_8 FILLER_58_3122 ();
 sg13g2_decap_8 FILLER_58_3129 ();
 sg13g2_decap_8 FILLER_58_3136 ();
 sg13g2_decap_8 FILLER_58_3143 ();
 sg13g2_decap_8 FILLER_58_3150 ();
 sg13g2_decap_8 FILLER_58_3157 ();
 sg13g2_decap_8 FILLER_58_3164 ();
 sg13g2_decap_8 FILLER_58_3171 ();
 sg13g2_decap_8 FILLER_58_3178 ();
 sg13g2_decap_8 FILLER_58_3185 ();
 sg13g2_decap_8 FILLER_58_3192 ();
 sg13g2_decap_8 FILLER_58_3199 ();
 sg13g2_decap_8 FILLER_58_3206 ();
 sg13g2_decap_8 FILLER_58_3213 ();
 sg13g2_decap_8 FILLER_58_3220 ();
 sg13g2_decap_8 FILLER_58_3227 ();
 sg13g2_decap_8 FILLER_58_3234 ();
 sg13g2_decap_8 FILLER_58_3241 ();
 sg13g2_decap_8 FILLER_58_3248 ();
 sg13g2_decap_8 FILLER_58_3255 ();
 sg13g2_decap_8 FILLER_58_3262 ();
 sg13g2_decap_8 FILLER_58_3269 ();
 sg13g2_decap_8 FILLER_58_3276 ();
 sg13g2_decap_8 FILLER_58_3283 ();
 sg13g2_decap_8 FILLER_58_3290 ();
 sg13g2_decap_8 FILLER_58_3297 ();
 sg13g2_decap_8 FILLER_58_3304 ();
 sg13g2_decap_8 FILLER_58_3311 ();
 sg13g2_decap_8 FILLER_58_3318 ();
 sg13g2_decap_8 FILLER_58_3325 ();
 sg13g2_decap_8 FILLER_58_3332 ();
 sg13g2_decap_8 FILLER_58_3339 ();
 sg13g2_decap_8 FILLER_58_3346 ();
 sg13g2_decap_8 FILLER_58_3353 ();
 sg13g2_decap_8 FILLER_58_3360 ();
 sg13g2_decap_8 FILLER_58_3367 ();
 sg13g2_decap_8 FILLER_58_3374 ();
 sg13g2_decap_8 FILLER_58_3381 ();
 sg13g2_decap_8 FILLER_58_3388 ();
 sg13g2_decap_8 FILLER_58_3395 ();
 sg13g2_decap_8 FILLER_58_3402 ();
 sg13g2_decap_8 FILLER_58_3409 ();
 sg13g2_decap_8 FILLER_58_3416 ();
 sg13g2_decap_8 FILLER_58_3423 ();
 sg13g2_decap_8 FILLER_58_3430 ();
 sg13g2_decap_8 FILLER_58_3437 ();
 sg13g2_decap_8 FILLER_58_3444 ();
 sg13g2_decap_8 FILLER_58_3451 ();
 sg13g2_decap_8 FILLER_58_3458 ();
 sg13g2_decap_8 FILLER_58_3465 ();
 sg13g2_decap_8 FILLER_58_3472 ();
 sg13g2_decap_8 FILLER_58_3479 ();
 sg13g2_decap_8 FILLER_58_3486 ();
 sg13g2_decap_8 FILLER_58_3493 ();
 sg13g2_decap_8 FILLER_58_3500 ();
 sg13g2_decap_8 FILLER_58_3507 ();
 sg13g2_decap_8 FILLER_58_3514 ();
 sg13g2_decap_8 FILLER_58_3521 ();
 sg13g2_decap_8 FILLER_58_3528 ();
 sg13g2_decap_8 FILLER_58_3535 ();
 sg13g2_decap_8 FILLER_58_3542 ();
 sg13g2_decap_8 FILLER_58_3549 ();
 sg13g2_decap_8 FILLER_58_3556 ();
 sg13g2_decap_8 FILLER_58_3563 ();
 sg13g2_decap_8 FILLER_58_3570 ();
 sg13g2_fill_2 FILLER_58_3577 ();
 sg13g2_fill_1 FILLER_58_3579 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_decap_8 FILLER_59_105 ();
 sg13g2_decap_8 FILLER_59_112 ();
 sg13g2_decap_8 FILLER_59_119 ();
 sg13g2_decap_8 FILLER_59_126 ();
 sg13g2_decap_8 FILLER_59_133 ();
 sg13g2_decap_8 FILLER_59_140 ();
 sg13g2_decap_8 FILLER_59_147 ();
 sg13g2_decap_8 FILLER_59_154 ();
 sg13g2_decap_8 FILLER_59_161 ();
 sg13g2_decap_8 FILLER_59_168 ();
 sg13g2_decap_8 FILLER_59_175 ();
 sg13g2_decap_8 FILLER_59_182 ();
 sg13g2_decap_8 FILLER_59_189 ();
 sg13g2_decap_8 FILLER_59_196 ();
 sg13g2_decap_8 FILLER_59_203 ();
 sg13g2_decap_8 FILLER_59_210 ();
 sg13g2_decap_8 FILLER_59_217 ();
 sg13g2_decap_8 FILLER_59_224 ();
 sg13g2_decap_8 FILLER_59_231 ();
 sg13g2_decap_8 FILLER_59_238 ();
 sg13g2_decap_8 FILLER_59_245 ();
 sg13g2_decap_8 FILLER_59_252 ();
 sg13g2_decap_8 FILLER_59_259 ();
 sg13g2_decap_8 FILLER_59_266 ();
 sg13g2_decap_8 FILLER_59_273 ();
 sg13g2_decap_8 FILLER_59_280 ();
 sg13g2_decap_8 FILLER_59_287 ();
 sg13g2_decap_8 FILLER_59_294 ();
 sg13g2_decap_8 FILLER_59_301 ();
 sg13g2_decap_8 FILLER_59_308 ();
 sg13g2_decap_8 FILLER_59_315 ();
 sg13g2_decap_8 FILLER_59_322 ();
 sg13g2_decap_8 FILLER_59_329 ();
 sg13g2_decap_8 FILLER_59_336 ();
 sg13g2_decap_8 FILLER_59_343 ();
 sg13g2_decap_8 FILLER_59_350 ();
 sg13g2_decap_8 FILLER_59_357 ();
 sg13g2_decap_8 FILLER_59_364 ();
 sg13g2_decap_8 FILLER_59_371 ();
 sg13g2_decap_8 FILLER_59_378 ();
 sg13g2_decap_8 FILLER_59_385 ();
 sg13g2_decap_8 FILLER_59_392 ();
 sg13g2_decap_8 FILLER_59_399 ();
 sg13g2_decap_8 FILLER_59_406 ();
 sg13g2_decap_8 FILLER_59_413 ();
 sg13g2_decap_8 FILLER_59_420 ();
 sg13g2_decap_8 FILLER_59_427 ();
 sg13g2_decap_8 FILLER_59_434 ();
 sg13g2_decap_8 FILLER_59_441 ();
 sg13g2_decap_8 FILLER_59_448 ();
 sg13g2_decap_8 FILLER_59_455 ();
 sg13g2_decap_8 FILLER_59_462 ();
 sg13g2_decap_8 FILLER_59_469 ();
 sg13g2_decap_8 FILLER_59_476 ();
 sg13g2_decap_8 FILLER_59_483 ();
 sg13g2_decap_8 FILLER_59_490 ();
 sg13g2_decap_8 FILLER_59_497 ();
 sg13g2_decap_8 FILLER_59_504 ();
 sg13g2_decap_8 FILLER_59_511 ();
 sg13g2_decap_8 FILLER_59_518 ();
 sg13g2_decap_8 FILLER_59_525 ();
 sg13g2_decap_8 FILLER_59_532 ();
 sg13g2_decap_8 FILLER_59_539 ();
 sg13g2_decap_8 FILLER_59_546 ();
 sg13g2_decap_8 FILLER_59_553 ();
 sg13g2_decap_8 FILLER_59_560 ();
 sg13g2_decap_8 FILLER_59_567 ();
 sg13g2_decap_8 FILLER_59_574 ();
 sg13g2_decap_8 FILLER_59_581 ();
 sg13g2_decap_8 FILLER_59_588 ();
 sg13g2_decap_8 FILLER_59_595 ();
 sg13g2_decap_8 FILLER_59_602 ();
 sg13g2_decap_8 FILLER_59_609 ();
 sg13g2_decap_8 FILLER_59_616 ();
 sg13g2_decap_8 FILLER_59_623 ();
 sg13g2_decap_8 FILLER_59_630 ();
 sg13g2_decap_8 FILLER_59_637 ();
 sg13g2_decap_8 FILLER_59_644 ();
 sg13g2_decap_8 FILLER_59_651 ();
 sg13g2_decap_8 FILLER_59_658 ();
 sg13g2_decap_8 FILLER_59_665 ();
 sg13g2_decap_8 FILLER_59_672 ();
 sg13g2_decap_8 FILLER_59_679 ();
 sg13g2_decap_8 FILLER_59_686 ();
 sg13g2_decap_8 FILLER_59_693 ();
 sg13g2_decap_8 FILLER_59_700 ();
 sg13g2_decap_8 FILLER_59_707 ();
 sg13g2_decap_8 FILLER_59_714 ();
 sg13g2_decap_8 FILLER_59_721 ();
 sg13g2_decap_8 FILLER_59_728 ();
 sg13g2_decap_8 FILLER_59_735 ();
 sg13g2_decap_8 FILLER_59_742 ();
 sg13g2_decap_8 FILLER_59_749 ();
 sg13g2_decap_8 FILLER_59_756 ();
 sg13g2_decap_8 FILLER_59_763 ();
 sg13g2_decap_8 FILLER_59_770 ();
 sg13g2_decap_8 FILLER_59_777 ();
 sg13g2_decap_8 FILLER_59_784 ();
 sg13g2_decap_8 FILLER_59_791 ();
 sg13g2_decap_8 FILLER_59_798 ();
 sg13g2_decap_8 FILLER_59_805 ();
 sg13g2_decap_8 FILLER_59_812 ();
 sg13g2_decap_8 FILLER_59_819 ();
 sg13g2_decap_8 FILLER_59_826 ();
 sg13g2_decap_8 FILLER_59_833 ();
 sg13g2_decap_8 FILLER_59_840 ();
 sg13g2_decap_8 FILLER_59_847 ();
 sg13g2_decap_8 FILLER_59_854 ();
 sg13g2_decap_8 FILLER_59_861 ();
 sg13g2_decap_8 FILLER_59_868 ();
 sg13g2_decap_8 FILLER_59_875 ();
 sg13g2_decap_8 FILLER_59_882 ();
 sg13g2_decap_8 FILLER_59_889 ();
 sg13g2_decap_8 FILLER_59_896 ();
 sg13g2_decap_8 FILLER_59_903 ();
 sg13g2_decap_8 FILLER_59_910 ();
 sg13g2_decap_8 FILLER_59_917 ();
 sg13g2_decap_8 FILLER_59_924 ();
 sg13g2_decap_8 FILLER_59_931 ();
 sg13g2_decap_8 FILLER_59_938 ();
 sg13g2_decap_8 FILLER_59_945 ();
 sg13g2_decap_8 FILLER_59_952 ();
 sg13g2_decap_8 FILLER_59_959 ();
 sg13g2_decap_8 FILLER_59_966 ();
 sg13g2_decap_8 FILLER_59_973 ();
 sg13g2_decap_8 FILLER_59_980 ();
 sg13g2_decap_8 FILLER_59_987 ();
 sg13g2_decap_8 FILLER_59_994 ();
 sg13g2_decap_8 FILLER_59_1001 ();
 sg13g2_decap_8 FILLER_59_1008 ();
 sg13g2_decap_8 FILLER_59_1015 ();
 sg13g2_decap_8 FILLER_59_1022 ();
 sg13g2_decap_8 FILLER_59_1029 ();
 sg13g2_decap_8 FILLER_59_1036 ();
 sg13g2_decap_8 FILLER_59_1043 ();
 sg13g2_decap_8 FILLER_59_1050 ();
 sg13g2_decap_8 FILLER_59_1057 ();
 sg13g2_decap_8 FILLER_59_1064 ();
 sg13g2_decap_8 FILLER_59_1071 ();
 sg13g2_decap_8 FILLER_59_1078 ();
 sg13g2_decap_8 FILLER_59_1085 ();
 sg13g2_decap_8 FILLER_59_1092 ();
 sg13g2_decap_8 FILLER_59_1099 ();
 sg13g2_decap_8 FILLER_59_1106 ();
 sg13g2_decap_8 FILLER_59_1113 ();
 sg13g2_decap_8 FILLER_59_1120 ();
 sg13g2_decap_8 FILLER_59_1127 ();
 sg13g2_decap_8 FILLER_59_1134 ();
 sg13g2_decap_8 FILLER_59_1141 ();
 sg13g2_decap_8 FILLER_59_1148 ();
 sg13g2_decap_8 FILLER_59_1155 ();
 sg13g2_decap_8 FILLER_59_1162 ();
 sg13g2_decap_8 FILLER_59_1169 ();
 sg13g2_decap_8 FILLER_59_1176 ();
 sg13g2_decap_8 FILLER_59_1183 ();
 sg13g2_decap_8 FILLER_59_1190 ();
 sg13g2_decap_8 FILLER_59_1197 ();
 sg13g2_decap_8 FILLER_59_1204 ();
 sg13g2_decap_8 FILLER_59_1211 ();
 sg13g2_decap_8 FILLER_59_1218 ();
 sg13g2_decap_8 FILLER_59_1225 ();
 sg13g2_decap_8 FILLER_59_1232 ();
 sg13g2_decap_8 FILLER_59_1239 ();
 sg13g2_decap_8 FILLER_59_1246 ();
 sg13g2_decap_8 FILLER_59_1253 ();
 sg13g2_decap_8 FILLER_59_1260 ();
 sg13g2_decap_8 FILLER_59_1267 ();
 sg13g2_decap_8 FILLER_59_1274 ();
 sg13g2_decap_8 FILLER_59_1281 ();
 sg13g2_decap_8 FILLER_59_1288 ();
 sg13g2_decap_8 FILLER_59_1295 ();
 sg13g2_decap_8 FILLER_59_1302 ();
 sg13g2_decap_8 FILLER_59_1309 ();
 sg13g2_decap_8 FILLER_59_1316 ();
 sg13g2_decap_8 FILLER_59_1323 ();
 sg13g2_decap_8 FILLER_59_1330 ();
 sg13g2_decap_8 FILLER_59_1337 ();
 sg13g2_decap_8 FILLER_59_1344 ();
 sg13g2_decap_8 FILLER_59_1351 ();
 sg13g2_decap_8 FILLER_59_1358 ();
 sg13g2_decap_8 FILLER_59_1365 ();
 sg13g2_decap_8 FILLER_59_1372 ();
 sg13g2_decap_8 FILLER_59_1379 ();
 sg13g2_decap_8 FILLER_59_1386 ();
 sg13g2_decap_8 FILLER_59_1393 ();
 sg13g2_decap_8 FILLER_59_1400 ();
 sg13g2_decap_8 FILLER_59_1407 ();
 sg13g2_decap_8 FILLER_59_1414 ();
 sg13g2_decap_8 FILLER_59_1421 ();
 sg13g2_decap_8 FILLER_59_1428 ();
 sg13g2_decap_8 FILLER_59_1435 ();
 sg13g2_decap_8 FILLER_59_1442 ();
 sg13g2_decap_8 FILLER_59_1449 ();
 sg13g2_decap_8 FILLER_59_1456 ();
 sg13g2_decap_8 FILLER_59_1463 ();
 sg13g2_decap_8 FILLER_59_1470 ();
 sg13g2_decap_8 FILLER_59_1477 ();
 sg13g2_decap_8 FILLER_59_1484 ();
 sg13g2_decap_8 FILLER_59_1491 ();
 sg13g2_decap_8 FILLER_59_1498 ();
 sg13g2_decap_8 FILLER_59_1505 ();
 sg13g2_decap_8 FILLER_59_1512 ();
 sg13g2_decap_8 FILLER_59_1519 ();
 sg13g2_decap_8 FILLER_59_1526 ();
 sg13g2_decap_8 FILLER_59_1533 ();
 sg13g2_decap_8 FILLER_59_1540 ();
 sg13g2_decap_8 FILLER_59_1547 ();
 sg13g2_decap_8 FILLER_59_1554 ();
 sg13g2_decap_8 FILLER_59_1561 ();
 sg13g2_decap_8 FILLER_59_1568 ();
 sg13g2_decap_8 FILLER_59_1575 ();
 sg13g2_decap_8 FILLER_59_1582 ();
 sg13g2_decap_8 FILLER_59_1589 ();
 sg13g2_decap_8 FILLER_59_1596 ();
 sg13g2_decap_8 FILLER_59_1603 ();
 sg13g2_decap_8 FILLER_59_1610 ();
 sg13g2_decap_8 FILLER_59_1617 ();
 sg13g2_decap_8 FILLER_59_1624 ();
 sg13g2_decap_8 FILLER_59_1631 ();
 sg13g2_decap_8 FILLER_59_1638 ();
 sg13g2_decap_8 FILLER_59_1645 ();
 sg13g2_decap_8 FILLER_59_1652 ();
 sg13g2_decap_8 FILLER_59_1659 ();
 sg13g2_decap_8 FILLER_59_1666 ();
 sg13g2_decap_8 FILLER_59_1673 ();
 sg13g2_decap_8 FILLER_59_1680 ();
 sg13g2_decap_8 FILLER_59_1687 ();
 sg13g2_decap_8 FILLER_59_1694 ();
 sg13g2_decap_8 FILLER_59_1701 ();
 sg13g2_decap_8 FILLER_59_1708 ();
 sg13g2_decap_8 FILLER_59_1715 ();
 sg13g2_decap_8 FILLER_59_1722 ();
 sg13g2_decap_8 FILLER_59_1729 ();
 sg13g2_decap_8 FILLER_59_1736 ();
 sg13g2_decap_8 FILLER_59_1743 ();
 sg13g2_decap_8 FILLER_59_1750 ();
 sg13g2_decap_8 FILLER_59_1757 ();
 sg13g2_decap_8 FILLER_59_1764 ();
 sg13g2_decap_8 FILLER_59_1771 ();
 sg13g2_decap_8 FILLER_59_1778 ();
 sg13g2_decap_8 FILLER_59_1785 ();
 sg13g2_decap_8 FILLER_59_1792 ();
 sg13g2_decap_8 FILLER_59_1799 ();
 sg13g2_decap_8 FILLER_59_1806 ();
 sg13g2_decap_8 FILLER_59_1813 ();
 sg13g2_decap_8 FILLER_59_1820 ();
 sg13g2_decap_8 FILLER_59_1827 ();
 sg13g2_decap_8 FILLER_59_1834 ();
 sg13g2_decap_8 FILLER_59_1841 ();
 sg13g2_decap_8 FILLER_59_1848 ();
 sg13g2_decap_8 FILLER_59_1855 ();
 sg13g2_decap_8 FILLER_59_1862 ();
 sg13g2_decap_8 FILLER_59_1869 ();
 sg13g2_decap_8 FILLER_59_1876 ();
 sg13g2_decap_8 FILLER_59_1883 ();
 sg13g2_decap_8 FILLER_59_1890 ();
 sg13g2_decap_8 FILLER_59_1897 ();
 sg13g2_decap_8 FILLER_59_1904 ();
 sg13g2_decap_8 FILLER_59_1911 ();
 sg13g2_decap_8 FILLER_59_1918 ();
 sg13g2_decap_8 FILLER_59_1925 ();
 sg13g2_decap_8 FILLER_59_1932 ();
 sg13g2_decap_8 FILLER_59_1939 ();
 sg13g2_decap_8 FILLER_59_1946 ();
 sg13g2_decap_8 FILLER_59_1953 ();
 sg13g2_decap_8 FILLER_59_1960 ();
 sg13g2_decap_8 FILLER_59_1967 ();
 sg13g2_decap_8 FILLER_59_1974 ();
 sg13g2_decap_8 FILLER_59_1981 ();
 sg13g2_decap_8 FILLER_59_1988 ();
 sg13g2_decap_8 FILLER_59_1995 ();
 sg13g2_decap_8 FILLER_59_2002 ();
 sg13g2_decap_8 FILLER_59_2009 ();
 sg13g2_decap_8 FILLER_59_2016 ();
 sg13g2_decap_8 FILLER_59_2023 ();
 sg13g2_decap_8 FILLER_59_2030 ();
 sg13g2_decap_8 FILLER_59_2037 ();
 sg13g2_decap_8 FILLER_59_2044 ();
 sg13g2_decap_8 FILLER_59_2051 ();
 sg13g2_decap_8 FILLER_59_2058 ();
 sg13g2_decap_8 FILLER_59_2065 ();
 sg13g2_decap_8 FILLER_59_2072 ();
 sg13g2_decap_8 FILLER_59_2079 ();
 sg13g2_decap_8 FILLER_59_2086 ();
 sg13g2_decap_8 FILLER_59_2093 ();
 sg13g2_decap_8 FILLER_59_2100 ();
 sg13g2_decap_8 FILLER_59_2107 ();
 sg13g2_decap_8 FILLER_59_2114 ();
 sg13g2_decap_8 FILLER_59_2121 ();
 sg13g2_decap_8 FILLER_59_2128 ();
 sg13g2_decap_8 FILLER_59_2135 ();
 sg13g2_decap_8 FILLER_59_2142 ();
 sg13g2_decap_8 FILLER_59_2149 ();
 sg13g2_decap_8 FILLER_59_2156 ();
 sg13g2_decap_8 FILLER_59_2163 ();
 sg13g2_decap_8 FILLER_59_2170 ();
 sg13g2_decap_8 FILLER_59_2177 ();
 sg13g2_decap_8 FILLER_59_2184 ();
 sg13g2_decap_8 FILLER_59_2191 ();
 sg13g2_decap_8 FILLER_59_2198 ();
 sg13g2_decap_8 FILLER_59_2205 ();
 sg13g2_decap_8 FILLER_59_2212 ();
 sg13g2_decap_8 FILLER_59_2219 ();
 sg13g2_decap_8 FILLER_59_2226 ();
 sg13g2_decap_8 FILLER_59_2233 ();
 sg13g2_decap_8 FILLER_59_2240 ();
 sg13g2_decap_8 FILLER_59_2247 ();
 sg13g2_decap_8 FILLER_59_2254 ();
 sg13g2_decap_8 FILLER_59_2261 ();
 sg13g2_decap_8 FILLER_59_2268 ();
 sg13g2_decap_8 FILLER_59_2275 ();
 sg13g2_decap_8 FILLER_59_2282 ();
 sg13g2_decap_8 FILLER_59_2289 ();
 sg13g2_decap_8 FILLER_59_2296 ();
 sg13g2_decap_8 FILLER_59_2303 ();
 sg13g2_decap_8 FILLER_59_2310 ();
 sg13g2_decap_8 FILLER_59_2317 ();
 sg13g2_decap_8 FILLER_59_2324 ();
 sg13g2_decap_8 FILLER_59_2331 ();
 sg13g2_decap_8 FILLER_59_2338 ();
 sg13g2_decap_8 FILLER_59_2345 ();
 sg13g2_decap_8 FILLER_59_2352 ();
 sg13g2_decap_8 FILLER_59_2359 ();
 sg13g2_decap_8 FILLER_59_2366 ();
 sg13g2_decap_8 FILLER_59_2373 ();
 sg13g2_decap_8 FILLER_59_2380 ();
 sg13g2_decap_8 FILLER_59_2387 ();
 sg13g2_decap_8 FILLER_59_2394 ();
 sg13g2_decap_8 FILLER_59_2401 ();
 sg13g2_decap_8 FILLER_59_2408 ();
 sg13g2_decap_8 FILLER_59_2415 ();
 sg13g2_decap_8 FILLER_59_2422 ();
 sg13g2_decap_8 FILLER_59_2429 ();
 sg13g2_decap_8 FILLER_59_2436 ();
 sg13g2_decap_8 FILLER_59_2443 ();
 sg13g2_decap_8 FILLER_59_2450 ();
 sg13g2_decap_8 FILLER_59_2457 ();
 sg13g2_decap_8 FILLER_59_2464 ();
 sg13g2_decap_8 FILLER_59_2471 ();
 sg13g2_decap_8 FILLER_59_2478 ();
 sg13g2_decap_8 FILLER_59_2485 ();
 sg13g2_decap_8 FILLER_59_2492 ();
 sg13g2_decap_8 FILLER_59_2499 ();
 sg13g2_decap_8 FILLER_59_2506 ();
 sg13g2_decap_8 FILLER_59_2513 ();
 sg13g2_decap_8 FILLER_59_2520 ();
 sg13g2_decap_8 FILLER_59_2527 ();
 sg13g2_decap_8 FILLER_59_2534 ();
 sg13g2_decap_8 FILLER_59_2541 ();
 sg13g2_decap_8 FILLER_59_2548 ();
 sg13g2_decap_8 FILLER_59_2555 ();
 sg13g2_decap_8 FILLER_59_2562 ();
 sg13g2_decap_8 FILLER_59_2569 ();
 sg13g2_decap_8 FILLER_59_2576 ();
 sg13g2_decap_8 FILLER_59_2583 ();
 sg13g2_decap_8 FILLER_59_2590 ();
 sg13g2_decap_8 FILLER_59_2597 ();
 sg13g2_decap_8 FILLER_59_2604 ();
 sg13g2_decap_8 FILLER_59_2611 ();
 sg13g2_decap_8 FILLER_59_2618 ();
 sg13g2_decap_8 FILLER_59_2625 ();
 sg13g2_decap_8 FILLER_59_2632 ();
 sg13g2_decap_8 FILLER_59_2639 ();
 sg13g2_decap_8 FILLER_59_2646 ();
 sg13g2_decap_8 FILLER_59_2653 ();
 sg13g2_decap_8 FILLER_59_2660 ();
 sg13g2_decap_8 FILLER_59_2667 ();
 sg13g2_decap_8 FILLER_59_2674 ();
 sg13g2_decap_8 FILLER_59_2681 ();
 sg13g2_decap_8 FILLER_59_2688 ();
 sg13g2_decap_8 FILLER_59_2695 ();
 sg13g2_decap_8 FILLER_59_2702 ();
 sg13g2_decap_8 FILLER_59_2709 ();
 sg13g2_decap_8 FILLER_59_2716 ();
 sg13g2_decap_8 FILLER_59_2723 ();
 sg13g2_decap_8 FILLER_59_2730 ();
 sg13g2_decap_8 FILLER_59_2737 ();
 sg13g2_decap_8 FILLER_59_2744 ();
 sg13g2_decap_8 FILLER_59_2751 ();
 sg13g2_decap_8 FILLER_59_2758 ();
 sg13g2_decap_8 FILLER_59_2765 ();
 sg13g2_decap_8 FILLER_59_2772 ();
 sg13g2_decap_8 FILLER_59_2779 ();
 sg13g2_decap_8 FILLER_59_2786 ();
 sg13g2_decap_8 FILLER_59_2793 ();
 sg13g2_decap_8 FILLER_59_2800 ();
 sg13g2_decap_8 FILLER_59_2807 ();
 sg13g2_decap_8 FILLER_59_2814 ();
 sg13g2_decap_8 FILLER_59_2821 ();
 sg13g2_decap_8 FILLER_59_2828 ();
 sg13g2_decap_8 FILLER_59_2835 ();
 sg13g2_decap_8 FILLER_59_2842 ();
 sg13g2_decap_8 FILLER_59_2849 ();
 sg13g2_decap_8 FILLER_59_2856 ();
 sg13g2_decap_8 FILLER_59_2863 ();
 sg13g2_decap_8 FILLER_59_2870 ();
 sg13g2_decap_8 FILLER_59_2877 ();
 sg13g2_decap_8 FILLER_59_2884 ();
 sg13g2_decap_8 FILLER_59_2891 ();
 sg13g2_decap_8 FILLER_59_2898 ();
 sg13g2_decap_8 FILLER_59_2905 ();
 sg13g2_decap_8 FILLER_59_2912 ();
 sg13g2_decap_8 FILLER_59_2919 ();
 sg13g2_decap_8 FILLER_59_2926 ();
 sg13g2_decap_8 FILLER_59_2933 ();
 sg13g2_decap_8 FILLER_59_2940 ();
 sg13g2_decap_8 FILLER_59_2947 ();
 sg13g2_decap_8 FILLER_59_2954 ();
 sg13g2_decap_8 FILLER_59_2961 ();
 sg13g2_decap_8 FILLER_59_2968 ();
 sg13g2_decap_8 FILLER_59_2975 ();
 sg13g2_decap_8 FILLER_59_2982 ();
 sg13g2_decap_8 FILLER_59_2989 ();
 sg13g2_decap_8 FILLER_59_2996 ();
 sg13g2_decap_8 FILLER_59_3003 ();
 sg13g2_decap_8 FILLER_59_3010 ();
 sg13g2_decap_8 FILLER_59_3017 ();
 sg13g2_decap_8 FILLER_59_3024 ();
 sg13g2_decap_8 FILLER_59_3031 ();
 sg13g2_decap_8 FILLER_59_3038 ();
 sg13g2_decap_8 FILLER_59_3045 ();
 sg13g2_decap_8 FILLER_59_3052 ();
 sg13g2_decap_8 FILLER_59_3059 ();
 sg13g2_decap_8 FILLER_59_3066 ();
 sg13g2_decap_8 FILLER_59_3073 ();
 sg13g2_decap_8 FILLER_59_3080 ();
 sg13g2_decap_8 FILLER_59_3087 ();
 sg13g2_decap_8 FILLER_59_3094 ();
 sg13g2_decap_8 FILLER_59_3101 ();
 sg13g2_decap_8 FILLER_59_3108 ();
 sg13g2_decap_8 FILLER_59_3115 ();
 sg13g2_decap_8 FILLER_59_3122 ();
 sg13g2_decap_8 FILLER_59_3129 ();
 sg13g2_decap_8 FILLER_59_3136 ();
 sg13g2_decap_8 FILLER_59_3143 ();
 sg13g2_decap_8 FILLER_59_3150 ();
 sg13g2_decap_8 FILLER_59_3157 ();
 sg13g2_decap_8 FILLER_59_3164 ();
 sg13g2_decap_8 FILLER_59_3171 ();
 sg13g2_decap_8 FILLER_59_3178 ();
 sg13g2_decap_8 FILLER_59_3185 ();
 sg13g2_decap_8 FILLER_59_3192 ();
 sg13g2_decap_8 FILLER_59_3199 ();
 sg13g2_decap_8 FILLER_59_3206 ();
 sg13g2_decap_8 FILLER_59_3213 ();
 sg13g2_decap_8 FILLER_59_3220 ();
 sg13g2_decap_8 FILLER_59_3227 ();
 sg13g2_decap_8 FILLER_59_3234 ();
 sg13g2_decap_8 FILLER_59_3241 ();
 sg13g2_decap_8 FILLER_59_3248 ();
 sg13g2_decap_8 FILLER_59_3255 ();
 sg13g2_decap_8 FILLER_59_3262 ();
 sg13g2_decap_8 FILLER_59_3269 ();
 sg13g2_decap_8 FILLER_59_3276 ();
 sg13g2_decap_8 FILLER_59_3283 ();
 sg13g2_decap_8 FILLER_59_3290 ();
 sg13g2_decap_8 FILLER_59_3297 ();
 sg13g2_decap_8 FILLER_59_3304 ();
 sg13g2_decap_8 FILLER_59_3311 ();
 sg13g2_decap_8 FILLER_59_3318 ();
 sg13g2_decap_8 FILLER_59_3325 ();
 sg13g2_decap_8 FILLER_59_3332 ();
 sg13g2_decap_8 FILLER_59_3339 ();
 sg13g2_decap_8 FILLER_59_3346 ();
 sg13g2_decap_8 FILLER_59_3353 ();
 sg13g2_decap_8 FILLER_59_3360 ();
 sg13g2_decap_8 FILLER_59_3367 ();
 sg13g2_decap_8 FILLER_59_3374 ();
 sg13g2_decap_8 FILLER_59_3381 ();
 sg13g2_decap_8 FILLER_59_3388 ();
 sg13g2_decap_8 FILLER_59_3395 ();
 sg13g2_decap_8 FILLER_59_3402 ();
 sg13g2_decap_8 FILLER_59_3409 ();
 sg13g2_decap_8 FILLER_59_3416 ();
 sg13g2_decap_8 FILLER_59_3423 ();
 sg13g2_decap_8 FILLER_59_3430 ();
 sg13g2_decap_8 FILLER_59_3437 ();
 sg13g2_decap_8 FILLER_59_3444 ();
 sg13g2_decap_8 FILLER_59_3451 ();
 sg13g2_decap_8 FILLER_59_3458 ();
 sg13g2_decap_8 FILLER_59_3465 ();
 sg13g2_decap_8 FILLER_59_3472 ();
 sg13g2_decap_8 FILLER_59_3479 ();
 sg13g2_decap_8 FILLER_59_3486 ();
 sg13g2_decap_8 FILLER_59_3493 ();
 sg13g2_decap_8 FILLER_59_3500 ();
 sg13g2_decap_8 FILLER_59_3507 ();
 sg13g2_decap_8 FILLER_59_3514 ();
 sg13g2_decap_8 FILLER_59_3521 ();
 sg13g2_decap_8 FILLER_59_3528 ();
 sg13g2_decap_8 FILLER_59_3535 ();
 sg13g2_decap_8 FILLER_59_3542 ();
 sg13g2_decap_8 FILLER_59_3549 ();
 sg13g2_decap_8 FILLER_59_3556 ();
 sg13g2_decap_8 FILLER_59_3563 ();
 sg13g2_decap_8 FILLER_59_3570 ();
 sg13g2_fill_2 FILLER_59_3577 ();
 sg13g2_fill_1 FILLER_59_3579 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_98 ();
 sg13g2_decap_8 FILLER_60_105 ();
 sg13g2_decap_8 FILLER_60_112 ();
 sg13g2_decap_8 FILLER_60_119 ();
 sg13g2_decap_8 FILLER_60_126 ();
 sg13g2_decap_8 FILLER_60_133 ();
 sg13g2_decap_8 FILLER_60_140 ();
 sg13g2_decap_8 FILLER_60_147 ();
 sg13g2_decap_8 FILLER_60_154 ();
 sg13g2_decap_8 FILLER_60_161 ();
 sg13g2_decap_8 FILLER_60_168 ();
 sg13g2_decap_8 FILLER_60_175 ();
 sg13g2_decap_8 FILLER_60_182 ();
 sg13g2_decap_8 FILLER_60_189 ();
 sg13g2_decap_8 FILLER_60_196 ();
 sg13g2_decap_8 FILLER_60_203 ();
 sg13g2_decap_8 FILLER_60_210 ();
 sg13g2_decap_8 FILLER_60_217 ();
 sg13g2_decap_8 FILLER_60_224 ();
 sg13g2_decap_8 FILLER_60_231 ();
 sg13g2_decap_8 FILLER_60_238 ();
 sg13g2_decap_8 FILLER_60_245 ();
 sg13g2_decap_8 FILLER_60_252 ();
 sg13g2_decap_8 FILLER_60_259 ();
 sg13g2_decap_8 FILLER_60_266 ();
 sg13g2_decap_8 FILLER_60_273 ();
 sg13g2_decap_8 FILLER_60_280 ();
 sg13g2_decap_8 FILLER_60_287 ();
 sg13g2_decap_8 FILLER_60_294 ();
 sg13g2_decap_8 FILLER_60_301 ();
 sg13g2_decap_8 FILLER_60_308 ();
 sg13g2_decap_8 FILLER_60_315 ();
 sg13g2_decap_8 FILLER_60_322 ();
 sg13g2_decap_8 FILLER_60_329 ();
 sg13g2_decap_8 FILLER_60_336 ();
 sg13g2_decap_8 FILLER_60_343 ();
 sg13g2_decap_8 FILLER_60_350 ();
 sg13g2_decap_8 FILLER_60_357 ();
 sg13g2_decap_8 FILLER_60_364 ();
 sg13g2_decap_8 FILLER_60_371 ();
 sg13g2_decap_8 FILLER_60_378 ();
 sg13g2_decap_8 FILLER_60_385 ();
 sg13g2_decap_8 FILLER_60_392 ();
 sg13g2_decap_8 FILLER_60_399 ();
 sg13g2_decap_8 FILLER_60_406 ();
 sg13g2_decap_8 FILLER_60_413 ();
 sg13g2_decap_8 FILLER_60_420 ();
 sg13g2_decap_8 FILLER_60_427 ();
 sg13g2_decap_8 FILLER_60_434 ();
 sg13g2_decap_8 FILLER_60_441 ();
 sg13g2_decap_8 FILLER_60_448 ();
 sg13g2_decap_8 FILLER_60_455 ();
 sg13g2_decap_8 FILLER_60_462 ();
 sg13g2_decap_8 FILLER_60_469 ();
 sg13g2_decap_8 FILLER_60_476 ();
 sg13g2_decap_8 FILLER_60_483 ();
 sg13g2_decap_8 FILLER_60_490 ();
 sg13g2_decap_8 FILLER_60_497 ();
 sg13g2_decap_8 FILLER_60_504 ();
 sg13g2_decap_8 FILLER_60_511 ();
 sg13g2_decap_8 FILLER_60_518 ();
 sg13g2_decap_8 FILLER_60_525 ();
 sg13g2_decap_8 FILLER_60_532 ();
 sg13g2_decap_8 FILLER_60_539 ();
 sg13g2_decap_8 FILLER_60_546 ();
 sg13g2_decap_8 FILLER_60_553 ();
 sg13g2_decap_8 FILLER_60_560 ();
 sg13g2_decap_8 FILLER_60_567 ();
 sg13g2_decap_8 FILLER_60_574 ();
 sg13g2_decap_8 FILLER_60_581 ();
 sg13g2_decap_8 FILLER_60_588 ();
 sg13g2_decap_8 FILLER_60_595 ();
 sg13g2_decap_8 FILLER_60_602 ();
 sg13g2_decap_8 FILLER_60_609 ();
 sg13g2_decap_8 FILLER_60_616 ();
 sg13g2_decap_8 FILLER_60_623 ();
 sg13g2_decap_8 FILLER_60_630 ();
 sg13g2_decap_8 FILLER_60_637 ();
 sg13g2_decap_8 FILLER_60_644 ();
 sg13g2_decap_8 FILLER_60_651 ();
 sg13g2_decap_8 FILLER_60_658 ();
 sg13g2_decap_8 FILLER_60_665 ();
 sg13g2_decap_8 FILLER_60_672 ();
 sg13g2_decap_8 FILLER_60_679 ();
 sg13g2_decap_8 FILLER_60_686 ();
 sg13g2_decap_8 FILLER_60_693 ();
 sg13g2_decap_8 FILLER_60_700 ();
 sg13g2_decap_8 FILLER_60_707 ();
 sg13g2_decap_8 FILLER_60_714 ();
 sg13g2_decap_8 FILLER_60_721 ();
 sg13g2_decap_8 FILLER_60_728 ();
 sg13g2_decap_8 FILLER_60_735 ();
 sg13g2_decap_8 FILLER_60_742 ();
 sg13g2_decap_8 FILLER_60_749 ();
 sg13g2_decap_8 FILLER_60_756 ();
 sg13g2_decap_8 FILLER_60_763 ();
 sg13g2_decap_8 FILLER_60_770 ();
 sg13g2_decap_8 FILLER_60_777 ();
 sg13g2_decap_8 FILLER_60_784 ();
 sg13g2_decap_8 FILLER_60_791 ();
 sg13g2_decap_8 FILLER_60_798 ();
 sg13g2_decap_8 FILLER_60_805 ();
 sg13g2_decap_8 FILLER_60_812 ();
 sg13g2_decap_8 FILLER_60_819 ();
 sg13g2_decap_8 FILLER_60_826 ();
 sg13g2_decap_8 FILLER_60_833 ();
 sg13g2_decap_8 FILLER_60_840 ();
 sg13g2_decap_8 FILLER_60_847 ();
 sg13g2_decap_8 FILLER_60_854 ();
 sg13g2_decap_8 FILLER_60_861 ();
 sg13g2_decap_8 FILLER_60_868 ();
 sg13g2_decap_8 FILLER_60_875 ();
 sg13g2_decap_8 FILLER_60_882 ();
 sg13g2_decap_8 FILLER_60_889 ();
 sg13g2_decap_8 FILLER_60_896 ();
 sg13g2_decap_8 FILLER_60_903 ();
 sg13g2_decap_8 FILLER_60_910 ();
 sg13g2_decap_8 FILLER_60_917 ();
 sg13g2_decap_8 FILLER_60_924 ();
 sg13g2_decap_8 FILLER_60_931 ();
 sg13g2_decap_8 FILLER_60_938 ();
 sg13g2_decap_8 FILLER_60_945 ();
 sg13g2_decap_8 FILLER_60_952 ();
 sg13g2_decap_8 FILLER_60_959 ();
 sg13g2_decap_8 FILLER_60_966 ();
 sg13g2_decap_8 FILLER_60_973 ();
 sg13g2_decap_8 FILLER_60_980 ();
 sg13g2_decap_8 FILLER_60_987 ();
 sg13g2_decap_8 FILLER_60_994 ();
 sg13g2_decap_8 FILLER_60_1001 ();
 sg13g2_decap_8 FILLER_60_1008 ();
 sg13g2_decap_8 FILLER_60_1015 ();
 sg13g2_decap_8 FILLER_60_1022 ();
 sg13g2_decap_8 FILLER_60_1029 ();
 sg13g2_decap_8 FILLER_60_1036 ();
 sg13g2_decap_8 FILLER_60_1043 ();
 sg13g2_decap_8 FILLER_60_1050 ();
 sg13g2_decap_8 FILLER_60_1057 ();
 sg13g2_decap_8 FILLER_60_1064 ();
 sg13g2_decap_8 FILLER_60_1071 ();
 sg13g2_decap_8 FILLER_60_1078 ();
 sg13g2_decap_8 FILLER_60_1085 ();
 sg13g2_decap_8 FILLER_60_1092 ();
 sg13g2_decap_8 FILLER_60_1099 ();
 sg13g2_decap_8 FILLER_60_1106 ();
 sg13g2_decap_8 FILLER_60_1113 ();
 sg13g2_decap_8 FILLER_60_1120 ();
 sg13g2_decap_8 FILLER_60_1127 ();
 sg13g2_decap_8 FILLER_60_1134 ();
 sg13g2_decap_8 FILLER_60_1141 ();
 sg13g2_decap_8 FILLER_60_1148 ();
 sg13g2_decap_8 FILLER_60_1155 ();
 sg13g2_decap_8 FILLER_60_1162 ();
 sg13g2_decap_8 FILLER_60_1169 ();
 sg13g2_decap_8 FILLER_60_1176 ();
 sg13g2_decap_8 FILLER_60_1183 ();
 sg13g2_decap_8 FILLER_60_1190 ();
 sg13g2_decap_8 FILLER_60_1197 ();
 sg13g2_decap_8 FILLER_60_1204 ();
 sg13g2_decap_8 FILLER_60_1211 ();
 sg13g2_decap_8 FILLER_60_1218 ();
 sg13g2_decap_8 FILLER_60_1225 ();
 sg13g2_decap_8 FILLER_60_1232 ();
 sg13g2_decap_8 FILLER_60_1239 ();
 sg13g2_decap_8 FILLER_60_1246 ();
 sg13g2_decap_8 FILLER_60_1253 ();
 sg13g2_decap_8 FILLER_60_1260 ();
 sg13g2_decap_8 FILLER_60_1267 ();
 sg13g2_decap_8 FILLER_60_1274 ();
 sg13g2_decap_8 FILLER_60_1281 ();
 sg13g2_decap_8 FILLER_60_1288 ();
 sg13g2_decap_8 FILLER_60_1295 ();
 sg13g2_decap_8 FILLER_60_1302 ();
 sg13g2_decap_8 FILLER_60_1309 ();
 sg13g2_decap_8 FILLER_60_1316 ();
 sg13g2_decap_8 FILLER_60_1323 ();
 sg13g2_decap_8 FILLER_60_1330 ();
 sg13g2_decap_8 FILLER_60_1337 ();
 sg13g2_decap_8 FILLER_60_1344 ();
 sg13g2_decap_8 FILLER_60_1351 ();
 sg13g2_decap_8 FILLER_60_1358 ();
 sg13g2_decap_8 FILLER_60_1365 ();
 sg13g2_decap_8 FILLER_60_1372 ();
 sg13g2_decap_8 FILLER_60_1379 ();
 sg13g2_decap_8 FILLER_60_1386 ();
 sg13g2_decap_8 FILLER_60_1393 ();
 sg13g2_decap_8 FILLER_60_1400 ();
 sg13g2_decap_8 FILLER_60_1407 ();
 sg13g2_decap_8 FILLER_60_1414 ();
 sg13g2_decap_8 FILLER_60_1421 ();
 sg13g2_decap_8 FILLER_60_1428 ();
 sg13g2_decap_8 FILLER_60_1435 ();
 sg13g2_decap_8 FILLER_60_1442 ();
 sg13g2_decap_8 FILLER_60_1449 ();
 sg13g2_decap_8 FILLER_60_1456 ();
 sg13g2_decap_8 FILLER_60_1463 ();
 sg13g2_decap_8 FILLER_60_1470 ();
 sg13g2_decap_8 FILLER_60_1477 ();
 sg13g2_decap_8 FILLER_60_1484 ();
 sg13g2_decap_8 FILLER_60_1491 ();
 sg13g2_decap_8 FILLER_60_1498 ();
 sg13g2_decap_8 FILLER_60_1505 ();
 sg13g2_decap_8 FILLER_60_1512 ();
 sg13g2_decap_8 FILLER_60_1519 ();
 sg13g2_decap_8 FILLER_60_1526 ();
 sg13g2_decap_8 FILLER_60_1533 ();
 sg13g2_decap_8 FILLER_60_1540 ();
 sg13g2_decap_8 FILLER_60_1547 ();
 sg13g2_decap_8 FILLER_60_1554 ();
 sg13g2_decap_8 FILLER_60_1561 ();
 sg13g2_decap_8 FILLER_60_1568 ();
 sg13g2_decap_8 FILLER_60_1575 ();
 sg13g2_decap_8 FILLER_60_1582 ();
 sg13g2_decap_8 FILLER_60_1589 ();
 sg13g2_decap_8 FILLER_60_1596 ();
 sg13g2_decap_8 FILLER_60_1603 ();
 sg13g2_decap_8 FILLER_60_1610 ();
 sg13g2_decap_8 FILLER_60_1617 ();
 sg13g2_decap_8 FILLER_60_1624 ();
 sg13g2_decap_8 FILLER_60_1631 ();
 sg13g2_decap_8 FILLER_60_1638 ();
 sg13g2_decap_8 FILLER_60_1645 ();
 sg13g2_decap_8 FILLER_60_1652 ();
 sg13g2_decap_8 FILLER_60_1659 ();
 sg13g2_decap_8 FILLER_60_1666 ();
 sg13g2_decap_8 FILLER_60_1673 ();
 sg13g2_decap_8 FILLER_60_1680 ();
 sg13g2_decap_8 FILLER_60_1687 ();
 sg13g2_decap_8 FILLER_60_1694 ();
 sg13g2_decap_8 FILLER_60_1701 ();
 sg13g2_decap_8 FILLER_60_1708 ();
 sg13g2_decap_8 FILLER_60_1715 ();
 sg13g2_decap_8 FILLER_60_1722 ();
 sg13g2_decap_8 FILLER_60_1729 ();
 sg13g2_decap_8 FILLER_60_1736 ();
 sg13g2_decap_8 FILLER_60_1743 ();
 sg13g2_decap_8 FILLER_60_1750 ();
 sg13g2_decap_8 FILLER_60_1757 ();
 sg13g2_decap_8 FILLER_60_1764 ();
 sg13g2_decap_8 FILLER_60_1771 ();
 sg13g2_decap_8 FILLER_60_1778 ();
 sg13g2_decap_8 FILLER_60_1785 ();
 sg13g2_decap_8 FILLER_60_1792 ();
 sg13g2_decap_8 FILLER_60_1799 ();
 sg13g2_decap_8 FILLER_60_1806 ();
 sg13g2_decap_8 FILLER_60_1813 ();
 sg13g2_decap_8 FILLER_60_1820 ();
 sg13g2_decap_8 FILLER_60_1827 ();
 sg13g2_decap_8 FILLER_60_1834 ();
 sg13g2_decap_8 FILLER_60_1841 ();
 sg13g2_decap_8 FILLER_60_1848 ();
 sg13g2_decap_8 FILLER_60_1855 ();
 sg13g2_decap_8 FILLER_60_1862 ();
 sg13g2_decap_8 FILLER_60_1869 ();
 sg13g2_decap_8 FILLER_60_1876 ();
 sg13g2_decap_8 FILLER_60_1883 ();
 sg13g2_decap_8 FILLER_60_1890 ();
 sg13g2_decap_8 FILLER_60_1897 ();
 sg13g2_decap_8 FILLER_60_1904 ();
 sg13g2_decap_8 FILLER_60_1911 ();
 sg13g2_decap_8 FILLER_60_1918 ();
 sg13g2_decap_8 FILLER_60_1925 ();
 sg13g2_decap_8 FILLER_60_1932 ();
 sg13g2_decap_8 FILLER_60_1939 ();
 sg13g2_decap_8 FILLER_60_1946 ();
 sg13g2_decap_8 FILLER_60_1953 ();
 sg13g2_decap_8 FILLER_60_1960 ();
 sg13g2_decap_8 FILLER_60_1967 ();
 sg13g2_decap_8 FILLER_60_1974 ();
 sg13g2_decap_8 FILLER_60_1981 ();
 sg13g2_decap_8 FILLER_60_1988 ();
 sg13g2_decap_8 FILLER_60_1995 ();
 sg13g2_decap_8 FILLER_60_2002 ();
 sg13g2_decap_8 FILLER_60_2009 ();
 sg13g2_decap_8 FILLER_60_2016 ();
 sg13g2_decap_8 FILLER_60_2023 ();
 sg13g2_decap_8 FILLER_60_2030 ();
 sg13g2_decap_8 FILLER_60_2037 ();
 sg13g2_decap_8 FILLER_60_2044 ();
 sg13g2_decap_8 FILLER_60_2051 ();
 sg13g2_decap_8 FILLER_60_2058 ();
 sg13g2_decap_8 FILLER_60_2065 ();
 sg13g2_decap_8 FILLER_60_2072 ();
 sg13g2_decap_8 FILLER_60_2079 ();
 sg13g2_decap_8 FILLER_60_2086 ();
 sg13g2_decap_8 FILLER_60_2093 ();
 sg13g2_decap_8 FILLER_60_2100 ();
 sg13g2_decap_8 FILLER_60_2107 ();
 sg13g2_decap_8 FILLER_60_2114 ();
 sg13g2_decap_8 FILLER_60_2121 ();
 sg13g2_decap_8 FILLER_60_2128 ();
 sg13g2_decap_8 FILLER_60_2135 ();
 sg13g2_decap_8 FILLER_60_2142 ();
 sg13g2_decap_8 FILLER_60_2149 ();
 sg13g2_decap_8 FILLER_60_2156 ();
 sg13g2_decap_8 FILLER_60_2163 ();
 sg13g2_decap_8 FILLER_60_2170 ();
 sg13g2_decap_8 FILLER_60_2177 ();
 sg13g2_decap_8 FILLER_60_2184 ();
 sg13g2_decap_8 FILLER_60_2191 ();
 sg13g2_decap_8 FILLER_60_2198 ();
 sg13g2_decap_8 FILLER_60_2205 ();
 sg13g2_decap_8 FILLER_60_2212 ();
 sg13g2_decap_8 FILLER_60_2219 ();
 sg13g2_decap_8 FILLER_60_2226 ();
 sg13g2_decap_8 FILLER_60_2233 ();
 sg13g2_decap_8 FILLER_60_2240 ();
 sg13g2_decap_8 FILLER_60_2247 ();
 sg13g2_decap_8 FILLER_60_2254 ();
 sg13g2_decap_8 FILLER_60_2261 ();
 sg13g2_decap_8 FILLER_60_2268 ();
 sg13g2_decap_8 FILLER_60_2275 ();
 sg13g2_decap_8 FILLER_60_2282 ();
 sg13g2_decap_8 FILLER_60_2289 ();
 sg13g2_decap_8 FILLER_60_2296 ();
 sg13g2_decap_8 FILLER_60_2303 ();
 sg13g2_decap_8 FILLER_60_2310 ();
 sg13g2_decap_8 FILLER_60_2317 ();
 sg13g2_decap_8 FILLER_60_2324 ();
 sg13g2_decap_8 FILLER_60_2331 ();
 sg13g2_decap_8 FILLER_60_2338 ();
 sg13g2_decap_8 FILLER_60_2345 ();
 sg13g2_decap_8 FILLER_60_2352 ();
 sg13g2_decap_8 FILLER_60_2359 ();
 sg13g2_decap_8 FILLER_60_2366 ();
 sg13g2_decap_8 FILLER_60_2373 ();
 sg13g2_decap_8 FILLER_60_2380 ();
 sg13g2_decap_8 FILLER_60_2387 ();
 sg13g2_decap_8 FILLER_60_2394 ();
 sg13g2_decap_8 FILLER_60_2401 ();
 sg13g2_decap_8 FILLER_60_2408 ();
 sg13g2_decap_8 FILLER_60_2415 ();
 sg13g2_decap_8 FILLER_60_2422 ();
 sg13g2_decap_8 FILLER_60_2429 ();
 sg13g2_decap_8 FILLER_60_2436 ();
 sg13g2_decap_8 FILLER_60_2443 ();
 sg13g2_decap_8 FILLER_60_2450 ();
 sg13g2_decap_8 FILLER_60_2457 ();
 sg13g2_decap_8 FILLER_60_2464 ();
 sg13g2_decap_8 FILLER_60_2471 ();
 sg13g2_decap_8 FILLER_60_2478 ();
 sg13g2_decap_8 FILLER_60_2485 ();
 sg13g2_decap_8 FILLER_60_2492 ();
 sg13g2_decap_8 FILLER_60_2499 ();
 sg13g2_decap_8 FILLER_60_2506 ();
 sg13g2_decap_8 FILLER_60_2513 ();
 sg13g2_decap_8 FILLER_60_2520 ();
 sg13g2_decap_8 FILLER_60_2527 ();
 sg13g2_decap_8 FILLER_60_2534 ();
 sg13g2_decap_8 FILLER_60_2541 ();
 sg13g2_decap_8 FILLER_60_2548 ();
 sg13g2_decap_8 FILLER_60_2555 ();
 sg13g2_decap_8 FILLER_60_2562 ();
 sg13g2_decap_8 FILLER_60_2569 ();
 sg13g2_decap_8 FILLER_60_2576 ();
 sg13g2_decap_8 FILLER_60_2583 ();
 sg13g2_decap_8 FILLER_60_2590 ();
 sg13g2_decap_8 FILLER_60_2597 ();
 sg13g2_decap_8 FILLER_60_2604 ();
 sg13g2_decap_8 FILLER_60_2611 ();
 sg13g2_decap_8 FILLER_60_2618 ();
 sg13g2_decap_8 FILLER_60_2625 ();
 sg13g2_decap_8 FILLER_60_2632 ();
 sg13g2_decap_8 FILLER_60_2639 ();
 sg13g2_decap_8 FILLER_60_2646 ();
 sg13g2_decap_8 FILLER_60_2653 ();
 sg13g2_decap_8 FILLER_60_2660 ();
 sg13g2_decap_8 FILLER_60_2667 ();
 sg13g2_decap_8 FILLER_60_2674 ();
 sg13g2_decap_8 FILLER_60_2681 ();
 sg13g2_decap_8 FILLER_60_2688 ();
 sg13g2_decap_8 FILLER_60_2695 ();
 sg13g2_decap_8 FILLER_60_2702 ();
 sg13g2_decap_8 FILLER_60_2709 ();
 sg13g2_decap_8 FILLER_60_2716 ();
 sg13g2_decap_8 FILLER_60_2723 ();
 sg13g2_decap_8 FILLER_60_2730 ();
 sg13g2_decap_8 FILLER_60_2737 ();
 sg13g2_decap_8 FILLER_60_2744 ();
 sg13g2_decap_8 FILLER_60_2751 ();
 sg13g2_decap_8 FILLER_60_2758 ();
 sg13g2_decap_8 FILLER_60_2765 ();
 sg13g2_decap_8 FILLER_60_2772 ();
 sg13g2_decap_8 FILLER_60_2779 ();
 sg13g2_decap_8 FILLER_60_2786 ();
 sg13g2_decap_8 FILLER_60_2793 ();
 sg13g2_decap_8 FILLER_60_2800 ();
 sg13g2_decap_8 FILLER_60_2807 ();
 sg13g2_decap_8 FILLER_60_2814 ();
 sg13g2_decap_8 FILLER_60_2821 ();
 sg13g2_decap_8 FILLER_60_2828 ();
 sg13g2_decap_8 FILLER_60_2835 ();
 sg13g2_decap_8 FILLER_60_2842 ();
 sg13g2_decap_8 FILLER_60_2849 ();
 sg13g2_decap_8 FILLER_60_2856 ();
 sg13g2_decap_8 FILLER_60_2863 ();
 sg13g2_decap_8 FILLER_60_2870 ();
 sg13g2_decap_8 FILLER_60_2877 ();
 sg13g2_decap_8 FILLER_60_2884 ();
 sg13g2_decap_8 FILLER_60_2891 ();
 sg13g2_decap_8 FILLER_60_2898 ();
 sg13g2_decap_8 FILLER_60_2905 ();
 sg13g2_decap_8 FILLER_60_2912 ();
 sg13g2_decap_8 FILLER_60_2919 ();
 sg13g2_decap_8 FILLER_60_2926 ();
 sg13g2_decap_8 FILLER_60_2933 ();
 sg13g2_decap_8 FILLER_60_2940 ();
 sg13g2_decap_8 FILLER_60_2947 ();
 sg13g2_decap_8 FILLER_60_2954 ();
 sg13g2_decap_8 FILLER_60_2961 ();
 sg13g2_decap_8 FILLER_60_2968 ();
 sg13g2_decap_8 FILLER_60_2975 ();
 sg13g2_decap_8 FILLER_60_2982 ();
 sg13g2_decap_8 FILLER_60_2989 ();
 sg13g2_decap_8 FILLER_60_2996 ();
 sg13g2_decap_8 FILLER_60_3003 ();
 sg13g2_decap_8 FILLER_60_3010 ();
 sg13g2_decap_8 FILLER_60_3017 ();
 sg13g2_decap_8 FILLER_60_3024 ();
 sg13g2_decap_8 FILLER_60_3031 ();
 sg13g2_decap_8 FILLER_60_3038 ();
 sg13g2_decap_8 FILLER_60_3045 ();
 sg13g2_decap_8 FILLER_60_3052 ();
 sg13g2_decap_8 FILLER_60_3059 ();
 sg13g2_decap_8 FILLER_60_3066 ();
 sg13g2_decap_8 FILLER_60_3073 ();
 sg13g2_decap_8 FILLER_60_3080 ();
 sg13g2_decap_8 FILLER_60_3087 ();
 sg13g2_decap_8 FILLER_60_3094 ();
 sg13g2_decap_8 FILLER_60_3101 ();
 sg13g2_decap_8 FILLER_60_3108 ();
 sg13g2_decap_8 FILLER_60_3115 ();
 sg13g2_decap_8 FILLER_60_3122 ();
 sg13g2_decap_8 FILLER_60_3129 ();
 sg13g2_decap_8 FILLER_60_3136 ();
 sg13g2_decap_8 FILLER_60_3143 ();
 sg13g2_decap_8 FILLER_60_3150 ();
 sg13g2_decap_8 FILLER_60_3157 ();
 sg13g2_decap_8 FILLER_60_3164 ();
 sg13g2_decap_8 FILLER_60_3171 ();
 sg13g2_decap_8 FILLER_60_3178 ();
 sg13g2_decap_8 FILLER_60_3185 ();
 sg13g2_decap_8 FILLER_60_3192 ();
 sg13g2_decap_8 FILLER_60_3199 ();
 sg13g2_decap_8 FILLER_60_3206 ();
 sg13g2_decap_8 FILLER_60_3213 ();
 sg13g2_decap_8 FILLER_60_3220 ();
 sg13g2_decap_8 FILLER_60_3227 ();
 sg13g2_decap_8 FILLER_60_3234 ();
 sg13g2_decap_8 FILLER_60_3241 ();
 sg13g2_decap_8 FILLER_60_3248 ();
 sg13g2_decap_8 FILLER_60_3255 ();
 sg13g2_decap_8 FILLER_60_3262 ();
 sg13g2_decap_8 FILLER_60_3269 ();
 sg13g2_decap_8 FILLER_60_3276 ();
 sg13g2_decap_8 FILLER_60_3283 ();
 sg13g2_decap_8 FILLER_60_3290 ();
 sg13g2_decap_8 FILLER_60_3297 ();
 sg13g2_decap_8 FILLER_60_3304 ();
 sg13g2_decap_8 FILLER_60_3311 ();
 sg13g2_decap_8 FILLER_60_3318 ();
 sg13g2_decap_8 FILLER_60_3325 ();
 sg13g2_decap_8 FILLER_60_3332 ();
 sg13g2_decap_8 FILLER_60_3339 ();
 sg13g2_decap_8 FILLER_60_3346 ();
 sg13g2_decap_8 FILLER_60_3353 ();
 sg13g2_decap_8 FILLER_60_3360 ();
 sg13g2_decap_8 FILLER_60_3367 ();
 sg13g2_decap_8 FILLER_60_3374 ();
 sg13g2_decap_8 FILLER_60_3381 ();
 sg13g2_decap_8 FILLER_60_3388 ();
 sg13g2_decap_8 FILLER_60_3395 ();
 sg13g2_decap_8 FILLER_60_3402 ();
 sg13g2_decap_8 FILLER_60_3409 ();
 sg13g2_decap_8 FILLER_60_3416 ();
 sg13g2_decap_8 FILLER_60_3423 ();
 sg13g2_decap_8 FILLER_60_3430 ();
 sg13g2_decap_8 FILLER_60_3437 ();
 sg13g2_decap_8 FILLER_60_3444 ();
 sg13g2_decap_8 FILLER_60_3451 ();
 sg13g2_decap_8 FILLER_60_3458 ();
 sg13g2_decap_8 FILLER_60_3465 ();
 sg13g2_decap_8 FILLER_60_3472 ();
 sg13g2_decap_8 FILLER_60_3479 ();
 sg13g2_decap_8 FILLER_60_3486 ();
 sg13g2_decap_8 FILLER_60_3493 ();
 sg13g2_decap_8 FILLER_60_3500 ();
 sg13g2_decap_8 FILLER_60_3507 ();
 sg13g2_decap_8 FILLER_60_3514 ();
 sg13g2_decap_8 FILLER_60_3521 ();
 sg13g2_decap_8 FILLER_60_3528 ();
 sg13g2_decap_8 FILLER_60_3535 ();
 sg13g2_decap_8 FILLER_60_3542 ();
 sg13g2_decap_8 FILLER_60_3549 ();
 sg13g2_decap_8 FILLER_60_3556 ();
 sg13g2_decap_8 FILLER_60_3563 ();
 sg13g2_decap_8 FILLER_60_3570 ();
 sg13g2_fill_2 FILLER_60_3577 ();
 sg13g2_fill_1 FILLER_60_3579 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_8 FILLER_61_91 ();
 sg13g2_decap_8 FILLER_61_98 ();
 sg13g2_decap_8 FILLER_61_105 ();
 sg13g2_decap_8 FILLER_61_112 ();
 sg13g2_decap_8 FILLER_61_119 ();
 sg13g2_decap_8 FILLER_61_126 ();
 sg13g2_decap_8 FILLER_61_133 ();
 sg13g2_decap_8 FILLER_61_140 ();
 sg13g2_decap_8 FILLER_61_147 ();
 sg13g2_decap_8 FILLER_61_154 ();
 sg13g2_decap_8 FILLER_61_161 ();
 sg13g2_decap_8 FILLER_61_168 ();
 sg13g2_decap_8 FILLER_61_175 ();
 sg13g2_decap_8 FILLER_61_182 ();
 sg13g2_decap_8 FILLER_61_189 ();
 sg13g2_decap_8 FILLER_61_196 ();
 sg13g2_decap_8 FILLER_61_203 ();
 sg13g2_decap_8 FILLER_61_210 ();
 sg13g2_decap_8 FILLER_61_217 ();
 sg13g2_decap_8 FILLER_61_224 ();
 sg13g2_decap_8 FILLER_61_231 ();
 sg13g2_decap_8 FILLER_61_238 ();
 sg13g2_decap_8 FILLER_61_245 ();
 sg13g2_decap_8 FILLER_61_252 ();
 sg13g2_decap_8 FILLER_61_259 ();
 sg13g2_decap_8 FILLER_61_266 ();
 sg13g2_decap_8 FILLER_61_273 ();
 sg13g2_decap_8 FILLER_61_280 ();
 sg13g2_decap_8 FILLER_61_287 ();
 sg13g2_decap_8 FILLER_61_294 ();
 sg13g2_decap_8 FILLER_61_301 ();
 sg13g2_decap_8 FILLER_61_308 ();
 sg13g2_decap_8 FILLER_61_315 ();
 sg13g2_decap_8 FILLER_61_322 ();
 sg13g2_decap_8 FILLER_61_329 ();
 sg13g2_decap_8 FILLER_61_336 ();
 sg13g2_decap_8 FILLER_61_343 ();
 sg13g2_decap_8 FILLER_61_350 ();
 sg13g2_decap_8 FILLER_61_357 ();
 sg13g2_decap_8 FILLER_61_364 ();
 sg13g2_decap_8 FILLER_61_371 ();
 sg13g2_decap_8 FILLER_61_378 ();
 sg13g2_decap_8 FILLER_61_385 ();
 sg13g2_decap_8 FILLER_61_392 ();
 sg13g2_decap_8 FILLER_61_399 ();
 sg13g2_decap_8 FILLER_61_406 ();
 sg13g2_decap_8 FILLER_61_413 ();
 sg13g2_decap_8 FILLER_61_420 ();
 sg13g2_decap_8 FILLER_61_427 ();
 sg13g2_decap_8 FILLER_61_434 ();
 sg13g2_decap_8 FILLER_61_441 ();
 sg13g2_decap_8 FILLER_61_448 ();
 sg13g2_decap_8 FILLER_61_455 ();
 sg13g2_decap_8 FILLER_61_462 ();
 sg13g2_decap_8 FILLER_61_469 ();
 sg13g2_decap_8 FILLER_61_476 ();
 sg13g2_decap_8 FILLER_61_483 ();
 sg13g2_decap_8 FILLER_61_490 ();
 sg13g2_decap_8 FILLER_61_497 ();
 sg13g2_decap_8 FILLER_61_504 ();
 sg13g2_decap_8 FILLER_61_511 ();
 sg13g2_decap_8 FILLER_61_518 ();
 sg13g2_decap_8 FILLER_61_525 ();
 sg13g2_decap_8 FILLER_61_532 ();
 sg13g2_decap_8 FILLER_61_539 ();
 sg13g2_decap_8 FILLER_61_546 ();
 sg13g2_decap_8 FILLER_61_553 ();
 sg13g2_decap_8 FILLER_61_560 ();
 sg13g2_decap_8 FILLER_61_567 ();
 sg13g2_decap_8 FILLER_61_574 ();
 sg13g2_decap_8 FILLER_61_581 ();
 sg13g2_decap_8 FILLER_61_588 ();
 sg13g2_decap_8 FILLER_61_595 ();
 sg13g2_decap_8 FILLER_61_602 ();
 sg13g2_decap_8 FILLER_61_609 ();
 sg13g2_decap_8 FILLER_61_616 ();
 sg13g2_decap_8 FILLER_61_623 ();
 sg13g2_decap_8 FILLER_61_630 ();
 sg13g2_decap_8 FILLER_61_637 ();
 sg13g2_decap_8 FILLER_61_644 ();
 sg13g2_decap_8 FILLER_61_651 ();
 sg13g2_decap_8 FILLER_61_658 ();
 sg13g2_decap_8 FILLER_61_665 ();
 sg13g2_decap_8 FILLER_61_672 ();
 sg13g2_decap_8 FILLER_61_679 ();
 sg13g2_decap_8 FILLER_61_686 ();
 sg13g2_decap_8 FILLER_61_693 ();
 sg13g2_decap_8 FILLER_61_700 ();
 sg13g2_decap_8 FILLER_61_707 ();
 sg13g2_decap_8 FILLER_61_714 ();
 sg13g2_decap_8 FILLER_61_721 ();
 sg13g2_decap_8 FILLER_61_728 ();
 sg13g2_decap_8 FILLER_61_735 ();
 sg13g2_decap_8 FILLER_61_742 ();
 sg13g2_decap_8 FILLER_61_749 ();
 sg13g2_decap_8 FILLER_61_756 ();
 sg13g2_decap_8 FILLER_61_763 ();
 sg13g2_decap_8 FILLER_61_770 ();
 sg13g2_decap_8 FILLER_61_777 ();
 sg13g2_decap_8 FILLER_61_784 ();
 sg13g2_decap_8 FILLER_61_791 ();
 sg13g2_decap_8 FILLER_61_798 ();
 sg13g2_decap_8 FILLER_61_805 ();
 sg13g2_decap_8 FILLER_61_812 ();
 sg13g2_decap_8 FILLER_61_819 ();
 sg13g2_decap_8 FILLER_61_826 ();
 sg13g2_decap_8 FILLER_61_833 ();
 sg13g2_decap_8 FILLER_61_840 ();
 sg13g2_decap_8 FILLER_61_847 ();
 sg13g2_decap_8 FILLER_61_854 ();
 sg13g2_decap_8 FILLER_61_861 ();
 sg13g2_decap_8 FILLER_61_868 ();
 sg13g2_decap_8 FILLER_61_875 ();
 sg13g2_decap_8 FILLER_61_882 ();
 sg13g2_decap_8 FILLER_61_889 ();
 sg13g2_decap_8 FILLER_61_896 ();
 sg13g2_decap_8 FILLER_61_903 ();
 sg13g2_decap_8 FILLER_61_910 ();
 sg13g2_decap_8 FILLER_61_917 ();
 sg13g2_decap_8 FILLER_61_924 ();
 sg13g2_decap_8 FILLER_61_931 ();
 sg13g2_decap_8 FILLER_61_938 ();
 sg13g2_decap_8 FILLER_61_945 ();
 sg13g2_decap_8 FILLER_61_952 ();
 sg13g2_decap_8 FILLER_61_959 ();
 sg13g2_decap_8 FILLER_61_966 ();
 sg13g2_decap_8 FILLER_61_973 ();
 sg13g2_decap_8 FILLER_61_980 ();
 sg13g2_decap_8 FILLER_61_987 ();
 sg13g2_decap_8 FILLER_61_994 ();
 sg13g2_decap_8 FILLER_61_1001 ();
 sg13g2_decap_8 FILLER_61_1008 ();
 sg13g2_decap_8 FILLER_61_1015 ();
 sg13g2_decap_8 FILLER_61_1022 ();
 sg13g2_decap_8 FILLER_61_1029 ();
 sg13g2_decap_8 FILLER_61_1036 ();
 sg13g2_decap_8 FILLER_61_1043 ();
 sg13g2_decap_8 FILLER_61_1050 ();
 sg13g2_decap_8 FILLER_61_1057 ();
 sg13g2_decap_8 FILLER_61_1064 ();
 sg13g2_decap_8 FILLER_61_1071 ();
 sg13g2_decap_8 FILLER_61_1078 ();
 sg13g2_decap_8 FILLER_61_1085 ();
 sg13g2_decap_8 FILLER_61_1092 ();
 sg13g2_decap_8 FILLER_61_1099 ();
 sg13g2_decap_8 FILLER_61_1106 ();
 sg13g2_decap_8 FILLER_61_1113 ();
 sg13g2_decap_8 FILLER_61_1120 ();
 sg13g2_decap_8 FILLER_61_1127 ();
 sg13g2_decap_8 FILLER_61_1134 ();
 sg13g2_decap_8 FILLER_61_1141 ();
 sg13g2_decap_8 FILLER_61_1148 ();
 sg13g2_decap_8 FILLER_61_1155 ();
 sg13g2_decap_8 FILLER_61_1162 ();
 sg13g2_decap_8 FILLER_61_1169 ();
 sg13g2_decap_8 FILLER_61_1176 ();
 sg13g2_decap_8 FILLER_61_1183 ();
 sg13g2_decap_8 FILLER_61_1190 ();
 sg13g2_decap_8 FILLER_61_1197 ();
 sg13g2_decap_8 FILLER_61_1204 ();
 sg13g2_decap_8 FILLER_61_1211 ();
 sg13g2_decap_8 FILLER_61_1218 ();
 sg13g2_decap_8 FILLER_61_1225 ();
 sg13g2_decap_8 FILLER_61_1232 ();
 sg13g2_decap_8 FILLER_61_1239 ();
 sg13g2_decap_8 FILLER_61_1246 ();
 sg13g2_decap_8 FILLER_61_1253 ();
 sg13g2_decap_8 FILLER_61_1260 ();
 sg13g2_decap_8 FILLER_61_1267 ();
 sg13g2_decap_8 FILLER_61_1274 ();
 sg13g2_decap_8 FILLER_61_1281 ();
 sg13g2_decap_8 FILLER_61_1288 ();
 sg13g2_decap_8 FILLER_61_1295 ();
 sg13g2_decap_8 FILLER_61_1302 ();
 sg13g2_decap_8 FILLER_61_1309 ();
 sg13g2_decap_8 FILLER_61_1316 ();
 sg13g2_decap_8 FILLER_61_1323 ();
 sg13g2_decap_8 FILLER_61_1330 ();
 sg13g2_decap_8 FILLER_61_1337 ();
 sg13g2_decap_8 FILLER_61_1344 ();
 sg13g2_decap_8 FILLER_61_1351 ();
 sg13g2_decap_8 FILLER_61_1358 ();
 sg13g2_decap_8 FILLER_61_1365 ();
 sg13g2_decap_8 FILLER_61_1372 ();
 sg13g2_decap_8 FILLER_61_1379 ();
 sg13g2_decap_8 FILLER_61_1386 ();
 sg13g2_decap_8 FILLER_61_1393 ();
 sg13g2_decap_8 FILLER_61_1400 ();
 sg13g2_decap_8 FILLER_61_1407 ();
 sg13g2_decap_8 FILLER_61_1414 ();
 sg13g2_decap_8 FILLER_61_1421 ();
 sg13g2_decap_8 FILLER_61_1428 ();
 sg13g2_decap_8 FILLER_61_1435 ();
 sg13g2_decap_8 FILLER_61_1442 ();
 sg13g2_decap_8 FILLER_61_1449 ();
 sg13g2_decap_8 FILLER_61_1456 ();
 sg13g2_decap_8 FILLER_61_1463 ();
 sg13g2_decap_8 FILLER_61_1470 ();
 sg13g2_decap_8 FILLER_61_1477 ();
 sg13g2_decap_8 FILLER_61_1484 ();
 sg13g2_decap_8 FILLER_61_1491 ();
 sg13g2_decap_8 FILLER_61_1498 ();
 sg13g2_decap_8 FILLER_61_1505 ();
 sg13g2_decap_8 FILLER_61_1512 ();
 sg13g2_decap_8 FILLER_61_1519 ();
 sg13g2_decap_8 FILLER_61_1526 ();
 sg13g2_decap_8 FILLER_61_1533 ();
 sg13g2_decap_8 FILLER_61_1540 ();
 sg13g2_decap_8 FILLER_61_1547 ();
 sg13g2_decap_8 FILLER_61_1554 ();
 sg13g2_decap_8 FILLER_61_1561 ();
 sg13g2_decap_8 FILLER_61_1568 ();
 sg13g2_decap_8 FILLER_61_1575 ();
 sg13g2_decap_8 FILLER_61_1582 ();
 sg13g2_decap_8 FILLER_61_1589 ();
 sg13g2_decap_8 FILLER_61_1596 ();
 sg13g2_decap_8 FILLER_61_1603 ();
 sg13g2_decap_8 FILLER_61_1610 ();
 sg13g2_decap_8 FILLER_61_1617 ();
 sg13g2_decap_8 FILLER_61_1624 ();
 sg13g2_decap_8 FILLER_61_1631 ();
 sg13g2_decap_8 FILLER_61_1638 ();
 sg13g2_decap_8 FILLER_61_1645 ();
 sg13g2_decap_8 FILLER_61_1652 ();
 sg13g2_decap_8 FILLER_61_1659 ();
 sg13g2_decap_8 FILLER_61_1666 ();
 sg13g2_decap_8 FILLER_61_1673 ();
 sg13g2_decap_8 FILLER_61_1680 ();
 sg13g2_decap_8 FILLER_61_1687 ();
 sg13g2_decap_8 FILLER_61_1694 ();
 sg13g2_decap_8 FILLER_61_1701 ();
 sg13g2_decap_8 FILLER_61_1708 ();
 sg13g2_decap_8 FILLER_61_1715 ();
 sg13g2_decap_8 FILLER_61_1722 ();
 sg13g2_decap_8 FILLER_61_1729 ();
 sg13g2_decap_8 FILLER_61_1736 ();
 sg13g2_decap_8 FILLER_61_1743 ();
 sg13g2_decap_8 FILLER_61_1750 ();
 sg13g2_decap_8 FILLER_61_1757 ();
 sg13g2_decap_8 FILLER_61_1764 ();
 sg13g2_decap_8 FILLER_61_1771 ();
 sg13g2_decap_8 FILLER_61_1778 ();
 sg13g2_decap_8 FILLER_61_1785 ();
 sg13g2_decap_8 FILLER_61_1792 ();
 sg13g2_decap_8 FILLER_61_1799 ();
 sg13g2_decap_8 FILLER_61_1806 ();
 sg13g2_decap_8 FILLER_61_1813 ();
 sg13g2_decap_8 FILLER_61_1820 ();
 sg13g2_decap_8 FILLER_61_1827 ();
 sg13g2_decap_8 FILLER_61_1834 ();
 sg13g2_decap_8 FILLER_61_1841 ();
 sg13g2_decap_8 FILLER_61_1848 ();
 sg13g2_decap_8 FILLER_61_1855 ();
 sg13g2_decap_8 FILLER_61_1862 ();
 sg13g2_decap_8 FILLER_61_1869 ();
 sg13g2_decap_8 FILLER_61_1876 ();
 sg13g2_decap_8 FILLER_61_1883 ();
 sg13g2_decap_8 FILLER_61_1890 ();
 sg13g2_decap_8 FILLER_61_1897 ();
 sg13g2_decap_8 FILLER_61_1904 ();
 sg13g2_decap_8 FILLER_61_1911 ();
 sg13g2_decap_8 FILLER_61_1918 ();
 sg13g2_decap_8 FILLER_61_1925 ();
 sg13g2_decap_8 FILLER_61_1932 ();
 sg13g2_decap_8 FILLER_61_1939 ();
 sg13g2_decap_8 FILLER_61_1946 ();
 sg13g2_decap_8 FILLER_61_1953 ();
 sg13g2_decap_8 FILLER_61_1960 ();
 sg13g2_decap_8 FILLER_61_1967 ();
 sg13g2_decap_8 FILLER_61_1974 ();
 sg13g2_decap_8 FILLER_61_1981 ();
 sg13g2_decap_8 FILLER_61_1988 ();
 sg13g2_decap_8 FILLER_61_1995 ();
 sg13g2_decap_8 FILLER_61_2002 ();
 sg13g2_decap_8 FILLER_61_2009 ();
 sg13g2_decap_8 FILLER_61_2016 ();
 sg13g2_decap_8 FILLER_61_2023 ();
 sg13g2_decap_8 FILLER_61_2030 ();
 sg13g2_decap_8 FILLER_61_2037 ();
 sg13g2_decap_8 FILLER_61_2044 ();
 sg13g2_decap_8 FILLER_61_2051 ();
 sg13g2_decap_8 FILLER_61_2058 ();
 sg13g2_decap_8 FILLER_61_2065 ();
 sg13g2_decap_8 FILLER_61_2072 ();
 sg13g2_decap_8 FILLER_61_2079 ();
 sg13g2_decap_8 FILLER_61_2086 ();
 sg13g2_decap_8 FILLER_61_2093 ();
 sg13g2_decap_8 FILLER_61_2100 ();
 sg13g2_decap_8 FILLER_61_2107 ();
 sg13g2_decap_8 FILLER_61_2114 ();
 sg13g2_decap_8 FILLER_61_2121 ();
 sg13g2_decap_8 FILLER_61_2128 ();
 sg13g2_decap_8 FILLER_61_2135 ();
 sg13g2_decap_8 FILLER_61_2142 ();
 sg13g2_decap_8 FILLER_61_2149 ();
 sg13g2_decap_8 FILLER_61_2156 ();
 sg13g2_decap_8 FILLER_61_2163 ();
 sg13g2_decap_8 FILLER_61_2170 ();
 sg13g2_decap_8 FILLER_61_2177 ();
 sg13g2_decap_8 FILLER_61_2184 ();
 sg13g2_decap_8 FILLER_61_2191 ();
 sg13g2_decap_8 FILLER_61_2198 ();
 sg13g2_decap_8 FILLER_61_2205 ();
 sg13g2_decap_8 FILLER_61_2212 ();
 sg13g2_decap_8 FILLER_61_2219 ();
 sg13g2_decap_8 FILLER_61_2226 ();
 sg13g2_decap_8 FILLER_61_2233 ();
 sg13g2_decap_8 FILLER_61_2240 ();
 sg13g2_decap_8 FILLER_61_2247 ();
 sg13g2_decap_8 FILLER_61_2254 ();
 sg13g2_decap_8 FILLER_61_2261 ();
 sg13g2_decap_8 FILLER_61_2268 ();
 sg13g2_decap_8 FILLER_61_2275 ();
 sg13g2_decap_8 FILLER_61_2282 ();
 sg13g2_decap_8 FILLER_61_2289 ();
 sg13g2_decap_8 FILLER_61_2296 ();
 sg13g2_decap_8 FILLER_61_2303 ();
 sg13g2_decap_8 FILLER_61_2310 ();
 sg13g2_decap_8 FILLER_61_2317 ();
 sg13g2_decap_8 FILLER_61_2324 ();
 sg13g2_decap_8 FILLER_61_2331 ();
 sg13g2_decap_8 FILLER_61_2338 ();
 sg13g2_decap_8 FILLER_61_2345 ();
 sg13g2_decap_8 FILLER_61_2352 ();
 sg13g2_decap_8 FILLER_61_2359 ();
 sg13g2_decap_8 FILLER_61_2366 ();
 sg13g2_decap_8 FILLER_61_2373 ();
 sg13g2_decap_8 FILLER_61_2380 ();
 sg13g2_decap_8 FILLER_61_2387 ();
 sg13g2_decap_8 FILLER_61_2394 ();
 sg13g2_decap_8 FILLER_61_2401 ();
 sg13g2_decap_8 FILLER_61_2408 ();
 sg13g2_decap_8 FILLER_61_2415 ();
 sg13g2_decap_8 FILLER_61_2422 ();
 sg13g2_decap_8 FILLER_61_2429 ();
 sg13g2_decap_8 FILLER_61_2436 ();
 sg13g2_decap_8 FILLER_61_2443 ();
 sg13g2_decap_8 FILLER_61_2450 ();
 sg13g2_decap_8 FILLER_61_2457 ();
 sg13g2_decap_8 FILLER_61_2464 ();
 sg13g2_decap_8 FILLER_61_2471 ();
 sg13g2_decap_8 FILLER_61_2478 ();
 sg13g2_decap_8 FILLER_61_2485 ();
 sg13g2_decap_8 FILLER_61_2492 ();
 sg13g2_decap_8 FILLER_61_2499 ();
 sg13g2_decap_8 FILLER_61_2506 ();
 sg13g2_decap_8 FILLER_61_2513 ();
 sg13g2_decap_8 FILLER_61_2520 ();
 sg13g2_decap_8 FILLER_61_2527 ();
 sg13g2_decap_8 FILLER_61_2534 ();
 sg13g2_decap_8 FILLER_61_2541 ();
 sg13g2_decap_8 FILLER_61_2548 ();
 sg13g2_decap_8 FILLER_61_2555 ();
 sg13g2_decap_8 FILLER_61_2562 ();
 sg13g2_decap_8 FILLER_61_2569 ();
 sg13g2_decap_8 FILLER_61_2576 ();
 sg13g2_decap_8 FILLER_61_2583 ();
 sg13g2_decap_8 FILLER_61_2590 ();
 sg13g2_decap_8 FILLER_61_2597 ();
 sg13g2_decap_8 FILLER_61_2604 ();
 sg13g2_decap_8 FILLER_61_2611 ();
 sg13g2_decap_8 FILLER_61_2618 ();
 sg13g2_decap_8 FILLER_61_2625 ();
 sg13g2_decap_8 FILLER_61_2632 ();
 sg13g2_decap_8 FILLER_61_2639 ();
 sg13g2_decap_8 FILLER_61_2646 ();
 sg13g2_decap_8 FILLER_61_2653 ();
 sg13g2_decap_8 FILLER_61_2660 ();
 sg13g2_decap_8 FILLER_61_2667 ();
 sg13g2_decap_8 FILLER_61_2674 ();
 sg13g2_decap_8 FILLER_61_2681 ();
 sg13g2_decap_8 FILLER_61_2688 ();
 sg13g2_decap_8 FILLER_61_2695 ();
 sg13g2_decap_8 FILLER_61_2702 ();
 sg13g2_decap_8 FILLER_61_2709 ();
 sg13g2_decap_8 FILLER_61_2716 ();
 sg13g2_decap_8 FILLER_61_2723 ();
 sg13g2_decap_8 FILLER_61_2730 ();
 sg13g2_decap_8 FILLER_61_2737 ();
 sg13g2_decap_8 FILLER_61_2744 ();
 sg13g2_decap_8 FILLER_61_2751 ();
 sg13g2_decap_8 FILLER_61_2758 ();
 sg13g2_decap_8 FILLER_61_2765 ();
 sg13g2_decap_8 FILLER_61_2772 ();
 sg13g2_decap_8 FILLER_61_2779 ();
 sg13g2_decap_8 FILLER_61_2786 ();
 sg13g2_decap_8 FILLER_61_2793 ();
 sg13g2_decap_8 FILLER_61_2800 ();
 sg13g2_decap_8 FILLER_61_2807 ();
 sg13g2_decap_8 FILLER_61_2814 ();
 sg13g2_decap_8 FILLER_61_2821 ();
 sg13g2_decap_8 FILLER_61_2828 ();
 sg13g2_decap_8 FILLER_61_2835 ();
 sg13g2_decap_8 FILLER_61_2842 ();
 sg13g2_decap_8 FILLER_61_2849 ();
 sg13g2_decap_8 FILLER_61_2856 ();
 sg13g2_decap_8 FILLER_61_2863 ();
 sg13g2_decap_8 FILLER_61_2870 ();
 sg13g2_decap_8 FILLER_61_2877 ();
 sg13g2_decap_8 FILLER_61_2884 ();
 sg13g2_decap_8 FILLER_61_2891 ();
 sg13g2_decap_8 FILLER_61_2898 ();
 sg13g2_decap_8 FILLER_61_2905 ();
 sg13g2_decap_8 FILLER_61_2912 ();
 sg13g2_decap_8 FILLER_61_2919 ();
 sg13g2_decap_8 FILLER_61_2926 ();
 sg13g2_decap_8 FILLER_61_2933 ();
 sg13g2_decap_8 FILLER_61_2940 ();
 sg13g2_decap_8 FILLER_61_2947 ();
 sg13g2_decap_8 FILLER_61_2954 ();
 sg13g2_decap_8 FILLER_61_2961 ();
 sg13g2_decap_8 FILLER_61_2968 ();
 sg13g2_decap_8 FILLER_61_2975 ();
 sg13g2_decap_8 FILLER_61_2982 ();
 sg13g2_decap_8 FILLER_61_2989 ();
 sg13g2_decap_8 FILLER_61_2996 ();
 sg13g2_decap_8 FILLER_61_3003 ();
 sg13g2_decap_8 FILLER_61_3010 ();
 sg13g2_decap_8 FILLER_61_3017 ();
 sg13g2_decap_8 FILLER_61_3024 ();
 sg13g2_decap_8 FILLER_61_3031 ();
 sg13g2_decap_8 FILLER_61_3038 ();
 sg13g2_decap_8 FILLER_61_3045 ();
 sg13g2_decap_8 FILLER_61_3052 ();
 sg13g2_decap_8 FILLER_61_3059 ();
 sg13g2_decap_8 FILLER_61_3066 ();
 sg13g2_decap_8 FILLER_61_3073 ();
 sg13g2_decap_8 FILLER_61_3080 ();
 sg13g2_decap_8 FILLER_61_3087 ();
 sg13g2_decap_8 FILLER_61_3094 ();
 sg13g2_decap_8 FILLER_61_3101 ();
 sg13g2_decap_8 FILLER_61_3108 ();
 sg13g2_decap_8 FILLER_61_3115 ();
 sg13g2_decap_8 FILLER_61_3122 ();
 sg13g2_decap_8 FILLER_61_3129 ();
 sg13g2_decap_8 FILLER_61_3136 ();
 sg13g2_decap_8 FILLER_61_3143 ();
 sg13g2_decap_8 FILLER_61_3150 ();
 sg13g2_decap_8 FILLER_61_3157 ();
 sg13g2_decap_8 FILLER_61_3164 ();
 sg13g2_decap_8 FILLER_61_3171 ();
 sg13g2_decap_8 FILLER_61_3178 ();
 sg13g2_decap_8 FILLER_61_3185 ();
 sg13g2_decap_8 FILLER_61_3192 ();
 sg13g2_decap_8 FILLER_61_3199 ();
 sg13g2_decap_8 FILLER_61_3206 ();
 sg13g2_decap_8 FILLER_61_3213 ();
 sg13g2_decap_8 FILLER_61_3220 ();
 sg13g2_decap_8 FILLER_61_3227 ();
 sg13g2_decap_8 FILLER_61_3234 ();
 sg13g2_decap_8 FILLER_61_3241 ();
 sg13g2_decap_8 FILLER_61_3248 ();
 sg13g2_decap_8 FILLER_61_3255 ();
 sg13g2_decap_8 FILLER_61_3262 ();
 sg13g2_decap_8 FILLER_61_3269 ();
 sg13g2_decap_8 FILLER_61_3276 ();
 sg13g2_decap_8 FILLER_61_3283 ();
 sg13g2_decap_8 FILLER_61_3290 ();
 sg13g2_decap_8 FILLER_61_3297 ();
 sg13g2_decap_8 FILLER_61_3304 ();
 sg13g2_decap_8 FILLER_61_3311 ();
 sg13g2_decap_8 FILLER_61_3318 ();
 sg13g2_decap_8 FILLER_61_3325 ();
 sg13g2_decap_8 FILLER_61_3332 ();
 sg13g2_decap_8 FILLER_61_3339 ();
 sg13g2_decap_8 FILLER_61_3346 ();
 sg13g2_decap_8 FILLER_61_3353 ();
 sg13g2_decap_8 FILLER_61_3360 ();
 sg13g2_decap_8 FILLER_61_3367 ();
 sg13g2_decap_8 FILLER_61_3374 ();
 sg13g2_decap_8 FILLER_61_3381 ();
 sg13g2_decap_8 FILLER_61_3388 ();
 sg13g2_decap_8 FILLER_61_3395 ();
 sg13g2_decap_8 FILLER_61_3402 ();
 sg13g2_decap_8 FILLER_61_3409 ();
 sg13g2_decap_8 FILLER_61_3416 ();
 sg13g2_decap_8 FILLER_61_3423 ();
 sg13g2_decap_8 FILLER_61_3430 ();
 sg13g2_decap_8 FILLER_61_3437 ();
 sg13g2_decap_8 FILLER_61_3444 ();
 sg13g2_decap_8 FILLER_61_3451 ();
 sg13g2_decap_8 FILLER_61_3458 ();
 sg13g2_decap_8 FILLER_61_3465 ();
 sg13g2_decap_8 FILLER_61_3472 ();
 sg13g2_decap_8 FILLER_61_3479 ();
 sg13g2_decap_8 FILLER_61_3486 ();
 sg13g2_decap_8 FILLER_61_3493 ();
 sg13g2_decap_8 FILLER_61_3500 ();
 sg13g2_decap_8 FILLER_61_3507 ();
 sg13g2_decap_8 FILLER_61_3514 ();
 sg13g2_decap_8 FILLER_61_3521 ();
 sg13g2_decap_8 FILLER_61_3528 ();
 sg13g2_decap_8 FILLER_61_3535 ();
 sg13g2_decap_8 FILLER_61_3542 ();
 sg13g2_decap_8 FILLER_61_3549 ();
 sg13g2_decap_8 FILLER_61_3556 ();
 sg13g2_decap_8 FILLER_61_3563 ();
 sg13g2_decap_8 FILLER_61_3570 ();
 sg13g2_fill_2 FILLER_61_3577 ();
 sg13g2_fill_1 FILLER_61_3579 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_8 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_decap_8 FILLER_62_112 ();
 sg13g2_decap_8 FILLER_62_119 ();
 sg13g2_decap_8 FILLER_62_126 ();
 sg13g2_decap_8 FILLER_62_133 ();
 sg13g2_decap_8 FILLER_62_140 ();
 sg13g2_decap_8 FILLER_62_147 ();
 sg13g2_decap_8 FILLER_62_154 ();
 sg13g2_decap_8 FILLER_62_161 ();
 sg13g2_decap_8 FILLER_62_168 ();
 sg13g2_decap_8 FILLER_62_175 ();
 sg13g2_decap_8 FILLER_62_182 ();
 sg13g2_decap_8 FILLER_62_189 ();
 sg13g2_decap_8 FILLER_62_196 ();
 sg13g2_decap_8 FILLER_62_203 ();
 sg13g2_decap_8 FILLER_62_210 ();
 sg13g2_decap_8 FILLER_62_217 ();
 sg13g2_decap_8 FILLER_62_224 ();
 sg13g2_decap_8 FILLER_62_231 ();
 sg13g2_decap_8 FILLER_62_238 ();
 sg13g2_decap_8 FILLER_62_245 ();
 sg13g2_decap_8 FILLER_62_252 ();
 sg13g2_decap_8 FILLER_62_259 ();
 sg13g2_decap_8 FILLER_62_266 ();
 sg13g2_decap_8 FILLER_62_273 ();
 sg13g2_decap_8 FILLER_62_280 ();
 sg13g2_decap_8 FILLER_62_287 ();
 sg13g2_decap_8 FILLER_62_294 ();
 sg13g2_decap_8 FILLER_62_301 ();
 sg13g2_decap_8 FILLER_62_308 ();
 sg13g2_decap_8 FILLER_62_315 ();
 sg13g2_decap_8 FILLER_62_322 ();
 sg13g2_decap_8 FILLER_62_329 ();
 sg13g2_decap_8 FILLER_62_336 ();
 sg13g2_decap_8 FILLER_62_343 ();
 sg13g2_decap_8 FILLER_62_350 ();
 sg13g2_decap_8 FILLER_62_357 ();
 sg13g2_decap_8 FILLER_62_364 ();
 sg13g2_decap_8 FILLER_62_371 ();
 sg13g2_decap_8 FILLER_62_378 ();
 sg13g2_decap_8 FILLER_62_385 ();
 sg13g2_decap_8 FILLER_62_392 ();
 sg13g2_decap_8 FILLER_62_399 ();
 sg13g2_decap_8 FILLER_62_406 ();
 sg13g2_decap_8 FILLER_62_413 ();
 sg13g2_decap_8 FILLER_62_420 ();
 sg13g2_decap_8 FILLER_62_427 ();
 sg13g2_decap_8 FILLER_62_434 ();
 sg13g2_decap_8 FILLER_62_441 ();
 sg13g2_decap_8 FILLER_62_448 ();
 sg13g2_decap_8 FILLER_62_455 ();
 sg13g2_decap_8 FILLER_62_462 ();
 sg13g2_decap_8 FILLER_62_469 ();
 sg13g2_decap_8 FILLER_62_476 ();
 sg13g2_decap_8 FILLER_62_483 ();
 sg13g2_decap_8 FILLER_62_490 ();
 sg13g2_decap_8 FILLER_62_497 ();
 sg13g2_decap_8 FILLER_62_504 ();
 sg13g2_decap_8 FILLER_62_511 ();
 sg13g2_decap_8 FILLER_62_518 ();
 sg13g2_decap_8 FILLER_62_525 ();
 sg13g2_decap_8 FILLER_62_532 ();
 sg13g2_decap_8 FILLER_62_539 ();
 sg13g2_decap_8 FILLER_62_546 ();
 sg13g2_decap_8 FILLER_62_553 ();
 sg13g2_decap_8 FILLER_62_560 ();
 sg13g2_decap_8 FILLER_62_567 ();
 sg13g2_decap_8 FILLER_62_574 ();
 sg13g2_decap_8 FILLER_62_581 ();
 sg13g2_decap_8 FILLER_62_588 ();
 sg13g2_decap_8 FILLER_62_595 ();
 sg13g2_decap_8 FILLER_62_602 ();
 sg13g2_decap_8 FILLER_62_609 ();
 sg13g2_decap_8 FILLER_62_616 ();
 sg13g2_decap_8 FILLER_62_623 ();
 sg13g2_decap_8 FILLER_62_630 ();
 sg13g2_decap_8 FILLER_62_637 ();
 sg13g2_decap_8 FILLER_62_644 ();
 sg13g2_decap_8 FILLER_62_651 ();
 sg13g2_decap_8 FILLER_62_658 ();
 sg13g2_decap_8 FILLER_62_665 ();
 sg13g2_decap_8 FILLER_62_672 ();
 sg13g2_decap_8 FILLER_62_679 ();
 sg13g2_decap_8 FILLER_62_686 ();
 sg13g2_decap_8 FILLER_62_693 ();
 sg13g2_decap_8 FILLER_62_700 ();
 sg13g2_decap_8 FILLER_62_707 ();
 sg13g2_decap_8 FILLER_62_714 ();
 sg13g2_decap_8 FILLER_62_721 ();
 sg13g2_decap_8 FILLER_62_728 ();
 sg13g2_decap_8 FILLER_62_735 ();
 sg13g2_decap_8 FILLER_62_742 ();
 sg13g2_decap_8 FILLER_62_749 ();
 sg13g2_decap_8 FILLER_62_756 ();
 sg13g2_decap_8 FILLER_62_763 ();
 sg13g2_decap_8 FILLER_62_770 ();
 sg13g2_decap_8 FILLER_62_777 ();
 sg13g2_decap_8 FILLER_62_784 ();
 sg13g2_decap_8 FILLER_62_791 ();
 sg13g2_decap_8 FILLER_62_798 ();
 sg13g2_decap_8 FILLER_62_805 ();
 sg13g2_decap_8 FILLER_62_812 ();
 sg13g2_decap_8 FILLER_62_819 ();
 sg13g2_decap_8 FILLER_62_826 ();
 sg13g2_decap_8 FILLER_62_833 ();
 sg13g2_decap_8 FILLER_62_840 ();
 sg13g2_decap_8 FILLER_62_847 ();
 sg13g2_decap_8 FILLER_62_854 ();
 sg13g2_decap_8 FILLER_62_861 ();
 sg13g2_decap_8 FILLER_62_868 ();
 sg13g2_decap_8 FILLER_62_875 ();
 sg13g2_decap_8 FILLER_62_882 ();
 sg13g2_decap_8 FILLER_62_889 ();
 sg13g2_decap_8 FILLER_62_896 ();
 sg13g2_decap_8 FILLER_62_903 ();
 sg13g2_decap_8 FILLER_62_910 ();
 sg13g2_decap_8 FILLER_62_917 ();
 sg13g2_decap_8 FILLER_62_924 ();
 sg13g2_decap_8 FILLER_62_931 ();
 sg13g2_decap_8 FILLER_62_938 ();
 sg13g2_decap_8 FILLER_62_945 ();
 sg13g2_decap_8 FILLER_62_952 ();
 sg13g2_decap_8 FILLER_62_959 ();
 sg13g2_decap_8 FILLER_62_966 ();
 sg13g2_decap_8 FILLER_62_973 ();
 sg13g2_decap_8 FILLER_62_980 ();
 sg13g2_decap_8 FILLER_62_987 ();
 sg13g2_decap_8 FILLER_62_994 ();
 sg13g2_decap_8 FILLER_62_1001 ();
 sg13g2_decap_8 FILLER_62_1008 ();
 sg13g2_decap_8 FILLER_62_1015 ();
 sg13g2_decap_8 FILLER_62_1022 ();
 sg13g2_decap_8 FILLER_62_1029 ();
 sg13g2_decap_8 FILLER_62_1036 ();
 sg13g2_decap_8 FILLER_62_1043 ();
 sg13g2_decap_8 FILLER_62_1050 ();
 sg13g2_decap_8 FILLER_62_1057 ();
 sg13g2_decap_8 FILLER_62_1064 ();
 sg13g2_decap_8 FILLER_62_1071 ();
 sg13g2_decap_8 FILLER_62_1078 ();
 sg13g2_decap_8 FILLER_62_1085 ();
 sg13g2_decap_8 FILLER_62_1092 ();
 sg13g2_decap_8 FILLER_62_1099 ();
 sg13g2_decap_8 FILLER_62_1106 ();
 sg13g2_decap_8 FILLER_62_1113 ();
 sg13g2_decap_8 FILLER_62_1120 ();
 sg13g2_decap_8 FILLER_62_1127 ();
 sg13g2_decap_8 FILLER_62_1134 ();
 sg13g2_decap_8 FILLER_62_1141 ();
 sg13g2_decap_8 FILLER_62_1148 ();
 sg13g2_decap_8 FILLER_62_1155 ();
 sg13g2_decap_8 FILLER_62_1162 ();
 sg13g2_decap_8 FILLER_62_1169 ();
 sg13g2_decap_8 FILLER_62_1176 ();
 sg13g2_decap_8 FILLER_62_1183 ();
 sg13g2_decap_8 FILLER_62_1190 ();
 sg13g2_decap_8 FILLER_62_1197 ();
 sg13g2_decap_8 FILLER_62_1204 ();
 sg13g2_decap_8 FILLER_62_1211 ();
 sg13g2_decap_8 FILLER_62_1218 ();
 sg13g2_decap_8 FILLER_62_1225 ();
 sg13g2_decap_8 FILLER_62_1232 ();
 sg13g2_decap_8 FILLER_62_1239 ();
 sg13g2_decap_8 FILLER_62_1246 ();
 sg13g2_decap_8 FILLER_62_1253 ();
 sg13g2_decap_8 FILLER_62_1260 ();
 sg13g2_decap_8 FILLER_62_1267 ();
 sg13g2_decap_8 FILLER_62_1274 ();
 sg13g2_decap_8 FILLER_62_1281 ();
 sg13g2_decap_8 FILLER_62_1288 ();
 sg13g2_decap_8 FILLER_62_1295 ();
 sg13g2_decap_8 FILLER_62_1302 ();
 sg13g2_decap_8 FILLER_62_1309 ();
 sg13g2_decap_8 FILLER_62_1316 ();
 sg13g2_decap_8 FILLER_62_1323 ();
 sg13g2_decap_8 FILLER_62_1330 ();
 sg13g2_decap_8 FILLER_62_1337 ();
 sg13g2_decap_8 FILLER_62_1344 ();
 sg13g2_decap_8 FILLER_62_1351 ();
 sg13g2_decap_8 FILLER_62_1358 ();
 sg13g2_decap_8 FILLER_62_1365 ();
 sg13g2_decap_8 FILLER_62_1372 ();
 sg13g2_decap_8 FILLER_62_1379 ();
 sg13g2_decap_8 FILLER_62_1386 ();
 sg13g2_decap_8 FILLER_62_1393 ();
 sg13g2_decap_8 FILLER_62_1400 ();
 sg13g2_decap_8 FILLER_62_1407 ();
 sg13g2_decap_8 FILLER_62_1414 ();
 sg13g2_decap_8 FILLER_62_1421 ();
 sg13g2_decap_8 FILLER_62_1428 ();
 sg13g2_decap_8 FILLER_62_1435 ();
 sg13g2_decap_8 FILLER_62_1442 ();
 sg13g2_decap_8 FILLER_62_1449 ();
 sg13g2_decap_8 FILLER_62_1456 ();
 sg13g2_decap_8 FILLER_62_1463 ();
 sg13g2_decap_8 FILLER_62_1470 ();
 sg13g2_decap_8 FILLER_62_1477 ();
 sg13g2_decap_8 FILLER_62_1484 ();
 sg13g2_decap_8 FILLER_62_1491 ();
 sg13g2_decap_8 FILLER_62_1498 ();
 sg13g2_decap_8 FILLER_62_1505 ();
 sg13g2_decap_8 FILLER_62_1512 ();
 sg13g2_decap_8 FILLER_62_1519 ();
 sg13g2_decap_8 FILLER_62_1526 ();
 sg13g2_decap_8 FILLER_62_1533 ();
 sg13g2_decap_8 FILLER_62_1540 ();
 sg13g2_decap_8 FILLER_62_1547 ();
 sg13g2_decap_8 FILLER_62_1554 ();
 sg13g2_decap_8 FILLER_62_1561 ();
 sg13g2_decap_8 FILLER_62_1568 ();
 sg13g2_decap_8 FILLER_62_1575 ();
 sg13g2_decap_8 FILLER_62_1582 ();
 sg13g2_decap_8 FILLER_62_1589 ();
 sg13g2_decap_8 FILLER_62_1596 ();
 sg13g2_decap_8 FILLER_62_1603 ();
 sg13g2_decap_8 FILLER_62_1610 ();
 sg13g2_decap_8 FILLER_62_1617 ();
 sg13g2_decap_8 FILLER_62_1624 ();
 sg13g2_decap_8 FILLER_62_1631 ();
 sg13g2_decap_8 FILLER_62_1638 ();
 sg13g2_decap_8 FILLER_62_1645 ();
 sg13g2_decap_8 FILLER_62_1652 ();
 sg13g2_decap_8 FILLER_62_1659 ();
 sg13g2_decap_8 FILLER_62_1666 ();
 sg13g2_decap_8 FILLER_62_1673 ();
 sg13g2_decap_8 FILLER_62_1680 ();
 sg13g2_decap_8 FILLER_62_1687 ();
 sg13g2_decap_8 FILLER_62_1694 ();
 sg13g2_decap_8 FILLER_62_1701 ();
 sg13g2_decap_8 FILLER_62_1708 ();
 sg13g2_decap_8 FILLER_62_1715 ();
 sg13g2_decap_8 FILLER_62_1722 ();
 sg13g2_decap_8 FILLER_62_1729 ();
 sg13g2_decap_8 FILLER_62_1736 ();
 sg13g2_decap_8 FILLER_62_1743 ();
 sg13g2_decap_8 FILLER_62_1750 ();
 sg13g2_decap_8 FILLER_62_1757 ();
 sg13g2_decap_8 FILLER_62_1764 ();
 sg13g2_decap_8 FILLER_62_1771 ();
 sg13g2_decap_8 FILLER_62_1778 ();
 sg13g2_decap_8 FILLER_62_1785 ();
 sg13g2_decap_8 FILLER_62_1792 ();
 sg13g2_decap_8 FILLER_62_1799 ();
 sg13g2_decap_8 FILLER_62_1806 ();
 sg13g2_decap_8 FILLER_62_1813 ();
 sg13g2_decap_8 FILLER_62_1820 ();
 sg13g2_decap_8 FILLER_62_1827 ();
 sg13g2_decap_8 FILLER_62_1834 ();
 sg13g2_decap_8 FILLER_62_1841 ();
 sg13g2_decap_8 FILLER_62_1848 ();
 sg13g2_decap_8 FILLER_62_1855 ();
 sg13g2_decap_8 FILLER_62_1862 ();
 sg13g2_decap_8 FILLER_62_1869 ();
 sg13g2_decap_8 FILLER_62_1876 ();
 sg13g2_decap_8 FILLER_62_1883 ();
 sg13g2_decap_8 FILLER_62_1890 ();
 sg13g2_decap_8 FILLER_62_1897 ();
 sg13g2_decap_8 FILLER_62_1904 ();
 sg13g2_decap_8 FILLER_62_1911 ();
 sg13g2_decap_8 FILLER_62_1918 ();
 sg13g2_decap_8 FILLER_62_1925 ();
 sg13g2_decap_8 FILLER_62_1932 ();
 sg13g2_decap_8 FILLER_62_1939 ();
 sg13g2_decap_8 FILLER_62_1946 ();
 sg13g2_decap_8 FILLER_62_1953 ();
 sg13g2_decap_8 FILLER_62_1960 ();
 sg13g2_decap_8 FILLER_62_1967 ();
 sg13g2_decap_8 FILLER_62_1974 ();
 sg13g2_decap_8 FILLER_62_1981 ();
 sg13g2_decap_8 FILLER_62_1988 ();
 sg13g2_decap_8 FILLER_62_1995 ();
 sg13g2_decap_8 FILLER_62_2002 ();
 sg13g2_decap_8 FILLER_62_2009 ();
 sg13g2_decap_8 FILLER_62_2016 ();
 sg13g2_decap_8 FILLER_62_2023 ();
 sg13g2_decap_8 FILLER_62_2030 ();
 sg13g2_decap_8 FILLER_62_2037 ();
 sg13g2_decap_8 FILLER_62_2044 ();
 sg13g2_decap_8 FILLER_62_2051 ();
 sg13g2_decap_8 FILLER_62_2058 ();
 sg13g2_decap_8 FILLER_62_2065 ();
 sg13g2_decap_8 FILLER_62_2072 ();
 sg13g2_decap_8 FILLER_62_2079 ();
 sg13g2_decap_8 FILLER_62_2086 ();
 sg13g2_decap_8 FILLER_62_2093 ();
 sg13g2_decap_8 FILLER_62_2100 ();
 sg13g2_decap_8 FILLER_62_2107 ();
 sg13g2_decap_8 FILLER_62_2114 ();
 sg13g2_decap_8 FILLER_62_2121 ();
 sg13g2_decap_8 FILLER_62_2128 ();
 sg13g2_decap_8 FILLER_62_2135 ();
 sg13g2_decap_8 FILLER_62_2142 ();
 sg13g2_decap_8 FILLER_62_2149 ();
 sg13g2_decap_8 FILLER_62_2156 ();
 sg13g2_decap_8 FILLER_62_2163 ();
 sg13g2_decap_8 FILLER_62_2170 ();
 sg13g2_decap_8 FILLER_62_2177 ();
 sg13g2_decap_8 FILLER_62_2184 ();
 sg13g2_decap_8 FILLER_62_2191 ();
 sg13g2_decap_8 FILLER_62_2198 ();
 sg13g2_decap_8 FILLER_62_2205 ();
 sg13g2_decap_8 FILLER_62_2212 ();
 sg13g2_decap_8 FILLER_62_2219 ();
 sg13g2_decap_8 FILLER_62_2226 ();
 sg13g2_decap_8 FILLER_62_2233 ();
 sg13g2_decap_8 FILLER_62_2240 ();
 sg13g2_decap_8 FILLER_62_2247 ();
 sg13g2_decap_8 FILLER_62_2254 ();
 sg13g2_decap_8 FILLER_62_2261 ();
 sg13g2_decap_8 FILLER_62_2268 ();
 sg13g2_decap_8 FILLER_62_2275 ();
 sg13g2_decap_8 FILLER_62_2282 ();
 sg13g2_decap_8 FILLER_62_2289 ();
 sg13g2_decap_8 FILLER_62_2296 ();
 sg13g2_decap_8 FILLER_62_2303 ();
 sg13g2_decap_8 FILLER_62_2310 ();
 sg13g2_decap_8 FILLER_62_2317 ();
 sg13g2_decap_8 FILLER_62_2324 ();
 sg13g2_decap_8 FILLER_62_2331 ();
 sg13g2_decap_8 FILLER_62_2338 ();
 sg13g2_decap_8 FILLER_62_2345 ();
 sg13g2_decap_8 FILLER_62_2352 ();
 sg13g2_decap_8 FILLER_62_2359 ();
 sg13g2_decap_8 FILLER_62_2366 ();
 sg13g2_decap_8 FILLER_62_2373 ();
 sg13g2_decap_8 FILLER_62_2380 ();
 sg13g2_decap_8 FILLER_62_2387 ();
 sg13g2_decap_8 FILLER_62_2394 ();
 sg13g2_decap_8 FILLER_62_2401 ();
 sg13g2_decap_8 FILLER_62_2408 ();
 sg13g2_decap_8 FILLER_62_2415 ();
 sg13g2_decap_8 FILLER_62_2422 ();
 sg13g2_decap_8 FILLER_62_2429 ();
 sg13g2_decap_8 FILLER_62_2436 ();
 sg13g2_decap_8 FILLER_62_2443 ();
 sg13g2_decap_8 FILLER_62_2450 ();
 sg13g2_decap_8 FILLER_62_2457 ();
 sg13g2_decap_8 FILLER_62_2464 ();
 sg13g2_decap_8 FILLER_62_2471 ();
 sg13g2_decap_8 FILLER_62_2478 ();
 sg13g2_decap_8 FILLER_62_2485 ();
 sg13g2_decap_8 FILLER_62_2492 ();
 sg13g2_decap_8 FILLER_62_2499 ();
 sg13g2_decap_8 FILLER_62_2506 ();
 sg13g2_decap_8 FILLER_62_2513 ();
 sg13g2_decap_8 FILLER_62_2520 ();
 sg13g2_decap_8 FILLER_62_2527 ();
 sg13g2_decap_8 FILLER_62_2534 ();
 sg13g2_decap_8 FILLER_62_2541 ();
 sg13g2_decap_8 FILLER_62_2548 ();
 sg13g2_decap_8 FILLER_62_2555 ();
 sg13g2_decap_8 FILLER_62_2562 ();
 sg13g2_decap_8 FILLER_62_2569 ();
 sg13g2_decap_8 FILLER_62_2576 ();
 sg13g2_decap_8 FILLER_62_2583 ();
 sg13g2_decap_8 FILLER_62_2590 ();
 sg13g2_decap_8 FILLER_62_2597 ();
 sg13g2_decap_8 FILLER_62_2604 ();
 sg13g2_decap_8 FILLER_62_2611 ();
 sg13g2_decap_8 FILLER_62_2618 ();
 sg13g2_decap_8 FILLER_62_2625 ();
 sg13g2_decap_8 FILLER_62_2632 ();
 sg13g2_decap_8 FILLER_62_2639 ();
 sg13g2_decap_8 FILLER_62_2646 ();
 sg13g2_decap_8 FILLER_62_2653 ();
 sg13g2_decap_8 FILLER_62_2660 ();
 sg13g2_decap_8 FILLER_62_2667 ();
 sg13g2_decap_8 FILLER_62_2674 ();
 sg13g2_decap_8 FILLER_62_2681 ();
 sg13g2_decap_8 FILLER_62_2688 ();
 sg13g2_decap_8 FILLER_62_2695 ();
 sg13g2_decap_8 FILLER_62_2702 ();
 sg13g2_decap_8 FILLER_62_2709 ();
 sg13g2_decap_8 FILLER_62_2716 ();
 sg13g2_decap_8 FILLER_62_2723 ();
 sg13g2_decap_8 FILLER_62_2730 ();
 sg13g2_decap_8 FILLER_62_2737 ();
 sg13g2_decap_8 FILLER_62_2744 ();
 sg13g2_decap_8 FILLER_62_2751 ();
 sg13g2_decap_8 FILLER_62_2758 ();
 sg13g2_decap_8 FILLER_62_2765 ();
 sg13g2_decap_8 FILLER_62_2772 ();
 sg13g2_decap_8 FILLER_62_2779 ();
 sg13g2_decap_8 FILLER_62_2786 ();
 sg13g2_decap_8 FILLER_62_2793 ();
 sg13g2_decap_8 FILLER_62_2800 ();
 sg13g2_decap_8 FILLER_62_2807 ();
 sg13g2_decap_8 FILLER_62_2814 ();
 sg13g2_decap_8 FILLER_62_2821 ();
 sg13g2_decap_8 FILLER_62_2828 ();
 sg13g2_decap_8 FILLER_62_2835 ();
 sg13g2_decap_8 FILLER_62_2842 ();
 sg13g2_decap_8 FILLER_62_2849 ();
 sg13g2_decap_8 FILLER_62_2856 ();
 sg13g2_decap_8 FILLER_62_2863 ();
 sg13g2_decap_8 FILLER_62_2870 ();
 sg13g2_decap_8 FILLER_62_2877 ();
 sg13g2_decap_8 FILLER_62_2884 ();
 sg13g2_decap_8 FILLER_62_2891 ();
 sg13g2_decap_8 FILLER_62_2898 ();
 sg13g2_decap_8 FILLER_62_2905 ();
 sg13g2_decap_8 FILLER_62_2912 ();
 sg13g2_decap_8 FILLER_62_2919 ();
 sg13g2_decap_8 FILLER_62_2926 ();
 sg13g2_decap_8 FILLER_62_2933 ();
 sg13g2_decap_8 FILLER_62_2940 ();
 sg13g2_decap_8 FILLER_62_2947 ();
 sg13g2_decap_8 FILLER_62_2954 ();
 sg13g2_decap_8 FILLER_62_2961 ();
 sg13g2_decap_8 FILLER_62_2968 ();
 sg13g2_decap_8 FILLER_62_2975 ();
 sg13g2_decap_8 FILLER_62_2982 ();
 sg13g2_decap_8 FILLER_62_2989 ();
 sg13g2_decap_8 FILLER_62_2996 ();
 sg13g2_decap_8 FILLER_62_3003 ();
 sg13g2_decap_8 FILLER_62_3010 ();
 sg13g2_decap_8 FILLER_62_3017 ();
 sg13g2_decap_8 FILLER_62_3024 ();
 sg13g2_decap_8 FILLER_62_3031 ();
 sg13g2_decap_8 FILLER_62_3038 ();
 sg13g2_decap_8 FILLER_62_3045 ();
 sg13g2_decap_8 FILLER_62_3052 ();
 sg13g2_decap_8 FILLER_62_3059 ();
 sg13g2_decap_8 FILLER_62_3066 ();
 sg13g2_decap_8 FILLER_62_3073 ();
 sg13g2_decap_8 FILLER_62_3080 ();
 sg13g2_decap_8 FILLER_62_3087 ();
 sg13g2_decap_8 FILLER_62_3094 ();
 sg13g2_decap_8 FILLER_62_3101 ();
 sg13g2_decap_8 FILLER_62_3108 ();
 sg13g2_decap_8 FILLER_62_3115 ();
 sg13g2_decap_8 FILLER_62_3122 ();
 sg13g2_decap_8 FILLER_62_3129 ();
 sg13g2_decap_8 FILLER_62_3136 ();
 sg13g2_decap_8 FILLER_62_3143 ();
 sg13g2_decap_8 FILLER_62_3150 ();
 sg13g2_decap_8 FILLER_62_3157 ();
 sg13g2_decap_8 FILLER_62_3164 ();
 sg13g2_decap_8 FILLER_62_3171 ();
 sg13g2_decap_8 FILLER_62_3178 ();
 sg13g2_decap_8 FILLER_62_3185 ();
 sg13g2_decap_8 FILLER_62_3192 ();
 sg13g2_decap_8 FILLER_62_3199 ();
 sg13g2_decap_8 FILLER_62_3206 ();
 sg13g2_decap_8 FILLER_62_3213 ();
 sg13g2_decap_8 FILLER_62_3220 ();
 sg13g2_decap_8 FILLER_62_3227 ();
 sg13g2_decap_8 FILLER_62_3234 ();
 sg13g2_decap_8 FILLER_62_3241 ();
 sg13g2_decap_8 FILLER_62_3248 ();
 sg13g2_decap_8 FILLER_62_3255 ();
 sg13g2_decap_8 FILLER_62_3262 ();
 sg13g2_decap_8 FILLER_62_3269 ();
 sg13g2_decap_8 FILLER_62_3276 ();
 sg13g2_decap_8 FILLER_62_3283 ();
 sg13g2_decap_8 FILLER_62_3290 ();
 sg13g2_decap_8 FILLER_62_3297 ();
 sg13g2_decap_8 FILLER_62_3304 ();
 sg13g2_decap_8 FILLER_62_3311 ();
 sg13g2_decap_8 FILLER_62_3318 ();
 sg13g2_decap_8 FILLER_62_3325 ();
 sg13g2_decap_8 FILLER_62_3332 ();
 sg13g2_decap_8 FILLER_62_3339 ();
 sg13g2_decap_8 FILLER_62_3346 ();
 sg13g2_decap_8 FILLER_62_3353 ();
 sg13g2_decap_8 FILLER_62_3360 ();
 sg13g2_decap_8 FILLER_62_3367 ();
 sg13g2_decap_8 FILLER_62_3374 ();
 sg13g2_decap_8 FILLER_62_3381 ();
 sg13g2_decap_8 FILLER_62_3388 ();
 sg13g2_decap_8 FILLER_62_3395 ();
 sg13g2_decap_8 FILLER_62_3402 ();
 sg13g2_decap_8 FILLER_62_3409 ();
 sg13g2_decap_8 FILLER_62_3416 ();
 sg13g2_decap_8 FILLER_62_3423 ();
 sg13g2_decap_8 FILLER_62_3430 ();
 sg13g2_decap_8 FILLER_62_3437 ();
 sg13g2_decap_8 FILLER_62_3444 ();
 sg13g2_decap_8 FILLER_62_3451 ();
 sg13g2_decap_8 FILLER_62_3458 ();
 sg13g2_decap_8 FILLER_62_3465 ();
 sg13g2_decap_8 FILLER_62_3472 ();
 sg13g2_decap_8 FILLER_62_3479 ();
 sg13g2_decap_8 FILLER_62_3486 ();
 sg13g2_decap_8 FILLER_62_3493 ();
 sg13g2_decap_8 FILLER_62_3500 ();
 sg13g2_decap_8 FILLER_62_3507 ();
 sg13g2_decap_8 FILLER_62_3514 ();
 sg13g2_decap_8 FILLER_62_3521 ();
 sg13g2_decap_8 FILLER_62_3528 ();
 sg13g2_decap_8 FILLER_62_3535 ();
 sg13g2_decap_8 FILLER_62_3542 ();
 sg13g2_decap_8 FILLER_62_3549 ();
 sg13g2_decap_8 FILLER_62_3556 ();
 sg13g2_decap_8 FILLER_62_3563 ();
 sg13g2_decap_8 FILLER_62_3570 ();
 sg13g2_fill_2 FILLER_62_3577 ();
 sg13g2_fill_1 FILLER_62_3579 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_decap_8 FILLER_63_105 ();
 sg13g2_decap_8 FILLER_63_112 ();
 sg13g2_decap_8 FILLER_63_119 ();
 sg13g2_decap_8 FILLER_63_126 ();
 sg13g2_decap_8 FILLER_63_133 ();
 sg13g2_decap_8 FILLER_63_140 ();
 sg13g2_decap_8 FILLER_63_147 ();
 sg13g2_decap_8 FILLER_63_154 ();
 sg13g2_decap_8 FILLER_63_161 ();
 sg13g2_decap_8 FILLER_63_168 ();
 sg13g2_decap_8 FILLER_63_175 ();
 sg13g2_decap_8 FILLER_63_182 ();
 sg13g2_decap_8 FILLER_63_189 ();
 sg13g2_decap_8 FILLER_63_196 ();
 sg13g2_decap_8 FILLER_63_203 ();
 sg13g2_decap_8 FILLER_63_210 ();
 sg13g2_decap_8 FILLER_63_217 ();
 sg13g2_decap_8 FILLER_63_224 ();
 sg13g2_decap_8 FILLER_63_231 ();
 sg13g2_decap_8 FILLER_63_238 ();
 sg13g2_decap_8 FILLER_63_245 ();
 sg13g2_decap_8 FILLER_63_252 ();
 sg13g2_decap_8 FILLER_63_259 ();
 sg13g2_decap_8 FILLER_63_266 ();
 sg13g2_decap_8 FILLER_63_273 ();
 sg13g2_decap_8 FILLER_63_280 ();
 sg13g2_decap_8 FILLER_63_287 ();
 sg13g2_decap_8 FILLER_63_294 ();
 sg13g2_decap_8 FILLER_63_301 ();
 sg13g2_decap_8 FILLER_63_308 ();
 sg13g2_decap_8 FILLER_63_315 ();
 sg13g2_decap_8 FILLER_63_322 ();
 sg13g2_decap_8 FILLER_63_329 ();
 sg13g2_decap_8 FILLER_63_336 ();
 sg13g2_decap_8 FILLER_63_343 ();
 sg13g2_decap_8 FILLER_63_350 ();
 sg13g2_decap_8 FILLER_63_357 ();
 sg13g2_decap_8 FILLER_63_364 ();
 sg13g2_decap_8 FILLER_63_371 ();
 sg13g2_decap_8 FILLER_63_378 ();
 sg13g2_decap_8 FILLER_63_385 ();
 sg13g2_decap_8 FILLER_63_392 ();
 sg13g2_decap_8 FILLER_63_399 ();
 sg13g2_decap_8 FILLER_63_406 ();
 sg13g2_decap_8 FILLER_63_413 ();
 sg13g2_decap_8 FILLER_63_420 ();
 sg13g2_decap_8 FILLER_63_427 ();
 sg13g2_decap_8 FILLER_63_434 ();
 sg13g2_decap_8 FILLER_63_441 ();
 sg13g2_decap_8 FILLER_63_448 ();
 sg13g2_decap_8 FILLER_63_455 ();
 sg13g2_decap_8 FILLER_63_462 ();
 sg13g2_decap_8 FILLER_63_469 ();
 sg13g2_decap_8 FILLER_63_476 ();
 sg13g2_decap_8 FILLER_63_483 ();
 sg13g2_decap_8 FILLER_63_490 ();
 sg13g2_decap_8 FILLER_63_497 ();
 sg13g2_decap_8 FILLER_63_504 ();
 sg13g2_decap_8 FILLER_63_511 ();
 sg13g2_decap_8 FILLER_63_518 ();
 sg13g2_decap_8 FILLER_63_525 ();
 sg13g2_decap_8 FILLER_63_532 ();
 sg13g2_decap_8 FILLER_63_539 ();
 sg13g2_decap_8 FILLER_63_546 ();
 sg13g2_decap_8 FILLER_63_553 ();
 sg13g2_decap_8 FILLER_63_560 ();
 sg13g2_decap_8 FILLER_63_567 ();
 sg13g2_decap_8 FILLER_63_574 ();
 sg13g2_decap_8 FILLER_63_581 ();
 sg13g2_decap_8 FILLER_63_588 ();
 sg13g2_decap_8 FILLER_63_595 ();
 sg13g2_decap_8 FILLER_63_602 ();
 sg13g2_decap_8 FILLER_63_609 ();
 sg13g2_decap_8 FILLER_63_616 ();
 sg13g2_decap_8 FILLER_63_623 ();
 sg13g2_decap_8 FILLER_63_630 ();
 sg13g2_decap_8 FILLER_63_637 ();
 sg13g2_decap_8 FILLER_63_644 ();
 sg13g2_decap_8 FILLER_63_651 ();
 sg13g2_decap_8 FILLER_63_658 ();
 sg13g2_decap_8 FILLER_63_665 ();
 sg13g2_decap_8 FILLER_63_672 ();
 sg13g2_decap_8 FILLER_63_679 ();
 sg13g2_decap_8 FILLER_63_686 ();
 sg13g2_decap_8 FILLER_63_693 ();
 sg13g2_decap_8 FILLER_63_700 ();
 sg13g2_decap_8 FILLER_63_707 ();
 sg13g2_decap_8 FILLER_63_714 ();
 sg13g2_decap_8 FILLER_63_721 ();
 sg13g2_decap_8 FILLER_63_728 ();
 sg13g2_decap_8 FILLER_63_735 ();
 sg13g2_decap_8 FILLER_63_742 ();
 sg13g2_decap_8 FILLER_63_749 ();
 sg13g2_decap_8 FILLER_63_756 ();
 sg13g2_decap_8 FILLER_63_763 ();
 sg13g2_decap_8 FILLER_63_770 ();
 sg13g2_decap_8 FILLER_63_777 ();
 sg13g2_decap_8 FILLER_63_784 ();
 sg13g2_decap_8 FILLER_63_791 ();
 sg13g2_decap_8 FILLER_63_798 ();
 sg13g2_decap_8 FILLER_63_805 ();
 sg13g2_decap_8 FILLER_63_812 ();
 sg13g2_decap_8 FILLER_63_819 ();
 sg13g2_decap_8 FILLER_63_826 ();
 sg13g2_decap_8 FILLER_63_833 ();
 sg13g2_decap_8 FILLER_63_840 ();
 sg13g2_decap_8 FILLER_63_847 ();
 sg13g2_decap_8 FILLER_63_854 ();
 sg13g2_decap_8 FILLER_63_861 ();
 sg13g2_decap_8 FILLER_63_868 ();
 sg13g2_decap_8 FILLER_63_875 ();
 sg13g2_decap_8 FILLER_63_882 ();
 sg13g2_decap_8 FILLER_63_889 ();
 sg13g2_decap_8 FILLER_63_896 ();
 sg13g2_decap_8 FILLER_63_903 ();
 sg13g2_decap_8 FILLER_63_910 ();
 sg13g2_decap_8 FILLER_63_917 ();
 sg13g2_decap_8 FILLER_63_924 ();
 sg13g2_decap_8 FILLER_63_931 ();
 sg13g2_decap_8 FILLER_63_938 ();
 sg13g2_decap_8 FILLER_63_945 ();
 sg13g2_decap_8 FILLER_63_952 ();
 sg13g2_decap_8 FILLER_63_959 ();
 sg13g2_decap_8 FILLER_63_966 ();
 sg13g2_decap_8 FILLER_63_973 ();
 sg13g2_decap_8 FILLER_63_980 ();
 sg13g2_decap_8 FILLER_63_987 ();
 sg13g2_decap_8 FILLER_63_994 ();
 sg13g2_decap_8 FILLER_63_1001 ();
 sg13g2_decap_8 FILLER_63_1008 ();
 sg13g2_decap_8 FILLER_63_1015 ();
 sg13g2_decap_8 FILLER_63_1022 ();
 sg13g2_decap_8 FILLER_63_1029 ();
 sg13g2_decap_8 FILLER_63_1036 ();
 sg13g2_decap_8 FILLER_63_1043 ();
 sg13g2_decap_8 FILLER_63_1050 ();
 sg13g2_decap_8 FILLER_63_1057 ();
 sg13g2_decap_8 FILLER_63_1064 ();
 sg13g2_decap_8 FILLER_63_1071 ();
 sg13g2_decap_8 FILLER_63_1078 ();
 sg13g2_decap_8 FILLER_63_1085 ();
 sg13g2_decap_8 FILLER_63_1092 ();
 sg13g2_decap_8 FILLER_63_1099 ();
 sg13g2_decap_8 FILLER_63_1106 ();
 sg13g2_decap_8 FILLER_63_1113 ();
 sg13g2_decap_8 FILLER_63_1120 ();
 sg13g2_decap_8 FILLER_63_1127 ();
 sg13g2_decap_8 FILLER_63_1134 ();
 sg13g2_decap_8 FILLER_63_1141 ();
 sg13g2_decap_8 FILLER_63_1148 ();
 sg13g2_decap_8 FILLER_63_1155 ();
 sg13g2_decap_8 FILLER_63_1162 ();
 sg13g2_decap_8 FILLER_63_1169 ();
 sg13g2_decap_8 FILLER_63_1176 ();
 sg13g2_decap_8 FILLER_63_1183 ();
 sg13g2_decap_8 FILLER_63_1190 ();
 sg13g2_decap_8 FILLER_63_1197 ();
 sg13g2_decap_8 FILLER_63_1204 ();
 sg13g2_decap_8 FILLER_63_1211 ();
 sg13g2_decap_8 FILLER_63_1218 ();
 sg13g2_decap_8 FILLER_63_1225 ();
 sg13g2_decap_8 FILLER_63_1232 ();
 sg13g2_decap_8 FILLER_63_1239 ();
 sg13g2_decap_8 FILLER_63_1246 ();
 sg13g2_decap_8 FILLER_63_1253 ();
 sg13g2_decap_8 FILLER_63_1260 ();
 sg13g2_decap_8 FILLER_63_1267 ();
 sg13g2_decap_8 FILLER_63_1274 ();
 sg13g2_decap_8 FILLER_63_1281 ();
 sg13g2_decap_8 FILLER_63_1288 ();
 sg13g2_decap_8 FILLER_63_1295 ();
 sg13g2_decap_8 FILLER_63_1302 ();
 sg13g2_decap_8 FILLER_63_1309 ();
 sg13g2_decap_8 FILLER_63_1316 ();
 sg13g2_decap_8 FILLER_63_1323 ();
 sg13g2_decap_8 FILLER_63_1330 ();
 sg13g2_decap_8 FILLER_63_1337 ();
 sg13g2_decap_8 FILLER_63_1344 ();
 sg13g2_decap_8 FILLER_63_1351 ();
 sg13g2_decap_8 FILLER_63_1358 ();
 sg13g2_decap_8 FILLER_63_1365 ();
 sg13g2_decap_8 FILLER_63_1372 ();
 sg13g2_decap_8 FILLER_63_1379 ();
 sg13g2_decap_8 FILLER_63_1386 ();
 sg13g2_decap_8 FILLER_63_1393 ();
 sg13g2_decap_8 FILLER_63_1400 ();
 sg13g2_decap_8 FILLER_63_1407 ();
 sg13g2_decap_8 FILLER_63_1414 ();
 sg13g2_decap_8 FILLER_63_1421 ();
 sg13g2_decap_8 FILLER_63_1428 ();
 sg13g2_decap_8 FILLER_63_1435 ();
 sg13g2_decap_8 FILLER_63_1442 ();
 sg13g2_decap_8 FILLER_63_1449 ();
 sg13g2_decap_8 FILLER_63_1456 ();
 sg13g2_decap_8 FILLER_63_1463 ();
 sg13g2_decap_8 FILLER_63_1470 ();
 sg13g2_decap_8 FILLER_63_1477 ();
 sg13g2_decap_8 FILLER_63_1484 ();
 sg13g2_decap_8 FILLER_63_1491 ();
 sg13g2_decap_8 FILLER_63_1498 ();
 sg13g2_decap_8 FILLER_63_1505 ();
 sg13g2_decap_8 FILLER_63_1512 ();
 sg13g2_decap_8 FILLER_63_1519 ();
 sg13g2_decap_8 FILLER_63_1526 ();
 sg13g2_decap_8 FILLER_63_1533 ();
 sg13g2_decap_8 FILLER_63_1540 ();
 sg13g2_decap_8 FILLER_63_1547 ();
 sg13g2_decap_8 FILLER_63_1554 ();
 sg13g2_decap_8 FILLER_63_1561 ();
 sg13g2_decap_8 FILLER_63_1568 ();
 sg13g2_decap_8 FILLER_63_1575 ();
 sg13g2_decap_8 FILLER_63_1582 ();
 sg13g2_decap_8 FILLER_63_1589 ();
 sg13g2_decap_8 FILLER_63_1596 ();
 sg13g2_decap_8 FILLER_63_1603 ();
 sg13g2_decap_8 FILLER_63_1610 ();
 sg13g2_decap_8 FILLER_63_1617 ();
 sg13g2_decap_8 FILLER_63_1624 ();
 sg13g2_decap_8 FILLER_63_1631 ();
 sg13g2_decap_8 FILLER_63_1638 ();
 sg13g2_decap_8 FILLER_63_1645 ();
 sg13g2_decap_8 FILLER_63_1652 ();
 sg13g2_decap_8 FILLER_63_1659 ();
 sg13g2_decap_8 FILLER_63_1666 ();
 sg13g2_decap_8 FILLER_63_1673 ();
 sg13g2_decap_8 FILLER_63_1680 ();
 sg13g2_decap_8 FILLER_63_1687 ();
 sg13g2_decap_8 FILLER_63_1694 ();
 sg13g2_decap_8 FILLER_63_1701 ();
 sg13g2_decap_8 FILLER_63_1708 ();
 sg13g2_decap_8 FILLER_63_1715 ();
 sg13g2_decap_8 FILLER_63_1722 ();
 sg13g2_decap_8 FILLER_63_1729 ();
 sg13g2_decap_8 FILLER_63_1736 ();
 sg13g2_decap_8 FILLER_63_1743 ();
 sg13g2_decap_8 FILLER_63_1750 ();
 sg13g2_decap_8 FILLER_63_1757 ();
 sg13g2_decap_8 FILLER_63_1764 ();
 sg13g2_decap_8 FILLER_63_1771 ();
 sg13g2_decap_8 FILLER_63_1778 ();
 sg13g2_decap_8 FILLER_63_1785 ();
 sg13g2_decap_8 FILLER_63_1792 ();
 sg13g2_decap_8 FILLER_63_1799 ();
 sg13g2_decap_8 FILLER_63_1806 ();
 sg13g2_decap_8 FILLER_63_1813 ();
 sg13g2_decap_8 FILLER_63_1820 ();
 sg13g2_decap_8 FILLER_63_1827 ();
 sg13g2_decap_8 FILLER_63_1834 ();
 sg13g2_decap_8 FILLER_63_1841 ();
 sg13g2_decap_8 FILLER_63_1848 ();
 sg13g2_decap_8 FILLER_63_1855 ();
 sg13g2_decap_8 FILLER_63_1862 ();
 sg13g2_decap_8 FILLER_63_1869 ();
 sg13g2_decap_8 FILLER_63_1876 ();
 sg13g2_decap_8 FILLER_63_1883 ();
 sg13g2_decap_8 FILLER_63_1890 ();
 sg13g2_decap_8 FILLER_63_1897 ();
 sg13g2_decap_8 FILLER_63_1904 ();
 sg13g2_decap_8 FILLER_63_1911 ();
 sg13g2_decap_8 FILLER_63_1918 ();
 sg13g2_decap_8 FILLER_63_1925 ();
 sg13g2_decap_8 FILLER_63_1932 ();
 sg13g2_decap_8 FILLER_63_1939 ();
 sg13g2_decap_8 FILLER_63_1946 ();
 sg13g2_decap_8 FILLER_63_1953 ();
 sg13g2_decap_8 FILLER_63_1960 ();
 sg13g2_decap_8 FILLER_63_1967 ();
 sg13g2_decap_8 FILLER_63_1974 ();
 sg13g2_decap_8 FILLER_63_1981 ();
 sg13g2_decap_8 FILLER_63_1988 ();
 sg13g2_decap_8 FILLER_63_1995 ();
 sg13g2_decap_8 FILLER_63_2002 ();
 sg13g2_decap_8 FILLER_63_2009 ();
 sg13g2_decap_8 FILLER_63_2016 ();
 sg13g2_decap_8 FILLER_63_2023 ();
 sg13g2_decap_8 FILLER_63_2030 ();
 sg13g2_decap_8 FILLER_63_2037 ();
 sg13g2_decap_8 FILLER_63_2044 ();
 sg13g2_decap_8 FILLER_63_2051 ();
 sg13g2_decap_8 FILLER_63_2058 ();
 sg13g2_decap_8 FILLER_63_2065 ();
 sg13g2_decap_8 FILLER_63_2072 ();
 sg13g2_decap_8 FILLER_63_2079 ();
 sg13g2_decap_8 FILLER_63_2086 ();
 sg13g2_decap_8 FILLER_63_2093 ();
 sg13g2_decap_8 FILLER_63_2100 ();
 sg13g2_decap_8 FILLER_63_2107 ();
 sg13g2_decap_8 FILLER_63_2114 ();
 sg13g2_decap_8 FILLER_63_2121 ();
 sg13g2_decap_8 FILLER_63_2128 ();
 sg13g2_decap_8 FILLER_63_2135 ();
 sg13g2_decap_8 FILLER_63_2142 ();
 sg13g2_decap_8 FILLER_63_2149 ();
 sg13g2_decap_8 FILLER_63_2156 ();
 sg13g2_decap_8 FILLER_63_2163 ();
 sg13g2_decap_8 FILLER_63_2170 ();
 sg13g2_decap_8 FILLER_63_2177 ();
 sg13g2_decap_8 FILLER_63_2184 ();
 sg13g2_decap_8 FILLER_63_2191 ();
 sg13g2_decap_8 FILLER_63_2198 ();
 sg13g2_decap_8 FILLER_63_2205 ();
 sg13g2_decap_8 FILLER_63_2212 ();
 sg13g2_decap_8 FILLER_63_2219 ();
 sg13g2_decap_8 FILLER_63_2226 ();
 sg13g2_decap_8 FILLER_63_2233 ();
 sg13g2_decap_8 FILLER_63_2240 ();
 sg13g2_decap_8 FILLER_63_2247 ();
 sg13g2_decap_8 FILLER_63_2254 ();
 sg13g2_decap_8 FILLER_63_2261 ();
 sg13g2_decap_8 FILLER_63_2268 ();
 sg13g2_decap_8 FILLER_63_2275 ();
 sg13g2_decap_8 FILLER_63_2282 ();
 sg13g2_decap_8 FILLER_63_2289 ();
 sg13g2_decap_8 FILLER_63_2296 ();
 sg13g2_decap_8 FILLER_63_2303 ();
 sg13g2_decap_8 FILLER_63_2310 ();
 sg13g2_decap_8 FILLER_63_2317 ();
 sg13g2_decap_8 FILLER_63_2324 ();
 sg13g2_decap_8 FILLER_63_2331 ();
 sg13g2_decap_8 FILLER_63_2338 ();
 sg13g2_decap_8 FILLER_63_2345 ();
 sg13g2_decap_8 FILLER_63_2352 ();
 sg13g2_decap_8 FILLER_63_2359 ();
 sg13g2_decap_8 FILLER_63_2366 ();
 sg13g2_decap_8 FILLER_63_2373 ();
 sg13g2_decap_8 FILLER_63_2380 ();
 sg13g2_decap_8 FILLER_63_2387 ();
 sg13g2_decap_8 FILLER_63_2394 ();
 sg13g2_decap_8 FILLER_63_2401 ();
 sg13g2_decap_8 FILLER_63_2408 ();
 sg13g2_decap_8 FILLER_63_2415 ();
 sg13g2_decap_8 FILLER_63_2422 ();
 sg13g2_decap_8 FILLER_63_2429 ();
 sg13g2_decap_8 FILLER_63_2436 ();
 sg13g2_decap_8 FILLER_63_2443 ();
 sg13g2_decap_8 FILLER_63_2450 ();
 sg13g2_decap_8 FILLER_63_2457 ();
 sg13g2_decap_8 FILLER_63_2464 ();
 sg13g2_decap_8 FILLER_63_2471 ();
 sg13g2_decap_8 FILLER_63_2478 ();
 sg13g2_decap_8 FILLER_63_2485 ();
 sg13g2_decap_8 FILLER_63_2492 ();
 sg13g2_decap_8 FILLER_63_2499 ();
 sg13g2_decap_8 FILLER_63_2506 ();
 sg13g2_decap_8 FILLER_63_2513 ();
 sg13g2_decap_8 FILLER_63_2520 ();
 sg13g2_decap_8 FILLER_63_2527 ();
 sg13g2_decap_8 FILLER_63_2534 ();
 sg13g2_decap_8 FILLER_63_2541 ();
 sg13g2_decap_8 FILLER_63_2548 ();
 sg13g2_decap_8 FILLER_63_2555 ();
 sg13g2_decap_8 FILLER_63_2562 ();
 sg13g2_decap_8 FILLER_63_2569 ();
 sg13g2_decap_8 FILLER_63_2576 ();
 sg13g2_decap_8 FILLER_63_2583 ();
 sg13g2_decap_8 FILLER_63_2590 ();
 sg13g2_decap_8 FILLER_63_2597 ();
 sg13g2_decap_8 FILLER_63_2604 ();
 sg13g2_decap_8 FILLER_63_2611 ();
 sg13g2_decap_8 FILLER_63_2618 ();
 sg13g2_decap_8 FILLER_63_2625 ();
 sg13g2_decap_8 FILLER_63_2632 ();
 sg13g2_decap_8 FILLER_63_2639 ();
 sg13g2_decap_8 FILLER_63_2646 ();
 sg13g2_decap_8 FILLER_63_2653 ();
 sg13g2_decap_8 FILLER_63_2660 ();
 sg13g2_decap_8 FILLER_63_2667 ();
 sg13g2_decap_8 FILLER_63_2674 ();
 sg13g2_decap_8 FILLER_63_2681 ();
 sg13g2_decap_8 FILLER_63_2688 ();
 sg13g2_decap_8 FILLER_63_2695 ();
 sg13g2_decap_8 FILLER_63_2702 ();
 sg13g2_decap_8 FILLER_63_2709 ();
 sg13g2_decap_8 FILLER_63_2716 ();
 sg13g2_decap_8 FILLER_63_2723 ();
 sg13g2_decap_8 FILLER_63_2730 ();
 sg13g2_decap_8 FILLER_63_2737 ();
 sg13g2_decap_8 FILLER_63_2744 ();
 sg13g2_decap_8 FILLER_63_2751 ();
 sg13g2_decap_8 FILLER_63_2758 ();
 sg13g2_decap_8 FILLER_63_2765 ();
 sg13g2_decap_8 FILLER_63_2772 ();
 sg13g2_decap_8 FILLER_63_2779 ();
 sg13g2_decap_8 FILLER_63_2786 ();
 sg13g2_decap_8 FILLER_63_2793 ();
 sg13g2_decap_8 FILLER_63_2800 ();
 sg13g2_decap_8 FILLER_63_2807 ();
 sg13g2_decap_8 FILLER_63_2814 ();
 sg13g2_decap_8 FILLER_63_2821 ();
 sg13g2_decap_8 FILLER_63_2828 ();
 sg13g2_decap_8 FILLER_63_2835 ();
 sg13g2_decap_8 FILLER_63_2842 ();
 sg13g2_decap_8 FILLER_63_2849 ();
 sg13g2_decap_8 FILLER_63_2856 ();
 sg13g2_decap_8 FILLER_63_2863 ();
 sg13g2_decap_8 FILLER_63_2870 ();
 sg13g2_decap_8 FILLER_63_2877 ();
 sg13g2_decap_8 FILLER_63_2884 ();
 sg13g2_decap_8 FILLER_63_2891 ();
 sg13g2_decap_8 FILLER_63_2898 ();
 sg13g2_decap_8 FILLER_63_2905 ();
 sg13g2_decap_8 FILLER_63_2912 ();
 sg13g2_decap_8 FILLER_63_2919 ();
 sg13g2_decap_8 FILLER_63_2926 ();
 sg13g2_decap_8 FILLER_63_2933 ();
 sg13g2_decap_8 FILLER_63_2940 ();
 sg13g2_decap_8 FILLER_63_2947 ();
 sg13g2_decap_8 FILLER_63_2954 ();
 sg13g2_decap_8 FILLER_63_2961 ();
 sg13g2_decap_8 FILLER_63_2968 ();
 sg13g2_decap_8 FILLER_63_2975 ();
 sg13g2_decap_8 FILLER_63_2982 ();
 sg13g2_decap_8 FILLER_63_2989 ();
 sg13g2_decap_8 FILLER_63_2996 ();
 sg13g2_decap_8 FILLER_63_3003 ();
 sg13g2_decap_8 FILLER_63_3010 ();
 sg13g2_decap_8 FILLER_63_3017 ();
 sg13g2_decap_8 FILLER_63_3024 ();
 sg13g2_decap_8 FILLER_63_3031 ();
 sg13g2_decap_8 FILLER_63_3038 ();
 sg13g2_decap_8 FILLER_63_3045 ();
 sg13g2_decap_8 FILLER_63_3052 ();
 sg13g2_decap_8 FILLER_63_3059 ();
 sg13g2_decap_8 FILLER_63_3066 ();
 sg13g2_decap_8 FILLER_63_3073 ();
 sg13g2_decap_8 FILLER_63_3080 ();
 sg13g2_decap_8 FILLER_63_3087 ();
 sg13g2_decap_8 FILLER_63_3094 ();
 sg13g2_decap_8 FILLER_63_3101 ();
 sg13g2_decap_8 FILLER_63_3108 ();
 sg13g2_decap_8 FILLER_63_3115 ();
 sg13g2_decap_8 FILLER_63_3122 ();
 sg13g2_decap_8 FILLER_63_3129 ();
 sg13g2_decap_8 FILLER_63_3136 ();
 sg13g2_decap_8 FILLER_63_3143 ();
 sg13g2_decap_8 FILLER_63_3150 ();
 sg13g2_decap_8 FILLER_63_3157 ();
 sg13g2_decap_8 FILLER_63_3164 ();
 sg13g2_decap_8 FILLER_63_3171 ();
 sg13g2_decap_8 FILLER_63_3178 ();
 sg13g2_decap_8 FILLER_63_3185 ();
 sg13g2_decap_8 FILLER_63_3192 ();
 sg13g2_decap_8 FILLER_63_3199 ();
 sg13g2_decap_8 FILLER_63_3206 ();
 sg13g2_decap_8 FILLER_63_3213 ();
 sg13g2_decap_8 FILLER_63_3220 ();
 sg13g2_decap_8 FILLER_63_3227 ();
 sg13g2_decap_8 FILLER_63_3234 ();
 sg13g2_decap_8 FILLER_63_3241 ();
 sg13g2_decap_8 FILLER_63_3248 ();
 sg13g2_decap_8 FILLER_63_3255 ();
 sg13g2_decap_8 FILLER_63_3262 ();
 sg13g2_decap_8 FILLER_63_3269 ();
 sg13g2_decap_8 FILLER_63_3276 ();
 sg13g2_decap_8 FILLER_63_3283 ();
 sg13g2_decap_8 FILLER_63_3290 ();
 sg13g2_decap_8 FILLER_63_3297 ();
 sg13g2_decap_8 FILLER_63_3304 ();
 sg13g2_decap_8 FILLER_63_3311 ();
 sg13g2_decap_8 FILLER_63_3318 ();
 sg13g2_decap_8 FILLER_63_3325 ();
 sg13g2_decap_8 FILLER_63_3332 ();
 sg13g2_decap_8 FILLER_63_3339 ();
 sg13g2_decap_8 FILLER_63_3346 ();
 sg13g2_decap_8 FILLER_63_3353 ();
 sg13g2_decap_8 FILLER_63_3360 ();
 sg13g2_decap_8 FILLER_63_3367 ();
 sg13g2_decap_8 FILLER_63_3374 ();
 sg13g2_decap_8 FILLER_63_3381 ();
 sg13g2_decap_8 FILLER_63_3388 ();
 sg13g2_decap_8 FILLER_63_3395 ();
 sg13g2_decap_8 FILLER_63_3402 ();
 sg13g2_decap_8 FILLER_63_3409 ();
 sg13g2_decap_8 FILLER_63_3416 ();
 sg13g2_decap_8 FILLER_63_3423 ();
 sg13g2_decap_8 FILLER_63_3430 ();
 sg13g2_decap_8 FILLER_63_3437 ();
 sg13g2_decap_8 FILLER_63_3444 ();
 sg13g2_decap_8 FILLER_63_3451 ();
 sg13g2_decap_8 FILLER_63_3458 ();
 sg13g2_decap_8 FILLER_63_3465 ();
 sg13g2_decap_8 FILLER_63_3472 ();
 sg13g2_decap_8 FILLER_63_3479 ();
 sg13g2_decap_8 FILLER_63_3486 ();
 sg13g2_decap_8 FILLER_63_3493 ();
 sg13g2_decap_8 FILLER_63_3500 ();
 sg13g2_decap_8 FILLER_63_3507 ();
 sg13g2_decap_8 FILLER_63_3514 ();
 sg13g2_decap_8 FILLER_63_3521 ();
 sg13g2_decap_8 FILLER_63_3528 ();
 sg13g2_decap_8 FILLER_63_3535 ();
 sg13g2_decap_8 FILLER_63_3542 ();
 sg13g2_decap_8 FILLER_63_3549 ();
 sg13g2_decap_8 FILLER_63_3556 ();
 sg13g2_decap_8 FILLER_63_3563 ();
 sg13g2_decap_8 FILLER_63_3570 ();
 sg13g2_fill_2 FILLER_63_3577 ();
 sg13g2_fill_1 FILLER_63_3579 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_decap_8 FILLER_64_112 ();
 sg13g2_decap_8 FILLER_64_119 ();
 sg13g2_decap_8 FILLER_64_126 ();
 sg13g2_decap_8 FILLER_64_133 ();
 sg13g2_decap_8 FILLER_64_140 ();
 sg13g2_decap_8 FILLER_64_147 ();
 sg13g2_decap_8 FILLER_64_154 ();
 sg13g2_decap_8 FILLER_64_161 ();
 sg13g2_decap_8 FILLER_64_168 ();
 sg13g2_decap_8 FILLER_64_175 ();
 sg13g2_decap_8 FILLER_64_182 ();
 sg13g2_decap_8 FILLER_64_189 ();
 sg13g2_decap_8 FILLER_64_196 ();
 sg13g2_decap_8 FILLER_64_203 ();
 sg13g2_decap_8 FILLER_64_210 ();
 sg13g2_decap_8 FILLER_64_217 ();
 sg13g2_decap_8 FILLER_64_224 ();
 sg13g2_decap_8 FILLER_64_231 ();
 sg13g2_decap_8 FILLER_64_238 ();
 sg13g2_decap_8 FILLER_64_245 ();
 sg13g2_decap_8 FILLER_64_252 ();
 sg13g2_decap_8 FILLER_64_259 ();
 sg13g2_decap_8 FILLER_64_266 ();
 sg13g2_decap_8 FILLER_64_273 ();
 sg13g2_decap_8 FILLER_64_280 ();
 sg13g2_decap_8 FILLER_64_287 ();
 sg13g2_decap_8 FILLER_64_294 ();
 sg13g2_decap_8 FILLER_64_301 ();
 sg13g2_decap_8 FILLER_64_308 ();
 sg13g2_decap_8 FILLER_64_315 ();
 sg13g2_decap_8 FILLER_64_322 ();
 sg13g2_decap_8 FILLER_64_329 ();
 sg13g2_decap_8 FILLER_64_336 ();
 sg13g2_decap_8 FILLER_64_343 ();
 sg13g2_decap_8 FILLER_64_350 ();
 sg13g2_decap_8 FILLER_64_357 ();
 sg13g2_decap_8 FILLER_64_364 ();
 sg13g2_decap_8 FILLER_64_371 ();
 sg13g2_decap_8 FILLER_64_378 ();
 sg13g2_decap_8 FILLER_64_385 ();
 sg13g2_decap_8 FILLER_64_392 ();
 sg13g2_decap_8 FILLER_64_399 ();
 sg13g2_decap_8 FILLER_64_406 ();
 sg13g2_decap_8 FILLER_64_413 ();
 sg13g2_decap_8 FILLER_64_420 ();
 sg13g2_decap_8 FILLER_64_427 ();
 sg13g2_decap_8 FILLER_64_434 ();
 sg13g2_decap_8 FILLER_64_441 ();
 sg13g2_decap_8 FILLER_64_448 ();
 sg13g2_decap_8 FILLER_64_455 ();
 sg13g2_decap_8 FILLER_64_462 ();
 sg13g2_decap_8 FILLER_64_469 ();
 sg13g2_decap_8 FILLER_64_476 ();
 sg13g2_decap_8 FILLER_64_483 ();
 sg13g2_decap_8 FILLER_64_490 ();
 sg13g2_decap_8 FILLER_64_497 ();
 sg13g2_decap_8 FILLER_64_504 ();
 sg13g2_decap_8 FILLER_64_511 ();
 sg13g2_decap_8 FILLER_64_518 ();
 sg13g2_decap_8 FILLER_64_525 ();
 sg13g2_decap_8 FILLER_64_532 ();
 sg13g2_decap_8 FILLER_64_539 ();
 sg13g2_decap_8 FILLER_64_546 ();
 sg13g2_decap_8 FILLER_64_553 ();
 sg13g2_decap_8 FILLER_64_560 ();
 sg13g2_decap_8 FILLER_64_567 ();
 sg13g2_decap_8 FILLER_64_574 ();
 sg13g2_decap_8 FILLER_64_581 ();
 sg13g2_decap_8 FILLER_64_588 ();
 sg13g2_decap_8 FILLER_64_595 ();
 sg13g2_decap_8 FILLER_64_602 ();
 sg13g2_decap_8 FILLER_64_609 ();
 sg13g2_decap_8 FILLER_64_616 ();
 sg13g2_decap_8 FILLER_64_623 ();
 sg13g2_decap_8 FILLER_64_630 ();
 sg13g2_decap_8 FILLER_64_637 ();
 sg13g2_decap_8 FILLER_64_644 ();
 sg13g2_decap_8 FILLER_64_651 ();
 sg13g2_decap_8 FILLER_64_658 ();
 sg13g2_decap_8 FILLER_64_665 ();
 sg13g2_decap_8 FILLER_64_672 ();
 sg13g2_decap_8 FILLER_64_679 ();
 sg13g2_decap_8 FILLER_64_686 ();
 sg13g2_decap_8 FILLER_64_693 ();
 sg13g2_decap_8 FILLER_64_700 ();
 sg13g2_decap_8 FILLER_64_707 ();
 sg13g2_decap_8 FILLER_64_714 ();
 sg13g2_decap_8 FILLER_64_721 ();
 sg13g2_decap_8 FILLER_64_728 ();
 sg13g2_decap_8 FILLER_64_735 ();
 sg13g2_decap_8 FILLER_64_742 ();
 sg13g2_decap_8 FILLER_64_749 ();
 sg13g2_decap_8 FILLER_64_756 ();
 sg13g2_decap_8 FILLER_64_763 ();
 sg13g2_decap_8 FILLER_64_770 ();
 sg13g2_decap_8 FILLER_64_777 ();
 sg13g2_decap_8 FILLER_64_784 ();
 sg13g2_decap_8 FILLER_64_791 ();
 sg13g2_decap_8 FILLER_64_798 ();
 sg13g2_decap_8 FILLER_64_805 ();
 sg13g2_decap_8 FILLER_64_812 ();
 sg13g2_decap_8 FILLER_64_819 ();
 sg13g2_decap_8 FILLER_64_826 ();
 sg13g2_decap_8 FILLER_64_833 ();
 sg13g2_decap_8 FILLER_64_840 ();
 sg13g2_decap_8 FILLER_64_847 ();
 sg13g2_decap_8 FILLER_64_854 ();
 sg13g2_decap_8 FILLER_64_861 ();
 sg13g2_decap_8 FILLER_64_868 ();
 sg13g2_decap_8 FILLER_64_875 ();
 sg13g2_decap_8 FILLER_64_882 ();
 sg13g2_decap_8 FILLER_64_889 ();
 sg13g2_decap_8 FILLER_64_896 ();
 sg13g2_decap_8 FILLER_64_903 ();
 sg13g2_decap_8 FILLER_64_910 ();
 sg13g2_decap_8 FILLER_64_917 ();
 sg13g2_decap_8 FILLER_64_924 ();
 sg13g2_decap_8 FILLER_64_931 ();
 sg13g2_decap_8 FILLER_64_938 ();
 sg13g2_decap_8 FILLER_64_945 ();
 sg13g2_decap_8 FILLER_64_952 ();
 sg13g2_decap_8 FILLER_64_959 ();
 sg13g2_decap_8 FILLER_64_966 ();
 sg13g2_decap_8 FILLER_64_973 ();
 sg13g2_decap_8 FILLER_64_980 ();
 sg13g2_decap_8 FILLER_64_987 ();
 sg13g2_decap_8 FILLER_64_994 ();
 sg13g2_decap_8 FILLER_64_1001 ();
 sg13g2_decap_8 FILLER_64_1008 ();
 sg13g2_decap_8 FILLER_64_1015 ();
 sg13g2_decap_8 FILLER_64_1022 ();
 sg13g2_decap_8 FILLER_64_1029 ();
 sg13g2_decap_8 FILLER_64_1036 ();
 sg13g2_decap_8 FILLER_64_1043 ();
 sg13g2_decap_8 FILLER_64_1050 ();
 sg13g2_decap_8 FILLER_64_1057 ();
 sg13g2_decap_8 FILLER_64_1064 ();
 sg13g2_decap_8 FILLER_64_1071 ();
 sg13g2_decap_8 FILLER_64_1078 ();
 sg13g2_decap_8 FILLER_64_1085 ();
 sg13g2_decap_8 FILLER_64_1092 ();
 sg13g2_decap_8 FILLER_64_1099 ();
 sg13g2_decap_8 FILLER_64_1106 ();
 sg13g2_decap_8 FILLER_64_1113 ();
 sg13g2_decap_8 FILLER_64_1120 ();
 sg13g2_decap_8 FILLER_64_1127 ();
 sg13g2_decap_8 FILLER_64_1134 ();
 sg13g2_decap_8 FILLER_64_1141 ();
 sg13g2_decap_8 FILLER_64_1148 ();
 sg13g2_decap_8 FILLER_64_1155 ();
 sg13g2_decap_8 FILLER_64_1162 ();
 sg13g2_decap_8 FILLER_64_1169 ();
 sg13g2_decap_8 FILLER_64_1176 ();
 sg13g2_decap_8 FILLER_64_1183 ();
 sg13g2_decap_8 FILLER_64_1190 ();
 sg13g2_decap_8 FILLER_64_1197 ();
 sg13g2_decap_8 FILLER_64_1204 ();
 sg13g2_decap_8 FILLER_64_1211 ();
 sg13g2_decap_8 FILLER_64_1218 ();
 sg13g2_decap_8 FILLER_64_1225 ();
 sg13g2_decap_8 FILLER_64_1232 ();
 sg13g2_decap_8 FILLER_64_1239 ();
 sg13g2_decap_8 FILLER_64_1246 ();
 sg13g2_decap_8 FILLER_64_1253 ();
 sg13g2_decap_8 FILLER_64_1260 ();
 sg13g2_decap_8 FILLER_64_1267 ();
 sg13g2_decap_8 FILLER_64_1274 ();
 sg13g2_decap_8 FILLER_64_1281 ();
 sg13g2_decap_8 FILLER_64_1288 ();
 sg13g2_decap_8 FILLER_64_1295 ();
 sg13g2_decap_8 FILLER_64_1302 ();
 sg13g2_decap_8 FILLER_64_1309 ();
 sg13g2_decap_8 FILLER_64_1316 ();
 sg13g2_decap_8 FILLER_64_1323 ();
 sg13g2_decap_8 FILLER_64_1330 ();
 sg13g2_decap_8 FILLER_64_1337 ();
 sg13g2_decap_8 FILLER_64_1344 ();
 sg13g2_decap_8 FILLER_64_1351 ();
 sg13g2_decap_8 FILLER_64_1358 ();
 sg13g2_decap_8 FILLER_64_1365 ();
 sg13g2_decap_8 FILLER_64_1372 ();
 sg13g2_decap_8 FILLER_64_1379 ();
 sg13g2_decap_8 FILLER_64_1386 ();
 sg13g2_decap_8 FILLER_64_1393 ();
 sg13g2_decap_8 FILLER_64_1400 ();
 sg13g2_decap_8 FILLER_64_1407 ();
 sg13g2_decap_8 FILLER_64_1414 ();
 sg13g2_decap_8 FILLER_64_1421 ();
 sg13g2_decap_8 FILLER_64_1428 ();
 sg13g2_decap_8 FILLER_64_1435 ();
 sg13g2_decap_8 FILLER_64_1442 ();
 sg13g2_decap_8 FILLER_64_1449 ();
 sg13g2_decap_8 FILLER_64_1456 ();
 sg13g2_decap_8 FILLER_64_1463 ();
 sg13g2_decap_8 FILLER_64_1470 ();
 sg13g2_decap_8 FILLER_64_1477 ();
 sg13g2_decap_8 FILLER_64_1484 ();
 sg13g2_decap_8 FILLER_64_1491 ();
 sg13g2_decap_8 FILLER_64_1498 ();
 sg13g2_decap_8 FILLER_64_1505 ();
 sg13g2_decap_8 FILLER_64_1512 ();
 sg13g2_decap_8 FILLER_64_1519 ();
 sg13g2_decap_8 FILLER_64_1526 ();
 sg13g2_decap_8 FILLER_64_1533 ();
 sg13g2_decap_8 FILLER_64_1540 ();
 sg13g2_decap_8 FILLER_64_1547 ();
 sg13g2_decap_8 FILLER_64_1554 ();
 sg13g2_decap_8 FILLER_64_1561 ();
 sg13g2_decap_8 FILLER_64_1568 ();
 sg13g2_decap_8 FILLER_64_1575 ();
 sg13g2_decap_8 FILLER_64_1582 ();
 sg13g2_decap_8 FILLER_64_1589 ();
 sg13g2_decap_8 FILLER_64_1596 ();
 sg13g2_decap_8 FILLER_64_1603 ();
 sg13g2_decap_8 FILLER_64_1610 ();
 sg13g2_decap_8 FILLER_64_1617 ();
 sg13g2_decap_8 FILLER_64_1624 ();
 sg13g2_decap_8 FILLER_64_1631 ();
 sg13g2_decap_8 FILLER_64_1638 ();
 sg13g2_decap_8 FILLER_64_1645 ();
 sg13g2_decap_8 FILLER_64_1652 ();
 sg13g2_decap_8 FILLER_64_1659 ();
 sg13g2_decap_8 FILLER_64_1666 ();
 sg13g2_decap_8 FILLER_64_1673 ();
 sg13g2_decap_8 FILLER_64_1680 ();
 sg13g2_decap_8 FILLER_64_1687 ();
 sg13g2_decap_8 FILLER_64_1694 ();
 sg13g2_decap_8 FILLER_64_1701 ();
 sg13g2_decap_8 FILLER_64_1708 ();
 sg13g2_decap_8 FILLER_64_1715 ();
 sg13g2_decap_8 FILLER_64_1722 ();
 sg13g2_decap_8 FILLER_64_1729 ();
 sg13g2_decap_8 FILLER_64_1736 ();
 sg13g2_decap_8 FILLER_64_1743 ();
 sg13g2_decap_8 FILLER_64_1750 ();
 sg13g2_decap_8 FILLER_64_1757 ();
 sg13g2_decap_8 FILLER_64_1764 ();
 sg13g2_decap_8 FILLER_64_1771 ();
 sg13g2_decap_8 FILLER_64_1778 ();
 sg13g2_decap_8 FILLER_64_1785 ();
 sg13g2_decap_8 FILLER_64_1792 ();
 sg13g2_decap_8 FILLER_64_1799 ();
 sg13g2_decap_8 FILLER_64_1806 ();
 sg13g2_decap_8 FILLER_64_1813 ();
 sg13g2_decap_8 FILLER_64_1820 ();
 sg13g2_decap_8 FILLER_64_1827 ();
 sg13g2_decap_8 FILLER_64_1834 ();
 sg13g2_decap_8 FILLER_64_1841 ();
 sg13g2_decap_8 FILLER_64_1848 ();
 sg13g2_decap_8 FILLER_64_1855 ();
 sg13g2_decap_8 FILLER_64_1862 ();
 sg13g2_decap_8 FILLER_64_1869 ();
 sg13g2_decap_8 FILLER_64_1876 ();
 sg13g2_decap_8 FILLER_64_1883 ();
 sg13g2_decap_8 FILLER_64_1890 ();
 sg13g2_decap_8 FILLER_64_1897 ();
 sg13g2_decap_8 FILLER_64_1904 ();
 sg13g2_decap_8 FILLER_64_1911 ();
 sg13g2_decap_8 FILLER_64_1918 ();
 sg13g2_decap_8 FILLER_64_1925 ();
 sg13g2_decap_8 FILLER_64_1932 ();
 sg13g2_decap_8 FILLER_64_1939 ();
 sg13g2_decap_8 FILLER_64_1946 ();
 sg13g2_decap_8 FILLER_64_1953 ();
 sg13g2_decap_8 FILLER_64_1960 ();
 sg13g2_decap_8 FILLER_64_1967 ();
 sg13g2_decap_8 FILLER_64_1974 ();
 sg13g2_decap_8 FILLER_64_1981 ();
 sg13g2_decap_8 FILLER_64_1988 ();
 sg13g2_decap_8 FILLER_64_1995 ();
 sg13g2_decap_8 FILLER_64_2002 ();
 sg13g2_decap_8 FILLER_64_2009 ();
 sg13g2_decap_8 FILLER_64_2016 ();
 sg13g2_decap_8 FILLER_64_2023 ();
 sg13g2_decap_8 FILLER_64_2030 ();
 sg13g2_decap_8 FILLER_64_2037 ();
 sg13g2_decap_8 FILLER_64_2044 ();
 sg13g2_decap_8 FILLER_64_2051 ();
 sg13g2_decap_8 FILLER_64_2058 ();
 sg13g2_decap_8 FILLER_64_2065 ();
 sg13g2_decap_8 FILLER_64_2072 ();
 sg13g2_decap_8 FILLER_64_2079 ();
 sg13g2_decap_8 FILLER_64_2086 ();
 sg13g2_decap_8 FILLER_64_2093 ();
 sg13g2_decap_8 FILLER_64_2100 ();
 sg13g2_decap_8 FILLER_64_2107 ();
 sg13g2_decap_8 FILLER_64_2114 ();
 sg13g2_decap_8 FILLER_64_2121 ();
 sg13g2_decap_8 FILLER_64_2128 ();
 sg13g2_decap_8 FILLER_64_2135 ();
 sg13g2_decap_8 FILLER_64_2142 ();
 sg13g2_decap_8 FILLER_64_2149 ();
 sg13g2_decap_8 FILLER_64_2156 ();
 sg13g2_decap_8 FILLER_64_2163 ();
 sg13g2_decap_8 FILLER_64_2170 ();
 sg13g2_decap_8 FILLER_64_2177 ();
 sg13g2_decap_8 FILLER_64_2184 ();
 sg13g2_decap_8 FILLER_64_2191 ();
 sg13g2_decap_8 FILLER_64_2198 ();
 sg13g2_decap_8 FILLER_64_2205 ();
 sg13g2_decap_8 FILLER_64_2212 ();
 sg13g2_decap_8 FILLER_64_2219 ();
 sg13g2_decap_8 FILLER_64_2226 ();
 sg13g2_decap_8 FILLER_64_2233 ();
 sg13g2_decap_8 FILLER_64_2240 ();
 sg13g2_decap_8 FILLER_64_2247 ();
 sg13g2_decap_8 FILLER_64_2254 ();
 sg13g2_decap_8 FILLER_64_2261 ();
 sg13g2_decap_8 FILLER_64_2268 ();
 sg13g2_decap_8 FILLER_64_2275 ();
 sg13g2_decap_8 FILLER_64_2282 ();
 sg13g2_decap_8 FILLER_64_2289 ();
 sg13g2_decap_8 FILLER_64_2296 ();
 sg13g2_decap_8 FILLER_64_2303 ();
 sg13g2_decap_8 FILLER_64_2310 ();
 sg13g2_decap_8 FILLER_64_2317 ();
 sg13g2_decap_8 FILLER_64_2324 ();
 sg13g2_decap_8 FILLER_64_2331 ();
 sg13g2_decap_8 FILLER_64_2338 ();
 sg13g2_decap_8 FILLER_64_2345 ();
 sg13g2_decap_8 FILLER_64_2352 ();
 sg13g2_decap_8 FILLER_64_2359 ();
 sg13g2_decap_8 FILLER_64_2366 ();
 sg13g2_decap_8 FILLER_64_2373 ();
 sg13g2_decap_8 FILLER_64_2380 ();
 sg13g2_decap_8 FILLER_64_2387 ();
 sg13g2_decap_8 FILLER_64_2394 ();
 sg13g2_decap_8 FILLER_64_2401 ();
 sg13g2_decap_8 FILLER_64_2408 ();
 sg13g2_decap_8 FILLER_64_2415 ();
 sg13g2_decap_8 FILLER_64_2422 ();
 sg13g2_decap_8 FILLER_64_2429 ();
 sg13g2_decap_8 FILLER_64_2436 ();
 sg13g2_decap_8 FILLER_64_2443 ();
 sg13g2_decap_8 FILLER_64_2450 ();
 sg13g2_decap_8 FILLER_64_2457 ();
 sg13g2_decap_8 FILLER_64_2464 ();
 sg13g2_decap_8 FILLER_64_2471 ();
 sg13g2_decap_8 FILLER_64_2478 ();
 sg13g2_decap_8 FILLER_64_2485 ();
 sg13g2_decap_8 FILLER_64_2492 ();
 sg13g2_decap_8 FILLER_64_2499 ();
 sg13g2_decap_8 FILLER_64_2506 ();
 sg13g2_decap_8 FILLER_64_2513 ();
 sg13g2_decap_8 FILLER_64_2520 ();
 sg13g2_decap_8 FILLER_64_2527 ();
 sg13g2_decap_8 FILLER_64_2534 ();
 sg13g2_decap_8 FILLER_64_2541 ();
 sg13g2_decap_8 FILLER_64_2548 ();
 sg13g2_decap_8 FILLER_64_2555 ();
 sg13g2_decap_8 FILLER_64_2562 ();
 sg13g2_decap_8 FILLER_64_2569 ();
 sg13g2_decap_8 FILLER_64_2576 ();
 sg13g2_decap_8 FILLER_64_2583 ();
 sg13g2_decap_8 FILLER_64_2590 ();
 sg13g2_decap_8 FILLER_64_2597 ();
 sg13g2_decap_8 FILLER_64_2604 ();
 sg13g2_decap_8 FILLER_64_2611 ();
 sg13g2_decap_8 FILLER_64_2618 ();
 sg13g2_decap_8 FILLER_64_2625 ();
 sg13g2_decap_8 FILLER_64_2632 ();
 sg13g2_decap_8 FILLER_64_2639 ();
 sg13g2_decap_8 FILLER_64_2646 ();
 sg13g2_decap_8 FILLER_64_2653 ();
 sg13g2_decap_8 FILLER_64_2660 ();
 sg13g2_decap_8 FILLER_64_2667 ();
 sg13g2_decap_8 FILLER_64_2674 ();
 sg13g2_decap_8 FILLER_64_2681 ();
 sg13g2_decap_8 FILLER_64_2688 ();
 sg13g2_decap_8 FILLER_64_2695 ();
 sg13g2_decap_8 FILLER_64_2702 ();
 sg13g2_decap_8 FILLER_64_2709 ();
 sg13g2_decap_8 FILLER_64_2716 ();
 sg13g2_decap_8 FILLER_64_2723 ();
 sg13g2_decap_8 FILLER_64_2730 ();
 sg13g2_decap_8 FILLER_64_2737 ();
 sg13g2_decap_8 FILLER_64_2744 ();
 sg13g2_decap_8 FILLER_64_2751 ();
 sg13g2_decap_8 FILLER_64_2758 ();
 sg13g2_decap_8 FILLER_64_2765 ();
 sg13g2_decap_8 FILLER_64_2772 ();
 sg13g2_decap_8 FILLER_64_2779 ();
 sg13g2_decap_8 FILLER_64_2786 ();
 sg13g2_decap_8 FILLER_64_2793 ();
 sg13g2_decap_8 FILLER_64_2800 ();
 sg13g2_decap_8 FILLER_64_2807 ();
 sg13g2_decap_8 FILLER_64_2814 ();
 sg13g2_decap_8 FILLER_64_2821 ();
 sg13g2_decap_8 FILLER_64_2828 ();
 sg13g2_decap_8 FILLER_64_2835 ();
 sg13g2_decap_8 FILLER_64_2842 ();
 sg13g2_decap_8 FILLER_64_2849 ();
 sg13g2_decap_8 FILLER_64_2856 ();
 sg13g2_decap_8 FILLER_64_2863 ();
 sg13g2_decap_8 FILLER_64_2870 ();
 sg13g2_decap_8 FILLER_64_2877 ();
 sg13g2_decap_8 FILLER_64_2884 ();
 sg13g2_decap_8 FILLER_64_2891 ();
 sg13g2_decap_8 FILLER_64_2898 ();
 sg13g2_decap_8 FILLER_64_2905 ();
 sg13g2_decap_8 FILLER_64_2912 ();
 sg13g2_decap_8 FILLER_64_2919 ();
 sg13g2_decap_8 FILLER_64_2926 ();
 sg13g2_decap_8 FILLER_64_2933 ();
 sg13g2_decap_8 FILLER_64_2940 ();
 sg13g2_decap_8 FILLER_64_2947 ();
 sg13g2_decap_8 FILLER_64_2954 ();
 sg13g2_decap_8 FILLER_64_2961 ();
 sg13g2_decap_8 FILLER_64_2968 ();
 sg13g2_decap_8 FILLER_64_2975 ();
 sg13g2_decap_8 FILLER_64_2982 ();
 sg13g2_decap_8 FILLER_64_2989 ();
 sg13g2_decap_8 FILLER_64_2996 ();
 sg13g2_decap_8 FILLER_64_3003 ();
 sg13g2_decap_8 FILLER_64_3010 ();
 sg13g2_decap_8 FILLER_64_3017 ();
 sg13g2_decap_8 FILLER_64_3024 ();
 sg13g2_decap_8 FILLER_64_3031 ();
 sg13g2_decap_8 FILLER_64_3038 ();
 sg13g2_decap_8 FILLER_64_3045 ();
 sg13g2_decap_8 FILLER_64_3052 ();
 sg13g2_decap_8 FILLER_64_3059 ();
 sg13g2_decap_8 FILLER_64_3066 ();
 sg13g2_decap_8 FILLER_64_3073 ();
 sg13g2_decap_8 FILLER_64_3080 ();
 sg13g2_decap_8 FILLER_64_3087 ();
 sg13g2_decap_8 FILLER_64_3094 ();
 sg13g2_decap_8 FILLER_64_3101 ();
 sg13g2_decap_8 FILLER_64_3108 ();
 sg13g2_decap_8 FILLER_64_3115 ();
 sg13g2_decap_8 FILLER_64_3122 ();
 sg13g2_decap_8 FILLER_64_3129 ();
 sg13g2_decap_8 FILLER_64_3136 ();
 sg13g2_decap_8 FILLER_64_3143 ();
 sg13g2_decap_8 FILLER_64_3150 ();
 sg13g2_decap_8 FILLER_64_3157 ();
 sg13g2_decap_8 FILLER_64_3164 ();
 sg13g2_decap_8 FILLER_64_3171 ();
 sg13g2_decap_8 FILLER_64_3178 ();
 sg13g2_decap_8 FILLER_64_3185 ();
 sg13g2_decap_8 FILLER_64_3192 ();
 sg13g2_decap_8 FILLER_64_3199 ();
 sg13g2_decap_8 FILLER_64_3206 ();
 sg13g2_decap_8 FILLER_64_3213 ();
 sg13g2_decap_8 FILLER_64_3220 ();
 sg13g2_decap_8 FILLER_64_3227 ();
 sg13g2_decap_8 FILLER_64_3234 ();
 sg13g2_decap_8 FILLER_64_3241 ();
 sg13g2_decap_8 FILLER_64_3248 ();
 sg13g2_decap_8 FILLER_64_3255 ();
 sg13g2_decap_8 FILLER_64_3262 ();
 sg13g2_decap_8 FILLER_64_3269 ();
 sg13g2_decap_8 FILLER_64_3276 ();
 sg13g2_decap_8 FILLER_64_3283 ();
 sg13g2_decap_8 FILLER_64_3290 ();
 sg13g2_decap_8 FILLER_64_3297 ();
 sg13g2_decap_8 FILLER_64_3304 ();
 sg13g2_decap_8 FILLER_64_3311 ();
 sg13g2_decap_8 FILLER_64_3318 ();
 sg13g2_decap_8 FILLER_64_3325 ();
 sg13g2_decap_8 FILLER_64_3332 ();
 sg13g2_decap_8 FILLER_64_3339 ();
 sg13g2_decap_8 FILLER_64_3346 ();
 sg13g2_decap_8 FILLER_64_3353 ();
 sg13g2_decap_8 FILLER_64_3360 ();
 sg13g2_decap_8 FILLER_64_3367 ();
 sg13g2_decap_8 FILLER_64_3374 ();
 sg13g2_decap_8 FILLER_64_3381 ();
 sg13g2_decap_8 FILLER_64_3388 ();
 sg13g2_decap_8 FILLER_64_3395 ();
 sg13g2_decap_8 FILLER_64_3402 ();
 sg13g2_decap_8 FILLER_64_3409 ();
 sg13g2_decap_8 FILLER_64_3416 ();
 sg13g2_decap_8 FILLER_64_3423 ();
 sg13g2_decap_8 FILLER_64_3430 ();
 sg13g2_decap_8 FILLER_64_3437 ();
 sg13g2_decap_8 FILLER_64_3444 ();
 sg13g2_decap_8 FILLER_64_3451 ();
 sg13g2_decap_8 FILLER_64_3458 ();
 sg13g2_decap_8 FILLER_64_3465 ();
 sg13g2_decap_8 FILLER_64_3472 ();
 sg13g2_decap_8 FILLER_64_3479 ();
 sg13g2_decap_8 FILLER_64_3486 ();
 sg13g2_decap_8 FILLER_64_3493 ();
 sg13g2_decap_8 FILLER_64_3500 ();
 sg13g2_decap_8 FILLER_64_3507 ();
 sg13g2_decap_8 FILLER_64_3514 ();
 sg13g2_decap_8 FILLER_64_3521 ();
 sg13g2_decap_8 FILLER_64_3528 ();
 sg13g2_decap_8 FILLER_64_3535 ();
 sg13g2_decap_8 FILLER_64_3542 ();
 sg13g2_decap_8 FILLER_64_3549 ();
 sg13g2_decap_8 FILLER_64_3556 ();
 sg13g2_decap_8 FILLER_64_3563 ();
 sg13g2_decap_8 FILLER_64_3570 ();
 sg13g2_fill_2 FILLER_64_3577 ();
 sg13g2_fill_1 FILLER_64_3579 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_decap_8 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_decap_8 FILLER_65_119 ();
 sg13g2_decap_8 FILLER_65_126 ();
 sg13g2_decap_8 FILLER_65_133 ();
 sg13g2_decap_8 FILLER_65_140 ();
 sg13g2_decap_8 FILLER_65_147 ();
 sg13g2_decap_8 FILLER_65_154 ();
 sg13g2_decap_8 FILLER_65_161 ();
 sg13g2_decap_8 FILLER_65_168 ();
 sg13g2_decap_8 FILLER_65_175 ();
 sg13g2_decap_8 FILLER_65_182 ();
 sg13g2_decap_8 FILLER_65_189 ();
 sg13g2_decap_8 FILLER_65_196 ();
 sg13g2_decap_8 FILLER_65_203 ();
 sg13g2_decap_8 FILLER_65_210 ();
 sg13g2_decap_8 FILLER_65_217 ();
 sg13g2_decap_8 FILLER_65_224 ();
 sg13g2_decap_8 FILLER_65_231 ();
 sg13g2_decap_8 FILLER_65_238 ();
 sg13g2_decap_8 FILLER_65_245 ();
 sg13g2_decap_8 FILLER_65_252 ();
 sg13g2_decap_8 FILLER_65_259 ();
 sg13g2_decap_8 FILLER_65_266 ();
 sg13g2_decap_8 FILLER_65_273 ();
 sg13g2_decap_8 FILLER_65_280 ();
 sg13g2_decap_8 FILLER_65_287 ();
 sg13g2_decap_8 FILLER_65_294 ();
 sg13g2_decap_8 FILLER_65_301 ();
 sg13g2_decap_8 FILLER_65_308 ();
 sg13g2_decap_8 FILLER_65_315 ();
 sg13g2_decap_8 FILLER_65_322 ();
 sg13g2_decap_8 FILLER_65_329 ();
 sg13g2_decap_8 FILLER_65_336 ();
 sg13g2_decap_8 FILLER_65_343 ();
 sg13g2_decap_8 FILLER_65_350 ();
 sg13g2_decap_8 FILLER_65_357 ();
 sg13g2_decap_8 FILLER_65_364 ();
 sg13g2_decap_8 FILLER_65_371 ();
 sg13g2_decap_8 FILLER_65_378 ();
 sg13g2_decap_8 FILLER_65_385 ();
 sg13g2_decap_8 FILLER_65_392 ();
 sg13g2_decap_8 FILLER_65_399 ();
 sg13g2_decap_8 FILLER_65_406 ();
 sg13g2_decap_8 FILLER_65_413 ();
 sg13g2_decap_8 FILLER_65_420 ();
 sg13g2_decap_8 FILLER_65_427 ();
 sg13g2_decap_8 FILLER_65_434 ();
 sg13g2_decap_8 FILLER_65_441 ();
 sg13g2_decap_8 FILLER_65_448 ();
 sg13g2_decap_8 FILLER_65_455 ();
 sg13g2_decap_8 FILLER_65_462 ();
 sg13g2_decap_8 FILLER_65_469 ();
 sg13g2_decap_8 FILLER_65_476 ();
 sg13g2_decap_8 FILLER_65_483 ();
 sg13g2_decap_8 FILLER_65_490 ();
 sg13g2_decap_8 FILLER_65_497 ();
 sg13g2_decap_8 FILLER_65_504 ();
 sg13g2_decap_8 FILLER_65_511 ();
 sg13g2_decap_8 FILLER_65_518 ();
 sg13g2_decap_8 FILLER_65_525 ();
 sg13g2_decap_8 FILLER_65_532 ();
 sg13g2_decap_8 FILLER_65_539 ();
 sg13g2_decap_8 FILLER_65_546 ();
 sg13g2_decap_8 FILLER_65_553 ();
 sg13g2_decap_8 FILLER_65_560 ();
 sg13g2_decap_8 FILLER_65_567 ();
 sg13g2_decap_8 FILLER_65_574 ();
 sg13g2_decap_8 FILLER_65_581 ();
 sg13g2_decap_8 FILLER_65_588 ();
 sg13g2_decap_8 FILLER_65_595 ();
 sg13g2_decap_8 FILLER_65_602 ();
 sg13g2_decap_8 FILLER_65_609 ();
 sg13g2_decap_8 FILLER_65_616 ();
 sg13g2_decap_8 FILLER_65_623 ();
 sg13g2_decap_8 FILLER_65_630 ();
 sg13g2_decap_8 FILLER_65_637 ();
 sg13g2_decap_8 FILLER_65_644 ();
 sg13g2_decap_8 FILLER_65_651 ();
 sg13g2_decap_8 FILLER_65_658 ();
 sg13g2_decap_8 FILLER_65_665 ();
 sg13g2_decap_8 FILLER_65_672 ();
 sg13g2_decap_8 FILLER_65_679 ();
 sg13g2_decap_8 FILLER_65_686 ();
 sg13g2_decap_8 FILLER_65_693 ();
 sg13g2_decap_8 FILLER_65_700 ();
 sg13g2_decap_8 FILLER_65_707 ();
 sg13g2_decap_8 FILLER_65_714 ();
 sg13g2_decap_8 FILLER_65_721 ();
 sg13g2_decap_8 FILLER_65_728 ();
 sg13g2_decap_8 FILLER_65_735 ();
 sg13g2_decap_8 FILLER_65_742 ();
 sg13g2_decap_8 FILLER_65_749 ();
 sg13g2_decap_8 FILLER_65_756 ();
 sg13g2_decap_8 FILLER_65_763 ();
 sg13g2_decap_8 FILLER_65_770 ();
 sg13g2_decap_8 FILLER_65_777 ();
 sg13g2_decap_8 FILLER_65_784 ();
 sg13g2_decap_8 FILLER_65_791 ();
 sg13g2_decap_8 FILLER_65_798 ();
 sg13g2_decap_8 FILLER_65_805 ();
 sg13g2_decap_8 FILLER_65_812 ();
 sg13g2_decap_8 FILLER_65_819 ();
 sg13g2_decap_8 FILLER_65_826 ();
 sg13g2_decap_8 FILLER_65_833 ();
 sg13g2_decap_8 FILLER_65_840 ();
 sg13g2_decap_8 FILLER_65_847 ();
 sg13g2_decap_8 FILLER_65_854 ();
 sg13g2_decap_8 FILLER_65_861 ();
 sg13g2_decap_8 FILLER_65_868 ();
 sg13g2_decap_8 FILLER_65_875 ();
 sg13g2_decap_8 FILLER_65_882 ();
 sg13g2_decap_8 FILLER_65_889 ();
 sg13g2_decap_8 FILLER_65_896 ();
 sg13g2_decap_8 FILLER_65_903 ();
 sg13g2_decap_8 FILLER_65_910 ();
 sg13g2_decap_8 FILLER_65_917 ();
 sg13g2_decap_8 FILLER_65_924 ();
 sg13g2_decap_8 FILLER_65_931 ();
 sg13g2_decap_8 FILLER_65_938 ();
 sg13g2_decap_8 FILLER_65_945 ();
 sg13g2_decap_8 FILLER_65_952 ();
 sg13g2_decap_8 FILLER_65_959 ();
 sg13g2_decap_8 FILLER_65_966 ();
 sg13g2_decap_8 FILLER_65_973 ();
 sg13g2_decap_8 FILLER_65_980 ();
 sg13g2_decap_8 FILLER_65_987 ();
 sg13g2_decap_8 FILLER_65_994 ();
 sg13g2_decap_8 FILLER_65_1001 ();
 sg13g2_decap_8 FILLER_65_1008 ();
 sg13g2_decap_8 FILLER_65_1015 ();
 sg13g2_decap_8 FILLER_65_1022 ();
 sg13g2_decap_8 FILLER_65_1029 ();
 sg13g2_decap_8 FILLER_65_1036 ();
 sg13g2_decap_8 FILLER_65_1043 ();
 sg13g2_decap_8 FILLER_65_1050 ();
 sg13g2_decap_8 FILLER_65_1057 ();
 sg13g2_decap_8 FILLER_65_1064 ();
 sg13g2_decap_8 FILLER_65_1071 ();
 sg13g2_decap_8 FILLER_65_1078 ();
 sg13g2_decap_8 FILLER_65_1085 ();
 sg13g2_decap_8 FILLER_65_1092 ();
 sg13g2_decap_8 FILLER_65_1099 ();
 sg13g2_decap_8 FILLER_65_1106 ();
 sg13g2_decap_8 FILLER_65_1113 ();
 sg13g2_decap_8 FILLER_65_1120 ();
 sg13g2_decap_8 FILLER_65_1127 ();
 sg13g2_decap_8 FILLER_65_1134 ();
 sg13g2_decap_8 FILLER_65_1141 ();
 sg13g2_decap_8 FILLER_65_1148 ();
 sg13g2_decap_8 FILLER_65_1155 ();
 sg13g2_decap_8 FILLER_65_1162 ();
 sg13g2_decap_8 FILLER_65_1169 ();
 sg13g2_decap_8 FILLER_65_1176 ();
 sg13g2_decap_8 FILLER_65_1183 ();
 sg13g2_decap_8 FILLER_65_1190 ();
 sg13g2_decap_8 FILLER_65_1197 ();
 sg13g2_decap_8 FILLER_65_1204 ();
 sg13g2_decap_8 FILLER_65_1211 ();
 sg13g2_decap_8 FILLER_65_1218 ();
 sg13g2_decap_8 FILLER_65_1225 ();
 sg13g2_decap_8 FILLER_65_1232 ();
 sg13g2_decap_8 FILLER_65_1239 ();
 sg13g2_decap_8 FILLER_65_1246 ();
 sg13g2_decap_8 FILLER_65_1253 ();
 sg13g2_decap_8 FILLER_65_1260 ();
 sg13g2_decap_8 FILLER_65_1267 ();
 sg13g2_decap_8 FILLER_65_1274 ();
 sg13g2_decap_8 FILLER_65_1281 ();
 sg13g2_decap_8 FILLER_65_1288 ();
 sg13g2_decap_8 FILLER_65_1295 ();
 sg13g2_decap_8 FILLER_65_1302 ();
 sg13g2_decap_8 FILLER_65_1309 ();
 sg13g2_decap_8 FILLER_65_1316 ();
 sg13g2_decap_8 FILLER_65_1323 ();
 sg13g2_decap_8 FILLER_65_1330 ();
 sg13g2_decap_8 FILLER_65_1337 ();
 sg13g2_decap_8 FILLER_65_1344 ();
 sg13g2_decap_8 FILLER_65_1351 ();
 sg13g2_decap_8 FILLER_65_1358 ();
 sg13g2_decap_8 FILLER_65_1365 ();
 sg13g2_decap_8 FILLER_65_1372 ();
 sg13g2_decap_8 FILLER_65_1379 ();
 sg13g2_decap_8 FILLER_65_1386 ();
 sg13g2_decap_8 FILLER_65_1393 ();
 sg13g2_decap_8 FILLER_65_1400 ();
 sg13g2_decap_8 FILLER_65_1407 ();
 sg13g2_decap_8 FILLER_65_1414 ();
 sg13g2_decap_8 FILLER_65_1421 ();
 sg13g2_decap_8 FILLER_65_1428 ();
 sg13g2_decap_8 FILLER_65_1435 ();
 sg13g2_decap_8 FILLER_65_1442 ();
 sg13g2_decap_8 FILLER_65_1449 ();
 sg13g2_decap_8 FILLER_65_1456 ();
 sg13g2_decap_8 FILLER_65_1463 ();
 sg13g2_decap_8 FILLER_65_1470 ();
 sg13g2_decap_8 FILLER_65_1477 ();
 sg13g2_decap_8 FILLER_65_1484 ();
 sg13g2_decap_8 FILLER_65_1491 ();
 sg13g2_decap_8 FILLER_65_1498 ();
 sg13g2_decap_8 FILLER_65_1505 ();
 sg13g2_decap_8 FILLER_65_1512 ();
 sg13g2_decap_8 FILLER_65_1519 ();
 sg13g2_decap_8 FILLER_65_1526 ();
 sg13g2_decap_8 FILLER_65_1533 ();
 sg13g2_decap_8 FILLER_65_1540 ();
 sg13g2_decap_8 FILLER_65_1547 ();
 sg13g2_decap_8 FILLER_65_1554 ();
 sg13g2_decap_8 FILLER_65_1561 ();
 sg13g2_decap_8 FILLER_65_1568 ();
 sg13g2_decap_8 FILLER_65_1575 ();
 sg13g2_decap_8 FILLER_65_1582 ();
 sg13g2_decap_8 FILLER_65_1589 ();
 sg13g2_decap_8 FILLER_65_1596 ();
 sg13g2_decap_8 FILLER_65_1603 ();
 sg13g2_decap_8 FILLER_65_1610 ();
 sg13g2_decap_8 FILLER_65_1617 ();
 sg13g2_decap_8 FILLER_65_1624 ();
 sg13g2_decap_8 FILLER_65_1631 ();
 sg13g2_decap_8 FILLER_65_1638 ();
 sg13g2_decap_8 FILLER_65_1645 ();
 sg13g2_decap_8 FILLER_65_1652 ();
 sg13g2_decap_8 FILLER_65_1659 ();
 sg13g2_decap_8 FILLER_65_1666 ();
 sg13g2_decap_8 FILLER_65_1673 ();
 sg13g2_decap_8 FILLER_65_1680 ();
 sg13g2_decap_8 FILLER_65_1687 ();
 sg13g2_decap_8 FILLER_65_1694 ();
 sg13g2_decap_8 FILLER_65_1701 ();
 sg13g2_decap_8 FILLER_65_1708 ();
 sg13g2_decap_8 FILLER_65_1715 ();
 sg13g2_decap_8 FILLER_65_1722 ();
 sg13g2_decap_8 FILLER_65_1729 ();
 sg13g2_decap_8 FILLER_65_1736 ();
 sg13g2_decap_8 FILLER_65_1743 ();
 sg13g2_decap_8 FILLER_65_1750 ();
 sg13g2_decap_8 FILLER_65_1757 ();
 sg13g2_decap_8 FILLER_65_1764 ();
 sg13g2_decap_8 FILLER_65_1771 ();
 sg13g2_decap_8 FILLER_65_1778 ();
 sg13g2_decap_8 FILLER_65_1785 ();
 sg13g2_decap_8 FILLER_65_1792 ();
 sg13g2_decap_8 FILLER_65_1799 ();
 sg13g2_decap_8 FILLER_65_1806 ();
 sg13g2_decap_8 FILLER_65_1813 ();
 sg13g2_decap_8 FILLER_65_1820 ();
 sg13g2_decap_8 FILLER_65_1827 ();
 sg13g2_decap_8 FILLER_65_1834 ();
 sg13g2_decap_8 FILLER_65_1841 ();
 sg13g2_decap_8 FILLER_65_1848 ();
 sg13g2_decap_8 FILLER_65_1855 ();
 sg13g2_decap_8 FILLER_65_1862 ();
 sg13g2_decap_8 FILLER_65_1869 ();
 sg13g2_decap_8 FILLER_65_1876 ();
 sg13g2_decap_8 FILLER_65_1883 ();
 sg13g2_decap_8 FILLER_65_1890 ();
 sg13g2_decap_8 FILLER_65_1897 ();
 sg13g2_decap_8 FILLER_65_1904 ();
 sg13g2_decap_8 FILLER_65_1911 ();
 sg13g2_decap_8 FILLER_65_1918 ();
 sg13g2_decap_8 FILLER_65_1925 ();
 sg13g2_decap_8 FILLER_65_1932 ();
 sg13g2_decap_8 FILLER_65_1939 ();
 sg13g2_decap_8 FILLER_65_1946 ();
 sg13g2_decap_8 FILLER_65_1953 ();
 sg13g2_decap_8 FILLER_65_1960 ();
 sg13g2_decap_8 FILLER_65_1967 ();
 sg13g2_decap_8 FILLER_65_1974 ();
 sg13g2_decap_8 FILLER_65_1981 ();
 sg13g2_decap_8 FILLER_65_1988 ();
 sg13g2_decap_8 FILLER_65_1995 ();
 sg13g2_decap_8 FILLER_65_2002 ();
 sg13g2_decap_8 FILLER_65_2009 ();
 sg13g2_decap_8 FILLER_65_2016 ();
 sg13g2_decap_8 FILLER_65_2023 ();
 sg13g2_decap_8 FILLER_65_2030 ();
 sg13g2_decap_8 FILLER_65_2037 ();
 sg13g2_decap_8 FILLER_65_2044 ();
 sg13g2_decap_8 FILLER_65_2051 ();
 sg13g2_decap_8 FILLER_65_2058 ();
 sg13g2_decap_8 FILLER_65_2065 ();
 sg13g2_decap_8 FILLER_65_2072 ();
 sg13g2_decap_8 FILLER_65_2079 ();
 sg13g2_decap_8 FILLER_65_2086 ();
 sg13g2_decap_8 FILLER_65_2093 ();
 sg13g2_decap_8 FILLER_65_2100 ();
 sg13g2_decap_8 FILLER_65_2107 ();
 sg13g2_decap_8 FILLER_65_2114 ();
 sg13g2_decap_8 FILLER_65_2121 ();
 sg13g2_decap_8 FILLER_65_2128 ();
 sg13g2_decap_8 FILLER_65_2135 ();
 sg13g2_decap_8 FILLER_65_2142 ();
 sg13g2_decap_8 FILLER_65_2149 ();
 sg13g2_decap_8 FILLER_65_2156 ();
 sg13g2_decap_8 FILLER_65_2163 ();
 sg13g2_decap_8 FILLER_65_2170 ();
 sg13g2_decap_8 FILLER_65_2177 ();
 sg13g2_decap_8 FILLER_65_2184 ();
 sg13g2_decap_8 FILLER_65_2191 ();
 sg13g2_decap_8 FILLER_65_2198 ();
 sg13g2_decap_8 FILLER_65_2205 ();
 sg13g2_decap_8 FILLER_65_2212 ();
 sg13g2_decap_8 FILLER_65_2219 ();
 sg13g2_decap_8 FILLER_65_2226 ();
 sg13g2_decap_8 FILLER_65_2233 ();
 sg13g2_decap_8 FILLER_65_2240 ();
 sg13g2_decap_8 FILLER_65_2247 ();
 sg13g2_decap_8 FILLER_65_2254 ();
 sg13g2_decap_8 FILLER_65_2261 ();
 sg13g2_decap_8 FILLER_65_2268 ();
 sg13g2_decap_8 FILLER_65_2275 ();
 sg13g2_decap_8 FILLER_65_2282 ();
 sg13g2_decap_8 FILLER_65_2289 ();
 sg13g2_decap_8 FILLER_65_2296 ();
 sg13g2_decap_8 FILLER_65_2303 ();
 sg13g2_decap_8 FILLER_65_2310 ();
 sg13g2_decap_8 FILLER_65_2317 ();
 sg13g2_decap_8 FILLER_65_2324 ();
 sg13g2_decap_8 FILLER_65_2331 ();
 sg13g2_decap_8 FILLER_65_2338 ();
 sg13g2_decap_8 FILLER_65_2345 ();
 sg13g2_decap_8 FILLER_65_2352 ();
 sg13g2_decap_8 FILLER_65_2359 ();
 sg13g2_decap_8 FILLER_65_2366 ();
 sg13g2_decap_8 FILLER_65_2373 ();
 sg13g2_decap_8 FILLER_65_2380 ();
 sg13g2_decap_8 FILLER_65_2387 ();
 sg13g2_decap_8 FILLER_65_2394 ();
 sg13g2_decap_8 FILLER_65_2401 ();
 sg13g2_decap_8 FILLER_65_2408 ();
 sg13g2_decap_8 FILLER_65_2415 ();
 sg13g2_decap_8 FILLER_65_2422 ();
 sg13g2_decap_8 FILLER_65_2429 ();
 sg13g2_decap_8 FILLER_65_2436 ();
 sg13g2_decap_8 FILLER_65_2443 ();
 sg13g2_decap_8 FILLER_65_2450 ();
 sg13g2_decap_8 FILLER_65_2457 ();
 sg13g2_decap_8 FILLER_65_2464 ();
 sg13g2_decap_8 FILLER_65_2471 ();
 sg13g2_decap_8 FILLER_65_2478 ();
 sg13g2_decap_8 FILLER_65_2485 ();
 sg13g2_decap_8 FILLER_65_2492 ();
 sg13g2_decap_8 FILLER_65_2499 ();
 sg13g2_decap_8 FILLER_65_2506 ();
 sg13g2_decap_8 FILLER_65_2513 ();
 sg13g2_decap_8 FILLER_65_2520 ();
 sg13g2_decap_8 FILLER_65_2527 ();
 sg13g2_decap_8 FILLER_65_2534 ();
 sg13g2_decap_8 FILLER_65_2541 ();
 sg13g2_decap_8 FILLER_65_2548 ();
 sg13g2_decap_8 FILLER_65_2555 ();
 sg13g2_decap_8 FILLER_65_2562 ();
 sg13g2_decap_8 FILLER_65_2569 ();
 sg13g2_decap_8 FILLER_65_2576 ();
 sg13g2_decap_8 FILLER_65_2583 ();
 sg13g2_decap_8 FILLER_65_2590 ();
 sg13g2_decap_8 FILLER_65_2597 ();
 sg13g2_decap_8 FILLER_65_2604 ();
 sg13g2_decap_8 FILLER_65_2611 ();
 sg13g2_decap_8 FILLER_65_2618 ();
 sg13g2_decap_8 FILLER_65_2625 ();
 sg13g2_decap_8 FILLER_65_2632 ();
 sg13g2_decap_8 FILLER_65_2639 ();
 sg13g2_decap_8 FILLER_65_2646 ();
 sg13g2_decap_8 FILLER_65_2653 ();
 sg13g2_decap_8 FILLER_65_2660 ();
 sg13g2_decap_8 FILLER_65_2667 ();
 sg13g2_decap_8 FILLER_65_2674 ();
 sg13g2_decap_8 FILLER_65_2681 ();
 sg13g2_decap_8 FILLER_65_2688 ();
 sg13g2_decap_8 FILLER_65_2695 ();
 sg13g2_decap_8 FILLER_65_2702 ();
 sg13g2_decap_8 FILLER_65_2709 ();
 sg13g2_decap_8 FILLER_65_2716 ();
 sg13g2_decap_8 FILLER_65_2723 ();
 sg13g2_decap_8 FILLER_65_2730 ();
 sg13g2_decap_8 FILLER_65_2737 ();
 sg13g2_decap_8 FILLER_65_2744 ();
 sg13g2_decap_8 FILLER_65_2751 ();
 sg13g2_decap_8 FILLER_65_2758 ();
 sg13g2_decap_8 FILLER_65_2765 ();
 sg13g2_decap_8 FILLER_65_2772 ();
 sg13g2_decap_8 FILLER_65_2779 ();
 sg13g2_decap_8 FILLER_65_2786 ();
 sg13g2_decap_8 FILLER_65_2793 ();
 sg13g2_decap_8 FILLER_65_2800 ();
 sg13g2_decap_8 FILLER_65_2807 ();
 sg13g2_decap_8 FILLER_65_2814 ();
 sg13g2_decap_8 FILLER_65_2821 ();
 sg13g2_decap_8 FILLER_65_2828 ();
 sg13g2_decap_8 FILLER_65_2835 ();
 sg13g2_decap_8 FILLER_65_2842 ();
 sg13g2_decap_8 FILLER_65_2849 ();
 sg13g2_decap_8 FILLER_65_2856 ();
 sg13g2_decap_8 FILLER_65_2863 ();
 sg13g2_decap_8 FILLER_65_2870 ();
 sg13g2_decap_8 FILLER_65_2877 ();
 sg13g2_decap_8 FILLER_65_2884 ();
 sg13g2_decap_8 FILLER_65_2891 ();
 sg13g2_decap_8 FILLER_65_2898 ();
 sg13g2_decap_8 FILLER_65_2905 ();
 sg13g2_decap_8 FILLER_65_2912 ();
 sg13g2_decap_8 FILLER_65_2919 ();
 sg13g2_decap_8 FILLER_65_2926 ();
 sg13g2_decap_8 FILLER_65_2933 ();
 sg13g2_decap_8 FILLER_65_2940 ();
 sg13g2_decap_8 FILLER_65_2947 ();
 sg13g2_decap_8 FILLER_65_2954 ();
 sg13g2_decap_8 FILLER_65_2961 ();
 sg13g2_decap_8 FILLER_65_2968 ();
 sg13g2_decap_8 FILLER_65_2975 ();
 sg13g2_decap_8 FILLER_65_2982 ();
 sg13g2_decap_8 FILLER_65_2989 ();
 sg13g2_decap_8 FILLER_65_2996 ();
 sg13g2_decap_8 FILLER_65_3003 ();
 sg13g2_decap_8 FILLER_65_3010 ();
 sg13g2_decap_8 FILLER_65_3017 ();
 sg13g2_decap_8 FILLER_65_3024 ();
 sg13g2_decap_8 FILLER_65_3031 ();
 sg13g2_decap_8 FILLER_65_3038 ();
 sg13g2_decap_8 FILLER_65_3045 ();
 sg13g2_decap_8 FILLER_65_3052 ();
 sg13g2_decap_8 FILLER_65_3059 ();
 sg13g2_decap_8 FILLER_65_3066 ();
 sg13g2_decap_8 FILLER_65_3073 ();
 sg13g2_decap_8 FILLER_65_3080 ();
 sg13g2_decap_8 FILLER_65_3087 ();
 sg13g2_decap_8 FILLER_65_3094 ();
 sg13g2_decap_8 FILLER_65_3101 ();
 sg13g2_decap_8 FILLER_65_3108 ();
 sg13g2_decap_8 FILLER_65_3115 ();
 sg13g2_decap_8 FILLER_65_3122 ();
 sg13g2_decap_8 FILLER_65_3129 ();
 sg13g2_decap_8 FILLER_65_3136 ();
 sg13g2_decap_8 FILLER_65_3143 ();
 sg13g2_decap_8 FILLER_65_3150 ();
 sg13g2_decap_8 FILLER_65_3157 ();
 sg13g2_decap_8 FILLER_65_3164 ();
 sg13g2_decap_8 FILLER_65_3171 ();
 sg13g2_decap_8 FILLER_65_3178 ();
 sg13g2_decap_8 FILLER_65_3185 ();
 sg13g2_decap_8 FILLER_65_3192 ();
 sg13g2_decap_8 FILLER_65_3199 ();
 sg13g2_decap_8 FILLER_65_3206 ();
 sg13g2_decap_8 FILLER_65_3213 ();
 sg13g2_decap_8 FILLER_65_3220 ();
 sg13g2_decap_8 FILLER_65_3227 ();
 sg13g2_decap_8 FILLER_65_3234 ();
 sg13g2_decap_8 FILLER_65_3241 ();
 sg13g2_decap_8 FILLER_65_3248 ();
 sg13g2_decap_8 FILLER_65_3255 ();
 sg13g2_decap_8 FILLER_65_3262 ();
 sg13g2_decap_8 FILLER_65_3269 ();
 sg13g2_decap_8 FILLER_65_3276 ();
 sg13g2_decap_8 FILLER_65_3283 ();
 sg13g2_decap_8 FILLER_65_3290 ();
 sg13g2_decap_8 FILLER_65_3297 ();
 sg13g2_decap_8 FILLER_65_3304 ();
 sg13g2_decap_8 FILLER_65_3311 ();
 sg13g2_decap_8 FILLER_65_3318 ();
 sg13g2_decap_8 FILLER_65_3325 ();
 sg13g2_decap_8 FILLER_65_3332 ();
 sg13g2_decap_8 FILLER_65_3339 ();
 sg13g2_decap_8 FILLER_65_3346 ();
 sg13g2_decap_8 FILLER_65_3353 ();
 sg13g2_decap_8 FILLER_65_3360 ();
 sg13g2_decap_8 FILLER_65_3367 ();
 sg13g2_decap_8 FILLER_65_3374 ();
 sg13g2_decap_8 FILLER_65_3381 ();
 sg13g2_decap_8 FILLER_65_3388 ();
 sg13g2_decap_8 FILLER_65_3395 ();
 sg13g2_decap_8 FILLER_65_3402 ();
 sg13g2_decap_8 FILLER_65_3409 ();
 sg13g2_decap_8 FILLER_65_3416 ();
 sg13g2_decap_8 FILLER_65_3423 ();
 sg13g2_decap_8 FILLER_65_3430 ();
 sg13g2_decap_8 FILLER_65_3437 ();
 sg13g2_decap_8 FILLER_65_3444 ();
 sg13g2_decap_8 FILLER_65_3451 ();
 sg13g2_decap_8 FILLER_65_3458 ();
 sg13g2_decap_8 FILLER_65_3465 ();
 sg13g2_decap_8 FILLER_65_3472 ();
 sg13g2_decap_8 FILLER_65_3479 ();
 sg13g2_decap_8 FILLER_65_3486 ();
 sg13g2_decap_8 FILLER_65_3493 ();
 sg13g2_decap_8 FILLER_65_3500 ();
 sg13g2_decap_8 FILLER_65_3507 ();
 sg13g2_decap_8 FILLER_65_3514 ();
 sg13g2_decap_8 FILLER_65_3521 ();
 sg13g2_decap_8 FILLER_65_3528 ();
 sg13g2_decap_8 FILLER_65_3535 ();
 sg13g2_decap_8 FILLER_65_3542 ();
 sg13g2_decap_8 FILLER_65_3549 ();
 sg13g2_decap_8 FILLER_65_3556 ();
 sg13g2_decap_8 FILLER_65_3563 ();
 sg13g2_decap_8 FILLER_65_3570 ();
 sg13g2_fill_2 FILLER_65_3577 ();
 sg13g2_fill_1 FILLER_65_3579 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_decap_8 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_decap_8 FILLER_66_112 ();
 sg13g2_decap_8 FILLER_66_119 ();
 sg13g2_decap_8 FILLER_66_126 ();
 sg13g2_decap_8 FILLER_66_133 ();
 sg13g2_decap_8 FILLER_66_140 ();
 sg13g2_decap_8 FILLER_66_147 ();
 sg13g2_decap_8 FILLER_66_154 ();
 sg13g2_decap_8 FILLER_66_161 ();
 sg13g2_decap_8 FILLER_66_168 ();
 sg13g2_decap_8 FILLER_66_175 ();
 sg13g2_decap_8 FILLER_66_182 ();
 sg13g2_decap_8 FILLER_66_189 ();
 sg13g2_decap_8 FILLER_66_196 ();
 sg13g2_decap_8 FILLER_66_203 ();
 sg13g2_decap_8 FILLER_66_210 ();
 sg13g2_decap_8 FILLER_66_217 ();
 sg13g2_decap_8 FILLER_66_224 ();
 sg13g2_decap_8 FILLER_66_231 ();
 sg13g2_decap_8 FILLER_66_238 ();
 sg13g2_decap_8 FILLER_66_245 ();
 sg13g2_decap_8 FILLER_66_252 ();
 sg13g2_decap_8 FILLER_66_259 ();
 sg13g2_decap_8 FILLER_66_266 ();
 sg13g2_decap_8 FILLER_66_273 ();
 sg13g2_decap_8 FILLER_66_280 ();
 sg13g2_decap_8 FILLER_66_287 ();
 sg13g2_decap_8 FILLER_66_294 ();
 sg13g2_decap_8 FILLER_66_301 ();
 sg13g2_decap_8 FILLER_66_308 ();
 sg13g2_decap_8 FILLER_66_315 ();
 sg13g2_decap_8 FILLER_66_322 ();
 sg13g2_decap_8 FILLER_66_329 ();
 sg13g2_decap_8 FILLER_66_336 ();
 sg13g2_decap_8 FILLER_66_343 ();
 sg13g2_decap_8 FILLER_66_350 ();
 sg13g2_decap_8 FILLER_66_357 ();
 sg13g2_decap_8 FILLER_66_364 ();
 sg13g2_decap_8 FILLER_66_371 ();
 sg13g2_decap_8 FILLER_66_378 ();
 sg13g2_decap_8 FILLER_66_385 ();
 sg13g2_decap_8 FILLER_66_392 ();
 sg13g2_decap_8 FILLER_66_399 ();
 sg13g2_decap_8 FILLER_66_406 ();
 sg13g2_decap_8 FILLER_66_413 ();
 sg13g2_decap_8 FILLER_66_420 ();
 sg13g2_decap_8 FILLER_66_427 ();
 sg13g2_decap_8 FILLER_66_434 ();
 sg13g2_decap_8 FILLER_66_441 ();
 sg13g2_decap_8 FILLER_66_448 ();
 sg13g2_decap_8 FILLER_66_455 ();
 sg13g2_decap_8 FILLER_66_462 ();
 sg13g2_decap_8 FILLER_66_469 ();
 sg13g2_decap_8 FILLER_66_476 ();
 sg13g2_decap_8 FILLER_66_483 ();
 sg13g2_decap_8 FILLER_66_490 ();
 sg13g2_decap_8 FILLER_66_497 ();
 sg13g2_decap_8 FILLER_66_504 ();
 sg13g2_decap_8 FILLER_66_511 ();
 sg13g2_decap_8 FILLER_66_518 ();
 sg13g2_decap_8 FILLER_66_525 ();
 sg13g2_decap_8 FILLER_66_532 ();
 sg13g2_decap_8 FILLER_66_539 ();
 sg13g2_decap_8 FILLER_66_546 ();
 sg13g2_decap_8 FILLER_66_553 ();
 sg13g2_decap_8 FILLER_66_560 ();
 sg13g2_decap_8 FILLER_66_567 ();
 sg13g2_decap_8 FILLER_66_574 ();
 sg13g2_decap_8 FILLER_66_581 ();
 sg13g2_decap_8 FILLER_66_588 ();
 sg13g2_decap_8 FILLER_66_595 ();
 sg13g2_decap_8 FILLER_66_602 ();
 sg13g2_decap_8 FILLER_66_609 ();
 sg13g2_decap_8 FILLER_66_616 ();
 sg13g2_decap_8 FILLER_66_623 ();
 sg13g2_decap_8 FILLER_66_630 ();
 sg13g2_decap_8 FILLER_66_637 ();
 sg13g2_decap_8 FILLER_66_644 ();
 sg13g2_decap_8 FILLER_66_651 ();
 sg13g2_decap_8 FILLER_66_658 ();
 sg13g2_decap_8 FILLER_66_665 ();
 sg13g2_decap_8 FILLER_66_672 ();
 sg13g2_decap_8 FILLER_66_679 ();
 sg13g2_decap_8 FILLER_66_686 ();
 sg13g2_decap_8 FILLER_66_693 ();
 sg13g2_decap_8 FILLER_66_700 ();
 sg13g2_decap_8 FILLER_66_707 ();
 sg13g2_decap_8 FILLER_66_714 ();
 sg13g2_decap_8 FILLER_66_721 ();
 sg13g2_decap_8 FILLER_66_728 ();
 sg13g2_decap_8 FILLER_66_735 ();
 sg13g2_decap_8 FILLER_66_742 ();
 sg13g2_decap_8 FILLER_66_749 ();
 sg13g2_decap_8 FILLER_66_756 ();
 sg13g2_decap_8 FILLER_66_763 ();
 sg13g2_decap_8 FILLER_66_770 ();
 sg13g2_decap_8 FILLER_66_777 ();
 sg13g2_decap_8 FILLER_66_784 ();
 sg13g2_decap_8 FILLER_66_791 ();
 sg13g2_decap_8 FILLER_66_798 ();
 sg13g2_decap_8 FILLER_66_805 ();
 sg13g2_decap_8 FILLER_66_812 ();
 sg13g2_decap_8 FILLER_66_819 ();
 sg13g2_decap_8 FILLER_66_826 ();
 sg13g2_decap_8 FILLER_66_833 ();
 sg13g2_decap_8 FILLER_66_840 ();
 sg13g2_decap_8 FILLER_66_847 ();
 sg13g2_decap_8 FILLER_66_854 ();
 sg13g2_decap_8 FILLER_66_861 ();
 sg13g2_decap_8 FILLER_66_868 ();
 sg13g2_decap_8 FILLER_66_875 ();
 sg13g2_decap_8 FILLER_66_882 ();
 sg13g2_decap_8 FILLER_66_889 ();
 sg13g2_decap_8 FILLER_66_896 ();
 sg13g2_decap_8 FILLER_66_903 ();
 sg13g2_decap_8 FILLER_66_910 ();
 sg13g2_decap_8 FILLER_66_917 ();
 sg13g2_decap_8 FILLER_66_924 ();
 sg13g2_decap_8 FILLER_66_931 ();
 sg13g2_decap_8 FILLER_66_938 ();
 sg13g2_decap_8 FILLER_66_945 ();
 sg13g2_decap_8 FILLER_66_952 ();
 sg13g2_decap_8 FILLER_66_959 ();
 sg13g2_decap_8 FILLER_66_966 ();
 sg13g2_decap_8 FILLER_66_973 ();
 sg13g2_decap_8 FILLER_66_980 ();
 sg13g2_decap_8 FILLER_66_987 ();
 sg13g2_decap_8 FILLER_66_994 ();
 sg13g2_decap_8 FILLER_66_1001 ();
 sg13g2_decap_8 FILLER_66_1008 ();
 sg13g2_decap_8 FILLER_66_1015 ();
 sg13g2_decap_8 FILLER_66_1022 ();
 sg13g2_decap_8 FILLER_66_1029 ();
 sg13g2_decap_8 FILLER_66_1036 ();
 sg13g2_decap_8 FILLER_66_1043 ();
 sg13g2_decap_8 FILLER_66_1050 ();
 sg13g2_decap_8 FILLER_66_1057 ();
 sg13g2_decap_8 FILLER_66_1064 ();
 sg13g2_decap_8 FILLER_66_1071 ();
 sg13g2_decap_8 FILLER_66_1078 ();
 sg13g2_decap_8 FILLER_66_1085 ();
 sg13g2_decap_8 FILLER_66_1092 ();
 sg13g2_decap_8 FILLER_66_1099 ();
 sg13g2_decap_8 FILLER_66_1106 ();
 sg13g2_decap_8 FILLER_66_1113 ();
 sg13g2_decap_8 FILLER_66_1120 ();
 sg13g2_decap_8 FILLER_66_1127 ();
 sg13g2_decap_8 FILLER_66_1134 ();
 sg13g2_decap_8 FILLER_66_1141 ();
 sg13g2_decap_8 FILLER_66_1148 ();
 sg13g2_decap_8 FILLER_66_1155 ();
 sg13g2_decap_8 FILLER_66_1162 ();
 sg13g2_decap_8 FILLER_66_1169 ();
 sg13g2_decap_8 FILLER_66_1176 ();
 sg13g2_decap_8 FILLER_66_1183 ();
 sg13g2_decap_8 FILLER_66_1190 ();
 sg13g2_decap_8 FILLER_66_1197 ();
 sg13g2_decap_8 FILLER_66_1204 ();
 sg13g2_decap_8 FILLER_66_1211 ();
 sg13g2_decap_8 FILLER_66_1218 ();
 sg13g2_decap_8 FILLER_66_1225 ();
 sg13g2_decap_8 FILLER_66_1232 ();
 sg13g2_decap_8 FILLER_66_1239 ();
 sg13g2_decap_8 FILLER_66_1246 ();
 sg13g2_decap_8 FILLER_66_1253 ();
 sg13g2_decap_8 FILLER_66_1260 ();
 sg13g2_decap_8 FILLER_66_1267 ();
 sg13g2_decap_8 FILLER_66_1274 ();
 sg13g2_decap_8 FILLER_66_1281 ();
 sg13g2_decap_8 FILLER_66_1288 ();
 sg13g2_decap_8 FILLER_66_1295 ();
 sg13g2_decap_8 FILLER_66_1302 ();
 sg13g2_decap_8 FILLER_66_1309 ();
 sg13g2_decap_8 FILLER_66_1316 ();
 sg13g2_decap_8 FILLER_66_1323 ();
 sg13g2_decap_8 FILLER_66_1330 ();
 sg13g2_decap_8 FILLER_66_1337 ();
 sg13g2_decap_8 FILLER_66_1344 ();
 sg13g2_decap_8 FILLER_66_1351 ();
 sg13g2_decap_8 FILLER_66_1358 ();
 sg13g2_decap_8 FILLER_66_1365 ();
 sg13g2_decap_8 FILLER_66_1372 ();
 sg13g2_decap_8 FILLER_66_1379 ();
 sg13g2_decap_8 FILLER_66_1386 ();
 sg13g2_decap_8 FILLER_66_1393 ();
 sg13g2_decap_8 FILLER_66_1400 ();
 sg13g2_decap_8 FILLER_66_1407 ();
 sg13g2_decap_8 FILLER_66_1414 ();
 sg13g2_decap_8 FILLER_66_1421 ();
 sg13g2_decap_8 FILLER_66_1428 ();
 sg13g2_decap_8 FILLER_66_1435 ();
 sg13g2_decap_8 FILLER_66_1442 ();
 sg13g2_decap_8 FILLER_66_1449 ();
 sg13g2_decap_8 FILLER_66_1456 ();
 sg13g2_decap_8 FILLER_66_1463 ();
 sg13g2_decap_8 FILLER_66_1470 ();
 sg13g2_decap_8 FILLER_66_1477 ();
 sg13g2_decap_8 FILLER_66_1484 ();
 sg13g2_decap_8 FILLER_66_1491 ();
 sg13g2_decap_8 FILLER_66_1498 ();
 sg13g2_decap_8 FILLER_66_1505 ();
 sg13g2_decap_8 FILLER_66_1512 ();
 sg13g2_decap_8 FILLER_66_1519 ();
 sg13g2_decap_8 FILLER_66_1526 ();
 sg13g2_decap_8 FILLER_66_1533 ();
 sg13g2_decap_8 FILLER_66_1540 ();
 sg13g2_decap_8 FILLER_66_1547 ();
 sg13g2_decap_8 FILLER_66_1554 ();
 sg13g2_decap_8 FILLER_66_1561 ();
 sg13g2_decap_8 FILLER_66_1568 ();
 sg13g2_decap_8 FILLER_66_1575 ();
 sg13g2_decap_8 FILLER_66_1582 ();
 sg13g2_decap_8 FILLER_66_1589 ();
 sg13g2_decap_8 FILLER_66_1596 ();
 sg13g2_decap_8 FILLER_66_1603 ();
 sg13g2_decap_8 FILLER_66_1610 ();
 sg13g2_decap_8 FILLER_66_1617 ();
 sg13g2_decap_8 FILLER_66_1624 ();
 sg13g2_decap_8 FILLER_66_1631 ();
 sg13g2_decap_8 FILLER_66_1638 ();
 sg13g2_decap_8 FILLER_66_1645 ();
 sg13g2_decap_8 FILLER_66_1652 ();
 sg13g2_decap_8 FILLER_66_1659 ();
 sg13g2_decap_8 FILLER_66_1666 ();
 sg13g2_decap_8 FILLER_66_1673 ();
 sg13g2_decap_8 FILLER_66_1680 ();
 sg13g2_decap_8 FILLER_66_1687 ();
 sg13g2_decap_8 FILLER_66_1694 ();
 sg13g2_decap_8 FILLER_66_1701 ();
 sg13g2_decap_8 FILLER_66_1708 ();
 sg13g2_decap_8 FILLER_66_1715 ();
 sg13g2_decap_8 FILLER_66_1722 ();
 sg13g2_decap_8 FILLER_66_1729 ();
 sg13g2_decap_8 FILLER_66_1736 ();
 sg13g2_decap_8 FILLER_66_1743 ();
 sg13g2_decap_8 FILLER_66_1750 ();
 sg13g2_decap_8 FILLER_66_1757 ();
 sg13g2_decap_8 FILLER_66_1764 ();
 sg13g2_decap_8 FILLER_66_1771 ();
 sg13g2_decap_8 FILLER_66_1778 ();
 sg13g2_decap_8 FILLER_66_1785 ();
 sg13g2_decap_8 FILLER_66_1792 ();
 sg13g2_decap_8 FILLER_66_1799 ();
 sg13g2_decap_8 FILLER_66_1806 ();
 sg13g2_decap_8 FILLER_66_1813 ();
 sg13g2_decap_8 FILLER_66_1820 ();
 sg13g2_decap_8 FILLER_66_1827 ();
 sg13g2_decap_8 FILLER_66_1834 ();
 sg13g2_decap_8 FILLER_66_1841 ();
 sg13g2_decap_8 FILLER_66_1848 ();
 sg13g2_decap_8 FILLER_66_1855 ();
 sg13g2_decap_8 FILLER_66_1862 ();
 sg13g2_decap_8 FILLER_66_1869 ();
 sg13g2_decap_8 FILLER_66_1876 ();
 sg13g2_decap_8 FILLER_66_1883 ();
 sg13g2_decap_8 FILLER_66_1890 ();
 sg13g2_decap_8 FILLER_66_1897 ();
 sg13g2_decap_8 FILLER_66_1904 ();
 sg13g2_decap_8 FILLER_66_1911 ();
 sg13g2_decap_8 FILLER_66_1918 ();
 sg13g2_decap_8 FILLER_66_1925 ();
 sg13g2_decap_8 FILLER_66_1932 ();
 sg13g2_decap_8 FILLER_66_1939 ();
 sg13g2_decap_8 FILLER_66_1946 ();
 sg13g2_decap_8 FILLER_66_1953 ();
 sg13g2_decap_8 FILLER_66_1960 ();
 sg13g2_decap_8 FILLER_66_1967 ();
 sg13g2_decap_8 FILLER_66_1974 ();
 sg13g2_decap_8 FILLER_66_1981 ();
 sg13g2_decap_8 FILLER_66_1988 ();
 sg13g2_decap_8 FILLER_66_1995 ();
 sg13g2_decap_8 FILLER_66_2002 ();
 sg13g2_decap_8 FILLER_66_2009 ();
 sg13g2_decap_8 FILLER_66_2016 ();
 sg13g2_decap_8 FILLER_66_2023 ();
 sg13g2_decap_8 FILLER_66_2030 ();
 sg13g2_decap_8 FILLER_66_2037 ();
 sg13g2_decap_8 FILLER_66_2044 ();
 sg13g2_decap_8 FILLER_66_2051 ();
 sg13g2_decap_8 FILLER_66_2058 ();
 sg13g2_decap_8 FILLER_66_2065 ();
 sg13g2_decap_8 FILLER_66_2072 ();
 sg13g2_decap_8 FILLER_66_2079 ();
 sg13g2_decap_8 FILLER_66_2086 ();
 sg13g2_decap_8 FILLER_66_2093 ();
 sg13g2_decap_8 FILLER_66_2100 ();
 sg13g2_decap_8 FILLER_66_2107 ();
 sg13g2_decap_8 FILLER_66_2114 ();
 sg13g2_decap_8 FILLER_66_2121 ();
 sg13g2_decap_8 FILLER_66_2128 ();
 sg13g2_decap_8 FILLER_66_2135 ();
 sg13g2_decap_8 FILLER_66_2142 ();
 sg13g2_decap_8 FILLER_66_2149 ();
 sg13g2_decap_8 FILLER_66_2156 ();
 sg13g2_decap_8 FILLER_66_2163 ();
 sg13g2_decap_8 FILLER_66_2170 ();
 sg13g2_decap_8 FILLER_66_2177 ();
 sg13g2_decap_8 FILLER_66_2184 ();
 sg13g2_decap_8 FILLER_66_2191 ();
 sg13g2_decap_8 FILLER_66_2198 ();
 sg13g2_decap_8 FILLER_66_2205 ();
 sg13g2_decap_8 FILLER_66_2212 ();
 sg13g2_decap_8 FILLER_66_2219 ();
 sg13g2_decap_8 FILLER_66_2226 ();
 sg13g2_decap_8 FILLER_66_2233 ();
 sg13g2_decap_8 FILLER_66_2240 ();
 sg13g2_decap_8 FILLER_66_2247 ();
 sg13g2_decap_8 FILLER_66_2254 ();
 sg13g2_decap_8 FILLER_66_2261 ();
 sg13g2_decap_8 FILLER_66_2268 ();
 sg13g2_decap_8 FILLER_66_2275 ();
 sg13g2_decap_8 FILLER_66_2282 ();
 sg13g2_decap_8 FILLER_66_2289 ();
 sg13g2_decap_8 FILLER_66_2296 ();
 sg13g2_decap_8 FILLER_66_2303 ();
 sg13g2_decap_8 FILLER_66_2310 ();
 sg13g2_decap_8 FILLER_66_2317 ();
 sg13g2_decap_8 FILLER_66_2324 ();
 sg13g2_decap_8 FILLER_66_2331 ();
 sg13g2_decap_8 FILLER_66_2338 ();
 sg13g2_decap_8 FILLER_66_2345 ();
 sg13g2_decap_8 FILLER_66_2352 ();
 sg13g2_decap_8 FILLER_66_2359 ();
 sg13g2_decap_8 FILLER_66_2366 ();
 sg13g2_decap_8 FILLER_66_2373 ();
 sg13g2_decap_8 FILLER_66_2380 ();
 sg13g2_decap_8 FILLER_66_2387 ();
 sg13g2_decap_8 FILLER_66_2394 ();
 sg13g2_decap_8 FILLER_66_2401 ();
 sg13g2_decap_8 FILLER_66_2408 ();
 sg13g2_decap_8 FILLER_66_2415 ();
 sg13g2_decap_8 FILLER_66_2422 ();
 sg13g2_decap_8 FILLER_66_2429 ();
 sg13g2_decap_8 FILLER_66_2436 ();
 sg13g2_decap_8 FILLER_66_2443 ();
 sg13g2_decap_8 FILLER_66_2450 ();
 sg13g2_decap_8 FILLER_66_2457 ();
 sg13g2_decap_8 FILLER_66_2464 ();
 sg13g2_decap_8 FILLER_66_2471 ();
 sg13g2_decap_8 FILLER_66_2478 ();
 sg13g2_decap_8 FILLER_66_2485 ();
 sg13g2_decap_8 FILLER_66_2492 ();
 sg13g2_decap_8 FILLER_66_2499 ();
 sg13g2_decap_8 FILLER_66_2506 ();
 sg13g2_decap_8 FILLER_66_2513 ();
 sg13g2_decap_8 FILLER_66_2520 ();
 sg13g2_decap_8 FILLER_66_2527 ();
 sg13g2_decap_8 FILLER_66_2534 ();
 sg13g2_decap_8 FILLER_66_2541 ();
 sg13g2_decap_8 FILLER_66_2548 ();
 sg13g2_decap_8 FILLER_66_2555 ();
 sg13g2_decap_8 FILLER_66_2562 ();
 sg13g2_decap_8 FILLER_66_2569 ();
 sg13g2_decap_8 FILLER_66_2576 ();
 sg13g2_decap_8 FILLER_66_2583 ();
 sg13g2_decap_8 FILLER_66_2590 ();
 sg13g2_decap_8 FILLER_66_2597 ();
 sg13g2_decap_8 FILLER_66_2604 ();
 sg13g2_decap_8 FILLER_66_2611 ();
 sg13g2_decap_8 FILLER_66_2618 ();
 sg13g2_decap_8 FILLER_66_2625 ();
 sg13g2_decap_8 FILLER_66_2632 ();
 sg13g2_decap_8 FILLER_66_2639 ();
 sg13g2_decap_8 FILLER_66_2646 ();
 sg13g2_decap_8 FILLER_66_2653 ();
 sg13g2_decap_8 FILLER_66_2660 ();
 sg13g2_decap_8 FILLER_66_2667 ();
 sg13g2_decap_8 FILLER_66_2674 ();
 sg13g2_decap_8 FILLER_66_2681 ();
 sg13g2_decap_8 FILLER_66_2688 ();
 sg13g2_decap_8 FILLER_66_2695 ();
 sg13g2_decap_8 FILLER_66_2702 ();
 sg13g2_decap_8 FILLER_66_2709 ();
 sg13g2_decap_8 FILLER_66_2716 ();
 sg13g2_decap_8 FILLER_66_2723 ();
 sg13g2_decap_8 FILLER_66_2730 ();
 sg13g2_decap_8 FILLER_66_2737 ();
 sg13g2_decap_8 FILLER_66_2744 ();
 sg13g2_decap_8 FILLER_66_2751 ();
 sg13g2_decap_8 FILLER_66_2758 ();
 sg13g2_decap_8 FILLER_66_2765 ();
 sg13g2_decap_8 FILLER_66_2772 ();
 sg13g2_decap_8 FILLER_66_2779 ();
 sg13g2_decap_8 FILLER_66_2786 ();
 sg13g2_decap_8 FILLER_66_2793 ();
 sg13g2_decap_8 FILLER_66_2800 ();
 sg13g2_decap_8 FILLER_66_2807 ();
 sg13g2_decap_8 FILLER_66_2814 ();
 sg13g2_decap_8 FILLER_66_2821 ();
 sg13g2_decap_8 FILLER_66_2828 ();
 sg13g2_decap_8 FILLER_66_2835 ();
 sg13g2_decap_8 FILLER_66_2842 ();
 sg13g2_decap_8 FILLER_66_2849 ();
 sg13g2_decap_8 FILLER_66_2856 ();
 sg13g2_decap_8 FILLER_66_2863 ();
 sg13g2_decap_8 FILLER_66_2870 ();
 sg13g2_decap_8 FILLER_66_2877 ();
 sg13g2_decap_8 FILLER_66_2884 ();
 sg13g2_decap_8 FILLER_66_2891 ();
 sg13g2_decap_8 FILLER_66_2898 ();
 sg13g2_decap_8 FILLER_66_2905 ();
 sg13g2_decap_8 FILLER_66_2912 ();
 sg13g2_decap_8 FILLER_66_2919 ();
 sg13g2_decap_8 FILLER_66_2926 ();
 sg13g2_decap_8 FILLER_66_2933 ();
 sg13g2_decap_8 FILLER_66_2940 ();
 sg13g2_decap_8 FILLER_66_2947 ();
 sg13g2_decap_8 FILLER_66_2954 ();
 sg13g2_decap_8 FILLER_66_2961 ();
 sg13g2_decap_8 FILLER_66_2968 ();
 sg13g2_decap_8 FILLER_66_2975 ();
 sg13g2_decap_8 FILLER_66_2982 ();
 sg13g2_decap_8 FILLER_66_2989 ();
 sg13g2_decap_8 FILLER_66_2996 ();
 sg13g2_decap_8 FILLER_66_3003 ();
 sg13g2_decap_8 FILLER_66_3010 ();
 sg13g2_decap_8 FILLER_66_3017 ();
 sg13g2_decap_8 FILLER_66_3024 ();
 sg13g2_decap_8 FILLER_66_3031 ();
 sg13g2_decap_8 FILLER_66_3038 ();
 sg13g2_decap_8 FILLER_66_3045 ();
 sg13g2_decap_8 FILLER_66_3052 ();
 sg13g2_decap_8 FILLER_66_3059 ();
 sg13g2_decap_8 FILLER_66_3066 ();
 sg13g2_decap_8 FILLER_66_3073 ();
 sg13g2_decap_8 FILLER_66_3080 ();
 sg13g2_decap_8 FILLER_66_3087 ();
 sg13g2_decap_8 FILLER_66_3094 ();
 sg13g2_decap_8 FILLER_66_3101 ();
 sg13g2_decap_8 FILLER_66_3108 ();
 sg13g2_decap_8 FILLER_66_3115 ();
 sg13g2_decap_8 FILLER_66_3122 ();
 sg13g2_decap_8 FILLER_66_3129 ();
 sg13g2_decap_8 FILLER_66_3136 ();
 sg13g2_decap_8 FILLER_66_3143 ();
 sg13g2_decap_8 FILLER_66_3150 ();
 sg13g2_decap_8 FILLER_66_3157 ();
 sg13g2_decap_8 FILLER_66_3164 ();
 sg13g2_decap_8 FILLER_66_3171 ();
 sg13g2_decap_8 FILLER_66_3178 ();
 sg13g2_decap_8 FILLER_66_3185 ();
 sg13g2_decap_8 FILLER_66_3192 ();
 sg13g2_decap_8 FILLER_66_3199 ();
 sg13g2_decap_8 FILLER_66_3206 ();
 sg13g2_decap_8 FILLER_66_3213 ();
 sg13g2_decap_8 FILLER_66_3220 ();
 sg13g2_decap_8 FILLER_66_3227 ();
 sg13g2_decap_8 FILLER_66_3234 ();
 sg13g2_decap_8 FILLER_66_3241 ();
 sg13g2_decap_8 FILLER_66_3248 ();
 sg13g2_decap_8 FILLER_66_3255 ();
 sg13g2_decap_8 FILLER_66_3262 ();
 sg13g2_decap_8 FILLER_66_3269 ();
 sg13g2_decap_8 FILLER_66_3276 ();
 sg13g2_decap_8 FILLER_66_3283 ();
 sg13g2_decap_8 FILLER_66_3290 ();
 sg13g2_decap_8 FILLER_66_3297 ();
 sg13g2_decap_8 FILLER_66_3304 ();
 sg13g2_decap_8 FILLER_66_3311 ();
 sg13g2_decap_8 FILLER_66_3318 ();
 sg13g2_decap_8 FILLER_66_3325 ();
 sg13g2_decap_8 FILLER_66_3332 ();
 sg13g2_decap_8 FILLER_66_3339 ();
 sg13g2_decap_8 FILLER_66_3346 ();
 sg13g2_decap_8 FILLER_66_3353 ();
 sg13g2_decap_8 FILLER_66_3360 ();
 sg13g2_decap_8 FILLER_66_3367 ();
 sg13g2_decap_8 FILLER_66_3374 ();
 sg13g2_decap_8 FILLER_66_3381 ();
 sg13g2_decap_8 FILLER_66_3388 ();
 sg13g2_decap_8 FILLER_66_3395 ();
 sg13g2_decap_8 FILLER_66_3402 ();
 sg13g2_decap_8 FILLER_66_3409 ();
 sg13g2_decap_8 FILLER_66_3416 ();
 sg13g2_decap_8 FILLER_66_3423 ();
 sg13g2_decap_8 FILLER_66_3430 ();
 sg13g2_decap_8 FILLER_66_3437 ();
 sg13g2_decap_8 FILLER_66_3444 ();
 sg13g2_decap_8 FILLER_66_3451 ();
 sg13g2_decap_8 FILLER_66_3458 ();
 sg13g2_decap_8 FILLER_66_3465 ();
 sg13g2_decap_8 FILLER_66_3472 ();
 sg13g2_decap_8 FILLER_66_3479 ();
 sg13g2_decap_8 FILLER_66_3486 ();
 sg13g2_decap_8 FILLER_66_3493 ();
 sg13g2_decap_8 FILLER_66_3500 ();
 sg13g2_decap_8 FILLER_66_3507 ();
 sg13g2_decap_8 FILLER_66_3514 ();
 sg13g2_decap_8 FILLER_66_3521 ();
 sg13g2_decap_8 FILLER_66_3528 ();
 sg13g2_decap_8 FILLER_66_3535 ();
 sg13g2_decap_8 FILLER_66_3542 ();
 sg13g2_decap_8 FILLER_66_3549 ();
 sg13g2_decap_8 FILLER_66_3556 ();
 sg13g2_decap_8 FILLER_66_3563 ();
 sg13g2_decap_8 FILLER_66_3570 ();
 sg13g2_fill_2 FILLER_66_3577 ();
 sg13g2_fill_1 FILLER_66_3579 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_decap_8 FILLER_67_112 ();
 sg13g2_decap_8 FILLER_67_119 ();
 sg13g2_decap_8 FILLER_67_126 ();
 sg13g2_decap_8 FILLER_67_133 ();
 sg13g2_decap_8 FILLER_67_140 ();
 sg13g2_decap_8 FILLER_67_147 ();
 sg13g2_decap_8 FILLER_67_154 ();
 sg13g2_decap_8 FILLER_67_161 ();
 sg13g2_decap_8 FILLER_67_168 ();
 sg13g2_decap_8 FILLER_67_175 ();
 sg13g2_decap_8 FILLER_67_182 ();
 sg13g2_decap_8 FILLER_67_189 ();
 sg13g2_decap_8 FILLER_67_196 ();
 sg13g2_decap_8 FILLER_67_203 ();
 sg13g2_decap_8 FILLER_67_210 ();
 sg13g2_decap_8 FILLER_67_217 ();
 sg13g2_decap_8 FILLER_67_224 ();
 sg13g2_decap_8 FILLER_67_231 ();
 sg13g2_decap_8 FILLER_67_238 ();
 sg13g2_decap_8 FILLER_67_245 ();
 sg13g2_decap_8 FILLER_67_252 ();
 sg13g2_decap_8 FILLER_67_259 ();
 sg13g2_decap_8 FILLER_67_266 ();
 sg13g2_decap_8 FILLER_67_273 ();
 sg13g2_decap_8 FILLER_67_280 ();
 sg13g2_decap_8 FILLER_67_287 ();
 sg13g2_decap_8 FILLER_67_294 ();
 sg13g2_decap_8 FILLER_67_301 ();
 sg13g2_decap_8 FILLER_67_308 ();
 sg13g2_decap_8 FILLER_67_315 ();
 sg13g2_decap_8 FILLER_67_322 ();
 sg13g2_decap_8 FILLER_67_329 ();
 sg13g2_decap_8 FILLER_67_336 ();
 sg13g2_decap_8 FILLER_67_343 ();
 sg13g2_decap_8 FILLER_67_350 ();
 sg13g2_decap_8 FILLER_67_357 ();
 sg13g2_decap_8 FILLER_67_364 ();
 sg13g2_decap_8 FILLER_67_371 ();
 sg13g2_decap_8 FILLER_67_378 ();
 sg13g2_decap_8 FILLER_67_385 ();
 sg13g2_decap_8 FILLER_67_392 ();
 sg13g2_decap_8 FILLER_67_399 ();
 sg13g2_decap_8 FILLER_67_406 ();
 sg13g2_decap_8 FILLER_67_413 ();
 sg13g2_decap_8 FILLER_67_420 ();
 sg13g2_decap_8 FILLER_67_427 ();
 sg13g2_decap_8 FILLER_67_434 ();
 sg13g2_decap_8 FILLER_67_441 ();
 sg13g2_decap_8 FILLER_67_448 ();
 sg13g2_decap_8 FILLER_67_455 ();
 sg13g2_decap_8 FILLER_67_462 ();
 sg13g2_decap_8 FILLER_67_469 ();
 sg13g2_decap_8 FILLER_67_476 ();
 sg13g2_decap_8 FILLER_67_483 ();
 sg13g2_decap_8 FILLER_67_490 ();
 sg13g2_decap_8 FILLER_67_497 ();
 sg13g2_decap_8 FILLER_67_504 ();
 sg13g2_decap_8 FILLER_67_511 ();
 sg13g2_decap_8 FILLER_67_518 ();
 sg13g2_decap_8 FILLER_67_525 ();
 sg13g2_decap_8 FILLER_67_532 ();
 sg13g2_decap_8 FILLER_67_539 ();
 sg13g2_decap_8 FILLER_67_546 ();
 sg13g2_decap_8 FILLER_67_553 ();
 sg13g2_decap_8 FILLER_67_560 ();
 sg13g2_decap_8 FILLER_67_567 ();
 sg13g2_decap_8 FILLER_67_574 ();
 sg13g2_decap_8 FILLER_67_581 ();
 sg13g2_decap_8 FILLER_67_588 ();
 sg13g2_decap_8 FILLER_67_595 ();
 sg13g2_decap_8 FILLER_67_602 ();
 sg13g2_decap_8 FILLER_67_609 ();
 sg13g2_decap_8 FILLER_67_616 ();
 sg13g2_decap_8 FILLER_67_623 ();
 sg13g2_decap_8 FILLER_67_630 ();
 sg13g2_decap_8 FILLER_67_637 ();
 sg13g2_decap_8 FILLER_67_644 ();
 sg13g2_decap_8 FILLER_67_651 ();
 sg13g2_decap_8 FILLER_67_658 ();
 sg13g2_decap_8 FILLER_67_665 ();
 sg13g2_decap_8 FILLER_67_672 ();
 sg13g2_decap_8 FILLER_67_679 ();
 sg13g2_decap_8 FILLER_67_686 ();
 sg13g2_decap_8 FILLER_67_693 ();
 sg13g2_decap_8 FILLER_67_700 ();
 sg13g2_decap_8 FILLER_67_707 ();
 sg13g2_decap_8 FILLER_67_714 ();
 sg13g2_decap_8 FILLER_67_721 ();
 sg13g2_decap_8 FILLER_67_728 ();
 sg13g2_decap_8 FILLER_67_735 ();
 sg13g2_decap_8 FILLER_67_742 ();
 sg13g2_decap_8 FILLER_67_749 ();
 sg13g2_decap_8 FILLER_67_756 ();
 sg13g2_decap_8 FILLER_67_763 ();
 sg13g2_decap_8 FILLER_67_770 ();
 sg13g2_decap_8 FILLER_67_777 ();
 sg13g2_decap_8 FILLER_67_784 ();
 sg13g2_decap_8 FILLER_67_791 ();
 sg13g2_decap_8 FILLER_67_798 ();
 sg13g2_decap_8 FILLER_67_805 ();
 sg13g2_decap_8 FILLER_67_812 ();
 sg13g2_decap_8 FILLER_67_819 ();
 sg13g2_decap_8 FILLER_67_826 ();
 sg13g2_decap_8 FILLER_67_833 ();
 sg13g2_decap_8 FILLER_67_840 ();
 sg13g2_decap_8 FILLER_67_847 ();
 sg13g2_decap_8 FILLER_67_854 ();
 sg13g2_decap_8 FILLER_67_861 ();
 sg13g2_decap_8 FILLER_67_868 ();
 sg13g2_decap_8 FILLER_67_875 ();
 sg13g2_decap_8 FILLER_67_882 ();
 sg13g2_decap_8 FILLER_67_889 ();
 sg13g2_decap_8 FILLER_67_896 ();
 sg13g2_decap_8 FILLER_67_903 ();
 sg13g2_decap_8 FILLER_67_910 ();
 sg13g2_decap_8 FILLER_67_917 ();
 sg13g2_decap_8 FILLER_67_924 ();
 sg13g2_decap_8 FILLER_67_931 ();
 sg13g2_decap_8 FILLER_67_938 ();
 sg13g2_decap_8 FILLER_67_945 ();
 sg13g2_decap_8 FILLER_67_952 ();
 sg13g2_decap_8 FILLER_67_959 ();
 sg13g2_decap_8 FILLER_67_966 ();
 sg13g2_decap_8 FILLER_67_973 ();
 sg13g2_decap_8 FILLER_67_980 ();
 sg13g2_decap_8 FILLER_67_987 ();
 sg13g2_decap_8 FILLER_67_994 ();
 sg13g2_decap_8 FILLER_67_1001 ();
 sg13g2_decap_8 FILLER_67_1008 ();
 sg13g2_decap_8 FILLER_67_1015 ();
 sg13g2_decap_8 FILLER_67_1022 ();
 sg13g2_decap_8 FILLER_67_1029 ();
 sg13g2_decap_8 FILLER_67_1036 ();
 sg13g2_decap_8 FILLER_67_1043 ();
 sg13g2_decap_8 FILLER_67_1050 ();
 sg13g2_decap_8 FILLER_67_1057 ();
 sg13g2_decap_8 FILLER_67_1064 ();
 sg13g2_decap_8 FILLER_67_1071 ();
 sg13g2_decap_8 FILLER_67_1078 ();
 sg13g2_decap_8 FILLER_67_1085 ();
 sg13g2_decap_8 FILLER_67_1092 ();
 sg13g2_decap_8 FILLER_67_1099 ();
 sg13g2_decap_8 FILLER_67_1106 ();
 sg13g2_decap_8 FILLER_67_1113 ();
 sg13g2_decap_8 FILLER_67_1120 ();
 sg13g2_decap_8 FILLER_67_1127 ();
 sg13g2_decap_8 FILLER_67_1134 ();
 sg13g2_decap_8 FILLER_67_1141 ();
 sg13g2_decap_8 FILLER_67_1148 ();
 sg13g2_decap_8 FILLER_67_1155 ();
 sg13g2_decap_8 FILLER_67_1162 ();
 sg13g2_decap_8 FILLER_67_1169 ();
 sg13g2_decap_8 FILLER_67_1176 ();
 sg13g2_decap_8 FILLER_67_1183 ();
 sg13g2_decap_8 FILLER_67_1190 ();
 sg13g2_decap_8 FILLER_67_1197 ();
 sg13g2_decap_8 FILLER_67_1204 ();
 sg13g2_decap_8 FILLER_67_1211 ();
 sg13g2_decap_8 FILLER_67_1218 ();
 sg13g2_decap_8 FILLER_67_1225 ();
 sg13g2_decap_8 FILLER_67_1232 ();
 sg13g2_decap_8 FILLER_67_1239 ();
 sg13g2_decap_8 FILLER_67_1246 ();
 sg13g2_decap_8 FILLER_67_1253 ();
 sg13g2_decap_8 FILLER_67_1260 ();
 sg13g2_decap_8 FILLER_67_1267 ();
 sg13g2_decap_8 FILLER_67_1274 ();
 sg13g2_decap_8 FILLER_67_1281 ();
 sg13g2_decap_8 FILLER_67_1288 ();
 sg13g2_decap_8 FILLER_67_1295 ();
 sg13g2_decap_8 FILLER_67_1302 ();
 sg13g2_decap_8 FILLER_67_1309 ();
 sg13g2_decap_8 FILLER_67_1316 ();
 sg13g2_decap_8 FILLER_67_1323 ();
 sg13g2_decap_8 FILLER_67_1330 ();
 sg13g2_decap_8 FILLER_67_1337 ();
 sg13g2_decap_8 FILLER_67_1344 ();
 sg13g2_decap_8 FILLER_67_1351 ();
 sg13g2_decap_8 FILLER_67_1358 ();
 sg13g2_decap_8 FILLER_67_1365 ();
 sg13g2_decap_8 FILLER_67_1372 ();
 sg13g2_decap_8 FILLER_67_1379 ();
 sg13g2_decap_8 FILLER_67_1386 ();
 sg13g2_decap_8 FILLER_67_1393 ();
 sg13g2_decap_8 FILLER_67_1400 ();
 sg13g2_decap_8 FILLER_67_1407 ();
 sg13g2_decap_8 FILLER_67_1414 ();
 sg13g2_decap_8 FILLER_67_1421 ();
 sg13g2_decap_8 FILLER_67_1428 ();
 sg13g2_decap_8 FILLER_67_1435 ();
 sg13g2_decap_8 FILLER_67_1442 ();
 sg13g2_decap_8 FILLER_67_1449 ();
 sg13g2_decap_8 FILLER_67_1456 ();
 sg13g2_decap_8 FILLER_67_1463 ();
 sg13g2_decap_8 FILLER_67_1470 ();
 sg13g2_decap_8 FILLER_67_1477 ();
 sg13g2_decap_8 FILLER_67_1484 ();
 sg13g2_decap_8 FILLER_67_1491 ();
 sg13g2_decap_8 FILLER_67_1498 ();
 sg13g2_decap_8 FILLER_67_1505 ();
 sg13g2_decap_8 FILLER_67_1512 ();
 sg13g2_decap_8 FILLER_67_1519 ();
 sg13g2_decap_8 FILLER_67_1526 ();
 sg13g2_decap_8 FILLER_67_1533 ();
 sg13g2_decap_8 FILLER_67_1540 ();
 sg13g2_decap_8 FILLER_67_1547 ();
 sg13g2_decap_8 FILLER_67_1554 ();
 sg13g2_decap_8 FILLER_67_1561 ();
 sg13g2_decap_8 FILLER_67_1568 ();
 sg13g2_decap_8 FILLER_67_1575 ();
 sg13g2_decap_8 FILLER_67_1582 ();
 sg13g2_decap_8 FILLER_67_1589 ();
 sg13g2_decap_8 FILLER_67_1596 ();
 sg13g2_decap_8 FILLER_67_1603 ();
 sg13g2_decap_8 FILLER_67_1610 ();
 sg13g2_decap_8 FILLER_67_1617 ();
 sg13g2_decap_8 FILLER_67_1624 ();
 sg13g2_decap_8 FILLER_67_1631 ();
 sg13g2_decap_8 FILLER_67_1638 ();
 sg13g2_decap_8 FILLER_67_1645 ();
 sg13g2_decap_8 FILLER_67_1652 ();
 sg13g2_decap_8 FILLER_67_1659 ();
 sg13g2_decap_8 FILLER_67_1666 ();
 sg13g2_decap_8 FILLER_67_1673 ();
 sg13g2_decap_8 FILLER_67_1680 ();
 sg13g2_decap_8 FILLER_67_1687 ();
 sg13g2_decap_8 FILLER_67_1694 ();
 sg13g2_decap_8 FILLER_67_1701 ();
 sg13g2_decap_8 FILLER_67_1708 ();
 sg13g2_decap_8 FILLER_67_1715 ();
 sg13g2_decap_8 FILLER_67_1722 ();
 sg13g2_decap_8 FILLER_67_1729 ();
 sg13g2_decap_8 FILLER_67_1736 ();
 sg13g2_decap_8 FILLER_67_1743 ();
 sg13g2_decap_8 FILLER_67_1750 ();
 sg13g2_decap_8 FILLER_67_1757 ();
 sg13g2_decap_8 FILLER_67_1764 ();
 sg13g2_decap_8 FILLER_67_1771 ();
 sg13g2_decap_8 FILLER_67_1778 ();
 sg13g2_decap_8 FILLER_67_1785 ();
 sg13g2_decap_8 FILLER_67_1792 ();
 sg13g2_decap_8 FILLER_67_1799 ();
 sg13g2_decap_8 FILLER_67_1806 ();
 sg13g2_decap_8 FILLER_67_1813 ();
 sg13g2_decap_8 FILLER_67_1820 ();
 sg13g2_decap_8 FILLER_67_1827 ();
 sg13g2_decap_8 FILLER_67_1834 ();
 sg13g2_decap_8 FILLER_67_1841 ();
 sg13g2_decap_8 FILLER_67_1848 ();
 sg13g2_decap_8 FILLER_67_1855 ();
 sg13g2_decap_8 FILLER_67_1862 ();
 sg13g2_decap_8 FILLER_67_1869 ();
 sg13g2_decap_8 FILLER_67_1876 ();
 sg13g2_decap_8 FILLER_67_1883 ();
 sg13g2_decap_8 FILLER_67_1890 ();
 sg13g2_decap_8 FILLER_67_1897 ();
 sg13g2_decap_8 FILLER_67_1904 ();
 sg13g2_decap_8 FILLER_67_1911 ();
 sg13g2_decap_8 FILLER_67_1918 ();
 sg13g2_decap_8 FILLER_67_1925 ();
 sg13g2_decap_8 FILLER_67_1932 ();
 sg13g2_decap_8 FILLER_67_1939 ();
 sg13g2_decap_8 FILLER_67_1946 ();
 sg13g2_decap_8 FILLER_67_1953 ();
 sg13g2_decap_8 FILLER_67_1960 ();
 sg13g2_decap_8 FILLER_67_1967 ();
 sg13g2_decap_8 FILLER_67_1974 ();
 sg13g2_decap_8 FILLER_67_1981 ();
 sg13g2_decap_8 FILLER_67_1988 ();
 sg13g2_decap_8 FILLER_67_1995 ();
 sg13g2_decap_8 FILLER_67_2002 ();
 sg13g2_decap_8 FILLER_67_2009 ();
 sg13g2_decap_8 FILLER_67_2016 ();
 sg13g2_decap_8 FILLER_67_2023 ();
 sg13g2_decap_8 FILLER_67_2030 ();
 sg13g2_decap_8 FILLER_67_2037 ();
 sg13g2_decap_8 FILLER_67_2044 ();
 sg13g2_decap_8 FILLER_67_2051 ();
 sg13g2_decap_8 FILLER_67_2058 ();
 sg13g2_decap_8 FILLER_67_2065 ();
 sg13g2_decap_8 FILLER_67_2072 ();
 sg13g2_decap_8 FILLER_67_2079 ();
 sg13g2_decap_8 FILLER_67_2086 ();
 sg13g2_decap_8 FILLER_67_2093 ();
 sg13g2_decap_8 FILLER_67_2100 ();
 sg13g2_decap_8 FILLER_67_2107 ();
 sg13g2_decap_8 FILLER_67_2114 ();
 sg13g2_decap_8 FILLER_67_2121 ();
 sg13g2_decap_8 FILLER_67_2128 ();
 sg13g2_decap_8 FILLER_67_2135 ();
 sg13g2_decap_8 FILLER_67_2142 ();
 sg13g2_decap_8 FILLER_67_2149 ();
 sg13g2_decap_8 FILLER_67_2156 ();
 sg13g2_decap_8 FILLER_67_2163 ();
 sg13g2_decap_8 FILLER_67_2170 ();
 sg13g2_decap_8 FILLER_67_2177 ();
 sg13g2_decap_8 FILLER_67_2184 ();
 sg13g2_decap_8 FILLER_67_2191 ();
 sg13g2_decap_8 FILLER_67_2198 ();
 sg13g2_decap_8 FILLER_67_2205 ();
 sg13g2_decap_8 FILLER_67_2212 ();
 sg13g2_decap_8 FILLER_67_2219 ();
 sg13g2_decap_8 FILLER_67_2226 ();
 sg13g2_decap_8 FILLER_67_2233 ();
 sg13g2_decap_8 FILLER_67_2240 ();
 sg13g2_decap_8 FILLER_67_2247 ();
 sg13g2_decap_8 FILLER_67_2254 ();
 sg13g2_decap_8 FILLER_67_2261 ();
 sg13g2_decap_8 FILLER_67_2268 ();
 sg13g2_decap_8 FILLER_67_2275 ();
 sg13g2_decap_8 FILLER_67_2282 ();
 sg13g2_decap_8 FILLER_67_2289 ();
 sg13g2_decap_8 FILLER_67_2296 ();
 sg13g2_decap_8 FILLER_67_2303 ();
 sg13g2_decap_8 FILLER_67_2310 ();
 sg13g2_decap_8 FILLER_67_2317 ();
 sg13g2_decap_8 FILLER_67_2324 ();
 sg13g2_decap_8 FILLER_67_2331 ();
 sg13g2_decap_8 FILLER_67_2338 ();
 sg13g2_decap_8 FILLER_67_2345 ();
 sg13g2_decap_8 FILLER_67_2352 ();
 sg13g2_decap_8 FILLER_67_2359 ();
 sg13g2_decap_8 FILLER_67_2366 ();
 sg13g2_decap_8 FILLER_67_2373 ();
 sg13g2_decap_8 FILLER_67_2380 ();
 sg13g2_decap_8 FILLER_67_2387 ();
 sg13g2_decap_8 FILLER_67_2394 ();
 sg13g2_decap_8 FILLER_67_2401 ();
 sg13g2_decap_8 FILLER_67_2408 ();
 sg13g2_decap_8 FILLER_67_2415 ();
 sg13g2_decap_8 FILLER_67_2422 ();
 sg13g2_decap_8 FILLER_67_2429 ();
 sg13g2_decap_8 FILLER_67_2436 ();
 sg13g2_decap_8 FILLER_67_2443 ();
 sg13g2_decap_8 FILLER_67_2450 ();
 sg13g2_decap_8 FILLER_67_2457 ();
 sg13g2_decap_8 FILLER_67_2464 ();
 sg13g2_decap_8 FILLER_67_2471 ();
 sg13g2_decap_8 FILLER_67_2478 ();
 sg13g2_decap_8 FILLER_67_2485 ();
 sg13g2_decap_8 FILLER_67_2492 ();
 sg13g2_decap_8 FILLER_67_2499 ();
 sg13g2_decap_8 FILLER_67_2506 ();
 sg13g2_decap_8 FILLER_67_2513 ();
 sg13g2_decap_8 FILLER_67_2520 ();
 sg13g2_decap_8 FILLER_67_2527 ();
 sg13g2_decap_8 FILLER_67_2534 ();
 sg13g2_decap_8 FILLER_67_2541 ();
 sg13g2_decap_8 FILLER_67_2548 ();
 sg13g2_decap_8 FILLER_67_2555 ();
 sg13g2_decap_8 FILLER_67_2562 ();
 sg13g2_decap_8 FILLER_67_2569 ();
 sg13g2_decap_8 FILLER_67_2576 ();
 sg13g2_decap_8 FILLER_67_2583 ();
 sg13g2_decap_8 FILLER_67_2590 ();
 sg13g2_decap_8 FILLER_67_2597 ();
 sg13g2_decap_8 FILLER_67_2604 ();
 sg13g2_decap_8 FILLER_67_2611 ();
 sg13g2_decap_8 FILLER_67_2618 ();
 sg13g2_decap_8 FILLER_67_2625 ();
 sg13g2_decap_8 FILLER_67_2632 ();
 sg13g2_decap_8 FILLER_67_2639 ();
 sg13g2_decap_8 FILLER_67_2646 ();
 sg13g2_decap_8 FILLER_67_2653 ();
 sg13g2_decap_8 FILLER_67_2660 ();
 sg13g2_decap_8 FILLER_67_2667 ();
 sg13g2_decap_8 FILLER_67_2674 ();
 sg13g2_decap_8 FILLER_67_2681 ();
 sg13g2_decap_8 FILLER_67_2688 ();
 sg13g2_decap_8 FILLER_67_2695 ();
 sg13g2_decap_8 FILLER_67_2702 ();
 sg13g2_decap_8 FILLER_67_2709 ();
 sg13g2_decap_8 FILLER_67_2716 ();
 sg13g2_decap_8 FILLER_67_2723 ();
 sg13g2_decap_8 FILLER_67_2730 ();
 sg13g2_decap_8 FILLER_67_2737 ();
 sg13g2_decap_8 FILLER_67_2744 ();
 sg13g2_decap_8 FILLER_67_2751 ();
 sg13g2_decap_8 FILLER_67_2758 ();
 sg13g2_decap_8 FILLER_67_2765 ();
 sg13g2_decap_8 FILLER_67_2772 ();
 sg13g2_decap_8 FILLER_67_2779 ();
 sg13g2_decap_8 FILLER_67_2786 ();
 sg13g2_decap_8 FILLER_67_2793 ();
 sg13g2_decap_8 FILLER_67_2800 ();
 sg13g2_decap_8 FILLER_67_2807 ();
 sg13g2_decap_8 FILLER_67_2814 ();
 sg13g2_decap_8 FILLER_67_2821 ();
 sg13g2_decap_8 FILLER_67_2828 ();
 sg13g2_decap_8 FILLER_67_2835 ();
 sg13g2_decap_8 FILLER_67_2842 ();
 sg13g2_decap_8 FILLER_67_2849 ();
 sg13g2_decap_8 FILLER_67_2856 ();
 sg13g2_decap_8 FILLER_67_2863 ();
 sg13g2_decap_8 FILLER_67_2870 ();
 sg13g2_decap_8 FILLER_67_2877 ();
 sg13g2_decap_8 FILLER_67_2884 ();
 sg13g2_decap_8 FILLER_67_2891 ();
 sg13g2_decap_8 FILLER_67_2898 ();
 sg13g2_decap_8 FILLER_67_2905 ();
 sg13g2_decap_8 FILLER_67_2912 ();
 sg13g2_decap_8 FILLER_67_2919 ();
 sg13g2_decap_8 FILLER_67_2926 ();
 sg13g2_decap_8 FILLER_67_2933 ();
 sg13g2_decap_8 FILLER_67_2940 ();
 sg13g2_decap_8 FILLER_67_2947 ();
 sg13g2_decap_8 FILLER_67_2954 ();
 sg13g2_decap_8 FILLER_67_2961 ();
 sg13g2_decap_8 FILLER_67_2968 ();
 sg13g2_decap_8 FILLER_67_2975 ();
 sg13g2_decap_8 FILLER_67_2982 ();
 sg13g2_decap_8 FILLER_67_2989 ();
 sg13g2_decap_8 FILLER_67_2996 ();
 sg13g2_decap_8 FILLER_67_3003 ();
 sg13g2_decap_8 FILLER_67_3010 ();
 sg13g2_decap_8 FILLER_67_3017 ();
 sg13g2_decap_8 FILLER_67_3024 ();
 sg13g2_decap_8 FILLER_67_3031 ();
 sg13g2_decap_8 FILLER_67_3038 ();
 sg13g2_decap_8 FILLER_67_3045 ();
 sg13g2_decap_8 FILLER_67_3052 ();
 sg13g2_decap_8 FILLER_67_3059 ();
 sg13g2_decap_8 FILLER_67_3066 ();
 sg13g2_decap_8 FILLER_67_3073 ();
 sg13g2_decap_8 FILLER_67_3080 ();
 sg13g2_decap_8 FILLER_67_3087 ();
 sg13g2_decap_8 FILLER_67_3094 ();
 sg13g2_decap_8 FILLER_67_3101 ();
 sg13g2_decap_8 FILLER_67_3108 ();
 sg13g2_decap_8 FILLER_67_3115 ();
 sg13g2_decap_8 FILLER_67_3122 ();
 sg13g2_decap_8 FILLER_67_3129 ();
 sg13g2_decap_8 FILLER_67_3136 ();
 sg13g2_decap_8 FILLER_67_3143 ();
 sg13g2_decap_8 FILLER_67_3150 ();
 sg13g2_decap_8 FILLER_67_3157 ();
 sg13g2_decap_8 FILLER_67_3164 ();
 sg13g2_decap_8 FILLER_67_3171 ();
 sg13g2_decap_8 FILLER_67_3178 ();
 sg13g2_decap_8 FILLER_67_3185 ();
 sg13g2_decap_8 FILLER_67_3192 ();
 sg13g2_decap_8 FILLER_67_3199 ();
 sg13g2_decap_8 FILLER_67_3206 ();
 sg13g2_decap_8 FILLER_67_3213 ();
 sg13g2_decap_8 FILLER_67_3220 ();
 sg13g2_decap_8 FILLER_67_3227 ();
 sg13g2_decap_8 FILLER_67_3234 ();
 sg13g2_decap_8 FILLER_67_3241 ();
 sg13g2_decap_8 FILLER_67_3248 ();
 sg13g2_decap_8 FILLER_67_3255 ();
 sg13g2_decap_8 FILLER_67_3262 ();
 sg13g2_decap_8 FILLER_67_3269 ();
 sg13g2_decap_8 FILLER_67_3276 ();
 sg13g2_decap_8 FILLER_67_3283 ();
 sg13g2_decap_8 FILLER_67_3290 ();
 sg13g2_decap_8 FILLER_67_3297 ();
 sg13g2_decap_8 FILLER_67_3304 ();
 sg13g2_decap_8 FILLER_67_3311 ();
 sg13g2_decap_8 FILLER_67_3318 ();
 sg13g2_decap_8 FILLER_67_3325 ();
 sg13g2_decap_8 FILLER_67_3332 ();
 sg13g2_decap_8 FILLER_67_3339 ();
 sg13g2_decap_8 FILLER_67_3346 ();
 sg13g2_decap_8 FILLER_67_3353 ();
 sg13g2_decap_8 FILLER_67_3360 ();
 sg13g2_decap_8 FILLER_67_3367 ();
 sg13g2_decap_8 FILLER_67_3374 ();
 sg13g2_decap_8 FILLER_67_3381 ();
 sg13g2_decap_8 FILLER_67_3388 ();
 sg13g2_decap_8 FILLER_67_3395 ();
 sg13g2_decap_8 FILLER_67_3402 ();
 sg13g2_decap_8 FILLER_67_3409 ();
 sg13g2_decap_8 FILLER_67_3416 ();
 sg13g2_decap_8 FILLER_67_3423 ();
 sg13g2_decap_8 FILLER_67_3430 ();
 sg13g2_decap_8 FILLER_67_3437 ();
 sg13g2_decap_8 FILLER_67_3444 ();
 sg13g2_decap_8 FILLER_67_3451 ();
 sg13g2_decap_8 FILLER_67_3458 ();
 sg13g2_decap_8 FILLER_67_3465 ();
 sg13g2_decap_8 FILLER_67_3472 ();
 sg13g2_decap_8 FILLER_67_3479 ();
 sg13g2_decap_8 FILLER_67_3486 ();
 sg13g2_decap_8 FILLER_67_3493 ();
 sg13g2_decap_8 FILLER_67_3500 ();
 sg13g2_decap_8 FILLER_67_3507 ();
 sg13g2_decap_8 FILLER_67_3514 ();
 sg13g2_decap_8 FILLER_67_3521 ();
 sg13g2_decap_8 FILLER_67_3528 ();
 sg13g2_decap_8 FILLER_67_3535 ();
 sg13g2_decap_8 FILLER_67_3542 ();
 sg13g2_decap_8 FILLER_67_3549 ();
 sg13g2_decap_8 FILLER_67_3556 ();
 sg13g2_decap_8 FILLER_67_3563 ();
 sg13g2_decap_8 FILLER_67_3570 ();
 sg13g2_fill_2 FILLER_67_3577 ();
 sg13g2_fill_1 FILLER_67_3579 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_decap_8 FILLER_68_119 ();
 sg13g2_decap_8 FILLER_68_126 ();
 sg13g2_decap_8 FILLER_68_133 ();
 sg13g2_decap_8 FILLER_68_140 ();
 sg13g2_decap_8 FILLER_68_147 ();
 sg13g2_decap_8 FILLER_68_154 ();
 sg13g2_decap_8 FILLER_68_161 ();
 sg13g2_decap_8 FILLER_68_168 ();
 sg13g2_decap_8 FILLER_68_175 ();
 sg13g2_decap_8 FILLER_68_182 ();
 sg13g2_decap_8 FILLER_68_189 ();
 sg13g2_decap_8 FILLER_68_196 ();
 sg13g2_decap_8 FILLER_68_203 ();
 sg13g2_decap_8 FILLER_68_210 ();
 sg13g2_fill_1 FILLER_68_217 ();
 sg13g2_decap_8 FILLER_68_222 ();
 sg13g2_decap_8 FILLER_68_229 ();
 sg13g2_decap_8 FILLER_68_236 ();
 sg13g2_decap_8 FILLER_68_243 ();
 sg13g2_decap_8 FILLER_68_250 ();
 sg13g2_decap_8 FILLER_68_257 ();
 sg13g2_decap_8 FILLER_68_264 ();
 sg13g2_decap_8 FILLER_68_271 ();
 sg13g2_decap_8 FILLER_68_278 ();
 sg13g2_decap_8 FILLER_68_285 ();
 sg13g2_decap_8 FILLER_68_292 ();
 sg13g2_decap_8 FILLER_68_299 ();
 sg13g2_decap_8 FILLER_68_306 ();
 sg13g2_decap_8 FILLER_68_313 ();
 sg13g2_decap_8 FILLER_68_320 ();
 sg13g2_decap_8 FILLER_68_327 ();
 sg13g2_decap_8 FILLER_68_334 ();
 sg13g2_decap_8 FILLER_68_341 ();
 sg13g2_decap_8 FILLER_68_348 ();
 sg13g2_decap_8 FILLER_68_355 ();
 sg13g2_decap_8 FILLER_68_362 ();
 sg13g2_decap_8 FILLER_68_369 ();
 sg13g2_decap_8 FILLER_68_376 ();
 sg13g2_decap_8 FILLER_68_383 ();
 sg13g2_decap_8 FILLER_68_390 ();
 sg13g2_decap_8 FILLER_68_397 ();
 sg13g2_decap_8 FILLER_68_404 ();
 sg13g2_decap_8 FILLER_68_411 ();
 sg13g2_decap_8 FILLER_68_418 ();
 sg13g2_decap_8 FILLER_68_425 ();
 sg13g2_decap_8 FILLER_68_432 ();
 sg13g2_decap_8 FILLER_68_439 ();
 sg13g2_decap_8 FILLER_68_446 ();
 sg13g2_decap_8 FILLER_68_453 ();
 sg13g2_decap_8 FILLER_68_460 ();
 sg13g2_decap_8 FILLER_68_467 ();
 sg13g2_decap_8 FILLER_68_474 ();
 sg13g2_decap_8 FILLER_68_481 ();
 sg13g2_decap_8 FILLER_68_488 ();
 sg13g2_decap_8 FILLER_68_495 ();
 sg13g2_decap_8 FILLER_68_502 ();
 sg13g2_decap_8 FILLER_68_509 ();
 sg13g2_decap_8 FILLER_68_516 ();
 sg13g2_decap_8 FILLER_68_523 ();
 sg13g2_decap_8 FILLER_68_530 ();
 sg13g2_decap_8 FILLER_68_537 ();
 sg13g2_decap_8 FILLER_68_544 ();
 sg13g2_decap_8 FILLER_68_551 ();
 sg13g2_decap_8 FILLER_68_558 ();
 sg13g2_decap_8 FILLER_68_565 ();
 sg13g2_decap_8 FILLER_68_572 ();
 sg13g2_decap_8 FILLER_68_579 ();
 sg13g2_decap_8 FILLER_68_586 ();
 sg13g2_decap_8 FILLER_68_593 ();
 sg13g2_decap_8 FILLER_68_600 ();
 sg13g2_decap_8 FILLER_68_607 ();
 sg13g2_decap_8 FILLER_68_614 ();
 sg13g2_decap_8 FILLER_68_621 ();
 sg13g2_decap_8 FILLER_68_628 ();
 sg13g2_decap_8 FILLER_68_635 ();
 sg13g2_decap_8 FILLER_68_642 ();
 sg13g2_decap_8 FILLER_68_649 ();
 sg13g2_decap_8 FILLER_68_656 ();
 sg13g2_decap_8 FILLER_68_663 ();
 sg13g2_decap_8 FILLER_68_670 ();
 sg13g2_decap_8 FILLER_68_677 ();
 sg13g2_decap_8 FILLER_68_684 ();
 sg13g2_decap_8 FILLER_68_691 ();
 sg13g2_decap_8 FILLER_68_698 ();
 sg13g2_decap_8 FILLER_68_705 ();
 sg13g2_decap_8 FILLER_68_712 ();
 sg13g2_decap_8 FILLER_68_719 ();
 sg13g2_decap_8 FILLER_68_726 ();
 sg13g2_decap_8 FILLER_68_733 ();
 sg13g2_decap_8 FILLER_68_740 ();
 sg13g2_decap_8 FILLER_68_747 ();
 sg13g2_decap_8 FILLER_68_754 ();
 sg13g2_decap_8 FILLER_68_761 ();
 sg13g2_decap_8 FILLER_68_768 ();
 sg13g2_decap_8 FILLER_68_775 ();
 sg13g2_decap_8 FILLER_68_782 ();
 sg13g2_decap_8 FILLER_68_789 ();
 sg13g2_decap_8 FILLER_68_796 ();
 sg13g2_decap_8 FILLER_68_803 ();
 sg13g2_decap_8 FILLER_68_810 ();
 sg13g2_decap_8 FILLER_68_817 ();
 sg13g2_decap_8 FILLER_68_824 ();
 sg13g2_decap_8 FILLER_68_831 ();
 sg13g2_decap_8 FILLER_68_838 ();
 sg13g2_decap_8 FILLER_68_845 ();
 sg13g2_decap_8 FILLER_68_852 ();
 sg13g2_decap_8 FILLER_68_859 ();
 sg13g2_decap_8 FILLER_68_866 ();
 sg13g2_decap_8 FILLER_68_873 ();
 sg13g2_decap_8 FILLER_68_880 ();
 sg13g2_decap_8 FILLER_68_887 ();
 sg13g2_decap_8 FILLER_68_894 ();
 sg13g2_decap_8 FILLER_68_901 ();
 sg13g2_decap_8 FILLER_68_908 ();
 sg13g2_decap_8 FILLER_68_915 ();
 sg13g2_decap_8 FILLER_68_922 ();
 sg13g2_decap_8 FILLER_68_929 ();
 sg13g2_decap_8 FILLER_68_936 ();
 sg13g2_decap_8 FILLER_68_943 ();
 sg13g2_decap_8 FILLER_68_950 ();
 sg13g2_decap_8 FILLER_68_957 ();
 sg13g2_decap_8 FILLER_68_964 ();
 sg13g2_decap_8 FILLER_68_971 ();
 sg13g2_decap_8 FILLER_68_978 ();
 sg13g2_decap_8 FILLER_68_985 ();
 sg13g2_decap_8 FILLER_68_992 ();
 sg13g2_decap_8 FILLER_68_999 ();
 sg13g2_decap_8 FILLER_68_1006 ();
 sg13g2_decap_8 FILLER_68_1013 ();
 sg13g2_decap_8 FILLER_68_1020 ();
 sg13g2_decap_8 FILLER_68_1027 ();
 sg13g2_decap_8 FILLER_68_1034 ();
 sg13g2_decap_8 FILLER_68_1041 ();
 sg13g2_decap_8 FILLER_68_1048 ();
 sg13g2_decap_8 FILLER_68_1055 ();
 sg13g2_decap_8 FILLER_68_1062 ();
 sg13g2_decap_8 FILLER_68_1069 ();
 sg13g2_decap_8 FILLER_68_1076 ();
 sg13g2_decap_8 FILLER_68_1083 ();
 sg13g2_decap_8 FILLER_68_1090 ();
 sg13g2_decap_8 FILLER_68_1097 ();
 sg13g2_decap_8 FILLER_68_1104 ();
 sg13g2_decap_8 FILLER_68_1111 ();
 sg13g2_decap_8 FILLER_68_1118 ();
 sg13g2_decap_8 FILLER_68_1125 ();
 sg13g2_decap_8 FILLER_68_1132 ();
 sg13g2_decap_8 FILLER_68_1139 ();
 sg13g2_decap_8 FILLER_68_1146 ();
 sg13g2_decap_8 FILLER_68_1153 ();
 sg13g2_decap_8 FILLER_68_1160 ();
 sg13g2_decap_8 FILLER_68_1167 ();
 sg13g2_decap_8 FILLER_68_1174 ();
 sg13g2_decap_8 FILLER_68_1181 ();
 sg13g2_decap_8 FILLER_68_1188 ();
 sg13g2_decap_8 FILLER_68_1195 ();
 sg13g2_decap_8 FILLER_68_1202 ();
 sg13g2_decap_8 FILLER_68_1209 ();
 sg13g2_decap_8 FILLER_68_1216 ();
 sg13g2_decap_8 FILLER_68_1223 ();
 sg13g2_decap_8 FILLER_68_1230 ();
 sg13g2_decap_8 FILLER_68_1237 ();
 sg13g2_decap_8 FILLER_68_1244 ();
 sg13g2_decap_8 FILLER_68_1251 ();
 sg13g2_decap_8 FILLER_68_1258 ();
 sg13g2_decap_8 FILLER_68_1265 ();
 sg13g2_decap_8 FILLER_68_1272 ();
 sg13g2_decap_8 FILLER_68_1279 ();
 sg13g2_decap_8 FILLER_68_1286 ();
 sg13g2_decap_8 FILLER_68_1293 ();
 sg13g2_decap_8 FILLER_68_1300 ();
 sg13g2_decap_8 FILLER_68_1307 ();
 sg13g2_decap_8 FILLER_68_1314 ();
 sg13g2_decap_8 FILLER_68_1321 ();
 sg13g2_decap_8 FILLER_68_1328 ();
 sg13g2_decap_8 FILLER_68_1335 ();
 sg13g2_decap_8 FILLER_68_1342 ();
 sg13g2_decap_8 FILLER_68_1349 ();
 sg13g2_decap_8 FILLER_68_1356 ();
 sg13g2_decap_8 FILLER_68_1363 ();
 sg13g2_decap_8 FILLER_68_1370 ();
 sg13g2_decap_8 FILLER_68_1377 ();
 sg13g2_decap_8 FILLER_68_1384 ();
 sg13g2_decap_8 FILLER_68_1391 ();
 sg13g2_decap_8 FILLER_68_1398 ();
 sg13g2_decap_8 FILLER_68_1405 ();
 sg13g2_decap_8 FILLER_68_1412 ();
 sg13g2_decap_8 FILLER_68_1419 ();
 sg13g2_decap_8 FILLER_68_1426 ();
 sg13g2_decap_8 FILLER_68_1433 ();
 sg13g2_decap_8 FILLER_68_1440 ();
 sg13g2_decap_8 FILLER_68_1447 ();
 sg13g2_decap_8 FILLER_68_1454 ();
 sg13g2_decap_8 FILLER_68_1461 ();
 sg13g2_decap_8 FILLER_68_1468 ();
 sg13g2_decap_8 FILLER_68_1475 ();
 sg13g2_decap_8 FILLER_68_1482 ();
 sg13g2_decap_8 FILLER_68_1489 ();
 sg13g2_decap_8 FILLER_68_1496 ();
 sg13g2_decap_8 FILLER_68_1503 ();
 sg13g2_decap_8 FILLER_68_1510 ();
 sg13g2_decap_8 FILLER_68_1517 ();
 sg13g2_decap_8 FILLER_68_1524 ();
 sg13g2_decap_8 FILLER_68_1531 ();
 sg13g2_decap_8 FILLER_68_1538 ();
 sg13g2_decap_8 FILLER_68_1545 ();
 sg13g2_decap_8 FILLER_68_1552 ();
 sg13g2_decap_8 FILLER_68_1559 ();
 sg13g2_decap_8 FILLER_68_1566 ();
 sg13g2_decap_8 FILLER_68_1573 ();
 sg13g2_decap_8 FILLER_68_1580 ();
 sg13g2_decap_8 FILLER_68_1587 ();
 sg13g2_decap_8 FILLER_68_1594 ();
 sg13g2_decap_8 FILLER_68_1601 ();
 sg13g2_decap_8 FILLER_68_1608 ();
 sg13g2_decap_8 FILLER_68_1615 ();
 sg13g2_decap_8 FILLER_68_1622 ();
 sg13g2_decap_8 FILLER_68_1629 ();
 sg13g2_decap_8 FILLER_68_1636 ();
 sg13g2_decap_8 FILLER_68_1643 ();
 sg13g2_decap_8 FILLER_68_1650 ();
 sg13g2_decap_8 FILLER_68_1657 ();
 sg13g2_decap_8 FILLER_68_1664 ();
 sg13g2_decap_8 FILLER_68_1671 ();
 sg13g2_decap_8 FILLER_68_1678 ();
 sg13g2_decap_8 FILLER_68_1685 ();
 sg13g2_decap_8 FILLER_68_1692 ();
 sg13g2_decap_8 FILLER_68_1699 ();
 sg13g2_decap_8 FILLER_68_1706 ();
 sg13g2_decap_8 FILLER_68_1713 ();
 sg13g2_decap_8 FILLER_68_1720 ();
 sg13g2_decap_8 FILLER_68_1727 ();
 sg13g2_decap_8 FILLER_68_1734 ();
 sg13g2_decap_8 FILLER_68_1741 ();
 sg13g2_decap_8 FILLER_68_1748 ();
 sg13g2_decap_8 FILLER_68_1755 ();
 sg13g2_decap_8 FILLER_68_1762 ();
 sg13g2_decap_8 FILLER_68_1769 ();
 sg13g2_decap_8 FILLER_68_1776 ();
 sg13g2_decap_8 FILLER_68_1783 ();
 sg13g2_decap_8 FILLER_68_1790 ();
 sg13g2_decap_8 FILLER_68_1797 ();
 sg13g2_decap_8 FILLER_68_1804 ();
 sg13g2_decap_8 FILLER_68_1811 ();
 sg13g2_decap_8 FILLER_68_1818 ();
 sg13g2_decap_8 FILLER_68_1825 ();
 sg13g2_decap_8 FILLER_68_1832 ();
 sg13g2_decap_8 FILLER_68_1839 ();
 sg13g2_decap_8 FILLER_68_1846 ();
 sg13g2_decap_8 FILLER_68_1853 ();
 sg13g2_decap_8 FILLER_68_1860 ();
 sg13g2_decap_8 FILLER_68_1867 ();
 sg13g2_decap_8 FILLER_68_1874 ();
 sg13g2_decap_8 FILLER_68_1881 ();
 sg13g2_decap_8 FILLER_68_1888 ();
 sg13g2_decap_8 FILLER_68_1895 ();
 sg13g2_decap_8 FILLER_68_1902 ();
 sg13g2_decap_8 FILLER_68_1909 ();
 sg13g2_decap_8 FILLER_68_1916 ();
 sg13g2_decap_8 FILLER_68_1923 ();
 sg13g2_decap_8 FILLER_68_1930 ();
 sg13g2_decap_8 FILLER_68_1937 ();
 sg13g2_decap_8 FILLER_68_1944 ();
 sg13g2_decap_8 FILLER_68_1951 ();
 sg13g2_decap_8 FILLER_68_1958 ();
 sg13g2_decap_8 FILLER_68_1965 ();
 sg13g2_decap_8 FILLER_68_1972 ();
 sg13g2_decap_8 FILLER_68_1979 ();
 sg13g2_decap_8 FILLER_68_1986 ();
 sg13g2_decap_8 FILLER_68_1993 ();
 sg13g2_decap_8 FILLER_68_2000 ();
 sg13g2_decap_8 FILLER_68_2007 ();
 sg13g2_decap_8 FILLER_68_2014 ();
 sg13g2_decap_8 FILLER_68_2021 ();
 sg13g2_decap_8 FILLER_68_2028 ();
 sg13g2_decap_8 FILLER_68_2035 ();
 sg13g2_decap_8 FILLER_68_2042 ();
 sg13g2_decap_8 FILLER_68_2049 ();
 sg13g2_decap_8 FILLER_68_2056 ();
 sg13g2_decap_8 FILLER_68_2063 ();
 sg13g2_decap_8 FILLER_68_2070 ();
 sg13g2_decap_8 FILLER_68_2077 ();
 sg13g2_decap_8 FILLER_68_2084 ();
 sg13g2_decap_8 FILLER_68_2091 ();
 sg13g2_decap_8 FILLER_68_2098 ();
 sg13g2_decap_8 FILLER_68_2105 ();
 sg13g2_decap_8 FILLER_68_2112 ();
 sg13g2_decap_8 FILLER_68_2119 ();
 sg13g2_decap_8 FILLER_68_2126 ();
 sg13g2_decap_8 FILLER_68_2133 ();
 sg13g2_decap_8 FILLER_68_2140 ();
 sg13g2_decap_8 FILLER_68_2147 ();
 sg13g2_decap_8 FILLER_68_2154 ();
 sg13g2_decap_8 FILLER_68_2161 ();
 sg13g2_decap_8 FILLER_68_2168 ();
 sg13g2_decap_8 FILLER_68_2175 ();
 sg13g2_decap_8 FILLER_68_2182 ();
 sg13g2_decap_8 FILLER_68_2189 ();
 sg13g2_decap_8 FILLER_68_2196 ();
 sg13g2_decap_8 FILLER_68_2203 ();
 sg13g2_decap_8 FILLER_68_2210 ();
 sg13g2_decap_8 FILLER_68_2217 ();
 sg13g2_decap_8 FILLER_68_2224 ();
 sg13g2_decap_8 FILLER_68_2231 ();
 sg13g2_decap_8 FILLER_68_2238 ();
 sg13g2_decap_8 FILLER_68_2245 ();
 sg13g2_decap_8 FILLER_68_2252 ();
 sg13g2_decap_8 FILLER_68_2259 ();
 sg13g2_decap_8 FILLER_68_2266 ();
 sg13g2_decap_8 FILLER_68_2273 ();
 sg13g2_decap_8 FILLER_68_2280 ();
 sg13g2_decap_8 FILLER_68_2287 ();
 sg13g2_decap_8 FILLER_68_2294 ();
 sg13g2_decap_8 FILLER_68_2301 ();
 sg13g2_decap_8 FILLER_68_2308 ();
 sg13g2_decap_8 FILLER_68_2315 ();
 sg13g2_decap_8 FILLER_68_2322 ();
 sg13g2_decap_8 FILLER_68_2329 ();
 sg13g2_decap_8 FILLER_68_2336 ();
 sg13g2_decap_8 FILLER_68_2343 ();
 sg13g2_decap_8 FILLER_68_2350 ();
 sg13g2_decap_8 FILLER_68_2357 ();
 sg13g2_decap_8 FILLER_68_2364 ();
 sg13g2_decap_8 FILLER_68_2371 ();
 sg13g2_decap_8 FILLER_68_2378 ();
 sg13g2_decap_8 FILLER_68_2385 ();
 sg13g2_decap_8 FILLER_68_2392 ();
 sg13g2_decap_8 FILLER_68_2399 ();
 sg13g2_decap_8 FILLER_68_2406 ();
 sg13g2_decap_8 FILLER_68_2413 ();
 sg13g2_decap_8 FILLER_68_2420 ();
 sg13g2_decap_8 FILLER_68_2427 ();
 sg13g2_decap_8 FILLER_68_2434 ();
 sg13g2_decap_8 FILLER_68_2441 ();
 sg13g2_decap_8 FILLER_68_2448 ();
 sg13g2_decap_8 FILLER_68_2455 ();
 sg13g2_decap_8 FILLER_68_2462 ();
 sg13g2_decap_8 FILLER_68_2469 ();
 sg13g2_decap_8 FILLER_68_2476 ();
 sg13g2_decap_8 FILLER_68_2483 ();
 sg13g2_decap_8 FILLER_68_2490 ();
 sg13g2_decap_8 FILLER_68_2497 ();
 sg13g2_decap_8 FILLER_68_2504 ();
 sg13g2_decap_8 FILLER_68_2511 ();
 sg13g2_decap_8 FILLER_68_2518 ();
 sg13g2_decap_8 FILLER_68_2525 ();
 sg13g2_decap_8 FILLER_68_2532 ();
 sg13g2_decap_8 FILLER_68_2539 ();
 sg13g2_decap_8 FILLER_68_2546 ();
 sg13g2_decap_8 FILLER_68_2553 ();
 sg13g2_decap_8 FILLER_68_2560 ();
 sg13g2_decap_8 FILLER_68_2567 ();
 sg13g2_decap_8 FILLER_68_2574 ();
 sg13g2_decap_8 FILLER_68_2581 ();
 sg13g2_decap_8 FILLER_68_2588 ();
 sg13g2_decap_8 FILLER_68_2595 ();
 sg13g2_decap_8 FILLER_68_2602 ();
 sg13g2_decap_8 FILLER_68_2609 ();
 sg13g2_decap_8 FILLER_68_2616 ();
 sg13g2_decap_8 FILLER_68_2623 ();
 sg13g2_decap_8 FILLER_68_2630 ();
 sg13g2_decap_8 FILLER_68_2637 ();
 sg13g2_decap_8 FILLER_68_2644 ();
 sg13g2_decap_8 FILLER_68_2651 ();
 sg13g2_decap_8 FILLER_68_2658 ();
 sg13g2_decap_8 FILLER_68_2665 ();
 sg13g2_decap_8 FILLER_68_2672 ();
 sg13g2_decap_8 FILLER_68_2679 ();
 sg13g2_decap_8 FILLER_68_2686 ();
 sg13g2_decap_8 FILLER_68_2693 ();
 sg13g2_decap_8 FILLER_68_2700 ();
 sg13g2_decap_8 FILLER_68_2707 ();
 sg13g2_decap_8 FILLER_68_2714 ();
 sg13g2_decap_8 FILLER_68_2721 ();
 sg13g2_decap_8 FILLER_68_2728 ();
 sg13g2_decap_8 FILLER_68_2735 ();
 sg13g2_decap_8 FILLER_68_2742 ();
 sg13g2_decap_8 FILLER_68_2749 ();
 sg13g2_decap_8 FILLER_68_2756 ();
 sg13g2_decap_8 FILLER_68_2763 ();
 sg13g2_decap_8 FILLER_68_2770 ();
 sg13g2_decap_8 FILLER_68_2777 ();
 sg13g2_decap_8 FILLER_68_2784 ();
 sg13g2_decap_8 FILLER_68_2791 ();
 sg13g2_decap_8 FILLER_68_2798 ();
 sg13g2_decap_8 FILLER_68_2805 ();
 sg13g2_decap_8 FILLER_68_2812 ();
 sg13g2_decap_8 FILLER_68_2819 ();
 sg13g2_decap_8 FILLER_68_2826 ();
 sg13g2_decap_8 FILLER_68_2833 ();
 sg13g2_decap_8 FILLER_68_2840 ();
 sg13g2_decap_8 FILLER_68_2847 ();
 sg13g2_decap_8 FILLER_68_2854 ();
 sg13g2_decap_8 FILLER_68_2861 ();
 sg13g2_decap_8 FILLER_68_2868 ();
 sg13g2_decap_8 FILLER_68_2875 ();
 sg13g2_decap_8 FILLER_68_2882 ();
 sg13g2_decap_8 FILLER_68_2889 ();
 sg13g2_decap_8 FILLER_68_2896 ();
 sg13g2_decap_8 FILLER_68_2903 ();
 sg13g2_decap_8 FILLER_68_2910 ();
 sg13g2_decap_8 FILLER_68_2917 ();
 sg13g2_decap_8 FILLER_68_2924 ();
 sg13g2_decap_8 FILLER_68_2931 ();
 sg13g2_decap_8 FILLER_68_2938 ();
 sg13g2_decap_8 FILLER_68_2945 ();
 sg13g2_decap_8 FILLER_68_2952 ();
 sg13g2_decap_8 FILLER_68_2959 ();
 sg13g2_decap_8 FILLER_68_2966 ();
 sg13g2_decap_8 FILLER_68_2973 ();
 sg13g2_decap_8 FILLER_68_2980 ();
 sg13g2_decap_8 FILLER_68_2987 ();
 sg13g2_decap_8 FILLER_68_2994 ();
 sg13g2_decap_8 FILLER_68_3001 ();
 sg13g2_decap_8 FILLER_68_3008 ();
 sg13g2_decap_8 FILLER_68_3015 ();
 sg13g2_decap_8 FILLER_68_3022 ();
 sg13g2_decap_8 FILLER_68_3029 ();
 sg13g2_decap_8 FILLER_68_3036 ();
 sg13g2_decap_8 FILLER_68_3043 ();
 sg13g2_decap_8 FILLER_68_3050 ();
 sg13g2_decap_8 FILLER_68_3057 ();
 sg13g2_decap_8 FILLER_68_3064 ();
 sg13g2_decap_8 FILLER_68_3071 ();
 sg13g2_decap_8 FILLER_68_3078 ();
 sg13g2_decap_8 FILLER_68_3085 ();
 sg13g2_decap_8 FILLER_68_3092 ();
 sg13g2_decap_8 FILLER_68_3099 ();
 sg13g2_decap_8 FILLER_68_3106 ();
 sg13g2_decap_8 FILLER_68_3113 ();
 sg13g2_decap_8 FILLER_68_3120 ();
 sg13g2_decap_8 FILLER_68_3127 ();
 sg13g2_decap_8 FILLER_68_3134 ();
 sg13g2_decap_8 FILLER_68_3141 ();
 sg13g2_decap_8 FILLER_68_3148 ();
 sg13g2_decap_8 FILLER_68_3155 ();
 sg13g2_decap_8 FILLER_68_3162 ();
 sg13g2_decap_8 FILLER_68_3169 ();
 sg13g2_decap_8 FILLER_68_3176 ();
 sg13g2_decap_8 FILLER_68_3183 ();
 sg13g2_decap_8 FILLER_68_3190 ();
 sg13g2_decap_8 FILLER_68_3197 ();
 sg13g2_decap_8 FILLER_68_3204 ();
 sg13g2_decap_8 FILLER_68_3211 ();
 sg13g2_decap_8 FILLER_68_3218 ();
 sg13g2_decap_8 FILLER_68_3225 ();
 sg13g2_decap_8 FILLER_68_3232 ();
 sg13g2_decap_8 FILLER_68_3239 ();
 sg13g2_decap_8 FILLER_68_3246 ();
 sg13g2_decap_8 FILLER_68_3253 ();
 sg13g2_decap_8 FILLER_68_3260 ();
 sg13g2_decap_8 FILLER_68_3267 ();
 sg13g2_decap_8 FILLER_68_3274 ();
 sg13g2_decap_8 FILLER_68_3281 ();
 sg13g2_decap_8 FILLER_68_3288 ();
 sg13g2_decap_8 FILLER_68_3295 ();
 sg13g2_decap_8 FILLER_68_3302 ();
 sg13g2_decap_8 FILLER_68_3309 ();
 sg13g2_decap_8 FILLER_68_3316 ();
 sg13g2_decap_8 FILLER_68_3323 ();
 sg13g2_decap_8 FILLER_68_3330 ();
 sg13g2_decap_8 FILLER_68_3337 ();
 sg13g2_decap_8 FILLER_68_3344 ();
 sg13g2_decap_8 FILLER_68_3351 ();
 sg13g2_decap_8 FILLER_68_3358 ();
 sg13g2_decap_8 FILLER_68_3365 ();
 sg13g2_decap_8 FILLER_68_3372 ();
 sg13g2_decap_8 FILLER_68_3379 ();
 sg13g2_decap_8 FILLER_68_3386 ();
 sg13g2_decap_8 FILLER_68_3393 ();
 sg13g2_decap_8 FILLER_68_3400 ();
 sg13g2_decap_8 FILLER_68_3407 ();
 sg13g2_decap_8 FILLER_68_3414 ();
 sg13g2_decap_8 FILLER_68_3421 ();
 sg13g2_decap_8 FILLER_68_3428 ();
 sg13g2_decap_8 FILLER_68_3435 ();
 sg13g2_decap_8 FILLER_68_3442 ();
 sg13g2_decap_8 FILLER_68_3449 ();
 sg13g2_decap_8 FILLER_68_3456 ();
 sg13g2_decap_8 FILLER_68_3463 ();
 sg13g2_decap_8 FILLER_68_3470 ();
 sg13g2_decap_8 FILLER_68_3477 ();
 sg13g2_decap_8 FILLER_68_3484 ();
 sg13g2_decap_8 FILLER_68_3491 ();
 sg13g2_decap_8 FILLER_68_3498 ();
 sg13g2_decap_8 FILLER_68_3505 ();
 sg13g2_decap_8 FILLER_68_3512 ();
 sg13g2_decap_8 FILLER_68_3519 ();
 sg13g2_decap_8 FILLER_68_3526 ();
 sg13g2_decap_8 FILLER_68_3533 ();
 sg13g2_decap_8 FILLER_68_3540 ();
 sg13g2_decap_8 FILLER_68_3547 ();
 sg13g2_decap_8 FILLER_68_3554 ();
 sg13g2_decap_8 FILLER_68_3561 ();
 sg13g2_decap_8 FILLER_68_3568 ();
 sg13g2_decap_4 FILLER_68_3575 ();
 sg13g2_fill_1 FILLER_68_3579 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_decap_8 FILLER_69_119 ();
 sg13g2_decap_8 FILLER_69_126 ();
 sg13g2_decap_8 FILLER_69_133 ();
 sg13g2_decap_8 FILLER_69_140 ();
 sg13g2_decap_8 FILLER_69_147 ();
 sg13g2_decap_4 FILLER_69_154 ();
 sg13g2_fill_1 FILLER_69_186 ();
 sg13g2_decap_8 FILLER_69_200 ();
 sg13g2_decap_4 FILLER_69_207 ();
 sg13g2_fill_1 FILLER_69_211 ();
 sg13g2_decap_8 FILLER_69_240 ();
 sg13g2_decap_8 FILLER_69_247 ();
 sg13g2_decap_8 FILLER_69_254 ();
 sg13g2_decap_8 FILLER_69_261 ();
 sg13g2_decap_8 FILLER_69_268 ();
 sg13g2_decap_8 FILLER_69_275 ();
 sg13g2_decap_8 FILLER_69_282 ();
 sg13g2_decap_8 FILLER_69_289 ();
 sg13g2_decap_8 FILLER_69_296 ();
 sg13g2_decap_8 FILLER_69_303 ();
 sg13g2_decap_8 FILLER_69_310 ();
 sg13g2_decap_8 FILLER_69_317 ();
 sg13g2_decap_8 FILLER_69_324 ();
 sg13g2_decap_8 FILLER_69_331 ();
 sg13g2_decap_8 FILLER_69_338 ();
 sg13g2_decap_8 FILLER_69_345 ();
 sg13g2_decap_8 FILLER_69_352 ();
 sg13g2_decap_8 FILLER_69_359 ();
 sg13g2_decap_8 FILLER_69_366 ();
 sg13g2_decap_8 FILLER_69_373 ();
 sg13g2_decap_8 FILLER_69_380 ();
 sg13g2_decap_8 FILLER_69_387 ();
 sg13g2_decap_8 FILLER_69_394 ();
 sg13g2_decap_8 FILLER_69_401 ();
 sg13g2_decap_8 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_69_415 ();
 sg13g2_decap_8 FILLER_69_422 ();
 sg13g2_decap_8 FILLER_69_429 ();
 sg13g2_decap_8 FILLER_69_436 ();
 sg13g2_decap_8 FILLER_69_443 ();
 sg13g2_decap_8 FILLER_69_450 ();
 sg13g2_decap_8 FILLER_69_457 ();
 sg13g2_decap_8 FILLER_69_464 ();
 sg13g2_decap_8 FILLER_69_471 ();
 sg13g2_decap_8 FILLER_69_478 ();
 sg13g2_decap_8 FILLER_69_485 ();
 sg13g2_decap_8 FILLER_69_492 ();
 sg13g2_decap_8 FILLER_69_499 ();
 sg13g2_decap_8 FILLER_69_506 ();
 sg13g2_decap_8 FILLER_69_513 ();
 sg13g2_decap_8 FILLER_69_520 ();
 sg13g2_decap_8 FILLER_69_527 ();
 sg13g2_decap_8 FILLER_69_534 ();
 sg13g2_decap_8 FILLER_69_541 ();
 sg13g2_decap_8 FILLER_69_548 ();
 sg13g2_decap_8 FILLER_69_555 ();
 sg13g2_decap_8 FILLER_69_562 ();
 sg13g2_decap_8 FILLER_69_569 ();
 sg13g2_decap_8 FILLER_69_576 ();
 sg13g2_decap_8 FILLER_69_583 ();
 sg13g2_decap_8 FILLER_69_590 ();
 sg13g2_decap_8 FILLER_69_597 ();
 sg13g2_decap_8 FILLER_69_604 ();
 sg13g2_decap_8 FILLER_69_611 ();
 sg13g2_decap_8 FILLER_69_618 ();
 sg13g2_decap_8 FILLER_69_625 ();
 sg13g2_decap_8 FILLER_69_632 ();
 sg13g2_decap_8 FILLER_69_639 ();
 sg13g2_decap_8 FILLER_69_646 ();
 sg13g2_decap_8 FILLER_69_653 ();
 sg13g2_decap_8 FILLER_69_660 ();
 sg13g2_decap_8 FILLER_69_667 ();
 sg13g2_decap_8 FILLER_69_674 ();
 sg13g2_decap_8 FILLER_69_681 ();
 sg13g2_decap_8 FILLER_69_688 ();
 sg13g2_decap_8 FILLER_69_695 ();
 sg13g2_decap_8 FILLER_69_702 ();
 sg13g2_decap_8 FILLER_69_709 ();
 sg13g2_decap_8 FILLER_69_716 ();
 sg13g2_decap_8 FILLER_69_723 ();
 sg13g2_decap_8 FILLER_69_730 ();
 sg13g2_decap_8 FILLER_69_737 ();
 sg13g2_decap_8 FILLER_69_744 ();
 sg13g2_decap_8 FILLER_69_751 ();
 sg13g2_decap_8 FILLER_69_758 ();
 sg13g2_decap_8 FILLER_69_765 ();
 sg13g2_decap_8 FILLER_69_772 ();
 sg13g2_decap_8 FILLER_69_779 ();
 sg13g2_decap_8 FILLER_69_786 ();
 sg13g2_decap_8 FILLER_69_793 ();
 sg13g2_decap_8 FILLER_69_800 ();
 sg13g2_decap_8 FILLER_69_807 ();
 sg13g2_decap_8 FILLER_69_814 ();
 sg13g2_decap_8 FILLER_69_821 ();
 sg13g2_decap_8 FILLER_69_828 ();
 sg13g2_decap_8 FILLER_69_835 ();
 sg13g2_decap_8 FILLER_69_842 ();
 sg13g2_decap_8 FILLER_69_849 ();
 sg13g2_decap_8 FILLER_69_856 ();
 sg13g2_decap_8 FILLER_69_863 ();
 sg13g2_decap_8 FILLER_69_870 ();
 sg13g2_decap_8 FILLER_69_877 ();
 sg13g2_decap_8 FILLER_69_884 ();
 sg13g2_decap_8 FILLER_69_891 ();
 sg13g2_decap_8 FILLER_69_898 ();
 sg13g2_decap_8 FILLER_69_905 ();
 sg13g2_decap_8 FILLER_69_912 ();
 sg13g2_decap_8 FILLER_69_919 ();
 sg13g2_decap_8 FILLER_69_926 ();
 sg13g2_decap_8 FILLER_69_933 ();
 sg13g2_decap_8 FILLER_69_940 ();
 sg13g2_decap_8 FILLER_69_947 ();
 sg13g2_decap_8 FILLER_69_954 ();
 sg13g2_decap_8 FILLER_69_961 ();
 sg13g2_decap_8 FILLER_69_968 ();
 sg13g2_decap_8 FILLER_69_975 ();
 sg13g2_decap_8 FILLER_69_982 ();
 sg13g2_decap_8 FILLER_69_989 ();
 sg13g2_decap_8 FILLER_69_996 ();
 sg13g2_decap_8 FILLER_69_1003 ();
 sg13g2_decap_8 FILLER_69_1010 ();
 sg13g2_decap_8 FILLER_69_1017 ();
 sg13g2_decap_8 FILLER_69_1024 ();
 sg13g2_decap_8 FILLER_69_1031 ();
 sg13g2_decap_8 FILLER_69_1038 ();
 sg13g2_decap_8 FILLER_69_1045 ();
 sg13g2_decap_8 FILLER_69_1052 ();
 sg13g2_decap_8 FILLER_69_1059 ();
 sg13g2_decap_8 FILLER_69_1066 ();
 sg13g2_decap_8 FILLER_69_1073 ();
 sg13g2_decap_8 FILLER_69_1080 ();
 sg13g2_decap_8 FILLER_69_1087 ();
 sg13g2_decap_8 FILLER_69_1094 ();
 sg13g2_decap_8 FILLER_69_1101 ();
 sg13g2_decap_8 FILLER_69_1108 ();
 sg13g2_decap_8 FILLER_69_1115 ();
 sg13g2_decap_8 FILLER_69_1122 ();
 sg13g2_decap_8 FILLER_69_1129 ();
 sg13g2_decap_8 FILLER_69_1136 ();
 sg13g2_decap_8 FILLER_69_1143 ();
 sg13g2_decap_8 FILLER_69_1150 ();
 sg13g2_decap_8 FILLER_69_1157 ();
 sg13g2_decap_8 FILLER_69_1164 ();
 sg13g2_decap_8 FILLER_69_1171 ();
 sg13g2_decap_8 FILLER_69_1178 ();
 sg13g2_decap_8 FILLER_69_1185 ();
 sg13g2_decap_8 FILLER_69_1192 ();
 sg13g2_decap_8 FILLER_69_1199 ();
 sg13g2_decap_8 FILLER_69_1206 ();
 sg13g2_decap_8 FILLER_69_1213 ();
 sg13g2_decap_8 FILLER_69_1220 ();
 sg13g2_decap_8 FILLER_69_1227 ();
 sg13g2_decap_8 FILLER_69_1234 ();
 sg13g2_decap_8 FILLER_69_1241 ();
 sg13g2_decap_8 FILLER_69_1248 ();
 sg13g2_decap_8 FILLER_69_1255 ();
 sg13g2_decap_8 FILLER_69_1262 ();
 sg13g2_decap_8 FILLER_69_1269 ();
 sg13g2_decap_8 FILLER_69_1276 ();
 sg13g2_decap_8 FILLER_69_1283 ();
 sg13g2_decap_8 FILLER_69_1290 ();
 sg13g2_decap_8 FILLER_69_1297 ();
 sg13g2_decap_8 FILLER_69_1304 ();
 sg13g2_decap_8 FILLER_69_1311 ();
 sg13g2_decap_8 FILLER_69_1318 ();
 sg13g2_decap_8 FILLER_69_1325 ();
 sg13g2_decap_8 FILLER_69_1332 ();
 sg13g2_decap_8 FILLER_69_1339 ();
 sg13g2_decap_8 FILLER_69_1346 ();
 sg13g2_decap_8 FILLER_69_1353 ();
 sg13g2_decap_8 FILLER_69_1360 ();
 sg13g2_decap_8 FILLER_69_1367 ();
 sg13g2_decap_8 FILLER_69_1374 ();
 sg13g2_decap_8 FILLER_69_1381 ();
 sg13g2_decap_8 FILLER_69_1388 ();
 sg13g2_decap_8 FILLER_69_1395 ();
 sg13g2_decap_8 FILLER_69_1402 ();
 sg13g2_decap_8 FILLER_69_1409 ();
 sg13g2_decap_8 FILLER_69_1416 ();
 sg13g2_decap_8 FILLER_69_1423 ();
 sg13g2_decap_8 FILLER_69_1430 ();
 sg13g2_decap_8 FILLER_69_1437 ();
 sg13g2_decap_8 FILLER_69_1444 ();
 sg13g2_decap_8 FILLER_69_1451 ();
 sg13g2_decap_8 FILLER_69_1458 ();
 sg13g2_decap_8 FILLER_69_1465 ();
 sg13g2_decap_8 FILLER_69_1472 ();
 sg13g2_decap_8 FILLER_69_1479 ();
 sg13g2_decap_8 FILLER_69_1486 ();
 sg13g2_decap_8 FILLER_69_1493 ();
 sg13g2_decap_8 FILLER_69_1500 ();
 sg13g2_decap_8 FILLER_69_1507 ();
 sg13g2_decap_8 FILLER_69_1514 ();
 sg13g2_decap_8 FILLER_69_1521 ();
 sg13g2_decap_8 FILLER_69_1528 ();
 sg13g2_decap_8 FILLER_69_1535 ();
 sg13g2_decap_8 FILLER_69_1542 ();
 sg13g2_decap_8 FILLER_69_1549 ();
 sg13g2_decap_8 FILLER_69_1556 ();
 sg13g2_decap_8 FILLER_69_1563 ();
 sg13g2_decap_8 FILLER_69_1570 ();
 sg13g2_decap_8 FILLER_69_1577 ();
 sg13g2_decap_8 FILLER_69_1584 ();
 sg13g2_decap_8 FILLER_69_1591 ();
 sg13g2_decap_8 FILLER_69_1598 ();
 sg13g2_decap_8 FILLER_69_1605 ();
 sg13g2_decap_8 FILLER_69_1612 ();
 sg13g2_decap_8 FILLER_69_1619 ();
 sg13g2_decap_8 FILLER_69_1626 ();
 sg13g2_decap_8 FILLER_69_1633 ();
 sg13g2_decap_8 FILLER_69_1640 ();
 sg13g2_decap_8 FILLER_69_1647 ();
 sg13g2_decap_8 FILLER_69_1654 ();
 sg13g2_decap_8 FILLER_69_1661 ();
 sg13g2_decap_8 FILLER_69_1668 ();
 sg13g2_decap_8 FILLER_69_1675 ();
 sg13g2_decap_8 FILLER_69_1682 ();
 sg13g2_decap_8 FILLER_69_1689 ();
 sg13g2_decap_8 FILLER_69_1696 ();
 sg13g2_decap_8 FILLER_69_1703 ();
 sg13g2_decap_8 FILLER_69_1710 ();
 sg13g2_decap_8 FILLER_69_1717 ();
 sg13g2_decap_8 FILLER_69_1724 ();
 sg13g2_decap_8 FILLER_69_1731 ();
 sg13g2_decap_8 FILLER_69_1738 ();
 sg13g2_decap_8 FILLER_69_1745 ();
 sg13g2_decap_8 FILLER_69_1752 ();
 sg13g2_decap_8 FILLER_69_1759 ();
 sg13g2_decap_8 FILLER_69_1766 ();
 sg13g2_decap_8 FILLER_69_1773 ();
 sg13g2_decap_8 FILLER_69_1780 ();
 sg13g2_decap_8 FILLER_69_1787 ();
 sg13g2_decap_8 FILLER_69_1794 ();
 sg13g2_decap_8 FILLER_69_1801 ();
 sg13g2_decap_8 FILLER_69_1808 ();
 sg13g2_decap_8 FILLER_69_1815 ();
 sg13g2_decap_8 FILLER_69_1822 ();
 sg13g2_decap_8 FILLER_69_1829 ();
 sg13g2_decap_8 FILLER_69_1836 ();
 sg13g2_decap_8 FILLER_69_1843 ();
 sg13g2_decap_8 FILLER_69_1850 ();
 sg13g2_decap_8 FILLER_69_1857 ();
 sg13g2_decap_8 FILLER_69_1864 ();
 sg13g2_decap_8 FILLER_69_1871 ();
 sg13g2_decap_8 FILLER_69_1878 ();
 sg13g2_decap_8 FILLER_69_1885 ();
 sg13g2_decap_8 FILLER_69_1892 ();
 sg13g2_decap_8 FILLER_69_1899 ();
 sg13g2_decap_8 FILLER_69_1906 ();
 sg13g2_decap_8 FILLER_69_1913 ();
 sg13g2_decap_8 FILLER_69_1920 ();
 sg13g2_decap_8 FILLER_69_1927 ();
 sg13g2_decap_8 FILLER_69_1934 ();
 sg13g2_decap_8 FILLER_69_1941 ();
 sg13g2_decap_8 FILLER_69_1948 ();
 sg13g2_decap_8 FILLER_69_1955 ();
 sg13g2_decap_8 FILLER_69_1962 ();
 sg13g2_decap_8 FILLER_69_1969 ();
 sg13g2_decap_8 FILLER_69_1976 ();
 sg13g2_decap_8 FILLER_69_1983 ();
 sg13g2_decap_8 FILLER_69_1990 ();
 sg13g2_decap_8 FILLER_69_1997 ();
 sg13g2_decap_8 FILLER_69_2004 ();
 sg13g2_decap_8 FILLER_69_2011 ();
 sg13g2_decap_8 FILLER_69_2018 ();
 sg13g2_decap_8 FILLER_69_2025 ();
 sg13g2_decap_8 FILLER_69_2032 ();
 sg13g2_decap_8 FILLER_69_2039 ();
 sg13g2_decap_8 FILLER_69_2046 ();
 sg13g2_decap_8 FILLER_69_2053 ();
 sg13g2_decap_8 FILLER_69_2060 ();
 sg13g2_decap_8 FILLER_69_2067 ();
 sg13g2_decap_8 FILLER_69_2074 ();
 sg13g2_decap_8 FILLER_69_2081 ();
 sg13g2_decap_8 FILLER_69_2088 ();
 sg13g2_decap_8 FILLER_69_2095 ();
 sg13g2_decap_8 FILLER_69_2102 ();
 sg13g2_decap_8 FILLER_69_2109 ();
 sg13g2_decap_8 FILLER_69_2116 ();
 sg13g2_decap_8 FILLER_69_2123 ();
 sg13g2_decap_8 FILLER_69_2130 ();
 sg13g2_decap_8 FILLER_69_2137 ();
 sg13g2_decap_8 FILLER_69_2144 ();
 sg13g2_decap_8 FILLER_69_2151 ();
 sg13g2_decap_8 FILLER_69_2158 ();
 sg13g2_decap_8 FILLER_69_2165 ();
 sg13g2_decap_8 FILLER_69_2172 ();
 sg13g2_decap_8 FILLER_69_2179 ();
 sg13g2_decap_8 FILLER_69_2186 ();
 sg13g2_decap_8 FILLER_69_2193 ();
 sg13g2_decap_8 FILLER_69_2200 ();
 sg13g2_decap_8 FILLER_69_2207 ();
 sg13g2_decap_8 FILLER_69_2214 ();
 sg13g2_decap_8 FILLER_69_2221 ();
 sg13g2_decap_8 FILLER_69_2228 ();
 sg13g2_decap_8 FILLER_69_2235 ();
 sg13g2_decap_8 FILLER_69_2242 ();
 sg13g2_decap_8 FILLER_69_2249 ();
 sg13g2_decap_8 FILLER_69_2256 ();
 sg13g2_decap_8 FILLER_69_2263 ();
 sg13g2_decap_8 FILLER_69_2270 ();
 sg13g2_decap_8 FILLER_69_2277 ();
 sg13g2_decap_8 FILLER_69_2284 ();
 sg13g2_decap_8 FILLER_69_2291 ();
 sg13g2_decap_8 FILLER_69_2298 ();
 sg13g2_decap_8 FILLER_69_2305 ();
 sg13g2_decap_8 FILLER_69_2312 ();
 sg13g2_decap_8 FILLER_69_2319 ();
 sg13g2_decap_8 FILLER_69_2326 ();
 sg13g2_decap_8 FILLER_69_2333 ();
 sg13g2_decap_8 FILLER_69_2340 ();
 sg13g2_decap_8 FILLER_69_2347 ();
 sg13g2_decap_8 FILLER_69_2354 ();
 sg13g2_decap_8 FILLER_69_2361 ();
 sg13g2_decap_8 FILLER_69_2368 ();
 sg13g2_decap_8 FILLER_69_2375 ();
 sg13g2_decap_8 FILLER_69_2382 ();
 sg13g2_decap_8 FILLER_69_2389 ();
 sg13g2_decap_8 FILLER_69_2396 ();
 sg13g2_decap_8 FILLER_69_2403 ();
 sg13g2_decap_8 FILLER_69_2410 ();
 sg13g2_decap_8 FILLER_69_2417 ();
 sg13g2_decap_8 FILLER_69_2424 ();
 sg13g2_decap_8 FILLER_69_2431 ();
 sg13g2_decap_8 FILLER_69_2438 ();
 sg13g2_decap_8 FILLER_69_2445 ();
 sg13g2_decap_8 FILLER_69_2452 ();
 sg13g2_decap_8 FILLER_69_2459 ();
 sg13g2_decap_8 FILLER_69_2466 ();
 sg13g2_decap_8 FILLER_69_2473 ();
 sg13g2_decap_8 FILLER_69_2480 ();
 sg13g2_decap_8 FILLER_69_2487 ();
 sg13g2_decap_8 FILLER_69_2494 ();
 sg13g2_decap_8 FILLER_69_2501 ();
 sg13g2_decap_8 FILLER_69_2508 ();
 sg13g2_decap_8 FILLER_69_2515 ();
 sg13g2_decap_8 FILLER_69_2522 ();
 sg13g2_decap_8 FILLER_69_2529 ();
 sg13g2_decap_8 FILLER_69_2536 ();
 sg13g2_decap_8 FILLER_69_2543 ();
 sg13g2_decap_8 FILLER_69_2550 ();
 sg13g2_decap_8 FILLER_69_2557 ();
 sg13g2_decap_8 FILLER_69_2564 ();
 sg13g2_decap_8 FILLER_69_2571 ();
 sg13g2_decap_8 FILLER_69_2578 ();
 sg13g2_decap_8 FILLER_69_2585 ();
 sg13g2_decap_8 FILLER_69_2592 ();
 sg13g2_decap_8 FILLER_69_2599 ();
 sg13g2_decap_8 FILLER_69_2606 ();
 sg13g2_decap_8 FILLER_69_2613 ();
 sg13g2_decap_8 FILLER_69_2620 ();
 sg13g2_decap_8 FILLER_69_2627 ();
 sg13g2_decap_8 FILLER_69_2634 ();
 sg13g2_decap_8 FILLER_69_2641 ();
 sg13g2_decap_8 FILLER_69_2648 ();
 sg13g2_decap_8 FILLER_69_2655 ();
 sg13g2_decap_8 FILLER_69_2662 ();
 sg13g2_decap_8 FILLER_69_2669 ();
 sg13g2_decap_8 FILLER_69_2676 ();
 sg13g2_decap_8 FILLER_69_2683 ();
 sg13g2_decap_8 FILLER_69_2690 ();
 sg13g2_decap_8 FILLER_69_2697 ();
 sg13g2_decap_8 FILLER_69_2704 ();
 sg13g2_decap_8 FILLER_69_2711 ();
 sg13g2_decap_8 FILLER_69_2718 ();
 sg13g2_decap_8 FILLER_69_2725 ();
 sg13g2_decap_8 FILLER_69_2732 ();
 sg13g2_decap_8 FILLER_69_2739 ();
 sg13g2_decap_8 FILLER_69_2746 ();
 sg13g2_decap_8 FILLER_69_2753 ();
 sg13g2_decap_8 FILLER_69_2760 ();
 sg13g2_decap_8 FILLER_69_2767 ();
 sg13g2_decap_8 FILLER_69_2774 ();
 sg13g2_decap_8 FILLER_69_2781 ();
 sg13g2_decap_8 FILLER_69_2788 ();
 sg13g2_decap_8 FILLER_69_2795 ();
 sg13g2_decap_8 FILLER_69_2802 ();
 sg13g2_decap_8 FILLER_69_2809 ();
 sg13g2_decap_8 FILLER_69_2816 ();
 sg13g2_decap_8 FILLER_69_2823 ();
 sg13g2_decap_8 FILLER_69_2830 ();
 sg13g2_decap_8 FILLER_69_2837 ();
 sg13g2_decap_8 FILLER_69_2844 ();
 sg13g2_decap_8 FILLER_69_2851 ();
 sg13g2_decap_8 FILLER_69_2858 ();
 sg13g2_decap_8 FILLER_69_2865 ();
 sg13g2_decap_8 FILLER_69_2872 ();
 sg13g2_decap_8 FILLER_69_2879 ();
 sg13g2_decap_8 FILLER_69_2886 ();
 sg13g2_decap_8 FILLER_69_2893 ();
 sg13g2_decap_8 FILLER_69_2900 ();
 sg13g2_decap_8 FILLER_69_2907 ();
 sg13g2_decap_8 FILLER_69_2914 ();
 sg13g2_decap_8 FILLER_69_2921 ();
 sg13g2_decap_8 FILLER_69_2928 ();
 sg13g2_decap_8 FILLER_69_2935 ();
 sg13g2_decap_8 FILLER_69_2942 ();
 sg13g2_decap_8 FILLER_69_2949 ();
 sg13g2_decap_8 FILLER_69_2956 ();
 sg13g2_decap_8 FILLER_69_2963 ();
 sg13g2_decap_8 FILLER_69_2970 ();
 sg13g2_decap_8 FILLER_69_2977 ();
 sg13g2_decap_8 FILLER_69_2984 ();
 sg13g2_decap_8 FILLER_69_2991 ();
 sg13g2_decap_8 FILLER_69_2998 ();
 sg13g2_decap_8 FILLER_69_3005 ();
 sg13g2_decap_8 FILLER_69_3012 ();
 sg13g2_decap_8 FILLER_69_3019 ();
 sg13g2_decap_8 FILLER_69_3026 ();
 sg13g2_decap_8 FILLER_69_3033 ();
 sg13g2_decap_8 FILLER_69_3040 ();
 sg13g2_decap_8 FILLER_69_3047 ();
 sg13g2_decap_8 FILLER_69_3054 ();
 sg13g2_decap_8 FILLER_69_3061 ();
 sg13g2_decap_8 FILLER_69_3068 ();
 sg13g2_decap_8 FILLER_69_3075 ();
 sg13g2_decap_8 FILLER_69_3082 ();
 sg13g2_decap_8 FILLER_69_3089 ();
 sg13g2_decap_8 FILLER_69_3096 ();
 sg13g2_decap_8 FILLER_69_3103 ();
 sg13g2_decap_8 FILLER_69_3110 ();
 sg13g2_decap_8 FILLER_69_3117 ();
 sg13g2_decap_8 FILLER_69_3124 ();
 sg13g2_decap_8 FILLER_69_3131 ();
 sg13g2_decap_8 FILLER_69_3138 ();
 sg13g2_decap_8 FILLER_69_3145 ();
 sg13g2_decap_8 FILLER_69_3152 ();
 sg13g2_decap_8 FILLER_69_3159 ();
 sg13g2_decap_8 FILLER_69_3166 ();
 sg13g2_decap_8 FILLER_69_3173 ();
 sg13g2_decap_8 FILLER_69_3180 ();
 sg13g2_decap_8 FILLER_69_3187 ();
 sg13g2_decap_8 FILLER_69_3194 ();
 sg13g2_decap_8 FILLER_69_3201 ();
 sg13g2_decap_8 FILLER_69_3208 ();
 sg13g2_decap_8 FILLER_69_3215 ();
 sg13g2_decap_8 FILLER_69_3222 ();
 sg13g2_decap_8 FILLER_69_3229 ();
 sg13g2_decap_8 FILLER_69_3236 ();
 sg13g2_decap_8 FILLER_69_3243 ();
 sg13g2_decap_8 FILLER_69_3250 ();
 sg13g2_decap_8 FILLER_69_3257 ();
 sg13g2_decap_8 FILLER_69_3264 ();
 sg13g2_decap_8 FILLER_69_3271 ();
 sg13g2_decap_8 FILLER_69_3278 ();
 sg13g2_decap_8 FILLER_69_3285 ();
 sg13g2_decap_8 FILLER_69_3292 ();
 sg13g2_decap_8 FILLER_69_3299 ();
 sg13g2_decap_8 FILLER_69_3306 ();
 sg13g2_decap_8 FILLER_69_3313 ();
 sg13g2_decap_8 FILLER_69_3320 ();
 sg13g2_decap_8 FILLER_69_3327 ();
 sg13g2_decap_8 FILLER_69_3334 ();
 sg13g2_decap_8 FILLER_69_3341 ();
 sg13g2_decap_8 FILLER_69_3348 ();
 sg13g2_decap_8 FILLER_69_3355 ();
 sg13g2_decap_8 FILLER_69_3362 ();
 sg13g2_decap_8 FILLER_69_3369 ();
 sg13g2_decap_8 FILLER_69_3376 ();
 sg13g2_decap_8 FILLER_69_3383 ();
 sg13g2_decap_8 FILLER_69_3390 ();
 sg13g2_decap_8 FILLER_69_3397 ();
 sg13g2_decap_8 FILLER_69_3404 ();
 sg13g2_decap_8 FILLER_69_3411 ();
 sg13g2_decap_8 FILLER_69_3418 ();
 sg13g2_decap_8 FILLER_69_3425 ();
 sg13g2_decap_8 FILLER_69_3432 ();
 sg13g2_decap_8 FILLER_69_3439 ();
 sg13g2_decap_8 FILLER_69_3446 ();
 sg13g2_decap_8 FILLER_69_3453 ();
 sg13g2_decap_8 FILLER_69_3460 ();
 sg13g2_decap_8 FILLER_69_3467 ();
 sg13g2_decap_8 FILLER_69_3474 ();
 sg13g2_decap_8 FILLER_69_3481 ();
 sg13g2_decap_8 FILLER_69_3488 ();
 sg13g2_decap_8 FILLER_69_3495 ();
 sg13g2_decap_8 FILLER_69_3502 ();
 sg13g2_decap_8 FILLER_69_3509 ();
 sg13g2_decap_8 FILLER_69_3516 ();
 sg13g2_decap_8 FILLER_69_3523 ();
 sg13g2_decap_8 FILLER_69_3530 ();
 sg13g2_decap_8 FILLER_69_3537 ();
 sg13g2_decap_8 FILLER_69_3544 ();
 sg13g2_decap_8 FILLER_69_3551 ();
 sg13g2_decap_8 FILLER_69_3558 ();
 sg13g2_decap_8 FILLER_69_3565 ();
 sg13g2_decap_8 FILLER_69_3572 ();
 sg13g2_fill_1 FILLER_69_3579 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_decap_8 FILLER_70_133 ();
 sg13g2_decap_8 FILLER_70_140 ();
 sg13g2_decap_8 FILLER_70_147 ();
 sg13g2_decap_8 FILLER_70_154 ();
 sg13g2_fill_2 FILLER_70_161 ();
 sg13g2_decap_8 FILLER_70_167 ();
 sg13g2_fill_2 FILLER_70_174 ();
 sg13g2_fill_1 FILLER_70_194 ();
 sg13g2_fill_2 FILLER_70_208 ();
 sg13g2_fill_1 FILLER_70_210 ();
 sg13g2_fill_2 FILLER_70_225 ();
 sg13g2_decap_8 FILLER_70_246 ();
 sg13g2_decap_4 FILLER_70_253 ();
 sg13g2_fill_1 FILLER_70_257 ();
 sg13g2_decap_8 FILLER_70_263 ();
 sg13g2_fill_2 FILLER_70_270 ();
 sg13g2_decap_8 FILLER_70_285 ();
 sg13g2_decap_8 FILLER_70_292 ();
 sg13g2_decap_8 FILLER_70_299 ();
 sg13g2_decap_8 FILLER_70_306 ();
 sg13g2_decap_8 FILLER_70_313 ();
 sg13g2_decap_8 FILLER_70_320 ();
 sg13g2_decap_8 FILLER_70_327 ();
 sg13g2_decap_8 FILLER_70_334 ();
 sg13g2_decap_8 FILLER_70_341 ();
 sg13g2_decap_8 FILLER_70_348 ();
 sg13g2_decap_8 FILLER_70_355 ();
 sg13g2_decap_8 FILLER_70_362 ();
 sg13g2_decap_8 FILLER_70_369 ();
 sg13g2_decap_8 FILLER_70_376 ();
 sg13g2_decap_8 FILLER_70_383 ();
 sg13g2_decap_8 FILLER_70_390 ();
 sg13g2_decap_8 FILLER_70_397 ();
 sg13g2_decap_8 FILLER_70_404 ();
 sg13g2_decap_8 FILLER_70_411 ();
 sg13g2_decap_8 FILLER_70_418 ();
 sg13g2_decap_8 FILLER_70_425 ();
 sg13g2_decap_8 FILLER_70_432 ();
 sg13g2_decap_8 FILLER_70_439 ();
 sg13g2_decap_8 FILLER_70_446 ();
 sg13g2_decap_8 FILLER_70_453 ();
 sg13g2_decap_8 FILLER_70_460 ();
 sg13g2_decap_8 FILLER_70_467 ();
 sg13g2_decap_8 FILLER_70_474 ();
 sg13g2_decap_8 FILLER_70_481 ();
 sg13g2_decap_8 FILLER_70_488 ();
 sg13g2_decap_8 FILLER_70_495 ();
 sg13g2_decap_8 FILLER_70_502 ();
 sg13g2_decap_8 FILLER_70_509 ();
 sg13g2_decap_8 FILLER_70_516 ();
 sg13g2_decap_8 FILLER_70_523 ();
 sg13g2_decap_8 FILLER_70_530 ();
 sg13g2_decap_8 FILLER_70_537 ();
 sg13g2_decap_8 FILLER_70_544 ();
 sg13g2_decap_8 FILLER_70_551 ();
 sg13g2_decap_8 FILLER_70_558 ();
 sg13g2_decap_8 FILLER_70_565 ();
 sg13g2_decap_8 FILLER_70_572 ();
 sg13g2_decap_8 FILLER_70_579 ();
 sg13g2_decap_8 FILLER_70_586 ();
 sg13g2_decap_8 FILLER_70_593 ();
 sg13g2_decap_8 FILLER_70_600 ();
 sg13g2_decap_8 FILLER_70_607 ();
 sg13g2_decap_8 FILLER_70_614 ();
 sg13g2_decap_8 FILLER_70_621 ();
 sg13g2_decap_8 FILLER_70_628 ();
 sg13g2_decap_8 FILLER_70_635 ();
 sg13g2_decap_8 FILLER_70_642 ();
 sg13g2_decap_8 FILLER_70_649 ();
 sg13g2_decap_8 FILLER_70_656 ();
 sg13g2_decap_8 FILLER_70_663 ();
 sg13g2_decap_8 FILLER_70_670 ();
 sg13g2_decap_8 FILLER_70_677 ();
 sg13g2_decap_8 FILLER_70_684 ();
 sg13g2_decap_8 FILLER_70_691 ();
 sg13g2_decap_8 FILLER_70_698 ();
 sg13g2_decap_8 FILLER_70_705 ();
 sg13g2_decap_8 FILLER_70_712 ();
 sg13g2_decap_8 FILLER_70_719 ();
 sg13g2_decap_8 FILLER_70_726 ();
 sg13g2_decap_8 FILLER_70_733 ();
 sg13g2_decap_8 FILLER_70_740 ();
 sg13g2_decap_8 FILLER_70_747 ();
 sg13g2_decap_8 FILLER_70_754 ();
 sg13g2_decap_8 FILLER_70_761 ();
 sg13g2_decap_8 FILLER_70_768 ();
 sg13g2_decap_8 FILLER_70_775 ();
 sg13g2_decap_8 FILLER_70_782 ();
 sg13g2_decap_8 FILLER_70_789 ();
 sg13g2_decap_8 FILLER_70_796 ();
 sg13g2_decap_8 FILLER_70_803 ();
 sg13g2_decap_8 FILLER_70_810 ();
 sg13g2_decap_8 FILLER_70_817 ();
 sg13g2_decap_8 FILLER_70_824 ();
 sg13g2_decap_8 FILLER_70_831 ();
 sg13g2_decap_8 FILLER_70_838 ();
 sg13g2_decap_8 FILLER_70_845 ();
 sg13g2_decap_8 FILLER_70_852 ();
 sg13g2_decap_8 FILLER_70_859 ();
 sg13g2_decap_8 FILLER_70_866 ();
 sg13g2_decap_8 FILLER_70_873 ();
 sg13g2_decap_8 FILLER_70_880 ();
 sg13g2_decap_8 FILLER_70_887 ();
 sg13g2_decap_8 FILLER_70_894 ();
 sg13g2_decap_8 FILLER_70_901 ();
 sg13g2_decap_8 FILLER_70_908 ();
 sg13g2_decap_8 FILLER_70_915 ();
 sg13g2_decap_8 FILLER_70_922 ();
 sg13g2_decap_8 FILLER_70_929 ();
 sg13g2_decap_8 FILLER_70_936 ();
 sg13g2_decap_8 FILLER_70_943 ();
 sg13g2_decap_8 FILLER_70_950 ();
 sg13g2_decap_8 FILLER_70_957 ();
 sg13g2_decap_8 FILLER_70_964 ();
 sg13g2_decap_8 FILLER_70_971 ();
 sg13g2_decap_8 FILLER_70_978 ();
 sg13g2_decap_8 FILLER_70_985 ();
 sg13g2_decap_8 FILLER_70_992 ();
 sg13g2_decap_8 FILLER_70_999 ();
 sg13g2_decap_8 FILLER_70_1006 ();
 sg13g2_decap_8 FILLER_70_1013 ();
 sg13g2_decap_8 FILLER_70_1020 ();
 sg13g2_decap_8 FILLER_70_1027 ();
 sg13g2_decap_8 FILLER_70_1034 ();
 sg13g2_decap_8 FILLER_70_1041 ();
 sg13g2_decap_8 FILLER_70_1048 ();
 sg13g2_decap_8 FILLER_70_1055 ();
 sg13g2_decap_8 FILLER_70_1062 ();
 sg13g2_decap_8 FILLER_70_1069 ();
 sg13g2_decap_8 FILLER_70_1076 ();
 sg13g2_decap_8 FILLER_70_1083 ();
 sg13g2_decap_8 FILLER_70_1090 ();
 sg13g2_decap_8 FILLER_70_1097 ();
 sg13g2_decap_8 FILLER_70_1104 ();
 sg13g2_decap_8 FILLER_70_1111 ();
 sg13g2_decap_8 FILLER_70_1118 ();
 sg13g2_decap_8 FILLER_70_1125 ();
 sg13g2_decap_8 FILLER_70_1132 ();
 sg13g2_decap_8 FILLER_70_1139 ();
 sg13g2_decap_8 FILLER_70_1146 ();
 sg13g2_decap_8 FILLER_70_1153 ();
 sg13g2_decap_8 FILLER_70_1160 ();
 sg13g2_decap_8 FILLER_70_1167 ();
 sg13g2_decap_8 FILLER_70_1174 ();
 sg13g2_decap_8 FILLER_70_1181 ();
 sg13g2_decap_8 FILLER_70_1188 ();
 sg13g2_decap_8 FILLER_70_1195 ();
 sg13g2_decap_8 FILLER_70_1202 ();
 sg13g2_decap_8 FILLER_70_1209 ();
 sg13g2_decap_8 FILLER_70_1216 ();
 sg13g2_decap_8 FILLER_70_1223 ();
 sg13g2_decap_8 FILLER_70_1230 ();
 sg13g2_decap_8 FILLER_70_1237 ();
 sg13g2_decap_8 FILLER_70_1244 ();
 sg13g2_decap_8 FILLER_70_1251 ();
 sg13g2_decap_8 FILLER_70_1258 ();
 sg13g2_decap_8 FILLER_70_1265 ();
 sg13g2_decap_8 FILLER_70_1272 ();
 sg13g2_decap_8 FILLER_70_1279 ();
 sg13g2_decap_8 FILLER_70_1286 ();
 sg13g2_decap_8 FILLER_70_1293 ();
 sg13g2_decap_8 FILLER_70_1300 ();
 sg13g2_decap_8 FILLER_70_1307 ();
 sg13g2_decap_8 FILLER_70_1314 ();
 sg13g2_decap_8 FILLER_70_1321 ();
 sg13g2_decap_8 FILLER_70_1328 ();
 sg13g2_decap_8 FILLER_70_1335 ();
 sg13g2_decap_8 FILLER_70_1342 ();
 sg13g2_decap_8 FILLER_70_1349 ();
 sg13g2_decap_8 FILLER_70_1356 ();
 sg13g2_decap_8 FILLER_70_1363 ();
 sg13g2_decap_8 FILLER_70_1370 ();
 sg13g2_decap_8 FILLER_70_1377 ();
 sg13g2_decap_8 FILLER_70_1384 ();
 sg13g2_decap_8 FILLER_70_1391 ();
 sg13g2_decap_8 FILLER_70_1398 ();
 sg13g2_decap_8 FILLER_70_1405 ();
 sg13g2_decap_8 FILLER_70_1412 ();
 sg13g2_decap_8 FILLER_70_1419 ();
 sg13g2_decap_8 FILLER_70_1426 ();
 sg13g2_decap_8 FILLER_70_1433 ();
 sg13g2_decap_8 FILLER_70_1440 ();
 sg13g2_decap_8 FILLER_70_1447 ();
 sg13g2_decap_8 FILLER_70_1454 ();
 sg13g2_decap_8 FILLER_70_1461 ();
 sg13g2_decap_8 FILLER_70_1468 ();
 sg13g2_decap_8 FILLER_70_1475 ();
 sg13g2_decap_8 FILLER_70_1482 ();
 sg13g2_decap_8 FILLER_70_1489 ();
 sg13g2_decap_8 FILLER_70_1496 ();
 sg13g2_decap_8 FILLER_70_1503 ();
 sg13g2_decap_8 FILLER_70_1510 ();
 sg13g2_decap_8 FILLER_70_1517 ();
 sg13g2_decap_8 FILLER_70_1524 ();
 sg13g2_decap_8 FILLER_70_1531 ();
 sg13g2_decap_8 FILLER_70_1538 ();
 sg13g2_decap_8 FILLER_70_1545 ();
 sg13g2_decap_8 FILLER_70_1552 ();
 sg13g2_decap_8 FILLER_70_1559 ();
 sg13g2_decap_8 FILLER_70_1566 ();
 sg13g2_decap_8 FILLER_70_1573 ();
 sg13g2_decap_8 FILLER_70_1580 ();
 sg13g2_decap_8 FILLER_70_1587 ();
 sg13g2_decap_8 FILLER_70_1594 ();
 sg13g2_decap_8 FILLER_70_1601 ();
 sg13g2_decap_8 FILLER_70_1608 ();
 sg13g2_decap_8 FILLER_70_1615 ();
 sg13g2_decap_8 FILLER_70_1622 ();
 sg13g2_decap_8 FILLER_70_1629 ();
 sg13g2_decap_8 FILLER_70_1636 ();
 sg13g2_decap_8 FILLER_70_1643 ();
 sg13g2_decap_8 FILLER_70_1650 ();
 sg13g2_decap_8 FILLER_70_1657 ();
 sg13g2_decap_8 FILLER_70_1664 ();
 sg13g2_decap_8 FILLER_70_1671 ();
 sg13g2_decap_8 FILLER_70_1678 ();
 sg13g2_decap_8 FILLER_70_1685 ();
 sg13g2_decap_8 FILLER_70_1692 ();
 sg13g2_decap_8 FILLER_70_1699 ();
 sg13g2_decap_8 FILLER_70_1706 ();
 sg13g2_decap_8 FILLER_70_1713 ();
 sg13g2_decap_8 FILLER_70_1720 ();
 sg13g2_decap_8 FILLER_70_1727 ();
 sg13g2_decap_8 FILLER_70_1734 ();
 sg13g2_decap_8 FILLER_70_1741 ();
 sg13g2_decap_8 FILLER_70_1748 ();
 sg13g2_decap_8 FILLER_70_1755 ();
 sg13g2_decap_8 FILLER_70_1762 ();
 sg13g2_decap_8 FILLER_70_1769 ();
 sg13g2_decap_8 FILLER_70_1776 ();
 sg13g2_decap_8 FILLER_70_1783 ();
 sg13g2_decap_8 FILLER_70_1790 ();
 sg13g2_decap_8 FILLER_70_1797 ();
 sg13g2_decap_8 FILLER_70_1804 ();
 sg13g2_decap_8 FILLER_70_1811 ();
 sg13g2_decap_8 FILLER_70_1818 ();
 sg13g2_decap_8 FILLER_70_1825 ();
 sg13g2_decap_8 FILLER_70_1832 ();
 sg13g2_decap_8 FILLER_70_1839 ();
 sg13g2_decap_8 FILLER_70_1846 ();
 sg13g2_decap_8 FILLER_70_1853 ();
 sg13g2_decap_8 FILLER_70_1860 ();
 sg13g2_decap_8 FILLER_70_1867 ();
 sg13g2_decap_8 FILLER_70_1874 ();
 sg13g2_decap_8 FILLER_70_1881 ();
 sg13g2_decap_8 FILLER_70_1888 ();
 sg13g2_decap_8 FILLER_70_1895 ();
 sg13g2_decap_8 FILLER_70_1902 ();
 sg13g2_decap_8 FILLER_70_1909 ();
 sg13g2_decap_8 FILLER_70_1916 ();
 sg13g2_decap_8 FILLER_70_1923 ();
 sg13g2_decap_8 FILLER_70_1930 ();
 sg13g2_decap_8 FILLER_70_1937 ();
 sg13g2_decap_8 FILLER_70_1944 ();
 sg13g2_decap_8 FILLER_70_1951 ();
 sg13g2_decap_8 FILLER_70_1958 ();
 sg13g2_decap_8 FILLER_70_1965 ();
 sg13g2_decap_8 FILLER_70_1972 ();
 sg13g2_decap_8 FILLER_70_1979 ();
 sg13g2_decap_8 FILLER_70_1986 ();
 sg13g2_decap_8 FILLER_70_1993 ();
 sg13g2_decap_8 FILLER_70_2000 ();
 sg13g2_decap_8 FILLER_70_2007 ();
 sg13g2_decap_8 FILLER_70_2014 ();
 sg13g2_decap_8 FILLER_70_2021 ();
 sg13g2_decap_8 FILLER_70_2028 ();
 sg13g2_decap_8 FILLER_70_2035 ();
 sg13g2_decap_8 FILLER_70_2042 ();
 sg13g2_decap_8 FILLER_70_2049 ();
 sg13g2_decap_8 FILLER_70_2056 ();
 sg13g2_decap_8 FILLER_70_2063 ();
 sg13g2_decap_8 FILLER_70_2070 ();
 sg13g2_decap_8 FILLER_70_2077 ();
 sg13g2_decap_8 FILLER_70_2084 ();
 sg13g2_decap_8 FILLER_70_2091 ();
 sg13g2_decap_8 FILLER_70_2098 ();
 sg13g2_decap_8 FILLER_70_2105 ();
 sg13g2_decap_8 FILLER_70_2112 ();
 sg13g2_decap_8 FILLER_70_2119 ();
 sg13g2_decap_8 FILLER_70_2126 ();
 sg13g2_decap_8 FILLER_70_2133 ();
 sg13g2_decap_8 FILLER_70_2140 ();
 sg13g2_decap_8 FILLER_70_2147 ();
 sg13g2_decap_8 FILLER_70_2154 ();
 sg13g2_decap_8 FILLER_70_2161 ();
 sg13g2_decap_8 FILLER_70_2168 ();
 sg13g2_decap_8 FILLER_70_2175 ();
 sg13g2_decap_8 FILLER_70_2182 ();
 sg13g2_decap_8 FILLER_70_2189 ();
 sg13g2_decap_8 FILLER_70_2196 ();
 sg13g2_decap_8 FILLER_70_2203 ();
 sg13g2_decap_8 FILLER_70_2210 ();
 sg13g2_decap_8 FILLER_70_2217 ();
 sg13g2_decap_8 FILLER_70_2224 ();
 sg13g2_decap_8 FILLER_70_2231 ();
 sg13g2_decap_8 FILLER_70_2238 ();
 sg13g2_decap_8 FILLER_70_2245 ();
 sg13g2_decap_8 FILLER_70_2252 ();
 sg13g2_decap_8 FILLER_70_2259 ();
 sg13g2_decap_8 FILLER_70_2266 ();
 sg13g2_decap_8 FILLER_70_2273 ();
 sg13g2_decap_8 FILLER_70_2280 ();
 sg13g2_decap_8 FILLER_70_2287 ();
 sg13g2_decap_8 FILLER_70_2294 ();
 sg13g2_decap_8 FILLER_70_2301 ();
 sg13g2_decap_8 FILLER_70_2308 ();
 sg13g2_decap_8 FILLER_70_2315 ();
 sg13g2_decap_8 FILLER_70_2322 ();
 sg13g2_decap_8 FILLER_70_2329 ();
 sg13g2_decap_8 FILLER_70_2336 ();
 sg13g2_decap_8 FILLER_70_2343 ();
 sg13g2_decap_8 FILLER_70_2350 ();
 sg13g2_decap_8 FILLER_70_2357 ();
 sg13g2_decap_8 FILLER_70_2364 ();
 sg13g2_decap_8 FILLER_70_2371 ();
 sg13g2_decap_8 FILLER_70_2378 ();
 sg13g2_decap_8 FILLER_70_2385 ();
 sg13g2_decap_8 FILLER_70_2392 ();
 sg13g2_decap_8 FILLER_70_2399 ();
 sg13g2_decap_8 FILLER_70_2406 ();
 sg13g2_decap_8 FILLER_70_2413 ();
 sg13g2_decap_8 FILLER_70_2420 ();
 sg13g2_decap_8 FILLER_70_2427 ();
 sg13g2_decap_8 FILLER_70_2434 ();
 sg13g2_decap_8 FILLER_70_2441 ();
 sg13g2_decap_8 FILLER_70_2448 ();
 sg13g2_decap_8 FILLER_70_2455 ();
 sg13g2_decap_8 FILLER_70_2462 ();
 sg13g2_decap_8 FILLER_70_2469 ();
 sg13g2_decap_8 FILLER_70_2476 ();
 sg13g2_decap_8 FILLER_70_2483 ();
 sg13g2_decap_8 FILLER_70_2490 ();
 sg13g2_decap_8 FILLER_70_2497 ();
 sg13g2_decap_8 FILLER_70_2504 ();
 sg13g2_decap_8 FILLER_70_2511 ();
 sg13g2_decap_8 FILLER_70_2518 ();
 sg13g2_decap_8 FILLER_70_2525 ();
 sg13g2_decap_8 FILLER_70_2532 ();
 sg13g2_decap_8 FILLER_70_2539 ();
 sg13g2_decap_8 FILLER_70_2546 ();
 sg13g2_decap_8 FILLER_70_2553 ();
 sg13g2_decap_8 FILLER_70_2560 ();
 sg13g2_decap_8 FILLER_70_2567 ();
 sg13g2_decap_8 FILLER_70_2574 ();
 sg13g2_decap_8 FILLER_70_2581 ();
 sg13g2_decap_8 FILLER_70_2588 ();
 sg13g2_decap_8 FILLER_70_2595 ();
 sg13g2_decap_8 FILLER_70_2602 ();
 sg13g2_decap_8 FILLER_70_2609 ();
 sg13g2_decap_8 FILLER_70_2616 ();
 sg13g2_decap_8 FILLER_70_2623 ();
 sg13g2_decap_8 FILLER_70_2630 ();
 sg13g2_decap_8 FILLER_70_2637 ();
 sg13g2_decap_8 FILLER_70_2644 ();
 sg13g2_decap_8 FILLER_70_2651 ();
 sg13g2_decap_8 FILLER_70_2658 ();
 sg13g2_decap_8 FILLER_70_2665 ();
 sg13g2_decap_8 FILLER_70_2672 ();
 sg13g2_decap_8 FILLER_70_2679 ();
 sg13g2_decap_8 FILLER_70_2686 ();
 sg13g2_decap_8 FILLER_70_2693 ();
 sg13g2_decap_8 FILLER_70_2700 ();
 sg13g2_decap_8 FILLER_70_2707 ();
 sg13g2_decap_8 FILLER_70_2714 ();
 sg13g2_decap_8 FILLER_70_2721 ();
 sg13g2_decap_8 FILLER_70_2728 ();
 sg13g2_decap_8 FILLER_70_2735 ();
 sg13g2_decap_8 FILLER_70_2742 ();
 sg13g2_decap_8 FILLER_70_2749 ();
 sg13g2_decap_8 FILLER_70_2756 ();
 sg13g2_decap_8 FILLER_70_2763 ();
 sg13g2_decap_8 FILLER_70_2770 ();
 sg13g2_decap_8 FILLER_70_2777 ();
 sg13g2_decap_8 FILLER_70_2784 ();
 sg13g2_decap_8 FILLER_70_2791 ();
 sg13g2_decap_8 FILLER_70_2798 ();
 sg13g2_decap_8 FILLER_70_2805 ();
 sg13g2_decap_8 FILLER_70_2812 ();
 sg13g2_decap_8 FILLER_70_2819 ();
 sg13g2_decap_8 FILLER_70_2826 ();
 sg13g2_decap_8 FILLER_70_2833 ();
 sg13g2_decap_8 FILLER_70_2840 ();
 sg13g2_decap_8 FILLER_70_2847 ();
 sg13g2_decap_8 FILLER_70_2854 ();
 sg13g2_decap_8 FILLER_70_2861 ();
 sg13g2_decap_8 FILLER_70_2868 ();
 sg13g2_decap_8 FILLER_70_2875 ();
 sg13g2_decap_8 FILLER_70_2882 ();
 sg13g2_decap_8 FILLER_70_2889 ();
 sg13g2_decap_8 FILLER_70_2896 ();
 sg13g2_decap_8 FILLER_70_2903 ();
 sg13g2_decap_8 FILLER_70_2910 ();
 sg13g2_decap_8 FILLER_70_2917 ();
 sg13g2_decap_8 FILLER_70_2924 ();
 sg13g2_decap_8 FILLER_70_2931 ();
 sg13g2_decap_8 FILLER_70_2938 ();
 sg13g2_decap_8 FILLER_70_2945 ();
 sg13g2_decap_8 FILLER_70_2952 ();
 sg13g2_decap_8 FILLER_70_2959 ();
 sg13g2_decap_8 FILLER_70_2966 ();
 sg13g2_decap_8 FILLER_70_2973 ();
 sg13g2_decap_8 FILLER_70_2980 ();
 sg13g2_decap_8 FILLER_70_2987 ();
 sg13g2_decap_8 FILLER_70_2994 ();
 sg13g2_decap_8 FILLER_70_3001 ();
 sg13g2_decap_8 FILLER_70_3008 ();
 sg13g2_decap_8 FILLER_70_3015 ();
 sg13g2_decap_8 FILLER_70_3022 ();
 sg13g2_decap_8 FILLER_70_3029 ();
 sg13g2_decap_8 FILLER_70_3036 ();
 sg13g2_decap_8 FILLER_70_3043 ();
 sg13g2_decap_8 FILLER_70_3050 ();
 sg13g2_decap_8 FILLER_70_3057 ();
 sg13g2_decap_8 FILLER_70_3064 ();
 sg13g2_decap_8 FILLER_70_3071 ();
 sg13g2_decap_8 FILLER_70_3078 ();
 sg13g2_decap_8 FILLER_70_3085 ();
 sg13g2_decap_8 FILLER_70_3092 ();
 sg13g2_decap_8 FILLER_70_3099 ();
 sg13g2_decap_8 FILLER_70_3106 ();
 sg13g2_decap_8 FILLER_70_3113 ();
 sg13g2_decap_8 FILLER_70_3120 ();
 sg13g2_decap_8 FILLER_70_3127 ();
 sg13g2_decap_8 FILLER_70_3134 ();
 sg13g2_decap_8 FILLER_70_3141 ();
 sg13g2_decap_8 FILLER_70_3148 ();
 sg13g2_decap_8 FILLER_70_3155 ();
 sg13g2_decap_8 FILLER_70_3162 ();
 sg13g2_decap_8 FILLER_70_3169 ();
 sg13g2_decap_8 FILLER_70_3176 ();
 sg13g2_decap_8 FILLER_70_3183 ();
 sg13g2_decap_8 FILLER_70_3190 ();
 sg13g2_decap_8 FILLER_70_3197 ();
 sg13g2_decap_8 FILLER_70_3204 ();
 sg13g2_decap_8 FILLER_70_3211 ();
 sg13g2_decap_8 FILLER_70_3218 ();
 sg13g2_decap_8 FILLER_70_3225 ();
 sg13g2_decap_8 FILLER_70_3232 ();
 sg13g2_decap_8 FILLER_70_3239 ();
 sg13g2_decap_8 FILLER_70_3246 ();
 sg13g2_decap_8 FILLER_70_3253 ();
 sg13g2_decap_8 FILLER_70_3260 ();
 sg13g2_decap_8 FILLER_70_3267 ();
 sg13g2_decap_8 FILLER_70_3274 ();
 sg13g2_decap_8 FILLER_70_3281 ();
 sg13g2_decap_8 FILLER_70_3288 ();
 sg13g2_decap_8 FILLER_70_3295 ();
 sg13g2_decap_8 FILLER_70_3302 ();
 sg13g2_decap_8 FILLER_70_3309 ();
 sg13g2_decap_8 FILLER_70_3316 ();
 sg13g2_decap_8 FILLER_70_3323 ();
 sg13g2_decap_8 FILLER_70_3330 ();
 sg13g2_decap_8 FILLER_70_3337 ();
 sg13g2_decap_8 FILLER_70_3344 ();
 sg13g2_decap_8 FILLER_70_3351 ();
 sg13g2_decap_8 FILLER_70_3358 ();
 sg13g2_decap_8 FILLER_70_3365 ();
 sg13g2_decap_8 FILLER_70_3372 ();
 sg13g2_decap_8 FILLER_70_3379 ();
 sg13g2_decap_8 FILLER_70_3386 ();
 sg13g2_decap_8 FILLER_70_3393 ();
 sg13g2_decap_8 FILLER_70_3400 ();
 sg13g2_decap_8 FILLER_70_3407 ();
 sg13g2_decap_8 FILLER_70_3414 ();
 sg13g2_decap_8 FILLER_70_3421 ();
 sg13g2_decap_8 FILLER_70_3428 ();
 sg13g2_decap_8 FILLER_70_3435 ();
 sg13g2_decap_8 FILLER_70_3442 ();
 sg13g2_decap_8 FILLER_70_3449 ();
 sg13g2_decap_8 FILLER_70_3456 ();
 sg13g2_decap_8 FILLER_70_3463 ();
 sg13g2_decap_8 FILLER_70_3470 ();
 sg13g2_decap_8 FILLER_70_3477 ();
 sg13g2_decap_8 FILLER_70_3484 ();
 sg13g2_decap_8 FILLER_70_3491 ();
 sg13g2_decap_8 FILLER_70_3498 ();
 sg13g2_decap_8 FILLER_70_3505 ();
 sg13g2_decap_8 FILLER_70_3512 ();
 sg13g2_decap_8 FILLER_70_3519 ();
 sg13g2_decap_8 FILLER_70_3526 ();
 sg13g2_decap_8 FILLER_70_3533 ();
 sg13g2_decap_8 FILLER_70_3540 ();
 sg13g2_decap_8 FILLER_70_3547 ();
 sg13g2_decap_8 FILLER_70_3554 ();
 sg13g2_decap_8 FILLER_70_3561 ();
 sg13g2_decap_8 FILLER_70_3568 ();
 sg13g2_decap_4 FILLER_70_3575 ();
 sg13g2_fill_1 FILLER_70_3579 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_133 ();
 sg13g2_decap_8 FILLER_71_140 ();
 sg13g2_decap_8 FILLER_71_147 ();
 sg13g2_decap_8 FILLER_71_154 ();
 sg13g2_fill_1 FILLER_71_165 ();
 sg13g2_fill_1 FILLER_71_201 ();
 sg13g2_fill_1 FILLER_71_242 ();
 sg13g2_fill_1 FILLER_71_251 ();
 sg13g2_fill_1 FILLER_71_265 ();
 sg13g2_decap_8 FILLER_71_294 ();
 sg13g2_decap_8 FILLER_71_301 ();
 sg13g2_decap_8 FILLER_71_308 ();
 sg13g2_decap_8 FILLER_71_315 ();
 sg13g2_decap_8 FILLER_71_322 ();
 sg13g2_decap_8 FILLER_71_329 ();
 sg13g2_decap_8 FILLER_71_336 ();
 sg13g2_decap_8 FILLER_71_343 ();
 sg13g2_decap_8 FILLER_71_350 ();
 sg13g2_decap_8 FILLER_71_357 ();
 sg13g2_decap_8 FILLER_71_364 ();
 sg13g2_decap_8 FILLER_71_371 ();
 sg13g2_decap_8 FILLER_71_378 ();
 sg13g2_decap_8 FILLER_71_385 ();
 sg13g2_decap_8 FILLER_71_392 ();
 sg13g2_decap_8 FILLER_71_399 ();
 sg13g2_decap_8 FILLER_71_406 ();
 sg13g2_decap_8 FILLER_71_413 ();
 sg13g2_decap_8 FILLER_71_420 ();
 sg13g2_decap_8 FILLER_71_427 ();
 sg13g2_decap_8 FILLER_71_434 ();
 sg13g2_decap_8 FILLER_71_441 ();
 sg13g2_decap_8 FILLER_71_448 ();
 sg13g2_decap_8 FILLER_71_455 ();
 sg13g2_decap_8 FILLER_71_462 ();
 sg13g2_decap_8 FILLER_71_469 ();
 sg13g2_decap_8 FILLER_71_476 ();
 sg13g2_decap_8 FILLER_71_483 ();
 sg13g2_decap_8 FILLER_71_490 ();
 sg13g2_decap_8 FILLER_71_497 ();
 sg13g2_decap_8 FILLER_71_504 ();
 sg13g2_decap_8 FILLER_71_511 ();
 sg13g2_decap_8 FILLER_71_518 ();
 sg13g2_decap_8 FILLER_71_525 ();
 sg13g2_decap_8 FILLER_71_532 ();
 sg13g2_decap_8 FILLER_71_539 ();
 sg13g2_decap_8 FILLER_71_546 ();
 sg13g2_decap_8 FILLER_71_553 ();
 sg13g2_decap_8 FILLER_71_560 ();
 sg13g2_decap_8 FILLER_71_567 ();
 sg13g2_decap_8 FILLER_71_574 ();
 sg13g2_decap_8 FILLER_71_581 ();
 sg13g2_decap_8 FILLER_71_588 ();
 sg13g2_decap_8 FILLER_71_595 ();
 sg13g2_decap_8 FILLER_71_602 ();
 sg13g2_decap_8 FILLER_71_609 ();
 sg13g2_decap_8 FILLER_71_616 ();
 sg13g2_decap_8 FILLER_71_623 ();
 sg13g2_decap_8 FILLER_71_630 ();
 sg13g2_decap_8 FILLER_71_637 ();
 sg13g2_decap_8 FILLER_71_644 ();
 sg13g2_decap_8 FILLER_71_651 ();
 sg13g2_decap_8 FILLER_71_658 ();
 sg13g2_decap_8 FILLER_71_665 ();
 sg13g2_decap_8 FILLER_71_672 ();
 sg13g2_decap_8 FILLER_71_679 ();
 sg13g2_decap_8 FILLER_71_686 ();
 sg13g2_decap_8 FILLER_71_693 ();
 sg13g2_decap_8 FILLER_71_700 ();
 sg13g2_decap_8 FILLER_71_707 ();
 sg13g2_decap_8 FILLER_71_714 ();
 sg13g2_decap_8 FILLER_71_721 ();
 sg13g2_decap_8 FILLER_71_728 ();
 sg13g2_decap_8 FILLER_71_735 ();
 sg13g2_decap_8 FILLER_71_742 ();
 sg13g2_decap_8 FILLER_71_749 ();
 sg13g2_decap_8 FILLER_71_756 ();
 sg13g2_decap_8 FILLER_71_763 ();
 sg13g2_decap_8 FILLER_71_770 ();
 sg13g2_decap_8 FILLER_71_777 ();
 sg13g2_decap_8 FILLER_71_784 ();
 sg13g2_decap_8 FILLER_71_791 ();
 sg13g2_decap_8 FILLER_71_798 ();
 sg13g2_decap_8 FILLER_71_805 ();
 sg13g2_decap_8 FILLER_71_812 ();
 sg13g2_decap_8 FILLER_71_819 ();
 sg13g2_decap_8 FILLER_71_826 ();
 sg13g2_decap_8 FILLER_71_833 ();
 sg13g2_decap_8 FILLER_71_840 ();
 sg13g2_decap_8 FILLER_71_847 ();
 sg13g2_decap_8 FILLER_71_854 ();
 sg13g2_decap_8 FILLER_71_861 ();
 sg13g2_decap_8 FILLER_71_868 ();
 sg13g2_decap_8 FILLER_71_875 ();
 sg13g2_decap_8 FILLER_71_882 ();
 sg13g2_decap_8 FILLER_71_889 ();
 sg13g2_decap_8 FILLER_71_896 ();
 sg13g2_decap_8 FILLER_71_903 ();
 sg13g2_decap_8 FILLER_71_910 ();
 sg13g2_decap_8 FILLER_71_917 ();
 sg13g2_decap_8 FILLER_71_924 ();
 sg13g2_decap_8 FILLER_71_931 ();
 sg13g2_decap_8 FILLER_71_938 ();
 sg13g2_decap_8 FILLER_71_945 ();
 sg13g2_decap_8 FILLER_71_952 ();
 sg13g2_decap_8 FILLER_71_959 ();
 sg13g2_decap_8 FILLER_71_966 ();
 sg13g2_decap_8 FILLER_71_973 ();
 sg13g2_decap_8 FILLER_71_980 ();
 sg13g2_decap_8 FILLER_71_987 ();
 sg13g2_decap_8 FILLER_71_994 ();
 sg13g2_decap_8 FILLER_71_1001 ();
 sg13g2_decap_8 FILLER_71_1008 ();
 sg13g2_decap_8 FILLER_71_1015 ();
 sg13g2_decap_8 FILLER_71_1022 ();
 sg13g2_decap_8 FILLER_71_1029 ();
 sg13g2_decap_8 FILLER_71_1036 ();
 sg13g2_decap_8 FILLER_71_1043 ();
 sg13g2_decap_8 FILLER_71_1050 ();
 sg13g2_decap_8 FILLER_71_1057 ();
 sg13g2_decap_8 FILLER_71_1064 ();
 sg13g2_decap_8 FILLER_71_1071 ();
 sg13g2_decap_8 FILLER_71_1078 ();
 sg13g2_decap_8 FILLER_71_1085 ();
 sg13g2_decap_8 FILLER_71_1092 ();
 sg13g2_decap_8 FILLER_71_1099 ();
 sg13g2_decap_8 FILLER_71_1106 ();
 sg13g2_decap_8 FILLER_71_1113 ();
 sg13g2_decap_8 FILLER_71_1120 ();
 sg13g2_decap_8 FILLER_71_1127 ();
 sg13g2_decap_8 FILLER_71_1134 ();
 sg13g2_decap_8 FILLER_71_1141 ();
 sg13g2_decap_8 FILLER_71_1148 ();
 sg13g2_decap_8 FILLER_71_1155 ();
 sg13g2_decap_8 FILLER_71_1162 ();
 sg13g2_decap_8 FILLER_71_1169 ();
 sg13g2_decap_8 FILLER_71_1176 ();
 sg13g2_decap_8 FILLER_71_1183 ();
 sg13g2_decap_8 FILLER_71_1190 ();
 sg13g2_decap_8 FILLER_71_1197 ();
 sg13g2_decap_8 FILLER_71_1204 ();
 sg13g2_decap_8 FILLER_71_1211 ();
 sg13g2_decap_8 FILLER_71_1218 ();
 sg13g2_decap_8 FILLER_71_1225 ();
 sg13g2_decap_8 FILLER_71_1232 ();
 sg13g2_decap_8 FILLER_71_1239 ();
 sg13g2_decap_8 FILLER_71_1246 ();
 sg13g2_decap_8 FILLER_71_1253 ();
 sg13g2_decap_8 FILLER_71_1260 ();
 sg13g2_decap_8 FILLER_71_1267 ();
 sg13g2_decap_8 FILLER_71_1274 ();
 sg13g2_decap_8 FILLER_71_1281 ();
 sg13g2_decap_8 FILLER_71_1288 ();
 sg13g2_decap_8 FILLER_71_1295 ();
 sg13g2_decap_8 FILLER_71_1302 ();
 sg13g2_decap_8 FILLER_71_1309 ();
 sg13g2_decap_8 FILLER_71_1316 ();
 sg13g2_decap_8 FILLER_71_1323 ();
 sg13g2_decap_8 FILLER_71_1330 ();
 sg13g2_decap_8 FILLER_71_1337 ();
 sg13g2_decap_8 FILLER_71_1344 ();
 sg13g2_decap_8 FILLER_71_1351 ();
 sg13g2_decap_8 FILLER_71_1358 ();
 sg13g2_decap_8 FILLER_71_1365 ();
 sg13g2_decap_8 FILLER_71_1372 ();
 sg13g2_decap_8 FILLER_71_1379 ();
 sg13g2_decap_8 FILLER_71_1386 ();
 sg13g2_decap_8 FILLER_71_1393 ();
 sg13g2_decap_8 FILLER_71_1400 ();
 sg13g2_decap_8 FILLER_71_1407 ();
 sg13g2_decap_8 FILLER_71_1414 ();
 sg13g2_decap_8 FILLER_71_1421 ();
 sg13g2_decap_8 FILLER_71_1428 ();
 sg13g2_decap_8 FILLER_71_1435 ();
 sg13g2_decap_8 FILLER_71_1442 ();
 sg13g2_decap_8 FILLER_71_1449 ();
 sg13g2_decap_8 FILLER_71_1456 ();
 sg13g2_decap_8 FILLER_71_1463 ();
 sg13g2_decap_8 FILLER_71_1470 ();
 sg13g2_decap_8 FILLER_71_1477 ();
 sg13g2_decap_8 FILLER_71_1484 ();
 sg13g2_decap_8 FILLER_71_1491 ();
 sg13g2_decap_8 FILLER_71_1498 ();
 sg13g2_decap_8 FILLER_71_1505 ();
 sg13g2_decap_8 FILLER_71_1512 ();
 sg13g2_decap_8 FILLER_71_1519 ();
 sg13g2_decap_8 FILLER_71_1526 ();
 sg13g2_decap_8 FILLER_71_1533 ();
 sg13g2_decap_8 FILLER_71_1540 ();
 sg13g2_decap_8 FILLER_71_1547 ();
 sg13g2_decap_8 FILLER_71_1554 ();
 sg13g2_decap_8 FILLER_71_1561 ();
 sg13g2_decap_8 FILLER_71_1568 ();
 sg13g2_decap_8 FILLER_71_1575 ();
 sg13g2_decap_8 FILLER_71_1582 ();
 sg13g2_decap_8 FILLER_71_1589 ();
 sg13g2_decap_8 FILLER_71_1596 ();
 sg13g2_decap_8 FILLER_71_1603 ();
 sg13g2_decap_8 FILLER_71_1610 ();
 sg13g2_decap_8 FILLER_71_1617 ();
 sg13g2_decap_8 FILLER_71_1624 ();
 sg13g2_decap_8 FILLER_71_1631 ();
 sg13g2_decap_8 FILLER_71_1638 ();
 sg13g2_decap_8 FILLER_71_1645 ();
 sg13g2_decap_8 FILLER_71_1652 ();
 sg13g2_decap_8 FILLER_71_1659 ();
 sg13g2_decap_8 FILLER_71_1666 ();
 sg13g2_decap_8 FILLER_71_1673 ();
 sg13g2_decap_8 FILLER_71_1680 ();
 sg13g2_decap_8 FILLER_71_1687 ();
 sg13g2_decap_8 FILLER_71_1694 ();
 sg13g2_decap_8 FILLER_71_1701 ();
 sg13g2_decap_8 FILLER_71_1708 ();
 sg13g2_decap_8 FILLER_71_1715 ();
 sg13g2_decap_8 FILLER_71_1722 ();
 sg13g2_decap_8 FILLER_71_1729 ();
 sg13g2_decap_8 FILLER_71_1736 ();
 sg13g2_decap_8 FILLER_71_1743 ();
 sg13g2_decap_8 FILLER_71_1750 ();
 sg13g2_decap_8 FILLER_71_1757 ();
 sg13g2_decap_8 FILLER_71_1764 ();
 sg13g2_decap_8 FILLER_71_1771 ();
 sg13g2_decap_8 FILLER_71_1778 ();
 sg13g2_decap_8 FILLER_71_1785 ();
 sg13g2_decap_8 FILLER_71_1792 ();
 sg13g2_decap_8 FILLER_71_1799 ();
 sg13g2_decap_8 FILLER_71_1806 ();
 sg13g2_decap_8 FILLER_71_1813 ();
 sg13g2_decap_8 FILLER_71_1820 ();
 sg13g2_decap_8 FILLER_71_1827 ();
 sg13g2_decap_8 FILLER_71_1834 ();
 sg13g2_decap_8 FILLER_71_1841 ();
 sg13g2_decap_8 FILLER_71_1848 ();
 sg13g2_decap_8 FILLER_71_1855 ();
 sg13g2_decap_8 FILLER_71_1862 ();
 sg13g2_decap_8 FILLER_71_1869 ();
 sg13g2_decap_8 FILLER_71_1876 ();
 sg13g2_decap_8 FILLER_71_1883 ();
 sg13g2_decap_8 FILLER_71_1890 ();
 sg13g2_decap_8 FILLER_71_1897 ();
 sg13g2_decap_8 FILLER_71_1904 ();
 sg13g2_decap_8 FILLER_71_1911 ();
 sg13g2_decap_8 FILLER_71_1918 ();
 sg13g2_decap_8 FILLER_71_1925 ();
 sg13g2_decap_8 FILLER_71_1932 ();
 sg13g2_decap_8 FILLER_71_1939 ();
 sg13g2_decap_8 FILLER_71_1946 ();
 sg13g2_decap_8 FILLER_71_1953 ();
 sg13g2_decap_8 FILLER_71_1960 ();
 sg13g2_decap_8 FILLER_71_1967 ();
 sg13g2_decap_8 FILLER_71_1974 ();
 sg13g2_decap_8 FILLER_71_1981 ();
 sg13g2_decap_8 FILLER_71_1988 ();
 sg13g2_decap_8 FILLER_71_1995 ();
 sg13g2_decap_8 FILLER_71_2002 ();
 sg13g2_decap_8 FILLER_71_2009 ();
 sg13g2_decap_8 FILLER_71_2016 ();
 sg13g2_decap_8 FILLER_71_2023 ();
 sg13g2_decap_8 FILLER_71_2030 ();
 sg13g2_decap_8 FILLER_71_2037 ();
 sg13g2_decap_8 FILLER_71_2044 ();
 sg13g2_decap_8 FILLER_71_2051 ();
 sg13g2_decap_8 FILLER_71_2058 ();
 sg13g2_decap_8 FILLER_71_2065 ();
 sg13g2_decap_8 FILLER_71_2072 ();
 sg13g2_decap_8 FILLER_71_2079 ();
 sg13g2_decap_8 FILLER_71_2086 ();
 sg13g2_decap_8 FILLER_71_2093 ();
 sg13g2_decap_8 FILLER_71_2100 ();
 sg13g2_decap_8 FILLER_71_2107 ();
 sg13g2_decap_8 FILLER_71_2114 ();
 sg13g2_decap_8 FILLER_71_2121 ();
 sg13g2_decap_8 FILLER_71_2128 ();
 sg13g2_decap_8 FILLER_71_2135 ();
 sg13g2_decap_8 FILLER_71_2142 ();
 sg13g2_decap_8 FILLER_71_2149 ();
 sg13g2_decap_8 FILLER_71_2156 ();
 sg13g2_decap_8 FILLER_71_2163 ();
 sg13g2_decap_8 FILLER_71_2170 ();
 sg13g2_decap_8 FILLER_71_2177 ();
 sg13g2_decap_8 FILLER_71_2184 ();
 sg13g2_decap_8 FILLER_71_2191 ();
 sg13g2_decap_8 FILLER_71_2198 ();
 sg13g2_decap_8 FILLER_71_2205 ();
 sg13g2_decap_8 FILLER_71_2212 ();
 sg13g2_decap_8 FILLER_71_2219 ();
 sg13g2_decap_8 FILLER_71_2226 ();
 sg13g2_decap_8 FILLER_71_2233 ();
 sg13g2_decap_8 FILLER_71_2240 ();
 sg13g2_decap_8 FILLER_71_2247 ();
 sg13g2_decap_8 FILLER_71_2254 ();
 sg13g2_decap_8 FILLER_71_2261 ();
 sg13g2_decap_8 FILLER_71_2268 ();
 sg13g2_decap_8 FILLER_71_2275 ();
 sg13g2_decap_8 FILLER_71_2282 ();
 sg13g2_decap_8 FILLER_71_2289 ();
 sg13g2_decap_8 FILLER_71_2296 ();
 sg13g2_decap_8 FILLER_71_2303 ();
 sg13g2_decap_8 FILLER_71_2310 ();
 sg13g2_decap_8 FILLER_71_2317 ();
 sg13g2_decap_8 FILLER_71_2324 ();
 sg13g2_decap_8 FILLER_71_2331 ();
 sg13g2_decap_8 FILLER_71_2338 ();
 sg13g2_decap_8 FILLER_71_2345 ();
 sg13g2_decap_8 FILLER_71_2352 ();
 sg13g2_decap_8 FILLER_71_2359 ();
 sg13g2_decap_8 FILLER_71_2366 ();
 sg13g2_decap_8 FILLER_71_2373 ();
 sg13g2_decap_8 FILLER_71_2380 ();
 sg13g2_decap_8 FILLER_71_2387 ();
 sg13g2_decap_8 FILLER_71_2394 ();
 sg13g2_decap_8 FILLER_71_2401 ();
 sg13g2_decap_8 FILLER_71_2408 ();
 sg13g2_decap_8 FILLER_71_2415 ();
 sg13g2_decap_8 FILLER_71_2422 ();
 sg13g2_decap_8 FILLER_71_2429 ();
 sg13g2_decap_8 FILLER_71_2436 ();
 sg13g2_decap_8 FILLER_71_2443 ();
 sg13g2_decap_8 FILLER_71_2450 ();
 sg13g2_decap_8 FILLER_71_2457 ();
 sg13g2_decap_8 FILLER_71_2464 ();
 sg13g2_decap_8 FILLER_71_2471 ();
 sg13g2_decap_8 FILLER_71_2478 ();
 sg13g2_decap_8 FILLER_71_2485 ();
 sg13g2_decap_8 FILLER_71_2492 ();
 sg13g2_decap_8 FILLER_71_2499 ();
 sg13g2_decap_8 FILLER_71_2506 ();
 sg13g2_decap_8 FILLER_71_2513 ();
 sg13g2_decap_8 FILLER_71_2520 ();
 sg13g2_decap_8 FILLER_71_2527 ();
 sg13g2_decap_8 FILLER_71_2534 ();
 sg13g2_decap_8 FILLER_71_2541 ();
 sg13g2_decap_8 FILLER_71_2548 ();
 sg13g2_decap_8 FILLER_71_2555 ();
 sg13g2_decap_8 FILLER_71_2562 ();
 sg13g2_decap_8 FILLER_71_2569 ();
 sg13g2_decap_8 FILLER_71_2576 ();
 sg13g2_decap_8 FILLER_71_2583 ();
 sg13g2_decap_8 FILLER_71_2590 ();
 sg13g2_decap_8 FILLER_71_2597 ();
 sg13g2_decap_8 FILLER_71_2604 ();
 sg13g2_decap_8 FILLER_71_2611 ();
 sg13g2_decap_8 FILLER_71_2618 ();
 sg13g2_decap_8 FILLER_71_2625 ();
 sg13g2_decap_8 FILLER_71_2632 ();
 sg13g2_decap_8 FILLER_71_2639 ();
 sg13g2_decap_8 FILLER_71_2646 ();
 sg13g2_decap_8 FILLER_71_2653 ();
 sg13g2_decap_8 FILLER_71_2660 ();
 sg13g2_decap_8 FILLER_71_2667 ();
 sg13g2_decap_8 FILLER_71_2674 ();
 sg13g2_decap_8 FILLER_71_2681 ();
 sg13g2_decap_8 FILLER_71_2688 ();
 sg13g2_decap_8 FILLER_71_2695 ();
 sg13g2_decap_8 FILLER_71_2702 ();
 sg13g2_decap_8 FILLER_71_2709 ();
 sg13g2_decap_8 FILLER_71_2716 ();
 sg13g2_decap_8 FILLER_71_2723 ();
 sg13g2_decap_8 FILLER_71_2730 ();
 sg13g2_decap_8 FILLER_71_2737 ();
 sg13g2_decap_8 FILLER_71_2744 ();
 sg13g2_decap_8 FILLER_71_2751 ();
 sg13g2_decap_8 FILLER_71_2758 ();
 sg13g2_decap_8 FILLER_71_2765 ();
 sg13g2_decap_8 FILLER_71_2772 ();
 sg13g2_decap_8 FILLER_71_2779 ();
 sg13g2_decap_8 FILLER_71_2786 ();
 sg13g2_decap_8 FILLER_71_2793 ();
 sg13g2_decap_8 FILLER_71_2800 ();
 sg13g2_decap_8 FILLER_71_2807 ();
 sg13g2_decap_8 FILLER_71_2814 ();
 sg13g2_decap_8 FILLER_71_2821 ();
 sg13g2_decap_8 FILLER_71_2828 ();
 sg13g2_decap_8 FILLER_71_2835 ();
 sg13g2_decap_8 FILLER_71_2842 ();
 sg13g2_decap_8 FILLER_71_2849 ();
 sg13g2_decap_8 FILLER_71_2856 ();
 sg13g2_decap_8 FILLER_71_2863 ();
 sg13g2_decap_8 FILLER_71_2870 ();
 sg13g2_decap_8 FILLER_71_2877 ();
 sg13g2_decap_8 FILLER_71_2884 ();
 sg13g2_decap_8 FILLER_71_2891 ();
 sg13g2_decap_8 FILLER_71_2898 ();
 sg13g2_decap_8 FILLER_71_2905 ();
 sg13g2_decap_8 FILLER_71_2912 ();
 sg13g2_decap_8 FILLER_71_2919 ();
 sg13g2_decap_8 FILLER_71_2926 ();
 sg13g2_decap_8 FILLER_71_2933 ();
 sg13g2_decap_8 FILLER_71_2940 ();
 sg13g2_decap_8 FILLER_71_2947 ();
 sg13g2_decap_8 FILLER_71_2954 ();
 sg13g2_decap_8 FILLER_71_2961 ();
 sg13g2_decap_8 FILLER_71_2968 ();
 sg13g2_decap_8 FILLER_71_2975 ();
 sg13g2_decap_8 FILLER_71_2982 ();
 sg13g2_decap_8 FILLER_71_2989 ();
 sg13g2_decap_8 FILLER_71_2996 ();
 sg13g2_decap_8 FILLER_71_3003 ();
 sg13g2_decap_8 FILLER_71_3010 ();
 sg13g2_decap_8 FILLER_71_3017 ();
 sg13g2_decap_8 FILLER_71_3024 ();
 sg13g2_decap_8 FILLER_71_3031 ();
 sg13g2_decap_8 FILLER_71_3038 ();
 sg13g2_decap_8 FILLER_71_3045 ();
 sg13g2_decap_8 FILLER_71_3052 ();
 sg13g2_decap_8 FILLER_71_3059 ();
 sg13g2_decap_8 FILLER_71_3066 ();
 sg13g2_decap_8 FILLER_71_3073 ();
 sg13g2_decap_8 FILLER_71_3080 ();
 sg13g2_decap_8 FILLER_71_3087 ();
 sg13g2_decap_8 FILLER_71_3094 ();
 sg13g2_decap_8 FILLER_71_3101 ();
 sg13g2_decap_8 FILLER_71_3108 ();
 sg13g2_decap_8 FILLER_71_3115 ();
 sg13g2_decap_8 FILLER_71_3122 ();
 sg13g2_decap_8 FILLER_71_3129 ();
 sg13g2_decap_8 FILLER_71_3136 ();
 sg13g2_decap_8 FILLER_71_3143 ();
 sg13g2_decap_8 FILLER_71_3150 ();
 sg13g2_decap_8 FILLER_71_3157 ();
 sg13g2_decap_8 FILLER_71_3164 ();
 sg13g2_decap_8 FILLER_71_3171 ();
 sg13g2_decap_8 FILLER_71_3178 ();
 sg13g2_decap_8 FILLER_71_3185 ();
 sg13g2_decap_8 FILLER_71_3192 ();
 sg13g2_decap_8 FILLER_71_3199 ();
 sg13g2_decap_8 FILLER_71_3206 ();
 sg13g2_decap_8 FILLER_71_3213 ();
 sg13g2_decap_8 FILLER_71_3220 ();
 sg13g2_decap_8 FILLER_71_3227 ();
 sg13g2_decap_8 FILLER_71_3234 ();
 sg13g2_decap_8 FILLER_71_3241 ();
 sg13g2_decap_8 FILLER_71_3248 ();
 sg13g2_decap_8 FILLER_71_3255 ();
 sg13g2_decap_8 FILLER_71_3262 ();
 sg13g2_decap_8 FILLER_71_3269 ();
 sg13g2_decap_8 FILLER_71_3276 ();
 sg13g2_decap_8 FILLER_71_3283 ();
 sg13g2_decap_8 FILLER_71_3290 ();
 sg13g2_decap_8 FILLER_71_3297 ();
 sg13g2_decap_8 FILLER_71_3304 ();
 sg13g2_decap_8 FILLER_71_3311 ();
 sg13g2_decap_8 FILLER_71_3318 ();
 sg13g2_decap_8 FILLER_71_3325 ();
 sg13g2_decap_8 FILLER_71_3332 ();
 sg13g2_decap_8 FILLER_71_3339 ();
 sg13g2_decap_8 FILLER_71_3346 ();
 sg13g2_decap_8 FILLER_71_3353 ();
 sg13g2_decap_8 FILLER_71_3360 ();
 sg13g2_decap_8 FILLER_71_3367 ();
 sg13g2_decap_8 FILLER_71_3374 ();
 sg13g2_decap_8 FILLER_71_3381 ();
 sg13g2_decap_8 FILLER_71_3388 ();
 sg13g2_decap_8 FILLER_71_3395 ();
 sg13g2_decap_8 FILLER_71_3402 ();
 sg13g2_decap_8 FILLER_71_3409 ();
 sg13g2_decap_8 FILLER_71_3416 ();
 sg13g2_decap_8 FILLER_71_3423 ();
 sg13g2_decap_8 FILLER_71_3430 ();
 sg13g2_decap_8 FILLER_71_3437 ();
 sg13g2_decap_8 FILLER_71_3444 ();
 sg13g2_decap_8 FILLER_71_3451 ();
 sg13g2_decap_8 FILLER_71_3458 ();
 sg13g2_decap_8 FILLER_71_3465 ();
 sg13g2_decap_8 FILLER_71_3472 ();
 sg13g2_decap_8 FILLER_71_3479 ();
 sg13g2_decap_8 FILLER_71_3486 ();
 sg13g2_decap_8 FILLER_71_3493 ();
 sg13g2_decap_8 FILLER_71_3500 ();
 sg13g2_decap_8 FILLER_71_3507 ();
 sg13g2_decap_8 FILLER_71_3514 ();
 sg13g2_decap_8 FILLER_71_3521 ();
 sg13g2_decap_8 FILLER_71_3528 ();
 sg13g2_decap_8 FILLER_71_3535 ();
 sg13g2_decap_8 FILLER_71_3542 ();
 sg13g2_decap_8 FILLER_71_3549 ();
 sg13g2_decap_8 FILLER_71_3556 ();
 sg13g2_decap_8 FILLER_71_3563 ();
 sg13g2_decap_8 FILLER_71_3570 ();
 sg13g2_fill_2 FILLER_71_3577 ();
 sg13g2_fill_1 FILLER_71_3579 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_decap_8 FILLER_72_140 ();
 sg13g2_decap_8 FILLER_72_147 ();
 sg13g2_fill_2 FILLER_72_154 ();
 sg13g2_fill_1 FILLER_72_184 ();
 sg13g2_fill_1 FILLER_72_208 ();
 sg13g2_fill_2 FILLER_72_214 ();
 sg13g2_fill_1 FILLER_72_216 ();
 sg13g2_fill_2 FILLER_72_234 ();
 sg13g2_fill_1 FILLER_72_246 ();
 sg13g2_decap_8 FILLER_72_282 ();
 sg13g2_decap_8 FILLER_72_289 ();
 sg13g2_decap_8 FILLER_72_296 ();
 sg13g2_decap_8 FILLER_72_303 ();
 sg13g2_decap_8 FILLER_72_310 ();
 sg13g2_decap_8 FILLER_72_317 ();
 sg13g2_decap_8 FILLER_72_324 ();
 sg13g2_decap_8 FILLER_72_331 ();
 sg13g2_decap_8 FILLER_72_338 ();
 sg13g2_decap_8 FILLER_72_345 ();
 sg13g2_decap_8 FILLER_72_352 ();
 sg13g2_decap_8 FILLER_72_359 ();
 sg13g2_decap_8 FILLER_72_366 ();
 sg13g2_decap_8 FILLER_72_373 ();
 sg13g2_decap_8 FILLER_72_380 ();
 sg13g2_decap_8 FILLER_72_387 ();
 sg13g2_decap_8 FILLER_72_394 ();
 sg13g2_decap_8 FILLER_72_401 ();
 sg13g2_decap_8 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_72_415 ();
 sg13g2_decap_8 FILLER_72_422 ();
 sg13g2_decap_8 FILLER_72_429 ();
 sg13g2_decap_8 FILLER_72_436 ();
 sg13g2_decap_8 FILLER_72_443 ();
 sg13g2_decap_8 FILLER_72_450 ();
 sg13g2_decap_8 FILLER_72_457 ();
 sg13g2_decap_8 FILLER_72_464 ();
 sg13g2_decap_8 FILLER_72_471 ();
 sg13g2_decap_8 FILLER_72_478 ();
 sg13g2_decap_8 FILLER_72_485 ();
 sg13g2_decap_8 FILLER_72_492 ();
 sg13g2_decap_8 FILLER_72_499 ();
 sg13g2_decap_8 FILLER_72_506 ();
 sg13g2_decap_8 FILLER_72_513 ();
 sg13g2_decap_8 FILLER_72_520 ();
 sg13g2_decap_8 FILLER_72_527 ();
 sg13g2_decap_8 FILLER_72_534 ();
 sg13g2_decap_8 FILLER_72_541 ();
 sg13g2_decap_8 FILLER_72_548 ();
 sg13g2_decap_8 FILLER_72_555 ();
 sg13g2_decap_8 FILLER_72_562 ();
 sg13g2_decap_8 FILLER_72_569 ();
 sg13g2_decap_8 FILLER_72_576 ();
 sg13g2_decap_8 FILLER_72_583 ();
 sg13g2_decap_8 FILLER_72_590 ();
 sg13g2_decap_8 FILLER_72_597 ();
 sg13g2_decap_8 FILLER_72_604 ();
 sg13g2_decap_8 FILLER_72_611 ();
 sg13g2_decap_8 FILLER_72_618 ();
 sg13g2_decap_8 FILLER_72_625 ();
 sg13g2_decap_8 FILLER_72_632 ();
 sg13g2_decap_8 FILLER_72_639 ();
 sg13g2_decap_8 FILLER_72_646 ();
 sg13g2_decap_8 FILLER_72_653 ();
 sg13g2_decap_8 FILLER_72_660 ();
 sg13g2_decap_8 FILLER_72_667 ();
 sg13g2_decap_8 FILLER_72_674 ();
 sg13g2_decap_8 FILLER_72_681 ();
 sg13g2_decap_8 FILLER_72_688 ();
 sg13g2_decap_8 FILLER_72_695 ();
 sg13g2_decap_8 FILLER_72_702 ();
 sg13g2_decap_8 FILLER_72_709 ();
 sg13g2_decap_8 FILLER_72_716 ();
 sg13g2_decap_8 FILLER_72_723 ();
 sg13g2_decap_8 FILLER_72_730 ();
 sg13g2_decap_8 FILLER_72_737 ();
 sg13g2_decap_8 FILLER_72_744 ();
 sg13g2_decap_8 FILLER_72_751 ();
 sg13g2_decap_8 FILLER_72_758 ();
 sg13g2_decap_8 FILLER_72_765 ();
 sg13g2_decap_8 FILLER_72_772 ();
 sg13g2_decap_8 FILLER_72_779 ();
 sg13g2_decap_8 FILLER_72_786 ();
 sg13g2_decap_8 FILLER_72_793 ();
 sg13g2_decap_8 FILLER_72_800 ();
 sg13g2_decap_8 FILLER_72_807 ();
 sg13g2_decap_8 FILLER_72_814 ();
 sg13g2_decap_8 FILLER_72_821 ();
 sg13g2_decap_8 FILLER_72_828 ();
 sg13g2_decap_8 FILLER_72_835 ();
 sg13g2_decap_8 FILLER_72_842 ();
 sg13g2_decap_8 FILLER_72_849 ();
 sg13g2_decap_8 FILLER_72_856 ();
 sg13g2_decap_8 FILLER_72_863 ();
 sg13g2_decap_8 FILLER_72_870 ();
 sg13g2_decap_8 FILLER_72_877 ();
 sg13g2_decap_8 FILLER_72_884 ();
 sg13g2_decap_8 FILLER_72_891 ();
 sg13g2_decap_8 FILLER_72_898 ();
 sg13g2_decap_8 FILLER_72_905 ();
 sg13g2_decap_8 FILLER_72_912 ();
 sg13g2_decap_8 FILLER_72_919 ();
 sg13g2_decap_8 FILLER_72_926 ();
 sg13g2_decap_8 FILLER_72_933 ();
 sg13g2_decap_8 FILLER_72_940 ();
 sg13g2_decap_8 FILLER_72_947 ();
 sg13g2_decap_8 FILLER_72_954 ();
 sg13g2_decap_8 FILLER_72_961 ();
 sg13g2_decap_8 FILLER_72_968 ();
 sg13g2_decap_8 FILLER_72_975 ();
 sg13g2_decap_8 FILLER_72_982 ();
 sg13g2_decap_8 FILLER_72_989 ();
 sg13g2_decap_8 FILLER_72_996 ();
 sg13g2_decap_8 FILLER_72_1003 ();
 sg13g2_decap_8 FILLER_72_1010 ();
 sg13g2_decap_8 FILLER_72_1017 ();
 sg13g2_decap_8 FILLER_72_1024 ();
 sg13g2_decap_8 FILLER_72_1031 ();
 sg13g2_decap_8 FILLER_72_1038 ();
 sg13g2_decap_8 FILLER_72_1045 ();
 sg13g2_decap_8 FILLER_72_1052 ();
 sg13g2_decap_8 FILLER_72_1059 ();
 sg13g2_decap_8 FILLER_72_1066 ();
 sg13g2_decap_8 FILLER_72_1073 ();
 sg13g2_decap_8 FILLER_72_1080 ();
 sg13g2_decap_8 FILLER_72_1087 ();
 sg13g2_decap_8 FILLER_72_1094 ();
 sg13g2_decap_8 FILLER_72_1101 ();
 sg13g2_decap_8 FILLER_72_1108 ();
 sg13g2_decap_8 FILLER_72_1115 ();
 sg13g2_decap_8 FILLER_72_1122 ();
 sg13g2_decap_8 FILLER_72_1129 ();
 sg13g2_decap_8 FILLER_72_1136 ();
 sg13g2_decap_8 FILLER_72_1143 ();
 sg13g2_decap_8 FILLER_72_1150 ();
 sg13g2_decap_8 FILLER_72_1157 ();
 sg13g2_decap_8 FILLER_72_1164 ();
 sg13g2_decap_8 FILLER_72_1171 ();
 sg13g2_decap_8 FILLER_72_1178 ();
 sg13g2_decap_8 FILLER_72_1185 ();
 sg13g2_decap_8 FILLER_72_1192 ();
 sg13g2_decap_8 FILLER_72_1199 ();
 sg13g2_decap_8 FILLER_72_1206 ();
 sg13g2_decap_8 FILLER_72_1213 ();
 sg13g2_decap_8 FILLER_72_1220 ();
 sg13g2_decap_8 FILLER_72_1227 ();
 sg13g2_decap_8 FILLER_72_1234 ();
 sg13g2_decap_8 FILLER_72_1241 ();
 sg13g2_decap_8 FILLER_72_1248 ();
 sg13g2_decap_8 FILLER_72_1255 ();
 sg13g2_decap_8 FILLER_72_1262 ();
 sg13g2_decap_8 FILLER_72_1269 ();
 sg13g2_decap_8 FILLER_72_1276 ();
 sg13g2_decap_8 FILLER_72_1283 ();
 sg13g2_decap_8 FILLER_72_1290 ();
 sg13g2_decap_8 FILLER_72_1297 ();
 sg13g2_decap_8 FILLER_72_1304 ();
 sg13g2_decap_8 FILLER_72_1311 ();
 sg13g2_decap_8 FILLER_72_1318 ();
 sg13g2_decap_8 FILLER_72_1325 ();
 sg13g2_decap_8 FILLER_72_1332 ();
 sg13g2_decap_8 FILLER_72_1339 ();
 sg13g2_decap_8 FILLER_72_1346 ();
 sg13g2_decap_8 FILLER_72_1353 ();
 sg13g2_decap_8 FILLER_72_1360 ();
 sg13g2_decap_8 FILLER_72_1367 ();
 sg13g2_decap_8 FILLER_72_1374 ();
 sg13g2_decap_8 FILLER_72_1381 ();
 sg13g2_decap_8 FILLER_72_1388 ();
 sg13g2_decap_8 FILLER_72_1395 ();
 sg13g2_decap_8 FILLER_72_1402 ();
 sg13g2_decap_8 FILLER_72_1409 ();
 sg13g2_decap_8 FILLER_72_1416 ();
 sg13g2_decap_8 FILLER_72_1423 ();
 sg13g2_decap_8 FILLER_72_1430 ();
 sg13g2_decap_8 FILLER_72_1437 ();
 sg13g2_decap_8 FILLER_72_1444 ();
 sg13g2_decap_8 FILLER_72_1451 ();
 sg13g2_decap_8 FILLER_72_1458 ();
 sg13g2_decap_8 FILLER_72_1465 ();
 sg13g2_decap_8 FILLER_72_1472 ();
 sg13g2_decap_8 FILLER_72_1479 ();
 sg13g2_decap_8 FILLER_72_1486 ();
 sg13g2_decap_8 FILLER_72_1493 ();
 sg13g2_decap_8 FILLER_72_1500 ();
 sg13g2_decap_8 FILLER_72_1507 ();
 sg13g2_decap_8 FILLER_72_1514 ();
 sg13g2_decap_8 FILLER_72_1521 ();
 sg13g2_decap_8 FILLER_72_1528 ();
 sg13g2_decap_8 FILLER_72_1535 ();
 sg13g2_decap_8 FILLER_72_1542 ();
 sg13g2_decap_8 FILLER_72_1549 ();
 sg13g2_decap_8 FILLER_72_1556 ();
 sg13g2_decap_8 FILLER_72_1563 ();
 sg13g2_decap_8 FILLER_72_1570 ();
 sg13g2_decap_8 FILLER_72_1577 ();
 sg13g2_decap_8 FILLER_72_1584 ();
 sg13g2_decap_8 FILLER_72_1591 ();
 sg13g2_decap_8 FILLER_72_1598 ();
 sg13g2_decap_8 FILLER_72_1605 ();
 sg13g2_decap_8 FILLER_72_1612 ();
 sg13g2_decap_8 FILLER_72_1619 ();
 sg13g2_decap_8 FILLER_72_1626 ();
 sg13g2_decap_8 FILLER_72_1633 ();
 sg13g2_decap_8 FILLER_72_1640 ();
 sg13g2_decap_8 FILLER_72_1647 ();
 sg13g2_decap_8 FILLER_72_1654 ();
 sg13g2_decap_8 FILLER_72_1661 ();
 sg13g2_decap_8 FILLER_72_1668 ();
 sg13g2_decap_8 FILLER_72_1675 ();
 sg13g2_decap_8 FILLER_72_1682 ();
 sg13g2_decap_8 FILLER_72_1689 ();
 sg13g2_decap_8 FILLER_72_1696 ();
 sg13g2_decap_8 FILLER_72_1703 ();
 sg13g2_decap_8 FILLER_72_1710 ();
 sg13g2_decap_8 FILLER_72_1717 ();
 sg13g2_decap_8 FILLER_72_1724 ();
 sg13g2_decap_8 FILLER_72_1731 ();
 sg13g2_decap_8 FILLER_72_1738 ();
 sg13g2_decap_8 FILLER_72_1745 ();
 sg13g2_decap_8 FILLER_72_1752 ();
 sg13g2_decap_8 FILLER_72_1759 ();
 sg13g2_decap_8 FILLER_72_1766 ();
 sg13g2_decap_8 FILLER_72_1773 ();
 sg13g2_decap_8 FILLER_72_1780 ();
 sg13g2_decap_8 FILLER_72_1787 ();
 sg13g2_decap_8 FILLER_72_1794 ();
 sg13g2_decap_8 FILLER_72_1801 ();
 sg13g2_decap_8 FILLER_72_1808 ();
 sg13g2_decap_8 FILLER_72_1815 ();
 sg13g2_decap_8 FILLER_72_1822 ();
 sg13g2_decap_8 FILLER_72_1829 ();
 sg13g2_decap_8 FILLER_72_1836 ();
 sg13g2_decap_8 FILLER_72_1843 ();
 sg13g2_decap_8 FILLER_72_1850 ();
 sg13g2_decap_8 FILLER_72_1857 ();
 sg13g2_decap_8 FILLER_72_1864 ();
 sg13g2_decap_8 FILLER_72_1871 ();
 sg13g2_decap_8 FILLER_72_1878 ();
 sg13g2_decap_8 FILLER_72_1885 ();
 sg13g2_decap_8 FILLER_72_1892 ();
 sg13g2_decap_8 FILLER_72_1899 ();
 sg13g2_decap_8 FILLER_72_1906 ();
 sg13g2_decap_8 FILLER_72_1913 ();
 sg13g2_decap_8 FILLER_72_1920 ();
 sg13g2_decap_8 FILLER_72_1927 ();
 sg13g2_decap_8 FILLER_72_1934 ();
 sg13g2_decap_8 FILLER_72_1941 ();
 sg13g2_decap_8 FILLER_72_1948 ();
 sg13g2_decap_8 FILLER_72_1955 ();
 sg13g2_decap_8 FILLER_72_1962 ();
 sg13g2_decap_8 FILLER_72_1969 ();
 sg13g2_decap_8 FILLER_72_1976 ();
 sg13g2_decap_8 FILLER_72_1983 ();
 sg13g2_decap_8 FILLER_72_1990 ();
 sg13g2_decap_8 FILLER_72_1997 ();
 sg13g2_decap_8 FILLER_72_2004 ();
 sg13g2_decap_8 FILLER_72_2011 ();
 sg13g2_decap_8 FILLER_72_2018 ();
 sg13g2_decap_8 FILLER_72_2025 ();
 sg13g2_decap_8 FILLER_72_2032 ();
 sg13g2_decap_8 FILLER_72_2039 ();
 sg13g2_decap_8 FILLER_72_2046 ();
 sg13g2_decap_8 FILLER_72_2053 ();
 sg13g2_decap_8 FILLER_72_2060 ();
 sg13g2_decap_8 FILLER_72_2067 ();
 sg13g2_decap_8 FILLER_72_2074 ();
 sg13g2_decap_8 FILLER_72_2081 ();
 sg13g2_decap_8 FILLER_72_2088 ();
 sg13g2_decap_8 FILLER_72_2095 ();
 sg13g2_decap_8 FILLER_72_2102 ();
 sg13g2_decap_8 FILLER_72_2109 ();
 sg13g2_decap_8 FILLER_72_2116 ();
 sg13g2_decap_8 FILLER_72_2123 ();
 sg13g2_decap_8 FILLER_72_2130 ();
 sg13g2_decap_8 FILLER_72_2137 ();
 sg13g2_decap_8 FILLER_72_2144 ();
 sg13g2_decap_8 FILLER_72_2151 ();
 sg13g2_decap_8 FILLER_72_2158 ();
 sg13g2_decap_8 FILLER_72_2165 ();
 sg13g2_decap_8 FILLER_72_2172 ();
 sg13g2_decap_8 FILLER_72_2179 ();
 sg13g2_decap_8 FILLER_72_2186 ();
 sg13g2_decap_8 FILLER_72_2193 ();
 sg13g2_decap_8 FILLER_72_2200 ();
 sg13g2_decap_8 FILLER_72_2207 ();
 sg13g2_decap_8 FILLER_72_2214 ();
 sg13g2_decap_8 FILLER_72_2221 ();
 sg13g2_decap_8 FILLER_72_2228 ();
 sg13g2_decap_8 FILLER_72_2235 ();
 sg13g2_decap_8 FILLER_72_2242 ();
 sg13g2_decap_8 FILLER_72_2249 ();
 sg13g2_decap_8 FILLER_72_2256 ();
 sg13g2_decap_8 FILLER_72_2263 ();
 sg13g2_decap_8 FILLER_72_2270 ();
 sg13g2_decap_8 FILLER_72_2277 ();
 sg13g2_decap_8 FILLER_72_2284 ();
 sg13g2_decap_8 FILLER_72_2291 ();
 sg13g2_decap_8 FILLER_72_2298 ();
 sg13g2_decap_8 FILLER_72_2305 ();
 sg13g2_decap_8 FILLER_72_2312 ();
 sg13g2_decap_8 FILLER_72_2319 ();
 sg13g2_decap_8 FILLER_72_2326 ();
 sg13g2_decap_8 FILLER_72_2333 ();
 sg13g2_decap_8 FILLER_72_2340 ();
 sg13g2_decap_8 FILLER_72_2347 ();
 sg13g2_decap_8 FILLER_72_2354 ();
 sg13g2_decap_8 FILLER_72_2361 ();
 sg13g2_decap_8 FILLER_72_2368 ();
 sg13g2_decap_8 FILLER_72_2375 ();
 sg13g2_decap_8 FILLER_72_2382 ();
 sg13g2_decap_8 FILLER_72_2389 ();
 sg13g2_decap_8 FILLER_72_2396 ();
 sg13g2_decap_8 FILLER_72_2403 ();
 sg13g2_decap_8 FILLER_72_2410 ();
 sg13g2_decap_8 FILLER_72_2417 ();
 sg13g2_decap_8 FILLER_72_2424 ();
 sg13g2_decap_8 FILLER_72_2431 ();
 sg13g2_decap_8 FILLER_72_2438 ();
 sg13g2_decap_8 FILLER_72_2445 ();
 sg13g2_decap_8 FILLER_72_2452 ();
 sg13g2_decap_8 FILLER_72_2459 ();
 sg13g2_decap_8 FILLER_72_2466 ();
 sg13g2_decap_8 FILLER_72_2473 ();
 sg13g2_decap_8 FILLER_72_2480 ();
 sg13g2_decap_8 FILLER_72_2487 ();
 sg13g2_decap_8 FILLER_72_2494 ();
 sg13g2_decap_8 FILLER_72_2501 ();
 sg13g2_decap_8 FILLER_72_2508 ();
 sg13g2_decap_8 FILLER_72_2515 ();
 sg13g2_decap_8 FILLER_72_2522 ();
 sg13g2_decap_8 FILLER_72_2529 ();
 sg13g2_decap_8 FILLER_72_2536 ();
 sg13g2_decap_8 FILLER_72_2543 ();
 sg13g2_decap_8 FILLER_72_2550 ();
 sg13g2_decap_8 FILLER_72_2557 ();
 sg13g2_decap_8 FILLER_72_2564 ();
 sg13g2_decap_8 FILLER_72_2571 ();
 sg13g2_decap_8 FILLER_72_2578 ();
 sg13g2_decap_8 FILLER_72_2585 ();
 sg13g2_decap_8 FILLER_72_2592 ();
 sg13g2_decap_8 FILLER_72_2599 ();
 sg13g2_decap_8 FILLER_72_2606 ();
 sg13g2_decap_8 FILLER_72_2613 ();
 sg13g2_decap_8 FILLER_72_2620 ();
 sg13g2_decap_8 FILLER_72_2627 ();
 sg13g2_decap_8 FILLER_72_2634 ();
 sg13g2_decap_8 FILLER_72_2641 ();
 sg13g2_decap_8 FILLER_72_2648 ();
 sg13g2_decap_8 FILLER_72_2655 ();
 sg13g2_decap_8 FILLER_72_2662 ();
 sg13g2_decap_8 FILLER_72_2669 ();
 sg13g2_decap_8 FILLER_72_2676 ();
 sg13g2_decap_8 FILLER_72_2683 ();
 sg13g2_decap_8 FILLER_72_2690 ();
 sg13g2_decap_8 FILLER_72_2697 ();
 sg13g2_decap_8 FILLER_72_2704 ();
 sg13g2_decap_8 FILLER_72_2711 ();
 sg13g2_decap_8 FILLER_72_2718 ();
 sg13g2_decap_8 FILLER_72_2725 ();
 sg13g2_decap_8 FILLER_72_2732 ();
 sg13g2_decap_8 FILLER_72_2739 ();
 sg13g2_decap_8 FILLER_72_2746 ();
 sg13g2_decap_8 FILLER_72_2753 ();
 sg13g2_decap_8 FILLER_72_2760 ();
 sg13g2_decap_8 FILLER_72_2767 ();
 sg13g2_decap_8 FILLER_72_2774 ();
 sg13g2_decap_8 FILLER_72_2781 ();
 sg13g2_decap_8 FILLER_72_2788 ();
 sg13g2_decap_8 FILLER_72_2795 ();
 sg13g2_decap_8 FILLER_72_2802 ();
 sg13g2_decap_8 FILLER_72_2809 ();
 sg13g2_decap_8 FILLER_72_2816 ();
 sg13g2_decap_8 FILLER_72_2823 ();
 sg13g2_decap_8 FILLER_72_2830 ();
 sg13g2_decap_8 FILLER_72_2837 ();
 sg13g2_decap_8 FILLER_72_2844 ();
 sg13g2_decap_8 FILLER_72_2851 ();
 sg13g2_decap_8 FILLER_72_2858 ();
 sg13g2_decap_8 FILLER_72_2865 ();
 sg13g2_decap_8 FILLER_72_2872 ();
 sg13g2_decap_8 FILLER_72_2879 ();
 sg13g2_decap_8 FILLER_72_2886 ();
 sg13g2_decap_8 FILLER_72_2893 ();
 sg13g2_decap_8 FILLER_72_2900 ();
 sg13g2_decap_8 FILLER_72_2907 ();
 sg13g2_decap_8 FILLER_72_2914 ();
 sg13g2_decap_8 FILLER_72_2921 ();
 sg13g2_decap_8 FILLER_72_2928 ();
 sg13g2_decap_8 FILLER_72_2935 ();
 sg13g2_decap_8 FILLER_72_2942 ();
 sg13g2_decap_8 FILLER_72_2949 ();
 sg13g2_decap_8 FILLER_72_2956 ();
 sg13g2_decap_8 FILLER_72_2963 ();
 sg13g2_decap_8 FILLER_72_2970 ();
 sg13g2_decap_8 FILLER_72_2977 ();
 sg13g2_decap_8 FILLER_72_2984 ();
 sg13g2_decap_8 FILLER_72_2991 ();
 sg13g2_decap_8 FILLER_72_2998 ();
 sg13g2_decap_8 FILLER_72_3005 ();
 sg13g2_decap_8 FILLER_72_3012 ();
 sg13g2_decap_8 FILLER_72_3019 ();
 sg13g2_decap_8 FILLER_72_3026 ();
 sg13g2_decap_8 FILLER_72_3033 ();
 sg13g2_decap_8 FILLER_72_3040 ();
 sg13g2_decap_8 FILLER_72_3047 ();
 sg13g2_decap_8 FILLER_72_3054 ();
 sg13g2_decap_8 FILLER_72_3061 ();
 sg13g2_decap_8 FILLER_72_3068 ();
 sg13g2_decap_8 FILLER_72_3075 ();
 sg13g2_decap_8 FILLER_72_3082 ();
 sg13g2_decap_8 FILLER_72_3089 ();
 sg13g2_decap_8 FILLER_72_3096 ();
 sg13g2_decap_8 FILLER_72_3103 ();
 sg13g2_decap_8 FILLER_72_3110 ();
 sg13g2_decap_8 FILLER_72_3117 ();
 sg13g2_decap_8 FILLER_72_3124 ();
 sg13g2_decap_8 FILLER_72_3131 ();
 sg13g2_decap_8 FILLER_72_3138 ();
 sg13g2_decap_8 FILLER_72_3145 ();
 sg13g2_decap_8 FILLER_72_3152 ();
 sg13g2_decap_8 FILLER_72_3159 ();
 sg13g2_decap_8 FILLER_72_3166 ();
 sg13g2_decap_8 FILLER_72_3173 ();
 sg13g2_decap_8 FILLER_72_3180 ();
 sg13g2_decap_8 FILLER_72_3187 ();
 sg13g2_decap_8 FILLER_72_3194 ();
 sg13g2_decap_8 FILLER_72_3201 ();
 sg13g2_decap_8 FILLER_72_3208 ();
 sg13g2_decap_8 FILLER_72_3215 ();
 sg13g2_decap_8 FILLER_72_3222 ();
 sg13g2_decap_8 FILLER_72_3229 ();
 sg13g2_decap_8 FILLER_72_3236 ();
 sg13g2_decap_8 FILLER_72_3243 ();
 sg13g2_decap_8 FILLER_72_3250 ();
 sg13g2_decap_8 FILLER_72_3257 ();
 sg13g2_decap_8 FILLER_72_3264 ();
 sg13g2_decap_8 FILLER_72_3271 ();
 sg13g2_decap_8 FILLER_72_3278 ();
 sg13g2_decap_8 FILLER_72_3285 ();
 sg13g2_decap_8 FILLER_72_3292 ();
 sg13g2_decap_8 FILLER_72_3299 ();
 sg13g2_decap_8 FILLER_72_3306 ();
 sg13g2_decap_8 FILLER_72_3313 ();
 sg13g2_decap_8 FILLER_72_3320 ();
 sg13g2_decap_8 FILLER_72_3327 ();
 sg13g2_decap_8 FILLER_72_3334 ();
 sg13g2_decap_8 FILLER_72_3341 ();
 sg13g2_decap_8 FILLER_72_3348 ();
 sg13g2_decap_8 FILLER_72_3355 ();
 sg13g2_decap_8 FILLER_72_3362 ();
 sg13g2_decap_8 FILLER_72_3369 ();
 sg13g2_decap_8 FILLER_72_3376 ();
 sg13g2_decap_8 FILLER_72_3383 ();
 sg13g2_decap_8 FILLER_72_3390 ();
 sg13g2_decap_8 FILLER_72_3397 ();
 sg13g2_decap_8 FILLER_72_3404 ();
 sg13g2_decap_8 FILLER_72_3411 ();
 sg13g2_decap_8 FILLER_72_3418 ();
 sg13g2_decap_8 FILLER_72_3425 ();
 sg13g2_decap_8 FILLER_72_3432 ();
 sg13g2_decap_8 FILLER_72_3439 ();
 sg13g2_decap_8 FILLER_72_3446 ();
 sg13g2_decap_8 FILLER_72_3453 ();
 sg13g2_decap_8 FILLER_72_3460 ();
 sg13g2_decap_8 FILLER_72_3467 ();
 sg13g2_decap_8 FILLER_72_3474 ();
 sg13g2_decap_8 FILLER_72_3481 ();
 sg13g2_decap_8 FILLER_72_3488 ();
 sg13g2_decap_8 FILLER_72_3495 ();
 sg13g2_decap_8 FILLER_72_3502 ();
 sg13g2_decap_8 FILLER_72_3509 ();
 sg13g2_decap_8 FILLER_72_3516 ();
 sg13g2_decap_8 FILLER_72_3523 ();
 sg13g2_decap_8 FILLER_72_3530 ();
 sg13g2_decap_8 FILLER_72_3537 ();
 sg13g2_decap_8 FILLER_72_3544 ();
 sg13g2_decap_8 FILLER_72_3551 ();
 sg13g2_decap_8 FILLER_72_3558 ();
 sg13g2_decap_8 FILLER_72_3565 ();
 sg13g2_decap_8 FILLER_72_3572 ();
 sg13g2_fill_1 FILLER_72_3579 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_8 FILLER_73_140 ();
 sg13g2_decap_8 FILLER_73_147 ();
 sg13g2_decap_8 FILLER_73_154 ();
 sg13g2_fill_2 FILLER_73_186 ();
 sg13g2_fill_1 FILLER_73_188 ();
 sg13g2_fill_1 FILLER_73_202 ();
 sg13g2_decap_8 FILLER_73_219 ();
 sg13g2_fill_2 FILLER_73_256 ();
 sg13g2_fill_2 FILLER_73_266 ();
 sg13g2_decap_8 FILLER_73_296 ();
 sg13g2_decap_8 FILLER_73_303 ();
 sg13g2_decap_8 FILLER_73_310 ();
 sg13g2_decap_8 FILLER_73_317 ();
 sg13g2_decap_8 FILLER_73_324 ();
 sg13g2_decap_8 FILLER_73_331 ();
 sg13g2_decap_8 FILLER_73_338 ();
 sg13g2_decap_8 FILLER_73_345 ();
 sg13g2_decap_8 FILLER_73_352 ();
 sg13g2_decap_8 FILLER_73_359 ();
 sg13g2_decap_8 FILLER_73_366 ();
 sg13g2_decap_8 FILLER_73_373 ();
 sg13g2_decap_8 FILLER_73_380 ();
 sg13g2_decap_8 FILLER_73_387 ();
 sg13g2_decap_8 FILLER_73_394 ();
 sg13g2_decap_8 FILLER_73_401 ();
 sg13g2_decap_8 FILLER_73_408 ();
 sg13g2_decap_8 FILLER_73_415 ();
 sg13g2_decap_8 FILLER_73_422 ();
 sg13g2_decap_8 FILLER_73_429 ();
 sg13g2_decap_8 FILLER_73_436 ();
 sg13g2_decap_8 FILLER_73_443 ();
 sg13g2_decap_8 FILLER_73_450 ();
 sg13g2_decap_8 FILLER_73_457 ();
 sg13g2_decap_8 FILLER_73_464 ();
 sg13g2_decap_8 FILLER_73_471 ();
 sg13g2_decap_8 FILLER_73_478 ();
 sg13g2_decap_8 FILLER_73_485 ();
 sg13g2_decap_8 FILLER_73_492 ();
 sg13g2_decap_8 FILLER_73_499 ();
 sg13g2_decap_8 FILLER_73_506 ();
 sg13g2_decap_8 FILLER_73_513 ();
 sg13g2_decap_8 FILLER_73_520 ();
 sg13g2_decap_8 FILLER_73_527 ();
 sg13g2_decap_8 FILLER_73_534 ();
 sg13g2_decap_8 FILLER_73_541 ();
 sg13g2_decap_8 FILLER_73_548 ();
 sg13g2_decap_8 FILLER_73_555 ();
 sg13g2_decap_8 FILLER_73_562 ();
 sg13g2_decap_8 FILLER_73_569 ();
 sg13g2_decap_8 FILLER_73_576 ();
 sg13g2_decap_8 FILLER_73_583 ();
 sg13g2_decap_8 FILLER_73_590 ();
 sg13g2_decap_8 FILLER_73_597 ();
 sg13g2_decap_8 FILLER_73_604 ();
 sg13g2_decap_8 FILLER_73_611 ();
 sg13g2_decap_8 FILLER_73_618 ();
 sg13g2_decap_8 FILLER_73_625 ();
 sg13g2_decap_8 FILLER_73_632 ();
 sg13g2_decap_8 FILLER_73_639 ();
 sg13g2_decap_8 FILLER_73_646 ();
 sg13g2_decap_8 FILLER_73_653 ();
 sg13g2_decap_8 FILLER_73_660 ();
 sg13g2_decap_8 FILLER_73_667 ();
 sg13g2_decap_8 FILLER_73_674 ();
 sg13g2_decap_8 FILLER_73_681 ();
 sg13g2_decap_8 FILLER_73_688 ();
 sg13g2_decap_8 FILLER_73_695 ();
 sg13g2_decap_8 FILLER_73_702 ();
 sg13g2_decap_8 FILLER_73_709 ();
 sg13g2_decap_8 FILLER_73_716 ();
 sg13g2_decap_8 FILLER_73_723 ();
 sg13g2_decap_8 FILLER_73_730 ();
 sg13g2_decap_8 FILLER_73_737 ();
 sg13g2_decap_8 FILLER_73_744 ();
 sg13g2_decap_8 FILLER_73_751 ();
 sg13g2_decap_8 FILLER_73_758 ();
 sg13g2_decap_8 FILLER_73_765 ();
 sg13g2_decap_8 FILLER_73_772 ();
 sg13g2_decap_8 FILLER_73_779 ();
 sg13g2_decap_8 FILLER_73_786 ();
 sg13g2_decap_8 FILLER_73_793 ();
 sg13g2_decap_8 FILLER_73_800 ();
 sg13g2_decap_8 FILLER_73_807 ();
 sg13g2_decap_8 FILLER_73_814 ();
 sg13g2_decap_8 FILLER_73_821 ();
 sg13g2_decap_8 FILLER_73_828 ();
 sg13g2_decap_8 FILLER_73_835 ();
 sg13g2_decap_8 FILLER_73_842 ();
 sg13g2_decap_8 FILLER_73_849 ();
 sg13g2_decap_8 FILLER_73_856 ();
 sg13g2_decap_8 FILLER_73_863 ();
 sg13g2_decap_8 FILLER_73_870 ();
 sg13g2_decap_8 FILLER_73_877 ();
 sg13g2_decap_8 FILLER_73_884 ();
 sg13g2_decap_8 FILLER_73_891 ();
 sg13g2_decap_8 FILLER_73_898 ();
 sg13g2_decap_8 FILLER_73_905 ();
 sg13g2_decap_8 FILLER_73_912 ();
 sg13g2_decap_8 FILLER_73_919 ();
 sg13g2_decap_8 FILLER_73_926 ();
 sg13g2_decap_8 FILLER_73_933 ();
 sg13g2_decap_8 FILLER_73_940 ();
 sg13g2_decap_8 FILLER_73_947 ();
 sg13g2_decap_8 FILLER_73_954 ();
 sg13g2_decap_8 FILLER_73_961 ();
 sg13g2_decap_8 FILLER_73_968 ();
 sg13g2_decap_8 FILLER_73_975 ();
 sg13g2_decap_8 FILLER_73_982 ();
 sg13g2_decap_8 FILLER_73_989 ();
 sg13g2_decap_8 FILLER_73_996 ();
 sg13g2_decap_8 FILLER_73_1003 ();
 sg13g2_decap_8 FILLER_73_1010 ();
 sg13g2_decap_8 FILLER_73_1017 ();
 sg13g2_decap_8 FILLER_73_1024 ();
 sg13g2_decap_8 FILLER_73_1031 ();
 sg13g2_decap_8 FILLER_73_1038 ();
 sg13g2_decap_8 FILLER_73_1045 ();
 sg13g2_decap_8 FILLER_73_1052 ();
 sg13g2_decap_8 FILLER_73_1059 ();
 sg13g2_decap_8 FILLER_73_1066 ();
 sg13g2_decap_8 FILLER_73_1073 ();
 sg13g2_decap_8 FILLER_73_1080 ();
 sg13g2_decap_8 FILLER_73_1087 ();
 sg13g2_decap_8 FILLER_73_1094 ();
 sg13g2_decap_8 FILLER_73_1101 ();
 sg13g2_decap_8 FILLER_73_1108 ();
 sg13g2_decap_8 FILLER_73_1115 ();
 sg13g2_decap_8 FILLER_73_1122 ();
 sg13g2_decap_8 FILLER_73_1129 ();
 sg13g2_decap_8 FILLER_73_1136 ();
 sg13g2_decap_8 FILLER_73_1143 ();
 sg13g2_decap_8 FILLER_73_1150 ();
 sg13g2_decap_8 FILLER_73_1157 ();
 sg13g2_decap_8 FILLER_73_1164 ();
 sg13g2_decap_8 FILLER_73_1171 ();
 sg13g2_decap_8 FILLER_73_1178 ();
 sg13g2_decap_8 FILLER_73_1185 ();
 sg13g2_decap_8 FILLER_73_1192 ();
 sg13g2_decap_8 FILLER_73_1199 ();
 sg13g2_decap_8 FILLER_73_1206 ();
 sg13g2_decap_8 FILLER_73_1213 ();
 sg13g2_decap_8 FILLER_73_1220 ();
 sg13g2_decap_8 FILLER_73_1227 ();
 sg13g2_decap_8 FILLER_73_1234 ();
 sg13g2_decap_8 FILLER_73_1241 ();
 sg13g2_decap_8 FILLER_73_1248 ();
 sg13g2_decap_8 FILLER_73_1255 ();
 sg13g2_decap_8 FILLER_73_1262 ();
 sg13g2_decap_8 FILLER_73_1269 ();
 sg13g2_decap_8 FILLER_73_1276 ();
 sg13g2_decap_8 FILLER_73_1283 ();
 sg13g2_decap_8 FILLER_73_1290 ();
 sg13g2_decap_8 FILLER_73_1297 ();
 sg13g2_decap_8 FILLER_73_1304 ();
 sg13g2_decap_8 FILLER_73_1311 ();
 sg13g2_decap_8 FILLER_73_1318 ();
 sg13g2_decap_8 FILLER_73_1325 ();
 sg13g2_decap_8 FILLER_73_1332 ();
 sg13g2_decap_8 FILLER_73_1339 ();
 sg13g2_decap_8 FILLER_73_1346 ();
 sg13g2_decap_8 FILLER_73_1353 ();
 sg13g2_decap_8 FILLER_73_1360 ();
 sg13g2_decap_8 FILLER_73_1367 ();
 sg13g2_decap_8 FILLER_73_1374 ();
 sg13g2_decap_8 FILLER_73_1381 ();
 sg13g2_decap_8 FILLER_73_1388 ();
 sg13g2_decap_8 FILLER_73_1395 ();
 sg13g2_decap_8 FILLER_73_1402 ();
 sg13g2_decap_8 FILLER_73_1409 ();
 sg13g2_decap_8 FILLER_73_1416 ();
 sg13g2_decap_8 FILLER_73_1423 ();
 sg13g2_decap_8 FILLER_73_1430 ();
 sg13g2_decap_8 FILLER_73_1437 ();
 sg13g2_decap_8 FILLER_73_1444 ();
 sg13g2_decap_8 FILLER_73_1451 ();
 sg13g2_decap_8 FILLER_73_1458 ();
 sg13g2_decap_8 FILLER_73_1465 ();
 sg13g2_decap_8 FILLER_73_1472 ();
 sg13g2_decap_8 FILLER_73_1479 ();
 sg13g2_decap_8 FILLER_73_1486 ();
 sg13g2_decap_8 FILLER_73_1493 ();
 sg13g2_decap_8 FILLER_73_1500 ();
 sg13g2_decap_8 FILLER_73_1507 ();
 sg13g2_decap_8 FILLER_73_1514 ();
 sg13g2_decap_8 FILLER_73_1521 ();
 sg13g2_decap_8 FILLER_73_1528 ();
 sg13g2_decap_8 FILLER_73_1535 ();
 sg13g2_decap_8 FILLER_73_1542 ();
 sg13g2_decap_8 FILLER_73_1549 ();
 sg13g2_decap_8 FILLER_73_1556 ();
 sg13g2_decap_8 FILLER_73_1563 ();
 sg13g2_decap_8 FILLER_73_1570 ();
 sg13g2_decap_8 FILLER_73_1577 ();
 sg13g2_decap_8 FILLER_73_1584 ();
 sg13g2_decap_8 FILLER_73_1591 ();
 sg13g2_decap_8 FILLER_73_1598 ();
 sg13g2_decap_8 FILLER_73_1605 ();
 sg13g2_decap_8 FILLER_73_1612 ();
 sg13g2_decap_8 FILLER_73_1619 ();
 sg13g2_decap_8 FILLER_73_1626 ();
 sg13g2_decap_8 FILLER_73_1633 ();
 sg13g2_decap_8 FILLER_73_1640 ();
 sg13g2_decap_8 FILLER_73_1647 ();
 sg13g2_decap_8 FILLER_73_1654 ();
 sg13g2_decap_8 FILLER_73_1661 ();
 sg13g2_decap_8 FILLER_73_1668 ();
 sg13g2_decap_8 FILLER_73_1675 ();
 sg13g2_decap_8 FILLER_73_1682 ();
 sg13g2_decap_8 FILLER_73_1689 ();
 sg13g2_decap_8 FILLER_73_1696 ();
 sg13g2_decap_8 FILLER_73_1703 ();
 sg13g2_decap_8 FILLER_73_1710 ();
 sg13g2_decap_8 FILLER_73_1717 ();
 sg13g2_decap_8 FILLER_73_1724 ();
 sg13g2_decap_8 FILLER_73_1731 ();
 sg13g2_decap_8 FILLER_73_1738 ();
 sg13g2_decap_8 FILLER_73_1745 ();
 sg13g2_decap_8 FILLER_73_1752 ();
 sg13g2_decap_8 FILLER_73_1759 ();
 sg13g2_decap_8 FILLER_73_1766 ();
 sg13g2_decap_8 FILLER_73_1773 ();
 sg13g2_decap_8 FILLER_73_1780 ();
 sg13g2_decap_8 FILLER_73_1787 ();
 sg13g2_decap_8 FILLER_73_1794 ();
 sg13g2_decap_8 FILLER_73_1801 ();
 sg13g2_decap_8 FILLER_73_1808 ();
 sg13g2_decap_8 FILLER_73_1815 ();
 sg13g2_decap_8 FILLER_73_1822 ();
 sg13g2_decap_8 FILLER_73_1829 ();
 sg13g2_decap_8 FILLER_73_1836 ();
 sg13g2_decap_8 FILLER_73_1843 ();
 sg13g2_decap_8 FILLER_73_1850 ();
 sg13g2_decap_8 FILLER_73_1857 ();
 sg13g2_decap_8 FILLER_73_1864 ();
 sg13g2_decap_8 FILLER_73_1871 ();
 sg13g2_decap_8 FILLER_73_1878 ();
 sg13g2_decap_8 FILLER_73_1885 ();
 sg13g2_decap_8 FILLER_73_1892 ();
 sg13g2_decap_8 FILLER_73_1899 ();
 sg13g2_decap_8 FILLER_73_1906 ();
 sg13g2_decap_8 FILLER_73_1913 ();
 sg13g2_decap_8 FILLER_73_1920 ();
 sg13g2_decap_8 FILLER_73_1927 ();
 sg13g2_decap_8 FILLER_73_1934 ();
 sg13g2_decap_8 FILLER_73_1941 ();
 sg13g2_decap_8 FILLER_73_1948 ();
 sg13g2_decap_8 FILLER_73_1955 ();
 sg13g2_decap_8 FILLER_73_1962 ();
 sg13g2_decap_8 FILLER_73_1969 ();
 sg13g2_decap_8 FILLER_73_1976 ();
 sg13g2_decap_8 FILLER_73_1983 ();
 sg13g2_decap_8 FILLER_73_1990 ();
 sg13g2_decap_8 FILLER_73_1997 ();
 sg13g2_decap_8 FILLER_73_2004 ();
 sg13g2_decap_8 FILLER_73_2011 ();
 sg13g2_decap_8 FILLER_73_2018 ();
 sg13g2_decap_8 FILLER_73_2025 ();
 sg13g2_decap_8 FILLER_73_2032 ();
 sg13g2_decap_8 FILLER_73_2039 ();
 sg13g2_decap_8 FILLER_73_2046 ();
 sg13g2_decap_8 FILLER_73_2053 ();
 sg13g2_decap_8 FILLER_73_2060 ();
 sg13g2_decap_8 FILLER_73_2067 ();
 sg13g2_decap_8 FILLER_73_2074 ();
 sg13g2_decap_8 FILLER_73_2081 ();
 sg13g2_decap_8 FILLER_73_2088 ();
 sg13g2_decap_8 FILLER_73_2095 ();
 sg13g2_decap_8 FILLER_73_2102 ();
 sg13g2_decap_8 FILLER_73_2109 ();
 sg13g2_decap_8 FILLER_73_2116 ();
 sg13g2_decap_8 FILLER_73_2123 ();
 sg13g2_decap_8 FILLER_73_2130 ();
 sg13g2_decap_8 FILLER_73_2137 ();
 sg13g2_decap_8 FILLER_73_2144 ();
 sg13g2_decap_8 FILLER_73_2151 ();
 sg13g2_decap_8 FILLER_73_2158 ();
 sg13g2_decap_8 FILLER_73_2165 ();
 sg13g2_decap_8 FILLER_73_2172 ();
 sg13g2_decap_8 FILLER_73_2179 ();
 sg13g2_decap_8 FILLER_73_2186 ();
 sg13g2_decap_8 FILLER_73_2193 ();
 sg13g2_decap_8 FILLER_73_2200 ();
 sg13g2_decap_8 FILLER_73_2207 ();
 sg13g2_decap_8 FILLER_73_2214 ();
 sg13g2_decap_8 FILLER_73_2221 ();
 sg13g2_decap_8 FILLER_73_2228 ();
 sg13g2_decap_8 FILLER_73_2235 ();
 sg13g2_decap_8 FILLER_73_2242 ();
 sg13g2_decap_8 FILLER_73_2249 ();
 sg13g2_decap_8 FILLER_73_2256 ();
 sg13g2_decap_8 FILLER_73_2263 ();
 sg13g2_decap_8 FILLER_73_2270 ();
 sg13g2_decap_8 FILLER_73_2277 ();
 sg13g2_decap_8 FILLER_73_2284 ();
 sg13g2_decap_8 FILLER_73_2291 ();
 sg13g2_decap_8 FILLER_73_2298 ();
 sg13g2_decap_8 FILLER_73_2305 ();
 sg13g2_decap_8 FILLER_73_2312 ();
 sg13g2_decap_8 FILLER_73_2319 ();
 sg13g2_decap_8 FILLER_73_2326 ();
 sg13g2_decap_8 FILLER_73_2333 ();
 sg13g2_decap_8 FILLER_73_2340 ();
 sg13g2_decap_8 FILLER_73_2347 ();
 sg13g2_decap_8 FILLER_73_2354 ();
 sg13g2_decap_8 FILLER_73_2361 ();
 sg13g2_decap_8 FILLER_73_2368 ();
 sg13g2_decap_8 FILLER_73_2375 ();
 sg13g2_decap_8 FILLER_73_2382 ();
 sg13g2_decap_8 FILLER_73_2389 ();
 sg13g2_decap_8 FILLER_73_2396 ();
 sg13g2_decap_8 FILLER_73_2403 ();
 sg13g2_decap_8 FILLER_73_2410 ();
 sg13g2_decap_8 FILLER_73_2417 ();
 sg13g2_decap_8 FILLER_73_2424 ();
 sg13g2_decap_8 FILLER_73_2431 ();
 sg13g2_decap_8 FILLER_73_2438 ();
 sg13g2_decap_8 FILLER_73_2445 ();
 sg13g2_decap_8 FILLER_73_2452 ();
 sg13g2_decap_8 FILLER_73_2459 ();
 sg13g2_decap_8 FILLER_73_2466 ();
 sg13g2_decap_8 FILLER_73_2473 ();
 sg13g2_decap_8 FILLER_73_2480 ();
 sg13g2_decap_8 FILLER_73_2487 ();
 sg13g2_decap_8 FILLER_73_2494 ();
 sg13g2_decap_8 FILLER_73_2501 ();
 sg13g2_decap_8 FILLER_73_2508 ();
 sg13g2_decap_8 FILLER_73_2515 ();
 sg13g2_decap_8 FILLER_73_2522 ();
 sg13g2_decap_8 FILLER_73_2529 ();
 sg13g2_decap_8 FILLER_73_2536 ();
 sg13g2_decap_8 FILLER_73_2543 ();
 sg13g2_decap_8 FILLER_73_2550 ();
 sg13g2_decap_8 FILLER_73_2557 ();
 sg13g2_decap_8 FILLER_73_2564 ();
 sg13g2_decap_8 FILLER_73_2571 ();
 sg13g2_decap_8 FILLER_73_2578 ();
 sg13g2_decap_8 FILLER_73_2585 ();
 sg13g2_decap_8 FILLER_73_2592 ();
 sg13g2_decap_8 FILLER_73_2599 ();
 sg13g2_decap_8 FILLER_73_2606 ();
 sg13g2_decap_8 FILLER_73_2613 ();
 sg13g2_decap_8 FILLER_73_2620 ();
 sg13g2_decap_8 FILLER_73_2627 ();
 sg13g2_decap_8 FILLER_73_2634 ();
 sg13g2_decap_8 FILLER_73_2641 ();
 sg13g2_decap_8 FILLER_73_2648 ();
 sg13g2_decap_8 FILLER_73_2655 ();
 sg13g2_decap_8 FILLER_73_2662 ();
 sg13g2_decap_8 FILLER_73_2669 ();
 sg13g2_decap_8 FILLER_73_2676 ();
 sg13g2_decap_8 FILLER_73_2683 ();
 sg13g2_decap_8 FILLER_73_2690 ();
 sg13g2_decap_8 FILLER_73_2697 ();
 sg13g2_decap_8 FILLER_73_2704 ();
 sg13g2_decap_8 FILLER_73_2711 ();
 sg13g2_decap_8 FILLER_73_2718 ();
 sg13g2_decap_8 FILLER_73_2725 ();
 sg13g2_decap_8 FILLER_73_2732 ();
 sg13g2_decap_8 FILLER_73_2739 ();
 sg13g2_decap_8 FILLER_73_2746 ();
 sg13g2_decap_8 FILLER_73_2753 ();
 sg13g2_decap_8 FILLER_73_2760 ();
 sg13g2_decap_8 FILLER_73_2767 ();
 sg13g2_decap_8 FILLER_73_2774 ();
 sg13g2_decap_8 FILLER_73_2781 ();
 sg13g2_decap_8 FILLER_73_2788 ();
 sg13g2_decap_8 FILLER_73_2795 ();
 sg13g2_decap_8 FILLER_73_2802 ();
 sg13g2_decap_8 FILLER_73_2809 ();
 sg13g2_decap_8 FILLER_73_2816 ();
 sg13g2_decap_8 FILLER_73_2823 ();
 sg13g2_decap_8 FILLER_73_2830 ();
 sg13g2_decap_8 FILLER_73_2837 ();
 sg13g2_decap_8 FILLER_73_2844 ();
 sg13g2_decap_8 FILLER_73_2851 ();
 sg13g2_decap_8 FILLER_73_2858 ();
 sg13g2_decap_8 FILLER_73_2865 ();
 sg13g2_decap_8 FILLER_73_2872 ();
 sg13g2_decap_8 FILLER_73_2879 ();
 sg13g2_decap_8 FILLER_73_2886 ();
 sg13g2_decap_8 FILLER_73_2893 ();
 sg13g2_decap_8 FILLER_73_2900 ();
 sg13g2_decap_8 FILLER_73_2907 ();
 sg13g2_decap_8 FILLER_73_2914 ();
 sg13g2_decap_8 FILLER_73_2921 ();
 sg13g2_decap_8 FILLER_73_2928 ();
 sg13g2_decap_8 FILLER_73_2935 ();
 sg13g2_decap_8 FILLER_73_2942 ();
 sg13g2_decap_8 FILLER_73_2949 ();
 sg13g2_decap_8 FILLER_73_2956 ();
 sg13g2_decap_8 FILLER_73_2963 ();
 sg13g2_decap_8 FILLER_73_2970 ();
 sg13g2_decap_8 FILLER_73_2977 ();
 sg13g2_decap_8 FILLER_73_2984 ();
 sg13g2_decap_8 FILLER_73_2991 ();
 sg13g2_decap_8 FILLER_73_2998 ();
 sg13g2_decap_8 FILLER_73_3005 ();
 sg13g2_decap_8 FILLER_73_3012 ();
 sg13g2_decap_8 FILLER_73_3019 ();
 sg13g2_decap_8 FILLER_73_3026 ();
 sg13g2_decap_8 FILLER_73_3033 ();
 sg13g2_decap_8 FILLER_73_3040 ();
 sg13g2_decap_8 FILLER_73_3047 ();
 sg13g2_decap_8 FILLER_73_3054 ();
 sg13g2_decap_8 FILLER_73_3061 ();
 sg13g2_decap_8 FILLER_73_3068 ();
 sg13g2_decap_8 FILLER_73_3075 ();
 sg13g2_decap_8 FILLER_73_3082 ();
 sg13g2_decap_8 FILLER_73_3089 ();
 sg13g2_decap_8 FILLER_73_3096 ();
 sg13g2_decap_8 FILLER_73_3103 ();
 sg13g2_decap_8 FILLER_73_3110 ();
 sg13g2_decap_8 FILLER_73_3117 ();
 sg13g2_decap_8 FILLER_73_3124 ();
 sg13g2_decap_8 FILLER_73_3131 ();
 sg13g2_decap_8 FILLER_73_3138 ();
 sg13g2_decap_8 FILLER_73_3145 ();
 sg13g2_decap_8 FILLER_73_3152 ();
 sg13g2_decap_8 FILLER_73_3159 ();
 sg13g2_decap_8 FILLER_73_3166 ();
 sg13g2_decap_8 FILLER_73_3173 ();
 sg13g2_decap_8 FILLER_73_3180 ();
 sg13g2_decap_8 FILLER_73_3187 ();
 sg13g2_decap_8 FILLER_73_3194 ();
 sg13g2_decap_8 FILLER_73_3201 ();
 sg13g2_decap_8 FILLER_73_3208 ();
 sg13g2_decap_8 FILLER_73_3215 ();
 sg13g2_decap_8 FILLER_73_3222 ();
 sg13g2_decap_8 FILLER_73_3229 ();
 sg13g2_decap_8 FILLER_73_3236 ();
 sg13g2_decap_8 FILLER_73_3243 ();
 sg13g2_decap_8 FILLER_73_3250 ();
 sg13g2_decap_8 FILLER_73_3257 ();
 sg13g2_decap_8 FILLER_73_3264 ();
 sg13g2_decap_8 FILLER_73_3271 ();
 sg13g2_decap_8 FILLER_73_3278 ();
 sg13g2_decap_8 FILLER_73_3285 ();
 sg13g2_decap_8 FILLER_73_3292 ();
 sg13g2_decap_8 FILLER_73_3299 ();
 sg13g2_decap_8 FILLER_73_3306 ();
 sg13g2_decap_8 FILLER_73_3313 ();
 sg13g2_decap_8 FILLER_73_3320 ();
 sg13g2_decap_8 FILLER_73_3327 ();
 sg13g2_decap_8 FILLER_73_3334 ();
 sg13g2_decap_8 FILLER_73_3341 ();
 sg13g2_decap_8 FILLER_73_3348 ();
 sg13g2_decap_8 FILLER_73_3355 ();
 sg13g2_decap_8 FILLER_73_3362 ();
 sg13g2_decap_8 FILLER_73_3369 ();
 sg13g2_decap_8 FILLER_73_3376 ();
 sg13g2_decap_8 FILLER_73_3383 ();
 sg13g2_decap_8 FILLER_73_3390 ();
 sg13g2_decap_8 FILLER_73_3397 ();
 sg13g2_decap_8 FILLER_73_3404 ();
 sg13g2_decap_8 FILLER_73_3411 ();
 sg13g2_decap_8 FILLER_73_3418 ();
 sg13g2_decap_8 FILLER_73_3425 ();
 sg13g2_decap_8 FILLER_73_3432 ();
 sg13g2_decap_8 FILLER_73_3439 ();
 sg13g2_decap_8 FILLER_73_3446 ();
 sg13g2_decap_8 FILLER_73_3453 ();
 sg13g2_decap_8 FILLER_73_3460 ();
 sg13g2_decap_8 FILLER_73_3467 ();
 sg13g2_decap_8 FILLER_73_3474 ();
 sg13g2_decap_8 FILLER_73_3481 ();
 sg13g2_decap_8 FILLER_73_3488 ();
 sg13g2_decap_8 FILLER_73_3495 ();
 sg13g2_decap_8 FILLER_73_3502 ();
 sg13g2_decap_8 FILLER_73_3509 ();
 sg13g2_decap_8 FILLER_73_3516 ();
 sg13g2_decap_8 FILLER_73_3523 ();
 sg13g2_decap_8 FILLER_73_3530 ();
 sg13g2_decap_8 FILLER_73_3537 ();
 sg13g2_decap_8 FILLER_73_3544 ();
 sg13g2_decap_8 FILLER_73_3551 ();
 sg13g2_decap_8 FILLER_73_3558 ();
 sg13g2_decap_8 FILLER_73_3565 ();
 sg13g2_decap_8 FILLER_73_3572 ();
 sg13g2_fill_1 FILLER_73_3579 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_8 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_147 ();
 sg13g2_decap_8 FILLER_74_154 ();
 sg13g2_fill_1 FILLER_74_161 ();
 sg13g2_decap_8 FILLER_74_217 ();
 sg13g2_decap_4 FILLER_74_224 ();
 sg13g2_fill_1 FILLER_74_246 ();
 sg13g2_decap_8 FILLER_74_269 ();
 sg13g2_fill_2 FILLER_74_276 ();
 sg13g2_decap_8 FILLER_74_287 ();
 sg13g2_decap_8 FILLER_74_294 ();
 sg13g2_decap_8 FILLER_74_301 ();
 sg13g2_decap_8 FILLER_74_308 ();
 sg13g2_decap_8 FILLER_74_315 ();
 sg13g2_decap_8 FILLER_74_322 ();
 sg13g2_decap_8 FILLER_74_329 ();
 sg13g2_decap_8 FILLER_74_336 ();
 sg13g2_decap_8 FILLER_74_343 ();
 sg13g2_decap_8 FILLER_74_350 ();
 sg13g2_decap_8 FILLER_74_357 ();
 sg13g2_decap_8 FILLER_74_364 ();
 sg13g2_decap_8 FILLER_74_371 ();
 sg13g2_decap_8 FILLER_74_378 ();
 sg13g2_decap_8 FILLER_74_385 ();
 sg13g2_decap_8 FILLER_74_392 ();
 sg13g2_decap_8 FILLER_74_399 ();
 sg13g2_decap_8 FILLER_74_406 ();
 sg13g2_decap_8 FILLER_74_413 ();
 sg13g2_decap_8 FILLER_74_420 ();
 sg13g2_decap_8 FILLER_74_427 ();
 sg13g2_decap_8 FILLER_74_434 ();
 sg13g2_decap_8 FILLER_74_441 ();
 sg13g2_decap_8 FILLER_74_448 ();
 sg13g2_decap_8 FILLER_74_455 ();
 sg13g2_decap_8 FILLER_74_462 ();
 sg13g2_decap_8 FILLER_74_469 ();
 sg13g2_decap_8 FILLER_74_476 ();
 sg13g2_decap_8 FILLER_74_483 ();
 sg13g2_decap_8 FILLER_74_490 ();
 sg13g2_decap_8 FILLER_74_497 ();
 sg13g2_decap_8 FILLER_74_504 ();
 sg13g2_decap_8 FILLER_74_511 ();
 sg13g2_decap_8 FILLER_74_518 ();
 sg13g2_decap_8 FILLER_74_525 ();
 sg13g2_decap_8 FILLER_74_532 ();
 sg13g2_decap_8 FILLER_74_539 ();
 sg13g2_decap_8 FILLER_74_546 ();
 sg13g2_decap_8 FILLER_74_553 ();
 sg13g2_decap_8 FILLER_74_560 ();
 sg13g2_decap_8 FILLER_74_567 ();
 sg13g2_decap_8 FILLER_74_574 ();
 sg13g2_decap_8 FILLER_74_581 ();
 sg13g2_decap_8 FILLER_74_588 ();
 sg13g2_decap_8 FILLER_74_595 ();
 sg13g2_decap_8 FILLER_74_602 ();
 sg13g2_decap_8 FILLER_74_609 ();
 sg13g2_decap_8 FILLER_74_616 ();
 sg13g2_decap_8 FILLER_74_623 ();
 sg13g2_decap_8 FILLER_74_630 ();
 sg13g2_decap_8 FILLER_74_637 ();
 sg13g2_decap_8 FILLER_74_644 ();
 sg13g2_decap_8 FILLER_74_651 ();
 sg13g2_decap_8 FILLER_74_658 ();
 sg13g2_decap_8 FILLER_74_665 ();
 sg13g2_decap_8 FILLER_74_672 ();
 sg13g2_decap_8 FILLER_74_679 ();
 sg13g2_decap_8 FILLER_74_686 ();
 sg13g2_decap_8 FILLER_74_693 ();
 sg13g2_decap_8 FILLER_74_700 ();
 sg13g2_decap_8 FILLER_74_707 ();
 sg13g2_decap_8 FILLER_74_714 ();
 sg13g2_decap_8 FILLER_74_721 ();
 sg13g2_decap_8 FILLER_74_728 ();
 sg13g2_decap_8 FILLER_74_735 ();
 sg13g2_decap_8 FILLER_74_742 ();
 sg13g2_decap_8 FILLER_74_749 ();
 sg13g2_decap_8 FILLER_74_756 ();
 sg13g2_decap_8 FILLER_74_763 ();
 sg13g2_decap_8 FILLER_74_770 ();
 sg13g2_decap_8 FILLER_74_777 ();
 sg13g2_decap_8 FILLER_74_784 ();
 sg13g2_decap_8 FILLER_74_791 ();
 sg13g2_decap_8 FILLER_74_798 ();
 sg13g2_decap_8 FILLER_74_805 ();
 sg13g2_decap_8 FILLER_74_812 ();
 sg13g2_decap_8 FILLER_74_819 ();
 sg13g2_decap_8 FILLER_74_826 ();
 sg13g2_decap_8 FILLER_74_833 ();
 sg13g2_decap_8 FILLER_74_840 ();
 sg13g2_decap_8 FILLER_74_847 ();
 sg13g2_decap_8 FILLER_74_854 ();
 sg13g2_decap_8 FILLER_74_861 ();
 sg13g2_decap_8 FILLER_74_868 ();
 sg13g2_decap_8 FILLER_74_875 ();
 sg13g2_decap_8 FILLER_74_882 ();
 sg13g2_decap_8 FILLER_74_889 ();
 sg13g2_decap_8 FILLER_74_896 ();
 sg13g2_decap_8 FILLER_74_903 ();
 sg13g2_decap_8 FILLER_74_910 ();
 sg13g2_decap_8 FILLER_74_917 ();
 sg13g2_decap_8 FILLER_74_924 ();
 sg13g2_decap_8 FILLER_74_931 ();
 sg13g2_decap_8 FILLER_74_938 ();
 sg13g2_decap_8 FILLER_74_945 ();
 sg13g2_decap_8 FILLER_74_952 ();
 sg13g2_decap_8 FILLER_74_959 ();
 sg13g2_decap_8 FILLER_74_966 ();
 sg13g2_decap_8 FILLER_74_973 ();
 sg13g2_decap_8 FILLER_74_980 ();
 sg13g2_decap_8 FILLER_74_987 ();
 sg13g2_decap_8 FILLER_74_994 ();
 sg13g2_decap_8 FILLER_74_1001 ();
 sg13g2_decap_8 FILLER_74_1008 ();
 sg13g2_decap_8 FILLER_74_1015 ();
 sg13g2_decap_8 FILLER_74_1022 ();
 sg13g2_decap_8 FILLER_74_1029 ();
 sg13g2_decap_8 FILLER_74_1036 ();
 sg13g2_decap_8 FILLER_74_1043 ();
 sg13g2_decap_8 FILLER_74_1050 ();
 sg13g2_decap_8 FILLER_74_1057 ();
 sg13g2_decap_8 FILLER_74_1064 ();
 sg13g2_decap_8 FILLER_74_1071 ();
 sg13g2_decap_8 FILLER_74_1078 ();
 sg13g2_decap_8 FILLER_74_1085 ();
 sg13g2_decap_8 FILLER_74_1092 ();
 sg13g2_decap_8 FILLER_74_1099 ();
 sg13g2_decap_8 FILLER_74_1106 ();
 sg13g2_decap_8 FILLER_74_1113 ();
 sg13g2_decap_8 FILLER_74_1120 ();
 sg13g2_decap_8 FILLER_74_1127 ();
 sg13g2_decap_8 FILLER_74_1134 ();
 sg13g2_decap_8 FILLER_74_1141 ();
 sg13g2_decap_8 FILLER_74_1148 ();
 sg13g2_decap_8 FILLER_74_1155 ();
 sg13g2_decap_8 FILLER_74_1162 ();
 sg13g2_decap_8 FILLER_74_1169 ();
 sg13g2_decap_8 FILLER_74_1176 ();
 sg13g2_decap_8 FILLER_74_1183 ();
 sg13g2_decap_8 FILLER_74_1190 ();
 sg13g2_decap_8 FILLER_74_1197 ();
 sg13g2_decap_8 FILLER_74_1204 ();
 sg13g2_decap_8 FILLER_74_1211 ();
 sg13g2_decap_8 FILLER_74_1218 ();
 sg13g2_decap_8 FILLER_74_1225 ();
 sg13g2_decap_8 FILLER_74_1232 ();
 sg13g2_decap_8 FILLER_74_1239 ();
 sg13g2_decap_8 FILLER_74_1246 ();
 sg13g2_decap_8 FILLER_74_1253 ();
 sg13g2_decap_8 FILLER_74_1260 ();
 sg13g2_decap_8 FILLER_74_1267 ();
 sg13g2_decap_8 FILLER_74_1274 ();
 sg13g2_decap_8 FILLER_74_1281 ();
 sg13g2_decap_8 FILLER_74_1288 ();
 sg13g2_decap_8 FILLER_74_1295 ();
 sg13g2_decap_8 FILLER_74_1302 ();
 sg13g2_decap_8 FILLER_74_1309 ();
 sg13g2_decap_8 FILLER_74_1316 ();
 sg13g2_decap_8 FILLER_74_1323 ();
 sg13g2_decap_8 FILLER_74_1330 ();
 sg13g2_decap_8 FILLER_74_1337 ();
 sg13g2_decap_8 FILLER_74_1344 ();
 sg13g2_decap_8 FILLER_74_1351 ();
 sg13g2_decap_8 FILLER_74_1358 ();
 sg13g2_decap_8 FILLER_74_1365 ();
 sg13g2_decap_8 FILLER_74_1372 ();
 sg13g2_decap_8 FILLER_74_1379 ();
 sg13g2_decap_8 FILLER_74_1386 ();
 sg13g2_decap_8 FILLER_74_1393 ();
 sg13g2_decap_8 FILLER_74_1400 ();
 sg13g2_decap_8 FILLER_74_1407 ();
 sg13g2_decap_8 FILLER_74_1414 ();
 sg13g2_decap_8 FILLER_74_1421 ();
 sg13g2_decap_8 FILLER_74_1428 ();
 sg13g2_decap_8 FILLER_74_1435 ();
 sg13g2_decap_8 FILLER_74_1442 ();
 sg13g2_decap_8 FILLER_74_1449 ();
 sg13g2_decap_8 FILLER_74_1456 ();
 sg13g2_decap_8 FILLER_74_1463 ();
 sg13g2_decap_8 FILLER_74_1470 ();
 sg13g2_decap_8 FILLER_74_1477 ();
 sg13g2_decap_8 FILLER_74_1484 ();
 sg13g2_decap_8 FILLER_74_1491 ();
 sg13g2_decap_8 FILLER_74_1498 ();
 sg13g2_decap_8 FILLER_74_1505 ();
 sg13g2_decap_8 FILLER_74_1512 ();
 sg13g2_decap_8 FILLER_74_1519 ();
 sg13g2_decap_8 FILLER_74_1526 ();
 sg13g2_decap_8 FILLER_74_1533 ();
 sg13g2_decap_8 FILLER_74_1540 ();
 sg13g2_decap_8 FILLER_74_1547 ();
 sg13g2_decap_8 FILLER_74_1554 ();
 sg13g2_decap_8 FILLER_74_1561 ();
 sg13g2_decap_8 FILLER_74_1568 ();
 sg13g2_decap_8 FILLER_74_1575 ();
 sg13g2_decap_8 FILLER_74_1582 ();
 sg13g2_decap_8 FILLER_74_1589 ();
 sg13g2_decap_8 FILLER_74_1596 ();
 sg13g2_decap_8 FILLER_74_1603 ();
 sg13g2_decap_8 FILLER_74_1610 ();
 sg13g2_decap_8 FILLER_74_1617 ();
 sg13g2_decap_8 FILLER_74_1624 ();
 sg13g2_decap_8 FILLER_74_1631 ();
 sg13g2_decap_8 FILLER_74_1638 ();
 sg13g2_decap_8 FILLER_74_1645 ();
 sg13g2_decap_8 FILLER_74_1652 ();
 sg13g2_decap_8 FILLER_74_1659 ();
 sg13g2_decap_8 FILLER_74_1666 ();
 sg13g2_decap_8 FILLER_74_1673 ();
 sg13g2_decap_8 FILLER_74_1680 ();
 sg13g2_decap_8 FILLER_74_1687 ();
 sg13g2_decap_8 FILLER_74_1694 ();
 sg13g2_decap_8 FILLER_74_1701 ();
 sg13g2_decap_8 FILLER_74_1708 ();
 sg13g2_decap_8 FILLER_74_1715 ();
 sg13g2_decap_8 FILLER_74_1722 ();
 sg13g2_decap_8 FILLER_74_1729 ();
 sg13g2_decap_8 FILLER_74_1736 ();
 sg13g2_decap_8 FILLER_74_1743 ();
 sg13g2_decap_8 FILLER_74_1750 ();
 sg13g2_decap_8 FILLER_74_1757 ();
 sg13g2_decap_8 FILLER_74_1764 ();
 sg13g2_decap_8 FILLER_74_1771 ();
 sg13g2_decap_8 FILLER_74_1778 ();
 sg13g2_decap_8 FILLER_74_1785 ();
 sg13g2_decap_8 FILLER_74_1792 ();
 sg13g2_decap_8 FILLER_74_1799 ();
 sg13g2_decap_8 FILLER_74_1806 ();
 sg13g2_decap_8 FILLER_74_1813 ();
 sg13g2_decap_8 FILLER_74_1820 ();
 sg13g2_decap_8 FILLER_74_1827 ();
 sg13g2_decap_8 FILLER_74_1834 ();
 sg13g2_decap_8 FILLER_74_1841 ();
 sg13g2_decap_8 FILLER_74_1848 ();
 sg13g2_decap_8 FILLER_74_1855 ();
 sg13g2_decap_8 FILLER_74_1862 ();
 sg13g2_decap_8 FILLER_74_1869 ();
 sg13g2_decap_8 FILLER_74_1876 ();
 sg13g2_decap_8 FILLER_74_1883 ();
 sg13g2_decap_8 FILLER_74_1890 ();
 sg13g2_decap_8 FILLER_74_1897 ();
 sg13g2_decap_8 FILLER_74_1904 ();
 sg13g2_decap_8 FILLER_74_1911 ();
 sg13g2_decap_8 FILLER_74_1918 ();
 sg13g2_decap_8 FILLER_74_1925 ();
 sg13g2_decap_8 FILLER_74_1932 ();
 sg13g2_decap_8 FILLER_74_1939 ();
 sg13g2_decap_8 FILLER_74_1946 ();
 sg13g2_decap_8 FILLER_74_1953 ();
 sg13g2_decap_8 FILLER_74_1960 ();
 sg13g2_decap_8 FILLER_74_1967 ();
 sg13g2_decap_8 FILLER_74_1974 ();
 sg13g2_decap_8 FILLER_74_1981 ();
 sg13g2_decap_8 FILLER_74_1988 ();
 sg13g2_decap_8 FILLER_74_1995 ();
 sg13g2_decap_8 FILLER_74_2002 ();
 sg13g2_decap_8 FILLER_74_2009 ();
 sg13g2_decap_8 FILLER_74_2016 ();
 sg13g2_decap_8 FILLER_74_2023 ();
 sg13g2_decap_8 FILLER_74_2030 ();
 sg13g2_decap_8 FILLER_74_2037 ();
 sg13g2_decap_8 FILLER_74_2044 ();
 sg13g2_decap_8 FILLER_74_2051 ();
 sg13g2_decap_8 FILLER_74_2058 ();
 sg13g2_decap_8 FILLER_74_2065 ();
 sg13g2_decap_8 FILLER_74_2072 ();
 sg13g2_decap_8 FILLER_74_2079 ();
 sg13g2_decap_8 FILLER_74_2086 ();
 sg13g2_decap_8 FILLER_74_2093 ();
 sg13g2_decap_8 FILLER_74_2100 ();
 sg13g2_decap_8 FILLER_74_2107 ();
 sg13g2_decap_8 FILLER_74_2114 ();
 sg13g2_decap_8 FILLER_74_2121 ();
 sg13g2_decap_8 FILLER_74_2128 ();
 sg13g2_decap_8 FILLER_74_2135 ();
 sg13g2_decap_8 FILLER_74_2142 ();
 sg13g2_decap_8 FILLER_74_2149 ();
 sg13g2_decap_8 FILLER_74_2156 ();
 sg13g2_decap_8 FILLER_74_2163 ();
 sg13g2_decap_8 FILLER_74_2170 ();
 sg13g2_decap_8 FILLER_74_2177 ();
 sg13g2_decap_8 FILLER_74_2184 ();
 sg13g2_decap_8 FILLER_74_2191 ();
 sg13g2_decap_8 FILLER_74_2198 ();
 sg13g2_decap_8 FILLER_74_2205 ();
 sg13g2_decap_8 FILLER_74_2212 ();
 sg13g2_decap_8 FILLER_74_2219 ();
 sg13g2_decap_8 FILLER_74_2226 ();
 sg13g2_decap_8 FILLER_74_2233 ();
 sg13g2_decap_8 FILLER_74_2240 ();
 sg13g2_decap_8 FILLER_74_2247 ();
 sg13g2_decap_8 FILLER_74_2254 ();
 sg13g2_decap_8 FILLER_74_2261 ();
 sg13g2_decap_8 FILLER_74_2268 ();
 sg13g2_decap_8 FILLER_74_2275 ();
 sg13g2_decap_8 FILLER_74_2282 ();
 sg13g2_decap_8 FILLER_74_2289 ();
 sg13g2_decap_8 FILLER_74_2296 ();
 sg13g2_decap_8 FILLER_74_2303 ();
 sg13g2_decap_8 FILLER_74_2310 ();
 sg13g2_decap_8 FILLER_74_2317 ();
 sg13g2_decap_8 FILLER_74_2324 ();
 sg13g2_decap_8 FILLER_74_2331 ();
 sg13g2_decap_8 FILLER_74_2338 ();
 sg13g2_decap_8 FILLER_74_2345 ();
 sg13g2_decap_8 FILLER_74_2352 ();
 sg13g2_decap_8 FILLER_74_2359 ();
 sg13g2_decap_8 FILLER_74_2366 ();
 sg13g2_decap_8 FILLER_74_2373 ();
 sg13g2_decap_8 FILLER_74_2380 ();
 sg13g2_decap_8 FILLER_74_2387 ();
 sg13g2_decap_8 FILLER_74_2394 ();
 sg13g2_decap_8 FILLER_74_2401 ();
 sg13g2_decap_8 FILLER_74_2408 ();
 sg13g2_decap_8 FILLER_74_2415 ();
 sg13g2_decap_8 FILLER_74_2422 ();
 sg13g2_decap_8 FILLER_74_2429 ();
 sg13g2_decap_8 FILLER_74_2436 ();
 sg13g2_decap_8 FILLER_74_2443 ();
 sg13g2_decap_8 FILLER_74_2450 ();
 sg13g2_decap_8 FILLER_74_2457 ();
 sg13g2_decap_8 FILLER_74_2464 ();
 sg13g2_decap_8 FILLER_74_2471 ();
 sg13g2_decap_8 FILLER_74_2478 ();
 sg13g2_decap_8 FILLER_74_2485 ();
 sg13g2_decap_8 FILLER_74_2492 ();
 sg13g2_decap_8 FILLER_74_2499 ();
 sg13g2_decap_8 FILLER_74_2506 ();
 sg13g2_decap_8 FILLER_74_2513 ();
 sg13g2_decap_8 FILLER_74_2520 ();
 sg13g2_decap_8 FILLER_74_2527 ();
 sg13g2_decap_8 FILLER_74_2534 ();
 sg13g2_decap_8 FILLER_74_2541 ();
 sg13g2_decap_8 FILLER_74_2548 ();
 sg13g2_decap_8 FILLER_74_2555 ();
 sg13g2_decap_8 FILLER_74_2562 ();
 sg13g2_decap_8 FILLER_74_2569 ();
 sg13g2_decap_8 FILLER_74_2576 ();
 sg13g2_decap_8 FILLER_74_2583 ();
 sg13g2_decap_8 FILLER_74_2590 ();
 sg13g2_decap_8 FILLER_74_2597 ();
 sg13g2_decap_8 FILLER_74_2604 ();
 sg13g2_decap_8 FILLER_74_2611 ();
 sg13g2_decap_8 FILLER_74_2618 ();
 sg13g2_decap_8 FILLER_74_2625 ();
 sg13g2_decap_8 FILLER_74_2632 ();
 sg13g2_decap_8 FILLER_74_2639 ();
 sg13g2_decap_8 FILLER_74_2646 ();
 sg13g2_decap_8 FILLER_74_2653 ();
 sg13g2_decap_8 FILLER_74_2660 ();
 sg13g2_decap_8 FILLER_74_2667 ();
 sg13g2_decap_8 FILLER_74_2674 ();
 sg13g2_decap_8 FILLER_74_2681 ();
 sg13g2_decap_8 FILLER_74_2688 ();
 sg13g2_decap_8 FILLER_74_2695 ();
 sg13g2_decap_8 FILLER_74_2702 ();
 sg13g2_decap_8 FILLER_74_2709 ();
 sg13g2_decap_8 FILLER_74_2716 ();
 sg13g2_decap_8 FILLER_74_2723 ();
 sg13g2_decap_8 FILLER_74_2730 ();
 sg13g2_decap_8 FILLER_74_2737 ();
 sg13g2_decap_8 FILLER_74_2744 ();
 sg13g2_decap_8 FILLER_74_2751 ();
 sg13g2_decap_8 FILLER_74_2758 ();
 sg13g2_decap_8 FILLER_74_2765 ();
 sg13g2_decap_8 FILLER_74_2772 ();
 sg13g2_decap_8 FILLER_74_2779 ();
 sg13g2_decap_8 FILLER_74_2786 ();
 sg13g2_decap_8 FILLER_74_2793 ();
 sg13g2_decap_8 FILLER_74_2800 ();
 sg13g2_decap_8 FILLER_74_2807 ();
 sg13g2_decap_8 FILLER_74_2814 ();
 sg13g2_decap_8 FILLER_74_2821 ();
 sg13g2_decap_8 FILLER_74_2828 ();
 sg13g2_decap_8 FILLER_74_2835 ();
 sg13g2_decap_8 FILLER_74_2842 ();
 sg13g2_decap_8 FILLER_74_2849 ();
 sg13g2_decap_8 FILLER_74_2856 ();
 sg13g2_decap_8 FILLER_74_2863 ();
 sg13g2_decap_8 FILLER_74_2870 ();
 sg13g2_decap_8 FILLER_74_2877 ();
 sg13g2_decap_8 FILLER_74_2884 ();
 sg13g2_decap_8 FILLER_74_2891 ();
 sg13g2_decap_8 FILLER_74_2898 ();
 sg13g2_decap_8 FILLER_74_2905 ();
 sg13g2_decap_8 FILLER_74_2912 ();
 sg13g2_decap_8 FILLER_74_2919 ();
 sg13g2_decap_8 FILLER_74_2926 ();
 sg13g2_decap_8 FILLER_74_2933 ();
 sg13g2_decap_8 FILLER_74_2940 ();
 sg13g2_decap_8 FILLER_74_2947 ();
 sg13g2_decap_8 FILLER_74_2954 ();
 sg13g2_decap_8 FILLER_74_2961 ();
 sg13g2_decap_8 FILLER_74_2968 ();
 sg13g2_decap_8 FILLER_74_2975 ();
 sg13g2_decap_8 FILLER_74_2982 ();
 sg13g2_decap_8 FILLER_74_2989 ();
 sg13g2_decap_8 FILLER_74_2996 ();
 sg13g2_decap_8 FILLER_74_3003 ();
 sg13g2_decap_8 FILLER_74_3010 ();
 sg13g2_decap_8 FILLER_74_3017 ();
 sg13g2_decap_8 FILLER_74_3024 ();
 sg13g2_decap_8 FILLER_74_3031 ();
 sg13g2_decap_8 FILLER_74_3038 ();
 sg13g2_decap_8 FILLER_74_3045 ();
 sg13g2_decap_8 FILLER_74_3052 ();
 sg13g2_decap_8 FILLER_74_3059 ();
 sg13g2_decap_8 FILLER_74_3066 ();
 sg13g2_decap_8 FILLER_74_3073 ();
 sg13g2_decap_8 FILLER_74_3080 ();
 sg13g2_decap_8 FILLER_74_3087 ();
 sg13g2_decap_8 FILLER_74_3094 ();
 sg13g2_decap_8 FILLER_74_3101 ();
 sg13g2_decap_8 FILLER_74_3108 ();
 sg13g2_decap_8 FILLER_74_3115 ();
 sg13g2_decap_8 FILLER_74_3122 ();
 sg13g2_decap_8 FILLER_74_3129 ();
 sg13g2_decap_8 FILLER_74_3136 ();
 sg13g2_decap_8 FILLER_74_3143 ();
 sg13g2_decap_8 FILLER_74_3150 ();
 sg13g2_decap_8 FILLER_74_3157 ();
 sg13g2_decap_8 FILLER_74_3164 ();
 sg13g2_decap_8 FILLER_74_3171 ();
 sg13g2_decap_8 FILLER_74_3178 ();
 sg13g2_decap_8 FILLER_74_3185 ();
 sg13g2_decap_8 FILLER_74_3192 ();
 sg13g2_decap_8 FILLER_74_3199 ();
 sg13g2_decap_8 FILLER_74_3206 ();
 sg13g2_decap_8 FILLER_74_3213 ();
 sg13g2_decap_8 FILLER_74_3220 ();
 sg13g2_decap_8 FILLER_74_3227 ();
 sg13g2_decap_8 FILLER_74_3234 ();
 sg13g2_decap_8 FILLER_74_3241 ();
 sg13g2_decap_8 FILLER_74_3248 ();
 sg13g2_decap_8 FILLER_74_3255 ();
 sg13g2_decap_8 FILLER_74_3262 ();
 sg13g2_decap_8 FILLER_74_3269 ();
 sg13g2_decap_8 FILLER_74_3276 ();
 sg13g2_decap_8 FILLER_74_3283 ();
 sg13g2_decap_8 FILLER_74_3290 ();
 sg13g2_decap_8 FILLER_74_3297 ();
 sg13g2_decap_8 FILLER_74_3304 ();
 sg13g2_decap_8 FILLER_74_3311 ();
 sg13g2_decap_8 FILLER_74_3318 ();
 sg13g2_decap_8 FILLER_74_3325 ();
 sg13g2_decap_8 FILLER_74_3332 ();
 sg13g2_decap_8 FILLER_74_3339 ();
 sg13g2_decap_8 FILLER_74_3346 ();
 sg13g2_decap_8 FILLER_74_3353 ();
 sg13g2_decap_8 FILLER_74_3360 ();
 sg13g2_decap_8 FILLER_74_3367 ();
 sg13g2_decap_8 FILLER_74_3374 ();
 sg13g2_decap_8 FILLER_74_3381 ();
 sg13g2_decap_8 FILLER_74_3388 ();
 sg13g2_decap_8 FILLER_74_3395 ();
 sg13g2_decap_8 FILLER_74_3402 ();
 sg13g2_decap_8 FILLER_74_3409 ();
 sg13g2_decap_8 FILLER_74_3416 ();
 sg13g2_decap_8 FILLER_74_3423 ();
 sg13g2_decap_8 FILLER_74_3430 ();
 sg13g2_decap_8 FILLER_74_3437 ();
 sg13g2_decap_8 FILLER_74_3444 ();
 sg13g2_decap_8 FILLER_74_3451 ();
 sg13g2_decap_8 FILLER_74_3458 ();
 sg13g2_decap_8 FILLER_74_3465 ();
 sg13g2_decap_8 FILLER_74_3472 ();
 sg13g2_decap_8 FILLER_74_3479 ();
 sg13g2_decap_8 FILLER_74_3486 ();
 sg13g2_decap_8 FILLER_74_3493 ();
 sg13g2_decap_8 FILLER_74_3500 ();
 sg13g2_decap_8 FILLER_74_3507 ();
 sg13g2_decap_8 FILLER_74_3514 ();
 sg13g2_decap_8 FILLER_74_3521 ();
 sg13g2_decap_8 FILLER_74_3528 ();
 sg13g2_decap_8 FILLER_74_3535 ();
 sg13g2_decap_8 FILLER_74_3542 ();
 sg13g2_decap_8 FILLER_74_3549 ();
 sg13g2_decap_8 FILLER_74_3556 ();
 sg13g2_decap_8 FILLER_74_3563 ();
 sg13g2_decap_8 FILLER_74_3570 ();
 sg13g2_fill_2 FILLER_74_3577 ();
 sg13g2_fill_1 FILLER_74_3579 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_decap_4 FILLER_75_161 ();
 sg13g2_fill_2 FILLER_75_165 ();
 sg13g2_decap_8 FILLER_75_171 ();
 sg13g2_decap_8 FILLER_75_178 ();
 sg13g2_fill_1 FILLER_75_185 ();
 sg13g2_decap_8 FILLER_75_191 ();
 sg13g2_decap_4 FILLER_75_235 ();
 sg13g2_decap_8 FILLER_75_267 ();
 sg13g2_decap_8 FILLER_75_274 ();
 sg13g2_decap_8 FILLER_75_281 ();
 sg13g2_decap_8 FILLER_75_288 ();
 sg13g2_decap_8 FILLER_75_295 ();
 sg13g2_decap_8 FILLER_75_302 ();
 sg13g2_decap_8 FILLER_75_309 ();
 sg13g2_decap_8 FILLER_75_316 ();
 sg13g2_decap_8 FILLER_75_323 ();
 sg13g2_decap_8 FILLER_75_330 ();
 sg13g2_decap_8 FILLER_75_337 ();
 sg13g2_decap_8 FILLER_75_344 ();
 sg13g2_decap_8 FILLER_75_351 ();
 sg13g2_decap_8 FILLER_75_358 ();
 sg13g2_decap_8 FILLER_75_365 ();
 sg13g2_decap_8 FILLER_75_372 ();
 sg13g2_decap_8 FILLER_75_379 ();
 sg13g2_decap_8 FILLER_75_386 ();
 sg13g2_decap_8 FILLER_75_393 ();
 sg13g2_decap_8 FILLER_75_400 ();
 sg13g2_decap_8 FILLER_75_407 ();
 sg13g2_decap_8 FILLER_75_414 ();
 sg13g2_decap_8 FILLER_75_421 ();
 sg13g2_decap_8 FILLER_75_428 ();
 sg13g2_decap_8 FILLER_75_435 ();
 sg13g2_decap_8 FILLER_75_442 ();
 sg13g2_decap_8 FILLER_75_449 ();
 sg13g2_decap_8 FILLER_75_456 ();
 sg13g2_decap_8 FILLER_75_463 ();
 sg13g2_decap_8 FILLER_75_470 ();
 sg13g2_decap_8 FILLER_75_477 ();
 sg13g2_decap_8 FILLER_75_484 ();
 sg13g2_decap_8 FILLER_75_491 ();
 sg13g2_decap_8 FILLER_75_498 ();
 sg13g2_decap_8 FILLER_75_505 ();
 sg13g2_decap_8 FILLER_75_512 ();
 sg13g2_decap_8 FILLER_75_519 ();
 sg13g2_decap_8 FILLER_75_526 ();
 sg13g2_decap_8 FILLER_75_533 ();
 sg13g2_decap_8 FILLER_75_540 ();
 sg13g2_decap_8 FILLER_75_547 ();
 sg13g2_decap_8 FILLER_75_554 ();
 sg13g2_decap_8 FILLER_75_561 ();
 sg13g2_decap_8 FILLER_75_568 ();
 sg13g2_decap_8 FILLER_75_575 ();
 sg13g2_decap_8 FILLER_75_582 ();
 sg13g2_decap_8 FILLER_75_589 ();
 sg13g2_decap_8 FILLER_75_596 ();
 sg13g2_decap_8 FILLER_75_603 ();
 sg13g2_decap_8 FILLER_75_610 ();
 sg13g2_decap_8 FILLER_75_617 ();
 sg13g2_decap_8 FILLER_75_624 ();
 sg13g2_decap_8 FILLER_75_631 ();
 sg13g2_decap_8 FILLER_75_638 ();
 sg13g2_decap_8 FILLER_75_645 ();
 sg13g2_decap_8 FILLER_75_652 ();
 sg13g2_decap_8 FILLER_75_659 ();
 sg13g2_decap_8 FILLER_75_666 ();
 sg13g2_decap_8 FILLER_75_673 ();
 sg13g2_decap_8 FILLER_75_680 ();
 sg13g2_decap_8 FILLER_75_687 ();
 sg13g2_decap_8 FILLER_75_694 ();
 sg13g2_decap_8 FILLER_75_701 ();
 sg13g2_decap_8 FILLER_75_708 ();
 sg13g2_decap_8 FILLER_75_715 ();
 sg13g2_decap_8 FILLER_75_722 ();
 sg13g2_decap_8 FILLER_75_729 ();
 sg13g2_decap_8 FILLER_75_736 ();
 sg13g2_decap_8 FILLER_75_743 ();
 sg13g2_decap_8 FILLER_75_750 ();
 sg13g2_decap_8 FILLER_75_757 ();
 sg13g2_decap_8 FILLER_75_764 ();
 sg13g2_decap_8 FILLER_75_771 ();
 sg13g2_decap_8 FILLER_75_778 ();
 sg13g2_decap_8 FILLER_75_785 ();
 sg13g2_decap_8 FILLER_75_792 ();
 sg13g2_decap_8 FILLER_75_799 ();
 sg13g2_decap_8 FILLER_75_806 ();
 sg13g2_decap_8 FILLER_75_813 ();
 sg13g2_decap_8 FILLER_75_820 ();
 sg13g2_decap_8 FILLER_75_827 ();
 sg13g2_decap_8 FILLER_75_834 ();
 sg13g2_decap_8 FILLER_75_841 ();
 sg13g2_decap_8 FILLER_75_848 ();
 sg13g2_decap_8 FILLER_75_855 ();
 sg13g2_decap_8 FILLER_75_862 ();
 sg13g2_decap_8 FILLER_75_869 ();
 sg13g2_decap_8 FILLER_75_876 ();
 sg13g2_decap_8 FILLER_75_883 ();
 sg13g2_decap_8 FILLER_75_890 ();
 sg13g2_decap_8 FILLER_75_897 ();
 sg13g2_decap_8 FILLER_75_904 ();
 sg13g2_decap_8 FILLER_75_911 ();
 sg13g2_decap_8 FILLER_75_918 ();
 sg13g2_decap_8 FILLER_75_925 ();
 sg13g2_decap_8 FILLER_75_932 ();
 sg13g2_decap_8 FILLER_75_939 ();
 sg13g2_decap_8 FILLER_75_946 ();
 sg13g2_decap_8 FILLER_75_953 ();
 sg13g2_decap_8 FILLER_75_960 ();
 sg13g2_decap_8 FILLER_75_967 ();
 sg13g2_decap_8 FILLER_75_974 ();
 sg13g2_decap_8 FILLER_75_981 ();
 sg13g2_decap_8 FILLER_75_988 ();
 sg13g2_decap_8 FILLER_75_995 ();
 sg13g2_decap_8 FILLER_75_1002 ();
 sg13g2_decap_8 FILLER_75_1009 ();
 sg13g2_decap_8 FILLER_75_1016 ();
 sg13g2_decap_8 FILLER_75_1023 ();
 sg13g2_decap_8 FILLER_75_1030 ();
 sg13g2_decap_8 FILLER_75_1037 ();
 sg13g2_decap_8 FILLER_75_1044 ();
 sg13g2_decap_8 FILLER_75_1051 ();
 sg13g2_decap_8 FILLER_75_1058 ();
 sg13g2_decap_8 FILLER_75_1065 ();
 sg13g2_decap_8 FILLER_75_1072 ();
 sg13g2_decap_8 FILLER_75_1079 ();
 sg13g2_decap_8 FILLER_75_1086 ();
 sg13g2_decap_8 FILLER_75_1093 ();
 sg13g2_decap_8 FILLER_75_1100 ();
 sg13g2_decap_8 FILLER_75_1107 ();
 sg13g2_decap_8 FILLER_75_1114 ();
 sg13g2_decap_8 FILLER_75_1121 ();
 sg13g2_decap_8 FILLER_75_1128 ();
 sg13g2_decap_8 FILLER_75_1135 ();
 sg13g2_decap_8 FILLER_75_1142 ();
 sg13g2_decap_8 FILLER_75_1149 ();
 sg13g2_decap_8 FILLER_75_1156 ();
 sg13g2_decap_8 FILLER_75_1163 ();
 sg13g2_decap_8 FILLER_75_1170 ();
 sg13g2_decap_8 FILLER_75_1177 ();
 sg13g2_decap_8 FILLER_75_1184 ();
 sg13g2_decap_8 FILLER_75_1191 ();
 sg13g2_decap_8 FILLER_75_1198 ();
 sg13g2_decap_8 FILLER_75_1205 ();
 sg13g2_decap_8 FILLER_75_1212 ();
 sg13g2_decap_8 FILLER_75_1219 ();
 sg13g2_decap_8 FILLER_75_1226 ();
 sg13g2_decap_8 FILLER_75_1233 ();
 sg13g2_decap_8 FILLER_75_1240 ();
 sg13g2_decap_8 FILLER_75_1247 ();
 sg13g2_decap_8 FILLER_75_1254 ();
 sg13g2_decap_8 FILLER_75_1261 ();
 sg13g2_decap_8 FILLER_75_1268 ();
 sg13g2_decap_8 FILLER_75_1275 ();
 sg13g2_decap_8 FILLER_75_1282 ();
 sg13g2_decap_8 FILLER_75_1289 ();
 sg13g2_decap_8 FILLER_75_1296 ();
 sg13g2_decap_8 FILLER_75_1303 ();
 sg13g2_decap_8 FILLER_75_1310 ();
 sg13g2_decap_8 FILLER_75_1317 ();
 sg13g2_decap_8 FILLER_75_1324 ();
 sg13g2_decap_8 FILLER_75_1331 ();
 sg13g2_decap_8 FILLER_75_1338 ();
 sg13g2_decap_8 FILLER_75_1345 ();
 sg13g2_decap_8 FILLER_75_1352 ();
 sg13g2_decap_8 FILLER_75_1359 ();
 sg13g2_decap_8 FILLER_75_1366 ();
 sg13g2_decap_8 FILLER_75_1373 ();
 sg13g2_decap_8 FILLER_75_1380 ();
 sg13g2_decap_8 FILLER_75_1387 ();
 sg13g2_decap_8 FILLER_75_1394 ();
 sg13g2_decap_8 FILLER_75_1401 ();
 sg13g2_decap_8 FILLER_75_1408 ();
 sg13g2_decap_8 FILLER_75_1415 ();
 sg13g2_decap_8 FILLER_75_1422 ();
 sg13g2_decap_8 FILLER_75_1429 ();
 sg13g2_decap_8 FILLER_75_1436 ();
 sg13g2_decap_8 FILLER_75_1443 ();
 sg13g2_decap_8 FILLER_75_1450 ();
 sg13g2_decap_8 FILLER_75_1457 ();
 sg13g2_decap_8 FILLER_75_1464 ();
 sg13g2_decap_8 FILLER_75_1471 ();
 sg13g2_decap_8 FILLER_75_1478 ();
 sg13g2_decap_8 FILLER_75_1485 ();
 sg13g2_decap_8 FILLER_75_1492 ();
 sg13g2_decap_8 FILLER_75_1499 ();
 sg13g2_decap_8 FILLER_75_1506 ();
 sg13g2_decap_8 FILLER_75_1513 ();
 sg13g2_decap_8 FILLER_75_1520 ();
 sg13g2_decap_8 FILLER_75_1527 ();
 sg13g2_decap_8 FILLER_75_1534 ();
 sg13g2_decap_8 FILLER_75_1541 ();
 sg13g2_decap_8 FILLER_75_1548 ();
 sg13g2_decap_8 FILLER_75_1555 ();
 sg13g2_decap_8 FILLER_75_1562 ();
 sg13g2_decap_8 FILLER_75_1569 ();
 sg13g2_decap_8 FILLER_75_1576 ();
 sg13g2_decap_8 FILLER_75_1583 ();
 sg13g2_decap_8 FILLER_75_1590 ();
 sg13g2_decap_8 FILLER_75_1597 ();
 sg13g2_decap_8 FILLER_75_1604 ();
 sg13g2_decap_8 FILLER_75_1611 ();
 sg13g2_decap_8 FILLER_75_1618 ();
 sg13g2_decap_8 FILLER_75_1625 ();
 sg13g2_decap_8 FILLER_75_1632 ();
 sg13g2_decap_8 FILLER_75_1639 ();
 sg13g2_decap_8 FILLER_75_1646 ();
 sg13g2_decap_8 FILLER_75_1653 ();
 sg13g2_decap_8 FILLER_75_1660 ();
 sg13g2_decap_8 FILLER_75_1667 ();
 sg13g2_decap_8 FILLER_75_1674 ();
 sg13g2_decap_8 FILLER_75_1681 ();
 sg13g2_decap_8 FILLER_75_1688 ();
 sg13g2_decap_8 FILLER_75_1695 ();
 sg13g2_decap_8 FILLER_75_1702 ();
 sg13g2_decap_8 FILLER_75_1709 ();
 sg13g2_decap_8 FILLER_75_1716 ();
 sg13g2_decap_8 FILLER_75_1723 ();
 sg13g2_decap_8 FILLER_75_1730 ();
 sg13g2_decap_8 FILLER_75_1737 ();
 sg13g2_decap_8 FILLER_75_1744 ();
 sg13g2_decap_8 FILLER_75_1751 ();
 sg13g2_decap_8 FILLER_75_1758 ();
 sg13g2_decap_8 FILLER_75_1765 ();
 sg13g2_decap_8 FILLER_75_1772 ();
 sg13g2_decap_8 FILLER_75_1779 ();
 sg13g2_decap_8 FILLER_75_1786 ();
 sg13g2_decap_8 FILLER_75_1793 ();
 sg13g2_decap_8 FILLER_75_1800 ();
 sg13g2_decap_8 FILLER_75_1807 ();
 sg13g2_decap_8 FILLER_75_1814 ();
 sg13g2_decap_8 FILLER_75_1821 ();
 sg13g2_decap_8 FILLER_75_1828 ();
 sg13g2_decap_8 FILLER_75_1835 ();
 sg13g2_decap_8 FILLER_75_1842 ();
 sg13g2_decap_8 FILLER_75_1849 ();
 sg13g2_decap_8 FILLER_75_1856 ();
 sg13g2_decap_8 FILLER_75_1863 ();
 sg13g2_decap_8 FILLER_75_1870 ();
 sg13g2_decap_8 FILLER_75_1877 ();
 sg13g2_decap_8 FILLER_75_1884 ();
 sg13g2_decap_8 FILLER_75_1891 ();
 sg13g2_decap_8 FILLER_75_1898 ();
 sg13g2_decap_8 FILLER_75_1905 ();
 sg13g2_decap_8 FILLER_75_1912 ();
 sg13g2_decap_8 FILLER_75_1919 ();
 sg13g2_decap_8 FILLER_75_1926 ();
 sg13g2_decap_8 FILLER_75_1933 ();
 sg13g2_decap_8 FILLER_75_1940 ();
 sg13g2_decap_8 FILLER_75_1947 ();
 sg13g2_decap_8 FILLER_75_1954 ();
 sg13g2_decap_8 FILLER_75_1961 ();
 sg13g2_decap_8 FILLER_75_1968 ();
 sg13g2_decap_8 FILLER_75_1975 ();
 sg13g2_decap_8 FILLER_75_1982 ();
 sg13g2_decap_8 FILLER_75_1989 ();
 sg13g2_decap_8 FILLER_75_1996 ();
 sg13g2_decap_8 FILLER_75_2003 ();
 sg13g2_decap_8 FILLER_75_2010 ();
 sg13g2_decap_8 FILLER_75_2017 ();
 sg13g2_decap_8 FILLER_75_2024 ();
 sg13g2_decap_8 FILLER_75_2031 ();
 sg13g2_decap_8 FILLER_75_2038 ();
 sg13g2_decap_8 FILLER_75_2045 ();
 sg13g2_decap_8 FILLER_75_2052 ();
 sg13g2_decap_8 FILLER_75_2059 ();
 sg13g2_decap_8 FILLER_75_2066 ();
 sg13g2_decap_8 FILLER_75_2073 ();
 sg13g2_decap_8 FILLER_75_2080 ();
 sg13g2_decap_8 FILLER_75_2087 ();
 sg13g2_decap_8 FILLER_75_2094 ();
 sg13g2_decap_8 FILLER_75_2101 ();
 sg13g2_decap_8 FILLER_75_2108 ();
 sg13g2_decap_8 FILLER_75_2115 ();
 sg13g2_decap_8 FILLER_75_2122 ();
 sg13g2_decap_8 FILLER_75_2129 ();
 sg13g2_decap_8 FILLER_75_2136 ();
 sg13g2_decap_8 FILLER_75_2143 ();
 sg13g2_decap_8 FILLER_75_2150 ();
 sg13g2_decap_8 FILLER_75_2157 ();
 sg13g2_decap_8 FILLER_75_2164 ();
 sg13g2_decap_8 FILLER_75_2171 ();
 sg13g2_decap_8 FILLER_75_2178 ();
 sg13g2_decap_8 FILLER_75_2185 ();
 sg13g2_decap_8 FILLER_75_2192 ();
 sg13g2_decap_8 FILLER_75_2199 ();
 sg13g2_decap_8 FILLER_75_2206 ();
 sg13g2_decap_8 FILLER_75_2213 ();
 sg13g2_decap_8 FILLER_75_2220 ();
 sg13g2_decap_8 FILLER_75_2227 ();
 sg13g2_decap_8 FILLER_75_2234 ();
 sg13g2_decap_8 FILLER_75_2241 ();
 sg13g2_decap_8 FILLER_75_2248 ();
 sg13g2_decap_8 FILLER_75_2255 ();
 sg13g2_decap_8 FILLER_75_2262 ();
 sg13g2_decap_8 FILLER_75_2269 ();
 sg13g2_decap_8 FILLER_75_2276 ();
 sg13g2_decap_8 FILLER_75_2283 ();
 sg13g2_decap_8 FILLER_75_2290 ();
 sg13g2_decap_8 FILLER_75_2297 ();
 sg13g2_decap_8 FILLER_75_2304 ();
 sg13g2_decap_8 FILLER_75_2311 ();
 sg13g2_decap_8 FILLER_75_2318 ();
 sg13g2_decap_8 FILLER_75_2325 ();
 sg13g2_decap_8 FILLER_75_2332 ();
 sg13g2_decap_8 FILLER_75_2339 ();
 sg13g2_decap_8 FILLER_75_2346 ();
 sg13g2_decap_8 FILLER_75_2353 ();
 sg13g2_decap_8 FILLER_75_2360 ();
 sg13g2_decap_8 FILLER_75_2367 ();
 sg13g2_decap_8 FILLER_75_2374 ();
 sg13g2_decap_8 FILLER_75_2381 ();
 sg13g2_decap_8 FILLER_75_2388 ();
 sg13g2_decap_8 FILLER_75_2395 ();
 sg13g2_decap_8 FILLER_75_2402 ();
 sg13g2_decap_8 FILLER_75_2409 ();
 sg13g2_decap_8 FILLER_75_2416 ();
 sg13g2_decap_8 FILLER_75_2423 ();
 sg13g2_decap_8 FILLER_75_2430 ();
 sg13g2_decap_8 FILLER_75_2437 ();
 sg13g2_decap_8 FILLER_75_2444 ();
 sg13g2_decap_8 FILLER_75_2451 ();
 sg13g2_decap_8 FILLER_75_2458 ();
 sg13g2_decap_8 FILLER_75_2465 ();
 sg13g2_decap_8 FILLER_75_2472 ();
 sg13g2_decap_8 FILLER_75_2479 ();
 sg13g2_decap_8 FILLER_75_2486 ();
 sg13g2_decap_8 FILLER_75_2493 ();
 sg13g2_decap_8 FILLER_75_2500 ();
 sg13g2_decap_8 FILLER_75_2507 ();
 sg13g2_decap_8 FILLER_75_2514 ();
 sg13g2_decap_8 FILLER_75_2521 ();
 sg13g2_decap_8 FILLER_75_2528 ();
 sg13g2_decap_8 FILLER_75_2535 ();
 sg13g2_decap_8 FILLER_75_2542 ();
 sg13g2_decap_8 FILLER_75_2549 ();
 sg13g2_decap_8 FILLER_75_2556 ();
 sg13g2_decap_8 FILLER_75_2563 ();
 sg13g2_decap_8 FILLER_75_2570 ();
 sg13g2_decap_8 FILLER_75_2577 ();
 sg13g2_decap_8 FILLER_75_2584 ();
 sg13g2_decap_8 FILLER_75_2591 ();
 sg13g2_decap_8 FILLER_75_2598 ();
 sg13g2_decap_8 FILLER_75_2605 ();
 sg13g2_decap_8 FILLER_75_2612 ();
 sg13g2_decap_8 FILLER_75_2619 ();
 sg13g2_decap_8 FILLER_75_2626 ();
 sg13g2_decap_8 FILLER_75_2633 ();
 sg13g2_decap_8 FILLER_75_2640 ();
 sg13g2_decap_8 FILLER_75_2647 ();
 sg13g2_decap_8 FILLER_75_2654 ();
 sg13g2_decap_8 FILLER_75_2661 ();
 sg13g2_decap_8 FILLER_75_2668 ();
 sg13g2_decap_8 FILLER_75_2675 ();
 sg13g2_decap_8 FILLER_75_2682 ();
 sg13g2_decap_8 FILLER_75_2689 ();
 sg13g2_decap_8 FILLER_75_2696 ();
 sg13g2_decap_8 FILLER_75_2703 ();
 sg13g2_decap_8 FILLER_75_2710 ();
 sg13g2_decap_8 FILLER_75_2717 ();
 sg13g2_decap_8 FILLER_75_2724 ();
 sg13g2_decap_8 FILLER_75_2731 ();
 sg13g2_decap_8 FILLER_75_2738 ();
 sg13g2_decap_8 FILLER_75_2745 ();
 sg13g2_decap_8 FILLER_75_2752 ();
 sg13g2_decap_8 FILLER_75_2759 ();
 sg13g2_decap_8 FILLER_75_2766 ();
 sg13g2_decap_8 FILLER_75_2773 ();
 sg13g2_decap_8 FILLER_75_2780 ();
 sg13g2_decap_8 FILLER_75_2787 ();
 sg13g2_decap_8 FILLER_75_2794 ();
 sg13g2_decap_8 FILLER_75_2801 ();
 sg13g2_decap_8 FILLER_75_2808 ();
 sg13g2_decap_8 FILLER_75_2815 ();
 sg13g2_decap_8 FILLER_75_2822 ();
 sg13g2_decap_8 FILLER_75_2829 ();
 sg13g2_decap_8 FILLER_75_2836 ();
 sg13g2_decap_8 FILLER_75_2843 ();
 sg13g2_decap_8 FILLER_75_2850 ();
 sg13g2_decap_8 FILLER_75_2857 ();
 sg13g2_decap_8 FILLER_75_2864 ();
 sg13g2_decap_8 FILLER_75_2871 ();
 sg13g2_decap_8 FILLER_75_2878 ();
 sg13g2_decap_8 FILLER_75_2885 ();
 sg13g2_decap_8 FILLER_75_2892 ();
 sg13g2_decap_8 FILLER_75_2899 ();
 sg13g2_decap_8 FILLER_75_2906 ();
 sg13g2_decap_8 FILLER_75_2913 ();
 sg13g2_decap_8 FILLER_75_2920 ();
 sg13g2_decap_8 FILLER_75_2927 ();
 sg13g2_decap_8 FILLER_75_2934 ();
 sg13g2_decap_8 FILLER_75_2941 ();
 sg13g2_decap_8 FILLER_75_2948 ();
 sg13g2_decap_8 FILLER_75_2955 ();
 sg13g2_decap_8 FILLER_75_2962 ();
 sg13g2_decap_8 FILLER_75_2969 ();
 sg13g2_decap_8 FILLER_75_2976 ();
 sg13g2_decap_8 FILLER_75_2983 ();
 sg13g2_decap_8 FILLER_75_2990 ();
 sg13g2_decap_8 FILLER_75_2997 ();
 sg13g2_decap_8 FILLER_75_3004 ();
 sg13g2_decap_8 FILLER_75_3011 ();
 sg13g2_decap_8 FILLER_75_3018 ();
 sg13g2_decap_8 FILLER_75_3025 ();
 sg13g2_decap_8 FILLER_75_3032 ();
 sg13g2_decap_8 FILLER_75_3039 ();
 sg13g2_decap_8 FILLER_75_3046 ();
 sg13g2_decap_8 FILLER_75_3053 ();
 sg13g2_decap_8 FILLER_75_3060 ();
 sg13g2_decap_8 FILLER_75_3067 ();
 sg13g2_decap_8 FILLER_75_3074 ();
 sg13g2_decap_8 FILLER_75_3081 ();
 sg13g2_decap_8 FILLER_75_3088 ();
 sg13g2_decap_8 FILLER_75_3095 ();
 sg13g2_decap_8 FILLER_75_3102 ();
 sg13g2_decap_8 FILLER_75_3109 ();
 sg13g2_decap_8 FILLER_75_3116 ();
 sg13g2_decap_8 FILLER_75_3123 ();
 sg13g2_decap_8 FILLER_75_3130 ();
 sg13g2_decap_8 FILLER_75_3137 ();
 sg13g2_decap_8 FILLER_75_3144 ();
 sg13g2_decap_8 FILLER_75_3151 ();
 sg13g2_decap_8 FILLER_75_3158 ();
 sg13g2_decap_8 FILLER_75_3165 ();
 sg13g2_decap_8 FILLER_75_3172 ();
 sg13g2_decap_8 FILLER_75_3179 ();
 sg13g2_decap_8 FILLER_75_3186 ();
 sg13g2_decap_8 FILLER_75_3193 ();
 sg13g2_decap_8 FILLER_75_3200 ();
 sg13g2_decap_8 FILLER_75_3207 ();
 sg13g2_decap_8 FILLER_75_3214 ();
 sg13g2_decap_8 FILLER_75_3221 ();
 sg13g2_decap_8 FILLER_75_3228 ();
 sg13g2_decap_8 FILLER_75_3235 ();
 sg13g2_decap_8 FILLER_75_3242 ();
 sg13g2_decap_8 FILLER_75_3249 ();
 sg13g2_decap_8 FILLER_75_3256 ();
 sg13g2_decap_8 FILLER_75_3263 ();
 sg13g2_decap_8 FILLER_75_3270 ();
 sg13g2_decap_8 FILLER_75_3277 ();
 sg13g2_decap_8 FILLER_75_3284 ();
 sg13g2_decap_8 FILLER_75_3291 ();
 sg13g2_decap_8 FILLER_75_3298 ();
 sg13g2_decap_8 FILLER_75_3305 ();
 sg13g2_decap_8 FILLER_75_3312 ();
 sg13g2_decap_8 FILLER_75_3319 ();
 sg13g2_decap_8 FILLER_75_3326 ();
 sg13g2_decap_8 FILLER_75_3333 ();
 sg13g2_decap_8 FILLER_75_3340 ();
 sg13g2_decap_8 FILLER_75_3347 ();
 sg13g2_decap_8 FILLER_75_3354 ();
 sg13g2_decap_8 FILLER_75_3361 ();
 sg13g2_decap_8 FILLER_75_3368 ();
 sg13g2_decap_8 FILLER_75_3375 ();
 sg13g2_decap_8 FILLER_75_3382 ();
 sg13g2_decap_8 FILLER_75_3389 ();
 sg13g2_decap_8 FILLER_75_3396 ();
 sg13g2_decap_8 FILLER_75_3403 ();
 sg13g2_decap_8 FILLER_75_3410 ();
 sg13g2_decap_8 FILLER_75_3417 ();
 sg13g2_decap_8 FILLER_75_3424 ();
 sg13g2_decap_8 FILLER_75_3431 ();
 sg13g2_decap_8 FILLER_75_3438 ();
 sg13g2_decap_8 FILLER_75_3445 ();
 sg13g2_decap_8 FILLER_75_3452 ();
 sg13g2_decap_8 FILLER_75_3459 ();
 sg13g2_decap_8 FILLER_75_3466 ();
 sg13g2_decap_8 FILLER_75_3473 ();
 sg13g2_decap_8 FILLER_75_3480 ();
 sg13g2_decap_8 FILLER_75_3487 ();
 sg13g2_decap_8 FILLER_75_3494 ();
 sg13g2_decap_8 FILLER_75_3501 ();
 sg13g2_decap_8 FILLER_75_3508 ();
 sg13g2_decap_8 FILLER_75_3515 ();
 sg13g2_decap_8 FILLER_75_3522 ();
 sg13g2_decap_8 FILLER_75_3529 ();
 sg13g2_decap_8 FILLER_75_3536 ();
 sg13g2_decap_8 FILLER_75_3543 ();
 sg13g2_decap_8 FILLER_75_3550 ();
 sg13g2_decap_8 FILLER_75_3557 ();
 sg13g2_decap_8 FILLER_75_3564 ();
 sg13g2_decap_8 FILLER_75_3571 ();
 sg13g2_fill_2 FILLER_75_3578 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_decap_8 FILLER_76_168 ();
 sg13g2_decap_8 FILLER_76_175 ();
 sg13g2_decap_8 FILLER_76_182 ();
 sg13g2_decap_8 FILLER_76_189 ();
 sg13g2_decap_8 FILLER_76_196 ();
 sg13g2_decap_8 FILLER_76_207 ();
 sg13g2_decap_8 FILLER_76_214 ();
 sg13g2_decap_8 FILLER_76_221 ();
 sg13g2_decap_8 FILLER_76_228 ();
 sg13g2_decap_8 FILLER_76_235 ();
 sg13g2_fill_2 FILLER_76_242 ();
 sg13g2_fill_1 FILLER_76_244 ();
 sg13g2_decap_8 FILLER_76_249 ();
 sg13g2_decap_8 FILLER_76_256 ();
 sg13g2_decap_8 FILLER_76_263 ();
 sg13g2_decap_8 FILLER_76_270 ();
 sg13g2_decap_8 FILLER_76_277 ();
 sg13g2_decap_8 FILLER_76_284 ();
 sg13g2_decap_8 FILLER_76_291 ();
 sg13g2_decap_8 FILLER_76_298 ();
 sg13g2_decap_8 FILLER_76_305 ();
 sg13g2_decap_8 FILLER_76_312 ();
 sg13g2_decap_8 FILLER_76_319 ();
 sg13g2_decap_8 FILLER_76_326 ();
 sg13g2_decap_8 FILLER_76_333 ();
 sg13g2_decap_8 FILLER_76_340 ();
 sg13g2_decap_8 FILLER_76_347 ();
 sg13g2_decap_8 FILLER_76_354 ();
 sg13g2_decap_8 FILLER_76_361 ();
 sg13g2_decap_8 FILLER_76_368 ();
 sg13g2_decap_8 FILLER_76_375 ();
 sg13g2_decap_8 FILLER_76_382 ();
 sg13g2_decap_8 FILLER_76_389 ();
 sg13g2_decap_8 FILLER_76_396 ();
 sg13g2_decap_8 FILLER_76_403 ();
 sg13g2_decap_8 FILLER_76_410 ();
 sg13g2_decap_8 FILLER_76_417 ();
 sg13g2_decap_8 FILLER_76_424 ();
 sg13g2_decap_8 FILLER_76_431 ();
 sg13g2_decap_8 FILLER_76_438 ();
 sg13g2_decap_8 FILLER_76_445 ();
 sg13g2_decap_8 FILLER_76_452 ();
 sg13g2_decap_8 FILLER_76_459 ();
 sg13g2_decap_8 FILLER_76_466 ();
 sg13g2_decap_8 FILLER_76_473 ();
 sg13g2_decap_8 FILLER_76_480 ();
 sg13g2_decap_8 FILLER_76_487 ();
 sg13g2_decap_8 FILLER_76_494 ();
 sg13g2_decap_8 FILLER_76_501 ();
 sg13g2_decap_8 FILLER_76_508 ();
 sg13g2_decap_8 FILLER_76_515 ();
 sg13g2_decap_8 FILLER_76_522 ();
 sg13g2_decap_8 FILLER_76_529 ();
 sg13g2_decap_8 FILLER_76_536 ();
 sg13g2_decap_8 FILLER_76_543 ();
 sg13g2_decap_8 FILLER_76_550 ();
 sg13g2_decap_8 FILLER_76_557 ();
 sg13g2_decap_8 FILLER_76_564 ();
 sg13g2_decap_8 FILLER_76_571 ();
 sg13g2_decap_8 FILLER_76_578 ();
 sg13g2_decap_8 FILLER_76_585 ();
 sg13g2_decap_8 FILLER_76_592 ();
 sg13g2_decap_8 FILLER_76_599 ();
 sg13g2_decap_8 FILLER_76_606 ();
 sg13g2_decap_8 FILLER_76_613 ();
 sg13g2_decap_8 FILLER_76_620 ();
 sg13g2_decap_8 FILLER_76_627 ();
 sg13g2_decap_8 FILLER_76_634 ();
 sg13g2_decap_8 FILLER_76_641 ();
 sg13g2_decap_8 FILLER_76_648 ();
 sg13g2_decap_8 FILLER_76_655 ();
 sg13g2_decap_8 FILLER_76_662 ();
 sg13g2_decap_8 FILLER_76_669 ();
 sg13g2_decap_8 FILLER_76_676 ();
 sg13g2_decap_8 FILLER_76_683 ();
 sg13g2_decap_8 FILLER_76_690 ();
 sg13g2_decap_8 FILLER_76_697 ();
 sg13g2_decap_8 FILLER_76_704 ();
 sg13g2_decap_8 FILLER_76_711 ();
 sg13g2_decap_8 FILLER_76_718 ();
 sg13g2_decap_8 FILLER_76_725 ();
 sg13g2_decap_8 FILLER_76_732 ();
 sg13g2_decap_8 FILLER_76_739 ();
 sg13g2_decap_8 FILLER_76_746 ();
 sg13g2_decap_8 FILLER_76_753 ();
 sg13g2_decap_8 FILLER_76_760 ();
 sg13g2_decap_8 FILLER_76_767 ();
 sg13g2_decap_8 FILLER_76_774 ();
 sg13g2_decap_8 FILLER_76_781 ();
 sg13g2_decap_8 FILLER_76_788 ();
 sg13g2_decap_8 FILLER_76_795 ();
 sg13g2_decap_8 FILLER_76_802 ();
 sg13g2_decap_8 FILLER_76_809 ();
 sg13g2_decap_8 FILLER_76_816 ();
 sg13g2_decap_8 FILLER_76_823 ();
 sg13g2_decap_8 FILLER_76_830 ();
 sg13g2_decap_8 FILLER_76_837 ();
 sg13g2_decap_8 FILLER_76_844 ();
 sg13g2_decap_8 FILLER_76_851 ();
 sg13g2_decap_8 FILLER_76_858 ();
 sg13g2_decap_8 FILLER_76_865 ();
 sg13g2_decap_8 FILLER_76_872 ();
 sg13g2_decap_8 FILLER_76_879 ();
 sg13g2_decap_8 FILLER_76_886 ();
 sg13g2_decap_8 FILLER_76_893 ();
 sg13g2_decap_8 FILLER_76_900 ();
 sg13g2_decap_8 FILLER_76_907 ();
 sg13g2_decap_8 FILLER_76_914 ();
 sg13g2_decap_8 FILLER_76_921 ();
 sg13g2_decap_8 FILLER_76_928 ();
 sg13g2_decap_8 FILLER_76_935 ();
 sg13g2_decap_8 FILLER_76_942 ();
 sg13g2_decap_8 FILLER_76_949 ();
 sg13g2_decap_8 FILLER_76_956 ();
 sg13g2_decap_8 FILLER_76_963 ();
 sg13g2_decap_8 FILLER_76_970 ();
 sg13g2_decap_8 FILLER_76_977 ();
 sg13g2_decap_8 FILLER_76_984 ();
 sg13g2_decap_8 FILLER_76_991 ();
 sg13g2_decap_8 FILLER_76_998 ();
 sg13g2_decap_8 FILLER_76_1005 ();
 sg13g2_decap_8 FILLER_76_1012 ();
 sg13g2_decap_8 FILLER_76_1019 ();
 sg13g2_decap_8 FILLER_76_1026 ();
 sg13g2_decap_8 FILLER_76_1033 ();
 sg13g2_decap_8 FILLER_76_1040 ();
 sg13g2_decap_8 FILLER_76_1047 ();
 sg13g2_decap_8 FILLER_76_1054 ();
 sg13g2_decap_8 FILLER_76_1061 ();
 sg13g2_decap_8 FILLER_76_1068 ();
 sg13g2_decap_8 FILLER_76_1075 ();
 sg13g2_decap_8 FILLER_76_1082 ();
 sg13g2_decap_8 FILLER_76_1089 ();
 sg13g2_decap_8 FILLER_76_1096 ();
 sg13g2_decap_8 FILLER_76_1103 ();
 sg13g2_decap_8 FILLER_76_1110 ();
 sg13g2_decap_8 FILLER_76_1117 ();
 sg13g2_decap_8 FILLER_76_1124 ();
 sg13g2_decap_8 FILLER_76_1131 ();
 sg13g2_decap_8 FILLER_76_1138 ();
 sg13g2_decap_8 FILLER_76_1145 ();
 sg13g2_decap_8 FILLER_76_1152 ();
 sg13g2_decap_8 FILLER_76_1159 ();
 sg13g2_decap_8 FILLER_76_1166 ();
 sg13g2_decap_8 FILLER_76_1173 ();
 sg13g2_decap_8 FILLER_76_1180 ();
 sg13g2_decap_8 FILLER_76_1187 ();
 sg13g2_decap_8 FILLER_76_1194 ();
 sg13g2_decap_8 FILLER_76_1201 ();
 sg13g2_decap_8 FILLER_76_1208 ();
 sg13g2_decap_8 FILLER_76_1215 ();
 sg13g2_decap_8 FILLER_76_1222 ();
 sg13g2_decap_8 FILLER_76_1229 ();
 sg13g2_decap_8 FILLER_76_1236 ();
 sg13g2_decap_8 FILLER_76_1243 ();
 sg13g2_decap_8 FILLER_76_1250 ();
 sg13g2_decap_8 FILLER_76_1257 ();
 sg13g2_decap_8 FILLER_76_1264 ();
 sg13g2_decap_8 FILLER_76_1271 ();
 sg13g2_decap_8 FILLER_76_1278 ();
 sg13g2_decap_8 FILLER_76_1285 ();
 sg13g2_decap_8 FILLER_76_1292 ();
 sg13g2_decap_8 FILLER_76_1299 ();
 sg13g2_decap_8 FILLER_76_1306 ();
 sg13g2_decap_8 FILLER_76_1313 ();
 sg13g2_decap_8 FILLER_76_1320 ();
 sg13g2_decap_8 FILLER_76_1327 ();
 sg13g2_decap_8 FILLER_76_1334 ();
 sg13g2_decap_8 FILLER_76_1341 ();
 sg13g2_decap_8 FILLER_76_1348 ();
 sg13g2_decap_8 FILLER_76_1355 ();
 sg13g2_decap_8 FILLER_76_1362 ();
 sg13g2_decap_8 FILLER_76_1369 ();
 sg13g2_decap_8 FILLER_76_1376 ();
 sg13g2_decap_8 FILLER_76_1383 ();
 sg13g2_decap_8 FILLER_76_1390 ();
 sg13g2_decap_8 FILLER_76_1397 ();
 sg13g2_decap_8 FILLER_76_1404 ();
 sg13g2_decap_8 FILLER_76_1411 ();
 sg13g2_decap_8 FILLER_76_1418 ();
 sg13g2_decap_8 FILLER_76_1425 ();
 sg13g2_decap_8 FILLER_76_1432 ();
 sg13g2_decap_8 FILLER_76_1439 ();
 sg13g2_decap_8 FILLER_76_1446 ();
 sg13g2_decap_8 FILLER_76_1453 ();
 sg13g2_decap_8 FILLER_76_1460 ();
 sg13g2_decap_8 FILLER_76_1467 ();
 sg13g2_decap_8 FILLER_76_1474 ();
 sg13g2_decap_8 FILLER_76_1481 ();
 sg13g2_decap_8 FILLER_76_1488 ();
 sg13g2_decap_8 FILLER_76_1495 ();
 sg13g2_decap_8 FILLER_76_1502 ();
 sg13g2_decap_8 FILLER_76_1509 ();
 sg13g2_decap_8 FILLER_76_1516 ();
 sg13g2_decap_8 FILLER_76_1523 ();
 sg13g2_decap_8 FILLER_76_1530 ();
 sg13g2_decap_8 FILLER_76_1537 ();
 sg13g2_decap_8 FILLER_76_1544 ();
 sg13g2_decap_8 FILLER_76_1551 ();
 sg13g2_decap_8 FILLER_76_1558 ();
 sg13g2_decap_8 FILLER_76_1565 ();
 sg13g2_decap_8 FILLER_76_1572 ();
 sg13g2_decap_8 FILLER_76_1579 ();
 sg13g2_decap_8 FILLER_76_1586 ();
 sg13g2_decap_8 FILLER_76_1593 ();
 sg13g2_decap_8 FILLER_76_1600 ();
 sg13g2_decap_8 FILLER_76_1607 ();
 sg13g2_decap_8 FILLER_76_1614 ();
 sg13g2_decap_8 FILLER_76_1621 ();
 sg13g2_decap_8 FILLER_76_1628 ();
 sg13g2_decap_8 FILLER_76_1635 ();
 sg13g2_decap_8 FILLER_76_1642 ();
 sg13g2_decap_8 FILLER_76_1649 ();
 sg13g2_decap_8 FILLER_76_1656 ();
 sg13g2_decap_8 FILLER_76_1663 ();
 sg13g2_decap_8 FILLER_76_1670 ();
 sg13g2_decap_8 FILLER_76_1677 ();
 sg13g2_decap_8 FILLER_76_1684 ();
 sg13g2_decap_8 FILLER_76_1691 ();
 sg13g2_decap_8 FILLER_76_1698 ();
 sg13g2_decap_8 FILLER_76_1705 ();
 sg13g2_decap_8 FILLER_76_1712 ();
 sg13g2_decap_8 FILLER_76_1719 ();
 sg13g2_decap_8 FILLER_76_1726 ();
 sg13g2_decap_8 FILLER_76_1733 ();
 sg13g2_decap_8 FILLER_76_1740 ();
 sg13g2_decap_8 FILLER_76_1747 ();
 sg13g2_decap_8 FILLER_76_1754 ();
 sg13g2_decap_8 FILLER_76_1761 ();
 sg13g2_decap_8 FILLER_76_1768 ();
 sg13g2_decap_8 FILLER_76_1775 ();
 sg13g2_decap_8 FILLER_76_1782 ();
 sg13g2_decap_8 FILLER_76_1789 ();
 sg13g2_decap_8 FILLER_76_1796 ();
 sg13g2_decap_8 FILLER_76_1803 ();
 sg13g2_decap_8 FILLER_76_1810 ();
 sg13g2_decap_8 FILLER_76_1817 ();
 sg13g2_decap_8 FILLER_76_1824 ();
 sg13g2_decap_8 FILLER_76_1831 ();
 sg13g2_decap_8 FILLER_76_1838 ();
 sg13g2_decap_8 FILLER_76_1845 ();
 sg13g2_decap_8 FILLER_76_1852 ();
 sg13g2_decap_8 FILLER_76_1859 ();
 sg13g2_decap_8 FILLER_76_1866 ();
 sg13g2_decap_8 FILLER_76_1873 ();
 sg13g2_decap_8 FILLER_76_1880 ();
 sg13g2_decap_8 FILLER_76_1887 ();
 sg13g2_decap_8 FILLER_76_1894 ();
 sg13g2_decap_8 FILLER_76_1901 ();
 sg13g2_decap_8 FILLER_76_1908 ();
 sg13g2_decap_8 FILLER_76_1915 ();
 sg13g2_decap_8 FILLER_76_1922 ();
 sg13g2_decap_8 FILLER_76_1929 ();
 sg13g2_decap_8 FILLER_76_1936 ();
 sg13g2_decap_8 FILLER_76_1943 ();
 sg13g2_decap_8 FILLER_76_1950 ();
 sg13g2_decap_8 FILLER_76_1957 ();
 sg13g2_decap_8 FILLER_76_1964 ();
 sg13g2_decap_8 FILLER_76_1971 ();
 sg13g2_decap_8 FILLER_76_1978 ();
 sg13g2_decap_8 FILLER_76_1985 ();
 sg13g2_decap_8 FILLER_76_1992 ();
 sg13g2_decap_8 FILLER_76_1999 ();
 sg13g2_decap_8 FILLER_76_2006 ();
 sg13g2_decap_8 FILLER_76_2013 ();
 sg13g2_decap_8 FILLER_76_2020 ();
 sg13g2_decap_8 FILLER_76_2027 ();
 sg13g2_decap_8 FILLER_76_2034 ();
 sg13g2_decap_8 FILLER_76_2041 ();
 sg13g2_decap_8 FILLER_76_2048 ();
 sg13g2_decap_8 FILLER_76_2055 ();
 sg13g2_decap_8 FILLER_76_2062 ();
 sg13g2_decap_8 FILLER_76_2069 ();
 sg13g2_decap_8 FILLER_76_2076 ();
 sg13g2_decap_8 FILLER_76_2083 ();
 sg13g2_decap_8 FILLER_76_2090 ();
 sg13g2_decap_8 FILLER_76_2097 ();
 sg13g2_decap_8 FILLER_76_2104 ();
 sg13g2_decap_8 FILLER_76_2111 ();
 sg13g2_decap_8 FILLER_76_2118 ();
 sg13g2_decap_8 FILLER_76_2125 ();
 sg13g2_decap_8 FILLER_76_2132 ();
 sg13g2_decap_8 FILLER_76_2139 ();
 sg13g2_decap_8 FILLER_76_2146 ();
 sg13g2_decap_8 FILLER_76_2153 ();
 sg13g2_decap_8 FILLER_76_2160 ();
 sg13g2_decap_8 FILLER_76_2167 ();
 sg13g2_decap_8 FILLER_76_2174 ();
 sg13g2_decap_8 FILLER_76_2181 ();
 sg13g2_decap_8 FILLER_76_2188 ();
 sg13g2_decap_8 FILLER_76_2195 ();
 sg13g2_decap_8 FILLER_76_2202 ();
 sg13g2_decap_8 FILLER_76_2209 ();
 sg13g2_decap_8 FILLER_76_2216 ();
 sg13g2_decap_8 FILLER_76_2223 ();
 sg13g2_decap_8 FILLER_76_2230 ();
 sg13g2_decap_8 FILLER_76_2237 ();
 sg13g2_decap_8 FILLER_76_2244 ();
 sg13g2_decap_8 FILLER_76_2251 ();
 sg13g2_decap_8 FILLER_76_2258 ();
 sg13g2_decap_8 FILLER_76_2265 ();
 sg13g2_decap_8 FILLER_76_2272 ();
 sg13g2_decap_8 FILLER_76_2279 ();
 sg13g2_decap_8 FILLER_76_2286 ();
 sg13g2_decap_8 FILLER_76_2293 ();
 sg13g2_decap_8 FILLER_76_2300 ();
 sg13g2_decap_8 FILLER_76_2307 ();
 sg13g2_decap_8 FILLER_76_2314 ();
 sg13g2_decap_8 FILLER_76_2321 ();
 sg13g2_decap_8 FILLER_76_2328 ();
 sg13g2_decap_8 FILLER_76_2335 ();
 sg13g2_decap_8 FILLER_76_2342 ();
 sg13g2_decap_8 FILLER_76_2349 ();
 sg13g2_decap_8 FILLER_76_2356 ();
 sg13g2_decap_8 FILLER_76_2363 ();
 sg13g2_decap_8 FILLER_76_2370 ();
 sg13g2_decap_8 FILLER_76_2377 ();
 sg13g2_decap_8 FILLER_76_2384 ();
 sg13g2_decap_8 FILLER_76_2391 ();
 sg13g2_decap_8 FILLER_76_2398 ();
 sg13g2_decap_8 FILLER_76_2405 ();
 sg13g2_decap_8 FILLER_76_2412 ();
 sg13g2_decap_8 FILLER_76_2419 ();
 sg13g2_decap_8 FILLER_76_2426 ();
 sg13g2_decap_8 FILLER_76_2433 ();
 sg13g2_decap_8 FILLER_76_2440 ();
 sg13g2_decap_8 FILLER_76_2447 ();
 sg13g2_decap_8 FILLER_76_2454 ();
 sg13g2_decap_8 FILLER_76_2461 ();
 sg13g2_decap_8 FILLER_76_2468 ();
 sg13g2_decap_8 FILLER_76_2475 ();
 sg13g2_decap_8 FILLER_76_2482 ();
 sg13g2_decap_8 FILLER_76_2489 ();
 sg13g2_decap_8 FILLER_76_2496 ();
 sg13g2_decap_8 FILLER_76_2503 ();
 sg13g2_decap_8 FILLER_76_2510 ();
 sg13g2_decap_8 FILLER_76_2517 ();
 sg13g2_decap_8 FILLER_76_2524 ();
 sg13g2_decap_8 FILLER_76_2531 ();
 sg13g2_decap_8 FILLER_76_2538 ();
 sg13g2_decap_8 FILLER_76_2545 ();
 sg13g2_decap_8 FILLER_76_2552 ();
 sg13g2_decap_8 FILLER_76_2559 ();
 sg13g2_decap_8 FILLER_76_2566 ();
 sg13g2_decap_8 FILLER_76_2573 ();
 sg13g2_decap_8 FILLER_76_2580 ();
 sg13g2_decap_8 FILLER_76_2587 ();
 sg13g2_decap_8 FILLER_76_2594 ();
 sg13g2_decap_8 FILLER_76_2601 ();
 sg13g2_decap_8 FILLER_76_2608 ();
 sg13g2_decap_8 FILLER_76_2615 ();
 sg13g2_decap_8 FILLER_76_2622 ();
 sg13g2_decap_8 FILLER_76_2629 ();
 sg13g2_decap_8 FILLER_76_2636 ();
 sg13g2_decap_8 FILLER_76_2643 ();
 sg13g2_decap_8 FILLER_76_2650 ();
 sg13g2_decap_8 FILLER_76_2657 ();
 sg13g2_decap_8 FILLER_76_2664 ();
 sg13g2_decap_8 FILLER_76_2671 ();
 sg13g2_decap_8 FILLER_76_2678 ();
 sg13g2_decap_8 FILLER_76_2685 ();
 sg13g2_decap_8 FILLER_76_2692 ();
 sg13g2_decap_8 FILLER_76_2699 ();
 sg13g2_decap_8 FILLER_76_2706 ();
 sg13g2_decap_8 FILLER_76_2713 ();
 sg13g2_decap_8 FILLER_76_2720 ();
 sg13g2_decap_8 FILLER_76_2727 ();
 sg13g2_decap_8 FILLER_76_2734 ();
 sg13g2_decap_8 FILLER_76_2741 ();
 sg13g2_decap_8 FILLER_76_2748 ();
 sg13g2_decap_8 FILLER_76_2755 ();
 sg13g2_decap_8 FILLER_76_2762 ();
 sg13g2_decap_8 FILLER_76_2769 ();
 sg13g2_decap_8 FILLER_76_2776 ();
 sg13g2_decap_8 FILLER_76_2783 ();
 sg13g2_decap_8 FILLER_76_2790 ();
 sg13g2_decap_8 FILLER_76_2797 ();
 sg13g2_decap_8 FILLER_76_2804 ();
 sg13g2_decap_8 FILLER_76_2811 ();
 sg13g2_decap_8 FILLER_76_2818 ();
 sg13g2_decap_8 FILLER_76_2825 ();
 sg13g2_decap_8 FILLER_76_2832 ();
 sg13g2_decap_8 FILLER_76_2839 ();
 sg13g2_decap_8 FILLER_76_2846 ();
 sg13g2_decap_8 FILLER_76_2853 ();
 sg13g2_decap_8 FILLER_76_2860 ();
 sg13g2_decap_8 FILLER_76_2867 ();
 sg13g2_decap_8 FILLER_76_2874 ();
 sg13g2_decap_8 FILLER_76_2881 ();
 sg13g2_decap_8 FILLER_76_2888 ();
 sg13g2_decap_8 FILLER_76_2895 ();
 sg13g2_decap_8 FILLER_76_2902 ();
 sg13g2_decap_8 FILLER_76_2909 ();
 sg13g2_decap_8 FILLER_76_2916 ();
 sg13g2_decap_8 FILLER_76_2923 ();
 sg13g2_decap_8 FILLER_76_2930 ();
 sg13g2_decap_8 FILLER_76_2937 ();
 sg13g2_decap_8 FILLER_76_2944 ();
 sg13g2_decap_8 FILLER_76_2951 ();
 sg13g2_decap_8 FILLER_76_2958 ();
 sg13g2_decap_8 FILLER_76_2965 ();
 sg13g2_decap_8 FILLER_76_2972 ();
 sg13g2_decap_8 FILLER_76_2979 ();
 sg13g2_decap_8 FILLER_76_2986 ();
 sg13g2_decap_8 FILLER_76_2993 ();
 sg13g2_decap_8 FILLER_76_3000 ();
 sg13g2_decap_8 FILLER_76_3007 ();
 sg13g2_decap_8 FILLER_76_3014 ();
 sg13g2_decap_8 FILLER_76_3021 ();
 sg13g2_decap_8 FILLER_76_3028 ();
 sg13g2_decap_8 FILLER_76_3035 ();
 sg13g2_decap_8 FILLER_76_3042 ();
 sg13g2_decap_8 FILLER_76_3049 ();
 sg13g2_decap_8 FILLER_76_3056 ();
 sg13g2_decap_8 FILLER_76_3063 ();
 sg13g2_decap_8 FILLER_76_3070 ();
 sg13g2_decap_8 FILLER_76_3077 ();
 sg13g2_decap_8 FILLER_76_3084 ();
 sg13g2_decap_8 FILLER_76_3091 ();
 sg13g2_decap_8 FILLER_76_3098 ();
 sg13g2_decap_8 FILLER_76_3105 ();
 sg13g2_decap_8 FILLER_76_3112 ();
 sg13g2_decap_8 FILLER_76_3119 ();
 sg13g2_decap_8 FILLER_76_3126 ();
 sg13g2_decap_8 FILLER_76_3133 ();
 sg13g2_decap_8 FILLER_76_3140 ();
 sg13g2_decap_8 FILLER_76_3147 ();
 sg13g2_decap_8 FILLER_76_3154 ();
 sg13g2_decap_8 FILLER_76_3161 ();
 sg13g2_decap_8 FILLER_76_3168 ();
 sg13g2_decap_8 FILLER_76_3175 ();
 sg13g2_decap_8 FILLER_76_3182 ();
 sg13g2_decap_8 FILLER_76_3189 ();
 sg13g2_decap_8 FILLER_76_3196 ();
 sg13g2_decap_8 FILLER_76_3203 ();
 sg13g2_decap_8 FILLER_76_3210 ();
 sg13g2_decap_8 FILLER_76_3217 ();
 sg13g2_decap_8 FILLER_76_3224 ();
 sg13g2_decap_8 FILLER_76_3231 ();
 sg13g2_decap_8 FILLER_76_3238 ();
 sg13g2_decap_8 FILLER_76_3245 ();
 sg13g2_decap_8 FILLER_76_3252 ();
 sg13g2_decap_8 FILLER_76_3259 ();
 sg13g2_decap_8 FILLER_76_3266 ();
 sg13g2_decap_8 FILLER_76_3273 ();
 sg13g2_decap_8 FILLER_76_3280 ();
 sg13g2_decap_8 FILLER_76_3287 ();
 sg13g2_decap_8 FILLER_76_3294 ();
 sg13g2_decap_8 FILLER_76_3301 ();
 sg13g2_decap_8 FILLER_76_3308 ();
 sg13g2_decap_8 FILLER_76_3315 ();
 sg13g2_decap_8 FILLER_76_3322 ();
 sg13g2_decap_8 FILLER_76_3329 ();
 sg13g2_decap_8 FILLER_76_3336 ();
 sg13g2_decap_8 FILLER_76_3343 ();
 sg13g2_decap_8 FILLER_76_3350 ();
 sg13g2_decap_8 FILLER_76_3357 ();
 sg13g2_decap_8 FILLER_76_3364 ();
 sg13g2_decap_8 FILLER_76_3371 ();
 sg13g2_decap_8 FILLER_76_3378 ();
 sg13g2_decap_8 FILLER_76_3385 ();
 sg13g2_decap_8 FILLER_76_3392 ();
 sg13g2_decap_8 FILLER_76_3399 ();
 sg13g2_decap_8 FILLER_76_3406 ();
 sg13g2_decap_8 FILLER_76_3413 ();
 sg13g2_decap_8 FILLER_76_3420 ();
 sg13g2_decap_8 FILLER_76_3427 ();
 sg13g2_decap_8 FILLER_76_3434 ();
 sg13g2_decap_8 FILLER_76_3441 ();
 sg13g2_decap_8 FILLER_76_3448 ();
 sg13g2_decap_8 FILLER_76_3455 ();
 sg13g2_decap_8 FILLER_76_3462 ();
 sg13g2_decap_8 FILLER_76_3469 ();
 sg13g2_decap_8 FILLER_76_3476 ();
 sg13g2_decap_8 FILLER_76_3483 ();
 sg13g2_decap_8 FILLER_76_3490 ();
 sg13g2_decap_8 FILLER_76_3497 ();
 sg13g2_decap_8 FILLER_76_3504 ();
 sg13g2_decap_8 FILLER_76_3511 ();
 sg13g2_decap_8 FILLER_76_3518 ();
 sg13g2_decap_8 FILLER_76_3525 ();
 sg13g2_decap_8 FILLER_76_3532 ();
 sg13g2_decap_8 FILLER_76_3539 ();
 sg13g2_decap_8 FILLER_76_3546 ();
 sg13g2_decap_8 FILLER_76_3553 ();
 sg13g2_decap_8 FILLER_76_3560 ();
 sg13g2_decap_8 FILLER_76_3567 ();
 sg13g2_decap_4 FILLER_76_3574 ();
 sg13g2_fill_2 FILLER_76_3578 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_161 ();
 sg13g2_decap_8 FILLER_77_168 ();
 sg13g2_decap_8 FILLER_77_175 ();
 sg13g2_decap_8 FILLER_77_182 ();
 sg13g2_decap_8 FILLER_77_189 ();
 sg13g2_decap_8 FILLER_77_196 ();
 sg13g2_decap_8 FILLER_77_203 ();
 sg13g2_decap_8 FILLER_77_210 ();
 sg13g2_decap_8 FILLER_77_217 ();
 sg13g2_decap_8 FILLER_77_224 ();
 sg13g2_decap_8 FILLER_77_231 ();
 sg13g2_decap_8 FILLER_77_238 ();
 sg13g2_decap_8 FILLER_77_245 ();
 sg13g2_decap_8 FILLER_77_252 ();
 sg13g2_decap_8 FILLER_77_259 ();
 sg13g2_decap_8 FILLER_77_266 ();
 sg13g2_decap_8 FILLER_77_273 ();
 sg13g2_decap_8 FILLER_77_280 ();
 sg13g2_decap_8 FILLER_77_287 ();
 sg13g2_decap_8 FILLER_77_294 ();
 sg13g2_decap_8 FILLER_77_301 ();
 sg13g2_decap_8 FILLER_77_308 ();
 sg13g2_decap_8 FILLER_77_315 ();
 sg13g2_decap_8 FILLER_77_322 ();
 sg13g2_decap_8 FILLER_77_329 ();
 sg13g2_decap_8 FILLER_77_336 ();
 sg13g2_decap_8 FILLER_77_343 ();
 sg13g2_decap_8 FILLER_77_350 ();
 sg13g2_decap_8 FILLER_77_357 ();
 sg13g2_decap_8 FILLER_77_364 ();
 sg13g2_decap_8 FILLER_77_371 ();
 sg13g2_decap_8 FILLER_77_378 ();
 sg13g2_decap_8 FILLER_77_385 ();
 sg13g2_decap_8 FILLER_77_392 ();
 sg13g2_decap_8 FILLER_77_399 ();
 sg13g2_decap_8 FILLER_77_406 ();
 sg13g2_decap_8 FILLER_77_413 ();
 sg13g2_decap_8 FILLER_77_420 ();
 sg13g2_decap_8 FILLER_77_427 ();
 sg13g2_decap_8 FILLER_77_434 ();
 sg13g2_decap_8 FILLER_77_441 ();
 sg13g2_decap_8 FILLER_77_448 ();
 sg13g2_decap_8 FILLER_77_455 ();
 sg13g2_decap_8 FILLER_77_462 ();
 sg13g2_decap_8 FILLER_77_469 ();
 sg13g2_decap_8 FILLER_77_476 ();
 sg13g2_decap_8 FILLER_77_483 ();
 sg13g2_decap_8 FILLER_77_490 ();
 sg13g2_decap_8 FILLER_77_497 ();
 sg13g2_decap_8 FILLER_77_504 ();
 sg13g2_decap_8 FILLER_77_511 ();
 sg13g2_decap_8 FILLER_77_518 ();
 sg13g2_decap_8 FILLER_77_525 ();
 sg13g2_decap_8 FILLER_77_532 ();
 sg13g2_decap_8 FILLER_77_539 ();
 sg13g2_decap_8 FILLER_77_546 ();
 sg13g2_decap_8 FILLER_77_553 ();
 sg13g2_decap_8 FILLER_77_560 ();
 sg13g2_decap_8 FILLER_77_567 ();
 sg13g2_decap_8 FILLER_77_574 ();
 sg13g2_decap_8 FILLER_77_581 ();
 sg13g2_decap_8 FILLER_77_588 ();
 sg13g2_decap_8 FILLER_77_595 ();
 sg13g2_decap_8 FILLER_77_602 ();
 sg13g2_decap_8 FILLER_77_609 ();
 sg13g2_decap_8 FILLER_77_616 ();
 sg13g2_decap_8 FILLER_77_623 ();
 sg13g2_decap_8 FILLER_77_630 ();
 sg13g2_decap_8 FILLER_77_637 ();
 sg13g2_decap_8 FILLER_77_644 ();
 sg13g2_decap_8 FILLER_77_651 ();
 sg13g2_decap_8 FILLER_77_658 ();
 sg13g2_decap_8 FILLER_77_665 ();
 sg13g2_decap_8 FILLER_77_672 ();
 sg13g2_decap_8 FILLER_77_679 ();
 sg13g2_decap_8 FILLER_77_686 ();
 sg13g2_decap_8 FILLER_77_693 ();
 sg13g2_decap_8 FILLER_77_700 ();
 sg13g2_decap_8 FILLER_77_707 ();
 sg13g2_decap_8 FILLER_77_714 ();
 sg13g2_decap_8 FILLER_77_721 ();
 sg13g2_decap_8 FILLER_77_728 ();
 sg13g2_decap_8 FILLER_77_735 ();
 sg13g2_decap_8 FILLER_77_742 ();
 sg13g2_decap_8 FILLER_77_749 ();
 sg13g2_decap_8 FILLER_77_756 ();
 sg13g2_decap_8 FILLER_77_763 ();
 sg13g2_decap_8 FILLER_77_770 ();
 sg13g2_decap_8 FILLER_77_777 ();
 sg13g2_decap_8 FILLER_77_784 ();
 sg13g2_decap_8 FILLER_77_791 ();
 sg13g2_decap_8 FILLER_77_798 ();
 sg13g2_decap_8 FILLER_77_805 ();
 sg13g2_decap_8 FILLER_77_812 ();
 sg13g2_decap_8 FILLER_77_819 ();
 sg13g2_decap_8 FILLER_77_826 ();
 sg13g2_decap_8 FILLER_77_833 ();
 sg13g2_decap_8 FILLER_77_840 ();
 sg13g2_decap_8 FILLER_77_847 ();
 sg13g2_decap_8 FILLER_77_854 ();
 sg13g2_decap_8 FILLER_77_861 ();
 sg13g2_decap_8 FILLER_77_868 ();
 sg13g2_decap_8 FILLER_77_875 ();
 sg13g2_decap_8 FILLER_77_882 ();
 sg13g2_decap_8 FILLER_77_889 ();
 sg13g2_decap_8 FILLER_77_896 ();
 sg13g2_decap_8 FILLER_77_903 ();
 sg13g2_decap_8 FILLER_77_910 ();
 sg13g2_decap_8 FILLER_77_917 ();
 sg13g2_decap_8 FILLER_77_924 ();
 sg13g2_decap_8 FILLER_77_931 ();
 sg13g2_decap_8 FILLER_77_938 ();
 sg13g2_decap_8 FILLER_77_945 ();
 sg13g2_decap_8 FILLER_77_952 ();
 sg13g2_decap_8 FILLER_77_959 ();
 sg13g2_decap_8 FILLER_77_966 ();
 sg13g2_decap_8 FILLER_77_973 ();
 sg13g2_decap_8 FILLER_77_980 ();
 sg13g2_decap_8 FILLER_77_987 ();
 sg13g2_decap_8 FILLER_77_994 ();
 sg13g2_decap_8 FILLER_77_1001 ();
 sg13g2_decap_8 FILLER_77_1008 ();
 sg13g2_decap_8 FILLER_77_1015 ();
 sg13g2_decap_8 FILLER_77_1022 ();
 sg13g2_decap_8 FILLER_77_1029 ();
 sg13g2_decap_8 FILLER_77_1036 ();
 sg13g2_decap_8 FILLER_77_1043 ();
 sg13g2_decap_8 FILLER_77_1050 ();
 sg13g2_decap_8 FILLER_77_1057 ();
 sg13g2_decap_8 FILLER_77_1064 ();
 sg13g2_decap_8 FILLER_77_1071 ();
 sg13g2_decap_8 FILLER_77_1078 ();
 sg13g2_decap_8 FILLER_77_1085 ();
 sg13g2_decap_8 FILLER_77_1092 ();
 sg13g2_decap_8 FILLER_77_1099 ();
 sg13g2_decap_8 FILLER_77_1106 ();
 sg13g2_decap_8 FILLER_77_1113 ();
 sg13g2_decap_8 FILLER_77_1120 ();
 sg13g2_decap_8 FILLER_77_1127 ();
 sg13g2_decap_8 FILLER_77_1134 ();
 sg13g2_decap_8 FILLER_77_1141 ();
 sg13g2_decap_8 FILLER_77_1148 ();
 sg13g2_decap_8 FILLER_77_1155 ();
 sg13g2_decap_8 FILLER_77_1162 ();
 sg13g2_decap_8 FILLER_77_1169 ();
 sg13g2_decap_8 FILLER_77_1176 ();
 sg13g2_decap_8 FILLER_77_1183 ();
 sg13g2_decap_8 FILLER_77_1190 ();
 sg13g2_decap_8 FILLER_77_1197 ();
 sg13g2_decap_8 FILLER_77_1204 ();
 sg13g2_decap_8 FILLER_77_1211 ();
 sg13g2_decap_8 FILLER_77_1218 ();
 sg13g2_decap_8 FILLER_77_1225 ();
 sg13g2_decap_8 FILLER_77_1232 ();
 sg13g2_decap_8 FILLER_77_1239 ();
 sg13g2_decap_8 FILLER_77_1246 ();
 sg13g2_decap_8 FILLER_77_1253 ();
 sg13g2_decap_8 FILLER_77_1260 ();
 sg13g2_decap_8 FILLER_77_1267 ();
 sg13g2_decap_8 FILLER_77_1274 ();
 sg13g2_decap_8 FILLER_77_1281 ();
 sg13g2_decap_8 FILLER_77_1288 ();
 sg13g2_decap_8 FILLER_77_1295 ();
 sg13g2_decap_8 FILLER_77_1302 ();
 sg13g2_decap_8 FILLER_77_1309 ();
 sg13g2_decap_8 FILLER_77_1316 ();
 sg13g2_decap_8 FILLER_77_1323 ();
 sg13g2_decap_8 FILLER_77_1330 ();
 sg13g2_decap_8 FILLER_77_1337 ();
 sg13g2_decap_8 FILLER_77_1344 ();
 sg13g2_decap_8 FILLER_77_1351 ();
 sg13g2_decap_8 FILLER_77_1358 ();
 sg13g2_decap_8 FILLER_77_1365 ();
 sg13g2_decap_8 FILLER_77_1372 ();
 sg13g2_decap_8 FILLER_77_1379 ();
 sg13g2_decap_8 FILLER_77_1386 ();
 sg13g2_decap_8 FILLER_77_1393 ();
 sg13g2_decap_8 FILLER_77_1400 ();
 sg13g2_decap_8 FILLER_77_1407 ();
 sg13g2_decap_8 FILLER_77_1414 ();
 sg13g2_decap_8 FILLER_77_1421 ();
 sg13g2_decap_8 FILLER_77_1428 ();
 sg13g2_decap_8 FILLER_77_1435 ();
 sg13g2_decap_8 FILLER_77_1442 ();
 sg13g2_decap_8 FILLER_77_1449 ();
 sg13g2_decap_8 FILLER_77_1456 ();
 sg13g2_decap_8 FILLER_77_1463 ();
 sg13g2_decap_8 FILLER_77_1470 ();
 sg13g2_decap_8 FILLER_77_1477 ();
 sg13g2_decap_8 FILLER_77_1484 ();
 sg13g2_decap_8 FILLER_77_1491 ();
 sg13g2_decap_8 FILLER_77_1498 ();
 sg13g2_decap_8 FILLER_77_1505 ();
 sg13g2_decap_8 FILLER_77_1512 ();
 sg13g2_decap_8 FILLER_77_1519 ();
 sg13g2_decap_8 FILLER_77_1526 ();
 sg13g2_decap_8 FILLER_77_1533 ();
 sg13g2_decap_8 FILLER_77_1540 ();
 sg13g2_decap_8 FILLER_77_1547 ();
 sg13g2_decap_8 FILLER_77_1554 ();
 sg13g2_decap_8 FILLER_77_1561 ();
 sg13g2_decap_8 FILLER_77_1568 ();
 sg13g2_decap_8 FILLER_77_1575 ();
 sg13g2_decap_8 FILLER_77_1582 ();
 sg13g2_decap_8 FILLER_77_1589 ();
 sg13g2_decap_8 FILLER_77_1596 ();
 sg13g2_decap_8 FILLER_77_1603 ();
 sg13g2_decap_8 FILLER_77_1610 ();
 sg13g2_decap_8 FILLER_77_1617 ();
 sg13g2_decap_8 FILLER_77_1624 ();
 sg13g2_decap_8 FILLER_77_1631 ();
 sg13g2_decap_8 FILLER_77_1638 ();
 sg13g2_decap_8 FILLER_77_1645 ();
 sg13g2_decap_8 FILLER_77_1652 ();
 sg13g2_decap_8 FILLER_77_1659 ();
 sg13g2_decap_8 FILLER_77_1666 ();
 sg13g2_decap_8 FILLER_77_1673 ();
 sg13g2_decap_8 FILLER_77_1680 ();
 sg13g2_decap_8 FILLER_77_1687 ();
 sg13g2_decap_8 FILLER_77_1694 ();
 sg13g2_decap_8 FILLER_77_1701 ();
 sg13g2_decap_8 FILLER_77_1708 ();
 sg13g2_decap_8 FILLER_77_1715 ();
 sg13g2_decap_8 FILLER_77_1722 ();
 sg13g2_decap_8 FILLER_77_1729 ();
 sg13g2_decap_8 FILLER_77_1736 ();
 sg13g2_decap_8 FILLER_77_1743 ();
 sg13g2_decap_8 FILLER_77_1750 ();
 sg13g2_decap_8 FILLER_77_1757 ();
 sg13g2_decap_8 FILLER_77_1764 ();
 sg13g2_decap_8 FILLER_77_1771 ();
 sg13g2_decap_8 FILLER_77_1778 ();
 sg13g2_decap_8 FILLER_77_1785 ();
 sg13g2_decap_8 FILLER_77_1792 ();
 sg13g2_decap_8 FILLER_77_1799 ();
 sg13g2_decap_8 FILLER_77_1806 ();
 sg13g2_decap_8 FILLER_77_1813 ();
 sg13g2_decap_8 FILLER_77_1820 ();
 sg13g2_decap_8 FILLER_77_1827 ();
 sg13g2_decap_8 FILLER_77_1834 ();
 sg13g2_decap_8 FILLER_77_1841 ();
 sg13g2_decap_8 FILLER_77_1848 ();
 sg13g2_decap_8 FILLER_77_1855 ();
 sg13g2_decap_8 FILLER_77_1862 ();
 sg13g2_decap_8 FILLER_77_1869 ();
 sg13g2_decap_8 FILLER_77_1876 ();
 sg13g2_decap_8 FILLER_77_1883 ();
 sg13g2_decap_8 FILLER_77_1890 ();
 sg13g2_decap_8 FILLER_77_1897 ();
 sg13g2_decap_8 FILLER_77_1904 ();
 sg13g2_decap_8 FILLER_77_1911 ();
 sg13g2_decap_8 FILLER_77_1918 ();
 sg13g2_decap_8 FILLER_77_1925 ();
 sg13g2_decap_8 FILLER_77_1932 ();
 sg13g2_decap_8 FILLER_77_1939 ();
 sg13g2_decap_8 FILLER_77_1946 ();
 sg13g2_decap_8 FILLER_77_1953 ();
 sg13g2_decap_8 FILLER_77_1960 ();
 sg13g2_decap_8 FILLER_77_1967 ();
 sg13g2_decap_8 FILLER_77_1974 ();
 sg13g2_decap_8 FILLER_77_1981 ();
 sg13g2_decap_8 FILLER_77_1988 ();
 sg13g2_decap_8 FILLER_77_1995 ();
 sg13g2_decap_8 FILLER_77_2002 ();
 sg13g2_decap_8 FILLER_77_2009 ();
 sg13g2_decap_8 FILLER_77_2016 ();
 sg13g2_decap_8 FILLER_77_2023 ();
 sg13g2_decap_8 FILLER_77_2030 ();
 sg13g2_decap_8 FILLER_77_2037 ();
 sg13g2_decap_8 FILLER_77_2044 ();
 sg13g2_decap_8 FILLER_77_2051 ();
 sg13g2_decap_8 FILLER_77_2058 ();
 sg13g2_decap_8 FILLER_77_2065 ();
 sg13g2_decap_8 FILLER_77_2072 ();
 sg13g2_decap_8 FILLER_77_2079 ();
 sg13g2_decap_8 FILLER_77_2086 ();
 sg13g2_decap_8 FILLER_77_2093 ();
 sg13g2_decap_8 FILLER_77_2100 ();
 sg13g2_decap_8 FILLER_77_2107 ();
 sg13g2_decap_8 FILLER_77_2114 ();
 sg13g2_decap_8 FILLER_77_2121 ();
 sg13g2_decap_8 FILLER_77_2128 ();
 sg13g2_decap_8 FILLER_77_2135 ();
 sg13g2_decap_8 FILLER_77_2142 ();
 sg13g2_decap_8 FILLER_77_2149 ();
 sg13g2_decap_8 FILLER_77_2156 ();
 sg13g2_decap_8 FILLER_77_2163 ();
 sg13g2_decap_8 FILLER_77_2170 ();
 sg13g2_decap_8 FILLER_77_2177 ();
 sg13g2_decap_8 FILLER_77_2184 ();
 sg13g2_decap_8 FILLER_77_2191 ();
 sg13g2_decap_8 FILLER_77_2198 ();
 sg13g2_decap_8 FILLER_77_2205 ();
 sg13g2_decap_8 FILLER_77_2212 ();
 sg13g2_decap_8 FILLER_77_2219 ();
 sg13g2_decap_8 FILLER_77_2226 ();
 sg13g2_decap_8 FILLER_77_2233 ();
 sg13g2_decap_8 FILLER_77_2240 ();
 sg13g2_decap_8 FILLER_77_2247 ();
 sg13g2_decap_8 FILLER_77_2254 ();
 sg13g2_decap_8 FILLER_77_2261 ();
 sg13g2_decap_8 FILLER_77_2268 ();
 sg13g2_decap_8 FILLER_77_2275 ();
 sg13g2_decap_8 FILLER_77_2282 ();
 sg13g2_decap_8 FILLER_77_2289 ();
 sg13g2_decap_8 FILLER_77_2296 ();
 sg13g2_decap_8 FILLER_77_2303 ();
 sg13g2_decap_8 FILLER_77_2310 ();
 sg13g2_decap_8 FILLER_77_2317 ();
 sg13g2_decap_8 FILLER_77_2324 ();
 sg13g2_decap_8 FILLER_77_2331 ();
 sg13g2_decap_8 FILLER_77_2338 ();
 sg13g2_decap_8 FILLER_77_2345 ();
 sg13g2_decap_8 FILLER_77_2352 ();
 sg13g2_decap_8 FILLER_77_2359 ();
 sg13g2_decap_8 FILLER_77_2366 ();
 sg13g2_decap_8 FILLER_77_2373 ();
 sg13g2_decap_8 FILLER_77_2380 ();
 sg13g2_decap_8 FILLER_77_2387 ();
 sg13g2_decap_8 FILLER_77_2394 ();
 sg13g2_decap_8 FILLER_77_2401 ();
 sg13g2_decap_8 FILLER_77_2408 ();
 sg13g2_decap_8 FILLER_77_2415 ();
 sg13g2_decap_8 FILLER_77_2422 ();
 sg13g2_decap_8 FILLER_77_2429 ();
 sg13g2_decap_8 FILLER_77_2436 ();
 sg13g2_decap_8 FILLER_77_2443 ();
 sg13g2_decap_8 FILLER_77_2450 ();
 sg13g2_decap_8 FILLER_77_2457 ();
 sg13g2_decap_8 FILLER_77_2464 ();
 sg13g2_decap_8 FILLER_77_2471 ();
 sg13g2_decap_8 FILLER_77_2478 ();
 sg13g2_decap_8 FILLER_77_2485 ();
 sg13g2_decap_8 FILLER_77_2492 ();
 sg13g2_decap_8 FILLER_77_2499 ();
 sg13g2_decap_8 FILLER_77_2506 ();
 sg13g2_decap_8 FILLER_77_2513 ();
 sg13g2_decap_8 FILLER_77_2520 ();
 sg13g2_decap_8 FILLER_77_2527 ();
 sg13g2_decap_8 FILLER_77_2534 ();
 sg13g2_decap_8 FILLER_77_2541 ();
 sg13g2_decap_8 FILLER_77_2548 ();
 sg13g2_decap_8 FILLER_77_2555 ();
 sg13g2_decap_8 FILLER_77_2562 ();
 sg13g2_decap_8 FILLER_77_2569 ();
 sg13g2_decap_8 FILLER_77_2576 ();
 sg13g2_decap_8 FILLER_77_2583 ();
 sg13g2_decap_8 FILLER_77_2590 ();
 sg13g2_decap_8 FILLER_77_2597 ();
 sg13g2_decap_8 FILLER_77_2604 ();
 sg13g2_decap_8 FILLER_77_2611 ();
 sg13g2_decap_8 FILLER_77_2618 ();
 sg13g2_decap_8 FILLER_77_2625 ();
 sg13g2_decap_8 FILLER_77_2632 ();
 sg13g2_decap_8 FILLER_77_2639 ();
 sg13g2_decap_8 FILLER_77_2646 ();
 sg13g2_decap_8 FILLER_77_2653 ();
 sg13g2_decap_8 FILLER_77_2660 ();
 sg13g2_decap_8 FILLER_77_2667 ();
 sg13g2_decap_8 FILLER_77_2674 ();
 sg13g2_decap_8 FILLER_77_2681 ();
 sg13g2_decap_8 FILLER_77_2688 ();
 sg13g2_decap_8 FILLER_77_2695 ();
 sg13g2_decap_8 FILLER_77_2702 ();
 sg13g2_decap_8 FILLER_77_2709 ();
 sg13g2_decap_8 FILLER_77_2716 ();
 sg13g2_decap_8 FILLER_77_2723 ();
 sg13g2_decap_8 FILLER_77_2730 ();
 sg13g2_decap_8 FILLER_77_2737 ();
 sg13g2_decap_8 FILLER_77_2744 ();
 sg13g2_decap_8 FILLER_77_2751 ();
 sg13g2_decap_8 FILLER_77_2758 ();
 sg13g2_decap_8 FILLER_77_2765 ();
 sg13g2_decap_8 FILLER_77_2772 ();
 sg13g2_decap_8 FILLER_77_2779 ();
 sg13g2_decap_8 FILLER_77_2786 ();
 sg13g2_decap_8 FILLER_77_2793 ();
 sg13g2_decap_8 FILLER_77_2800 ();
 sg13g2_decap_8 FILLER_77_2807 ();
 sg13g2_decap_8 FILLER_77_2814 ();
 sg13g2_decap_8 FILLER_77_2821 ();
 sg13g2_decap_8 FILLER_77_2828 ();
 sg13g2_decap_8 FILLER_77_2835 ();
 sg13g2_decap_8 FILLER_77_2842 ();
 sg13g2_decap_8 FILLER_77_2849 ();
 sg13g2_decap_8 FILLER_77_2856 ();
 sg13g2_decap_8 FILLER_77_2863 ();
 sg13g2_decap_8 FILLER_77_2870 ();
 sg13g2_decap_8 FILLER_77_2877 ();
 sg13g2_decap_8 FILLER_77_2884 ();
 sg13g2_decap_8 FILLER_77_2891 ();
 sg13g2_decap_8 FILLER_77_2898 ();
 sg13g2_decap_8 FILLER_77_2905 ();
 sg13g2_decap_8 FILLER_77_2912 ();
 sg13g2_decap_8 FILLER_77_2919 ();
 sg13g2_decap_8 FILLER_77_2926 ();
 sg13g2_decap_8 FILLER_77_2933 ();
 sg13g2_decap_8 FILLER_77_2940 ();
 sg13g2_decap_8 FILLER_77_2947 ();
 sg13g2_decap_8 FILLER_77_2954 ();
 sg13g2_decap_8 FILLER_77_2961 ();
 sg13g2_decap_8 FILLER_77_2968 ();
 sg13g2_decap_8 FILLER_77_2975 ();
 sg13g2_decap_8 FILLER_77_2982 ();
 sg13g2_decap_8 FILLER_77_2989 ();
 sg13g2_decap_8 FILLER_77_2996 ();
 sg13g2_decap_8 FILLER_77_3003 ();
 sg13g2_decap_8 FILLER_77_3010 ();
 sg13g2_decap_8 FILLER_77_3017 ();
 sg13g2_decap_8 FILLER_77_3024 ();
 sg13g2_decap_8 FILLER_77_3031 ();
 sg13g2_decap_8 FILLER_77_3038 ();
 sg13g2_decap_8 FILLER_77_3045 ();
 sg13g2_decap_8 FILLER_77_3052 ();
 sg13g2_decap_8 FILLER_77_3059 ();
 sg13g2_decap_8 FILLER_77_3066 ();
 sg13g2_decap_8 FILLER_77_3073 ();
 sg13g2_decap_8 FILLER_77_3080 ();
 sg13g2_decap_8 FILLER_77_3087 ();
 sg13g2_decap_8 FILLER_77_3094 ();
 sg13g2_decap_8 FILLER_77_3101 ();
 sg13g2_decap_8 FILLER_77_3108 ();
 sg13g2_decap_8 FILLER_77_3115 ();
 sg13g2_decap_8 FILLER_77_3122 ();
 sg13g2_decap_8 FILLER_77_3129 ();
 sg13g2_decap_8 FILLER_77_3136 ();
 sg13g2_decap_8 FILLER_77_3143 ();
 sg13g2_decap_8 FILLER_77_3150 ();
 sg13g2_decap_8 FILLER_77_3157 ();
 sg13g2_decap_8 FILLER_77_3164 ();
 sg13g2_decap_8 FILLER_77_3171 ();
 sg13g2_decap_8 FILLER_77_3178 ();
 sg13g2_decap_8 FILLER_77_3185 ();
 sg13g2_decap_8 FILLER_77_3192 ();
 sg13g2_decap_8 FILLER_77_3199 ();
 sg13g2_decap_8 FILLER_77_3206 ();
 sg13g2_decap_8 FILLER_77_3213 ();
 sg13g2_decap_8 FILLER_77_3220 ();
 sg13g2_decap_8 FILLER_77_3227 ();
 sg13g2_decap_8 FILLER_77_3234 ();
 sg13g2_decap_8 FILLER_77_3241 ();
 sg13g2_decap_8 FILLER_77_3248 ();
 sg13g2_decap_8 FILLER_77_3255 ();
 sg13g2_decap_8 FILLER_77_3262 ();
 sg13g2_decap_8 FILLER_77_3269 ();
 sg13g2_decap_8 FILLER_77_3276 ();
 sg13g2_decap_8 FILLER_77_3283 ();
 sg13g2_decap_8 FILLER_77_3290 ();
 sg13g2_decap_8 FILLER_77_3297 ();
 sg13g2_decap_8 FILLER_77_3304 ();
 sg13g2_decap_8 FILLER_77_3311 ();
 sg13g2_decap_8 FILLER_77_3318 ();
 sg13g2_decap_8 FILLER_77_3325 ();
 sg13g2_decap_8 FILLER_77_3332 ();
 sg13g2_decap_8 FILLER_77_3339 ();
 sg13g2_decap_8 FILLER_77_3346 ();
 sg13g2_decap_8 FILLER_77_3353 ();
 sg13g2_decap_8 FILLER_77_3360 ();
 sg13g2_decap_8 FILLER_77_3367 ();
 sg13g2_decap_8 FILLER_77_3374 ();
 sg13g2_decap_8 FILLER_77_3381 ();
 sg13g2_decap_8 FILLER_77_3388 ();
 sg13g2_decap_8 FILLER_77_3395 ();
 sg13g2_decap_8 FILLER_77_3402 ();
 sg13g2_decap_8 FILLER_77_3409 ();
 sg13g2_decap_8 FILLER_77_3416 ();
 sg13g2_decap_8 FILLER_77_3423 ();
 sg13g2_decap_8 FILLER_77_3430 ();
 sg13g2_decap_8 FILLER_77_3437 ();
 sg13g2_decap_8 FILLER_77_3444 ();
 sg13g2_decap_8 FILLER_77_3451 ();
 sg13g2_decap_8 FILLER_77_3458 ();
 sg13g2_decap_8 FILLER_77_3465 ();
 sg13g2_decap_8 FILLER_77_3472 ();
 sg13g2_decap_8 FILLER_77_3479 ();
 sg13g2_decap_8 FILLER_77_3486 ();
 sg13g2_decap_8 FILLER_77_3493 ();
 sg13g2_decap_8 FILLER_77_3500 ();
 sg13g2_decap_8 FILLER_77_3507 ();
 sg13g2_decap_8 FILLER_77_3514 ();
 sg13g2_decap_8 FILLER_77_3521 ();
 sg13g2_decap_8 FILLER_77_3528 ();
 sg13g2_decap_8 FILLER_77_3535 ();
 sg13g2_decap_8 FILLER_77_3542 ();
 sg13g2_decap_8 FILLER_77_3549 ();
 sg13g2_decap_8 FILLER_77_3556 ();
 sg13g2_decap_8 FILLER_77_3563 ();
 sg13g2_decap_8 FILLER_77_3570 ();
 sg13g2_fill_2 FILLER_77_3577 ();
 sg13g2_fill_1 FILLER_77_3579 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_8 FILLER_78_154 ();
 sg13g2_decap_8 FILLER_78_161 ();
 sg13g2_decap_8 FILLER_78_168 ();
 sg13g2_decap_8 FILLER_78_175 ();
 sg13g2_decap_8 FILLER_78_182 ();
 sg13g2_decap_8 FILLER_78_189 ();
 sg13g2_decap_8 FILLER_78_196 ();
 sg13g2_decap_8 FILLER_78_203 ();
 sg13g2_decap_8 FILLER_78_210 ();
 sg13g2_decap_8 FILLER_78_217 ();
 sg13g2_decap_8 FILLER_78_224 ();
 sg13g2_decap_8 FILLER_78_231 ();
 sg13g2_decap_8 FILLER_78_238 ();
 sg13g2_decap_8 FILLER_78_245 ();
 sg13g2_decap_8 FILLER_78_252 ();
 sg13g2_decap_8 FILLER_78_259 ();
 sg13g2_decap_8 FILLER_78_266 ();
 sg13g2_decap_8 FILLER_78_273 ();
 sg13g2_decap_8 FILLER_78_280 ();
 sg13g2_decap_8 FILLER_78_287 ();
 sg13g2_decap_8 FILLER_78_294 ();
 sg13g2_decap_8 FILLER_78_301 ();
 sg13g2_decap_8 FILLER_78_308 ();
 sg13g2_decap_8 FILLER_78_315 ();
 sg13g2_decap_8 FILLER_78_322 ();
 sg13g2_decap_8 FILLER_78_329 ();
 sg13g2_decap_8 FILLER_78_336 ();
 sg13g2_decap_8 FILLER_78_343 ();
 sg13g2_decap_8 FILLER_78_350 ();
 sg13g2_decap_8 FILLER_78_357 ();
 sg13g2_decap_8 FILLER_78_364 ();
 sg13g2_decap_8 FILLER_78_371 ();
 sg13g2_decap_8 FILLER_78_378 ();
 sg13g2_decap_8 FILLER_78_385 ();
 sg13g2_decap_8 FILLER_78_392 ();
 sg13g2_decap_8 FILLER_78_399 ();
 sg13g2_decap_8 FILLER_78_406 ();
 sg13g2_decap_8 FILLER_78_413 ();
 sg13g2_decap_8 FILLER_78_420 ();
 sg13g2_decap_8 FILLER_78_427 ();
 sg13g2_decap_8 FILLER_78_434 ();
 sg13g2_decap_8 FILLER_78_441 ();
 sg13g2_decap_8 FILLER_78_448 ();
 sg13g2_decap_8 FILLER_78_455 ();
 sg13g2_decap_8 FILLER_78_462 ();
 sg13g2_decap_8 FILLER_78_469 ();
 sg13g2_decap_8 FILLER_78_476 ();
 sg13g2_decap_8 FILLER_78_483 ();
 sg13g2_decap_8 FILLER_78_490 ();
 sg13g2_decap_8 FILLER_78_497 ();
 sg13g2_decap_8 FILLER_78_504 ();
 sg13g2_decap_8 FILLER_78_511 ();
 sg13g2_decap_8 FILLER_78_518 ();
 sg13g2_decap_8 FILLER_78_525 ();
 sg13g2_decap_8 FILLER_78_532 ();
 sg13g2_decap_8 FILLER_78_539 ();
 sg13g2_decap_8 FILLER_78_546 ();
 sg13g2_decap_8 FILLER_78_553 ();
 sg13g2_decap_8 FILLER_78_560 ();
 sg13g2_decap_8 FILLER_78_567 ();
 sg13g2_decap_8 FILLER_78_574 ();
 sg13g2_decap_8 FILLER_78_581 ();
 sg13g2_decap_8 FILLER_78_588 ();
 sg13g2_decap_8 FILLER_78_595 ();
 sg13g2_decap_8 FILLER_78_602 ();
 sg13g2_decap_8 FILLER_78_609 ();
 sg13g2_decap_8 FILLER_78_616 ();
 sg13g2_decap_8 FILLER_78_623 ();
 sg13g2_decap_8 FILLER_78_630 ();
 sg13g2_decap_8 FILLER_78_637 ();
 sg13g2_decap_8 FILLER_78_644 ();
 sg13g2_decap_8 FILLER_78_651 ();
 sg13g2_decap_8 FILLER_78_658 ();
 sg13g2_decap_8 FILLER_78_665 ();
 sg13g2_decap_8 FILLER_78_672 ();
 sg13g2_decap_8 FILLER_78_679 ();
 sg13g2_decap_8 FILLER_78_686 ();
 sg13g2_decap_8 FILLER_78_693 ();
 sg13g2_decap_8 FILLER_78_700 ();
 sg13g2_decap_8 FILLER_78_707 ();
 sg13g2_decap_8 FILLER_78_714 ();
 sg13g2_decap_8 FILLER_78_721 ();
 sg13g2_decap_8 FILLER_78_728 ();
 sg13g2_decap_8 FILLER_78_735 ();
 sg13g2_decap_8 FILLER_78_742 ();
 sg13g2_decap_8 FILLER_78_749 ();
 sg13g2_decap_8 FILLER_78_756 ();
 sg13g2_decap_8 FILLER_78_763 ();
 sg13g2_decap_8 FILLER_78_770 ();
 sg13g2_decap_8 FILLER_78_777 ();
 sg13g2_decap_8 FILLER_78_784 ();
 sg13g2_decap_8 FILLER_78_791 ();
 sg13g2_decap_8 FILLER_78_798 ();
 sg13g2_decap_8 FILLER_78_805 ();
 sg13g2_decap_8 FILLER_78_812 ();
 sg13g2_decap_8 FILLER_78_819 ();
 sg13g2_decap_8 FILLER_78_826 ();
 sg13g2_decap_8 FILLER_78_833 ();
 sg13g2_decap_8 FILLER_78_840 ();
 sg13g2_decap_8 FILLER_78_847 ();
 sg13g2_decap_8 FILLER_78_854 ();
 sg13g2_decap_8 FILLER_78_861 ();
 sg13g2_decap_8 FILLER_78_868 ();
 sg13g2_decap_8 FILLER_78_875 ();
 sg13g2_decap_8 FILLER_78_882 ();
 sg13g2_decap_8 FILLER_78_889 ();
 sg13g2_decap_8 FILLER_78_896 ();
 sg13g2_decap_8 FILLER_78_903 ();
 sg13g2_decap_8 FILLER_78_910 ();
 sg13g2_decap_8 FILLER_78_917 ();
 sg13g2_decap_8 FILLER_78_924 ();
 sg13g2_decap_8 FILLER_78_931 ();
 sg13g2_decap_8 FILLER_78_938 ();
 sg13g2_decap_8 FILLER_78_945 ();
 sg13g2_decap_8 FILLER_78_952 ();
 sg13g2_decap_8 FILLER_78_959 ();
 sg13g2_decap_8 FILLER_78_966 ();
 sg13g2_decap_8 FILLER_78_973 ();
 sg13g2_decap_8 FILLER_78_980 ();
 sg13g2_decap_8 FILLER_78_987 ();
 sg13g2_decap_8 FILLER_78_994 ();
 sg13g2_decap_8 FILLER_78_1001 ();
 sg13g2_decap_8 FILLER_78_1008 ();
 sg13g2_decap_8 FILLER_78_1015 ();
 sg13g2_decap_8 FILLER_78_1022 ();
 sg13g2_decap_8 FILLER_78_1029 ();
 sg13g2_decap_8 FILLER_78_1036 ();
 sg13g2_decap_8 FILLER_78_1043 ();
 sg13g2_decap_8 FILLER_78_1050 ();
 sg13g2_decap_8 FILLER_78_1057 ();
 sg13g2_decap_8 FILLER_78_1064 ();
 sg13g2_decap_8 FILLER_78_1071 ();
 sg13g2_decap_8 FILLER_78_1078 ();
 sg13g2_decap_8 FILLER_78_1085 ();
 sg13g2_decap_8 FILLER_78_1092 ();
 sg13g2_decap_8 FILLER_78_1099 ();
 sg13g2_decap_8 FILLER_78_1106 ();
 sg13g2_decap_8 FILLER_78_1113 ();
 sg13g2_decap_8 FILLER_78_1120 ();
 sg13g2_decap_8 FILLER_78_1127 ();
 sg13g2_decap_8 FILLER_78_1134 ();
 sg13g2_decap_8 FILLER_78_1141 ();
 sg13g2_decap_8 FILLER_78_1148 ();
 sg13g2_decap_8 FILLER_78_1155 ();
 sg13g2_decap_8 FILLER_78_1162 ();
 sg13g2_decap_8 FILLER_78_1169 ();
 sg13g2_decap_8 FILLER_78_1176 ();
 sg13g2_decap_8 FILLER_78_1183 ();
 sg13g2_decap_8 FILLER_78_1190 ();
 sg13g2_decap_8 FILLER_78_1197 ();
 sg13g2_decap_8 FILLER_78_1204 ();
 sg13g2_decap_8 FILLER_78_1211 ();
 sg13g2_decap_8 FILLER_78_1218 ();
 sg13g2_decap_8 FILLER_78_1225 ();
 sg13g2_decap_8 FILLER_78_1232 ();
 sg13g2_decap_8 FILLER_78_1239 ();
 sg13g2_decap_8 FILLER_78_1246 ();
 sg13g2_decap_8 FILLER_78_1253 ();
 sg13g2_decap_8 FILLER_78_1260 ();
 sg13g2_decap_8 FILLER_78_1267 ();
 sg13g2_decap_8 FILLER_78_1274 ();
 sg13g2_decap_8 FILLER_78_1281 ();
 sg13g2_decap_8 FILLER_78_1288 ();
 sg13g2_decap_8 FILLER_78_1295 ();
 sg13g2_decap_8 FILLER_78_1302 ();
 sg13g2_decap_8 FILLER_78_1309 ();
 sg13g2_decap_8 FILLER_78_1316 ();
 sg13g2_decap_8 FILLER_78_1323 ();
 sg13g2_decap_8 FILLER_78_1330 ();
 sg13g2_decap_8 FILLER_78_1337 ();
 sg13g2_decap_8 FILLER_78_1344 ();
 sg13g2_decap_8 FILLER_78_1351 ();
 sg13g2_decap_8 FILLER_78_1358 ();
 sg13g2_decap_8 FILLER_78_1365 ();
 sg13g2_decap_8 FILLER_78_1372 ();
 sg13g2_decap_8 FILLER_78_1379 ();
 sg13g2_decap_8 FILLER_78_1386 ();
 sg13g2_decap_8 FILLER_78_1393 ();
 sg13g2_decap_8 FILLER_78_1400 ();
 sg13g2_decap_8 FILLER_78_1407 ();
 sg13g2_decap_8 FILLER_78_1414 ();
 sg13g2_decap_8 FILLER_78_1421 ();
 sg13g2_decap_8 FILLER_78_1428 ();
 sg13g2_decap_8 FILLER_78_1435 ();
 sg13g2_decap_8 FILLER_78_1442 ();
 sg13g2_decap_8 FILLER_78_1449 ();
 sg13g2_decap_8 FILLER_78_1456 ();
 sg13g2_decap_8 FILLER_78_1463 ();
 sg13g2_decap_8 FILLER_78_1470 ();
 sg13g2_decap_8 FILLER_78_1477 ();
 sg13g2_decap_8 FILLER_78_1484 ();
 sg13g2_decap_8 FILLER_78_1491 ();
 sg13g2_decap_8 FILLER_78_1498 ();
 sg13g2_decap_8 FILLER_78_1505 ();
 sg13g2_decap_8 FILLER_78_1512 ();
 sg13g2_decap_8 FILLER_78_1519 ();
 sg13g2_decap_8 FILLER_78_1526 ();
 sg13g2_decap_8 FILLER_78_1533 ();
 sg13g2_decap_8 FILLER_78_1540 ();
 sg13g2_decap_8 FILLER_78_1547 ();
 sg13g2_decap_8 FILLER_78_1554 ();
 sg13g2_decap_8 FILLER_78_1561 ();
 sg13g2_decap_8 FILLER_78_1568 ();
 sg13g2_decap_8 FILLER_78_1575 ();
 sg13g2_decap_8 FILLER_78_1582 ();
 sg13g2_decap_8 FILLER_78_1589 ();
 sg13g2_decap_8 FILLER_78_1596 ();
 sg13g2_decap_8 FILLER_78_1603 ();
 sg13g2_decap_8 FILLER_78_1610 ();
 sg13g2_decap_8 FILLER_78_1617 ();
 sg13g2_decap_8 FILLER_78_1624 ();
 sg13g2_decap_8 FILLER_78_1631 ();
 sg13g2_decap_8 FILLER_78_1638 ();
 sg13g2_decap_8 FILLER_78_1645 ();
 sg13g2_decap_8 FILLER_78_1652 ();
 sg13g2_decap_8 FILLER_78_1659 ();
 sg13g2_decap_8 FILLER_78_1666 ();
 sg13g2_decap_8 FILLER_78_1673 ();
 sg13g2_decap_8 FILLER_78_1680 ();
 sg13g2_decap_8 FILLER_78_1687 ();
 sg13g2_decap_8 FILLER_78_1694 ();
 sg13g2_decap_8 FILLER_78_1701 ();
 sg13g2_decap_8 FILLER_78_1708 ();
 sg13g2_decap_8 FILLER_78_1715 ();
 sg13g2_decap_8 FILLER_78_1722 ();
 sg13g2_decap_8 FILLER_78_1729 ();
 sg13g2_decap_8 FILLER_78_1736 ();
 sg13g2_decap_8 FILLER_78_1743 ();
 sg13g2_decap_8 FILLER_78_1750 ();
 sg13g2_decap_8 FILLER_78_1757 ();
 sg13g2_decap_8 FILLER_78_1764 ();
 sg13g2_decap_8 FILLER_78_1771 ();
 sg13g2_decap_8 FILLER_78_1778 ();
 sg13g2_decap_8 FILLER_78_1785 ();
 sg13g2_decap_8 FILLER_78_1792 ();
 sg13g2_decap_8 FILLER_78_1799 ();
 sg13g2_decap_8 FILLER_78_1806 ();
 sg13g2_decap_8 FILLER_78_1813 ();
 sg13g2_decap_8 FILLER_78_1820 ();
 sg13g2_decap_8 FILLER_78_1827 ();
 sg13g2_decap_8 FILLER_78_1834 ();
 sg13g2_decap_8 FILLER_78_1841 ();
 sg13g2_decap_8 FILLER_78_1848 ();
 sg13g2_decap_8 FILLER_78_1855 ();
 sg13g2_decap_8 FILLER_78_1862 ();
 sg13g2_decap_8 FILLER_78_1869 ();
 sg13g2_decap_8 FILLER_78_1876 ();
 sg13g2_decap_8 FILLER_78_1883 ();
 sg13g2_decap_8 FILLER_78_1890 ();
 sg13g2_decap_8 FILLER_78_1897 ();
 sg13g2_decap_8 FILLER_78_1904 ();
 sg13g2_decap_8 FILLER_78_1911 ();
 sg13g2_decap_8 FILLER_78_1918 ();
 sg13g2_decap_8 FILLER_78_1925 ();
 sg13g2_decap_8 FILLER_78_1932 ();
 sg13g2_decap_8 FILLER_78_1939 ();
 sg13g2_decap_8 FILLER_78_1946 ();
 sg13g2_decap_8 FILLER_78_1953 ();
 sg13g2_decap_8 FILLER_78_1960 ();
 sg13g2_decap_8 FILLER_78_1967 ();
 sg13g2_decap_8 FILLER_78_1974 ();
 sg13g2_decap_8 FILLER_78_1981 ();
 sg13g2_decap_8 FILLER_78_1988 ();
 sg13g2_decap_8 FILLER_78_1995 ();
 sg13g2_decap_8 FILLER_78_2002 ();
 sg13g2_decap_8 FILLER_78_2009 ();
 sg13g2_decap_8 FILLER_78_2016 ();
 sg13g2_decap_8 FILLER_78_2023 ();
 sg13g2_decap_8 FILLER_78_2030 ();
 sg13g2_decap_8 FILLER_78_2037 ();
 sg13g2_decap_8 FILLER_78_2044 ();
 sg13g2_decap_8 FILLER_78_2051 ();
 sg13g2_decap_8 FILLER_78_2058 ();
 sg13g2_decap_8 FILLER_78_2065 ();
 sg13g2_decap_8 FILLER_78_2072 ();
 sg13g2_decap_8 FILLER_78_2079 ();
 sg13g2_decap_8 FILLER_78_2086 ();
 sg13g2_decap_8 FILLER_78_2093 ();
 sg13g2_decap_8 FILLER_78_2100 ();
 sg13g2_decap_8 FILLER_78_2107 ();
 sg13g2_decap_8 FILLER_78_2114 ();
 sg13g2_decap_8 FILLER_78_2121 ();
 sg13g2_decap_8 FILLER_78_2128 ();
 sg13g2_decap_8 FILLER_78_2135 ();
 sg13g2_decap_8 FILLER_78_2142 ();
 sg13g2_decap_8 FILLER_78_2149 ();
 sg13g2_decap_8 FILLER_78_2156 ();
 sg13g2_decap_8 FILLER_78_2163 ();
 sg13g2_decap_8 FILLER_78_2170 ();
 sg13g2_decap_8 FILLER_78_2177 ();
 sg13g2_decap_8 FILLER_78_2184 ();
 sg13g2_decap_8 FILLER_78_2191 ();
 sg13g2_decap_8 FILLER_78_2198 ();
 sg13g2_decap_8 FILLER_78_2205 ();
 sg13g2_decap_8 FILLER_78_2212 ();
 sg13g2_decap_8 FILLER_78_2219 ();
 sg13g2_decap_8 FILLER_78_2226 ();
 sg13g2_decap_8 FILLER_78_2233 ();
 sg13g2_decap_8 FILLER_78_2240 ();
 sg13g2_decap_8 FILLER_78_2247 ();
 sg13g2_decap_8 FILLER_78_2254 ();
 sg13g2_decap_8 FILLER_78_2261 ();
 sg13g2_decap_8 FILLER_78_2268 ();
 sg13g2_decap_8 FILLER_78_2275 ();
 sg13g2_decap_8 FILLER_78_2282 ();
 sg13g2_decap_8 FILLER_78_2289 ();
 sg13g2_decap_8 FILLER_78_2296 ();
 sg13g2_decap_8 FILLER_78_2303 ();
 sg13g2_decap_8 FILLER_78_2310 ();
 sg13g2_decap_8 FILLER_78_2317 ();
 sg13g2_decap_8 FILLER_78_2324 ();
 sg13g2_decap_8 FILLER_78_2331 ();
 sg13g2_decap_8 FILLER_78_2338 ();
 sg13g2_decap_8 FILLER_78_2345 ();
 sg13g2_decap_8 FILLER_78_2352 ();
 sg13g2_decap_8 FILLER_78_2359 ();
 sg13g2_decap_8 FILLER_78_2366 ();
 sg13g2_decap_8 FILLER_78_2373 ();
 sg13g2_decap_8 FILLER_78_2380 ();
 sg13g2_decap_8 FILLER_78_2387 ();
 sg13g2_decap_8 FILLER_78_2394 ();
 sg13g2_decap_8 FILLER_78_2401 ();
 sg13g2_decap_8 FILLER_78_2408 ();
 sg13g2_decap_8 FILLER_78_2415 ();
 sg13g2_decap_8 FILLER_78_2422 ();
 sg13g2_decap_8 FILLER_78_2429 ();
 sg13g2_decap_8 FILLER_78_2436 ();
 sg13g2_decap_8 FILLER_78_2443 ();
 sg13g2_decap_8 FILLER_78_2450 ();
 sg13g2_decap_8 FILLER_78_2457 ();
 sg13g2_decap_8 FILLER_78_2464 ();
 sg13g2_decap_8 FILLER_78_2471 ();
 sg13g2_decap_8 FILLER_78_2478 ();
 sg13g2_decap_8 FILLER_78_2485 ();
 sg13g2_decap_8 FILLER_78_2492 ();
 sg13g2_decap_8 FILLER_78_2499 ();
 sg13g2_decap_8 FILLER_78_2506 ();
 sg13g2_decap_8 FILLER_78_2513 ();
 sg13g2_decap_8 FILLER_78_2520 ();
 sg13g2_decap_8 FILLER_78_2527 ();
 sg13g2_decap_8 FILLER_78_2534 ();
 sg13g2_decap_8 FILLER_78_2541 ();
 sg13g2_decap_8 FILLER_78_2548 ();
 sg13g2_decap_8 FILLER_78_2555 ();
 sg13g2_decap_8 FILLER_78_2562 ();
 sg13g2_decap_8 FILLER_78_2569 ();
 sg13g2_decap_8 FILLER_78_2576 ();
 sg13g2_decap_8 FILLER_78_2583 ();
 sg13g2_decap_8 FILLER_78_2590 ();
 sg13g2_decap_8 FILLER_78_2597 ();
 sg13g2_decap_8 FILLER_78_2604 ();
 sg13g2_decap_8 FILLER_78_2611 ();
 sg13g2_decap_8 FILLER_78_2618 ();
 sg13g2_decap_8 FILLER_78_2625 ();
 sg13g2_decap_8 FILLER_78_2632 ();
 sg13g2_decap_8 FILLER_78_2639 ();
 sg13g2_decap_8 FILLER_78_2646 ();
 sg13g2_decap_8 FILLER_78_2653 ();
 sg13g2_decap_8 FILLER_78_2660 ();
 sg13g2_decap_8 FILLER_78_2667 ();
 sg13g2_decap_8 FILLER_78_2674 ();
 sg13g2_decap_8 FILLER_78_2681 ();
 sg13g2_decap_8 FILLER_78_2688 ();
 sg13g2_decap_8 FILLER_78_2695 ();
 sg13g2_decap_8 FILLER_78_2702 ();
 sg13g2_decap_8 FILLER_78_2709 ();
 sg13g2_decap_8 FILLER_78_2716 ();
 sg13g2_decap_8 FILLER_78_2723 ();
 sg13g2_decap_8 FILLER_78_2730 ();
 sg13g2_decap_8 FILLER_78_2737 ();
 sg13g2_decap_8 FILLER_78_2744 ();
 sg13g2_decap_8 FILLER_78_2751 ();
 sg13g2_decap_8 FILLER_78_2758 ();
 sg13g2_decap_8 FILLER_78_2765 ();
 sg13g2_decap_8 FILLER_78_2772 ();
 sg13g2_decap_8 FILLER_78_2779 ();
 sg13g2_decap_8 FILLER_78_2786 ();
 sg13g2_decap_8 FILLER_78_2793 ();
 sg13g2_decap_8 FILLER_78_2800 ();
 sg13g2_decap_8 FILLER_78_2807 ();
 sg13g2_decap_8 FILLER_78_2814 ();
 sg13g2_decap_8 FILLER_78_2821 ();
 sg13g2_decap_8 FILLER_78_2828 ();
 sg13g2_decap_8 FILLER_78_2835 ();
 sg13g2_decap_8 FILLER_78_2842 ();
 sg13g2_decap_8 FILLER_78_2849 ();
 sg13g2_decap_8 FILLER_78_2856 ();
 sg13g2_decap_8 FILLER_78_2863 ();
 sg13g2_decap_8 FILLER_78_2870 ();
 sg13g2_decap_8 FILLER_78_2877 ();
 sg13g2_decap_8 FILLER_78_2884 ();
 sg13g2_decap_8 FILLER_78_2891 ();
 sg13g2_decap_8 FILLER_78_2898 ();
 sg13g2_decap_8 FILLER_78_2905 ();
 sg13g2_decap_8 FILLER_78_2912 ();
 sg13g2_decap_8 FILLER_78_2919 ();
 sg13g2_decap_8 FILLER_78_2926 ();
 sg13g2_decap_8 FILLER_78_2933 ();
 sg13g2_decap_8 FILLER_78_2940 ();
 sg13g2_decap_8 FILLER_78_2947 ();
 sg13g2_decap_8 FILLER_78_2954 ();
 sg13g2_decap_8 FILLER_78_2961 ();
 sg13g2_decap_8 FILLER_78_2968 ();
 sg13g2_decap_8 FILLER_78_2975 ();
 sg13g2_decap_8 FILLER_78_2982 ();
 sg13g2_decap_8 FILLER_78_2989 ();
 sg13g2_decap_8 FILLER_78_2996 ();
 sg13g2_decap_8 FILLER_78_3003 ();
 sg13g2_decap_8 FILLER_78_3010 ();
 sg13g2_decap_8 FILLER_78_3017 ();
 sg13g2_decap_8 FILLER_78_3024 ();
 sg13g2_decap_8 FILLER_78_3031 ();
 sg13g2_decap_8 FILLER_78_3038 ();
 sg13g2_decap_8 FILLER_78_3045 ();
 sg13g2_decap_8 FILLER_78_3052 ();
 sg13g2_decap_8 FILLER_78_3059 ();
 sg13g2_decap_8 FILLER_78_3066 ();
 sg13g2_decap_8 FILLER_78_3073 ();
 sg13g2_decap_8 FILLER_78_3080 ();
 sg13g2_decap_8 FILLER_78_3087 ();
 sg13g2_decap_8 FILLER_78_3094 ();
 sg13g2_decap_8 FILLER_78_3101 ();
 sg13g2_decap_8 FILLER_78_3108 ();
 sg13g2_decap_8 FILLER_78_3115 ();
 sg13g2_decap_8 FILLER_78_3122 ();
 sg13g2_decap_8 FILLER_78_3129 ();
 sg13g2_decap_8 FILLER_78_3136 ();
 sg13g2_decap_8 FILLER_78_3143 ();
 sg13g2_decap_8 FILLER_78_3150 ();
 sg13g2_decap_8 FILLER_78_3157 ();
 sg13g2_decap_8 FILLER_78_3164 ();
 sg13g2_decap_8 FILLER_78_3171 ();
 sg13g2_decap_8 FILLER_78_3178 ();
 sg13g2_decap_8 FILLER_78_3185 ();
 sg13g2_decap_8 FILLER_78_3192 ();
 sg13g2_decap_8 FILLER_78_3199 ();
 sg13g2_decap_8 FILLER_78_3206 ();
 sg13g2_decap_8 FILLER_78_3213 ();
 sg13g2_decap_8 FILLER_78_3220 ();
 sg13g2_decap_8 FILLER_78_3227 ();
 sg13g2_decap_8 FILLER_78_3234 ();
 sg13g2_decap_8 FILLER_78_3241 ();
 sg13g2_decap_8 FILLER_78_3248 ();
 sg13g2_decap_8 FILLER_78_3255 ();
 sg13g2_decap_8 FILLER_78_3262 ();
 sg13g2_decap_8 FILLER_78_3269 ();
 sg13g2_decap_8 FILLER_78_3276 ();
 sg13g2_decap_8 FILLER_78_3283 ();
 sg13g2_decap_8 FILLER_78_3290 ();
 sg13g2_decap_8 FILLER_78_3297 ();
 sg13g2_decap_8 FILLER_78_3304 ();
 sg13g2_decap_8 FILLER_78_3311 ();
 sg13g2_decap_8 FILLER_78_3318 ();
 sg13g2_decap_8 FILLER_78_3325 ();
 sg13g2_decap_8 FILLER_78_3332 ();
 sg13g2_decap_8 FILLER_78_3339 ();
 sg13g2_decap_8 FILLER_78_3346 ();
 sg13g2_decap_8 FILLER_78_3353 ();
 sg13g2_decap_8 FILLER_78_3360 ();
 sg13g2_decap_8 FILLER_78_3367 ();
 sg13g2_decap_8 FILLER_78_3374 ();
 sg13g2_decap_8 FILLER_78_3381 ();
 sg13g2_decap_8 FILLER_78_3388 ();
 sg13g2_decap_8 FILLER_78_3395 ();
 sg13g2_decap_8 FILLER_78_3402 ();
 sg13g2_decap_8 FILLER_78_3409 ();
 sg13g2_decap_8 FILLER_78_3416 ();
 sg13g2_decap_8 FILLER_78_3423 ();
 sg13g2_decap_8 FILLER_78_3430 ();
 sg13g2_decap_8 FILLER_78_3437 ();
 sg13g2_decap_8 FILLER_78_3444 ();
 sg13g2_decap_8 FILLER_78_3451 ();
 sg13g2_decap_8 FILLER_78_3458 ();
 sg13g2_decap_8 FILLER_78_3465 ();
 sg13g2_decap_8 FILLER_78_3472 ();
 sg13g2_decap_8 FILLER_78_3479 ();
 sg13g2_decap_8 FILLER_78_3486 ();
 sg13g2_decap_8 FILLER_78_3493 ();
 sg13g2_decap_8 FILLER_78_3500 ();
 sg13g2_decap_8 FILLER_78_3507 ();
 sg13g2_decap_8 FILLER_78_3514 ();
 sg13g2_decap_8 FILLER_78_3521 ();
 sg13g2_decap_8 FILLER_78_3528 ();
 sg13g2_decap_8 FILLER_78_3535 ();
 sg13g2_decap_8 FILLER_78_3542 ();
 sg13g2_decap_8 FILLER_78_3549 ();
 sg13g2_decap_8 FILLER_78_3556 ();
 sg13g2_decap_8 FILLER_78_3563 ();
 sg13g2_decap_8 FILLER_78_3570 ();
 sg13g2_fill_2 FILLER_78_3577 ();
 sg13g2_fill_1 FILLER_78_3579 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_168 ();
 sg13g2_decap_8 FILLER_79_175 ();
 sg13g2_decap_8 FILLER_79_182 ();
 sg13g2_decap_8 FILLER_79_189 ();
 sg13g2_decap_8 FILLER_79_196 ();
 sg13g2_decap_8 FILLER_79_203 ();
 sg13g2_decap_8 FILLER_79_210 ();
 sg13g2_decap_8 FILLER_79_217 ();
 sg13g2_decap_8 FILLER_79_224 ();
 sg13g2_decap_8 FILLER_79_231 ();
 sg13g2_decap_8 FILLER_79_238 ();
 sg13g2_decap_8 FILLER_79_245 ();
 sg13g2_decap_8 FILLER_79_252 ();
 sg13g2_decap_8 FILLER_79_259 ();
 sg13g2_decap_8 FILLER_79_266 ();
 sg13g2_decap_8 FILLER_79_273 ();
 sg13g2_decap_8 FILLER_79_280 ();
 sg13g2_decap_8 FILLER_79_287 ();
 sg13g2_decap_8 FILLER_79_294 ();
 sg13g2_decap_8 FILLER_79_301 ();
 sg13g2_decap_8 FILLER_79_308 ();
 sg13g2_decap_8 FILLER_79_315 ();
 sg13g2_decap_8 FILLER_79_322 ();
 sg13g2_decap_8 FILLER_79_329 ();
 sg13g2_decap_8 FILLER_79_336 ();
 sg13g2_decap_8 FILLER_79_343 ();
 sg13g2_decap_8 FILLER_79_350 ();
 sg13g2_decap_8 FILLER_79_357 ();
 sg13g2_decap_8 FILLER_79_364 ();
 sg13g2_decap_8 FILLER_79_371 ();
 sg13g2_decap_8 FILLER_79_378 ();
 sg13g2_decap_8 FILLER_79_385 ();
 sg13g2_decap_8 FILLER_79_392 ();
 sg13g2_decap_8 FILLER_79_399 ();
 sg13g2_decap_8 FILLER_79_406 ();
 sg13g2_decap_8 FILLER_79_413 ();
 sg13g2_decap_8 FILLER_79_420 ();
 sg13g2_decap_8 FILLER_79_427 ();
 sg13g2_decap_8 FILLER_79_434 ();
 sg13g2_decap_8 FILLER_79_441 ();
 sg13g2_decap_8 FILLER_79_448 ();
 sg13g2_decap_8 FILLER_79_455 ();
 sg13g2_decap_8 FILLER_79_462 ();
 sg13g2_decap_8 FILLER_79_469 ();
 sg13g2_decap_8 FILLER_79_476 ();
 sg13g2_decap_8 FILLER_79_483 ();
 sg13g2_decap_8 FILLER_79_490 ();
 sg13g2_decap_8 FILLER_79_497 ();
 sg13g2_decap_8 FILLER_79_504 ();
 sg13g2_decap_8 FILLER_79_511 ();
 sg13g2_decap_8 FILLER_79_518 ();
 sg13g2_decap_8 FILLER_79_525 ();
 sg13g2_decap_8 FILLER_79_532 ();
 sg13g2_decap_8 FILLER_79_539 ();
 sg13g2_decap_8 FILLER_79_546 ();
 sg13g2_decap_8 FILLER_79_553 ();
 sg13g2_decap_8 FILLER_79_560 ();
 sg13g2_decap_8 FILLER_79_567 ();
 sg13g2_decap_8 FILLER_79_574 ();
 sg13g2_decap_8 FILLER_79_581 ();
 sg13g2_decap_8 FILLER_79_588 ();
 sg13g2_decap_8 FILLER_79_595 ();
 sg13g2_decap_8 FILLER_79_602 ();
 sg13g2_decap_8 FILLER_79_609 ();
 sg13g2_decap_8 FILLER_79_616 ();
 sg13g2_decap_8 FILLER_79_623 ();
 sg13g2_decap_8 FILLER_79_630 ();
 sg13g2_decap_8 FILLER_79_637 ();
 sg13g2_decap_8 FILLER_79_644 ();
 sg13g2_decap_8 FILLER_79_651 ();
 sg13g2_decap_8 FILLER_79_658 ();
 sg13g2_decap_8 FILLER_79_665 ();
 sg13g2_decap_8 FILLER_79_672 ();
 sg13g2_decap_8 FILLER_79_679 ();
 sg13g2_decap_8 FILLER_79_686 ();
 sg13g2_decap_8 FILLER_79_693 ();
 sg13g2_decap_8 FILLER_79_700 ();
 sg13g2_decap_8 FILLER_79_707 ();
 sg13g2_decap_8 FILLER_79_714 ();
 sg13g2_decap_8 FILLER_79_721 ();
 sg13g2_decap_8 FILLER_79_728 ();
 sg13g2_decap_8 FILLER_79_735 ();
 sg13g2_decap_8 FILLER_79_742 ();
 sg13g2_decap_8 FILLER_79_749 ();
 sg13g2_decap_8 FILLER_79_756 ();
 sg13g2_decap_8 FILLER_79_763 ();
 sg13g2_decap_8 FILLER_79_770 ();
 sg13g2_decap_8 FILLER_79_777 ();
 sg13g2_decap_8 FILLER_79_784 ();
 sg13g2_decap_8 FILLER_79_791 ();
 sg13g2_decap_8 FILLER_79_798 ();
 sg13g2_decap_8 FILLER_79_805 ();
 sg13g2_decap_8 FILLER_79_812 ();
 sg13g2_decap_8 FILLER_79_819 ();
 sg13g2_decap_8 FILLER_79_826 ();
 sg13g2_decap_8 FILLER_79_833 ();
 sg13g2_decap_8 FILLER_79_840 ();
 sg13g2_decap_8 FILLER_79_847 ();
 sg13g2_decap_8 FILLER_79_854 ();
 sg13g2_decap_8 FILLER_79_861 ();
 sg13g2_decap_8 FILLER_79_868 ();
 sg13g2_decap_8 FILLER_79_875 ();
 sg13g2_decap_8 FILLER_79_882 ();
 sg13g2_decap_8 FILLER_79_889 ();
 sg13g2_decap_8 FILLER_79_896 ();
 sg13g2_decap_8 FILLER_79_903 ();
 sg13g2_decap_8 FILLER_79_910 ();
 sg13g2_decap_8 FILLER_79_917 ();
 sg13g2_decap_8 FILLER_79_924 ();
 sg13g2_decap_8 FILLER_79_931 ();
 sg13g2_decap_8 FILLER_79_938 ();
 sg13g2_decap_8 FILLER_79_945 ();
 sg13g2_decap_8 FILLER_79_952 ();
 sg13g2_decap_8 FILLER_79_959 ();
 sg13g2_decap_8 FILLER_79_966 ();
 sg13g2_decap_8 FILLER_79_973 ();
 sg13g2_decap_8 FILLER_79_980 ();
 sg13g2_decap_8 FILLER_79_987 ();
 sg13g2_decap_8 FILLER_79_994 ();
 sg13g2_decap_8 FILLER_79_1001 ();
 sg13g2_decap_8 FILLER_79_1008 ();
 sg13g2_decap_8 FILLER_79_1015 ();
 sg13g2_decap_8 FILLER_79_1022 ();
 sg13g2_decap_8 FILLER_79_1029 ();
 sg13g2_decap_8 FILLER_79_1036 ();
 sg13g2_decap_8 FILLER_79_1043 ();
 sg13g2_decap_8 FILLER_79_1050 ();
 sg13g2_decap_8 FILLER_79_1057 ();
 sg13g2_decap_8 FILLER_79_1064 ();
 sg13g2_decap_8 FILLER_79_1071 ();
 sg13g2_decap_8 FILLER_79_1078 ();
 sg13g2_decap_8 FILLER_79_1085 ();
 sg13g2_decap_8 FILLER_79_1092 ();
 sg13g2_decap_8 FILLER_79_1099 ();
 sg13g2_decap_8 FILLER_79_1106 ();
 sg13g2_decap_8 FILLER_79_1113 ();
 sg13g2_decap_8 FILLER_79_1120 ();
 sg13g2_decap_8 FILLER_79_1127 ();
 sg13g2_decap_8 FILLER_79_1134 ();
 sg13g2_decap_8 FILLER_79_1141 ();
 sg13g2_decap_8 FILLER_79_1148 ();
 sg13g2_decap_8 FILLER_79_1155 ();
 sg13g2_decap_8 FILLER_79_1162 ();
 sg13g2_decap_8 FILLER_79_1169 ();
 sg13g2_decap_8 FILLER_79_1176 ();
 sg13g2_decap_8 FILLER_79_1183 ();
 sg13g2_decap_8 FILLER_79_1190 ();
 sg13g2_decap_8 FILLER_79_1197 ();
 sg13g2_decap_8 FILLER_79_1204 ();
 sg13g2_decap_8 FILLER_79_1211 ();
 sg13g2_decap_8 FILLER_79_1218 ();
 sg13g2_decap_8 FILLER_79_1225 ();
 sg13g2_decap_8 FILLER_79_1232 ();
 sg13g2_decap_8 FILLER_79_1239 ();
 sg13g2_decap_8 FILLER_79_1246 ();
 sg13g2_decap_8 FILLER_79_1253 ();
 sg13g2_decap_8 FILLER_79_1260 ();
 sg13g2_decap_8 FILLER_79_1267 ();
 sg13g2_decap_8 FILLER_79_1274 ();
 sg13g2_decap_8 FILLER_79_1281 ();
 sg13g2_decap_8 FILLER_79_1288 ();
 sg13g2_decap_8 FILLER_79_1295 ();
 sg13g2_decap_8 FILLER_79_1302 ();
 sg13g2_decap_8 FILLER_79_1309 ();
 sg13g2_decap_8 FILLER_79_1316 ();
 sg13g2_decap_8 FILLER_79_1323 ();
 sg13g2_decap_8 FILLER_79_1330 ();
 sg13g2_decap_8 FILLER_79_1337 ();
 sg13g2_decap_8 FILLER_79_1344 ();
 sg13g2_decap_8 FILLER_79_1351 ();
 sg13g2_decap_8 FILLER_79_1358 ();
 sg13g2_decap_8 FILLER_79_1365 ();
 sg13g2_decap_8 FILLER_79_1372 ();
 sg13g2_decap_8 FILLER_79_1379 ();
 sg13g2_decap_8 FILLER_79_1386 ();
 sg13g2_decap_8 FILLER_79_1393 ();
 sg13g2_decap_8 FILLER_79_1400 ();
 sg13g2_decap_8 FILLER_79_1407 ();
 sg13g2_decap_8 FILLER_79_1414 ();
 sg13g2_decap_8 FILLER_79_1421 ();
 sg13g2_decap_8 FILLER_79_1428 ();
 sg13g2_decap_8 FILLER_79_1435 ();
 sg13g2_decap_8 FILLER_79_1442 ();
 sg13g2_decap_8 FILLER_79_1449 ();
 sg13g2_decap_8 FILLER_79_1456 ();
 sg13g2_decap_8 FILLER_79_1463 ();
 sg13g2_decap_8 FILLER_79_1470 ();
 sg13g2_decap_8 FILLER_79_1477 ();
 sg13g2_decap_8 FILLER_79_1484 ();
 sg13g2_decap_8 FILLER_79_1491 ();
 sg13g2_decap_8 FILLER_79_1498 ();
 sg13g2_decap_8 FILLER_79_1505 ();
 sg13g2_decap_8 FILLER_79_1512 ();
 sg13g2_decap_8 FILLER_79_1519 ();
 sg13g2_decap_8 FILLER_79_1526 ();
 sg13g2_decap_8 FILLER_79_1533 ();
 sg13g2_decap_8 FILLER_79_1540 ();
 sg13g2_decap_8 FILLER_79_1547 ();
 sg13g2_decap_8 FILLER_79_1554 ();
 sg13g2_decap_8 FILLER_79_1561 ();
 sg13g2_decap_8 FILLER_79_1568 ();
 sg13g2_decap_8 FILLER_79_1575 ();
 sg13g2_decap_8 FILLER_79_1582 ();
 sg13g2_decap_8 FILLER_79_1589 ();
 sg13g2_decap_8 FILLER_79_1596 ();
 sg13g2_decap_8 FILLER_79_1603 ();
 sg13g2_decap_8 FILLER_79_1610 ();
 sg13g2_decap_8 FILLER_79_1617 ();
 sg13g2_decap_8 FILLER_79_1624 ();
 sg13g2_decap_8 FILLER_79_1631 ();
 sg13g2_decap_8 FILLER_79_1638 ();
 sg13g2_decap_8 FILLER_79_1645 ();
 sg13g2_decap_8 FILLER_79_1652 ();
 sg13g2_decap_8 FILLER_79_1659 ();
 sg13g2_decap_8 FILLER_79_1666 ();
 sg13g2_decap_8 FILLER_79_1673 ();
 sg13g2_decap_8 FILLER_79_1680 ();
 sg13g2_decap_8 FILLER_79_1687 ();
 sg13g2_decap_8 FILLER_79_1694 ();
 sg13g2_decap_8 FILLER_79_1701 ();
 sg13g2_decap_8 FILLER_79_1708 ();
 sg13g2_decap_8 FILLER_79_1715 ();
 sg13g2_decap_8 FILLER_79_1722 ();
 sg13g2_decap_8 FILLER_79_1729 ();
 sg13g2_decap_8 FILLER_79_1736 ();
 sg13g2_decap_8 FILLER_79_1743 ();
 sg13g2_decap_8 FILLER_79_1750 ();
 sg13g2_decap_8 FILLER_79_1757 ();
 sg13g2_decap_8 FILLER_79_1764 ();
 sg13g2_decap_8 FILLER_79_1771 ();
 sg13g2_decap_8 FILLER_79_1778 ();
 sg13g2_decap_8 FILLER_79_1785 ();
 sg13g2_decap_8 FILLER_79_1792 ();
 sg13g2_decap_8 FILLER_79_1799 ();
 sg13g2_decap_8 FILLER_79_1806 ();
 sg13g2_decap_8 FILLER_79_1813 ();
 sg13g2_decap_8 FILLER_79_1820 ();
 sg13g2_decap_8 FILLER_79_1827 ();
 sg13g2_decap_8 FILLER_79_1834 ();
 sg13g2_decap_8 FILLER_79_1841 ();
 sg13g2_decap_8 FILLER_79_1848 ();
 sg13g2_decap_8 FILLER_79_1855 ();
 sg13g2_decap_8 FILLER_79_1862 ();
 sg13g2_decap_8 FILLER_79_1869 ();
 sg13g2_decap_8 FILLER_79_1876 ();
 sg13g2_decap_8 FILLER_79_1883 ();
 sg13g2_decap_8 FILLER_79_1890 ();
 sg13g2_decap_8 FILLER_79_1897 ();
 sg13g2_decap_8 FILLER_79_1904 ();
 sg13g2_decap_8 FILLER_79_1911 ();
 sg13g2_decap_8 FILLER_79_1918 ();
 sg13g2_decap_8 FILLER_79_1925 ();
 sg13g2_decap_8 FILLER_79_1932 ();
 sg13g2_decap_8 FILLER_79_1939 ();
 sg13g2_decap_8 FILLER_79_1946 ();
 sg13g2_decap_8 FILLER_79_1953 ();
 sg13g2_decap_8 FILLER_79_1960 ();
 sg13g2_decap_8 FILLER_79_1967 ();
 sg13g2_decap_8 FILLER_79_1974 ();
 sg13g2_decap_8 FILLER_79_1981 ();
 sg13g2_decap_8 FILLER_79_1988 ();
 sg13g2_decap_8 FILLER_79_1995 ();
 sg13g2_decap_8 FILLER_79_2002 ();
 sg13g2_decap_8 FILLER_79_2009 ();
 sg13g2_decap_8 FILLER_79_2016 ();
 sg13g2_decap_8 FILLER_79_2023 ();
 sg13g2_decap_8 FILLER_79_2030 ();
 sg13g2_decap_8 FILLER_79_2037 ();
 sg13g2_decap_8 FILLER_79_2044 ();
 sg13g2_decap_8 FILLER_79_2051 ();
 sg13g2_decap_8 FILLER_79_2058 ();
 sg13g2_decap_8 FILLER_79_2065 ();
 sg13g2_decap_8 FILLER_79_2072 ();
 sg13g2_decap_8 FILLER_79_2079 ();
 sg13g2_decap_8 FILLER_79_2086 ();
 sg13g2_decap_8 FILLER_79_2093 ();
 sg13g2_decap_8 FILLER_79_2100 ();
 sg13g2_decap_8 FILLER_79_2107 ();
 sg13g2_decap_8 FILLER_79_2114 ();
 sg13g2_decap_8 FILLER_79_2121 ();
 sg13g2_decap_8 FILLER_79_2128 ();
 sg13g2_decap_8 FILLER_79_2135 ();
 sg13g2_decap_8 FILLER_79_2142 ();
 sg13g2_decap_8 FILLER_79_2149 ();
 sg13g2_decap_8 FILLER_79_2156 ();
 sg13g2_decap_8 FILLER_79_2163 ();
 sg13g2_decap_8 FILLER_79_2170 ();
 sg13g2_decap_8 FILLER_79_2177 ();
 sg13g2_decap_8 FILLER_79_2184 ();
 sg13g2_decap_8 FILLER_79_2191 ();
 sg13g2_decap_8 FILLER_79_2198 ();
 sg13g2_decap_8 FILLER_79_2205 ();
 sg13g2_decap_8 FILLER_79_2212 ();
 sg13g2_decap_8 FILLER_79_2219 ();
 sg13g2_decap_8 FILLER_79_2226 ();
 sg13g2_decap_8 FILLER_79_2233 ();
 sg13g2_decap_8 FILLER_79_2240 ();
 sg13g2_decap_8 FILLER_79_2247 ();
 sg13g2_decap_8 FILLER_79_2254 ();
 sg13g2_decap_8 FILLER_79_2261 ();
 sg13g2_decap_8 FILLER_79_2268 ();
 sg13g2_decap_8 FILLER_79_2275 ();
 sg13g2_decap_8 FILLER_79_2282 ();
 sg13g2_decap_8 FILLER_79_2289 ();
 sg13g2_decap_8 FILLER_79_2296 ();
 sg13g2_decap_8 FILLER_79_2303 ();
 sg13g2_decap_8 FILLER_79_2310 ();
 sg13g2_decap_8 FILLER_79_2317 ();
 sg13g2_decap_8 FILLER_79_2324 ();
 sg13g2_decap_8 FILLER_79_2331 ();
 sg13g2_decap_8 FILLER_79_2338 ();
 sg13g2_decap_8 FILLER_79_2345 ();
 sg13g2_decap_8 FILLER_79_2352 ();
 sg13g2_decap_8 FILLER_79_2359 ();
 sg13g2_decap_8 FILLER_79_2366 ();
 sg13g2_decap_8 FILLER_79_2373 ();
 sg13g2_decap_8 FILLER_79_2380 ();
 sg13g2_decap_8 FILLER_79_2387 ();
 sg13g2_decap_8 FILLER_79_2394 ();
 sg13g2_decap_8 FILLER_79_2401 ();
 sg13g2_decap_8 FILLER_79_2408 ();
 sg13g2_decap_8 FILLER_79_2415 ();
 sg13g2_decap_8 FILLER_79_2422 ();
 sg13g2_decap_8 FILLER_79_2429 ();
 sg13g2_decap_8 FILLER_79_2436 ();
 sg13g2_decap_8 FILLER_79_2443 ();
 sg13g2_decap_8 FILLER_79_2450 ();
 sg13g2_decap_8 FILLER_79_2457 ();
 sg13g2_decap_8 FILLER_79_2464 ();
 sg13g2_decap_8 FILLER_79_2471 ();
 sg13g2_decap_8 FILLER_79_2478 ();
 sg13g2_decap_8 FILLER_79_2485 ();
 sg13g2_decap_8 FILLER_79_2492 ();
 sg13g2_decap_8 FILLER_79_2499 ();
 sg13g2_decap_8 FILLER_79_2506 ();
 sg13g2_decap_8 FILLER_79_2513 ();
 sg13g2_decap_8 FILLER_79_2520 ();
 sg13g2_decap_8 FILLER_79_2527 ();
 sg13g2_decap_8 FILLER_79_2534 ();
 sg13g2_decap_8 FILLER_79_2541 ();
 sg13g2_decap_8 FILLER_79_2548 ();
 sg13g2_decap_8 FILLER_79_2555 ();
 sg13g2_decap_8 FILLER_79_2562 ();
 sg13g2_decap_8 FILLER_79_2569 ();
 sg13g2_decap_8 FILLER_79_2576 ();
 sg13g2_decap_8 FILLER_79_2583 ();
 sg13g2_decap_8 FILLER_79_2590 ();
 sg13g2_decap_8 FILLER_79_2597 ();
 sg13g2_decap_8 FILLER_79_2604 ();
 sg13g2_decap_8 FILLER_79_2611 ();
 sg13g2_decap_8 FILLER_79_2618 ();
 sg13g2_decap_8 FILLER_79_2625 ();
 sg13g2_decap_8 FILLER_79_2632 ();
 sg13g2_decap_8 FILLER_79_2639 ();
 sg13g2_decap_8 FILLER_79_2646 ();
 sg13g2_decap_8 FILLER_79_2653 ();
 sg13g2_decap_8 FILLER_79_2660 ();
 sg13g2_decap_8 FILLER_79_2667 ();
 sg13g2_decap_8 FILLER_79_2674 ();
 sg13g2_decap_8 FILLER_79_2681 ();
 sg13g2_decap_8 FILLER_79_2688 ();
 sg13g2_decap_8 FILLER_79_2695 ();
 sg13g2_decap_8 FILLER_79_2702 ();
 sg13g2_decap_8 FILLER_79_2709 ();
 sg13g2_decap_8 FILLER_79_2716 ();
 sg13g2_decap_8 FILLER_79_2723 ();
 sg13g2_decap_8 FILLER_79_2730 ();
 sg13g2_decap_8 FILLER_79_2737 ();
 sg13g2_decap_8 FILLER_79_2744 ();
 sg13g2_decap_8 FILLER_79_2751 ();
 sg13g2_decap_8 FILLER_79_2758 ();
 sg13g2_decap_8 FILLER_79_2765 ();
 sg13g2_decap_8 FILLER_79_2772 ();
 sg13g2_decap_8 FILLER_79_2779 ();
 sg13g2_decap_8 FILLER_79_2786 ();
 sg13g2_decap_8 FILLER_79_2793 ();
 sg13g2_decap_8 FILLER_79_2800 ();
 sg13g2_decap_8 FILLER_79_2807 ();
 sg13g2_decap_8 FILLER_79_2814 ();
 sg13g2_decap_8 FILLER_79_2821 ();
 sg13g2_decap_8 FILLER_79_2828 ();
 sg13g2_decap_8 FILLER_79_2835 ();
 sg13g2_decap_8 FILLER_79_2842 ();
 sg13g2_decap_8 FILLER_79_2849 ();
 sg13g2_decap_8 FILLER_79_2856 ();
 sg13g2_decap_8 FILLER_79_2863 ();
 sg13g2_decap_8 FILLER_79_2870 ();
 sg13g2_decap_8 FILLER_79_2877 ();
 sg13g2_decap_8 FILLER_79_2884 ();
 sg13g2_decap_8 FILLER_79_2891 ();
 sg13g2_decap_8 FILLER_79_2898 ();
 sg13g2_decap_8 FILLER_79_2905 ();
 sg13g2_decap_8 FILLER_79_2912 ();
 sg13g2_decap_8 FILLER_79_2919 ();
 sg13g2_decap_8 FILLER_79_2926 ();
 sg13g2_decap_8 FILLER_79_2933 ();
 sg13g2_decap_8 FILLER_79_2940 ();
 sg13g2_decap_8 FILLER_79_2947 ();
 sg13g2_decap_8 FILLER_79_2954 ();
 sg13g2_decap_8 FILLER_79_2961 ();
 sg13g2_decap_8 FILLER_79_2968 ();
 sg13g2_decap_8 FILLER_79_2975 ();
 sg13g2_decap_8 FILLER_79_2982 ();
 sg13g2_decap_8 FILLER_79_2989 ();
 sg13g2_decap_8 FILLER_79_2996 ();
 sg13g2_decap_8 FILLER_79_3003 ();
 sg13g2_decap_8 FILLER_79_3010 ();
 sg13g2_decap_8 FILLER_79_3017 ();
 sg13g2_decap_8 FILLER_79_3024 ();
 sg13g2_decap_8 FILLER_79_3031 ();
 sg13g2_decap_8 FILLER_79_3038 ();
 sg13g2_decap_8 FILLER_79_3045 ();
 sg13g2_decap_8 FILLER_79_3052 ();
 sg13g2_decap_8 FILLER_79_3059 ();
 sg13g2_decap_8 FILLER_79_3066 ();
 sg13g2_decap_8 FILLER_79_3073 ();
 sg13g2_decap_8 FILLER_79_3080 ();
 sg13g2_decap_8 FILLER_79_3087 ();
 sg13g2_decap_8 FILLER_79_3094 ();
 sg13g2_decap_8 FILLER_79_3101 ();
 sg13g2_decap_8 FILLER_79_3108 ();
 sg13g2_decap_8 FILLER_79_3115 ();
 sg13g2_decap_8 FILLER_79_3122 ();
 sg13g2_decap_8 FILLER_79_3129 ();
 sg13g2_decap_8 FILLER_79_3136 ();
 sg13g2_decap_8 FILLER_79_3143 ();
 sg13g2_decap_8 FILLER_79_3150 ();
 sg13g2_decap_8 FILLER_79_3157 ();
 sg13g2_decap_8 FILLER_79_3164 ();
 sg13g2_decap_8 FILLER_79_3171 ();
 sg13g2_decap_8 FILLER_79_3178 ();
 sg13g2_decap_8 FILLER_79_3185 ();
 sg13g2_decap_8 FILLER_79_3192 ();
 sg13g2_decap_8 FILLER_79_3199 ();
 sg13g2_decap_8 FILLER_79_3206 ();
 sg13g2_decap_8 FILLER_79_3213 ();
 sg13g2_decap_8 FILLER_79_3220 ();
 sg13g2_decap_8 FILLER_79_3227 ();
 sg13g2_decap_8 FILLER_79_3234 ();
 sg13g2_decap_8 FILLER_79_3241 ();
 sg13g2_decap_8 FILLER_79_3248 ();
 sg13g2_decap_8 FILLER_79_3255 ();
 sg13g2_decap_8 FILLER_79_3262 ();
 sg13g2_decap_8 FILLER_79_3269 ();
 sg13g2_decap_8 FILLER_79_3276 ();
 sg13g2_decap_8 FILLER_79_3283 ();
 sg13g2_decap_8 FILLER_79_3290 ();
 sg13g2_decap_8 FILLER_79_3297 ();
 sg13g2_decap_8 FILLER_79_3304 ();
 sg13g2_decap_8 FILLER_79_3311 ();
 sg13g2_decap_8 FILLER_79_3318 ();
 sg13g2_decap_8 FILLER_79_3325 ();
 sg13g2_decap_8 FILLER_79_3332 ();
 sg13g2_decap_8 FILLER_79_3339 ();
 sg13g2_decap_8 FILLER_79_3346 ();
 sg13g2_decap_8 FILLER_79_3353 ();
 sg13g2_decap_8 FILLER_79_3360 ();
 sg13g2_decap_8 FILLER_79_3367 ();
 sg13g2_decap_8 FILLER_79_3374 ();
 sg13g2_decap_8 FILLER_79_3381 ();
 sg13g2_decap_8 FILLER_79_3388 ();
 sg13g2_decap_8 FILLER_79_3395 ();
 sg13g2_decap_8 FILLER_79_3402 ();
 sg13g2_decap_8 FILLER_79_3409 ();
 sg13g2_decap_8 FILLER_79_3416 ();
 sg13g2_decap_8 FILLER_79_3423 ();
 sg13g2_decap_8 FILLER_79_3430 ();
 sg13g2_decap_8 FILLER_79_3437 ();
 sg13g2_decap_8 FILLER_79_3444 ();
 sg13g2_decap_8 FILLER_79_3451 ();
 sg13g2_decap_8 FILLER_79_3458 ();
 sg13g2_decap_8 FILLER_79_3465 ();
 sg13g2_decap_8 FILLER_79_3472 ();
 sg13g2_decap_8 FILLER_79_3479 ();
 sg13g2_decap_8 FILLER_79_3486 ();
 sg13g2_decap_8 FILLER_79_3493 ();
 sg13g2_decap_8 FILLER_79_3500 ();
 sg13g2_decap_8 FILLER_79_3507 ();
 sg13g2_decap_8 FILLER_79_3514 ();
 sg13g2_decap_8 FILLER_79_3521 ();
 sg13g2_decap_8 FILLER_79_3528 ();
 sg13g2_decap_8 FILLER_79_3535 ();
 sg13g2_decap_8 FILLER_79_3542 ();
 sg13g2_decap_8 FILLER_79_3549 ();
 sg13g2_decap_8 FILLER_79_3556 ();
 sg13g2_decap_8 FILLER_79_3563 ();
 sg13g2_decap_8 FILLER_79_3570 ();
 sg13g2_fill_2 FILLER_79_3577 ();
 sg13g2_fill_1 FILLER_79_3579 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_201 ();
 sg13g2_decap_8 FILLER_80_208 ();
 sg13g2_decap_8 FILLER_80_215 ();
 sg13g2_decap_8 FILLER_80_222 ();
 sg13g2_decap_8 FILLER_80_229 ();
 sg13g2_decap_8 FILLER_80_236 ();
 sg13g2_decap_8 FILLER_80_243 ();
 sg13g2_decap_8 FILLER_80_250 ();
 sg13g2_decap_8 FILLER_80_257 ();
 sg13g2_decap_8 FILLER_80_264 ();
 sg13g2_decap_8 FILLER_80_271 ();
 sg13g2_decap_8 FILLER_80_278 ();
 sg13g2_decap_8 FILLER_80_285 ();
 sg13g2_decap_8 FILLER_80_292 ();
 sg13g2_decap_8 FILLER_80_299 ();
 sg13g2_decap_8 FILLER_80_306 ();
 sg13g2_decap_8 FILLER_80_313 ();
 sg13g2_decap_8 FILLER_80_320 ();
 sg13g2_decap_8 FILLER_80_327 ();
 sg13g2_decap_8 FILLER_80_334 ();
 sg13g2_decap_8 FILLER_80_341 ();
 sg13g2_decap_8 FILLER_80_348 ();
 sg13g2_decap_4 FILLER_80_355 ();
 sg13g2_fill_1 FILLER_80_359 ();
 sg13g2_fill_2 FILLER_80_365 ();
 sg13g2_fill_1 FILLER_80_367 ();
 sg13g2_decap_4 FILLER_80_372 ();
 sg13g2_decap_8 FILLER_80_381 ();
 sg13g2_decap_8 FILLER_80_388 ();
 sg13g2_decap_8 FILLER_80_395 ();
 sg13g2_decap_8 FILLER_80_402 ();
 sg13g2_decap_8 FILLER_80_409 ();
 sg13g2_decap_8 FILLER_80_416 ();
 sg13g2_decap_8 FILLER_80_423 ();
 sg13g2_decap_8 FILLER_80_430 ();
 sg13g2_decap_8 FILLER_80_437 ();
 sg13g2_decap_8 FILLER_80_444 ();
 sg13g2_decap_8 FILLER_80_451 ();
 sg13g2_decap_8 FILLER_80_458 ();
 sg13g2_decap_8 FILLER_80_465 ();
 sg13g2_decap_8 FILLER_80_472 ();
 sg13g2_decap_8 FILLER_80_479 ();
 sg13g2_decap_8 FILLER_80_486 ();
 sg13g2_decap_8 FILLER_80_493 ();
 sg13g2_decap_8 FILLER_80_500 ();
 sg13g2_decap_8 FILLER_80_507 ();
 sg13g2_decap_8 FILLER_80_514 ();
 sg13g2_decap_8 FILLER_80_521 ();
 sg13g2_decap_8 FILLER_80_528 ();
 sg13g2_decap_8 FILLER_80_535 ();
 sg13g2_decap_8 FILLER_80_542 ();
 sg13g2_decap_8 FILLER_80_549 ();
 sg13g2_decap_8 FILLER_80_556 ();
 sg13g2_decap_8 FILLER_80_563 ();
 sg13g2_decap_8 FILLER_80_570 ();
 sg13g2_decap_8 FILLER_80_577 ();
 sg13g2_decap_8 FILLER_80_584 ();
 sg13g2_decap_8 FILLER_80_591 ();
 sg13g2_decap_8 FILLER_80_598 ();
 sg13g2_decap_8 FILLER_80_605 ();
 sg13g2_decap_8 FILLER_80_612 ();
 sg13g2_decap_8 FILLER_80_619 ();
 sg13g2_decap_8 FILLER_80_626 ();
 sg13g2_decap_8 FILLER_80_633 ();
 sg13g2_decap_8 FILLER_80_640 ();
 sg13g2_decap_8 FILLER_80_647 ();
 sg13g2_decap_8 FILLER_80_654 ();
 sg13g2_decap_8 FILLER_80_661 ();
 sg13g2_decap_8 FILLER_80_668 ();
 sg13g2_decap_8 FILLER_80_675 ();
 sg13g2_decap_8 FILLER_80_682 ();
 sg13g2_decap_8 FILLER_80_689 ();
 sg13g2_decap_8 FILLER_80_696 ();
 sg13g2_decap_8 FILLER_80_703 ();
 sg13g2_decap_8 FILLER_80_710 ();
 sg13g2_decap_8 FILLER_80_717 ();
 sg13g2_decap_8 FILLER_80_724 ();
 sg13g2_decap_8 FILLER_80_731 ();
 sg13g2_decap_8 FILLER_80_738 ();
 sg13g2_decap_8 FILLER_80_745 ();
 sg13g2_decap_8 FILLER_80_752 ();
 sg13g2_decap_8 FILLER_80_759 ();
 sg13g2_decap_8 FILLER_80_766 ();
 sg13g2_decap_8 FILLER_80_773 ();
 sg13g2_decap_8 FILLER_80_780 ();
 sg13g2_decap_8 FILLER_80_787 ();
 sg13g2_decap_8 FILLER_80_794 ();
 sg13g2_decap_8 FILLER_80_801 ();
 sg13g2_decap_8 FILLER_80_808 ();
 sg13g2_decap_8 FILLER_80_815 ();
 sg13g2_decap_8 FILLER_80_822 ();
 sg13g2_decap_8 FILLER_80_829 ();
 sg13g2_decap_8 FILLER_80_836 ();
 sg13g2_decap_8 FILLER_80_843 ();
 sg13g2_decap_8 FILLER_80_850 ();
 sg13g2_decap_8 FILLER_80_857 ();
 sg13g2_decap_8 FILLER_80_864 ();
 sg13g2_decap_8 FILLER_80_871 ();
 sg13g2_decap_8 FILLER_80_878 ();
 sg13g2_decap_8 FILLER_80_885 ();
 sg13g2_decap_8 FILLER_80_892 ();
 sg13g2_decap_8 FILLER_80_899 ();
 sg13g2_decap_8 FILLER_80_906 ();
 sg13g2_decap_8 FILLER_80_913 ();
 sg13g2_decap_8 FILLER_80_920 ();
 sg13g2_decap_8 FILLER_80_927 ();
 sg13g2_decap_8 FILLER_80_934 ();
 sg13g2_decap_8 FILLER_80_941 ();
 sg13g2_decap_8 FILLER_80_948 ();
 sg13g2_decap_8 FILLER_80_955 ();
 sg13g2_decap_8 FILLER_80_962 ();
 sg13g2_decap_8 FILLER_80_969 ();
 sg13g2_decap_8 FILLER_80_976 ();
 sg13g2_decap_8 FILLER_80_983 ();
 sg13g2_decap_8 FILLER_80_990 ();
 sg13g2_decap_8 FILLER_80_997 ();
 sg13g2_decap_8 FILLER_80_1004 ();
 sg13g2_decap_8 FILLER_80_1011 ();
 sg13g2_decap_8 FILLER_80_1018 ();
 sg13g2_decap_8 FILLER_80_1025 ();
 sg13g2_decap_8 FILLER_80_1032 ();
 sg13g2_decap_8 FILLER_80_1039 ();
 sg13g2_decap_8 FILLER_80_1046 ();
 sg13g2_decap_8 FILLER_80_1053 ();
 sg13g2_decap_8 FILLER_80_1060 ();
 sg13g2_decap_8 FILLER_80_1067 ();
 sg13g2_decap_8 FILLER_80_1074 ();
 sg13g2_decap_8 FILLER_80_1081 ();
 sg13g2_decap_8 FILLER_80_1088 ();
 sg13g2_decap_8 FILLER_80_1095 ();
 sg13g2_decap_8 FILLER_80_1102 ();
 sg13g2_decap_8 FILLER_80_1109 ();
 sg13g2_decap_8 FILLER_80_1116 ();
 sg13g2_decap_8 FILLER_80_1123 ();
 sg13g2_decap_8 FILLER_80_1130 ();
 sg13g2_decap_8 FILLER_80_1137 ();
 sg13g2_decap_8 FILLER_80_1144 ();
 sg13g2_decap_8 FILLER_80_1151 ();
 sg13g2_decap_8 FILLER_80_1158 ();
 sg13g2_decap_8 FILLER_80_1165 ();
 sg13g2_decap_8 FILLER_80_1172 ();
 sg13g2_decap_8 FILLER_80_1179 ();
 sg13g2_decap_8 FILLER_80_1186 ();
 sg13g2_decap_8 FILLER_80_1193 ();
 sg13g2_decap_8 FILLER_80_1200 ();
 sg13g2_decap_8 FILLER_80_1207 ();
 sg13g2_decap_8 FILLER_80_1214 ();
 sg13g2_decap_8 FILLER_80_1221 ();
 sg13g2_decap_8 FILLER_80_1228 ();
 sg13g2_decap_8 FILLER_80_1235 ();
 sg13g2_decap_8 FILLER_80_1242 ();
 sg13g2_decap_8 FILLER_80_1249 ();
 sg13g2_decap_8 FILLER_80_1256 ();
 sg13g2_decap_8 FILLER_80_1263 ();
 sg13g2_decap_8 FILLER_80_1270 ();
 sg13g2_decap_8 FILLER_80_1277 ();
 sg13g2_decap_8 FILLER_80_1284 ();
 sg13g2_decap_8 FILLER_80_1291 ();
 sg13g2_decap_8 FILLER_80_1298 ();
 sg13g2_decap_8 FILLER_80_1305 ();
 sg13g2_decap_8 FILLER_80_1312 ();
 sg13g2_decap_8 FILLER_80_1319 ();
 sg13g2_decap_8 FILLER_80_1326 ();
 sg13g2_decap_8 FILLER_80_1333 ();
 sg13g2_decap_8 FILLER_80_1340 ();
 sg13g2_decap_8 FILLER_80_1347 ();
 sg13g2_decap_8 FILLER_80_1354 ();
 sg13g2_decap_8 FILLER_80_1361 ();
 sg13g2_decap_8 FILLER_80_1368 ();
 sg13g2_decap_8 FILLER_80_1375 ();
 sg13g2_decap_8 FILLER_80_1382 ();
 sg13g2_decap_8 FILLER_80_1389 ();
 sg13g2_decap_8 FILLER_80_1396 ();
 sg13g2_decap_8 FILLER_80_1403 ();
 sg13g2_decap_8 FILLER_80_1410 ();
 sg13g2_decap_8 FILLER_80_1417 ();
 sg13g2_decap_8 FILLER_80_1424 ();
 sg13g2_decap_8 FILLER_80_1431 ();
 sg13g2_decap_8 FILLER_80_1438 ();
 sg13g2_decap_8 FILLER_80_1445 ();
 sg13g2_decap_8 FILLER_80_1452 ();
 sg13g2_decap_8 FILLER_80_1459 ();
 sg13g2_decap_8 FILLER_80_1466 ();
 sg13g2_decap_8 FILLER_80_1473 ();
 sg13g2_decap_8 FILLER_80_1480 ();
 sg13g2_decap_8 FILLER_80_1487 ();
 sg13g2_decap_8 FILLER_80_1494 ();
 sg13g2_decap_8 FILLER_80_1501 ();
 sg13g2_decap_8 FILLER_80_1508 ();
 sg13g2_decap_8 FILLER_80_1515 ();
 sg13g2_decap_8 FILLER_80_1522 ();
 sg13g2_decap_8 FILLER_80_1529 ();
 sg13g2_decap_8 FILLER_80_1536 ();
 sg13g2_decap_8 FILLER_80_1543 ();
 sg13g2_decap_8 FILLER_80_1550 ();
 sg13g2_decap_8 FILLER_80_1557 ();
 sg13g2_decap_8 FILLER_80_1564 ();
 sg13g2_decap_8 FILLER_80_1571 ();
 sg13g2_decap_8 FILLER_80_1578 ();
 sg13g2_decap_8 FILLER_80_1585 ();
 sg13g2_decap_8 FILLER_80_1592 ();
 sg13g2_decap_8 FILLER_80_1599 ();
 sg13g2_decap_8 FILLER_80_1606 ();
 sg13g2_decap_8 FILLER_80_1613 ();
 sg13g2_decap_8 FILLER_80_1620 ();
 sg13g2_decap_8 FILLER_80_1627 ();
 sg13g2_decap_8 FILLER_80_1634 ();
 sg13g2_decap_8 FILLER_80_1641 ();
 sg13g2_decap_8 FILLER_80_1648 ();
 sg13g2_decap_8 FILLER_80_1655 ();
 sg13g2_decap_8 FILLER_80_1662 ();
 sg13g2_decap_8 FILLER_80_1669 ();
 sg13g2_decap_8 FILLER_80_1676 ();
 sg13g2_decap_8 FILLER_80_1683 ();
 sg13g2_decap_8 FILLER_80_1690 ();
 sg13g2_decap_8 FILLER_80_1697 ();
 sg13g2_decap_8 FILLER_80_1704 ();
 sg13g2_decap_8 FILLER_80_1711 ();
 sg13g2_decap_8 FILLER_80_1718 ();
 sg13g2_decap_8 FILLER_80_1725 ();
 sg13g2_decap_8 FILLER_80_1732 ();
 sg13g2_decap_8 FILLER_80_1739 ();
 sg13g2_decap_8 FILLER_80_1746 ();
 sg13g2_decap_8 FILLER_80_1753 ();
 sg13g2_decap_8 FILLER_80_1760 ();
 sg13g2_decap_8 FILLER_80_1767 ();
 sg13g2_decap_8 FILLER_80_1774 ();
 sg13g2_decap_8 FILLER_80_1781 ();
 sg13g2_decap_8 FILLER_80_1788 ();
 sg13g2_decap_8 FILLER_80_1795 ();
 sg13g2_decap_8 FILLER_80_1802 ();
 sg13g2_decap_8 FILLER_80_1809 ();
 sg13g2_decap_8 FILLER_80_1816 ();
 sg13g2_decap_8 FILLER_80_1823 ();
 sg13g2_decap_8 FILLER_80_1830 ();
 sg13g2_decap_8 FILLER_80_1837 ();
 sg13g2_decap_8 FILLER_80_1844 ();
 sg13g2_decap_8 FILLER_80_1851 ();
 sg13g2_decap_8 FILLER_80_1858 ();
 sg13g2_decap_8 FILLER_80_1865 ();
 sg13g2_decap_8 FILLER_80_1872 ();
 sg13g2_decap_8 FILLER_80_1879 ();
 sg13g2_decap_8 FILLER_80_1886 ();
 sg13g2_decap_8 FILLER_80_1893 ();
 sg13g2_decap_8 FILLER_80_1900 ();
 sg13g2_decap_8 FILLER_80_1907 ();
 sg13g2_decap_8 FILLER_80_1914 ();
 sg13g2_decap_8 FILLER_80_1921 ();
 sg13g2_decap_8 FILLER_80_1928 ();
 sg13g2_decap_8 FILLER_80_1935 ();
 sg13g2_decap_8 FILLER_80_1942 ();
 sg13g2_decap_8 FILLER_80_1949 ();
 sg13g2_decap_8 FILLER_80_1956 ();
 sg13g2_decap_8 FILLER_80_1963 ();
 sg13g2_decap_8 FILLER_80_1970 ();
 sg13g2_decap_8 FILLER_80_1977 ();
 sg13g2_decap_8 FILLER_80_1984 ();
 sg13g2_decap_8 FILLER_80_1991 ();
 sg13g2_decap_8 FILLER_80_1998 ();
 sg13g2_decap_8 FILLER_80_2005 ();
 sg13g2_decap_8 FILLER_80_2012 ();
 sg13g2_decap_8 FILLER_80_2019 ();
 sg13g2_decap_8 FILLER_80_2026 ();
 sg13g2_decap_8 FILLER_80_2033 ();
 sg13g2_decap_8 FILLER_80_2040 ();
 sg13g2_decap_8 FILLER_80_2047 ();
 sg13g2_decap_8 FILLER_80_2054 ();
 sg13g2_decap_8 FILLER_80_2061 ();
 sg13g2_decap_8 FILLER_80_2068 ();
 sg13g2_decap_8 FILLER_80_2075 ();
 sg13g2_decap_8 FILLER_80_2082 ();
 sg13g2_decap_8 FILLER_80_2089 ();
 sg13g2_decap_8 FILLER_80_2096 ();
 sg13g2_decap_8 FILLER_80_2103 ();
 sg13g2_decap_8 FILLER_80_2110 ();
 sg13g2_decap_8 FILLER_80_2117 ();
 sg13g2_decap_8 FILLER_80_2124 ();
 sg13g2_decap_8 FILLER_80_2131 ();
 sg13g2_decap_8 FILLER_80_2138 ();
 sg13g2_decap_8 FILLER_80_2145 ();
 sg13g2_decap_8 FILLER_80_2152 ();
 sg13g2_decap_8 FILLER_80_2159 ();
 sg13g2_decap_8 FILLER_80_2166 ();
 sg13g2_decap_8 FILLER_80_2173 ();
 sg13g2_decap_8 FILLER_80_2180 ();
 sg13g2_decap_8 FILLER_80_2187 ();
 sg13g2_decap_8 FILLER_80_2194 ();
 sg13g2_decap_8 FILLER_80_2201 ();
 sg13g2_decap_8 FILLER_80_2208 ();
 sg13g2_decap_8 FILLER_80_2215 ();
 sg13g2_decap_8 FILLER_80_2222 ();
 sg13g2_decap_8 FILLER_80_2229 ();
 sg13g2_decap_8 FILLER_80_2236 ();
 sg13g2_decap_8 FILLER_80_2243 ();
 sg13g2_decap_8 FILLER_80_2250 ();
 sg13g2_decap_8 FILLER_80_2257 ();
 sg13g2_decap_8 FILLER_80_2264 ();
 sg13g2_decap_8 FILLER_80_2271 ();
 sg13g2_decap_8 FILLER_80_2278 ();
 sg13g2_decap_8 FILLER_80_2285 ();
 sg13g2_decap_8 FILLER_80_2292 ();
 sg13g2_decap_8 FILLER_80_2299 ();
 sg13g2_decap_8 FILLER_80_2306 ();
 sg13g2_decap_8 FILLER_80_2313 ();
 sg13g2_decap_8 FILLER_80_2320 ();
 sg13g2_decap_8 FILLER_80_2327 ();
 sg13g2_decap_8 FILLER_80_2334 ();
 sg13g2_decap_8 FILLER_80_2341 ();
 sg13g2_decap_8 FILLER_80_2348 ();
 sg13g2_decap_8 FILLER_80_2355 ();
 sg13g2_decap_8 FILLER_80_2362 ();
 sg13g2_decap_8 FILLER_80_2369 ();
 sg13g2_decap_8 FILLER_80_2376 ();
 sg13g2_decap_8 FILLER_80_2383 ();
 sg13g2_decap_8 FILLER_80_2390 ();
 sg13g2_decap_8 FILLER_80_2397 ();
 sg13g2_decap_8 FILLER_80_2404 ();
 sg13g2_decap_8 FILLER_80_2411 ();
 sg13g2_decap_8 FILLER_80_2418 ();
 sg13g2_decap_8 FILLER_80_2425 ();
 sg13g2_decap_8 FILLER_80_2432 ();
 sg13g2_decap_8 FILLER_80_2439 ();
 sg13g2_decap_8 FILLER_80_2446 ();
 sg13g2_decap_8 FILLER_80_2453 ();
 sg13g2_decap_8 FILLER_80_2460 ();
 sg13g2_decap_8 FILLER_80_2467 ();
 sg13g2_decap_8 FILLER_80_2474 ();
 sg13g2_decap_8 FILLER_80_2481 ();
 sg13g2_decap_8 FILLER_80_2488 ();
 sg13g2_decap_8 FILLER_80_2495 ();
 sg13g2_decap_8 FILLER_80_2502 ();
 sg13g2_decap_8 FILLER_80_2509 ();
 sg13g2_decap_8 FILLER_80_2516 ();
 sg13g2_decap_8 FILLER_80_2523 ();
 sg13g2_decap_8 FILLER_80_2530 ();
 sg13g2_decap_8 FILLER_80_2537 ();
 sg13g2_decap_8 FILLER_80_2544 ();
 sg13g2_decap_8 FILLER_80_2551 ();
 sg13g2_decap_8 FILLER_80_2558 ();
 sg13g2_decap_8 FILLER_80_2565 ();
 sg13g2_decap_8 FILLER_80_2572 ();
 sg13g2_decap_8 FILLER_80_2579 ();
 sg13g2_decap_8 FILLER_80_2586 ();
 sg13g2_decap_8 FILLER_80_2593 ();
 sg13g2_decap_8 FILLER_80_2600 ();
 sg13g2_decap_8 FILLER_80_2607 ();
 sg13g2_decap_8 FILLER_80_2614 ();
 sg13g2_decap_8 FILLER_80_2621 ();
 sg13g2_decap_8 FILLER_80_2628 ();
 sg13g2_decap_8 FILLER_80_2635 ();
 sg13g2_decap_8 FILLER_80_2642 ();
 sg13g2_decap_8 FILLER_80_2649 ();
 sg13g2_decap_8 FILLER_80_2656 ();
 sg13g2_decap_8 FILLER_80_2663 ();
 sg13g2_decap_8 FILLER_80_2670 ();
 sg13g2_decap_8 FILLER_80_2677 ();
 sg13g2_decap_8 FILLER_80_2684 ();
 sg13g2_decap_8 FILLER_80_2691 ();
 sg13g2_decap_8 FILLER_80_2698 ();
 sg13g2_decap_8 FILLER_80_2705 ();
 sg13g2_decap_8 FILLER_80_2712 ();
 sg13g2_decap_8 FILLER_80_2719 ();
 sg13g2_decap_8 FILLER_80_2726 ();
 sg13g2_decap_8 FILLER_80_2733 ();
 sg13g2_decap_8 FILLER_80_2740 ();
 sg13g2_decap_8 FILLER_80_2747 ();
 sg13g2_decap_8 FILLER_80_2754 ();
 sg13g2_decap_8 FILLER_80_2761 ();
 sg13g2_decap_8 FILLER_80_2768 ();
 sg13g2_decap_8 FILLER_80_2775 ();
 sg13g2_decap_8 FILLER_80_2782 ();
 sg13g2_decap_8 FILLER_80_2789 ();
 sg13g2_decap_8 FILLER_80_2796 ();
 sg13g2_decap_8 FILLER_80_2803 ();
 sg13g2_decap_8 FILLER_80_2810 ();
 sg13g2_decap_8 FILLER_80_2817 ();
 sg13g2_decap_8 FILLER_80_2824 ();
 sg13g2_decap_8 FILLER_80_2831 ();
 sg13g2_decap_8 FILLER_80_2838 ();
 sg13g2_decap_8 FILLER_80_2845 ();
 sg13g2_decap_8 FILLER_80_2852 ();
 sg13g2_decap_8 FILLER_80_2859 ();
 sg13g2_decap_8 FILLER_80_2866 ();
 sg13g2_decap_8 FILLER_80_2873 ();
 sg13g2_decap_8 FILLER_80_2880 ();
 sg13g2_decap_8 FILLER_80_2887 ();
 sg13g2_decap_8 FILLER_80_2894 ();
 sg13g2_decap_8 FILLER_80_2901 ();
 sg13g2_decap_8 FILLER_80_2908 ();
 sg13g2_decap_8 FILLER_80_2915 ();
 sg13g2_decap_8 FILLER_80_2922 ();
 sg13g2_decap_8 FILLER_80_2929 ();
 sg13g2_decap_8 FILLER_80_2936 ();
 sg13g2_decap_8 FILLER_80_2943 ();
 sg13g2_decap_8 FILLER_80_2950 ();
 sg13g2_decap_8 FILLER_80_2957 ();
 sg13g2_decap_8 FILLER_80_2964 ();
 sg13g2_decap_8 FILLER_80_2971 ();
 sg13g2_decap_8 FILLER_80_2978 ();
 sg13g2_decap_8 FILLER_80_2985 ();
 sg13g2_decap_8 FILLER_80_2992 ();
 sg13g2_decap_8 FILLER_80_2999 ();
 sg13g2_decap_8 FILLER_80_3006 ();
 sg13g2_decap_8 FILLER_80_3013 ();
 sg13g2_decap_8 FILLER_80_3020 ();
 sg13g2_decap_8 FILLER_80_3027 ();
 sg13g2_decap_8 FILLER_80_3034 ();
 sg13g2_decap_8 FILLER_80_3041 ();
 sg13g2_decap_8 FILLER_80_3048 ();
 sg13g2_decap_8 FILLER_80_3055 ();
 sg13g2_decap_8 FILLER_80_3062 ();
 sg13g2_decap_8 FILLER_80_3069 ();
 sg13g2_decap_8 FILLER_80_3076 ();
 sg13g2_decap_8 FILLER_80_3083 ();
 sg13g2_decap_8 FILLER_80_3090 ();
 sg13g2_decap_8 FILLER_80_3097 ();
 sg13g2_decap_8 FILLER_80_3104 ();
 sg13g2_decap_8 FILLER_80_3111 ();
 sg13g2_decap_8 FILLER_80_3118 ();
 sg13g2_decap_8 FILLER_80_3125 ();
 sg13g2_decap_8 FILLER_80_3132 ();
 sg13g2_decap_8 FILLER_80_3139 ();
 sg13g2_decap_8 FILLER_80_3146 ();
 sg13g2_decap_8 FILLER_80_3153 ();
 sg13g2_decap_8 FILLER_80_3160 ();
 sg13g2_decap_8 FILLER_80_3167 ();
 sg13g2_decap_8 FILLER_80_3174 ();
 sg13g2_decap_8 FILLER_80_3181 ();
 sg13g2_decap_8 FILLER_80_3188 ();
 sg13g2_decap_8 FILLER_80_3195 ();
 sg13g2_decap_8 FILLER_80_3202 ();
 sg13g2_decap_8 FILLER_80_3209 ();
 sg13g2_decap_8 FILLER_80_3216 ();
 sg13g2_decap_8 FILLER_80_3223 ();
 sg13g2_decap_8 FILLER_80_3230 ();
 sg13g2_decap_8 FILLER_80_3237 ();
 sg13g2_decap_8 FILLER_80_3244 ();
 sg13g2_decap_8 FILLER_80_3251 ();
 sg13g2_decap_8 FILLER_80_3258 ();
 sg13g2_decap_8 FILLER_80_3265 ();
 sg13g2_decap_8 FILLER_80_3272 ();
 sg13g2_decap_8 FILLER_80_3279 ();
 sg13g2_decap_8 FILLER_80_3286 ();
 sg13g2_decap_8 FILLER_80_3293 ();
 sg13g2_decap_8 FILLER_80_3300 ();
 sg13g2_decap_8 FILLER_80_3307 ();
 sg13g2_decap_8 FILLER_80_3314 ();
 sg13g2_decap_8 FILLER_80_3321 ();
 sg13g2_decap_8 FILLER_80_3328 ();
 sg13g2_decap_8 FILLER_80_3335 ();
 sg13g2_decap_8 FILLER_80_3342 ();
 sg13g2_decap_8 FILLER_80_3349 ();
 sg13g2_decap_8 FILLER_80_3356 ();
 sg13g2_decap_8 FILLER_80_3363 ();
 sg13g2_decap_8 FILLER_80_3370 ();
 sg13g2_decap_8 FILLER_80_3377 ();
 sg13g2_decap_8 FILLER_80_3384 ();
 sg13g2_decap_8 FILLER_80_3391 ();
 sg13g2_decap_8 FILLER_80_3398 ();
 sg13g2_decap_8 FILLER_80_3405 ();
 sg13g2_decap_8 FILLER_80_3412 ();
 sg13g2_decap_8 FILLER_80_3419 ();
 sg13g2_decap_8 FILLER_80_3426 ();
 sg13g2_decap_8 FILLER_80_3433 ();
 sg13g2_decap_8 FILLER_80_3440 ();
 sg13g2_decap_8 FILLER_80_3447 ();
 sg13g2_decap_8 FILLER_80_3454 ();
 sg13g2_decap_8 FILLER_80_3461 ();
 sg13g2_decap_8 FILLER_80_3468 ();
 sg13g2_decap_8 FILLER_80_3475 ();
 sg13g2_decap_8 FILLER_80_3482 ();
 sg13g2_decap_8 FILLER_80_3489 ();
 sg13g2_decap_8 FILLER_80_3496 ();
 sg13g2_decap_8 FILLER_80_3503 ();
 sg13g2_decap_8 FILLER_80_3510 ();
 sg13g2_decap_8 FILLER_80_3517 ();
 sg13g2_decap_8 FILLER_80_3524 ();
 sg13g2_decap_8 FILLER_80_3531 ();
 sg13g2_decap_8 FILLER_80_3538 ();
 sg13g2_decap_8 FILLER_80_3545 ();
 sg13g2_decap_8 FILLER_80_3552 ();
 sg13g2_decap_8 FILLER_80_3559 ();
 sg13g2_decap_8 FILLER_80_3566 ();
 sg13g2_decap_8 FILLER_80_3573 ();
 assign uio_oe[0] = net7;
 assign uio_oe[1] = net8;
 assign uio_oe[2] = net9;
 assign uio_oe[3] = net10;
 assign uio_oe[4] = net11;
 assign uio_oe[5] = net12;
 assign uio_oe[6] = net13;
 assign uio_oe[7] = net14;
 assign uio_out[0] = net15;
 assign uio_out[1] = net16;
 assign uio_out[2] = net17;
 assign uio_out[3] = net18;
 assign uio_out[4] = net19;
 assign uio_out[5] = net20;
 assign uio_out[6] = net21;
 assign uio_out[7] = net22;
endmodule
