module tt_um_ebeam_pixel_core (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire cfg_miso;
 wire \cfg_wr_addr_ff1[0] ;
 wire \cfg_wr_addr_ff1[1] ;
 wire \cfg_wr_addr_ff1[2] ;
 wire \cfg_wr_addr_ff2[0] ;
 wire \cfg_wr_addr_ff2[1] ;
 wire \cfg_wr_addr_ff2[2] ;
 wire \cfg_wr_data_ff1[0] ;
 wire \cfg_wr_data_ff1[1] ;
 wire \cfg_wr_data_ff1[2] ;
 wire \cfg_wr_data_ff1[3] ;
 wire \cfg_wr_data_ff1[4] ;
 wire \cfg_wr_data_ff1[5] ;
 wire \cfg_wr_data_ff1[6] ;
 wire \cfg_wr_data_ff1[7] ;
 wire \cfg_wr_data_ff2[0] ;
 wire \cfg_wr_data_ff2[1] ;
 wire \cfg_wr_data_ff2[2] ;
 wire \cfg_wr_data_ff2[3] ;
 wire \cfg_wr_data_ff2[4] ;
 wire \cfg_wr_data_ff2[5] ;
 wire \cfg_wr_data_ff2[6] ;
 wire \cfg_wr_data_ff2[7] ;
 wire cfg_wr_toggle_ff1;
 wire cfg_wr_toggle_ff2;
 wire cfg_wr_toggle_ff2_d;
 wire \mean_q[0] ;
 wire \mean_q[1] ;
 wire \mean_q[2] ;
 wire \mean_q[3] ;
 wire \mean_q[4] ;
 wire \mean_q[5] ;
 wire \mean_q[6] ;
 wire \mean_q[7] ;
 wire \pixel_q[0] ;
 wire \pixel_q[1] ;
 wire \pixel_q[2] ;
 wire \pixel_q[3] ;
 wire \pixel_q[4] ;
 wire \pixel_q[5] ;
 wire \pixel_q[6] ;
 wire \pixel_q[7] ;
 wire \prev_pixel[0] ;
 wire \prev_pixel[1] ;
 wire \prev_pixel[2] ;
 wire \prev_pixel[3] ;
 wire \prev_pixel[4] ;
 wire \prev_pixel[5] ;
 wire \prev_pixel[6] ;
 wire \prev_pixel[7] ;
 wire \reg_absdiff_rdback[0] ;
 wire \reg_absdiff_rdback[1] ;
 wire \reg_absdiff_rdback[2] ;
 wire \reg_absdiff_rdback[3] ;
 wire \reg_absdiff_rdback[4] ;
 wire \reg_absdiff_rdback[5] ;
 wire \reg_absdiff_rdback[6] ;
 wire \reg_absdiff_rdback[7] ;
 wire \reg_alpha_shift[2] ;
 wire \reg_contrast_thr[0] ;
 wire \reg_contrast_thr[1] ;
 wire \reg_contrast_thr[4] ;
 wire \reg_contrast_thr[5] ;
 wire \reg_contrast_thr[6] ;
 wire \reg_contrast_thr[7] ;
 wire \reg_edge_thr[0] ;
 wire \reg_edge_thr[1] ;
 wire \reg_edge_thr[4] ;
 wire \reg_edge_thr[5] ;
 wire \reg_edge_thr[6] ;
 wire \reg_edge_thr[7] ;
 wire \reg_mode[0] ;
 wire \reg_mode[1] ;
 wire \reg_mode[2] ;
 wire \reg_mode[3] ;
 wire \reg_mode[4] ;
 wire \reg_mode[5] ;
 wire \reg_mode[6] ;
 wire \reg_mode[7] ;
 wire \reg_status[4] ;
 wire \reg_status[5] ;
 wire \reg_status[6] ;
 wire \reg_status[7] ;
 wire \reg_thresh[0] ;
 wire \reg_thresh[1] ;
 wire \reg_thresh[2] ;
 wire \reg_thresh[3] ;
 wire \reg_thresh[4] ;
 wire \reg_thresh[5] ;
 wire \reg_thresh[6] ;
 wire \spi_bitcnt[0] ;
 wire \spi_bitcnt[1] ;
 wire \spi_bitcnt[2] ;
 wire \spi_bitcnt[3] ;
 wire \spi_cmd_addr[0] ;
 wire \spi_cmd_addr[1] ;
 wire \spi_cmd_addr[2] ;
 wire spi_cmd_wr;
 wire \spi_rd_bus_ff1[0] ;
 wire \spi_rd_bus_ff1[10] ;
 wire \spi_rd_bus_ff1[11] ;
 wire \spi_rd_bus_ff1[12] ;
 wire \spi_rd_bus_ff1[13] ;
 wire \spi_rd_bus_ff1[14] ;
 wire \spi_rd_bus_ff1[15] ;
 wire \spi_rd_bus_ff1[16] ;
 wire \spi_rd_bus_ff1[17] ;
 wire \spi_rd_bus_ff1[18] ;
 wire \spi_rd_bus_ff1[19] ;
 wire \spi_rd_bus_ff1[1] ;
 wire \spi_rd_bus_ff1[20] ;
 wire \spi_rd_bus_ff1[21] ;
 wire \spi_rd_bus_ff1[22] ;
 wire \spi_rd_bus_ff1[23] ;
 wire \spi_rd_bus_ff1[24] ;
 wire \spi_rd_bus_ff1[25] ;
 wire \spi_rd_bus_ff1[26] ;
 wire \spi_rd_bus_ff1[2] ;
 wire \spi_rd_bus_ff1[32] ;
 wire \spi_rd_bus_ff1[33] ;
 wire \spi_rd_bus_ff1[34] ;
 wire \spi_rd_bus_ff1[35] ;
 wire \spi_rd_bus_ff1[36] ;
 wire \spi_rd_bus_ff1[37] ;
 wire \spi_rd_bus_ff1[38] ;
 wire \spi_rd_bus_ff1[39] ;
 wire \spi_rd_bus_ff1[3] ;
 wire \spi_rd_bus_ff1[44] ;
 wire \spi_rd_bus_ff1[45] ;
 wire \spi_rd_bus_ff1[46] ;
 wire \spi_rd_bus_ff1[47] ;
 wire \spi_rd_bus_ff1[48] ;
 wire \spi_rd_bus_ff1[49] ;
 wire \spi_rd_bus_ff1[4] ;
 wire \spi_rd_bus_ff1[50] ;
 wire \spi_rd_bus_ff1[51] ;
 wire \spi_rd_bus_ff1[52] ;
 wire \spi_rd_bus_ff1[53] ;
 wire \spi_rd_bus_ff1[54] ;
 wire \spi_rd_bus_ff1[55] ;
 wire \spi_rd_bus_ff1[56] ;
 wire \spi_rd_bus_ff1[57] ;
 wire \spi_rd_bus_ff1[58] ;
 wire \spi_rd_bus_ff1[59] ;
 wire \spi_rd_bus_ff1[5] ;
 wire \spi_rd_bus_ff1[60] ;
 wire \spi_rd_bus_ff1[61] ;
 wire \spi_rd_bus_ff1[62] ;
 wire \spi_rd_bus_ff1[63] ;
 wire \spi_rd_bus_ff1[6] ;
 wire \spi_rd_bus_ff1[7] ;
 wire \spi_rd_bus_ff1[8] ;
 wire \spi_rd_bus_ff1[9] ;
 wire \spi_rd_bus_ff2[0] ;
 wire \spi_rd_bus_ff2[10] ;
 wire \spi_rd_bus_ff2[11] ;
 wire \spi_rd_bus_ff2[12] ;
 wire \spi_rd_bus_ff2[13] ;
 wire \spi_rd_bus_ff2[14] ;
 wire \spi_rd_bus_ff2[15] ;
 wire \spi_rd_bus_ff2[16] ;
 wire \spi_rd_bus_ff2[17] ;
 wire \spi_rd_bus_ff2[18] ;
 wire \spi_rd_bus_ff2[19] ;
 wire \spi_rd_bus_ff2[1] ;
 wire \spi_rd_bus_ff2[20] ;
 wire \spi_rd_bus_ff2[21] ;
 wire \spi_rd_bus_ff2[22] ;
 wire \spi_rd_bus_ff2[23] ;
 wire \spi_rd_bus_ff2[24] ;
 wire \spi_rd_bus_ff2[25] ;
 wire \spi_rd_bus_ff2[26] ;
 wire \spi_rd_bus_ff2[2] ;
 wire \spi_rd_bus_ff2[32] ;
 wire \spi_rd_bus_ff2[33] ;
 wire \spi_rd_bus_ff2[34] ;
 wire \spi_rd_bus_ff2[35] ;
 wire \spi_rd_bus_ff2[36] ;
 wire \spi_rd_bus_ff2[37] ;
 wire \spi_rd_bus_ff2[38] ;
 wire \spi_rd_bus_ff2[39] ;
 wire \spi_rd_bus_ff2[3] ;
 wire \spi_rd_bus_ff2[44] ;
 wire \spi_rd_bus_ff2[45] ;
 wire \spi_rd_bus_ff2[46] ;
 wire \spi_rd_bus_ff2[47] ;
 wire \spi_rd_bus_ff2[48] ;
 wire \spi_rd_bus_ff2[49] ;
 wire \spi_rd_bus_ff2[4] ;
 wire \spi_rd_bus_ff2[50] ;
 wire \spi_rd_bus_ff2[51] ;
 wire \spi_rd_bus_ff2[52] ;
 wire \spi_rd_bus_ff2[53] ;
 wire \spi_rd_bus_ff2[54] ;
 wire \spi_rd_bus_ff2[55] ;
 wire \spi_rd_bus_ff2[56] ;
 wire \spi_rd_bus_ff2[57] ;
 wire \spi_rd_bus_ff2[58] ;
 wire \spi_rd_bus_ff2[59] ;
 wire \spi_rd_bus_ff2[5] ;
 wire \spi_rd_bus_ff2[60] ;
 wire \spi_rd_bus_ff2[61] ;
 wire \spi_rd_bus_ff2[62] ;
 wire \spi_rd_bus_ff2[63] ;
 wire \spi_rd_bus_ff2[6] ;
 wire \spi_rd_bus_ff2[7] ;
 wire \spi_rd_bus_ff2[8] ;
 wire \spi_rd_bus_ff2[9] ;
 wire \spi_shift_in[0] ;
 wire \spi_shift_in[1] ;
 wire \spi_shift_in[2] ;
 wire \spi_shift_in[3] ;
 wire \spi_shift_in[4] ;
 wire \spi_shift_in[5] ;
 wire \spi_shift_in[6] ;
 wire \spi_shift_out[1] ;
 wire \spi_shift_out[2] ;
 wire \spi_shift_out[3] ;
 wire \spi_shift_out[4] ;
 wire \spi_shift_out[5] ;
 wire \spi_shift_out[6] ;
 wire \spi_shift_out[7] ;
 wire \spi_shift_out_load[0] ;
 wire \spi_shift_out_load[1] ;
 wire \spi_shift_out_load[2] ;
 wire \spi_shift_out_load[3] ;
 wire \spi_shift_out_load[4] ;
 wire \spi_shift_out_load[5] ;
 wire \spi_shift_out_load[6] ;
 wire \spi_shift_out_load[7] ;
 wire spi_shift_out_load_pending;
 wire \spi_wr_addr[0] ;
 wire \spi_wr_addr[1] ;
 wire \spi_wr_addr[2] ;
 wire \spi_wr_data[0] ;
 wire \spi_wr_data[1] ;
 wire \spi_wr_data[2] ;
 wire \spi_wr_data[3] ;
 wire \spi_wr_data[4] ;
 wire \spi_wr_data[5] ;
 wire \spi_wr_data[6] ;
 wire \spi_wr_data[7] ;
 wire spi_wr_toggle;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire clknet_0_clk;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;

 sg13g2_inv_2 _0858_ (.Y(_0367_),
    .A(net254));
 sg13g2_inv_2 _0859_ (.Y(_0368_),
    .A(net255));
 sg13g2_inv_1 _0860_ (.Y(_0369_),
    .A(_0019_));
 sg13g2_inv_2 _0861_ (.Y(_0030_),
    .A(net302));
 sg13g2_inv_1 _0862_ (.Y(_0370_),
    .A(\mean_q[0] ));
 sg13g2_inv_2 _0863_ (.Y(_0371_),
    .A(net379));
 sg13g2_inv_1 _0864_ (.Y(_0372_),
    .A(net204));
 sg13g2_inv_1 _0865_ (.Y(_0373_),
    .A(net216));
 sg13g2_inv_1 _0866_ (.Y(_0374_),
    .A(net394));
 sg13g2_inv_1 _0867_ (.Y(_0375_),
    .A(net375));
 sg13g2_inv_1 _0868_ (.Y(_0376_),
    .A(net208));
 sg13g2_inv_1 _0869_ (.Y(_0377_),
    .A(net381));
 sg13g2_inv_1 _0870_ (.Y(_0378_),
    .A(net399));
 sg13g2_inv_1 _0871_ (.Y(_0379_),
    .A(net220));
 sg13g2_inv_2 _0872_ (.Y(_0380_),
    .A(net397));
 sg13g2_inv_1 _0873_ (.Y(_0381_),
    .A(net234));
 sg13g2_inv_2 _0874_ (.Y(_0382_),
    .A(net403));
 sg13g2_inv_1 _0875_ (.Y(_0383_),
    .A(net214));
 sg13g2_inv_1 _0876_ (.Y(_0384_),
    .A(net395));
 sg13g2_inv_2 _0877_ (.Y(_0385_),
    .A(net163));
 sg13g2_inv_2 _0878_ (.Y(_0386_),
    .A(net179));
 sg13g2_inv_1 _0879_ (.Y(_0387_),
    .A(net385));
 sg13g2_inv_1 _0880_ (.Y(_0388_),
    .A(net398));
 sg13g2_inv_2 _0881_ (.Y(_0389_),
    .A(net380));
 sg13g2_inv_1 _0882_ (.Y(_0390_),
    .A(net400));
 sg13g2_inv_1 _0883_ (.Y(_0391_),
    .A(net401));
 sg13g2_inv_1 _0884_ (.Y(_0392_),
    .A(net391));
 sg13g2_inv_1 _0885_ (.Y(_0393_),
    .A(net202));
 sg13g2_inv_4 _0886_ (.A(net259),
    .Y(_0394_));
 sg13g2_inv_4 _0887_ (.A(\spi_shift_in[3] ),
    .Y(_0395_));
 sg13g2_inv_4 _0888_ (.A(\spi_shift_in[4] ),
    .Y(_0396_));
 sg13g2_inv_1 _0889_ (.Y(_0397_),
    .A(net303));
 sg13g2_inv_1 _0890_ (.Y(_0398_),
    .A(\reg_mode[1] ));
 sg13g2_inv_4 _0891_ (.A(\reg_thresh[6] ),
    .Y(_0399_));
 sg13g2_inv_1 _0892_ (.Y(_0400_),
    .A(\reg_thresh[5] ));
 sg13g2_inv_2 _0893_ (.Y(_0401_),
    .A(\reg_thresh[4] ));
 sg13g2_inv_1 _0894_ (.Y(_0402_),
    .A(net224));
 sg13g2_inv_1 _0895_ (.Y(_0403_),
    .A(net206));
 sg13g2_inv_1 _0896_ (.Y(_0404_),
    .A(\reg_thresh[1] ));
 sg13g2_inv_1 _0897_ (.Y(_0405_),
    .A(\spi_shift_out_load[1] ));
 sg13g2_inv_1 _0898_ (.Y(_0406_),
    .A(\spi_shift_out_load[2] ));
 sg13g2_inv_1 _0899_ (.Y(_0407_),
    .A(\spi_shift_out_load[3] ));
 sg13g2_inv_1 _0900_ (.Y(_0408_),
    .A(\spi_shift_out_load[4] ));
 sg13g2_inv_1 _0901_ (.Y(_0409_),
    .A(\spi_shift_out_load[5] ));
 sg13g2_inv_1 _0902_ (.Y(_0410_),
    .A(\spi_shift_out_load[6] ));
 sg13g2_inv_1 _0903_ (.Y(_0411_),
    .A(\spi_shift_out_load[7] ));
 sg13g2_inv_1 _0904_ (.Y(_0022_),
    .A(net286));
 sg13g2_inv_1 _0905_ (.Y(_0412_),
    .A(net212));
 sg13g2_inv_1 _0906_ (.Y(_0413_),
    .A(net230));
 sg13g2_inv_1 _0907_ (.Y(_0414_),
    .A(net210));
 sg13g2_inv_1 _0908_ (.Y(_0415_),
    .A(net359));
 sg13g2_inv_1 _0909_ (.Y(_0416_),
    .A(net228));
 sg13g2_inv_1 _0910_ (.Y(_0417_),
    .A(net226));
 sg13g2_inv_1 _0911_ (.Y(_0418_),
    .A(net222));
 sg13g2_and3_1 _0912_ (.X(_0005_),
    .A(net275),
    .B(net258),
    .C(\spi_shift_out_load[0] ));
 sg13g2_o21ai_1 _0913_ (.B1(net275),
    .Y(_0419_),
    .A1(net258),
    .A2(\spi_shift_out[1] ));
 sg13g2_a21oi_1 _0914_ (.A1(net258),
    .A2(_0405_),
    .Y(_0006_),
    .B1(_0419_));
 sg13g2_o21ai_1 _0915_ (.B1(net275),
    .Y(_0420_),
    .A1(net258),
    .A2(\spi_shift_out[2] ));
 sg13g2_a21oi_1 _0916_ (.A1(net258),
    .A2(_0406_),
    .Y(_0007_),
    .B1(_0420_));
 sg13g2_o21ai_1 _0917_ (.B1(net275),
    .Y(_0421_),
    .A1(net258),
    .A2(\spi_shift_out[3] ));
 sg13g2_a21oi_1 _0918_ (.A1(net258),
    .A2(_0407_),
    .Y(_0008_),
    .B1(_0421_));
 sg13g2_o21ai_1 _0919_ (.B1(net275),
    .Y(_0422_),
    .A1(net257),
    .A2(\spi_shift_out[4] ));
 sg13g2_a21oi_1 _0920_ (.A1(net257),
    .A2(_0408_),
    .Y(_0009_),
    .B1(_0422_));
 sg13g2_o21ai_1 _0921_ (.B1(net275),
    .Y(_0423_),
    .A1(net257),
    .A2(\spi_shift_out[5] ));
 sg13g2_a21oi_1 _0922_ (.A1(net257),
    .A2(_0409_),
    .Y(_0010_),
    .B1(_0423_));
 sg13g2_o21ai_1 _0923_ (.B1(_0030_),
    .Y(_0424_),
    .A1(net257),
    .A2(\spi_shift_out[6] ));
 sg13g2_a21oi_1 _0924_ (.A1(net257),
    .A2(_0410_),
    .Y(_0011_),
    .B1(_0424_));
 sg13g2_o21ai_1 _0925_ (.B1(_0030_),
    .Y(_0425_),
    .A1(net257),
    .A2(\spi_shift_out[7] ));
 sg13g2_a21oi_1 _0926_ (.A1(net257),
    .A2(_0411_),
    .Y(_0000_),
    .B1(_0425_));
 sg13g2_a21oi_1 _0927_ (.A1(\spi_bitcnt[0] ),
    .A2(_0014_),
    .Y(_0001_),
    .B1(net302));
 sg13g2_nor2b_2 _0928_ (.A(net302),
    .B_N(_0014_),
    .Y(_0426_));
 sg13g2_nand2_1 _0929_ (.Y(_0427_),
    .A(net275),
    .B(_0014_));
 sg13g2_xnor2_1 _0930_ (.Y(_0428_),
    .A(\spi_bitcnt[1] ),
    .B(\spi_bitcnt[0] ));
 sg13g2_nor2_1 _0931_ (.A(_0427_),
    .B(_0428_),
    .Y(_0002_));
 sg13g2_nand3_1 _0932_ (.B(\spi_bitcnt[0] ),
    .C(\spi_bitcnt[2] ),
    .A(\spi_bitcnt[1] ),
    .Y(_0429_));
 sg13g2_nand2_1 _0933_ (.Y(_0430_),
    .A(net247),
    .B(_0429_));
 sg13g2_a21oi_1 _0934_ (.A1(\spi_bitcnt[1] ),
    .A2(\spi_bitcnt[0] ),
    .Y(_0431_),
    .B1(\spi_bitcnt[2] ));
 sg13g2_nor2_1 _0935_ (.A(_0430_),
    .B(_0431_),
    .Y(_0003_));
 sg13g2_and3_1 _0936_ (.X(_0004_),
    .A(\spi_bitcnt[3] ),
    .B(net247),
    .C(_0429_));
 sg13g2_nor2_1 _0937_ (.A(\spi_bitcnt[3] ),
    .B(_0429_),
    .Y(_0432_));
 sg13g2_nand2b_2 _0938_ (.Y(_0433_),
    .B(_0432_),
    .A_N(_0013_));
 sg13g2_nor2_1 _0939_ (.A(\spi_shift_in[6] ),
    .B(_0433_),
    .Y(_0434_));
 sg13g2_nand2_2 _0940_ (.Y(_0435_),
    .A(net247),
    .B(_0434_));
 sg13g2_inv_1 _0941_ (.Y(_0012_),
    .A(net237));
 sg13g2_and2_1 _0942_ (.A(net10),
    .B(net1),
    .X(_0436_));
 sg13g2_nand2_2 _0943_ (.Y(_0437_),
    .A(net10),
    .B(net1));
 sg13g2_nand2_2 _0944_ (.Y(_0438_),
    .A(\pixel_q[7] ),
    .B(_0375_));
 sg13g2_xnor2_1 _0945_ (.Y(_0439_),
    .A(\pixel_q[7] ),
    .B(\prev_pixel[7] ));
 sg13g2_nor2b_1 _0946_ (.A(\prev_pixel[6] ),
    .B_N(net260),
    .Y(_0440_));
 sg13g2_xor2_1 _0947_ (.B(net260),
    .A(\prev_pixel[6] ),
    .X(_0441_));
 sg13g2_nor2_1 _0948_ (.A(_0377_),
    .B(\pixel_q[5] ),
    .Y(_0442_));
 sg13g2_nor2_1 _0949_ (.A(\prev_pixel[4] ),
    .B(_0380_),
    .Y(_0443_));
 sg13g2_xnor2_1 _0950_ (.Y(_0444_),
    .A(\prev_pixel[4] ),
    .B(\pixel_q[4] ));
 sg13g2_nand2_1 _0951_ (.Y(_0445_),
    .A(\prev_pixel[3] ),
    .B(_0382_));
 sg13g2_nor2_1 _0952_ (.A(\prev_pixel[3] ),
    .B(_0382_),
    .Y(_0446_));
 sg13g2_nand2_1 _0953_ (.Y(_0447_),
    .A(_0383_),
    .B(\pixel_q[2] ));
 sg13g2_xnor2_1 _0954_ (.Y(_0448_),
    .A(\prev_pixel[2] ),
    .B(\pixel_q[2] ));
 sg13g2_inv_1 _0955_ (.Y(_0449_),
    .A(_0448_));
 sg13g2_nor2b_1 _0956_ (.A(\prev_pixel[1] ),
    .B_N(\pixel_q[1] ),
    .Y(_0450_));
 sg13g2_nand2b_2 _0957_ (.Y(_0451_),
    .B(\prev_pixel[0] ),
    .A_N(\pixel_q[0] ));
 sg13g2_xnor2_1 _0958_ (.Y(_0452_),
    .A(\prev_pixel[1] ),
    .B(\pixel_q[1] ));
 sg13g2_a21oi_1 _0959_ (.A1(_0451_),
    .A2(_0452_),
    .Y(_0453_),
    .B1(_0450_));
 sg13g2_o21ai_1 _0960_ (.B1(_0447_),
    .Y(_0454_),
    .A1(_0449_),
    .A2(_0453_));
 sg13g2_a21o_2 _0961_ (.A2(_0454_),
    .A1(_0445_),
    .B1(_0446_),
    .X(_0455_));
 sg13g2_a21oi_1 _0962_ (.A1(_0444_),
    .A2(_0455_),
    .Y(_0456_),
    .B1(_0443_));
 sg13g2_a221oi_1 _0963_ (.B2(_0455_),
    .C1(_0443_),
    .B1(_0444_),
    .A1(_0377_),
    .Y(_0457_),
    .A2(\pixel_q[5] ));
 sg13g2_nor3_1 _0964_ (.A(_0441_),
    .B(_0442_),
    .C(_0457_),
    .Y(_0458_));
 sg13g2_o21ai_1 _0965_ (.B1(_0439_),
    .Y(_0459_),
    .A1(_0440_),
    .A2(_0458_));
 sg13g2_or3_1 _0966_ (.A(_0439_),
    .B(_0440_),
    .C(_0458_),
    .X(_0460_));
 sg13g2_nand2_1 _0967_ (.Y(_0461_),
    .A(_0459_),
    .B(_0460_));
 sg13g2_and2_1 _0968_ (.A(_0438_),
    .B(_0459_),
    .X(_0462_));
 sg13g2_xnor2_1 _0969_ (.Y(_0463_),
    .A(\pixel_q[0] ),
    .B(\prev_pixel[0] ));
 sg13g2_inv_1 _0970_ (.Y(_0464_),
    .A(_0463_));
 sg13g2_and2_1 _0971_ (.A(_0452_),
    .B(_0463_),
    .X(_0465_));
 sg13g2_nand2_1 _0972_ (.Y(_0466_),
    .A(_0452_),
    .B(_0463_));
 sg13g2_xnor2_1 _0973_ (.Y(_0467_),
    .A(\prev_pixel[3] ),
    .B(\pixel_q[3] ));
 sg13g2_xnor2_1 _0974_ (.Y(_0468_),
    .A(_0448_),
    .B(_0453_));
 sg13g2_nand2_1 _0975_ (.Y(_0469_),
    .A(_0448_),
    .B(_0465_));
 sg13g2_and3_1 _0976_ (.X(_0470_),
    .A(_0448_),
    .B(_0465_),
    .C(_0467_));
 sg13g2_inv_1 _0977_ (.Y(_0471_),
    .A(_0470_));
 sg13g2_xnor2_1 _0978_ (.Y(_0472_),
    .A(\prev_pixel[5] ),
    .B(\pixel_q[5] ));
 sg13g2_nand3_1 _0979_ (.B(_0470_),
    .C(_0472_),
    .A(_0444_),
    .Y(_0473_));
 sg13g2_nand2_1 _0980_ (.Y(_0474_),
    .A(_0462_),
    .B(_0473_));
 sg13g2_o21ai_1 _0981_ (.B1(_0462_),
    .Y(_0475_),
    .A1(_0441_),
    .A2(_0473_));
 sg13g2_xor2_1 _0982_ (.B(_0475_),
    .A(_0461_),
    .X(_0476_));
 sg13g2_a21oi_1 _0983_ (.A1(\reg_edge_thr[0] ),
    .A2(_0463_),
    .Y(_0477_),
    .B1(\reg_edge_thr[1] ));
 sg13g2_xnor2_1 _0984_ (.Y(_0478_),
    .A(_0451_),
    .B(_0452_));
 sg13g2_nand3_1 _0985_ (.B(_0459_),
    .C(_0464_),
    .A(_0438_),
    .Y(_0479_));
 sg13g2_xor2_1 _0986_ (.B(_0479_),
    .A(_0478_),
    .X(_0480_));
 sg13g2_nand3_1 _0987_ (.B(_0459_),
    .C(_0466_),
    .A(_0438_),
    .Y(_0481_));
 sg13g2_xor2_1 _0988_ (.B(_0481_),
    .A(_0468_),
    .X(_0482_));
 sg13g2_xnor2_1 _0989_ (.Y(_0483_),
    .A(_0468_),
    .B(_0481_));
 sg13g2_nor2_1 _0990_ (.A(_0018_),
    .B(_0483_),
    .Y(_0484_));
 sg13g2_nand3_1 _0991_ (.B(\reg_edge_thr[1] ),
    .C(_0463_),
    .A(\reg_edge_thr[0] ),
    .Y(_0485_));
 sg13g2_a21oi_1 _0992_ (.A1(_0480_),
    .A2(_0485_),
    .Y(_0486_),
    .B1(_0477_));
 sg13g2_xor2_1 _0993_ (.B(_0467_),
    .A(_0454_),
    .X(_0487_));
 sg13g2_nand3_1 _0994_ (.B(_0459_),
    .C(_0469_),
    .A(_0438_),
    .Y(_0488_));
 sg13g2_xor2_1 _0995_ (.B(_0488_),
    .A(_0487_),
    .X(_0489_));
 sg13g2_xnor2_1 _0996_ (.Y(_0490_),
    .A(_0487_),
    .B(_0488_));
 sg13g2_a22oi_1 _0997_ (.Y(_0491_),
    .B1(_0490_),
    .B2(_0019_),
    .A2(_0483_),
    .A1(_0018_));
 sg13g2_o21ai_1 _0998_ (.B1(_0491_),
    .Y(_0492_),
    .A1(_0484_),
    .A2(_0486_));
 sg13g2_xnor2_1 _0999_ (.Y(_0493_),
    .A(_0444_),
    .B(_0455_));
 sg13g2_nand3_1 _1000_ (.B(_0459_),
    .C(_0471_),
    .A(_0438_),
    .Y(_0494_));
 sg13g2_xnor2_1 _1001_ (.Y(_0495_),
    .A(_0493_),
    .B(_0494_));
 sg13g2_inv_1 _1002_ (.Y(_0496_),
    .A(_0495_));
 sg13g2_a22oi_1 _1003_ (.Y(_0497_),
    .B1(_0495_),
    .B2(\reg_edge_thr[4] ),
    .A2(_0489_),
    .A1(_0369_));
 sg13g2_nand2_1 _1004_ (.Y(_0498_),
    .A(_0470_),
    .B(_0493_));
 sg13g2_nand3_1 _1005_ (.B(_0459_),
    .C(_0498_),
    .A(_0438_),
    .Y(_0499_));
 sg13g2_xor2_1 _1006_ (.B(_0472_),
    .A(_0456_),
    .X(_0500_));
 sg13g2_xnor2_1 _1007_ (.Y(_0501_),
    .A(_0499_),
    .B(_0500_));
 sg13g2_or2_1 _1008_ (.X(_0502_),
    .B(_0501_),
    .A(\reg_edge_thr[5] ));
 sg13g2_o21ai_1 _1009_ (.B1(_0502_),
    .Y(_0503_),
    .A1(\reg_edge_thr[4] ),
    .A2(_0495_));
 sg13g2_a21oi_1 _1010_ (.A1(_0492_),
    .A2(_0497_),
    .Y(_0504_),
    .B1(_0503_));
 sg13g2_o21ai_1 _1011_ (.B1(_0441_),
    .Y(_0505_),
    .A1(_0442_),
    .A2(_0457_));
 sg13g2_nor2b_1 _1012_ (.A(_0458_),
    .B_N(_0505_),
    .Y(_0506_));
 sg13g2_xnor2_1 _1013_ (.Y(_0507_),
    .A(_0474_),
    .B(_0506_));
 sg13g2_nand2_1 _1014_ (.Y(_0508_),
    .A(\reg_edge_thr[5] ),
    .B(_0501_));
 sg13g2_o21ai_1 _1015_ (.B1(_0508_),
    .Y(_0509_),
    .A1(_0386_),
    .A2(_0507_));
 sg13g2_a22oi_1 _1016_ (.Y(_0510_),
    .B1(_0507_),
    .B2(_0386_),
    .A2(_0476_),
    .A1(_0385_));
 sg13g2_o21ai_1 _1017_ (.B1(_0510_),
    .Y(_0511_),
    .A1(_0504_),
    .A2(_0509_));
 sg13g2_o21ai_1 _1018_ (.B1(_0511_),
    .Y(_0512_),
    .A1(_0385_),
    .A2(_0476_));
 sg13g2_nand2_1 _1019_ (.Y(_0513_),
    .A(net158),
    .B(net261));
 sg13g2_o21ai_1 _1020_ (.B1(_0513_),
    .Y(_0031_),
    .A1(net261),
    .A2(_0512_));
 sg13g2_nor2b_2 _1021_ (.A(\mean_q[7] ),
    .B_N(\pixel_q[7] ),
    .Y(_0514_));
 sg13g2_xnor2_1 _1022_ (.Y(_0515_),
    .A(\pixel_q[7] ),
    .B(\mean_q[7] ));
 sg13g2_nand2_1 _1023_ (.Y(_0516_),
    .A(net260),
    .B(_0388_));
 sg13g2_nor2_1 _1024_ (.A(net260),
    .B(_0388_),
    .Y(_0517_));
 sg13g2_xnor2_1 _1025_ (.Y(_0518_),
    .A(net260),
    .B(\mean_q[6] ));
 sg13g2_nor2b_1 _1026_ (.A(\mean_q[3] ),
    .B_N(\pixel_q[3] ),
    .Y(_0519_));
 sg13g2_nand2b_1 _1027_ (.Y(_0520_),
    .B(\mean_q[3] ),
    .A_N(\pixel_q[3] ));
 sg13g2_xor2_1 _1028_ (.B(\mean_q[3] ),
    .A(\pixel_q[3] ),
    .X(_0521_));
 sg13g2_nor2b_1 _1029_ (.A(\mean_q[2] ),
    .B_N(\pixel_q[2] ),
    .Y(_0522_));
 sg13g2_xnor2_1 _1030_ (.Y(_0523_),
    .A(\pixel_q[2] ),
    .B(\mean_q[2] ));
 sg13g2_nand2b_1 _1031_ (.Y(_0524_),
    .B(_0523_),
    .A_N(_0521_));
 sg13g2_nor2b_1 _1032_ (.A(\mean_q[1] ),
    .B_N(\pixel_q[1] ),
    .Y(_0525_));
 sg13g2_nand2b_2 _1033_ (.Y(_0526_),
    .B(\mean_q[0] ),
    .A_N(\pixel_q[0] ));
 sg13g2_xnor2_1 _1034_ (.Y(_0527_),
    .A(\pixel_q[1] ),
    .B(\mean_q[1] ));
 sg13g2_a21oi_1 _1035_ (.A1(_0526_),
    .A2(_0527_),
    .Y(_0528_),
    .B1(_0525_));
 sg13g2_a21oi_1 _1036_ (.A1(_0520_),
    .A2(_0522_),
    .Y(_0529_),
    .B1(_0519_));
 sg13g2_o21ai_1 _1037_ (.B1(_0529_),
    .Y(_0530_),
    .A1(_0524_),
    .A2(_0528_));
 sg13g2_nor2_1 _1038_ (.A(_0380_),
    .B(\mean_q[4] ),
    .Y(_0531_));
 sg13g2_xnor2_1 _1039_ (.Y(_0532_),
    .A(\pixel_q[4] ),
    .B(\mean_q[4] ));
 sg13g2_nor2b_1 _1040_ (.A(\mean_q[5] ),
    .B_N(\pixel_q[5] ),
    .Y(_0533_));
 sg13g2_nand2b_1 _1041_ (.Y(_0534_),
    .B(\mean_q[5] ),
    .A_N(\pixel_q[5] ));
 sg13g2_nor2b_1 _1042_ (.A(_0533_),
    .B_N(_0534_),
    .Y(_0535_));
 sg13g2_and2_1 _1043_ (.A(_0532_),
    .B(_0535_),
    .X(_0536_));
 sg13g2_a221oi_1 _1044_ (.B2(_0530_),
    .C1(_0533_),
    .B1(_0536_),
    .A1(_0531_),
    .Y(_0537_),
    .A2(_0534_));
 sg13g2_o21ai_1 _1045_ (.B1(_0516_),
    .Y(_0538_),
    .A1(_0517_),
    .A2(_0537_));
 sg13g2_a21oi_2 _1046_ (.B1(_0514_),
    .Y(_0539_),
    .A2(_0538_),
    .A1(_0515_));
 sg13g2_a21o_2 _1047_ (.A2(_0538_),
    .A1(_0515_),
    .B1(_0514_),
    .X(_0540_));
 sg13g2_xor2_1 _1048_ (.B(_0538_),
    .A(_0515_),
    .X(_0541_));
 sg13g2_xnor2_1 _1049_ (.Y(_0542_),
    .A(_0515_),
    .B(_0538_));
 sg13g2_nand2_1 _1050_ (.Y(_0543_),
    .A(_0370_),
    .B(\pixel_q[0] ));
 sg13g2_and2_1 _1051_ (.A(_0526_),
    .B(_0543_),
    .X(_0544_));
 sg13g2_nand2_1 _1052_ (.Y(_0545_),
    .A(_0527_),
    .B(_0544_));
 sg13g2_or2_1 _1053_ (.X(_0546_),
    .B(_0545_),
    .A(_0524_));
 sg13g2_inv_1 _1054_ (.Y(_0547_),
    .A(_0546_));
 sg13g2_nand2_1 _1055_ (.Y(_0548_),
    .A(_0536_),
    .B(_0547_));
 sg13g2_xnor2_1 _1056_ (.Y(_0549_),
    .A(_0518_),
    .B(_0537_));
 sg13g2_o21ai_1 _1057_ (.B1(_0539_),
    .Y(_0550_),
    .A1(_0548_),
    .A2(_0549_));
 sg13g2_xnor2_1 _1058_ (.Y(_0551_),
    .A(_0541_),
    .B(_0550_));
 sg13g2_xnor2_1 _1059_ (.Y(_0552_),
    .A(_0542_),
    .B(_0550_));
 sg13g2_nand2_1 _1060_ (.Y(_0553_),
    .A(net404),
    .B(_0552_));
 sg13g2_nand2b_1 _1061_ (.Y(_0554_),
    .B(_0523_),
    .A_N(_0528_));
 sg13g2_xnor2_1 _1062_ (.Y(_0555_),
    .A(_0523_),
    .B(_0528_));
 sg13g2_nand2_1 _1063_ (.Y(_0556_),
    .A(_0539_),
    .B(_0545_));
 sg13g2_xnor2_1 _1064_ (.Y(_0557_),
    .A(_0555_),
    .B(_0556_));
 sg13g2_a21o_1 _1065_ (.A2(_0544_),
    .A1(\reg_contrast_thr[0] ),
    .B1(\reg_contrast_thr[1] ),
    .X(_0558_));
 sg13g2_and3_1 _1066_ (.X(_0559_),
    .A(\reg_contrast_thr[1] ),
    .B(\reg_contrast_thr[0] ),
    .C(_0544_));
 sg13g2_xor2_1 _1067_ (.B(_0527_),
    .A(_0526_),
    .X(_0560_));
 sg13g2_a221oi_1 _1068_ (.B2(_0526_),
    .C1(_0514_),
    .B1(_0543_),
    .A1(_0515_),
    .Y(_0561_),
    .A2(_0538_));
 sg13g2_xnor2_1 _1069_ (.Y(_0562_),
    .A(_0560_),
    .B(_0561_));
 sg13g2_a21oi_1 _1070_ (.A1(_0558_),
    .A2(_0562_),
    .Y(_0563_),
    .B1(_0559_));
 sg13g2_o21ai_1 _1071_ (.B1(_0563_),
    .Y(_0564_),
    .A1(_0016_),
    .A2(_0557_));
 sg13g2_nor2b_1 _1072_ (.A(_0522_),
    .B_N(_0554_),
    .Y(_0565_));
 sg13g2_xnor2_1 _1073_ (.Y(_0566_),
    .A(_0521_),
    .B(_0565_));
 sg13g2_o21ai_1 _1074_ (.B1(_0539_),
    .Y(_0567_),
    .A1(_0545_),
    .A2(_0555_));
 sg13g2_xnor2_1 _1075_ (.Y(_0568_),
    .A(_0566_),
    .B(_0567_));
 sg13g2_xor2_1 _1076_ (.B(_0567_),
    .A(_0566_),
    .X(_0569_));
 sg13g2_a22oi_1 _1077_ (.Y(_0570_),
    .B1(_0569_),
    .B2(_0017_),
    .A2(_0557_),
    .A1(_0016_));
 sg13g2_nand2_1 _1078_ (.Y(_0571_),
    .A(_0539_),
    .B(_0546_));
 sg13g2_xnor2_1 _1079_ (.Y(_0572_),
    .A(_0530_),
    .B(_0532_));
 sg13g2_xnor2_1 _1080_ (.Y(_0573_),
    .A(_0571_),
    .B(_0572_));
 sg13g2_inv_1 _1081_ (.Y(_0574_),
    .A(_0573_));
 sg13g2_nor2_1 _1082_ (.A(_0017_),
    .B(_0569_),
    .Y(_0575_));
 sg13g2_a221oi_1 _1083_ (.B2(\reg_contrast_thr[4] ),
    .C1(_0575_),
    .B1(_0573_),
    .A1(_0564_),
    .Y(_0576_),
    .A2(_0570_));
 sg13g2_nor2_1 _1084_ (.A(\reg_contrast_thr[4] ),
    .B(_0573_),
    .Y(_0577_));
 sg13g2_a21o_1 _1085_ (.A2(_0547_),
    .A1(_0532_),
    .B1(_0540_),
    .X(_0578_));
 sg13g2_a21oi_1 _1086_ (.A1(_0530_),
    .A2(_0532_),
    .Y(_0579_),
    .B1(_0531_));
 sg13g2_xor2_1 _1087_ (.B(_0579_),
    .A(_0535_),
    .X(_0580_));
 sg13g2_inv_1 _1088_ (.Y(_0581_),
    .A(_0580_));
 sg13g2_xnor2_1 _1089_ (.Y(_0582_),
    .A(_0578_),
    .B(_0580_));
 sg13g2_inv_1 _1090_ (.Y(_0583_),
    .A(_0582_));
 sg13g2_nor2_1 _1091_ (.A(\reg_contrast_thr[5] ),
    .B(_0582_),
    .Y(_0584_));
 sg13g2_nor3_1 _1092_ (.A(_0576_),
    .B(_0577_),
    .C(_0584_),
    .Y(_0585_));
 sg13g2_nand2_1 _1093_ (.Y(_0586_),
    .A(_0539_),
    .B(_0548_));
 sg13g2_xor2_1 _1094_ (.B(_0586_),
    .A(_0549_),
    .X(_0587_));
 sg13g2_a221oi_1 _1095_ (.B2(\reg_contrast_thr[6] ),
    .C1(_0585_),
    .B1(_0587_),
    .A1(\reg_contrast_thr[5] ),
    .Y(_0588_),
    .A2(_0582_));
 sg13g2_nand2_1 _1096_ (.Y(_0589_),
    .A(_0393_),
    .B(_0551_));
 sg13g2_o21ai_1 _1097_ (.B1(_0589_),
    .Y(_0590_),
    .A1(\reg_contrast_thr[6] ),
    .A2(_0587_));
 sg13g2_o21ai_1 _1098_ (.B1(_0553_),
    .Y(_0591_),
    .A1(_0588_),
    .A2(_0590_));
 sg13g2_or2_1 _1099_ (.X(_0592_),
    .B(_0591_),
    .A(_0540_));
 sg13g2_nand2_1 _1100_ (.Y(_0593_),
    .A(net160),
    .B(net273));
 sg13g2_o21ai_1 _1101_ (.B1(_0593_),
    .Y(_0032_),
    .A1(net273),
    .A2(_0592_));
 sg13g2_nand2b_1 _1102_ (.Y(_0594_),
    .B(_0540_),
    .A_N(_0591_));
 sg13g2_nand2_1 _1103_ (.Y(_0595_),
    .A(net157),
    .B(net273));
 sg13g2_o21ai_1 _1104_ (.B1(_0595_),
    .Y(_0033_),
    .A1(net273),
    .A2(_0594_));
 sg13g2_a21oi_1 _1105_ (.A1(_0512_),
    .A2(_0591_),
    .Y(_0596_),
    .B1(net261));
 sg13g2_a21o_1 _1106_ (.A2(net261),
    .A1(net178),
    .B1(_0596_),
    .X(_0034_));
 sg13g2_and2_1 _1107_ (.A(\reg_thresh[0] ),
    .B(net327),
    .X(_0035_));
 sg13g2_and2_1 _1108_ (.A(\reg_thresh[1] ),
    .B(net327),
    .X(_0036_));
 sg13g2_and2_1 _1109_ (.A(\reg_thresh[2] ),
    .B(net341),
    .X(_0037_));
 sg13g2_and2_1 _1110_ (.A(\reg_thresh[3] ),
    .B(net327),
    .X(_0038_));
 sg13g2_and2_1 _1111_ (.A(\reg_thresh[4] ),
    .B(net322),
    .X(_0039_));
 sg13g2_and2_1 _1112_ (.A(\reg_thresh[5] ),
    .B(net320),
    .X(_0040_));
 sg13g2_and2_1 _1113_ (.A(\reg_thresh[6] ),
    .B(net320),
    .X(_0041_));
 sg13g2_nor2b_1 _1114_ (.A(_0015_),
    .B_N(net308),
    .Y(_0042_));
 sg13g2_and2_1 _1115_ (.A(\reg_contrast_thr[0] ),
    .B(net339),
    .X(_0043_));
 sg13g2_and2_1 _1116_ (.A(\reg_contrast_thr[1] ),
    .B(net339),
    .X(_0044_));
 sg13g2_nor2b_1 _1117_ (.A(_0016_),
    .B_N(net327),
    .Y(_0045_));
 sg13g2_nor2b_1 _1118_ (.A(_0017_),
    .B_N(net330),
    .Y(_0046_));
 sg13g2_and2_1 _1119_ (.A(\reg_contrast_thr[4] ),
    .B(net321),
    .X(_0047_));
 sg13g2_and2_1 _1120_ (.A(\reg_contrast_thr[5] ),
    .B(net308),
    .X(_0048_));
 sg13g2_and2_1 _1121_ (.A(\reg_contrast_thr[6] ),
    .B(net305),
    .X(_0049_));
 sg13g2_and2_1 _1122_ (.A(\reg_contrast_thr[7] ),
    .B(net317),
    .X(_0050_));
 sg13g2_and2_1 _1123_ (.A(\reg_edge_thr[0] ),
    .B(net340),
    .X(_0051_));
 sg13g2_and2_1 _1124_ (.A(\reg_edge_thr[1] ),
    .B(net340),
    .X(_0052_));
 sg13g2_nor2b_1 _1125_ (.A(_0018_),
    .B_N(net340),
    .Y(_0053_));
 sg13g2_nor2b_1 _1126_ (.A(_0019_),
    .B_N(net330),
    .Y(_0054_));
 sg13g2_and2_1 _1127_ (.A(\reg_edge_thr[4] ),
    .B(net308),
    .X(_0055_));
 sg13g2_and2_1 _1128_ (.A(\reg_edge_thr[5] ),
    .B(net308),
    .X(_0056_));
 sg13g2_and2_1 _1129_ (.A(\reg_edge_thr[6] ),
    .B(net309),
    .X(_0057_));
 sg13g2_and2_1 _1130_ (.A(\reg_edge_thr[7] ),
    .B(net309),
    .X(_0058_));
 sg13g2_nor2b_1 _1131_ (.A(net256),
    .B_N(net345),
    .Y(_0059_));
 sg13g2_nor2b_1 _1132_ (.A(net254),
    .B_N(net341),
    .Y(_0060_));
 sg13g2_and2_1 _1133_ (.A(net253),
    .B(net345),
    .X(_0061_));
 sg13g2_and2_1 _1134_ (.A(net250),
    .B(net341),
    .X(_0062_));
 sg13g2_and2_1 _1135_ (.A(\reg_mode[1] ),
    .B(net335),
    .X(_0063_));
 sg13g2_and2_1 _1136_ (.A(net318),
    .B(\reg_mode[2] ),
    .X(_0064_));
 sg13g2_and2_1 _1137_ (.A(net320),
    .B(\reg_mode[3] ),
    .X(_0065_));
 sg13g2_and2_1 _1138_ (.A(net306),
    .B(\reg_mode[4] ),
    .X(_0066_));
 sg13g2_and2_1 _1139_ (.A(net306),
    .B(\reg_mode[5] ),
    .X(_0067_));
 sg13g2_and2_1 _1140_ (.A(net306),
    .B(\reg_mode[6] ),
    .X(_0068_));
 sg13g2_and2_1 _1141_ (.A(net307),
    .B(\reg_mode[7] ),
    .X(_0069_));
 sg13g2_and2_1 _1142_ (.A(\reg_status[4] ),
    .B(net316),
    .X(_0070_));
 sg13g2_and2_1 _1143_ (.A(\reg_status[5] ),
    .B(net337),
    .X(_0071_));
 sg13g2_and2_1 _1144_ (.A(\reg_status[6] ),
    .B(net335),
    .X(_0072_));
 sg13g2_and2_1 _1145_ (.A(\reg_status[7] ),
    .B(net316),
    .X(_0073_));
 sg13g2_and2_1 _1146_ (.A(\mean_q[0] ),
    .B(net347),
    .X(_0074_));
 sg13g2_and2_1 _1147_ (.A(\mean_q[1] ),
    .B(net347),
    .X(_0075_));
 sg13g2_and2_1 _1148_ (.A(\mean_q[2] ),
    .B(net346),
    .X(_0076_));
 sg13g2_and2_1 _1149_ (.A(\mean_q[3] ),
    .B(net346),
    .X(_0077_));
 sg13g2_and2_1 _1150_ (.A(\mean_q[4] ),
    .B(net341),
    .X(_0078_));
 sg13g2_and2_1 _1151_ (.A(\mean_q[5] ),
    .B(net348),
    .X(_0079_));
 sg13g2_and2_1 _1152_ (.A(\mean_q[6] ),
    .B(net348),
    .X(_0080_));
 sg13g2_and2_1 _1153_ (.A(\mean_q[7] ),
    .B(net345),
    .X(_0081_));
 sg13g2_and2_1 _1154_ (.A(net343),
    .B(\reg_absdiff_rdback[0] ),
    .X(_0082_));
 sg13g2_and2_1 _1155_ (.A(net344),
    .B(\reg_absdiff_rdback[1] ),
    .X(_0083_));
 sg13g2_and2_1 _1156_ (.A(net346),
    .B(\reg_absdiff_rdback[2] ),
    .X(_0084_));
 sg13g2_and2_1 _1157_ (.A(net327),
    .B(\reg_absdiff_rdback[3] ),
    .X(_0085_));
 sg13g2_and2_1 _1158_ (.A(net320),
    .B(\reg_absdiff_rdback[4] ),
    .X(_0086_));
 sg13g2_and2_1 _1159_ (.A(net326),
    .B(\reg_absdiff_rdback[5] ),
    .X(_0087_));
 sg13g2_and2_1 _1160_ (.A(net308),
    .B(\reg_absdiff_rdback[6] ),
    .X(_0088_));
 sg13g2_and2_1 _1161_ (.A(net317),
    .B(\reg_absdiff_rdback[7] ),
    .X(_0089_));
 sg13g2_nand2_1 _1162_ (.Y(_0597_),
    .A(net161),
    .B(net264));
 sg13g2_o21ai_1 _1163_ (.B1(_0597_),
    .Y(_0090_),
    .A1(net264),
    .A2(_0544_));
 sg13g2_nand2_1 _1164_ (.Y(_0598_),
    .A(net155),
    .B(net264));
 sg13g2_o21ai_1 _1165_ (.B1(_0598_),
    .Y(_0091_),
    .A1(net264),
    .A2(_0562_));
 sg13g2_mux2_1 _1166_ (.A0(net188),
    .A1(_0557_),
    .S(_0436_),
    .X(_0092_));
 sg13g2_nand2_1 _1167_ (.Y(_0599_),
    .A(net156),
    .B(net263));
 sg13g2_o21ai_1 _1168_ (.B1(_0599_),
    .Y(_0093_),
    .A1(net263),
    .A2(_0568_));
 sg13g2_nand2_1 _1169_ (.Y(_0600_),
    .A(net170),
    .B(net262));
 sg13g2_o21ai_1 _1170_ (.B1(_0600_),
    .Y(_0094_),
    .A1(net262),
    .A2(_0573_));
 sg13g2_nand2_1 _1171_ (.Y(_0601_),
    .A(net154),
    .B(net263));
 sg13g2_o21ai_1 _1172_ (.B1(_0601_),
    .Y(_0095_),
    .A1(net262),
    .A2(_0582_));
 sg13g2_nand2_1 _1173_ (.Y(_0602_),
    .A(net162),
    .B(net261));
 sg13g2_o21ai_1 _1174_ (.B1(_0602_),
    .Y(_0096_),
    .A1(net261),
    .A2(_0587_));
 sg13g2_nand2_1 _1175_ (.Y(_0603_),
    .A(net159),
    .B(net261));
 sg13g2_o21ai_1 _1176_ (.B1(_0603_),
    .Y(_0097_),
    .A1(net261),
    .A2(_0552_));
 sg13g2_nor2_1 _1177_ (.A(net2),
    .B(net269),
    .Y(_0604_));
 sg13g2_a21oi_1 _1178_ (.A1(_0371_),
    .A2(net270),
    .Y(_0098_),
    .B1(_0604_));
 sg13g2_nor2_1 _1179_ (.A(net3),
    .B(net273),
    .Y(_0605_));
 sg13g2_a21oi_1 _1180_ (.A1(_0374_),
    .A2(net273),
    .Y(_0099_),
    .B1(_0605_));
 sg13g2_nor2_1 _1181_ (.A(net4),
    .B(net273),
    .Y(_0606_));
 sg13g2_a21oi_1 _1182_ (.A1(_0384_),
    .A2(net273),
    .Y(_0100_),
    .B1(_0606_));
 sg13g2_nor2_1 _1183_ (.A(net5),
    .B(net269),
    .Y(_0607_));
 sg13g2_a21oi_1 _1184_ (.A1(_0382_),
    .A2(net269),
    .Y(_0101_),
    .B1(_0607_));
 sg13g2_nor2_1 _1185_ (.A(net6),
    .B(net267),
    .Y(_0608_));
 sg13g2_a21oi_1 _1186_ (.A1(_0380_),
    .A2(net267),
    .Y(_0102_),
    .B1(_0608_));
 sg13g2_nor2_1 _1187_ (.A(net7),
    .B(net267),
    .Y(_0609_));
 sg13g2_a21oi_1 _1188_ (.A1(_0378_),
    .A2(net265),
    .Y(_0103_),
    .B1(_0609_));
 sg13g2_mux2_1 _1189_ (.A0(net352),
    .A1(net8),
    .S(_0436_),
    .X(_0104_));
 sg13g2_mux2_1 _1190_ (.A0(net402),
    .A1(net9),
    .S(_0436_),
    .X(_0105_));
 sg13g2_a21oi_1 _1191_ (.A1(net2),
    .A2(net303),
    .Y(_0610_),
    .B1(net270));
 sg13g2_nand2_1 _1192_ (.Y(_0611_),
    .A(\pixel_q[0] ),
    .B(net274));
 sg13g2_a22oi_1 _1193_ (.Y(_0106_),
    .B1(_0610_),
    .B2(_0611_),
    .A2(net270),
    .A1(_0372_));
 sg13g2_a21oi_1 _1194_ (.A1(net303),
    .A2(net3),
    .Y(_0612_),
    .B1(net271));
 sg13g2_nand2_1 _1195_ (.Y(_0613_),
    .A(\pixel_q[1] ),
    .B(net274));
 sg13g2_a22oi_1 _1196_ (.Y(_0107_),
    .B1(_0612_),
    .B2(_0613_),
    .A2(net271),
    .A1(_0373_));
 sg13g2_a21oi_1 _1197_ (.A1(net303),
    .A2(net4),
    .Y(_0614_),
    .B1(net271));
 sg13g2_nand2_1 _1198_ (.Y(_0615_),
    .A(\pixel_q[2] ),
    .B(net274));
 sg13g2_a22oi_1 _1199_ (.Y(_0108_),
    .B1(_0614_),
    .B2(_0615_),
    .A2(net271),
    .A1(_0383_));
 sg13g2_a21oi_1 _1200_ (.A1(net303),
    .A2(net5),
    .Y(_0616_),
    .B1(net270));
 sg13g2_nand2_1 _1201_ (.Y(_0617_),
    .A(\pixel_q[3] ),
    .B(net274));
 sg13g2_a22oi_1 _1202_ (.Y(_0109_),
    .B1(_0616_),
    .B2(_0617_),
    .A2(net270),
    .A1(_0381_));
 sg13g2_a21oi_1 _1203_ (.A1(net304),
    .A2(net6),
    .Y(_0618_),
    .B1(net269));
 sg13g2_nand2_1 _1204_ (.Y(_0619_),
    .A(\pixel_q[4] ),
    .B(net274));
 sg13g2_a22oi_1 _1205_ (.Y(_0110_),
    .B1(_0618_),
    .B2(_0619_),
    .A2(net269),
    .A1(_0379_));
 sg13g2_a21oi_1 _1206_ (.A1(net304),
    .A2(net7),
    .Y(_0620_),
    .B1(net269));
 sg13g2_nand2_1 _1207_ (.Y(_0621_),
    .A(\pixel_q[5] ),
    .B(net274));
 sg13g2_a22oi_1 _1208_ (.Y(_0111_),
    .B1(_0620_),
    .B2(_0621_),
    .A2(net265),
    .A1(_0377_));
 sg13g2_a21oi_1 _1209_ (.A1(net304),
    .A2(net8),
    .Y(_0622_),
    .B1(net267));
 sg13g2_nand2_1 _1210_ (.Y(_0623_),
    .A(net260),
    .B(net274));
 sg13g2_a22oi_1 _1211_ (.Y(_0112_),
    .B1(_0622_),
    .B2(_0623_),
    .A2(net265),
    .A1(_0376_));
 sg13g2_a21oi_1 _1212_ (.A1(net304),
    .A2(net9),
    .Y(_0624_),
    .B1(net265));
 sg13g2_nand2_1 _1213_ (.Y(_0625_),
    .A(\pixel_q[7] ),
    .B(net274));
 sg13g2_a22oi_1 _1214_ (.Y(_0113_),
    .B1(_0624_),
    .B2(_0625_),
    .A2(net265),
    .A1(_0375_));
 sg13g2_and2_1 _1215_ (.A(net255),
    .B(_0549_),
    .X(_0626_));
 sg13g2_a21oi_1 _1216_ (.A1(_0368_),
    .A2(_0541_),
    .Y(_0627_),
    .B1(_0626_));
 sg13g2_a21o_1 _1217_ (.A2(_0541_),
    .A1(_0368_),
    .B1(_0626_),
    .X(_0628_));
 sg13g2_or2_1 _1218_ (.X(_0629_),
    .B(_0572_),
    .A(_0368_));
 sg13g2_o21ai_1 _1219_ (.B1(_0629_),
    .Y(_0630_),
    .A1(net255),
    .A2(_0580_));
 sg13g2_or2_1 _1220_ (.X(_0631_),
    .B(_0630_),
    .A(_0367_));
 sg13g2_o21ai_1 _1221_ (.B1(_0631_),
    .Y(_0632_),
    .A1(net254),
    .A2(_0628_));
 sg13g2_nand2_1 _1222_ (.Y(_0633_),
    .A(net255),
    .B(_0555_));
 sg13g2_o21ai_1 _1223_ (.B1(_0633_),
    .Y(_0634_),
    .A1(net255),
    .A2(_0566_));
 sg13g2_nand2_1 _1224_ (.Y(_0635_),
    .A(_0367_),
    .B(_0634_));
 sg13g2_o21ai_1 _1225_ (.B1(net254),
    .Y(_0636_),
    .A1(net255),
    .A2(_0560_));
 sg13g2_a21oi_1 _1226_ (.A1(net256),
    .A2(_0544_),
    .Y(_0637_),
    .B1(_0636_));
 sg13g2_nor2_1 _1227_ (.A(net251),
    .B(_0637_),
    .Y(_0638_));
 sg13g2_a22oi_1 _1228_ (.Y(_0639_),
    .B1(_0635_),
    .B2(_0638_),
    .A2(_0632_),
    .A1(net252));
 sg13g2_a221oi_1 _1229_ (.B2(_0638_),
    .C1(_0370_),
    .B1(_0635_),
    .A1(net252),
    .Y(_0640_),
    .A2(_0632_));
 sg13g2_o21ai_1 _1230_ (.B1(_0397_),
    .Y(_0641_),
    .A1(net393),
    .A2(_0639_));
 sg13g2_o21ai_1 _1231_ (.B1(_0610_),
    .Y(_0642_),
    .A1(_0640_),
    .A2(_0641_));
 sg13g2_o21ai_1 _1232_ (.B1(_0642_),
    .Y(_0643_),
    .A1(net393),
    .A2(_0436_));
 sg13g2_inv_1 _1233_ (.Y(_0114_),
    .A(_0643_));
 sg13g2_mux2_1 _1234_ (.A0(_0566_),
    .A1(_0572_),
    .S(_0368_),
    .X(_0644_));
 sg13g2_nand2_1 _1235_ (.Y(_0645_),
    .A(_0368_),
    .B(_0555_));
 sg13g2_a21oi_1 _1236_ (.A1(net256),
    .A2(_0560_),
    .Y(_0646_),
    .B1(_0367_));
 sg13g2_a221oi_1 _1237_ (.B2(_0646_),
    .C1(net252),
    .B1(_0645_),
    .A1(_0367_),
    .Y(_0647_),
    .A2(_0644_));
 sg13g2_mux2_1 _1238_ (.A0(_0540_),
    .A1(_0542_),
    .S(net255),
    .X(_0648_));
 sg13g2_nor2_1 _1239_ (.A(_0368_),
    .B(_0580_),
    .Y(_0649_));
 sg13g2_a21oi_1 _1240_ (.A1(_0368_),
    .A2(_0549_),
    .Y(_0650_),
    .B1(_0649_));
 sg13g2_mux4_1 _1241_ (.S0(net255),
    .A0(_0539_),
    .A1(_0541_),
    .A2(_0549_),
    .A3(_0581_),
    .S1(net254),
    .X(_0651_));
 sg13g2_a21oi_1 _1242_ (.A1(net252),
    .A2(_0651_),
    .Y(_0652_),
    .B1(_0647_));
 sg13g2_nor2_1 _1243_ (.A(_0392_),
    .B(_0652_),
    .Y(_0653_));
 sg13g2_xnor2_1 _1244_ (.Y(_0654_),
    .A(net391),
    .B(_0652_));
 sg13g2_a21oi_1 _1245_ (.A1(_0640_),
    .A2(_0654_),
    .Y(_0655_),
    .B1(net303));
 sg13g2_o21ai_1 _1246_ (.B1(_0655_),
    .Y(_0656_),
    .A1(_0640_),
    .A2(_0654_));
 sg13g2_a22oi_1 _1247_ (.Y(_0115_),
    .B1(_0612_),
    .B2(_0656_),
    .A2(net271),
    .A1(_0392_));
 sg13g2_nor2_1 _1248_ (.A(net254),
    .B(_0539_),
    .Y(_0657_));
 sg13g2_a21oi_1 _1249_ (.A1(net254),
    .A2(_0627_),
    .Y(_0658_),
    .B1(_0657_));
 sg13g2_mux4_1 _1250_ (.S0(_0021_),
    .A0(_0630_),
    .A1(_0634_),
    .A2(_0539_),
    .A3(_0628_),
    .S1(net252),
    .X(_0659_));
 sg13g2_and2_1 _1251_ (.A(\mean_q[2] ),
    .B(_0659_),
    .X(_0660_));
 sg13g2_xor2_1 _1252_ (.B(_0659_),
    .A(\mean_q[2] ),
    .X(_0661_));
 sg13g2_a21oi_1 _1253_ (.A1(_0640_),
    .A2(_0654_),
    .Y(_0662_),
    .B1(_0653_));
 sg13g2_nand2b_1 _1254_ (.Y(_0663_),
    .B(_0661_),
    .A_N(_0662_));
 sg13g2_xor2_1 _1255_ (.B(_0662_),
    .A(_0661_),
    .X(_0664_));
 sg13g2_o21ai_1 _1256_ (.B1(_0614_),
    .Y(_0665_),
    .A1(net303),
    .A2(_0664_));
 sg13g2_o21ai_1 _1257_ (.B1(_0665_),
    .Y(_0666_),
    .A1(net396),
    .A2(_0436_));
 sg13g2_inv_1 _1258_ (.Y(_0116_),
    .A(_0666_));
 sg13g2_a21oi_1 _1259_ (.A1(_0021_),
    .A2(_0648_),
    .Y(_0667_),
    .B1(_0657_));
 sg13g2_mux4_1 _1260_ (.S0(net251),
    .A0(_0644_),
    .A1(_0648_),
    .A2(_0650_),
    .A3(_0540_),
    .S1(_0367_),
    .X(_0668_));
 sg13g2_nor2_1 _1261_ (.A(_0391_),
    .B(_0668_),
    .Y(_0669_));
 sg13g2_nand2_1 _1262_ (.Y(_0670_),
    .A(_0391_),
    .B(_0668_));
 sg13g2_xnor2_1 _1263_ (.Y(_0671_),
    .A(net401),
    .B(_0668_));
 sg13g2_nor2b_1 _1264_ (.A(_0660_),
    .B_N(_0663_),
    .Y(_0672_));
 sg13g2_xnor2_1 _1265_ (.Y(_0673_),
    .A(_0671_),
    .B(_0672_));
 sg13g2_nand2b_1 _1266_ (.Y(_0674_),
    .B(_0673_),
    .A_N(net303));
 sg13g2_a22oi_1 _1267_ (.Y(_0117_),
    .B1(_0616_),
    .B2(_0674_),
    .A2(net271),
    .A1(_0391_));
 sg13g2_nand2_1 _1268_ (.Y(_0675_),
    .A(net251),
    .B(_0540_));
 sg13g2_mux2_1 _1269_ (.A0(_0632_),
    .A1(_0540_),
    .S(net251),
    .X(_0676_));
 sg13g2_or2_1 _1270_ (.X(_0677_),
    .B(_0676_),
    .A(_0390_));
 sg13g2_xnor2_1 _1271_ (.Y(_0678_),
    .A(_0390_),
    .B(_0676_));
 sg13g2_nand2_1 _1272_ (.Y(_0679_),
    .A(_0661_),
    .B(_0671_));
 sg13g2_a21oi_1 _1273_ (.A1(_0660_),
    .A2(_0670_),
    .Y(_0680_),
    .B1(_0669_));
 sg13g2_o21ai_1 _1274_ (.B1(_0680_),
    .Y(_0681_),
    .A1(_0662_),
    .A2(_0679_));
 sg13g2_nand2b_1 _1275_ (.Y(_0682_),
    .B(_0681_),
    .A_N(_0678_));
 sg13g2_nand2b_1 _1276_ (.Y(_0683_),
    .B(_0678_),
    .A_N(_0681_));
 sg13g2_nand3b_1 _1277_ (.B(_0682_),
    .C(_0683_),
    .Y(_0684_),
    .A_N(net11));
 sg13g2_a22oi_1 _1278_ (.Y(_0118_),
    .B1(_0618_),
    .B2(_0684_),
    .A2(net269),
    .A1(_0390_));
 sg13g2_o21ai_1 _1279_ (.B1(_0675_),
    .Y(_0685_),
    .A1(net251),
    .A2(_0651_));
 sg13g2_nand2_1 _1280_ (.Y(_0686_),
    .A(_0389_),
    .B(_0685_));
 sg13g2_xnor2_1 _1281_ (.Y(_0687_),
    .A(_0389_),
    .B(_0685_));
 sg13g2_nand2_1 _1282_ (.Y(_0688_),
    .A(_0677_),
    .B(_0682_));
 sg13g2_xnor2_1 _1283_ (.Y(_0689_),
    .A(_0687_),
    .B(_0688_));
 sg13g2_nand2b_1 _1284_ (.Y(_0690_),
    .B(_0689_),
    .A_N(net304));
 sg13g2_a22oi_1 _1285_ (.Y(_0119_),
    .B1(_0620_),
    .B2(_0690_),
    .A2(net269),
    .A1(_0389_));
 sg13g2_nor2_1 _1286_ (.A(_0678_),
    .B(_0687_),
    .Y(_0691_));
 sg13g2_o21ai_1 _1287_ (.B1(_0677_),
    .Y(_0692_),
    .A1(_0389_),
    .A2(_0685_));
 sg13g2_a22oi_1 _1288_ (.Y(_0693_),
    .B1(_0692_),
    .B2(_0686_),
    .A2(_0691_),
    .A1(_0681_));
 sg13g2_nor2_1 _1289_ (.A(net251),
    .B(_0658_),
    .Y(_0694_));
 sg13g2_a21oi_1 _1290_ (.A1(net251),
    .A2(_0540_),
    .Y(_0695_),
    .B1(_0694_));
 sg13g2_nand2_1 _1291_ (.Y(_0696_),
    .A(\mean_q[6] ),
    .B(_0695_));
 sg13g2_xnor2_1 _1292_ (.Y(_0697_),
    .A(net398),
    .B(_0695_));
 sg13g2_a21oi_1 _1293_ (.A1(_0693_),
    .A2(_0697_),
    .Y(_0698_),
    .B1(net304));
 sg13g2_o21ai_1 _1294_ (.B1(_0698_),
    .Y(_0699_),
    .A1(_0693_),
    .A2(_0697_));
 sg13g2_a22oi_1 _1295_ (.Y(_0120_),
    .B1(_0622_),
    .B2(_0699_),
    .A2(net266),
    .A1(_0388_));
 sg13g2_o21ai_1 _1296_ (.B1(_0696_),
    .Y(_0700_),
    .A1(_0693_),
    .A2(_0697_));
 sg13g2_o21ai_1 _1297_ (.B1(_0675_),
    .Y(_0701_),
    .A1(net251),
    .A2(_0667_));
 sg13g2_xnor2_1 _1298_ (.Y(_0702_),
    .A(net385),
    .B(_0701_));
 sg13g2_a21oi_1 _1299_ (.A1(_0700_),
    .A2(_0702_),
    .Y(_0703_),
    .B1(net304));
 sg13g2_o21ai_1 _1300_ (.B1(_0703_),
    .Y(_0704_),
    .A1(_0700_),
    .A2(_0702_));
 sg13g2_a22oi_1 _1301_ (.Y(_0121_),
    .B1(_0624_),
    .B2(_0704_),
    .A2(net265),
    .A1(_0387_));
 sg13g2_nand2b_1 _1302_ (.Y(_0705_),
    .B(_0551_),
    .A_N(_0476_));
 sg13g2_and2_1 _1303_ (.A(_0464_),
    .B(_0544_),
    .X(_0706_));
 sg13g2_nor2_1 _1304_ (.A(_0562_),
    .B(_0706_),
    .Y(_0707_));
 sg13g2_nor2b_1 _1305_ (.A(_0707_),
    .B_N(_0480_),
    .Y(_0708_));
 sg13g2_nand2_1 _1306_ (.Y(_0709_),
    .A(_0527_),
    .B(_0706_));
 sg13g2_o21ai_1 _1307_ (.B1(_0709_),
    .Y(_0710_),
    .A1(_0482_),
    .A2(_0557_));
 sg13g2_a22oi_1 _1308_ (.Y(_0711_),
    .B1(_0569_),
    .B2(_0489_),
    .A2(_0557_),
    .A1(_0482_));
 sg13g2_o21ai_1 _1309_ (.B1(_0711_),
    .Y(_0712_),
    .A1(_0708_),
    .A2(_0710_));
 sg13g2_nand2_1 _1310_ (.Y(_0713_),
    .A(_0501_),
    .B(_0583_));
 sg13g2_a22oi_1 _1311_ (.Y(_0714_),
    .B1(_0583_),
    .B2(_0501_),
    .A2(_0574_),
    .A1(_0495_));
 sg13g2_o21ai_1 _1312_ (.B1(_0713_),
    .Y(_0715_),
    .A1(_0496_),
    .A2(_0573_));
 sg13g2_nand2b_1 _1313_ (.Y(_0716_),
    .B(_0573_),
    .A_N(_0495_));
 sg13g2_nand2_1 _1314_ (.Y(_0717_),
    .A(_0490_),
    .B(_0568_));
 sg13g2_nand2b_1 _1315_ (.Y(_0718_),
    .B(_0582_),
    .A_N(_0501_));
 sg13g2_and4_1 _1316_ (.A(_0714_),
    .B(_0716_),
    .C(_0717_),
    .D(_0718_),
    .X(_0719_));
 sg13g2_nor2_1 _1317_ (.A(_0507_),
    .B(_0587_),
    .Y(_0720_));
 sg13g2_a221oi_1 _1318_ (.B2(_0712_),
    .C1(_0720_),
    .B1(_0719_),
    .A1(_0715_),
    .Y(_0721_),
    .A2(_0718_));
 sg13g2_a22oi_1 _1319_ (.Y(_0722_),
    .B1(_0587_),
    .B2(_0507_),
    .A2(_0552_),
    .A1(_0476_));
 sg13g2_inv_1 _1320_ (.Y(_0723_),
    .A(_0722_));
 sg13g2_o21ai_1 _1321_ (.B1(_0705_),
    .Y(_0724_),
    .A1(_0721_),
    .A2(_0723_));
 sg13g2_nand2b_1 _1322_ (.Y(_0725_),
    .B(_0463_),
    .A_N(_0724_));
 sg13g2_nor2_2 _1323_ (.A(\reg_mode[1] ),
    .B(net249),
    .Y(_0726_));
 sg13g2_inv_1 _1324_ (.Y(_0727_),
    .A(_0726_));
 sg13g2_a21oi_1 _1325_ (.A1(_0544_),
    .A2(_0724_),
    .Y(_0728_),
    .B1(_0727_));
 sg13g2_nand2_1 _1326_ (.Y(_0729_),
    .A(net2),
    .B(net249));
 sg13g2_a21oi_1 _1327_ (.A1(_0725_),
    .A2(_0728_),
    .Y(_0730_),
    .B1(net265));
 sg13g2_a22oi_1 _1328_ (.Y(_0122_),
    .B1(_0729_),
    .B2(_0730_),
    .A2(net267),
    .A1(_0412_));
 sg13g2_nor2_1 _1329_ (.A(net218),
    .B(_0436_),
    .Y(_0731_));
 sg13g2_and2_1 _1330_ (.A(_0562_),
    .B(_0724_),
    .X(_0732_));
 sg13g2_o21ai_1 _1331_ (.B1(_0726_),
    .Y(_0733_),
    .A1(_0480_),
    .A2(_0724_));
 sg13g2_a21oi_1 _1332_ (.A1(net3),
    .A2(net249),
    .Y(_0734_),
    .B1(net271));
 sg13g2_o21ai_1 _1333_ (.B1(_0734_),
    .Y(_0735_),
    .A1(_0732_),
    .A2(_0733_));
 sg13g2_nor2b_1 _1334_ (.A(_0731_),
    .B_N(_0735_),
    .Y(_0123_));
 sg13g2_mux2_1 _1335_ (.A0(_0483_),
    .A1(_0557_),
    .S(_0724_),
    .X(_0736_));
 sg13g2_a221oi_1 _1336_ (.B2(_0736_),
    .C1(net267),
    .B1(_0726_),
    .A1(net4),
    .Y(_0737_),
    .A2(net249));
 sg13g2_a21oi_1 _1337_ (.A1(_0413_),
    .A2(net267),
    .Y(_0124_),
    .B1(_0737_));
 sg13g2_mux2_1 _1338_ (.A0(_0490_),
    .A1(_0569_),
    .S(_0724_),
    .X(_0738_));
 sg13g2_nand2_1 _1339_ (.Y(_0739_),
    .A(net5),
    .B(net249));
 sg13g2_a21oi_1 _1340_ (.A1(_0726_),
    .A2(_0738_),
    .Y(_0740_),
    .B1(net265));
 sg13g2_a22oi_1 _1341_ (.Y(_0125_),
    .B1(_0739_),
    .B2(_0740_),
    .A2(net267),
    .A1(_0414_));
 sg13g2_nand2b_1 _1342_ (.Y(_0741_),
    .B(_0726_),
    .A_N(_0512_));
 sg13g2_a21oi_1 _1343_ (.A1(net6),
    .A2(net249),
    .Y(_0742_),
    .B1(net268));
 sg13g2_a22oi_1 _1344_ (.Y(_0126_),
    .B1(_0741_),
    .B2(_0742_),
    .A2(net268),
    .A1(_0415_));
 sg13g2_nand2b_1 _1345_ (.Y(_0743_),
    .B(_0726_),
    .A_N(_0592_));
 sg13g2_a21oi_1 _1346_ (.A1(net7),
    .A2(net250),
    .Y(_0744_),
    .B1(net268));
 sg13g2_a22oi_1 _1347_ (.Y(_0127_),
    .B1(_0743_),
    .B2(_0744_),
    .A2(net268),
    .A1(_0416_));
 sg13g2_nand2b_1 _1348_ (.Y(_0745_),
    .B(_0726_),
    .A_N(_0594_));
 sg13g2_a21oi_1 _1349_ (.A1(net8),
    .A2(net250),
    .Y(_0746_),
    .B1(net268));
 sg13g2_a22oi_1 _1350_ (.Y(_0128_),
    .B1(_0745_),
    .B2(_0746_),
    .A2(net268),
    .A1(_0417_));
 sg13g2_a21o_1 _1351_ (.A2(_0591_),
    .A1(_0512_),
    .B1(_0727_),
    .X(_0747_));
 sg13g2_nor2_1 _1352_ (.A(net260),
    .B(_0399_),
    .Y(_0252_));
 sg13g2_a22oi_1 _1353_ (.Y(_0253_),
    .B1(\reg_thresh[0] ),
    .B2(_0371_),
    .A2(\reg_thresh[1] ),
    .A1(_0374_));
 sg13g2_a221oi_1 _1354_ (.B2(\pixel_q[1] ),
    .C1(_0253_),
    .B1(_0404_),
    .A1(\pixel_q[2] ),
    .Y(_0254_),
    .A2(_0403_));
 sg13g2_a221oi_1 _1355_ (.B2(_0384_),
    .C1(_0254_),
    .B1(\reg_thresh[2] ),
    .A1(_0382_),
    .Y(_0255_),
    .A2(\reg_thresh[3] ));
 sg13g2_a221oi_1 _1356_ (.B2(\pixel_q[3] ),
    .C1(_0255_),
    .B1(_0402_),
    .A1(\pixel_q[4] ),
    .Y(_0256_),
    .A2(_0401_));
 sg13g2_a221oi_1 _1357_ (.B2(_0380_),
    .C1(_0256_),
    .B1(\reg_thresh[4] ),
    .A1(_0378_),
    .Y(_0257_),
    .A2(\reg_thresh[5] ));
 sg13g2_a21oi_1 _1358_ (.A1(\pixel_q[5] ),
    .A2(_0400_),
    .Y(_0258_),
    .B1(_0257_));
 sg13g2_a22oi_1 _1359_ (.Y(_0259_),
    .B1(net260),
    .B2(_0399_),
    .A2(\pixel_q[7] ),
    .A1(_0015_));
 sg13g2_o21ai_1 _1360_ (.B1(_0259_),
    .Y(_0260_),
    .A1(_0252_),
    .A2(_0258_));
 sg13g2_nor2_1 _1361_ (.A(_0015_),
    .B(\pixel_q[7] ),
    .Y(_0261_));
 sg13g2_nor3_1 _1362_ (.A(_0398_),
    .B(net249),
    .C(_0261_),
    .Y(_0262_));
 sg13g2_a221oi_1 _1363_ (.B2(_0262_),
    .C1(net266),
    .B1(_0260_),
    .A1(net9),
    .Y(_0263_),
    .A2(net249));
 sg13g2_a22oi_1 _1364_ (.Y(_0129_),
    .B1(_0747_),
    .B2(_0263_),
    .A2(net266),
    .A1(_0418_));
 sg13g2_and4_1 _1365_ (.A(_0013_),
    .B(spi_cmd_wr),
    .C(net247),
    .D(_0432_),
    .X(_0264_));
 sg13g2_xor2_1 _1366_ (.B(net244),
    .A(spi_wr_toggle),
    .X(_0130_));
 sg13g2_mux2_1 _1367_ (.A0(\spi_wr_addr[0] ),
    .A1(\spi_cmd_addr[0] ),
    .S(net244),
    .X(_0131_));
 sg13g2_mux2_1 _1368_ (.A0(\spi_wr_addr[1] ),
    .A1(\spi_cmd_addr[1] ),
    .S(net244),
    .X(_0132_));
 sg13g2_mux2_1 _1369_ (.A0(\spi_wr_addr[2] ),
    .A1(\spi_cmd_addr[2] ),
    .S(net244),
    .X(_0133_));
 sg13g2_mux2_1 _1370_ (.A0(\spi_wr_data[0] ),
    .A1(net13),
    .S(net244),
    .X(_0134_));
 sg13g2_mux2_1 _1371_ (.A0(\spi_wr_data[1] ),
    .A1(\spi_shift_in[0] ),
    .S(net243),
    .X(_0135_));
 sg13g2_mux2_1 _1372_ (.A0(\spi_wr_data[2] ),
    .A1(\spi_shift_in[1] ),
    .S(net244),
    .X(_0136_));
 sg13g2_mux2_1 _1373_ (.A0(\spi_wr_data[3] ),
    .A1(\spi_shift_in[2] ),
    .S(net244),
    .X(_0137_));
 sg13g2_nor2_1 _1374_ (.A(\spi_wr_data[4] ),
    .B(net243),
    .Y(_0265_));
 sg13g2_a21oi_1 _1375_ (.A1(_0395_),
    .A2(net243),
    .Y(_0138_),
    .B1(_0265_));
 sg13g2_nor2_1 _1376_ (.A(\spi_wr_data[5] ),
    .B(net243),
    .Y(_0266_));
 sg13g2_a21oi_1 _1377_ (.A1(_0396_),
    .A2(net243),
    .Y(_0139_),
    .B1(_0266_));
 sg13g2_nor2_1 _1378_ (.A(\spi_wr_data[6] ),
    .B(net243),
    .Y(_0267_));
 sg13g2_a21oi_1 _1379_ (.A1(_0394_),
    .A2(net243),
    .Y(_0140_),
    .B1(_0267_));
 sg13g2_mux2_1 _1380_ (.A0(\spi_wr_data[7] ),
    .A1(\spi_shift_in[6] ),
    .S(net243),
    .X(_0141_));
 sg13g2_mux2_1 _1381_ (.A0(net13),
    .A1(\spi_shift_in[0] ),
    .S(net302),
    .X(_0142_));
 sg13g2_a22oi_1 _1382_ (.Y(_0268_),
    .B1(net248),
    .B2(\spi_shift_in[0] ),
    .A2(\spi_shift_in[1] ),
    .A1(net12));
 sg13g2_inv_1 _1383_ (.Y(_0143_),
    .A(_0268_));
 sg13g2_a22oi_1 _1384_ (.Y(_0269_),
    .B1(net248),
    .B2(\spi_shift_in[1] ),
    .A2(\spi_shift_in[2] ),
    .A1(net12));
 sg13g2_inv_1 _1385_ (.Y(_0144_),
    .A(_0269_));
 sg13g2_a22oi_1 _1386_ (.Y(_0270_),
    .B1(\spi_shift_in[2] ),
    .B2(net248),
    .A2(\spi_shift_in[3] ),
    .A1(net302));
 sg13g2_inv_1 _1387_ (.Y(_0145_),
    .A(_0270_));
 sg13g2_nand2_1 _1388_ (.Y(_0271_),
    .A(\spi_shift_in[3] ),
    .B(net248));
 sg13g2_a22oi_1 _1389_ (.Y(_0272_),
    .B1(net247),
    .B2(\spi_shift_in[3] ),
    .A2(\spi_shift_in[4] ),
    .A1(net302));
 sg13g2_inv_1 _1390_ (.Y(_0146_),
    .A(_0272_));
 sg13g2_nand2_1 _1391_ (.Y(_0273_),
    .A(\spi_shift_in[4] ),
    .B(net247));
 sg13g2_a22oi_1 _1392_ (.Y(_0274_),
    .B1(\spi_shift_in[4] ),
    .B2(net247),
    .A2(net259),
    .A1(net302));
 sg13g2_inv_1 _1393_ (.Y(_0147_),
    .A(_0274_));
 sg13g2_nand2_1 _1394_ (.Y(_0275_),
    .A(net259),
    .B(net248));
 sg13g2_a22oi_1 _1395_ (.Y(_0276_),
    .B1(net259),
    .B2(net247),
    .A2(\spi_shift_in[6] ),
    .A1(net302));
 sg13g2_inv_1 _1396_ (.Y(_0148_),
    .A(_0276_));
 sg13g2_o21ai_1 _1397_ (.B1(_0013_),
    .Y(_0277_),
    .A1(\spi_bitcnt[3] ),
    .A2(_0429_));
 sg13g2_a21oi_1 _1398_ (.A1(_0433_),
    .A2(_0277_),
    .Y(_0149_),
    .B1(_0427_));
 sg13g2_nor2b_1 _1399_ (.A(spi_cmd_wr),
    .B_N(_0433_),
    .Y(_0278_));
 sg13g2_nor3_1 _1400_ (.A(_0427_),
    .B(_0434_),
    .C(_0278_),
    .Y(_0150_));
 sg13g2_and2_1 _1401_ (.A(net248),
    .B(_0433_),
    .X(_0279_));
 sg13g2_nand2_1 _1402_ (.Y(_0280_),
    .A(\spi_cmd_addr[0] ),
    .B(_0279_));
 sg13g2_o21ai_1 _1403_ (.B1(_0280_),
    .Y(_0151_),
    .A1(_0433_),
    .A2(_0271_));
 sg13g2_nand2_1 _1404_ (.Y(_0281_),
    .A(\spi_cmd_addr[1] ),
    .B(_0279_));
 sg13g2_o21ai_1 _1405_ (.B1(_0281_),
    .Y(_0152_),
    .A1(_0433_),
    .A2(_0273_));
 sg13g2_nand2_1 _1406_ (.Y(_0282_),
    .A(\spi_cmd_addr[2] ),
    .B(_0279_));
 sg13g2_o21ai_1 _1407_ (.B1(_0282_),
    .Y(_0153_),
    .A1(_0433_),
    .A2(_0275_));
 sg13g2_nand2_1 _1408_ (.Y(_0283_),
    .A(\spi_shift_out_load[0] ),
    .B(net237));
 sg13g2_nor2_2 _1409_ (.A(\spi_shift_in[3] ),
    .B(\spi_shift_in[4] ),
    .Y(_0284_));
 sg13g2_nor3_2 _1410_ (.A(net259),
    .B(\spi_shift_in[3] ),
    .C(\spi_shift_in[4] ),
    .Y(_0285_));
 sg13g2_nand2_2 _1411_ (.Y(_0286_),
    .A(_0394_),
    .B(net246));
 sg13g2_nor3_2 _1412_ (.A(net259),
    .B(\spi_shift_in[3] ),
    .C(_0396_),
    .Y(_0287_));
 sg13g2_nor3_2 _1413_ (.A(_0394_),
    .B(_0395_),
    .C(_0396_),
    .Y(_0288_));
 sg13g2_nor3_2 _1414_ (.A(net259),
    .B(_0395_),
    .C(_0396_),
    .Y(_0289_));
 sg13g2_a22oi_1 _1415_ (.Y(_0290_),
    .B1(_0289_),
    .B2(\spi_rd_bus_ff2[24] ),
    .A2(_0288_),
    .A1(\spi_rd_bus_ff2[56] ));
 sg13g2_nor3_2 _1416_ (.A(_0394_),
    .B(\spi_shift_in[3] ),
    .C(_0396_),
    .Y(_0291_));
 sg13g2_nor3_2 _1417_ (.A(net259),
    .B(_0395_),
    .C(\spi_shift_in[4] ),
    .Y(_0292_));
 sg13g2_a221oi_1 _1418_ (.B2(\spi_rd_bus_ff2[48] ),
    .C1(_0285_),
    .B1(_0291_),
    .A1(\spi_rd_bus_ff2[32] ),
    .Y(_0293_),
    .A2(net246));
 sg13g2_a22oi_1 _1419_ (.Y(_0294_),
    .B1(_0292_),
    .B2(\spi_rd_bus_ff2[8] ),
    .A2(_0287_),
    .A1(\spi_rd_bus_ff2[16] ));
 sg13g2_and3_1 _1420_ (.X(_0295_),
    .A(_0290_),
    .B(_0293_),
    .C(_0294_));
 sg13g2_o21ai_1 _1421_ (.B1(net236),
    .Y(_0296_),
    .A1(\spi_rd_bus_ff2[0] ),
    .A2(net245));
 sg13g2_o21ai_1 _1422_ (.B1(_0283_),
    .Y(_0154_),
    .A1(_0295_),
    .A2(_0296_));
 sg13g2_nand2_1 _1423_ (.Y(_0297_),
    .A(\spi_shift_out_load[1] ),
    .B(net237));
 sg13g2_nand3_1 _1424_ (.B(\spi_rd_bus_ff2[33] ),
    .C(net246),
    .A(\spi_shift_in[5] ),
    .Y(_0298_));
 sg13g2_a22oi_1 _1425_ (.Y(_0299_),
    .B1(_0291_),
    .B2(\spi_rd_bus_ff2[49] ),
    .A2(_0288_),
    .A1(\spi_rd_bus_ff2[57] ));
 sg13g2_a22oi_1 _1426_ (.Y(_0300_),
    .B1(_0292_),
    .B2(\spi_rd_bus_ff2[9] ),
    .A2(_0287_),
    .A1(\spi_rd_bus_ff2[17] ));
 sg13g2_a21oi_1 _1427_ (.A1(\spi_rd_bus_ff2[25] ),
    .A2(_0289_),
    .Y(_0301_),
    .B1(_0285_));
 sg13g2_and4_1 _1428_ (.A(_0298_),
    .B(_0299_),
    .C(_0300_),
    .D(_0301_),
    .X(_0302_));
 sg13g2_o21ai_1 _1429_ (.B1(net236),
    .Y(_0303_),
    .A1(\spi_rd_bus_ff2[1] ),
    .A2(net245));
 sg13g2_o21ai_1 _1430_ (.B1(_0297_),
    .Y(_0155_),
    .A1(_0302_),
    .A2(_0303_));
 sg13g2_nand2_1 _1431_ (.Y(_0304_),
    .A(\spi_shift_out_load[2] ),
    .B(net237));
 sg13g2_a22oi_1 _1432_ (.Y(_0305_),
    .B1(_0291_),
    .B2(\spi_rd_bus_ff2[50] ),
    .A2(_0287_),
    .A1(\spi_rd_bus_ff2[18] ));
 sg13g2_a221oi_1 _1433_ (.B2(\spi_rd_bus_ff2[58] ),
    .C1(_0285_),
    .B1(_0288_),
    .A1(\spi_rd_bus_ff2[34] ),
    .Y(_0306_),
    .A2(_0284_));
 sg13g2_a22oi_1 _1434_ (.Y(_0307_),
    .B1(_0292_),
    .B2(\spi_rd_bus_ff2[10] ),
    .A2(_0289_),
    .A1(\spi_rd_bus_ff2[26] ));
 sg13g2_and3_1 _1435_ (.X(_0308_),
    .A(_0305_),
    .B(_0306_),
    .C(_0307_));
 sg13g2_o21ai_1 _1436_ (.B1(net236),
    .Y(_0309_),
    .A1(\spi_rd_bus_ff2[2] ),
    .A2(net245));
 sg13g2_o21ai_1 _1437_ (.B1(_0304_),
    .Y(_0156_),
    .A1(_0308_),
    .A2(_0309_));
 sg13g2_nand2_1 _1438_ (.Y(_0310_),
    .A(\spi_shift_out_load[3] ),
    .B(_0435_));
 sg13g2_nand2_1 _1439_ (.Y(_0311_),
    .A(\spi_rd_bus_ff2[19] ),
    .B(_0287_));
 sg13g2_a22oi_1 _1440_ (.Y(_0312_),
    .B1(_0288_),
    .B2(\spi_rd_bus_ff2[59] ),
    .A2(net246),
    .A1(\spi_rd_bus_ff2[35] ));
 sg13g2_nand3_1 _1441_ (.B(_0311_),
    .C(_0312_),
    .A(_0286_),
    .Y(_0313_));
 sg13g2_a221oi_1 _1442_ (.B2(\spi_rd_bus_ff2[11] ),
    .C1(_0313_),
    .B1(_0292_),
    .A1(\spi_rd_bus_ff2[51] ),
    .Y(_0314_),
    .A2(_0291_));
 sg13g2_o21ai_1 _1443_ (.B1(_0012_),
    .Y(_0315_),
    .A1(\spi_rd_bus_ff2[3] ),
    .A2(net245));
 sg13g2_o21ai_1 _1444_ (.B1(_0310_),
    .Y(_0157_),
    .A1(_0314_),
    .A2(_0315_));
 sg13g2_nand2_1 _1445_ (.Y(_0316_),
    .A(\spi_shift_out_load[4] ),
    .B(net237));
 sg13g2_nand2_1 _1446_ (.Y(_0317_),
    .A(\spi_rd_bus_ff2[20] ),
    .B(_0287_));
 sg13g2_nor3_2 _1447_ (.A(_0394_),
    .B(_0395_),
    .C(\spi_shift_in[4] ),
    .Y(_0318_));
 sg13g2_a22oi_1 _1448_ (.Y(_0319_),
    .B1(_0292_),
    .B2(\spi_rd_bus_ff2[12] ),
    .A2(_0288_),
    .A1(\spi_rd_bus_ff2[60] ));
 sg13g2_o21ai_1 _1449_ (.B1(net246),
    .Y(_0320_),
    .A1(_0394_),
    .A2(\spi_rd_bus_ff2[36] ));
 sg13g2_a22oi_1 _1450_ (.Y(_0321_),
    .B1(_0318_),
    .B2(\spi_rd_bus_ff2[44] ),
    .A2(_0291_),
    .A1(\spi_rd_bus_ff2[52] ));
 sg13g2_and4_1 _1451_ (.A(_0317_),
    .B(_0319_),
    .C(_0320_),
    .D(_0321_),
    .X(_0322_));
 sg13g2_o21ai_1 _1452_ (.B1(net236),
    .Y(_0323_),
    .A1(\spi_rd_bus_ff2[4] ),
    .A2(net245));
 sg13g2_o21ai_1 _1453_ (.B1(_0316_),
    .Y(_0158_),
    .A1(_0322_),
    .A2(_0323_));
 sg13g2_nand2_1 _1454_ (.Y(_0324_),
    .A(\spi_shift_out_load[5] ),
    .B(net237));
 sg13g2_nand3_1 _1455_ (.B(\spi_rd_bus_ff2[37] ),
    .C(net246),
    .A(\spi_shift_in[5] ),
    .Y(_0325_));
 sg13g2_a21oi_1 _1456_ (.A1(\spi_rd_bus_ff2[45] ),
    .A2(_0318_),
    .Y(_0326_),
    .B1(_0285_));
 sg13g2_a22oi_1 _1457_ (.Y(_0327_),
    .B1(_0291_),
    .B2(\spi_rd_bus_ff2[53] ),
    .A2(_0288_),
    .A1(\spi_rd_bus_ff2[61] ));
 sg13g2_a22oi_1 _1458_ (.Y(_0328_),
    .B1(_0292_),
    .B2(\spi_rd_bus_ff2[13] ),
    .A2(_0287_),
    .A1(\spi_rd_bus_ff2[21] ));
 sg13g2_and4_1 _1459_ (.A(_0325_),
    .B(_0326_),
    .C(_0327_),
    .D(_0328_),
    .X(_0329_));
 sg13g2_o21ai_1 _1460_ (.B1(net236),
    .Y(_0330_),
    .A1(\spi_rd_bus_ff2[5] ),
    .A2(net245));
 sg13g2_o21ai_1 _1461_ (.B1(_0324_),
    .Y(_0159_),
    .A1(_0329_),
    .A2(_0330_));
 sg13g2_nand2_1 _1462_ (.Y(_0331_),
    .A(\spi_shift_out_load[6] ),
    .B(net237));
 sg13g2_a22oi_1 _1463_ (.Y(_0332_),
    .B1(_0318_),
    .B2(\spi_rd_bus_ff2[46] ),
    .A2(_0287_),
    .A1(\spi_rd_bus_ff2[22] ));
 sg13g2_a221oi_1 _1464_ (.B2(\spi_rd_bus_ff2[54] ),
    .C1(_0285_),
    .B1(_0291_),
    .A1(\spi_rd_bus_ff2[38] ),
    .Y(_0333_),
    .A2(net246));
 sg13g2_a22oi_1 _1465_ (.Y(_0334_),
    .B1(_0292_),
    .B2(\spi_rd_bus_ff2[14] ),
    .A2(_0288_),
    .A1(\spi_rd_bus_ff2[62] ));
 sg13g2_and3_1 _1466_ (.X(_0335_),
    .A(_0332_),
    .B(_0333_),
    .C(_0334_));
 sg13g2_o21ai_1 _1467_ (.B1(net236),
    .Y(_0336_),
    .A1(\spi_rd_bus_ff2[6] ),
    .A2(net245));
 sg13g2_o21ai_1 _1468_ (.B1(_0331_),
    .Y(_0160_),
    .A1(_0335_),
    .A2(_0336_));
 sg13g2_nand2_1 _1469_ (.Y(_0337_),
    .A(\spi_shift_out_load[7] ),
    .B(net237));
 sg13g2_a22oi_1 _1470_ (.Y(_0338_),
    .B1(_0318_),
    .B2(\spi_rd_bus_ff2[47] ),
    .A2(_0292_),
    .A1(\spi_rd_bus_ff2[15] ));
 sg13g2_a221oi_1 _1471_ (.B2(\spi_rd_bus_ff2[55] ),
    .C1(_0285_),
    .B1(_0291_),
    .A1(\spi_rd_bus_ff2[39] ),
    .Y(_0339_),
    .A2(net246));
 sg13g2_a22oi_1 _1472_ (.Y(_0340_),
    .B1(_0288_),
    .B2(\spi_rd_bus_ff2[63] ),
    .A2(_0287_),
    .A1(\spi_rd_bus_ff2[23] ));
 sg13g2_and3_1 _1473_ (.X(_0341_),
    .A(_0338_),
    .B(_0339_),
    .C(_0340_));
 sg13g2_o21ai_1 _1474_ (.B1(net236),
    .Y(_0342_),
    .A1(\spi_rd_bus_ff2[7] ),
    .A2(net245));
 sg13g2_o21ai_1 _1475_ (.B1(_0337_),
    .Y(_0161_),
    .A1(_0341_),
    .A2(_0342_));
 sg13g2_xnor2_1 _1476_ (.Y(_0343_),
    .A(cfg_wr_toggle_ff2_d),
    .B(cfg_wr_toggle_ff2));
 sg13g2_nor3_1 _1477_ (.A(\cfg_wr_addr_ff2[0] ),
    .B(\cfg_wr_addr_ff2[1] ),
    .C(_0343_),
    .Y(_0344_));
 sg13g2_nor2_1 _1478_ (.A(\cfg_wr_addr_ff2[2] ),
    .B(_0343_),
    .Y(_0345_));
 sg13g2_nor2b_2 _1479_ (.A(\cfg_wr_addr_ff2[2] ),
    .B_N(_0344_),
    .Y(_0346_));
 sg13g2_mux2_1 _1480_ (.A0(net371),
    .A1(net176),
    .S(net241),
    .X(_0162_));
 sg13g2_mux2_1 _1481_ (.A0(net232),
    .A1(net171),
    .S(net242),
    .X(_0163_));
 sg13g2_nand2_1 _1482_ (.Y(_0347_),
    .A(net165),
    .B(net242));
 sg13g2_o21ai_1 _1483_ (.B1(_0347_),
    .Y(_0164_),
    .A1(_0403_),
    .A2(net242));
 sg13g2_nand2_1 _1484_ (.Y(_0348_),
    .A(net186),
    .B(net242));
 sg13g2_o21ai_1 _1485_ (.B1(_0348_),
    .Y(_0165_),
    .A1(_0402_),
    .A2(net242));
 sg13g2_nand2_1 _1486_ (.Y(_0349_),
    .A(net181),
    .B(net241));
 sg13g2_o21ai_1 _1487_ (.B1(net182),
    .Y(_0166_),
    .A1(_0401_),
    .A2(net241));
 sg13g2_mux2_1 _1488_ (.A0(\reg_thresh[5] ),
    .A1(net353),
    .S(net241),
    .X(_0167_));
 sg13g2_nand2_1 _1489_ (.Y(_0350_),
    .A(net173),
    .B(net241));
 sg13g2_o21ai_1 _1490_ (.B1(net174),
    .Y(_0168_),
    .A1(_0399_),
    .A2(net241));
 sg13g2_nor2_1 _1491_ (.A(_0015_),
    .B(net241),
    .Y(_0351_));
 sg13g2_a21oi_1 _1492_ (.A1(net152),
    .A2(net241),
    .Y(_0169_),
    .B1(_0351_));
 sg13g2_nand2_1 _1493_ (.Y(_0352_),
    .A(\cfg_wr_addr_ff2[0] ),
    .B(_0345_));
 sg13g2_nor2_2 _1494_ (.A(\cfg_wr_addr_ff2[1] ),
    .B(_0352_),
    .Y(_0353_));
 sg13g2_mux2_1 _1495_ (.A0(net363),
    .A1(net176),
    .S(net240),
    .X(_0170_));
 sg13g2_mux2_1 _1496_ (.A0(net357),
    .A1(net171),
    .S(_0353_),
    .X(_0171_));
 sg13g2_nor2_1 _1497_ (.A(net167),
    .B(net240),
    .Y(_0354_));
 sg13g2_a21oi_1 _1498_ (.A1(net165),
    .A2(net240),
    .Y(_0172_),
    .B1(net168));
 sg13g2_nor2_1 _1499_ (.A(_0017_),
    .B(_0353_),
    .Y(_0355_));
 sg13g2_a21oi_1 _1500_ (.A1(net186),
    .A2(_0353_),
    .Y(_0173_),
    .B1(_0355_));
 sg13g2_mux2_1 _1501_ (.A0(net383),
    .A1(net181),
    .S(net240),
    .X(_0174_));
 sg13g2_mux2_1 _1502_ (.A0(net369),
    .A1(net353),
    .S(net240),
    .X(_0175_));
 sg13g2_mux2_1 _1503_ (.A0(net365),
    .A1(net173),
    .S(net240),
    .X(_0176_));
 sg13g2_nand2_1 _1504_ (.Y(_0356_),
    .A(net152),
    .B(net240));
 sg13g2_o21ai_1 _1505_ (.B1(_0356_),
    .Y(_0177_),
    .A1(_0393_),
    .A2(net240));
 sg13g2_nand2_1 _1506_ (.Y(_0357_),
    .A(\cfg_wr_addr_ff2[1] ),
    .B(_0345_));
 sg13g2_nor2_1 _1507_ (.A(\cfg_wr_addr_ff2[0] ),
    .B(_0357_),
    .Y(_0358_));
 sg13g2_mux2_1 _1508_ (.A0(net373),
    .A1(net176),
    .S(net238),
    .X(_0178_));
 sg13g2_mux2_1 _1509_ (.A0(net361),
    .A1(net171),
    .S(net238),
    .X(_0179_));
 sg13g2_nor2_1 _1510_ (.A(_0018_),
    .B(net239),
    .Y(_0359_));
 sg13g2_a21oi_1 _1511_ (.A1(net165),
    .A2(net239),
    .Y(_0180_),
    .B1(_0359_));
 sg13g2_nor2_1 _1512_ (.A(net191),
    .B(net239),
    .Y(_0360_));
 sg13g2_a21oi_1 _1513_ (.A1(net186),
    .A2(net239),
    .Y(_0181_),
    .B1(net192));
 sg13g2_mux2_1 _1514_ (.A0(net377),
    .A1(net181),
    .S(net238),
    .X(_0182_));
 sg13g2_mux2_1 _1515_ (.A0(net355),
    .A1(net353),
    .S(net238),
    .X(_0183_));
 sg13g2_nand2_1 _1516_ (.Y(_0361_),
    .A(net173),
    .B(net238));
 sg13g2_o21ai_1 _1517_ (.B1(_0361_),
    .Y(_0184_),
    .A1(_0386_),
    .A2(net238));
 sg13g2_nand2_1 _1518_ (.Y(_0362_),
    .A(net152),
    .B(net238));
 sg13g2_o21ai_1 _1519_ (.B1(_0362_),
    .Y(_0185_),
    .A1(_0385_),
    .A2(net238));
 sg13g2_nand3_1 _1520_ (.B(\cfg_wr_addr_ff2[1] ),
    .C(_0345_),
    .A(\cfg_wr_addr_ff2[0] ),
    .Y(_0363_));
 sg13g2_nand2_1 _1521_ (.Y(_0364_),
    .A(net256),
    .B(_0363_));
 sg13g2_o21ai_1 _1522_ (.B1(_0364_),
    .Y(_0186_),
    .A1(net176),
    .A2(_0363_));
 sg13g2_nand2_1 _1523_ (.Y(_0365_),
    .A(net254),
    .B(_0363_));
 sg13g2_o21ai_1 _1524_ (.B1(_0365_),
    .Y(_0187_),
    .A1(net171),
    .A2(_0363_));
 sg13g2_mux2_1 _1525_ (.A0(net165),
    .A1(net253),
    .S(_0363_),
    .X(_0188_));
 sg13g2_and2_1 _1526_ (.A(net329),
    .B(\spi_rd_bus_ff1[0] ),
    .X(_0189_));
 sg13g2_and2_1 _1527_ (.A(net329),
    .B(\spi_rd_bus_ff1[1] ),
    .X(_0190_));
 sg13g2_and2_1 _1528_ (.A(net329),
    .B(\spi_rd_bus_ff1[2] ),
    .X(_0191_));
 sg13g2_and2_1 _1529_ (.A(net328),
    .B(\spi_rd_bus_ff1[3] ),
    .X(_0192_));
 sg13g2_and2_1 _1530_ (.A(net325),
    .B(\spi_rd_bus_ff1[4] ),
    .X(_0193_));
 sg13g2_and2_1 _1531_ (.A(net321),
    .B(\spi_rd_bus_ff1[5] ),
    .X(_0194_));
 sg13g2_and2_1 _1532_ (.A(net321),
    .B(\spi_rd_bus_ff1[6] ),
    .X(_0195_));
 sg13g2_and2_1 _1533_ (.A(net321),
    .B(\spi_rd_bus_ff1[7] ),
    .X(_0196_));
 sg13g2_and2_1 _1534_ (.A(net342),
    .B(\spi_rd_bus_ff1[8] ),
    .X(_0197_));
 sg13g2_and2_1 _1535_ (.A(net329),
    .B(\spi_rd_bus_ff1[9] ),
    .X(_0198_));
 sg13g2_and2_1 _1536_ (.A(net329),
    .B(\spi_rd_bus_ff1[10] ),
    .X(_0199_));
 sg13g2_and2_1 _1537_ (.A(net328),
    .B(\spi_rd_bus_ff1[11] ),
    .X(_0200_));
 sg13g2_and2_1 _1538_ (.A(net321),
    .B(\spi_rd_bus_ff1[12] ),
    .X(_0201_));
 sg13g2_and2_1 _1539_ (.A(net322),
    .B(\spi_rd_bus_ff1[13] ),
    .X(_0202_));
 sg13g2_and2_1 _1540_ (.A(net320),
    .B(\spi_rd_bus_ff1[14] ),
    .X(_0203_));
 sg13g2_and2_1 _1541_ (.A(net326),
    .B(\spi_rd_bus_ff1[15] ),
    .X(_0204_));
 sg13g2_and2_1 _1542_ (.A(net342),
    .B(\spi_rd_bus_ff1[16] ),
    .X(_0205_));
 sg13g2_and2_1 _1543_ (.A(net342),
    .B(\spi_rd_bus_ff1[17] ),
    .X(_0206_));
 sg13g2_and2_1 _1544_ (.A(net342),
    .B(\spi_rd_bus_ff1[18] ),
    .X(_0207_));
 sg13g2_and2_1 _1545_ (.A(net327),
    .B(\spi_rd_bus_ff1[19] ),
    .X(_0208_));
 sg13g2_and2_1 _1546_ (.A(net322),
    .B(\spi_rd_bus_ff1[20] ),
    .X(_0209_));
 sg13g2_and2_1 _1547_ (.A(net322),
    .B(\spi_rd_bus_ff1[21] ),
    .X(_0210_));
 sg13g2_and2_1 _1548_ (.A(net308),
    .B(\spi_rd_bus_ff1[22] ),
    .X(_0211_));
 sg13g2_and2_1 _1549_ (.A(net322),
    .B(\spi_rd_bus_ff1[23] ),
    .X(_0212_));
 sg13g2_and2_1 _1550_ (.A(net344),
    .B(\spi_rd_bus_ff1[24] ),
    .X(_0213_));
 sg13g2_and2_1 _1551_ (.A(net343),
    .B(\spi_rd_bus_ff1[25] ),
    .X(_0214_));
 sg13g2_and2_1 _1552_ (.A(net343),
    .B(\spi_rd_bus_ff1[26] ),
    .X(_0215_));
 sg13g2_and2_1 _1553_ (.A(net342),
    .B(\spi_rd_bus_ff1[32] ),
    .X(_0216_));
 sg13g2_and2_1 _1554_ (.A(net330),
    .B(\spi_rd_bus_ff1[33] ),
    .X(_0217_));
 sg13g2_and2_1 _1555_ (.A(net329),
    .B(\spi_rd_bus_ff1[34] ),
    .X(_0218_));
 sg13g2_and2_1 _1556_ (.A(net321),
    .B(\spi_rd_bus_ff1[35] ),
    .X(_0219_));
 sg13g2_and2_1 _1557_ (.A(net320),
    .B(\spi_rd_bus_ff1[36] ),
    .X(_0220_));
 sg13g2_and2_1 _1558_ (.A(net320),
    .B(\spi_rd_bus_ff1[37] ),
    .X(_0221_));
 sg13g2_and2_1 _1559_ (.A(net320),
    .B(\spi_rd_bus_ff1[38] ),
    .X(_0222_));
 sg13g2_and2_1 _1560_ (.A(net322),
    .B(\spi_rd_bus_ff1[39] ),
    .X(_0223_));
 sg13g2_and2_1 _1561_ (.A(net326),
    .B(\spi_rd_bus_ff1[44] ),
    .X(_0224_));
 sg13g2_and2_1 _1562_ (.A(net316),
    .B(\spi_rd_bus_ff1[45] ),
    .X(_0225_));
 sg13g2_and2_1 _1563_ (.A(net335),
    .B(\spi_rd_bus_ff1[46] ),
    .X(_0226_));
 sg13g2_and2_1 _1564_ (.A(net317),
    .B(\spi_rd_bus_ff1[47] ),
    .X(_0227_));
 sg13g2_and2_1 _1565_ (.A(net349),
    .B(\spi_rd_bus_ff1[48] ),
    .X(_0228_));
 sg13g2_and2_1 _1566_ (.A(net349),
    .B(\spi_rd_bus_ff1[49] ),
    .X(_0229_));
 sg13g2_and2_1 _1567_ (.A(net347),
    .B(\spi_rd_bus_ff1[50] ),
    .X(_0230_));
 sg13g2_and2_1 _1568_ (.A(net342),
    .B(\spi_rd_bus_ff1[51] ),
    .X(_0231_));
 sg13g2_and2_1 _1569_ (.A(net327),
    .B(\spi_rd_bus_ff1[52] ),
    .X(_0232_));
 sg13g2_and2_1 _1570_ (.A(net344),
    .B(\spi_rd_bus_ff1[53] ),
    .X(_0233_));
 sg13g2_and2_1 _1571_ (.A(net326),
    .B(\spi_rd_bus_ff1[54] ),
    .X(_0234_));
 sg13g2_and2_1 _1572_ (.A(net326),
    .B(\spi_rd_bus_ff1[55] ),
    .X(_0235_));
 sg13g2_and2_1 _1573_ (.A(net343),
    .B(\spi_rd_bus_ff1[56] ),
    .X(_0236_));
 sg13g2_and2_1 _1574_ (.A(net342),
    .B(\spi_rd_bus_ff1[57] ),
    .X(_0237_));
 sg13g2_and2_1 _1575_ (.A(net347),
    .B(\spi_rd_bus_ff1[58] ),
    .X(_0238_));
 sg13g2_and2_1 _1576_ (.A(net328),
    .B(\spi_rd_bus_ff1[59] ),
    .X(_0239_));
 sg13g2_and2_1 _1577_ (.A(net321),
    .B(\spi_rd_bus_ff1[60] ),
    .X(_0240_));
 sg13g2_and2_1 _1578_ (.A(net328),
    .B(\spi_rd_bus_ff1[61] ),
    .X(_0241_));
 sg13g2_and2_1 _1579_ (.A(net322),
    .B(\spi_rd_bus_ff1[62] ),
    .X(_0242_));
 sg13g2_and2_1 _1580_ (.A(net326),
    .B(\spi_rd_bus_ff1[63] ),
    .X(_0243_));
 sg13g2_nand2_2 _1581_ (.Y(_0366_),
    .A(\cfg_wr_addr_ff2[2] ),
    .B(_0344_));
 sg13g2_mux2_1 _1582_ (.A0(net176),
    .A1(net250),
    .S(_0366_),
    .X(_0244_));
 sg13g2_mux2_1 _1583_ (.A0(net171),
    .A1(net367),
    .S(_0366_),
    .X(_0245_));
 sg13g2_mux2_1 _1584_ (.A0(net165),
    .A1(net200),
    .S(_0366_),
    .X(_0246_));
 sg13g2_mux2_1 _1585_ (.A0(net186),
    .A1(net198),
    .S(_0366_),
    .X(_0247_));
 sg13g2_mux2_1 _1586_ (.A0(net181),
    .A1(net196),
    .S(_0366_),
    .X(_0248_));
 sg13g2_mux2_1 _1587_ (.A0(\cfg_wr_data_ff2[5] ),
    .A1(net184),
    .S(_0366_),
    .X(_0249_));
 sg13g2_mux2_1 _1588_ (.A0(net173),
    .A1(net194),
    .S(_0366_),
    .X(_0250_));
 sg13g2_mux2_1 _1589_ (.A0(net152),
    .A1(net189),
    .S(_0366_),
    .X(_0251_));
 sg13g2_inv_1 _1590_ (.Y(_0023_),
    .A(net286));
 sg13g2_inv_1 _1591_ (.Y(_0024_),
    .A(net287));
 sg13g2_inv_1 _1592_ (.Y(_0025_),
    .A(net286));
 sg13g2_inv_1 _1593_ (.Y(_0026_),
    .A(net286));
 sg13g2_inv_1 _1594_ (.Y(_0027_),
    .A(net286));
 sg13g2_inv_1 _1595_ (.Y(_0028_),
    .A(net286));
 sg13g2_inv_1 _1596_ (.Y(_0029_),
    .A(net301));
 sg13g2_dfrbpq_1 _1597_ (.RESET_B(net323),
    .D(_0005_),
    .Q(\spi_shift_out[1] ),
    .CLK(_0022_));
 sg13g2_dfrbpq_1 _1598_ (.RESET_B(net323),
    .D(_0006_),
    .Q(\spi_shift_out[2] ),
    .CLK(_0023_));
 sg13g2_dfrbpq_1 _1599_ (.RESET_B(net324),
    .D(_0007_),
    .Q(\spi_shift_out[3] ),
    .CLK(_0024_));
 sg13g2_dfrbpq_1 _1600_ (.RESET_B(net323),
    .D(_0008_),
    .Q(\spi_shift_out[4] ),
    .CLK(_0025_));
 sg13g2_dfrbpq_1 _1601_ (.RESET_B(net323),
    .D(_0009_),
    .Q(\spi_shift_out[5] ),
    .CLK(_0026_));
 sg13g2_dfrbpq_1 _1602_ (.RESET_B(net323),
    .D(_0010_),
    .Q(\spi_shift_out[6] ),
    .CLK(_0027_));
 sg13g2_dfrbpq_1 _1603_ (.RESET_B(net323),
    .D(_0011_),
    .Q(\spi_shift_out[7] ),
    .CLK(_0028_));
 sg13g2_dfrbpq_1 _1604_ (.RESET_B(net316),
    .D(_0031_),
    .Q(\reg_status[4] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _1605_ (.RESET_B(net338),
    .D(_0032_),
    .Q(\reg_status[5] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _1606_ (.RESET_B(net338),
    .D(_0033_),
    .Q(\reg_status[6] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_1 _1607_ (.RESET_B(net312),
    .D(_0034_),
    .Q(\reg_status[7] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_1 _1608_ (.RESET_B(net82),
    .D(_0035_),
    .Q(\spi_rd_bus_ff1[0] ),
    .CLK(net293));
 sg13g2_dfrbpq_1 _1609_ (.RESET_B(net81),
    .D(_0036_),
    .Q(\spi_rd_bus_ff1[1] ),
    .CLK(net293));
 sg13g2_dfrbpq_1 _1610_ (.RESET_B(net80),
    .D(_0037_),
    .Q(\spi_rd_bus_ff1[2] ),
    .CLK(net296));
 sg13g2_dfrbpq_1 _1611_ (.RESET_B(net79),
    .D(_0038_),
    .Q(\spi_rd_bus_ff1[3] ),
    .CLK(net291));
 sg13g2_dfrbpq_1 _1612_ (.RESET_B(net78),
    .D(_0039_),
    .Q(\spi_rd_bus_ff1[4] ),
    .CLK(net282));
 sg13g2_dfrbpq_1 _1613_ (.RESET_B(net77),
    .D(_0040_),
    .Q(\spi_rd_bus_ff1[5] ),
    .CLK(net282));
 sg13g2_dfrbpq_1 _1614_ (.RESET_B(net76),
    .D(_0041_),
    .Q(\spi_rd_bus_ff1[6] ),
    .CLK(net282));
 sg13g2_dfrbpq_1 _1615_ (.RESET_B(net75),
    .D(_0042_),
    .Q(\spi_rd_bus_ff1[7] ),
    .CLK(net282));
 sg13g2_dfrbpq_1 _1616_ (.RESET_B(net74),
    .D(_0043_),
    .Q(\spi_rd_bus_ff1[8] ),
    .CLK(net299));
 sg13g2_dfrbpq_1 _1617_ (.RESET_B(net73),
    .D(_0044_),
    .Q(\spi_rd_bus_ff1[9] ),
    .CLK(net299));
 sg13g2_dfrbpq_1 _1618_ (.RESET_B(net72),
    .D(_0045_),
    .Q(\spi_rd_bus_ff1[10] ),
    .CLK(net290));
 sg13g2_dfrbpq_1 _1619_ (.RESET_B(net71),
    .D(_0046_),
    .Q(\spi_rd_bus_ff1[11] ),
    .CLK(net290));
 sg13g2_dfrbpq_1 _1620_ (.RESET_B(net70),
    .D(_0047_),
    .Q(\spi_rd_bus_ff1[12] ),
    .CLK(net282));
 sg13g2_dfrbpq_1 _1621_ (.RESET_B(net69),
    .D(_0048_),
    .Q(\spi_rd_bus_ff1[13] ),
    .CLK(net283));
 sg13g2_dfrbpq_1 _1622_ (.RESET_B(net68),
    .D(_0049_),
    .Q(\spi_rd_bus_ff1[14] ),
    .CLK(net276));
 sg13g2_dfrbpq_1 _1623_ (.RESET_B(net67),
    .D(_0050_),
    .Q(\spi_rd_bus_ff1[15] ),
    .CLK(net280));
 sg13g2_dfrbpq_1 _1624_ (.RESET_B(net66),
    .D(_0051_),
    .Q(\spi_rd_bus_ff1[16] ),
    .CLK(net299));
 sg13g2_dfrbpq_1 _1625_ (.RESET_B(net65),
    .D(_0052_),
    .Q(\spi_rd_bus_ff1[17] ),
    .CLK(net299));
 sg13g2_dfrbpq_1 _1626_ (.RESET_B(net64),
    .D(_0053_),
    .Q(\spi_rd_bus_ff1[18] ),
    .CLK(net299));
 sg13g2_dfrbpq_1 _1627_ (.RESET_B(net63),
    .D(_0054_),
    .Q(\spi_rd_bus_ff1[19] ),
    .CLK(net290));
 sg13g2_dfrbpq_1 _1628_ (.RESET_B(net62),
    .D(_0055_),
    .Q(\spi_rd_bus_ff1[20] ),
    .CLK(net283));
 sg13g2_dfrbpq_1 _1629_ (.RESET_B(net61),
    .D(_0056_),
    .Q(\spi_rd_bus_ff1[21] ),
    .CLK(net283));
 sg13g2_dfrbpq_1 _1630_ (.RESET_B(net60),
    .D(_0057_),
    .Q(\spi_rd_bus_ff1[22] ),
    .CLK(net281));
 sg13g2_dfrbpq_1 _1631_ (.RESET_B(net59),
    .D(_0058_),
    .Q(\spi_rd_bus_ff1[23] ),
    .CLK(net281));
 sg13g2_dfrbpq_1 _1632_ (.RESET_B(net58),
    .D(_0059_),
    .Q(\spi_rd_bus_ff1[24] ),
    .CLK(net298));
 sg13g2_dfrbpq_1 _1633_ (.RESET_B(net57),
    .D(_0060_),
    .Q(\spi_rd_bus_ff1[25] ),
    .CLK(net296));
 sg13g2_dfrbpq_1 _1634_ (.RESET_B(net56),
    .D(_0061_),
    .Q(\spi_rd_bus_ff1[26] ),
    .CLK(net298));
 sg13g2_dfrbpq_1 _1635_ (.RESET_B(net55),
    .D(_0062_),
    .Q(\spi_rd_bus_ff1[32] ),
    .CLK(net296));
 sg13g2_dfrbpq_1 _1636_ (.RESET_B(net54),
    .D(_0063_),
    .Q(\spi_rd_bus_ff1[33] ),
    .CLK(net280));
 sg13g2_dfrbpq_1 _1637_ (.RESET_B(net53),
    .D(_0064_),
    .Q(\spi_rd_bus_ff1[34] ),
    .CLK(net290));
 sg13g2_dfrbpq_1 _1638_ (.RESET_B(net52),
    .D(_0065_),
    .Q(\spi_rd_bus_ff1[35] ),
    .CLK(net282));
 sg13g2_dfrbpq_1 _1639_ (.RESET_B(net51),
    .D(_0066_),
    .Q(\spi_rd_bus_ff1[36] ),
    .CLK(net282));
 sg13g2_dfrbpq_1 _1640_ (.RESET_B(net50),
    .D(_0067_),
    .Q(\spi_rd_bus_ff1[37] ),
    .CLK(net281));
 sg13g2_dfrbpq_1 _1641_ (.RESET_B(net49),
    .D(_0068_),
    .Q(\spi_rd_bus_ff1[38] ),
    .CLK(net276));
 sg13g2_dfrbpq_1 _1642_ (.RESET_B(net48),
    .D(_0069_),
    .Q(\spi_rd_bus_ff1[39] ),
    .CLK(net276));
 sg13g2_dfrbpq_1 _1643_ (.RESET_B(net47),
    .D(_0070_),
    .Q(\spi_rd_bus_ff1[44] ),
    .CLK(net280));
 sg13g2_dfrbpq_1 _1644_ (.RESET_B(net46),
    .D(_0071_),
    .Q(\spi_rd_bus_ff1[45] ),
    .CLK(net295));
 sg13g2_dfrbpq_1 _1645_ (.RESET_B(net45),
    .D(_0072_),
    .Q(\spi_rd_bus_ff1[46] ),
    .CLK(net301));
 sg13g2_dfrbpq_1 _1646_ (.RESET_B(net44),
    .D(_0073_),
    .Q(\spi_rd_bus_ff1[47] ),
    .CLK(net280));
 sg13g2_dfrbpq_1 _1647_ (.RESET_B(net43),
    .D(_0074_),
    .Q(\spi_rd_bus_ff1[48] ),
    .CLK(net300));
 sg13g2_dfrbpq_1 _1648_ (.RESET_B(net42),
    .D(_0075_),
    .Q(\spi_rd_bus_ff1[49] ),
    .CLK(net300));
 sg13g2_dfrbpq_1 _1649_ (.RESET_B(net41),
    .D(_0076_),
    .Q(\spi_rd_bus_ff1[50] ),
    .CLK(net300));
 sg13g2_dfrbpq_1 _1650_ (.RESET_B(net40),
    .D(_0077_),
    .Q(\spi_rd_bus_ff1[51] ),
    .CLK(net298));
 sg13g2_dfrbpq_1 _1651_ (.RESET_B(net39),
    .D(_0078_),
    .Q(\spi_rd_bus_ff1[52] ),
    .CLK(net299));
 sg13g2_dfrbpq_1 _1652_ (.RESET_B(net38),
    .D(_0079_),
    .Q(\spi_rd_bus_ff1[53] ),
    .CLK(net298));
 sg13g2_dfrbpq_1 _1653_ (.RESET_B(net37),
    .D(_0080_),
    .Q(\spi_rd_bus_ff1[54] ),
    .CLK(net289));
 sg13g2_dfrbpq_1 _1654_ (.RESET_B(net36),
    .D(_0081_),
    .Q(\spi_rd_bus_ff1[55] ),
    .CLK(net289));
 sg13g2_dfrbpq_1 _1655_ (.RESET_B(net35),
    .D(_0082_),
    .Q(\spi_rd_bus_ff1[56] ),
    .CLK(net297));
 sg13g2_dfrbpq_1 _1656_ (.RESET_B(net34),
    .D(_0083_),
    .Q(\spi_rd_bus_ff1[57] ),
    .CLK(net298));
 sg13g2_dfrbpq_1 _1657_ (.RESET_B(net33),
    .D(_0084_),
    .Q(\spi_rd_bus_ff1[58] ),
    .CLK(net300));
 sg13g2_dfrbpq_1 _1658_ (.RESET_B(net32),
    .D(_0085_),
    .Q(\spi_rd_bus_ff1[59] ),
    .CLK(net291));
 sg13g2_dfrbpq_1 _1659_ (.RESET_B(net31),
    .D(_0086_),
    .Q(\spi_rd_bus_ff1[60] ),
    .CLK(net282));
 sg13g2_dfrbpq_1 _1660_ (.RESET_B(net30),
    .D(_0087_),
    .Q(\spi_rd_bus_ff1[61] ),
    .CLK(net290));
 sg13g2_dfrbpq_1 _1661_ (.RESET_B(net29),
    .D(_0088_),
    .Q(\spi_rd_bus_ff1[62] ),
    .CLK(net276));
 sg13g2_dfrbpq_1 _1662_ (.RESET_B(net28),
    .D(_0089_),
    .Q(\spi_rd_bus_ff1[63] ),
    .CLK(net280));
 sg13g2_dfrbpq_1 _1663_ (.RESET_B(net342),
    .D(_0090_),
    .Q(\reg_absdiff_rdback[0] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_1 _1664_ (.RESET_B(net344),
    .D(_0091_),
    .Q(\reg_absdiff_rdback[1] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_1 _1665_ (.RESET_B(net346),
    .D(_0092_),
    .Q(\reg_absdiff_rdback[2] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_1 _1666_ (.RESET_B(net326),
    .D(_0093_),
    .Q(\reg_absdiff_rdback[3] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _1667_ (.RESET_B(net317),
    .D(_0094_),
    .Q(\reg_absdiff_rdback[4] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _1668_ (.RESET_B(net326),
    .D(_0095_),
    .Q(\reg_absdiff_rdback[5] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_1 _1669_ (.RESET_B(net316),
    .D(_0096_),
    .Q(\reg_absdiff_rdback[6] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_1 _1670_ (.RESET_B(net316),
    .D(_0097_),
    .Q(\reg_absdiff_rdback[7] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_2 _1671_ (.RESET_B(net348),
    .D(_0098_),
    .Q(\pixel_q[0] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _1672_ (.RESET_B(net344),
    .D(_0099_),
    .Q(\pixel_q[1] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _1673_ (.RESET_B(net344),
    .D(_0100_),
    .Q(\pixel_q[2] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _1674_ (.RESET_B(net348),
    .D(_0101_),
    .Q(\pixel_q[3] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _1675_ (.RESET_B(net348),
    .D(_0102_),
    .Q(\pixel_q[4] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_2 _1676_ (.RESET_B(net336),
    .D(_0103_),
    .Q(\pixel_q[5] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _1677_ (.RESET_B(net336),
    .D(_0104_),
    .Q(\pixel_q[6] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_2 _1678_ (.RESET_B(net337),
    .D(_0105_),
    .Q(\pixel_q[7] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _1679_ (.RESET_B(net347),
    .D(net205),
    .Q(\prev_pixel[0] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_1 _1680_ (.RESET_B(net346),
    .D(net217),
    .Q(\prev_pixel[1] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_1 _1681_ (.RESET_B(net346),
    .D(net215),
    .Q(\prev_pixel[2] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _1682_ (.RESET_B(net347),
    .D(net235),
    .Q(\prev_pixel[3] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _1683_ (.RESET_B(net348),
    .D(net221),
    .Q(\prev_pixel[4] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_1 _1684_ (.RESET_B(net336),
    .D(net382),
    .Q(\prev_pixel[5] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _1685_ (.RESET_B(net337),
    .D(net209),
    .Q(\prev_pixel[6] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _1686_ (.RESET_B(net337),
    .D(net376),
    .Q(\prev_pixel[7] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _1687_ (.RESET_B(net349),
    .D(_0114_),
    .Q(\mean_q[0] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _1688_ (.RESET_B(net346),
    .D(net392),
    .Q(\mean_q[1] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _1689_ (.RESET_B(net346),
    .D(_0116_),
    .Q(\mean_q[2] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _1690_ (.RESET_B(net347),
    .D(_0117_),
    .Q(\mean_q[3] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _1691_ (.RESET_B(net348),
    .D(_0118_),
    .Q(\mean_q[4] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _1692_ (.RESET_B(net348),
    .D(_0119_),
    .Q(\mean_q[5] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _1693_ (.RESET_B(net336),
    .D(_0120_),
    .Q(\mean_q[6] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_2 _1694_ (.RESET_B(net337),
    .D(net386),
    .Q(\mean_q[7] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _1695_ (.RESET_B(net338),
    .D(_0000_),
    .Q(cfg_miso),
    .CLK(_0029_));
 sg13g2_dfrbpq_2 _1696_ (.RESET_B(net337),
    .D(net213),
    .Q(uo_out[0]),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _1697_ (.RESET_B(net337),
    .D(net219),
    .Q(uo_out[1]),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_2 _1698_ (.RESET_B(net336),
    .D(net231),
    .Q(uo_out[2]),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_2 _1699_ (.RESET_B(net336),
    .D(net211),
    .Q(uo_out[3]),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_2 _1700_ (.RESET_B(net336),
    .D(net360),
    .Q(uo_out[4]),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_2 _1701_ (.RESET_B(net336),
    .D(net229),
    .Q(uo_out[5]),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_2 _1702_ (.RESET_B(net338),
    .D(net227),
    .Q(uo_out[6]),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _1703_ (.RESET_B(net338),
    .D(net223),
    .Q(uo_out[7]),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_1 _1704_ (.RESET_B(net331),
    .D(_0130_),
    .Q(spi_wr_toggle),
    .CLK(net295));
 sg13g2_dfrbpq_1 _1705_ (.RESET_B(net313),
    .D(_0131_),
    .Q(\spi_wr_addr[0] ),
    .CLK(net278));
 sg13g2_dfrbpq_1 _1706_ (.RESET_B(net313),
    .D(_0132_),
    .Q(\spi_wr_addr[1] ),
    .CLK(net278));
 sg13g2_dfrbpq_1 _1707_ (.RESET_B(net313),
    .D(_0133_),
    .Q(\spi_wr_addr[2] ),
    .CLK(net278));
 sg13g2_dfrbpq_1 _1708_ (.RESET_B(net333),
    .D(_0134_),
    .Q(\spi_wr_data[0] ),
    .CLK(net295));
 sg13g2_dfrbpq_1 _1709_ (.RESET_B(net331),
    .D(_0135_),
    .Q(\spi_wr_data[1] ),
    .CLK(net295));
 sg13g2_dfrbpq_1 _1710_ (.RESET_B(net331),
    .D(_0136_),
    .Q(\spi_wr_data[2] ),
    .CLK(net295));
 sg13g2_dfrbpq_1 _1711_ (.RESET_B(net313),
    .D(_0137_),
    .Q(\spi_wr_data[3] ),
    .CLK(net278));
 sg13g2_dfrbpq_1 _1712_ (.RESET_B(net310),
    .D(_0138_),
    .Q(\spi_wr_data[4] ),
    .CLK(net276));
 sg13g2_dfrbpq_1 _1713_ (.RESET_B(net310),
    .D(_0139_),
    .Q(\spi_wr_data[5] ),
    .CLK(net276));
 sg13g2_dfrbpq_1 _1714_ (.RESET_B(net310),
    .D(_0140_),
    .Q(\spi_wr_data[6] ),
    .CLK(net276));
 sg13g2_dfrbpq_1 _1715_ (.RESET_B(net311),
    .D(_0141_),
    .Q(\spi_wr_data[7] ),
    .CLK(net277));
 sg13g2_dfrbpq_2 _1716_ (.RESET_B(net311),
    .D(_0001_),
    .Q(\spi_bitcnt[0] ),
    .CLK(net277));
 sg13g2_dfrbpq_1 _1717_ (.RESET_B(net311),
    .D(_0002_),
    .Q(\spi_bitcnt[1] ),
    .CLK(net277));
 sg13g2_dfrbpq_1 _1718_ (.RESET_B(net311),
    .D(_0003_),
    .Q(\spi_bitcnt[2] ),
    .CLK(net277));
 sg13g2_dfrbpq_1 _1719_ (.RESET_B(net311),
    .D(_0004_),
    .Q(\spi_bitcnt[3] ),
    .CLK(net277));
 sg13g2_dfrbpq_1 _1720_ (.RESET_B(net333),
    .D(_0142_),
    .Q(\spi_shift_in[0] ),
    .CLK(net295));
 sg13g2_dfrbpq_1 _1721_ (.RESET_B(net331),
    .D(_0143_),
    .Q(\spi_shift_in[1] ),
    .CLK(net295));
 sg13g2_dfrbpq_1 _1722_ (.RESET_B(net331),
    .D(_0144_),
    .Q(\spi_shift_in[2] ),
    .CLK(net295));
 sg13g2_dfrbpq_2 _1723_ (.RESET_B(net314),
    .D(_0145_),
    .Q(\spi_shift_in[3] ),
    .CLK(net279));
 sg13g2_dfrbpq_2 _1724_ (.RESET_B(net312),
    .D(_0146_),
    .Q(\spi_shift_in[4] ),
    .CLK(net279));
 sg13g2_dfrbpq_2 _1725_ (.RESET_B(net314),
    .D(_0147_),
    .Q(\spi_shift_in[5] ),
    .CLK(net278));
 sg13g2_dfrbpq_1 _1726_ (.RESET_B(net311),
    .D(_0148_),
    .Q(\spi_shift_in[6] ),
    .CLK(net277));
 sg13g2_dfrbpq_1 _1727_ (.RESET_B(net311),
    .D(_0149_),
    .Q(_0013_),
    .CLK(net277));
 sg13g2_dfrbpq_1 _1728_ (.RESET_B(net311),
    .D(_0150_),
    .Q(spi_cmd_wr),
    .CLK(net277));
 sg13g2_dfrbpq_1 _1729_ (.RESET_B(net313),
    .D(_0151_),
    .Q(\spi_cmd_addr[0] ),
    .CLK(net278));
 sg13g2_dfrbpq_1 _1730_ (.RESET_B(net313),
    .D(_0152_),
    .Q(\spi_cmd_addr[1] ),
    .CLK(net278));
 sg13g2_dfrbpq_1 _1731_ (.RESET_B(net313),
    .D(_0153_),
    .Q(\spi_cmd_addr[2] ),
    .CLK(net278));
 sg13g2_dfrbpq_2 _1732_ (.RESET_B(net325),
    .D(net236),
    .Q(spi_shift_out_load_pending),
    .CLK(net288));
 sg13g2_dfrbpq_1 _1733_ (.RESET_B(net310),
    .D(net275),
    .Q(_0014_),
    .CLK(net276));
 sg13g2_dfrbpq_1 _1734_ (.RESET_B(net328),
    .D(_0154_),
    .Q(\spi_shift_out_load[0] ),
    .CLK(net292));
 sg13g2_dfrbpq_1 _1735_ (.RESET_B(net328),
    .D(_0155_),
    .Q(\spi_shift_out_load[1] ),
    .CLK(net292));
 sg13g2_dfrbpq_1 _1736_ (.RESET_B(net328),
    .D(_0156_),
    .Q(\spi_shift_out_load[2] ),
    .CLK(net292));
 sg13g2_dfrbpq_1 _1737_ (.RESET_B(net328),
    .D(_0157_),
    .Q(\spi_shift_out_load[3] ),
    .CLK(net292));
 sg13g2_dfrbpq_1 _1738_ (.RESET_B(net323),
    .D(_0158_),
    .Q(\spi_shift_out_load[4] ),
    .CLK(net286));
 sg13g2_dfrbpq_1 _1739_ (.RESET_B(net323),
    .D(_0159_),
    .Q(\spi_shift_out_load[5] ),
    .CLK(net286));
 sg13g2_dfrbpq_1 _1740_ (.RESET_B(net324),
    .D(_0160_),
    .Q(\spi_shift_out_load[6] ),
    .CLK(net287));
 sg13g2_dfrbpq_1 _1741_ (.RESET_B(net324),
    .D(_0161_),
    .Q(\spi_shift_out_load[7] ),
    .CLK(net287));
 sg13g2_dfrbpq_1 _1742_ (.RESET_B(net339),
    .D(net372),
    .Q(\reg_thresh[0] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_2 _1743_ (.RESET_B(net339),
    .D(net233),
    .Q(\reg_thresh[1] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_1 _1744_ (.RESET_B(net339),
    .D(net207),
    .Q(\reg_thresh[2] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_1 _1745_ (.RESET_B(net339),
    .D(net225),
    .Q(\reg_thresh[3] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _1746_ (.RESET_B(net316),
    .D(net183),
    .Q(\reg_thresh[4] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _1747_ (.RESET_B(net305),
    .D(net354),
    .Q(\reg_thresh[5] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_2 _1748_ (.RESET_B(net305),
    .D(net175),
    .Q(\reg_thresh[6] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_2 _1749_ (.RESET_B(net307),
    .D(net153),
    .Q(_0015_),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _1750_ (.RESET_B(net335),
    .D(net364),
    .Q(\reg_contrast_thr[0] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _1751_ (.RESET_B(net334),
    .D(net358),
    .Q(\reg_contrast_thr[1] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _1752_ (.RESET_B(net318),
    .D(net169),
    .Q(_0016_),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _1753_ (.RESET_B(net318),
    .D(net187),
    .Q(_0017_),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_2 _1754_ (.RESET_B(net305),
    .D(net384),
    .Q(\reg_contrast_thr[4] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_2 _1755_ (.RESET_B(net308),
    .D(net370),
    .Q(\reg_contrast_thr[5] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_2 _1756_ (.RESET_B(net305),
    .D(net366),
    .Q(\reg_contrast_thr[6] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_1 _1757_ (.RESET_B(net316),
    .D(net203),
    .Q(\reg_contrast_thr[7] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_2 _1758_ (.RESET_B(net335),
    .D(net374),
    .Q(\reg_edge_thr[0] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _1759_ (.RESET_B(net334),
    .D(net362),
    .Q(\reg_edge_thr[1] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _1760_ (.RESET_B(net334),
    .D(net166),
    .Q(_0018_),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _1761_ (.RESET_B(net318),
    .D(net193),
    .Q(_0019_),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _1762_ (.RESET_B(net308),
    .D(net378),
    .Q(\reg_edge_thr[4] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_2 _1763_ (.RESET_B(net307),
    .D(net356),
    .Q(\reg_edge_thr[5] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_1 _1764_ (.RESET_B(net307),
    .D(net180),
    .Q(\reg_edge_thr[6] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_1 _1765_ (.RESET_B(net307),
    .D(net164),
    .Q(\reg_edge_thr[7] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_1 _1766_ (.RESET_B(net339),
    .D(net177),
    .Q(_0020_),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_2 _1767_ (.RESET_B(net339),
    .D(net172),
    .Q(_0021_),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_1 _1768_ (.RESET_B(net340),
    .D(net390),
    .Q(\reg_alpha_shift[2] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_1 _1769_ (.RESET_B(net331),
    .D(spi_wr_toggle),
    .Q(cfg_wr_toggle_ff1),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _1770_ (.RESET_B(net332),
    .D(net142),
    .Q(cfg_wr_toggle_ff2),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _1771_ (.RESET_B(net332),
    .D(net151),
    .Q(cfg_wr_toggle_ff2_d),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_1 _1772_ (.RESET_B(net332),
    .D(\spi_wr_addr[0] ),
    .Q(\cfg_wr_addr_ff1[0] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _1773_ (.RESET_B(net314),
    .D(\spi_wr_addr[1] ),
    .Q(\cfg_wr_addr_ff1[1] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _1774_ (.RESET_B(net314),
    .D(\spi_wr_addr[2] ),
    .Q(\cfg_wr_addr_ff1[2] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _1775_ (.RESET_B(net332),
    .D(net144),
    .Q(\cfg_wr_addr_ff2[0] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_2 _1776_ (.RESET_B(net313),
    .D(net147),
    .Q(\cfg_wr_addr_ff2[1] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_2 _1777_ (.RESET_B(net332),
    .D(net150),
    .Q(\cfg_wr_addr_ff2[2] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _1778_ (.RESET_B(net333),
    .D(\spi_wr_data[0] ),
    .Q(\cfg_wr_data_ff1[0] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _1779_ (.RESET_B(net331),
    .D(\spi_wr_data[1] ),
    .Q(\cfg_wr_data_ff1[1] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _1780_ (.RESET_B(net331),
    .D(\spi_wr_data[2] ),
    .Q(\cfg_wr_data_ff1[2] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _1781_ (.RESET_B(net314),
    .D(\spi_wr_data[3] ),
    .Q(\cfg_wr_data_ff1[3] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_1 _1782_ (.RESET_B(net310),
    .D(\spi_wr_data[4] ),
    .Q(\cfg_wr_data_ff1[4] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_1 _1783_ (.RESET_B(net310),
    .D(\spi_wr_data[5] ),
    .Q(\cfg_wr_data_ff1[5] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_1 _1784_ (.RESET_B(net310),
    .D(\spi_wr_data[6] ),
    .Q(\cfg_wr_data_ff1[6] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_1 _1785_ (.RESET_B(net312),
    .D(\spi_wr_data[7] ),
    .Q(\cfg_wr_data_ff1[7] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _1786_ (.RESET_B(net334),
    .D(net145),
    .Q(\cfg_wr_data_ff2[0] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_2 _1787_ (.RESET_B(net334),
    .D(net146),
    .Q(\cfg_wr_data_ff2[1] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _1788_ (.RESET_B(net334),
    .D(net148),
    .Q(\cfg_wr_data_ff2[2] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_2 _1789_ (.RESET_B(net318),
    .D(net139),
    .Q(\cfg_wr_data_ff2[3] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_2 _1790_ (.RESET_B(net307),
    .D(net143),
    .Q(\cfg_wr_data_ff2[4] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_2 _1791_ (.RESET_B(net307),
    .D(net140),
    .Q(\cfg_wr_data_ff2[5] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_2 _1792_ (.RESET_B(net310),
    .D(net141),
    .Q(\cfg_wr_data_ff2[6] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_2 _1793_ (.RESET_B(net312),
    .D(net149),
    .Q(\cfg_wr_data_ff2[7] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_1 _1794_ (.RESET_B(net129),
    .D(_0189_),
    .Q(\spi_rd_bus_ff2[0] ),
    .CLK(net291));
 sg13g2_dfrbpq_1 _1795_ (.RESET_B(net128),
    .D(_0190_),
    .Q(\spi_rd_bus_ff2[1] ),
    .CLK(net293));
 sg13g2_dfrbpq_1 _1796_ (.RESET_B(net127),
    .D(_0191_),
    .Q(\spi_rd_bus_ff2[2] ),
    .CLK(net293));
 sg13g2_dfrbpq_1 _1797_ (.RESET_B(net126),
    .D(_0192_),
    .Q(\spi_rd_bus_ff2[3] ),
    .CLK(net292));
 sg13g2_dfrbpq_1 _1798_ (.RESET_B(net125),
    .D(_0193_),
    .Q(\spi_rd_bus_ff2[4] ),
    .CLK(net288));
 sg13g2_dfrbpq_1 _1799_ (.RESET_B(net124),
    .D(_0194_),
    .Q(\spi_rd_bus_ff2[5] ),
    .CLK(net288));
 sg13g2_dfrbpq_1 _1800_ (.RESET_B(net123),
    .D(_0195_),
    .Q(\spi_rd_bus_ff2[6] ),
    .CLK(net288));
 sg13g2_dfrbpq_1 _1801_ (.RESET_B(net122),
    .D(_0196_),
    .Q(\spi_rd_bus_ff2[7] ),
    .CLK(net283));
 sg13g2_dfrbpq_1 _1802_ (.RESET_B(net121),
    .D(_0197_),
    .Q(\spi_rd_bus_ff2[8] ),
    .CLK(net296));
 sg13g2_dfrbpq_1 _1803_ (.RESET_B(net120),
    .D(_0198_),
    .Q(\spi_rd_bus_ff2[9] ),
    .CLK(net296));
 sg13g2_dfrbpq_1 _1804_ (.RESET_B(net119),
    .D(_0199_),
    .Q(\spi_rd_bus_ff2[10] ),
    .CLK(net293));
 sg13g2_dfrbpq_1 _1805_ (.RESET_B(net118),
    .D(_0200_),
    .Q(\spi_rd_bus_ff2[11] ),
    .CLK(net291));
 sg13g2_dfrbpq_1 _1806_ (.RESET_B(net117),
    .D(_0201_),
    .Q(\spi_rd_bus_ff2[12] ),
    .CLK(net288));
 sg13g2_dfrbpq_1 _1807_ (.RESET_B(net116),
    .D(_0202_),
    .Q(\spi_rd_bus_ff2[13] ),
    .CLK(net284));
 sg13g2_dfrbpq_1 _1808_ (.RESET_B(net115),
    .D(_0203_),
    .Q(\spi_rd_bus_ff2[14] ),
    .CLK(net284));
 sg13g2_dfrbpq_1 _1809_ (.RESET_B(net114),
    .D(_0204_),
    .Q(\spi_rd_bus_ff2[15] ),
    .CLK(net289));
 sg13g2_dfrbpq_1 _1810_ (.RESET_B(net113),
    .D(_0205_),
    .Q(\spi_rd_bus_ff2[16] ),
    .CLK(net296));
 sg13g2_dfrbpq_1 _1811_ (.RESET_B(net112),
    .D(_0206_),
    .Q(\spi_rd_bus_ff2[17] ),
    .CLK(net296));
 sg13g2_dfrbpq_1 _1812_ (.RESET_B(net111),
    .D(_0207_),
    .Q(\spi_rd_bus_ff2[18] ),
    .CLK(net297));
 sg13g2_dfrbpq_1 _1813_ (.RESET_B(net110),
    .D(_0208_),
    .Q(\spi_rd_bus_ff2[19] ),
    .CLK(net291));
 sg13g2_dfrbpq_1 _1814_ (.RESET_B(net109),
    .D(_0209_),
    .Q(\spi_rd_bus_ff2[20] ),
    .CLK(net284));
 sg13g2_dfrbpq_1 _1815_ (.RESET_B(net108),
    .D(_0210_),
    .Q(\spi_rd_bus_ff2[21] ),
    .CLK(net284));
 sg13g2_dfrbpq_1 _1816_ (.RESET_B(net107),
    .D(_0211_),
    .Q(\spi_rd_bus_ff2[22] ),
    .CLK(net283));
 sg13g2_dfrbpq_1 _1817_ (.RESET_B(net106),
    .D(_0212_),
    .Q(\spi_rd_bus_ff2[23] ),
    .CLK(net283));
 sg13g2_dfrbpq_1 _1818_ (.RESET_B(net105),
    .D(_0213_),
    .Q(\spi_rd_bus_ff2[24] ),
    .CLK(net298));
 sg13g2_dfrbpq_1 _1819_ (.RESET_B(net104),
    .D(_0214_),
    .Q(\spi_rd_bus_ff2[25] ),
    .CLK(net297));
 sg13g2_dfrbpq_1 _1820_ (.RESET_B(net103),
    .D(_0215_),
    .Q(\spi_rd_bus_ff2[26] ),
    .CLK(net297));
 sg13g2_dfrbpq_1 _1821_ (.RESET_B(net102),
    .D(_0216_),
    .Q(\spi_rd_bus_ff2[32] ),
    .CLK(net297));
 sg13g2_dfrbpq_1 _1822_ (.RESET_B(net101),
    .D(_0217_),
    .Q(\spi_rd_bus_ff2[33] ),
    .CLK(net290));
 sg13g2_dfrbpq_1 _1823_ (.RESET_B(net100),
    .D(_0218_),
    .Q(\spi_rd_bus_ff2[34] ),
    .CLK(net296));
 sg13g2_dfrbpq_2 _1824_ (.RESET_B(net99),
    .D(_0219_),
    .Q(\spi_rd_bus_ff2[35] ),
    .CLK(net288));
 sg13g2_dfrbpq_1 _1825_ (.RESET_B(net98),
    .D(_0220_),
    .Q(\spi_rd_bus_ff2[36] ),
    .CLK(net285));
 sg13g2_dfrbpq_1 _1826_ (.RESET_B(net97),
    .D(_0221_),
    .Q(\spi_rd_bus_ff2[37] ),
    .CLK(net285));
 sg13g2_dfrbpq_1 _1827_ (.RESET_B(net96),
    .D(_0222_),
    .Q(\spi_rd_bus_ff2[38] ),
    .CLK(net285));
 sg13g2_dfrbpq_1 _1828_ (.RESET_B(net95),
    .D(_0223_),
    .Q(\spi_rd_bus_ff2[39] ),
    .CLK(net283));
 sg13g2_dfrbpq_1 _1829_ (.RESET_B(net94),
    .D(_0224_),
    .Q(\spi_rd_bus_ff2[44] ),
    .CLK(net289));
 sg13g2_dfrbpq_1 _1830_ (.RESET_B(net93),
    .D(_0225_),
    .Q(\spi_rd_bus_ff2[45] ),
    .CLK(net289));
 sg13g2_dfrbpq_1 _1831_ (.RESET_B(net92),
    .D(_0226_),
    .Q(\spi_rd_bus_ff2[46] ),
    .CLK(net280));
 sg13g2_dfrbpq_1 _1832_ (.RESET_B(net91),
    .D(_0227_),
    .Q(\spi_rd_bus_ff2[47] ),
    .CLK(net289));
 sg13g2_dfrbpq_1 _1833_ (.RESET_B(net90),
    .D(_0228_),
    .Q(\spi_rd_bus_ff2[48] ),
    .CLK(net300));
 sg13g2_dfrbpq_1 _1834_ (.RESET_B(net89),
    .D(_0229_),
    .Q(\spi_rd_bus_ff2[49] ),
    .CLK(net300));
 sg13g2_dfrbpq_1 _1835_ (.RESET_B(net88),
    .D(_0230_),
    .Q(\spi_rd_bus_ff2[50] ),
    .CLK(net300));
 sg13g2_dfrbpq_1 _1836_ (.RESET_B(net87),
    .D(_0231_),
    .Q(\spi_rd_bus_ff2[51] ),
    .CLK(net293));
 sg13g2_dfrbpq_1 _1837_ (.RESET_B(net86),
    .D(_0232_),
    .Q(\spi_rd_bus_ff2[52] ),
    .CLK(net290));
 sg13g2_dfrbpq_1 _1838_ (.RESET_B(net85),
    .D(_0233_),
    .Q(\spi_rd_bus_ff2[53] ),
    .CLK(net291));
 sg13g2_dfrbpq_1 _1839_ (.RESET_B(net84),
    .D(_0234_),
    .Q(\spi_rd_bus_ff2[54] ),
    .CLK(net289));
 sg13g2_dfrbpq_1 _1840_ (.RESET_B(net83),
    .D(_0235_),
    .Q(\spi_rd_bus_ff2[55] ),
    .CLK(net284));
 sg13g2_dfrbpq_1 _1841_ (.RESET_B(net137),
    .D(_0236_),
    .Q(\spi_rd_bus_ff2[56] ),
    .CLK(net297));
 sg13g2_dfrbpq_1 _1842_ (.RESET_B(net136),
    .D(_0237_),
    .Q(\spi_rd_bus_ff2[57] ),
    .CLK(net297));
 sg13g2_dfrbpq_1 _1843_ (.RESET_B(net135),
    .D(_0238_),
    .Q(\spi_rd_bus_ff2[58] ),
    .CLK(net301));
 sg13g2_dfrbpq_1 _1844_ (.RESET_B(net134),
    .D(_0239_),
    .Q(\spi_rd_bus_ff2[59] ),
    .CLK(net291));
 sg13g2_dfrbpq_1 _1845_ (.RESET_B(net133),
    .D(_0240_),
    .Q(\spi_rd_bus_ff2[60] ),
    .CLK(net288));
 sg13g2_dfrbpq_1 _1846_ (.RESET_B(net132),
    .D(_0241_),
    .Q(\spi_rd_bus_ff2[61] ),
    .CLK(net291));
 sg13g2_dfrbpq_1 _1847_ (.RESET_B(net131),
    .D(_0242_),
    .Q(\spi_rd_bus_ff2[62] ),
    .CLK(net283));
 sg13g2_dfrbpq_1 _1848_ (.RESET_B(net130),
    .D(_0243_),
    .Q(\spi_rd_bus_ff2[63] ),
    .CLK(net289));
 sg13g2_dfrbpq_1 _1849_ (.RESET_B(net334),
    .D(net388),
    .Q(\reg_mode[0] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _1850_ (.RESET_B(net334),
    .D(net368),
    .Q(\reg_mode[1] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_1 _1851_ (.RESET_B(net318),
    .D(net201),
    .Q(\reg_mode[2] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_1 _1852_ (.RESET_B(net306),
    .D(net199),
    .Q(\reg_mode[3] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_1 _1853_ (.RESET_B(net305),
    .D(net197),
    .Q(\reg_mode[4] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_1 _1854_ (.RESET_B(net305),
    .D(net185),
    .Q(\reg_mode[5] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_1 _1855_ (.RESET_B(net305),
    .D(net195),
    .Q(\reg_mode[6] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_1 _1856_ (.RESET_B(net307),
    .D(net190),
    .Q(\reg_mode[7] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_tiehi _1661__29 (.L_HI(net29));
 sg13g2_tiehi _1660__30 (.L_HI(net30));
 sg13g2_tiehi _1659__31 (.L_HI(net31));
 sg13g2_tiehi _1658__32 (.L_HI(net32));
 sg13g2_tiehi _1657__33 (.L_HI(net33));
 sg13g2_tiehi _1656__34 (.L_HI(net34));
 sg13g2_tiehi _1655__35 (.L_HI(net35));
 sg13g2_tiehi _1654__36 (.L_HI(net36));
 sg13g2_tiehi _1653__37 (.L_HI(net37));
 sg13g2_tiehi _1652__38 (.L_HI(net38));
 sg13g2_tiehi _1651__39 (.L_HI(net39));
 sg13g2_tiehi _1650__40 (.L_HI(net40));
 sg13g2_tiehi _1649__41 (.L_HI(net41));
 sg13g2_tiehi _1648__42 (.L_HI(net42));
 sg13g2_tiehi _1647__43 (.L_HI(net43));
 sg13g2_tiehi _1646__44 (.L_HI(net44));
 sg13g2_tiehi _1645__45 (.L_HI(net45));
 sg13g2_tiehi _1644__46 (.L_HI(net46));
 sg13g2_tiehi _1643__47 (.L_HI(net47));
 sg13g2_tiehi _1642__48 (.L_HI(net48));
 sg13g2_tiehi _1641__49 (.L_HI(net49));
 sg13g2_tiehi _1640__50 (.L_HI(net50));
 sg13g2_tiehi _1639__51 (.L_HI(net51));
 sg13g2_tiehi _1638__52 (.L_HI(net52));
 sg13g2_tiehi _1637__53 (.L_HI(net53));
 sg13g2_tiehi _1636__54 (.L_HI(net54));
 sg13g2_tiehi _1635__55 (.L_HI(net55));
 sg13g2_tiehi _1634__56 (.L_HI(net56));
 sg13g2_tiehi _1633__57 (.L_HI(net57));
 sg13g2_tiehi _1632__58 (.L_HI(net58));
 sg13g2_tiehi _1631__59 (.L_HI(net59));
 sg13g2_tiehi _1630__60 (.L_HI(net60));
 sg13g2_tiehi _1629__61 (.L_HI(net61));
 sg13g2_tiehi _1628__62 (.L_HI(net62));
 sg13g2_tiehi _1627__63 (.L_HI(net63));
 sg13g2_tiehi _1626__64 (.L_HI(net64));
 sg13g2_tiehi _1625__65 (.L_HI(net65));
 sg13g2_tiehi _1624__66 (.L_HI(net66));
 sg13g2_tiehi _1623__67 (.L_HI(net67));
 sg13g2_tiehi _1622__68 (.L_HI(net68));
 sg13g2_tiehi _1621__69 (.L_HI(net69));
 sg13g2_tiehi _1620__70 (.L_HI(net70));
 sg13g2_tiehi _1619__71 (.L_HI(net71));
 sg13g2_tiehi _1618__72 (.L_HI(net72));
 sg13g2_tiehi _1617__73 (.L_HI(net73));
 sg13g2_tiehi _1616__74 (.L_HI(net74));
 sg13g2_tiehi _1615__75 (.L_HI(net75));
 sg13g2_tiehi _1614__76 (.L_HI(net76));
 sg13g2_tiehi _1613__77 (.L_HI(net77));
 sg13g2_tiehi _1612__78 (.L_HI(net78));
 sg13g2_tiehi _1611__79 (.L_HI(net79));
 sg13g2_tiehi _1610__80 (.L_HI(net80));
 sg13g2_tiehi _1609__81 (.L_HI(net81));
 sg13g2_tiehi _1608__82 (.L_HI(net82));
 sg13g2_tiehi _1840__83 (.L_HI(net83));
 sg13g2_tiehi _1839__84 (.L_HI(net84));
 sg13g2_tiehi _1838__85 (.L_HI(net85));
 sg13g2_tiehi _1837__86 (.L_HI(net86));
 sg13g2_tiehi _1836__87 (.L_HI(net87));
 sg13g2_tiehi _1835__88 (.L_HI(net88));
 sg13g2_tiehi _1834__89 (.L_HI(net89));
 sg13g2_tiehi _1833__90 (.L_HI(net90));
 sg13g2_tiehi _1832__91 (.L_HI(net91));
 sg13g2_tiehi _1831__92 (.L_HI(net92));
 sg13g2_tiehi _1830__93 (.L_HI(net93));
 sg13g2_tiehi _1829__94 (.L_HI(net94));
 sg13g2_tiehi _1828__95 (.L_HI(net95));
 sg13g2_tiehi _1827__96 (.L_HI(net96));
 sg13g2_tiehi _1826__97 (.L_HI(net97));
 sg13g2_tiehi _1825__98 (.L_HI(net98));
 sg13g2_tiehi _1824__99 (.L_HI(net99));
 sg13g2_tiehi _1823__100 (.L_HI(net100));
 sg13g2_tiehi _1822__101 (.L_HI(net101));
 sg13g2_tiehi _1821__102 (.L_HI(net102));
 sg13g2_tiehi _1820__103 (.L_HI(net103));
 sg13g2_tiehi _1819__104 (.L_HI(net104));
 sg13g2_tiehi _1818__105 (.L_HI(net105));
 sg13g2_tiehi _1817__106 (.L_HI(net106));
 sg13g2_tiehi _1816__107 (.L_HI(net107));
 sg13g2_tiehi _1815__108 (.L_HI(net108));
 sg13g2_tiehi _1814__109 (.L_HI(net109));
 sg13g2_tiehi _1813__110 (.L_HI(net110));
 sg13g2_tiehi _1812__111 (.L_HI(net111));
 sg13g2_tiehi _1811__112 (.L_HI(net112));
 sg13g2_tiehi _1810__113 (.L_HI(net113));
 sg13g2_tiehi _1809__114 (.L_HI(net114));
 sg13g2_tiehi _1808__115 (.L_HI(net115));
 sg13g2_tiehi _1807__116 (.L_HI(net116));
 sg13g2_tiehi _1806__117 (.L_HI(net117));
 sg13g2_tiehi _1805__118 (.L_HI(net118));
 sg13g2_tiehi _1804__119 (.L_HI(net119));
 sg13g2_tiehi _1803__120 (.L_HI(net120));
 sg13g2_tiehi _1802__121 (.L_HI(net121));
 sg13g2_tiehi _1801__122 (.L_HI(net122));
 sg13g2_tiehi _1800__123 (.L_HI(net123));
 sg13g2_tiehi _1799__124 (.L_HI(net124));
 sg13g2_tiehi _1798__125 (.L_HI(net125));
 sg13g2_tiehi _1797__126 (.L_HI(net126));
 sg13g2_tiehi _1796__127 (.L_HI(net127));
 sg13g2_tiehi _1795__128 (.L_HI(net128));
 sg13g2_tiehi _1794__129 (.L_HI(net129));
 sg13g2_tiehi _1848__130 (.L_HI(net130));
 sg13g2_tiehi _1847__131 (.L_HI(net131));
 sg13g2_tiehi _1846__132 (.L_HI(net132));
 sg13g2_tiehi _1845__133 (.L_HI(net133));
 sg13g2_tiehi _1844__134 (.L_HI(net134));
 sg13g2_tiehi _1843__135 (.L_HI(net135));
 sg13g2_tiehi _1842__136 (.L_HI(net136));
 sg13g2_tiehi _1841__137 (.L_HI(net137));
 sg13g2_tiehi tt_um_ebeam_pixel_core_138 (.L_HI(net138));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_ebeam_pixel_core_15 (.L_LO(net15));
 sg13g2_tielo tt_um_ebeam_pixel_core_16 (.L_LO(net16));
 sg13g2_tielo tt_um_ebeam_pixel_core_17 (.L_LO(net17));
 sg13g2_tielo tt_um_ebeam_pixel_core_18 (.L_LO(net18));
 sg13g2_tielo tt_um_ebeam_pixel_core_19 (.L_LO(net19));
 sg13g2_tielo tt_um_ebeam_pixel_core_20 (.L_LO(net20));
 sg13g2_tielo tt_um_ebeam_pixel_core_21 (.L_LO(net21));
 sg13g2_tielo tt_um_ebeam_pixel_core_22 (.L_LO(net22));
 sg13g2_tielo tt_um_ebeam_pixel_core_23 (.L_LO(net23));
 sg13g2_tielo tt_um_ebeam_pixel_core_24 (.L_LO(net24));
 sg13g2_tielo tt_um_ebeam_pixel_core_25 (.L_LO(net25));
 sg13g2_tielo tt_um_ebeam_pixel_core_26 (.L_LO(net26));
 sg13g2_tielo tt_um_ebeam_pixel_core_27 (.L_LO(net27));
 sg13g2_tiehi _1662__28 (.L_HI(net28));
 sg13g2_buf_8 _1982_ (.A(cfg_miso),
    .X(uio_out[5]));
 sg13g2_buf_8 fanout236 (.A(_0012_),
    .X(net236));
 sg13g2_buf_8 fanout237 (.A(_0435_),
    .X(net237));
 sg13g2_buf_8 fanout238 (.A(_0358_),
    .X(net238));
 sg13g2_buf_1 fanout239 (.A(_0358_),
    .X(net239));
 sg13g2_buf_8 fanout240 (.A(_0353_),
    .X(net240));
 sg13g2_buf_8 fanout241 (.A(_0346_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_0346_),
    .X(net242));
 sg13g2_buf_8 fanout243 (.A(_0264_),
    .X(net243));
 sg13g2_buf_8 fanout244 (.A(_0264_),
    .X(net244));
 sg13g2_buf_8 fanout245 (.A(_0286_),
    .X(net245));
 sg13g2_buf_8 fanout246 (.A(_0284_),
    .X(net246));
 sg13g2_buf_8 fanout247 (.A(_0426_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_0426_),
    .X(net248));
 sg13g2_buf_8 fanout249 (.A(net250),
    .X(net249));
 sg13g2_buf_8 fanout250 (.A(net387),
    .X(net250));
 sg13g2_buf_8 fanout251 (.A(net253),
    .X(net251));
 sg13g2_buf_1 fanout252 (.A(net253),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(net389),
    .X(net253));
 sg13g2_buf_8 fanout254 (.A(_0021_),
    .X(net254));
 sg13g2_buf_8 fanout255 (.A(net256),
    .X(net255));
 sg13g2_buf_8 fanout256 (.A(_0020_),
    .X(net256));
 sg13g2_buf_8 fanout257 (.A(spi_shift_out_load_pending),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(spi_shift_out_load_pending),
    .X(net258));
 sg13g2_buf_8 fanout259 (.A(\spi_shift_in[5] ),
    .X(net259));
 sg13g2_buf_8 fanout260 (.A(\pixel_q[6] ),
    .X(net260));
 sg13g2_buf_8 fanout261 (.A(net262),
    .X(net261));
 sg13g2_buf_1 fanout262 (.A(net263),
    .X(net262));
 sg13g2_buf_1 fanout263 (.A(net264),
    .X(net263));
 sg13g2_buf_1 fanout264 (.A(_0437_),
    .X(net264));
 sg13g2_buf_8 fanout265 (.A(net266),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(net272),
    .X(net266));
 sg13g2_buf_8 fanout267 (.A(net268),
    .X(net267));
 sg13g2_buf_8 fanout268 (.A(net272),
    .X(net268));
 sg13g2_buf_8 fanout269 (.A(net272),
    .X(net269));
 sg13g2_buf_1 fanout270 (.A(net271),
    .X(net270));
 sg13g2_buf_8 fanout271 (.A(net272),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_0437_),
    .X(net272));
 sg13g2_buf_8 fanout273 (.A(_0437_),
    .X(net273));
 sg13g2_buf_8 fanout274 (.A(_0397_),
    .X(net274));
 sg13g2_buf_8 fanout275 (.A(_0030_),
    .X(net275));
 sg13g2_buf_8 fanout276 (.A(net281),
    .X(net276));
 sg13g2_buf_8 fanout277 (.A(net279),
    .X(net277));
 sg13g2_buf_8 fanout278 (.A(net279),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(net280),
    .X(net279));
 sg13g2_buf_8 fanout280 (.A(net281),
    .X(net280));
 sg13g2_buf_8 fanout281 (.A(uio_in[3]),
    .X(net281));
 sg13g2_buf_8 fanout282 (.A(net285),
    .X(net282));
 sg13g2_buf_8 fanout283 (.A(net285),
    .X(net283));
 sg13g2_buf_1 fanout284 (.A(net285),
    .X(net284));
 sg13g2_buf_8 fanout285 (.A(net294),
    .X(net285));
 sg13g2_buf_8 fanout286 (.A(net287),
    .X(net286));
 sg13g2_buf_1 fanout287 (.A(net288),
    .X(net287));
 sg13g2_buf_8 fanout288 (.A(net294),
    .X(net288));
 sg13g2_buf_8 fanout289 (.A(net290),
    .X(net289));
 sg13g2_buf_8 fanout290 (.A(net294),
    .X(net290));
 sg13g2_buf_8 fanout291 (.A(net293),
    .X(net291));
 sg13g2_buf_1 fanout292 (.A(net293),
    .X(net292));
 sg13g2_buf_8 fanout293 (.A(net294),
    .X(net293));
 sg13g2_buf_8 fanout294 (.A(uio_in[3]),
    .X(net294));
 sg13g2_buf_8 fanout295 (.A(net301),
    .X(net295));
 sg13g2_buf_8 fanout296 (.A(net298),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(net298),
    .X(net297));
 sg13g2_buf_8 fanout298 (.A(net299),
    .X(net298));
 sg13g2_buf_8 fanout299 (.A(net300),
    .X(net299));
 sg13g2_buf_8 fanout300 (.A(net301),
    .X(net300));
 sg13g2_buf_8 fanout301 (.A(uio_in[3]),
    .X(net301));
 sg13g2_buf_8 fanout302 (.A(net12),
    .X(net302));
 sg13g2_buf_8 fanout303 (.A(net304),
    .X(net303));
 sg13g2_buf_8 fanout304 (.A(net11),
    .X(net304));
 sg13g2_buf_8 fanout305 (.A(net319),
    .X(net305));
 sg13g2_buf_1 fanout306 (.A(net319),
    .X(net306));
 sg13g2_buf_8 fanout307 (.A(net309),
    .X(net307));
 sg13g2_buf_8 fanout308 (.A(net309),
    .X(net308));
 sg13g2_buf_1 fanout309 (.A(net319),
    .X(net309));
 sg13g2_buf_8 fanout310 (.A(net319),
    .X(net310));
 sg13g2_buf_8 fanout311 (.A(net315),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(net315),
    .X(net312));
 sg13g2_buf_8 fanout313 (.A(net315),
    .X(net313));
 sg13g2_buf_8 fanout314 (.A(net315),
    .X(net314));
 sg13g2_buf_8 fanout315 (.A(net319),
    .X(net315));
 sg13g2_buf_8 fanout316 (.A(net318),
    .X(net316));
 sg13g2_buf_1 fanout317 (.A(net318),
    .X(net317));
 sg13g2_buf_8 fanout318 (.A(net319),
    .X(net318));
 sg13g2_buf_8 fanout319 (.A(net351),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(net321),
    .X(net320));
 sg13g2_buf_8 fanout321 (.A(net322),
    .X(net321));
 sg13g2_buf_8 fanout322 (.A(net325),
    .X(net322));
 sg13g2_buf_8 fanout323 (.A(net324),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(net325),
    .X(net324));
 sg13g2_buf_8 fanout325 (.A(net351),
    .X(net325));
 sg13g2_buf_8 fanout326 (.A(net327),
    .X(net326));
 sg13g2_buf_8 fanout327 (.A(net330),
    .X(net327));
 sg13g2_buf_8 fanout328 (.A(net330),
    .X(net328));
 sg13g2_buf_1 fanout329 (.A(net330),
    .X(net329));
 sg13g2_buf_8 fanout330 (.A(net351),
    .X(net330));
 sg13g2_buf_8 fanout331 (.A(net333),
    .X(net331));
 sg13g2_buf_8 fanout332 (.A(net333),
    .X(net332));
 sg13g2_buf_8 fanout333 (.A(net350),
    .X(net333));
 sg13g2_buf_8 fanout334 (.A(net335),
    .X(net334));
 sg13g2_buf_8 fanout335 (.A(net350),
    .X(net335));
 sg13g2_buf_8 fanout336 (.A(net337),
    .X(net336));
 sg13g2_buf_8 fanout337 (.A(net338),
    .X(net337));
 sg13g2_buf_8 fanout338 (.A(net350),
    .X(net338));
 sg13g2_buf_8 fanout339 (.A(net341),
    .X(net339));
 sg13g2_buf_1 fanout340 (.A(net341),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(net345),
    .X(net341));
 sg13g2_buf_8 fanout342 (.A(net344),
    .X(net342));
 sg13g2_buf_1 fanout343 (.A(net344),
    .X(net343));
 sg13g2_buf_8 fanout344 (.A(net345),
    .X(net344));
 sg13g2_buf_1 fanout345 (.A(net350),
    .X(net345));
 sg13g2_buf_8 fanout346 (.A(net347),
    .X(net346));
 sg13g2_buf_8 fanout347 (.A(net349),
    .X(net347));
 sg13g2_buf_8 fanout348 (.A(net350),
    .X(net348));
 sg13g2_buf_1 fanout349 (.A(net350),
    .X(net349));
 sg13g2_buf_8 fanout350 (.A(net351),
    .X(net350));
 sg13g2_buf_8 fanout351 (.A(rst_n),
    .X(net351));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[0]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[1]),
    .X(net11));
 sg13g2_buf_2 input12 (.A(uio_in[2]),
    .X(net12));
 sg13g2_buf_2 input13 (.A(uio_in[4]),
    .X(net13));
 sg13g2_tielo tt_um_ebeam_pixel_core_14 (.L_LO(net14));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_4_0_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_1_0_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_4_2_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_3_0_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_4_4_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_5_0_clk));
 sg13g2_buf_1 clkload6 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_7_0_clk));
 sg13g2_buf_1 clkload8 (.A(clknet_4_8_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_11_0_clk));
 sg13g2_buf_1 clkload11 (.A(clknet_4_12_0_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_4_13_0_clk));
 sg13g2_buf_1 clkload13 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\cfg_wr_data_ff1[3] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold2 (.A(\cfg_wr_data_ff1[5] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold3 (.A(\cfg_wr_data_ff1[6] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold4 (.A(cfg_wr_toggle_ff1),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold5 (.A(\cfg_wr_data_ff1[4] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold6 (.A(\cfg_wr_addr_ff1[0] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold7 (.A(\cfg_wr_data_ff1[0] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold8 (.A(\cfg_wr_data_ff1[1] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold9 (.A(\cfg_wr_addr_ff1[1] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold10 (.A(\cfg_wr_data_ff1[2] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold11 (.A(\cfg_wr_data_ff1[7] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold12 (.A(\cfg_wr_addr_ff1[2] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold13 (.A(cfg_wr_toggle_ff2),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold14 (.A(\cfg_wr_data_ff2[7] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0169_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold16 (.A(\reg_absdiff_rdback[5] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold17 (.A(\reg_absdiff_rdback[1] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold18 (.A(\reg_absdiff_rdback[3] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold19 (.A(\reg_status[6] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold20 (.A(\reg_status[4] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold21 (.A(\reg_absdiff_rdback[7] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold22 (.A(\reg_status[5] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold23 (.A(\reg_absdiff_rdback[0] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold24 (.A(\reg_absdiff_rdback[6] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold25 (.A(\reg_edge_thr[7] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0185_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold27 (.A(\cfg_wr_data_ff2[2] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0180_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0016_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0354_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0172_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold32 (.A(\reg_absdiff_rdback[4] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold33 (.A(\cfg_wr_data_ff2[1] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0187_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold35 (.A(\cfg_wr_data_ff2[6] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0350_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0168_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold38 (.A(\cfg_wr_data_ff2[0] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0186_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold40 (.A(\reg_status[7] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold41 (.A(\reg_edge_thr[6] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0184_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold43 (.A(\cfg_wr_data_ff2[4] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0349_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0166_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold46 (.A(\reg_mode[5] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0249_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold48 (.A(\cfg_wr_data_ff2[3] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0173_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold50 (.A(\reg_absdiff_rdback[2] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold51 (.A(\reg_mode[7] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0251_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0019_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0360_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0181_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold56 (.A(\reg_mode[6] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0250_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold58 (.A(\reg_mode[4] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0248_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold60 (.A(\reg_mode[3] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0247_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold62 (.A(\reg_mode[2] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0246_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold64 (.A(\reg_contrast_thr[7] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0177_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold66 (.A(\prev_pixel[0] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0106_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold68 (.A(\reg_thresh[2] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0164_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold70 (.A(\prev_pixel[6] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0112_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold72 (.A(uo_out[3]),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0125_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold74 (.A(uo_out[0]),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0122_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold76 (.A(\prev_pixel[2] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0108_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold78 (.A(\prev_pixel[1] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0107_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold80 (.A(uo_out[1]),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0123_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold82 (.A(\prev_pixel[4] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0110_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold84 (.A(uo_out[7]),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0129_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold86 (.A(\reg_thresh[3] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0165_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold88 (.A(uo_out[6]),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0128_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold90 (.A(uo_out[5]),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0127_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold92 (.A(uo_out[2]),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0124_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold94 (.A(\reg_thresh[1] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0163_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold96 (.A(\prev_pixel[3] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0109_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold98 (.A(\pixel_q[6] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold99 (.A(\cfg_wr_data_ff2[5] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0167_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold101 (.A(\reg_edge_thr[5] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0183_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold103 (.A(\reg_contrast_thr[1] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0171_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold105 (.A(uo_out[4]),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0126_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold107 (.A(\reg_edge_thr[1] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0179_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold109 (.A(\reg_contrast_thr[0] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0170_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold111 (.A(\reg_contrast_thr[6] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0176_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold113 (.A(\reg_mode[1] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0245_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold115 (.A(\reg_contrast_thr[5] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0175_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold117 (.A(\reg_thresh[0] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0162_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold119 (.A(\reg_edge_thr[0] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0178_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold121 (.A(\prev_pixel[7] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0113_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold123 (.A(\reg_edge_thr[4] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0182_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold125 (.A(\pixel_q[0] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold126 (.A(\mean_q[5] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold127 (.A(\prev_pixel[5] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0111_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold129 (.A(\reg_contrast_thr[4] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0174_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold131 (.A(\mean_q[7] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0121_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold133 (.A(\reg_mode[0] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0244_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold135 (.A(\reg_alpha_shift[2] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0188_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold137 (.A(\mean_q[1] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0115_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold139 (.A(\mean_q[0] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold140 (.A(\pixel_q[1] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold141 (.A(\pixel_q[2] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold142 (.A(\mean_q[2] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold143 (.A(\pixel_q[4] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold144 (.A(\mean_q[6] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold145 (.A(\pixel_q[5] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold146 (.A(\mean_q[4] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold147 (.A(\mean_q[3] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold148 (.A(\pixel_q[7] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold149 (.A(\pixel_q[3] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold150 (.A(\reg_contrast_thr[7] ),
    .X(net404));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_fill_2 FILLER_0_245 ();
 sg13g2_decap_4 FILLER_0_256 ();
 sg13g2_fill_2 FILLER_0_260 ();
 sg13g2_fill_1 FILLER_0_271 ();
 sg13g2_decap_8 FILLER_0_277 ();
 sg13g2_decap_8 FILLER_0_284 ();
 sg13g2_decap_8 FILLER_0_291 ();
 sg13g2_decap_8 FILLER_0_298 ();
 sg13g2_decap_8 FILLER_0_305 ();
 sg13g2_decap_8 FILLER_0_312 ();
 sg13g2_decap_8 FILLER_0_319 ();
 sg13g2_decap_8 FILLER_0_326 ();
 sg13g2_decap_8 FILLER_0_333 ();
 sg13g2_decap_8 FILLER_0_340 ();
 sg13g2_decap_8 FILLER_0_347 ();
 sg13g2_decap_8 FILLER_0_354 ();
 sg13g2_decap_8 FILLER_0_361 ();
 sg13g2_decap_8 FILLER_0_368 ();
 sg13g2_decap_8 FILLER_0_375 ();
 sg13g2_decap_8 FILLER_0_382 ();
 sg13g2_decap_8 FILLER_0_389 ();
 sg13g2_decap_8 FILLER_0_396 ();
 sg13g2_decap_4 FILLER_0_403 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_4 FILLER_1_231 ();
 sg13g2_fill_1 FILLER_1_235 ();
 sg13g2_fill_2 FILLER_1_272 ();
 sg13g2_fill_1 FILLER_1_274 ();
 sg13g2_fill_2 FILLER_1_292 ();
 sg13g2_decap_4 FILLER_1_299 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_fill_1 FILLER_2_231 ();
 sg13g2_fill_2 FILLER_2_259 ();
 sg13g2_fill_2 FILLER_2_320 ();
 sg13g2_decap_8 FILLER_2_349 ();
 sg13g2_decap_8 FILLER_2_356 ();
 sg13g2_decap_8 FILLER_2_363 ();
 sg13g2_decap_8 FILLER_2_370 ();
 sg13g2_decap_8 FILLER_2_377 ();
 sg13g2_decap_8 FILLER_2_384 ();
 sg13g2_decap_8 FILLER_2_391 ();
 sg13g2_decap_8 FILLER_2_398 ();
 sg13g2_decap_4 FILLER_2_405 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_fill_1 FILLER_3_182 ();
 sg13g2_fill_2 FILLER_3_268 ();
 sg13g2_decap_4 FILLER_3_297 ();
 sg13g2_fill_2 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_312 ();
 sg13g2_fill_2 FILLER_3_319 ();
 sg13g2_decap_8 FILLER_3_352 ();
 sg13g2_decap_8 FILLER_3_359 ();
 sg13g2_decap_8 FILLER_3_366 ();
 sg13g2_decap_8 FILLER_3_373 ();
 sg13g2_decap_8 FILLER_3_380 ();
 sg13g2_decap_8 FILLER_3_387 ();
 sg13g2_decap_8 FILLER_3_394 ();
 sg13g2_decap_8 FILLER_3_401 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_fill_2 FILLER_4_189 ();
 sg13g2_fill_2 FILLER_4_231 ();
 sg13g2_fill_1 FILLER_4_246 ();
 sg13g2_fill_1 FILLER_4_260 ();
 sg13g2_decap_8 FILLER_4_289 ();
 sg13g2_decap_8 FILLER_4_296 ();
 sg13g2_fill_2 FILLER_4_303 ();
 sg13g2_fill_1 FILLER_4_305 ();
 sg13g2_decap_8 FILLER_4_311 ();
 sg13g2_decap_8 FILLER_4_318 ();
 sg13g2_decap_4 FILLER_4_325 ();
 sg13g2_fill_1 FILLER_4_329 ();
 sg13g2_fill_1 FILLER_4_334 ();
 sg13g2_decap_8 FILLER_4_340 ();
 sg13g2_decap_8 FILLER_4_347 ();
 sg13g2_decap_8 FILLER_4_354 ();
 sg13g2_decap_8 FILLER_4_361 ();
 sg13g2_decap_8 FILLER_4_368 ();
 sg13g2_decap_8 FILLER_4_375 ();
 sg13g2_decap_8 FILLER_4_382 ();
 sg13g2_decap_8 FILLER_4_389 ();
 sg13g2_decap_8 FILLER_4_396 ();
 sg13g2_decap_4 FILLER_4_403 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_4 FILLER_5_189 ();
 sg13g2_fill_2 FILLER_5_193 ();
 sg13g2_decap_4 FILLER_5_204 ();
 sg13g2_fill_2 FILLER_5_208 ();
 sg13g2_fill_1 FILLER_5_219 ();
 sg13g2_fill_2 FILLER_5_244 ();
 sg13g2_fill_1 FILLER_5_246 ();
 sg13g2_fill_2 FILLER_5_274 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_fill_2 FILLER_6_210 ();
 sg13g2_fill_1 FILLER_6_212 ();
 sg13g2_decap_4 FILLER_6_273 ();
 sg13g2_fill_2 FILLER_6_304 ();
 sg13g2_decap_8 FILLER_6_310 ();
 sg13g2_decap_8 FILLER_6_317 ();
 sg13g2_decap_4 FILLER_6_324 ();
 sg13g2_fill_1 FILLER_6_332 ();
 sg13g2_decap_8 FILLER_6_338 ();
 sg13g2_decap_4 FILLER_6_345 ();
 sg13g2_fill_1 FILLER_6_349 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_fill_1 FILLER_7_168 ();
 sg13g2_fill_1 FILLER_7_181 ();
 sg13g2_fill_2 FILLER_7_222 ();
 sg13g2_fill_2 FILLER_7_242 ();
 sg13g2_decap_8 FILLER_7_282 ();
 sg13g2_fill_2 FILLER_7_289 ();
 sg13g2_decap_4 FILLER_7_296 ();
 sg13g2_decap_4 FILLER_7_327 ();
 sg13g2_fill_1 FILLER_7_331 ();
 sg13g2_fill_2 FILLER_7_337 ();
 sg13g2_fill_1 FILLER_7_339 ();
 sg13g2_decap_8 FILLER_7_375 ();
 sg13g2_decap_8 FILLER_7_382 ();
 sg13g2_decap_8 FILLER_7_389 ();
 sg13g2_decap_8 FILLER_7_396 ();
 sg13g2_decap_4 FILLER_7_403 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_fill_2 FILLER_8_140 ();
 sg13g2_fill_1 FILLER_8_142 ();
 sg13g2_fill_1 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_4 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_309 ();
 sg13g2_decap_8 FILLER_8_316 ();
 sg13g2_decap_8 FILLER_8_323 ();
 sg13g2_decap_8 FILLER_8_330 ();
 sg13g2_fill_2 FILLER_8_337 ();
 sg13g2_fill_1 FILLER_8_339 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_fill_2 FILLER_9_161 ();
 sg13g2_fill_1 FILLER_9_163 ();
 sg13g2_decap_4 FILLER_9_198 ();
 sg13g2_fill_1 FILLER_9_202 ();
 sg13g2_decap_8 FILLER_9_212 ();
 sg13g2_fill_1 FILLER_9_219 ();
 sg13g2_fill_2 FILLER_9_243 ();
 sg13g2_fill_1 FILLER_9_245 ();
 sg13g2_fill_2 FILLER_9_267 ();
 sg13g2_fill_1 FILLER_9_269 ();
 sg13g2_decap_8 FILLER_9_356 ();
 sg13g2_decap_8 FILLER_9_363 ();
 sg13g2_decap_8 FILLER_9_370 ();
 sg13g2_decap_8 FILLER_9_377 ();
 sg13g2_decap_8 FILLER_9_384 ();
 sg13g2_decap_8 FILLER_9_391 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_fill_2 FILLER_10_147 ();
 sg13g2_fill_1 FILLER_10_185 ();
 sg13g2_decap_8 FILLER_10_191 ();
 sg13g2_decap_8 FILLER_10_198 ();
 sg13g2_decap_8 FILLER_10_205 ();
 sg13g2_decap_8 FILLER_10_212 ();
 sg13g2_decap_4 FILLER_10_219 ();
 sg13g2_fill_2 FILLER_10_223 ();
 sg13g2_fill_1 FILLER_10_300 ();
 sg13g2_fill_1 FILLER_10_328 ();
 sg13g2_decap_4 FILLER_10_343 ();
 sg13g2_fill_1 FILLER_10_347 ();
 sg13g2_decap_8 FILLER_10_375 ();
 sg13g2_decap_8 FILLER_10_382 ();
 sg13g2_decap_8 FILLER_10_389 ();
 sg13g2_decap_8 FILLER_10_396 ();
 sg13g2_decap_4 FILLER_10_403 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_fill_1 FILLER_11_166 ();
 sg13g2_decap_4 FILLER_11_175 ();
 sg13g2_fill_1 FILLER_11_179 ();
 sg13g2_decap_8 FILLER_11_185 ();
 sg13g2_decap_8 FILLER_11_192 ();
 sg13g2_decap_4 FILLER_11_199 ();
 sg13g2_decap_8 FILLER_11_239 ();
 sg13g2_decap_4 FILLER_11_246 ();
 sg13g2_fill_1 FILLER_11_260 ();
 sg13g2_fill_2 FILLER_11_270 ();
 sg13g2_decap_8 FILLER_11_285 ();
 sg13g2_decap_8 FILLER_11_292 ();
 sg13g2_decap_8 FILLER_11_299 ();
 sg13g2_decap_8 FILLER_11_314 ();
 sg13g2_decap_8 FILLER_11_321 ();
 sg13g2_fill_1 FILLER_11_328 ();
 sg13g2_decap_8 FILLER_11_333 ();
 sg13g2_decap_4 FILLER_11_340 ();
 sg13g2_fill_1 FILLER_11_344 ();
 sg13g2_decap_8 FILLER_11_376 ();
 sg13g2_decap_8 FILLER_11_383 ();
 sg13g2_decap_8 FILLER_11_390 ();
 sg13g2_decap_8 FILLER_11_397 ();
 sg13g2_decap_4 FILLER_11_404 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_4 FILLER_12_161 ();
 sg13g2_fill_2 FILLER_12_201 ();
 sg13g2_decap_8 FILLER_12_212 ();
 sg13g2_decap_4 FILLER_12_219 ();
 sg13g2_fill_1 FILLER_12_223 ();
 sg13g2_fill_1 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_258 ();
 sg13g2_fill_1 FILLER_12_265 ();
 sg13g2_decap_8 FILLER_12_293 ();
 sg13g2_decap_8 FILLER_12_300 ();
 sg13g2_decap_8 FILLER_12_312 ();
 sg13g2_decap_8 FILLER_12_319 ();
 sg13g2_decap_4 FILLER_12_326 ();
 sg13g2_fill_2 FILLER_12_330 ();
 sg13g2_decap_8 FILLER_12_345 ();
 sg13g2_fill_2 FILLER_12_352 ();
 sg13g2_fill_1 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_359 ();
 sg13g2_decap_8 FILLER_12_366 ();
 sg13g2_decap_8 FILLER_12_373 ();
 sg13g2_decap_8 FILLER_12_380 ();
 sg13g2_decap_8 FILLER_12_387 ();
 sg13g2_decap_8 FILLER_12_394 ();
 sg13g2_decap_8 FILLER_12_401 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_fill_2 FILLER_13_147 ();
 sg13g2_fill_1 FILLER_13_149 ();
 sg13g2_fill_2 FILLER_13_182 ();
 sg13g2_fill_1 FILLER_13_184 ();
 sg13g2_decap_4 FILLER_13_189 ();
 sg13g2_fill_1 FILLER_13_193 ();
 sg13g2_decap_8 FILLER_13_221 ();
 sg13g2_fill_1 FILLER_13_228 ();
 sg13g2_decap_8 FILLER_13_256 ();
 sg13g2_decap_8 FILLER_13_263 ();
 sg13g2_fill_2 FILLER_13_301 ();
 sg13g2_fill_1 FILLER_13_303 ();
 sg13g2_fill_2 FILLER_13_317 ();
 sg13g2_fill_1 FILLER_13_368 ();
 sg13g2_decap_8 FILLER_13_375 ();
 sg13g2_decap_8 FILLER_13_382 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_decap_4 FILLER_13_403 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_fill_2 FILLER_14_179 ();
 sg13g2_fill_2 FILLER_14_188 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_4 FILLER_14_224 ();
 sg13g2_decap_4 FILLER_14_247 ();
 sg13g2_decap_8 FILLER_14_269 ();
 sg13g2_decap_4 FILLER_14_276 ();
 sg13g2_fill_1 FILLER_14_284 ();
 sg13g2_fill_2 FILLER_14_321 ();
 sg13g2_fill_1 FILLER_14_323 ();
 sg13g2_decap_8 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_4 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_201 ();
 sg13g2_decap_8 FILLER_15_208 ();
 sg13g2_fill_1 FILLER_15_215 ();
 sg13g2_decap_8 FILLER_15_234 ();
 sg13g2_fill_1 FILLER_15_241 ();
 sg13g2_fill_2 FILLER_15_252 ();
 sg13g2_fill_1 FILLER_15_254 ();
 sg13g2_fill_2 FILLER_15_288 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_fill_2 FILLER_15_306 ();
 sg13g2_fill_1 FILLER_15_308 ();
 sg13g2_decap_4 FILLER_15_340 ();
 sg13g2_decap_8 FILLER_15_382 ();
 sg13g2_decap_8 FILLER_15_389 ();
 sg13g2_decap_8 FILLER_15_396 ();
 sg13g2_decap_4 FILLER_15_403 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_4 FILLER_16_154 ();
 sg13g2_decap_4 FILLER_16_161 ();
 sg13g2_fill_1 FILLER_16_165 ();
 sg13g2_fill_1 FILLER_16_172 ();
 sg13g2_decap_8 FILLER_16_183 ();
 sg13g2_fill_1 FILLER_16_190 ();
 sg13g2_fill_2 FILLER_16_218 ();
 sg13g2_fill_1 FILLER_16_220 ();
 sg13g2_fill_2 FILLER_16_286 ();
 sg13g2_decap_8 FILLER_16_328 ();
 sg13g2_decap_8 FILLER_16_335 ();
 sg13g2_decap_8 FILLER_16_342 ();
 sg13g2_decap_8 FILLER_16_349 ();
 sg13g2_decap_4 FILLER_16_356 ();
 sg13g2_decap_4 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_396 ();
 sg13g2_decap_4 FILLER_16_403 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_4 FILLER_17_147 ();
 sg13g2_decap_4 FILLER_17_204 ();
 sg13g2_decap_4 FILLER_17_240 ();
 sg13g2_decap_8 FILLER_17_314 ();
 sg13g2_decap_8 FILLER_17_321 ();
 sg13g2_fill_1 FILLER_17_328 ();
 sg13g2_decap_8 FILLER_17_356 ();
 sg13g2_decap_4 FILLER_17_363 ();
 sg13g2_fill_2 FILLER_17_367 ();
 sg13g2_decap_8 FILLER_17_383 ();
 sg13g2_decap_8 FILLER_17_390 ();
 sg13g2_decap_8 FILLER_17_397 ();
 sg13g2_decap_4 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_fill_1 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_173 ();
 sg13g2_decap_4 FILLER_18_180 ();
 sg13g2_fill_2 FILLER_18_184 ();
 sg13g2_fill_2 FILLER_18_199 ();
 sg13g2_fill_2 FILLER_18_206 ();
 sg13g2_decap_4 FILLER_18_221 ();
 sg13g2_fill_1 FILLER_18_285 ();
 sg13g2_fill_2 FILLER_18_313 ();
 sg13g2_fill_1 FILLER_18_315 ();
 sg13g2_decap_4 FILLER_18_352 ();
 sg13g2_fill_1 FILLER_18_356 ();
 sg13g2_fill_1 FILLER_18_362 ();
 sg13g2_decap_8 FILLER_18_381 ();
 sg13g2_decap_4 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_4 FILLER_19_154 ();
 sg13g2_fill_1 FILLER_19_158 ();
 sg13g2_decap_4 FILLER_19_171 ();
 sg13g2_decap_8 FILLER_19_180 ();
 sg13g2_decap_8 FILLER_19_187 ();
 sg13g2_decap_8 FILLER_19_194 ();
 sg13g2_decap_4 FILLER_19_201 ();
 sg13g2_fill_2 FILLER_19_205 ();
 sg13g2_decap_4 FILLER_19_222 ();
 sg13g2_fill_1 FILLER_19_226 ();
 sg13g2_fill_2 FILLER_19_263 ();
 sg13g2_fill_2 FILLER_19_289 ();
 sg13g2_decap_8 FILLER_19_303 ();
 sg13g2_decap_4 FILLER_19_310 ();
 sg13g2_fill_2 FILLER_19_351 ();
 sg13g2_fill_1 FILLER_19_359 ();
 sg13g2_fill_1 FILLER_19_372 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_4 FILLER_20_133 ();
 sg13g2_fill_1 FILLER_20_137 ();
 sg13g2_fill_2 FILLER_20_170 ();
 sg13g2_decap_4 FILLER_20_184 ();
 sg13g2_fill_1 FILLER_20_188 ();
 sg13g2_decap_4 FILLER_20_192 ();
 sg13g2_decap_8 FILLER_20_209 ();
 sg13g2_decap_8 FILLER_20_216 ();
 sg13g2_decap_8 FILLER_20_223 ();
 sg13g2_fill_1 FILLER_20_230 ();
 sg13g2_fill_1 FILLER_20_235 ();
 sg13g2_fill_1 FILLER_20_240 ();
 sg13g2_decap_8 FILLER_20_283 ();
 sg13g2_decap_8 FILLER_20_290 ();
 sg13g2_decap_8 FILLER_20_297 ();
 sg13g2_decap_8 FILLER_20_304 ();
 sg13g2_decap_8 FILLER_20_311 ();
 sg13g2_decap_8 FILLER_20_318 ();
 sg13g2_decap_4 FILLER_20_325 ();
 sg13g2_decap_8 FILLER_20_337 ();
 sg13g2_fill_2 FILLER_20_344 ();
 sg13g2_fill_2 FILLER_20_364 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_291 ();
 sg13g2_decap_4 FILLER_21_298 ();
 sg13g2_fill_2 FILLER_21_302 ();
 sg13g2_decap_8 FILLER_21_309 ();
 sg13g2_decap_4 FILLER_21_316 ();
 sg13g2_decap_8 FILLER_21_324 ();
 sg13g2_decap_8 FILLER_21_331 ();
 sg13g2_decap_8 FILLER_21_338 ();
 sg13g2_decap_8 FILLER_21_345 ();
 sg13g2_fill_1 FILLER_21_352 ();
 sg13g2_decap_8 FILLER_21_362 ();
 sg13g2_decap_8 FILLER_21_369 ();
 sg13g2_fill_2 FILLER_21_376 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_4 FILLER_22_133 ();
 sg13g2_fill_1 FILLER_22_137 ();
 sg13g2_fill_2 FILLER_22_170 ();
 sg13g2_decap_4 FILLER_22_176 ();
 sg13g2_fill_1 FILLER_22_180 ();
 sg13g2_fill_2 FILLER_22_212 ();
 sg13g2_fill_1 FILLER_22_226 ();
 sg13g2_fill_2 FILLER_22_236 ();
 sg13g2_fill_1 FILLER_22_238 ();
 sg13g2_fill_2 FILLER_22_243 ();
 sg13g2_decap_8 FILLER_22_298 ();
 sg13g2_decap_4 FILLER_22_310 ();
 sg13g2_fill_1 FILLER_22_314 ();
 sg13g2_fill_1 FILLER_22_342 ();
 sg13g2_decap_8 FILLER_22_361 ();
 sg13g2_decap_8 FILLER_22_368 ();
 sg13g2_decap_8 FILLER_22_375 ();
 sg13g2_fill_1 FILLER_22_382 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_4 FILLER_23_154 ();
 sg13g2_fill_2 FILLER_23_158 ();
 sg13g2_decap_8 FILLER_23_169 ();
 sg13g2_decap_4 FILLER_23_176 ();
 sg13g2_fill_1 FILLER_23_180 ();
 sg13g2_decap_4 FILLER_23_209 ();
 sg13g2_decap_8 FILLER_23_218 ();
 sg13g2_decap_4 FILLER_23_225 ();
 sg13g2_fill_2 FILLER_23_248 ();
 sg13g2_fill_1 FILLER_23_250 ();
 sg13g2_fill_1 FILLER_23_264 ();
 sg13g2_decap_4 FILLER_23_282 ();
 sg13g2_fill_2 FILLER_23_286 ();
 sg13g2_fill_1 FILLER_23_293 ();
 sg13g2_decap_4 FILLER_23_338 ();
 sg13g2_fill_2 FILLER_23_342 ();
 sg13g2_fill_2 FILLER_23_350 ();
 sg13g2_fill_1 FILLER_23_352 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_fill_1 FILLER_23_392 ();
 sg13g2_fill_1 FILLER_23_396 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_fill_2 FILLER_24_154 ();
 sg13g2_fill_1 FILLER_24_156 ();
 sg13g2_decap_4 FILLER_24_167 ();
 sg13g2_decap_8 FILLER_24_180 ();
 sg13g2_decap_8 FILLER_24_187 ();
 sg13g2_fill_2 FILLER_24_207 ();
 sg13g2_fill_2 FILLER_24_245 ();
 sg13g2_fill_1 FILLER_24_247 ();
 sg13g2_fill_2 FILLER_24_275 ();
 sg13g2_fill_2 FILLER_24_281 ();
 sg13g2_fill_1 FILLER_24_283 ();
 sg13g2_fill_1 FILLER_24_297 ();
 sg13g2_fill_1 FILLER_24_311 ();
 sg13g2_decap_4 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_375 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_4 FILLER_25_167 ();
 sg13g2_decap_8 FILLER_25_207 ();
 sg13g2_decap_8 FILLER_25_214 ();
 sg13g2_fill_1 FILLER_25_221 ();
 sg13g2_decap_4 FILLER_25_325 ();
 sg13g2_fill_1 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_334 ();
 sg13g2_decap_8 FILLER_25_341 ();
 sg13g2_decap_4 FILLER_25_348 ();
 sg13g2_decap_4 FILLER_25_359 ();
 sg13g2_fill_2 FILLER_25_363 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_4 FILLER_26_154 ();
 sg13g2_fill_1 FILLER_26_158 ();
 sg13g2_decap_8 FILLER_26_169 ();
 sg13g2_decap_8 FILLER_26_176 ();
 sg13g2_decap_8 FILLER_26_183 ();
 sg13g2_fill_2 FILLER_26_190 ();
 sg13g2_fill_2 FILLER_26_231 ();
 sg13g2_fill_1 FILLER_26_233 ();
 sg13g2_decap_8 FILLER_26_283 ();
 sg13g2_decap_8 FILLER_26_290 ();
 sg13g2_decap_8 FILLER_26_297 ();
 sg13g2_decap_8 FILLER_26_304 ();
 sg13g2_fill_1 FILLER_26_311 ();
 sg13g2_decap_8 FILLER_26_360 ();
 sg13g2_fill_1 FILLER_26_367 ();
 sg13g2_decap_4 FILLER_26_373 ();
 sg13g2_fill_2 FILLER_26_377 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_fill_1 FILLER_27_140 ();
 sg13g2_fill_2 FILLER_27_168 ();
 sg13g2_fill_2 FILLER_27_197 ();
 sg13g2_decap_8 FILLER_27_226 ();
 sg13g2_fill_2 FILLER_27_233 ();
 sg13g2_fill_1 FILLER_27_235 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_256 ();
 sg13g2_decap_8 FILLER_27_263 ();
 sg13g2_decap_4 FILLER_27_270 ();
 sg13g2_fill_2 FILLER_27_274 ();
 sg13g2_decap_8 FILLER_27_281 ();
 sg13g2_decap_8 FILLER_27_288 ();
 sg13g2_fill_2 FILLER_27_295 ();
 sg13g2_fill_1 FILLER_27_297 ();
 sg13g2_decap_8 FILLER_27_325 ();
 sg13g2_decap_8 FILLER_27_332 ();
 sg13g2_decap_8 FILLER_27_339 ();
 sg13g2_decap_4 FILLER_27_359 ();
 sg13g2_fill_2 FILLER_27_363 ();
 sg13g2_decap_8 FILLER_27_370 ();
 sg13g2_fill_2 FILLER_27_377 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_4 FILLER_28_140 ();
 sg13g2_decap_4 FILLER_28_181 ();
 sg13g2_fill_2 FILLER_28_185 ();
 sg13g2_fill_1 FILLER_28_217 ();
 sg13g2_fill_2 FILLER_28_246 ();
 sg13g2_fill_2 FILLER_28_279 ();
 sg13g2_fill_1 FILLER_28_281 ();
 sg13g2_fill_1 FILLER_28_309 ();
 sg13g2_fill_2 FILLER_28_315 ();
 sg13g2_fill_1 FILLER_28_317 ();
 sg13g2_decap_8 FILLER_28_351 ();
 sg13g2_fill_2 FILLER_28_363 ();
 sg13g2_decap_8 FILLER_28_400 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_fill_2 FILLER_29_154 ();
 sg13g2_fill_1 FILLER_29_156 ();
 sg13g2_decap_4 FILLER_29_167 ();
 sg13g2_decap_8 FILLER_29_198 ();
 sg13g2_decap_8 FILLER_29_205 ();
 sg13g2_fill_2 FILLER_29_212 ();
 sg13g2_decap_4 FILLER_29_236 ();
 sg13g2_fill_2 FILLER_29_267 ();
 sg13g2_decap_4 FILLER_29_296 ();
 sg13g2_fill_2 FILLER_29_300 ();
 sg13g2_fill_2 FILLER_29_311 ();
 sg13g2_fill_1 FILLER_29_313 ();
 sg13g2_decap_8 FILLER_29_368 ();
 sg13g2_decap_4 FILLER_29_375 ();
 sg13g2_fill_1 FILLER_29_379 ();
 sg13g2_decap_8 FILLER_29_384 ();
 sg13g2_decap_8 FILLER_29_391 ();
 sg13g2_decap_8 FILLER_29_398 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_fill_2 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_211 ();
 sg13g2_decap_8 FILLER_30_218 ();
 sg13g2_fill_2 FILLER_30_225 ();
 sg13g2_fill_1 FILLER_30_227 ();
 sg13g2_decap_8 FILLER_30_297 ();
 sg13g2_fill_2 FILLER_30_304 ();
 sg13g2_fill_1 FILLER_30_306 ();
 sg13g2_decap_8 FILLER_30_312 ();
 sg13g2_decap_8 FILLER_30_327 ();
 sg13g2_decap_4 FILLER_30_334 ();
 sg13g2_fill_1 FILLER_30_338 ();
 sg13g2_decap_8 FILLER_30_347 ();
 sg13g2_decap_4 FILLER_30_354 ();
 sg13g2_fill_2 FILLER_30_358 ();
 sg13g2_decap_4 FILLER_30_366 ();
 sg13g2_fill_2 FILLER_30_370 ();
 sg13g2_decap_4 FILLER_30_403 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_4 FILLER_31_133 ();
 sg13g2_fill_1 FILLER_31_137 ();
 sg13g2_decap_8 FILLER_31_171 ();
 sg13g2_decap_8 FILLER_31_178 ();
 sg13g2_decap_4 FILLER_31_185 ();
 sg13g2_fill_2 FILLER_31_225 ();
 sg13g2_fill_1 FILLER_31_227 ();
 sg13g2_fill_1 FILLER_31_238 ();
 sg13g2_fill_2 FILLER_31_276 ();
 sg13g2_fill_1 FILLER_31_278 ();
 sg13g2_fill_2 FILLER_31_306 ();
 sg13g2_decap_8 FILLER_31_326 ();
 sg13g2_fill_1 FILLER_31_333 ();
 sg13g2_fill_2 FILLER_31_361 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_fill_1 FILLER_32_140 ();
 sg13g2_fill_2 FILLER_32_228 ();
 sg13g2_fill_2 FILLER_32_262 ();
 sg13g2_fill_1 FILLER_32_264 ();
 sg13g2_decap_8 FILLER_32_287 ();
 sg13g2_decap_4 FILLER_32_294 ();
 sg13g2_fill_2 FILLER_32_298 ();
 sg13g2_decap_8 FILLER_32_327 ();
 sg13g2_decap_8 FILLER_32_334 ();
 sg13g2_decap_8 FILLER_32_341 ();
 sg13g2_decap_8 FILLER_32_348 ();
 sg13g2_decap_8 FILLER_32_355 ();
 sg13g2_decap_8 FILLER_32_362 ();
 sg13g2_decap_4 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_4 FILLER_33_147 ();
 sg13g2_fill_1 FILLER_33_151 ();
 sg13g2_fill_1 FILLER_33_155 ();
 sg13g2_fill_2 FILLER_33_175 ();
 sg13g2_fill_2 FILLER_33_194 ();
 sg13g2_fill_2 FILLER_33_236 ();
 sg13g2_decap_8 FILLER_33_310 ();
 sg13g2_decap_8 FILLER_33_317 ();
 sg13g2_fill_1 FILLER_33_324 ();
 sg13g2_decap_8 FILLER_33_352 ();
 sg13g2_decap_8 FILLER_33_359 ();
 sg13g2_decap_8 FILLER_33_366 ();
 sg13g2_decap_8 FILLER_33_373 ();
 sg13g2_decap_8 FILLER_33_383 ();
 sg13g2_fill_2 FILLER_33_390 ();
 sg13g2_fill_1 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_398 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_fill_2 FILLER_34_194 ();
 sg13g2_fill_1 FILLER_34_196 ();
 sg13g2_fill_1 FILLER_34_225 ();
 sg13g2_fill_1 FILLER_34_231 ();
 sg13g2_decap_4 FILLER_34_241 ();
 sg13g2_fill_1 FILLER_34_245 ();
 sg13g2_fill_2 FILLER_34_258 ();
 sg13g2_decap_8 FILLER_34_281 ();
 sg13g2_decap_4 FILLER_34_288 ();
 sg13g2_fill_1 FILLER_34_292 ();
 sg13g2_decap_4 FILLER_34_325 ();
 sg13g2_fill_1 FILLER_34_329 ();
 sg13g2_decap_8 FILLER_34_365 ();
 sg13g2_decap_8 FILLER_34_372 ();
 sg13g2_decap_8 FILLER_34_379 ();
 sg13g2_fill_2 FILLER_34_386 ();
 sg13g2_decap_4 FILLER_34_404 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_fill_2 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_162 ();
 sg13g2_fill_1 FILLER_35_169 ();
 sg13g2_fill_2 FILLER_35_223 ();
 sg13g2_fill_2 FILLER_35_244 ();
 sg13g2_fill_1 FILLER_35_246 ();
 sg13g2_fill_2 FILLER_35_260 ();
 sg13g2_fill_1 FILLER_35_262 ();
 sg13g2_fill_1 FILLER_35_272 ();
 sg13g2_fill_2 FILLER_35_291 ();
 sg13g2_fill_1 FILLER_35_293 ();
 sg13g2_decap_8 FILLER_35_302 ();
 sg13g2_decap_8 FILLER_35_323 ();
 sg13g2_decap_8 FILLER_35_330 ();
 sg13g2_fill_1 FILLER_35_355 ();
 sg13g2_decap_8 FILLER_35_360 ();
 sg13g2_decap_4 FILLER_35_367 ();
 sg13g2_decap_4 FILLER_35_377 ();
 sg13g2_fill_1 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_fill_2 FILLER_36_155 ();
 sg13g2_fill_1 FILLER_36_157 ();
 sg13g2_decap_8 FILLER_36_195 ();
 sg13g2_decap_8 FILLER_36_202 ();
 sg13g2_decap_8 FILLER_36_209 ();
 sg13g2_decap_8 FILLER_36_216 ();
 sg13g2_fill_2 FILLER_36_223 ();
 sg13g2_fill_2 FILLER_36_259 ();
 sg13g2_fill_1 FILLER_36_261 ();
 sg13g2_fill_2 FILLER_36_317 ();
 sg13g2_fill_1 FILLER_36_319 ();
 sg13g2_decap_4 FILLER_36_347 ();
 sg13g2_decap_4 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_4 FILLER_37_147 ();
 sg13g2_fill_2 FILLER_37_151 ();
 sg13g2_decap_8 FILLER_37_173 ();
 sg13g2_decap_8 FILLER_37_180 ();
 sg13g2_decap_8 FILLER_37_187 ();
 sg13g2_decap_8 FILLER_37_194 ();
 sg13g2_decap_8 FILLER_37_201 ();
 sg13g2_fill_2 FILLER_37_208 ();
 sg13g2_decap_8 FILLER_37_223 ();
 sg13g2_fill_2 FILLER_37_230 ();
 sg13g2_fill_2 FILLER_37_236 ();
 sg13g2_fill_2 FILLER_37_242 ();
 sg13g2_fill_1 FILLER_37_244 ();
 sg13g2_fill_2 FILLER_37_258 ();
 sg13g2_fill_1 FILLER_37_260 ();
 sg13g2_decap_8 FILLER_37_296 ();
 sg13g2_decap_8 FILLER_37_303 ();
 sg13g2_fill_2 FILLER_37_323 ();
 sg13g2_decap_4 FILLER_37_329 ();
 sg13g2_fill_2 FILLER_37_333 ();
 sg13g2_fill_1 FILLER_37_389 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_4 FILLER_38_133 ();
 sg13g2_fill_1 FILLER_38_137 ();
 sg13g2_fill_2 FILLER_38_165 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_222 ();
 sg13g2_decap_8 FILLER_38_229 ();
 sg13g2_fill_1 FILLER_38_236 ();
 sg13g2_fill_1 FILLER_38_250 ();
 sg13g2_decap_4 FILLER_38_294 ();
 sg13g2_fill_2 FILLER_38_298 ();
 sg13g2_fill_1 FILLER_38_318 ();
 sg13g2_decap_8 FILLER_38_346 ();
 sg13g2_decap_4 FILLER_38_353 ();
 sg13g2_decap_8 FILLER_38_366 ();
 sg13g2_fill_1 FILLER_38_373 ();
 sg13g2_decap_8 FILLER_38_380 ();
 sg13g2_decap_8 FILLER_38_387 ();
 sg13g2_decap_8 FILLER_38_394 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_4 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_164 ();
 sg13g2_fill_2 FILLER_39_171 ();
 sg13g2_fill_1 FILLER_39_173 ();
 sg13g2_fill_1 FILLER_39_339 ();
 sg13g2_decap_4 FILLER_39_344 ();
 sg13g2_fill_1 FILLER_39_353 ();
 sg13g2_decap_8 FILLER_39_402 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_decap_4 FILLER_40_147 ();
 sg13g2_fill_1 FILLER_40_151 ();
 sg13g2_fill_2 FILLER_40_162 ();
 sg13g2_fill_1 FILLER_40_164 ();
 sg13g2_fill_2 FILLER_40_178 ();
 sg13g2_fill_1 FILLER_40_180 ();
 sg13g2_fill_2 FILLER_40_234 ();
 sg13g2_fill_1 FILLER_40_301 ();
 sg13g2_decap_8 FILLER_40_306 ();
 sg13g2_decap_4 FILLER_40_313 ();
 sg13g2_fill_1 FILLER_40_317 ();
 sg13g2_decap_8 FILLER_40_331 ();
 sg13g2_decap_8 FILLER_40_338 ();
 sg13g2_decap_8 FILLER_40_345 ();
 sg13g2_decap_8 FILLER_40_352 ();
 sg13g2_decap_4 FILLER_40_363 ();
 sg13g2_fill_2 FILLER_40_367 ();
 sg13g2_fill_1 FILLER_40_386 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_8 FILLER_41_147 ();
 sg13g2_decap_4 FILLER_41_154 ();
 sg13g2_fill_2 FILLER_41_158 ();
 sg13g2_fill_1 FILLER_41_187 ();
 sg13g2_fill_2 FILLER_41_225 ();
 sg13g2_fill_1 FILLER_41_259 ();
 sg13g2_fill_1 FILLER_41_265 ();
 sg13g2_decap_8 FILLER_41_280 ();
 sg13g2_fill_2 FILLER_41_314 ();
 sg13g2_fill_1 FILLER_41_316 ();
 sg13g2_decap_8 FILLER_41_326 ();
 sg13g2_fill_1 FILLER_41_346 ();
 sg13g2_decap_4 FILLER_41_374 ();
 sg13g2_fill_1 FILLER_41_378 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_decap_8 FILLER_42_154 ();
 sg13g2_fill_1 FILLER_42_161 ();
 sg13g2_decap_8 FILLER_42_189 ();
 sg13g2_fill_1 FILLER_42_224 ();
 sg13g2_fill_1 FILLER_42_260 ();
 sg13g2_decap_8 FILLER_42_299 ();
 sg13g2_decap_8 FILLER_42_306 ();
 sg13g2_fill_2 FILLER_42_313 ();
 sg13g2_fill_1 FILLER_42_315 ();
 sg13g2_fill_2 FILLER_42_321 ();
 sg13g2_fill_1 FILLER_42_323 ();
 sg13g2_decap_8 FILLER_42_360 ();
 sg13g2_decap_8 FILLER_42_367 ();
 sg13g2_decap_8 FILLER_42_401 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_decap_8 FILLER_43_133 ();
 sg13g2_decap_8 FILLER_43_140 ();
 sg13g2_decap_8 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_154 ();
 sg13g2_decap_8 FILLER_43_161 ();
 sg13g2_decap_8 FILLER_43_168 ();
 sg13g2_decap_8 FILLER_43_175 ();
 sg13g2_decap_8 FILLER_43_182 ();
 sg13g2_fill_2 FILLER_43_189 ();
 sg13g2_fill_1 FILLER_43_191 ();
 sg13g2_decap_4 FILLER_43_206 ();
 sg13g2_decap_4 FILLER_43_214 ();
 sg13g2_decap_4 FILLER_43_227 ();
 sg13g2_fill_1 FILLER_43_231 ();
 sg13g2_decap_4 FILLER_43_250 ();
 sg13g2_fill_2 FILLER_43_269 ();
 sg13g2_fill_1 FILLER_43_271 ();
 sg13g2_decap_8 FILLER_43_300 ();
 sg13g2_fill_1 FILLER_43_307 ();
 sg13g2_fill_2 FILLER_43_345 ();
 sg13g2_decap_8 FILLER_43_360 ();
 sg13g2_fill_1 FILLER_43_367 ();
 sg13g2_decap_4 FILLER_43_373 ();
 sg13g2_fill_2 FILLER_43_377 ();
 sg13g2_decap_4 FILLER_43_383 ();
 sg13g2_fill_2 FILLER_43_387 ();
 sg13g2_decap_8 FILLER_43_393 ();
 sg13g2_decap_8 FILLER_43_400 ();
 sg13g2_fill_2 FILLER_43_407 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_decap_8 FILLER_44_133 ();
 sg13g2_decap_8 FILLER_44_140 ();
 sg13g2_decap_8 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_154 ();
 sg13g2_decap_8 FILLER_44_161 ();
 sg13g2_fill_1 FILLER_44_168 ();
 sg13g2_fill_2 FILLER_44_269 ();
 sg13g2_fill_2 FILLER_44_280 ();
 sg13g2_decap_8 FILLER_44_304 ();
 sg13g2_decap_8 FILLER_44_311 ();
 sg13g2_decap_8 FILLER_44_322 ();
 sg13g2_decap_8 FILLER_44_333 ();
 sg13g2_fill_1 FILLER_44_340 ();
 sg13g2_fill_1 FILLER_44_381 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_decap_8 FILLER_45_133 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_decap_8 FILLER_45_147 ();
 sg13g2_decap_8 FILLER_45_154 ();
 sg13g2_decap_8 FILLER_45_161 ();
 sg13g2_decap_8 FILLER_45_181 ();
 sg13g2_decap_4 FILLER_45_211 ();
 sg13g2_fill_1 FILLER_45_215 ();
 sg13g2_decap_4 FILLER_45_295 ();
 sg13g2_decap_8 FILLER_45_308 ();
 sg13g2_decap_8 FILLER_45_315 ();
 sg13g2_fill_2 FILLER_45_322 ();
 sg13g2_decap_8 FILLER_45_337 ();
 sg13g2_decap_4 FILLER_45_344 ();
 sg13g2_fill_2 FILLER_45_352 ();
 sg13g2_decap_8 FILLER_45_385 ();
 sg13g2_fill_1 FILLER_45_392 ();
 sg13g2_decap_8 FILLER_45_397 ();
 sg13g2_decap_4 FILLER_45_404 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_8 FILLER_46_133 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_decap_8 FILLER_46_147 ();
 sg13g2_decap_8 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_161 ();
 sg13g2_decap_8 FILLER_46_168 ();
 sg13g2_decap_4 FILLER_46_190 ();
 sg13g2_fill_1 FILLER_46_194 ();
 sg13g2_decap_4 FILLER_46_200 ();
 sg13g2_fill_1 FILLER_46_204 ();
 sg13g2_decap_8 FILLER_46_210 ();
 sg13g2_decap_4 FILLER_46_217 ();
 sg13g2_fill_2 FILLER_46_240 ();
 sg13g2_fill_1 FILLER_46_242 ();
 sg13g2_fill_2 FILLER_46_338 ();
 sg13g2_decap_4 FILLER_46_380 ();
 sg13g2_fill_1 FILLER_46_384 ();
 sg13g2_fill_1 FILLER_46_395 ();
 sg13g2_fill_2 FILLER_46_406 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_fill_2 FILLER_47_161 ();
 sg13g2_fill_1 FILLER_47_222 ();
 sg13g2_decap_4 FILLER_47_232 ();
 sg13g2_fill_2 FILLER_47_245 ();
 sg13g2_fill_2 FILLER_47_325 ();
 sg13g2_fill_1 FILLER_47_327 ();
 sg13g2_fill_2 FILLER_47_360 ();
 sg13g2_fill_1 FILLER_47_362 ();
 sg13g2_decap_8 FILLER_47_367 ();
 sg13g2_decap_8 FILLER_47_374 ();
 sg13g2_fill_1 FILLER_47_381 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_4 FILLER_48_147 ();
 sg13g2_fill_2 FILLER_48_151 ();
 sg13g2_fill_1 FILLER_48_181 ();
 sg13g2_fill_1 FILLER_48_212 ();
 sg13g2_decap_4 FILLER_48_229 ();
 sg13g2_fill_2 FILLER_48_233 ();
 sg13g2_decap_8 FILLER_48_240 ();
 sg13g2_fill_2 FILLER_48_247 ();
 sg13g2_decap_4 FILLER_48_258 ();
 sg13g2_fill_2 FILLER_48_262 ();
 sg13g2_decap_8 FILLER_48_349 ();
 sg13g2_decap_8 FILLER_48_356 ();
 sg13g2_decap_8 FILLER_48_363 ();
 sg13g2_decap_8 FILLER_48_370 ();
 sg13g2_decap_4 FILLER_48_377 ();
 sg13g2_fill_1 FILLER_48_381 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_decap_8 FILLER_49_133 ();
 sg13g2_decap_8 FILLER_49_140 ();
 sg13g2_decap_4 FILLER_49_147 ();
 sg13g2_fill_2 FILLER_49_151 ();
 sg13g2_fill_1 FILLER_49_216 ();
 sg13g2_decap_4 FILLER_49_228 ();
 sg13g2_fill_1 FILLER_49_253 ();
 sg13g2_fill_2 FILLER_49_260 ();
 sg13g2_fill_1 FILLER_49_270 ();
 sg13g2_fill_1 FILLER_49_298 ();
 sg13g2_fill_1 FILLER_49_315 ();
 sg13g2_decap_4 FILLER_49_330 ();
 sg13g2_fill_2 FILLER_49_334 ();
 sg13g2_decap_8 FILLER_49_341 ();
 sg13g2_decap_8 FILLER_49_348 ();
 sg13g2_decap_8 FILLER_49_355 ();
 sg13g2_fill_2 FILLER_49_362 ();
 sg13g2_decap_8 FILLER_49_368 ();
 sg13g2_decap_8 FILLER_49_375 ();
 sg13g2_decap_4 FILLER_49_382 ();
 sg13g2_fill_2 FILLER_49_406 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_98 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_decap_8 FILLER_50_112 ();
 sg13g2_decap_8 FILLER_50_119 ();
 sg13g2_decap_8 FILLER_50_126 ();
 sg13g2_decap_8 FILLER_50_133 ();
 sg13g2_decap_8 FILLER_50_140 ();
 sg13g2_decap_8 FILLER_50_147 ();
 sg13g2_decap_4 FILLER_50_154 ();
 sg13g2_fill_2 FILLER_50_233 ();
 sg13g2_fill_1 FILLER_50_235 ();
 sg13g2_fill_1 FILLER_50_292 ();
 sg13g2_fill_1 FILLER_50_321 ();
 sg13g2_decap_4 FILLER_50_327 ();
 sg13g2_fill_1 FILLER_50_358 ();
 sg13g2_decap_8 FILLER_50_386 ();
 sg13g2_fill_2 FILLER_50_393 ();
 sg13g2_decap_8 FILLER_50_399 ();
 sg13g2_fill_2 FILLER_50_406 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_98 ();
 sg13g2_decap_8 FILLER_51_105 ();
 sg13g2_decap_8 FILLER_51_112 ();
 sg13g2_decap_8 FILLER_51_119 ();
 sg13g2_decap_8 FILLER_51_126 ();
 sg13g2_decap_8 FILLER_51_133 ();
 sg13g2_decap_8 FILLER_51_140 ();
 sg13g2_decap_8 FILLER_51_147 ();
 sg13g2_decap_8 FILLER_51_154 ();
 sg13g2_decap_4 FILLER_51_161 ();
 sg13g2_fill_2 FILLER_51_192 ();
 sg13g2_fill_1 FILLER_51_214 ();
 sg13g2_fill_1 FILLER_51_242 ();
 sg13g2_fill_1 FILLER_51_274 ();
 sg13g2_decap_8 FILLER_51_317 ();
 sg13g2_fill_1 FILLER_51_324 ();
 sg13g2_fill_2 FILLER_51_366 ();
 sg13g2_fill_1 FILLER_51_368 ();
 sg13g2_decap_8 FILLER_51_396 ();
 sg13g2_decap_4 FILLER_51_403 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_decap_8 FILLER_52_112 ();
 sg13g2_decap_8 FILLER_52_119 ();
 sg13g2_decap_8 FILLER_52_126 ();
 sg13g2_decap_8 FILLER_52_133 ();
 sg13g2_decap_8 FILLER_52_140 ();
 sg13g2_decap_8 FILLER_52_147 ();
 sg13g2_decap_8 FILLER_52_154 ();
 sg13g2_decap_4 FILLER_52_161 ();
 sg13g2_fill_2 FILLER_52_165 ();
 sg13g2_fill_2 FILLER_52_234 ();
 sg13g2_fill_2 FILLER_52_246 ();
 sg13g2_fill_1 FILLER_52_270 ();
 sg13g2_fill_2 FILLER_52_279 ();
 sg13g2_fill_1 FILLER_52_300 ();
 sg13g2_decap_8 FILLER_52_314 ();
 sg13g2_decap_8 FILLER_52_321 ();
 sg13g2_decap_8 FILLER_52_328 ();
 sg13g2_fill_1 FILLER_52_335 ();
 sg13g2_decap_8 FILLER_52_340 ();
 sg13g2_decap_8 FILLER_52_347 ();
 sg13g2_fill_2 FILLER_52_354 ();
 sg13g2_fill_1 FILLER_52_383 ();
 sg13g2_decap_8 FILLER_52_388 ();
 sg13g2_decap_8 FILLER_52_395 ();
 sg13g2_decap_8 FILLER_52_402 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_8 FILLER_53_105 ();
 sg13g2_decap_8 FILLER_53_112 ();
 sg13g2_decap_8 FILLER_53_119 ();
 sg13g2_decap_8 FILLER_53_126 ();
 sg13g2_decap_8 FILLER_53_133 ();
 sg13g2_decap_8 FILLER_53_140 ();
 sg13g2_decap_8 FILLER_53_147 ();
 sg13g2_decap_8 FILLER_53_154 ();
 sg13g2_fill_1 FILLER_53_161 ();
 sg13g2_fill_2 FILLER_53_190 ();
 sg13g2_fill_2 FILLER_53_212 ();
 sg13g2_fill_1 FILLER_53_214 ();
 sg13g2_decap_4 FILLER_53_220 ();
 sg13g2_fill_1 FILLER_53_224 ();
 sg13g2_decap_8 FILLER_53_233 ();
 sg13g2_decap_4 FILLER_53_240 ();
 sg13g2_fill_2 FILLER_53_244 ();
 sg13g2_fill_1 FILLER_53_249 ();
 sg13g2_decap_8 FILLER_53_259 ();
 sg13g2_decap_8 FILLER_53_266 ();
 sg13g2_fill_2 FILLER_53_273 ();
 sg13g2_decap_4 FILLER_53_289 ();
 sg13g2_decap_8 FILLER_53_334 ();
 sg13g2_decap_8 FILLER_53_341 ();
 sg13g2_decap_8 FILLER_53_348 ();
 sg13g2_decap_4 FILLER_53_355 ();
 sg13g2_fill_2 FILLER_53_359 ();
 sg13g2_decap_8 FILLER_53_365 ();
 sg13g2_fill_2 FILLER_53_372 ();
 sg13g2_fill_1 FILLER_53_378 ();
 sg13g2_fill_2 FILLER_53_406 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_decap_8 FILLER_54_105 ();
 sg13g2_decap_8 FILLER_54_112 ();
 sg13g2_decap_8 FILLER_54_119 ();
 sg13g2_decap_8 FILLER_54_126 ();
 sg13g2_decap_8 FILLER_54_133 ();
 sg13g2_decap_8 FILLER_54_140 ();
 sg13g2_decap_4 FILLER_54_147 ();
 sg13g2_fill_2 FILLER_54_179 ();
 sg13g2_fill_1 FILLER_54_181 ();
 sg13g2_decap_4 FILLER_54_195 ();
 sg13g2_decap_8 FILLER_54_208 ();
 sg13g2_decap_8 FILLER_54_215 ();
 sg13g2_decap_8 FILLER_54_222 ();
 sg13g2_fill_2 FILLER_54_229 ();
 sg13g2_fill_1 FILLER_54_231 ();
 sg13g2_decap_8 FILLER_54_240 ();
 sg13g2_fill_2 FILLER_54_247 ();
 sg13g2_decap_8 FILLER_54_259 ();
 sg13g2_fill_2 FILLER_54_266 ();
 sg13g2_decap_4 FILLER_54_321 ();
 sg13g2_fill_1 FILLER_54_325 ();
 sg13g2_decap_8 FILLER_54_372 ();
 sg13g2_decap_8 FILLER_54_379 ();
 sg13g2_decap_8 FILLER_54_386 ();
 sg13g2_fill_2 FILLER_54_393 ();
 sg13g2_fill_1 FILLER_54_395 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_98 ();
 sg13g2_decap_8 FILLER_55_105 ();
 sg13g2_decap_8 FILLER_55_112 ();
 sg13g2_decap_8 FILLER_55_119 ();
 sg13g2_decap_8 FILLER_55_126 ();
 sg13g2_decap_8 FILLER_55_133 ();
 sg13g2_decap_8 FILLER_55_140 ();
 sg13g2_decap_8 FILLER_55_147 ();
 sg13g2_decap_4 FILLER_55_191 ();
 sg13g2_fill_2 FILLER_55_213 ();
 sg13g2_fill_1 FILLER_55_220 ();
 sg13g2_decap_8 FILLER_55_225 ();
 sg13g2_decap_8 FILLER_55_232 ();
 sg13g2_decap_8 FILLER_55_239 ();
 sg13g2_decap_8 FILLER_55_246 ();
 sg13g2_fill_2 FILLER_55_253 ();
 sg13g2_decap_8 FILLER_55_270 ();
 sg13g2_fill_2 FILLER_55_277 ();
 sg13g2_fill_1 FILLER_55_294 ();
 sg13g2_decap_4 FILLER_55_322 ();
 sg13g2_fill_2 FILLER_55_353 ();
 sg13g2_fill_1 FILLER_55_355 ();
 sg13g2_decap_8 FILLER_55_361 ();
 sg13g2_fill_2 FILLER_55_368 ();
 sg13g2_fill_1 FILLER_55_370 ();
 sg13g2_fill_2 FILLER_55_406 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_decap_8 FILLER_56_105 ();
 sg13g2_decap_8 FILLER_56_112 ();
 sg13g2_decap_8 FILLER_56_119 ();
 sg13g2_decap_8 FILLER_56_126 ();
 sg13g2_decap_8 FILLER_56_133 ();
 sg13g2_decap_8 FILLER_56_140 ();
 sg13g2_decap_8 FILLER_56_147 ();
 sg13g2_decap_8 FILLER_56_154 ();
 sg13g2_fill_2 FILLER_56_175 ();
 sg13g2_decap_4 FILLER_56_218 ();
 sg13g2_decap_8 FILLER_56_238 ();
 sg13g2_fill_2 FILLER_56_245 ();
 sg13g2_decap_8 FILLER_56_260 ();
 sg13g2_decap_8 FILLER_56_267 ();
 sg13g2_decap_8 FILLER_56_297 ();
 sg13g2_fill_2 FILLER_56_324 ();
 sg13g2_fill_1 FILLER_56_326 ();
 sg13g2_decap_4 FILLER_56_335 ();
 sg13g2_fill_1 FILLER_56_339 ();
 sg13g2_decap_8 FILLER_56_344 ();
 sg13g2_decap_8 FILLER_56_351 ();
 sg13g2_decap_8 FILLER_56_358 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_98 ();
 sg13g2_decap_8 FILLER_57_105 ();
 sg13g2_decap_8 FILLER_57_112 ();
 sg13g2_decap_8 FILLER_57_119 ();
 sg13g2_decap_8 FILLER_57_126 ();
 sg13g2_decap_8 FILLER_57_133 ();
 sg13g2_decap_8 FILLER_57_140 ();
 sg13g2_decap_8 FILLER_57_147 ();
 sg13g2_decap_8 FILLER_57_154 ();
 sg13g2_decap_8 FILLER_57_161 ();
 sg13g2_decap_4 FILLER_57_168 ();
 sg13g2_fill_1 FILLER_57_181 ();
 sg13g2_fill_1 FILLER_57_194 ();
 sg13g2_fill_2 FILLER_57_204 ();
 sg13g2_fill_1 FILLER_57_206 ();
 sg13g2_fill_1 FILLER_57_233 ();
 sg13g2_decap_4 FILLER_57_272 ();
 sg13g2_fill_2 FILLER_57_276 ();
 sg13g2_decap_8 FILLER_57_290 ();
 sg13g2_decap_4 FILLER_57_297 ();
 sg13g2_fill_2 FILLER_57_310 ();
 sg13g2_decap_8 FILLER_57_316 ();
 sg13g2_decap_8 FILLER_57_350 ();
 sg13g2_fill_2 FILLER_57_357 ();
 sg13g2_fill_1 FILLER_57_359 ();
 sg13g2_fill_2 FILLER_57_387 ();
 sg13g2_fill_1 FILLER_57_389 ();
 sg13g2_decap_4 FILLER_57_403 ();
 sg13g2_fill_2 FILLER_57_407 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_decap_8 FILLER_58_112 ();
 sg13g2_decap_8 FILLER_58_119 ();
 sg13g2_decap_8 FILLER_58_126 ();
 sg13g2_decap_8 FILLER_58_133 ();
 sg13g2_decap_8 FILLER_58_140 ();
 sg13g2_decap_4 FILLER_58_147 ();
 sg13g2_fill_2 FILLER_58_151 ();
 sg13g2_fill_1 FILLER_58_213 ();
 sg13g2_fill_2 FILLER_58_220 ();
 sg13g2_fill_1 FILLER_58_222 ();
 sg13g2_fill_2 FILLER_58_228 ();
 sg13g2_decap_4 FILLER_58_281 ();
 sg13g2_decap_8 FILLER_58_313 ();
 sg13g2_fill_1 FILLER_58_320 ();
 sg13g2_decap_4 FILLER_58_348 ();
 sg13g2_decap_8 FILLER_58_357 ();
 sg13g2_fill_1 FILLER_58_364 ();
 sg13g2_fill_1 FILLER_58_369 ();
 sg13g2_decap_8 FILLER_58_374 ();
 sg13g2_decap_8 FILLER_58_381 ();
 sg13g2_fill_2 FILLER_58_394 ();
 sg13g2_fill_1 FILLER_58_396 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_decap_8 FILLER_59_105 ();
 sg13g2_decap_8 FILLER_59_112 ();
 sg13g2_decap_8 FILLER_59_119 ();
 sg13g2_decap_8 FILLER_59_126 ();
 sg13g2_decap_8 FILLER_59_133 ();
 sg13g2_decap_8 FILLER_59_140 ();
 sg13g2_decap_8 FILLER_59_147 ();
 sg13g2_decap_8 FILLER_59_154 ();
 sg13g2_decap_8 FILLER_59_161 ();
 sg13g2_decap_8 FILLER_59_168 ();
 sg13g2_decap_4 FILLER_59_175 ();
 sg13g2_fill_1 FILLER_59_206 ();
 sg13g2_fill_2 FILLER_59_215 ();
 sg13g2_fill_2 FILLER_59_233 ();
 sg13g2_decap_4 FILLER_59_243 ();
 sg13g2_decap_8 FILLER_59_318 ();
 sg13g2_fill_1 FILLER_59_325 ();
 sg13g2_decap_8 FILLER_59_330 ();
 sg13g2_decap_8 FILLER_59_337 ();
 sg13g2_decap_4 FILLER_59_344 ();
 sg13g2_fill_1 FILLER_59_348 ();
 sg13g2_fill_2 FILLER_59_354 ();
 sg13g2_fill_1 FILLER_59_356 ();
 sg13g2_decap_4 FILLER_59_384 ();
 sg13g2_fill_1 FILLER_59_388 ();
 sg13g2_decap_4 FILLER_59_404 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_98 ();
 sg13g2_decap_8 FILLER_60_105 ();
 sg13g2_decap_8 FILLER_60_112 ();
 sg13g2_decap_8 FILLER_60_119 ();
 sg13g2_decap_8 FILLER_60_126 ();
 sg13g2_decap_8 FILLER_60_133 ();
 sg13g2_decap_8 FILLER_60_140 ();
 sg13g2_decap_8 FILLER_60_147 ();
 sg13g2_decap_4 FILLER_60_154 ();
 sg13g2_fill_2 FILLER_60_158 ();
 sg13g2_fill_2 FILLER_60_187 ();
 sg13g2_decap_4 FILLER_60_227 ();
 sg13g2_decap_4 FILLER_60_235 ();
 sg13g2_fill_2 FILLER_60_239 ();
 sg13g2_decap_8 FILLER_60_259 ();
 sg13g2_decap_8 FILLER_60_266 ();
 sg13g2_decap_8 FILLER_60_273 ();
 sg13g2_decap_4 FILLER_60_280 ();
 sg13g2_fill_2 FILLER_60_347 ();
 sg13g2_fill_1 FILLER_60_349 ();
 sg13g2_decap_8 FILLER_60_355 ();
 sg13g2_decap_8 FILLER_60_370 ();
 sg13g2_decap_8 FILLER_60_377 ();
 sg13g2_fill_2 FILLER_60_384 ();
 sg13g2_decap_4 FILLER_60_392 ();
 sg13g2_fill_1 FILLER_60_396 ();
 sg13g2_decap_4 FILLER_60_403 ();
 sg13g2_fill_2 FILLER_60_407 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_8 FILLER_61_91 ();
 sg13g2_decap_8 FILLER_61_98 ();
 sg13g2_decap_8 FILLER_61_105 ();
 sg13g2_decap_8 FILLER_61_112 ();
 sg13g2_decap_8 FILLER_61_119 ();
 sg13g2_decap_8 FILLER_61_126 ();
 sg13g2_decap_8 FILLER_61_133 ();
 sg13g2_decap_8 FILLER_61_140 ();
 sg13g2_decap_8 FILLER_61_147 ();
 sg13g2_fill_1 FILLER_61_182 ();
 sg13g2_fill_2 FILLER_61_198 ();
 sg13g2_fill_1 FILLER_61_200 ();
 sg13g2_decap_8 FILLER_61_214 ();
 sg13g2_decap_8 FILLER_61_221 ();
 sg13g2_fill_1 FILLER_61_228 ();
 sg13g2_fill_1 FILLER_61_273 ();
 sg13g2_decap_4 FILLER_61_279 ();
 sg13g2_fill_2 FILLER_61_283 ();
 sg13g2_decap_8 FILLER_61_293 ();
 sg13g2_fill_2 FILLER_61_300 ();
 sg13g2_fill_1 FILLER_61_302 ();
 sg13g2_decap_8 FILLER_61_309 ();
 sg13g2_fill_1 FILLER_61_316 ();
 sg13g2_fill_2 FILLER_61_322 ();
 sg13g2_fill_1 FILLER_61_324 ();
 sg13g2_decap_4 FILLER_61_356 ();
 sg13g2_decap_8 FILLER_61_387 ();
 sg13g2_decap_8 FILLER_61_394 ();
 sg13g2_decap_8 FILLER_61_401 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_8 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_decap_8 FILLER_62_112 ();
 sg13g2_decap_8 FILLER_62_119 ();
 sg13g2_decap_8 FILLER_62_126 ();
 sg13g2_decap_8 FILLER_62_133 ();
 sg13g2_decap_8 FILLER_62_140 ();
 sg13g2_decap_8 FILLER_62_147 ();
 sg13g2_decap_4 FILLER_62_154 ();
 sg13g2_fill_1 FILLER_62_158 ();
 sg13g2_fill_1 FILLER_62_172 ();
 sg13g2_fill_1 FILLER_62_191 ();
 sg13g2_fill_2 FILLER_62_205 ();
 sg13g2_fill_1 FILLER_62_222 ();
 sg13g2_fill_2 FILLER_62_236 ();
 sg13g2_fill_2 FILLER_62_246 ();
 sg13g2_fill_1 FILLER_62_258 ();
 sg13g2_fill_1 FILLER_62_267 ();
 sg13g2_fill_1 FILLER_62_281 ();
 sg13g2_decap_8 FILLER_62_298 ();
 sg13g2_decap_8 FILLER_62_305 ();
 sg13g2_decap_8 FILLER_62_312 ();
 sg13g2_decap_8 FILLER_62_319 ();
 sg13g2_decap_8 FILLER_62_326 ();
 sg13g2_fill_1 FILLER_62_333 ();
 sg13g2_fill_1 FILLER_62_338 ();
 sg13g2_fill_2 FILLER_62_376 ();
 sg13g2_decap_4 FILLER_62_405 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_decap_8 FILLER_63_105 ();
 sg13g2_decap_8 FILLER_63_112 ();
 sg13g2_decap_8 FILLER_63_119 ();
 sg13g2_decap_8 FILLER_63_126 ();
 sg13g2_decap_8 FILLER_63_133 ();
 sg13g2_decap_8 FILLER_63_140 ();
 sg13g2_decap_8 FILLER_63_147 ();
 sg13g2_decap_8 FILLER_63_154 ();
 sg13g2_decap_8 FILLER_63_161 ();
 sg13g2_fill_1 FILLER_63_168 ();
 sg13g2_fill_2 FILLER_63_192 ();
 sg13g2_fill_1 FILLER_63_194 ();
 sg13g2_decap_8 FILLER_63_226 ();
 sg13g2_decap_8 FILLER_63_233 ();
 sg13g2_decap_8 FILLER_63_240 ();
 sg13g2_decap_8 FILLER_63_247 ();
 sg13g2_decap_8 FILLER_63_254 ();
 sg13g2_decap_4 FILLER_63_261 ();
 sg13g2_fill_1 FILLER_63_273 ();
 sg13g2_fill_2 FILLER_63_288 ();
 sg13g2_decap_8 FILLER_63_323 ();
 sg13g2_decap_8 FILLER_63_330 ();
 sg13g2_decap_8 FILLER_63_337 ();
 sg13g2_decap_8 FILLER_63_348 ();
 sg13g2_decap_8 FILLER_63_355 ();
 sg13g2_decap_8 FILLER_63_362 ();
 sg13g2_decap_8 FILLER_63_369 ();
 sg13g2_fill_2 FILLER_63_407 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_decap_8 FILLER_64_112 ();
 sg13g2_decap_8 FILLER_64_119 ();
 sg13g2_decap_8 FILLER_64_126 ();
 sg13g2_decap_8 FILLER_64_133 ();
 sg13g2_decap_8 FILLER_64_140 ();
 sg13g2_decap_8 FILLER_64_147 ();
 sg13g2_fill_2 FILLER_64_154 ();
 sg13g2_fill_1 FILLER_64_156 ();
 sg13g2_fill_1 FILLER_64_207 ();
 sg13g2_decap_4 FILLER_64_211 ();
 sg13g2_fill_1 FILLER_64_215 ();
 sg13g2_fill_2 FILLER_64_220 ();
 sg13g2_fill_1 FILLER_64_222 ();
 sg13g2_decap_8 FILLER_64_239 ();
 sg13g2_decap_8 FILLER_64_246 ();
 sg13g2_decap_8 FILLER_64_253 ();
 sg13g2_fill_2 FILLER_64_260 ();
 sg13g2_fill_2 FILLER_64_278 ();
 sg13g2_decap_4 FILLER_64_349 ();
 sg13g2_fill_2 FILLER_64_358 ();
 sg13g2_fill_1 FILLER_64_360 ();
 sg13g2_decap_8 FILLER_64_374 ();
 sg13g2_decap_4 FILLER_64_381 ();
 sg13g2_decap_8 FILLER_64_393 ();
 sg13g2_decap_8 FILLER_64_400 ();
 sg13g2_fill_2 FILLER_64_407 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_decap_8 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_decap_8 FILLER_65_119 ();
 sg13g2_decap_8 FILLER_65_126 ();
 sg13g2_decap_8 FILLER_65_133 ();
 sg13g2_decap_8 FILLER_65_140 ();
 sg13g2_decap_8 FILLER_65_147 ();
 sg13g2_decap_8 FILLER_65_154 ();
 sg13g2_decap_8 FILLER_65_174 ();
 sg13g2_fill_2 FILLER_65_181 ();
 sg13g2_fill_1 FILLER_65_183 ();
 sg13g2_decap_4 FILLER_65_231 ();
 sg13g2_fill_1 FILLER_65_235 ();
 sg13g2_decap_8 FILLER_65_244 ();
 sg13g2_decap_8 FILLER_65_251 ();
 sg13g2_decap_8 FILLER_65_258 ();
 sg13g2_fill_1 FILLER_65_265 ();
 sg13g2_decap_8 FILLER_65_271 ();
 sg13g2_decap_4 FILLER_65_278 ();
 sg13g2_fill_2 FILLER_65_282 ();
 sg13g2_decap_8 FILLER_65_328 ();
 sg13g2_decap_8 FILLER_65_335 ();
 sg13g2_decap_8 FILLER_65_342 ();
 sg13g2_decap_4 FILLER_65_349 ();
 sg13g2_fill_1 FILLER_65_353 ();
 sg13g2_decap_8 FILLER_65_358 ();
 sg13g2_decap_8 FILLER_65_365 ();
 sg13g2_fill_2 FILLER_65_372 ();
 sg13g2_fill_1 FILLER_65_374 ();
 sg13g2_fill_2 FILLER_65_407 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_decap_8 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_decap_8 FILLER_66_112 ();
 sg13g2_decap_8 FILLER_66_119 ();
 sg13g2_decap_8 FILLER_66_126 ();
 sg13g2_decap_8 FILLER_66_133 ();
 sg13g2_decap_8 FILLER_66_140 ();
 sg13g2_decap_8 FILLER_66_147 ();
 sg13g2_decap_8 FILLER_66_154 ();
 sg13g2_fill_1 FILLER_66_161 ();
 sg13g2_fill_2 FILLER_66_190 ();
 sg13g2_fill_2 FILLER_66_214 ();
 sg13g2_decap_4 FILLER_66_220 ();
 sg13g2_fill_2 FILLER_66_224 ();
 sg13g2_fill_2 FILLER_66_234 ();
 sg13g2_decap_4 FILLER_66_252 ();
 sg13g2_fill_2 FILLER_66_264 ();
 sg13g2_fill_1 FILLER_66_274 ();
 sg13g2_fill_2 FILLER_66_285 ();
 sg13g2_fill_1 FILLER_66_287 ();
 sg13g2_fill_2 FILLER_66_296 ();
 sg13g2_fill_1 FILLER_66_298 ();
 sg13g2_fill_2 FILLER_66_304 ();
 sg13g2_fill_1 FILLER_66_306 ();
 sg13g2_fill_2 FILLER_66_347 ();
 sg13g2_fill_1 FILLER_66_381 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_decap_8 FILLER_67_112 ();
 sg13g2_decap_8 FILLER_67_119 ();
 sg13g2_decap_8 FILLER_67_126 ();
 sg13g2_decap_8 FILLER_67_133 ();
 sg13g2_decap_8 FILLER_67_140 ();
 sg13g2_decap_8 FILLER_67_147 ();
 sg13g2_decap_8 FILLER_67_154 ();
 sg13g2_decap_4 FILLER_67_161 ();
 sg13g2_fill_1 FILLER_67_165 ();
 sg13g2_fill_1 FILLER_67_193 ();
 sg13g2_fill_2 FILLER_67_203 ();
 sg13g2_fill_2 FILLER_67_231 ();
 sg13g2_decap_8 FILLER_67_294 ();
 sg13g2_fill_2 FILLER_67_301 ();
 sg13g2_fill_1 FILLER_67_327 ();
 sg13g2_fill_2 FILLER_67_342 ();
 sg13g2_decap_8 FILLER_67_371 ();
 sg13g2_decap_8 FILLER_67_395 ();
 sg13g2_decap_8 FILLER_67_402 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_decap_8 FILLER_68_119 ();
 sg13g2_decap_8 FILLER_68_126 ();
 sg13g2_decap_8 FILLER_68_133 ();
 sg13g2_decap_8 FILLER_68_140 ();
 sg13g2_decap_8 FILLER_68_147 ();
 sg13g2_decap_8 FILLER_68_154 ();
 sg13g2_decap_8 FILLER_68_161 ();
 sg13g2_fill_2 FILLER_68_168 ();
 sg13g2_fill_2 FILLER_68_230 ();
 sg13g2_fill_1 FILLER_68_267 ();
 sg13g2_fill_1 FILLER_68_277 ();
 sg13g2_fill_2 FILLER_68_286 ();
 sg13g2_fill_1 FILLER_68_301 ();
 sg13g2_fill_1 FILLER_68_305 ();
 sg13g2_fill_2 FILLER_68_346 ();
 sg13g2_decap_8 FILLER_68_357 ();
 sg13g2_fill_1 FILLER_68_364 ();
 sg13g2_decap_4 FILLER_68_370 ();
 sg13g2_fill_1 FILLER_68_374 ();
 sg13g2_fill_2 FILLER_68_379 ();
 sg13g2_fill_1 FILLER_68_381 ();
 sg13g2_fill_1 FILLER_68_387 ();
 sg13g2_decap_8 FILLER_68_393 ();
 sg13g2_decap_8 FILLER_68_400 ();
 sg13g2_fill_2 FILLER_68_407 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_decap_8 FILLER_69_119 ();
 sg13g2_decap_8 FILLER_69_126 ();
 sg13g2_decap_8 FILLER_69_133 ();
 sg13g2_decap_8 FILLER_69_140 ();
 sg13g2_decap_8 FILLER_69_147 ();
 sg13g2_decap_8 FILLER_69_154 ();
 sg13g2_decap_8 FILLER_69_161 ();
 sg13g2_fill_1 FILLER_69_168 ();
 sg13g2_fill_2 FILLER_69_197 ();
 sg13g2_fill_2 FILLER_69_222 ();
 sg13g2_decap_8 FILLER_69_253 ();
 sg13g2_decap_8 FILLER_69_260 ();
 sg13g2_fill_2 FILLER_69_267 ();
 sg13g2_decap_8 FILLER_69_273 ();
 sg13g2_fill_1 FILLER_69_280 ();
 sg13g2_decap_8 FILLER_69_315 ();
 sg13g2_decap_4 FILLER_69_322 ();
 sg13g2_fill_1 FILLER_69_326 ();
 sg13g2_decap_8 FILLER_69_354 ();
 sg13g2_decap_4 FILLER_69_361 ();
 sg13g2_fill_1 FILLER_69_365 ();
 sg13g2_decap_8 FILLER_69_397 ();
 sg13g2_decap_4 FILLER_69_404 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_decap_8 FILLER_70_133 ();
 sg13g2_decap_8 FILLER_70_140 ();
 sg13g2_decap_8 FILLER_70_147 ();
 sg13g2_decap_8 FILLER_70_154 ();
 sg13g2_decap_8 FILLER_70_161 ();
 sg13g2_decap_8 FILLER_70_168 ();
 sg13g2_fill_2 FILLER_70_175 ();
 sg13g2_fill_1 FILLER_70_177 ();
 sg13g2_decap_4 FILLER_70_193 ();
 sg13g2_fill_1 FILLER_70_197 ();
 sg13g2_fill_1 FILLER_70_210 ();
 sg13g2_fill_2 FILLER_70_221 ();
 sg13g2_decap_8 FILLER_70_228 ();
 sg13g2_decap_8 FILLER_70_235 ();
 sg13g2_decap_8 FILLER_70_242 ();
 sg13g2_decap_8 FILLER_70_249 ();
 sg13g2_decap_8 FILLER_70_256 ();
 sg13g2_decap_8 FILLER_70_263 ();
 sg13g2_decap_4 FILLER_70_270 ();
 sg13g2_decap_8 FILLER_70_279 ();
 sg13g2_fill_1 FILLER_70_286 ();
 sg13g2_fill_1 FILLER_70_312 ();
 sg13g2_fill_2 FILLER_70_326 ();
 sg13g2_fill_1 FILLER_70_328 ();
 sg13g2_decap_8 FILLER_70_356 ();
 sg13g2_decap_8 FILLER_70_363 ();
 sg13g2_fill_1 FILLER_70_370 ();
 sg13g2_fill_2 FILLER_70_380 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_133 ();
 sg13g2_decap_8 FILLER_71_140 ();
 sg13g2_decap_8 FILLER_71_147 ();
 sg13g2_decap_8 FILLER_71_154 ();
 sg13g2_decap_8 FILLER_71_161 ();
 sg13g2_decap_8 FILLER_71_168 ();
 sg13g2_decap_4 FILLER_71_175 ();
 sg13g2_decap_4 FILLER_71_185 ();
 sg13g2_fill_1 FILLER_71_189 ();
 sg13g2_fill_2 FILLER_71_194 ();
 sg13g2_fill_2 FILLER_71_201 ();
 sg13g2_fill_1 FILLER_71_203 ();
 sg13g2_decap_8 FILLER_71_209 ();
 sg13g2_decap_8 FILLER_71_216 ();
 sg13g2_decap_8 FILLER_71_223 ();
 sg13g2_decap_4 FILLER_71_230 ();
 sg13g2_fill_1 FILLER_71_234 ();
 sg13g2_fill_2 FILLER_71_250 ();
 sg13g2_fill_1 FILLER_71_266 ();
 sg13g2_decap_8 FILLER_71_285 ();
 sg13g2_decap_8 FILLER_71_292 ();
 sg13g2_decap_8 FILLER_71_299 ();
 sg13g2_fill_2 FILLER_71_306 ();
 sg13g2_fill_1 FILLER_71_308 ();
 sg13g2_decap_4 FILLER_71_313 ();
 sg13g2_fill_1 FILLER_71_317 ();
 sg13g2_fill_2 FILLER_71_333 ();
 sg13g2_fill_1 FILLER_71_335 ();
 sg13g2_fill_2 FILLER_71_363 ();
 sg13g2_decap_8 FILLER_71_370 ();
 sg13g2_fill_1 FILLER_71_377 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_decap_8 FILLER_72_140 ();
 sg13g2_decap_8 FILLER_72_147 ();
 sg13g2_decap_8 FILLER_72_154 ();
 sg13g2_decap_8 FILLER_72_161 ();
 sg13g2_decap_4 FILLER_72_205 ();
 sg13g2_decap_8 FILLER_72_221 ();
 sg13g2_fill_2 FILLER_72_228 ();
 sg13g2_decap_8 FILLER_72_285 ();
 sg13g2_fill_1 FILLER_72_292 ();
 sg13g2_fill_1 FILLER_72_298 ();
 sg13g2_decap_8 FILLER_72_307 ();
 sg13g2_decap_8 FILLER_72_314 ();
 sg13g2_fill_2 FILLER_72_330 ();
 sg13g2_decap_4 FILLER_72_403 ();
 sg13g2_fill_2 FILLER_72_407 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_8 FILLER_73_140 ();
 sg13g2_decap_8 FILLER_73_147 ();
 sg13g2_decap_8 FILLER_73_154 ();
 sg13g2_decap_8 FILLER_73_161 ();
 sg13g2_decap_8 FILLER_73_168 ();
 sg13g2_decap_4 FILLER_73_175 ();
 sg13g2_fill_1 FILLER_73_179 ();
 sg13g2_fill_2 FILLER_73_257 ();
 sg13g2_decap_4 FILLER_73_337 ();
 sg13g2_decap_8 FILLER_73_345 ();
 sg13g2_fill_2 FILLER_73_352 ();
 sg13g2_decap_8 FILLER_73_358 ();
 sg13g2_decap_8 FILLER_73_365 ();
 sg13g2_decap_8 FILLER_73_372 ();
 sg13g2_fill_1 FILLER_73_379 ();
 sg13g2_decap_8 FILLER_73_384 ();
 sg13g2_decap_8 FILLER_73_391 ();
 sg13g2_decap_8 FILLER_73_398 ();
 sg13g2_decap_4 FILLER_73_405 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_8 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_147 ();
 sg13g2_decap_8 FILLER_74_154 ();
 sg13g2_decap_8 FILLER_74_161 ();
 sg13g2_decap_4 FILLER_74_168 ();
 sg13g2_decap_4 FILLER_74_199 ();
 sg13g2_fill_2 FILLER_74_207 ();
 sg13g2_fill_1 FILLER_74_209 ();
 sg13g2_decap_8 FILLER_74_220 ();
 sg13g2_fill_1 FILLER_74_227 ();
 sg13g2_fill_2 FILLER_74_250 ();
 sg13g2_fill_1 FILLER_74_252 ();
 sg13g2_fill_1 FILLER_74_263 ();
 sg13g2_decap_4 FILLER_74_285 ();
 sg13g2_fill_2 FILLER_74_289 ();
 sg13g2_decap_8 FILLER_74_300 ();
 sg13g2_decap_8 FILLER_74_317 ();
 sg13g2_fill_2 FILLER_74_324 ();
 sg13g2_fill_1 FILLER_74_335 ();
 sg13g2_decap_8 FILLER_74_341 ();
 sg13g2_fill_2 FILLER_74_348 ();
 sg13g2_decap_8 FILLER_74_363 ();
 sg13g2_fill_2 FILLER_74_370 ();
 sg13g2_decap_4 FILLER_74_377 ();
 sg13g2_fill_2 FILLER_74_381 ();
 sg13g2_decap_8 FILLER_74_400 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_decap_8 FILLER_75_161 ();
 sg13g2_decap_4 FILLER_75_202 ();
 sg13g2_fill_1 FILLER_75_206 ();
 sg13g2_decap_8 FILLER_75_220 ();
 sg13g2_decap_8 FILLER_75_227 ();
 sg13g2_fill_1 FILLER_75_234 ();
 sg13g2_decap_8 FILLER_75_240 ();
 sg13g2_decap_8 FILLER_75_247 ();
 sg13g2_decap_8 FILLER_75_254 ();
 sg13g2_fill_2 FILLER_75_261 ();
 sg13g2_fill_2 FILLER_75_267 ();
 sg13g2_fill_1 FILLER_75_269 ();
 sg13g2_fill_2 FILLER_75_280 ();
 sg13g2_fill_1 FILLER_75_282 ();
 sg13g2_fill_2 FILLER_75_311 ();
 sg13g2_fill_1 FILLER_75_313 ();
 sg13g2_fill_2 FILLER_75_346 ();
 sg13g2_fill_2 FILLER_75_375 ();
 sg13g2_fill_1 FILLER_75_377 ();
 sg13g2_decap_4 FILLER_75_405 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_decap_8 FILLER_76_168 ();
 sg13g2_fill_1 FILLER_76_175 ();
 sg13g2_fill_1 FILLER_76_198 ();
 sg13g2_decap_8 FILLER_76_212 ();
 sg13g2_fill_1 FILLER_76_219 ();
 sg13g2_decap_4 FILLER_76_236 ();
 sg13g2_fill_2 FILLER_76_240 ();
 sg13g2_decap_8 FILLER_76_251 ();
 sg13g2_decap_8 FILLER_76_258 ();
 sg13g2_fill_2 FILLER_76_265 ();
 sg13g2_decap_8 FILLER_76_314 ();
 sg13g2_decap_8 FILLER_76_321 ();
 sg13g2_decap_4 FILLER_76_328 ();
 sg13g2_fill_2 FILLER_76_345 ();
 sg13g2_fill_2 FILLER_76_379 ();
 sg13g2_fill_1 FILLER_76_381 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_161 ();
 sg13g2_decap_8 FILLER_77_168 ();
 sg13g2_decap_4 FILLER_77_175 ();
 sg13g2_fill_2 FILLER_77_179 ();
 sg13g2_fill_2 FILLER_77_185 ();
 sg13g2_fill_1 FILLER_77_200 ();
 sg13g2_fill_2 FILLER_77_210 ();
 sg13g2_fill_2 FILLER_77_274 ();
 sg13g2_fill_2 FILLER_77_289 ();
 sg13g2_decap_4 FILLER_77_343 ();
 sg13g2_fill_2 FILLER_77_347 ();
 sg13g2_decap_8 FILLER_77_357 ();
 sg13g2_decap_4 FILLER_77_364 ();
 sg13g2_decap_4 FILLER_77_381 ();
 sg13g2_fill_2 FILLER_77_385 ();
 sg13g2_decap_8 FILLER_77_391 ();
 sg13g2_decap_8 FILLER_77_398 ();
 sg13g2_decap_4 FILLER_77_405 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_8 FILLER_78_154 ();
 sg13g2_decap_8 FILLER_78_161 ();
 sg13g2_decap_8 FILLER_78_168 ();
 sg13g2_fill_2 FILLER_78_175 ();
 sg13g2_fill_1 FILLER_78_177 ();
 sg13g2_decap_4 FILLER_78_206 ();
 sg13g2_fill_1 FILLER_78_210 ();
 sg13g2_fill_2 FILLER_78_239 ();
 sg13g2_fill_1 FILLER_78_247 ();
 sg13g2_fill_2 FILLER_78_273 ();
 sg13g2_fill_1 FILLER_78_275 ();
 sg13g2_fill_1 FILLER_78_294 ();
 sg13g2_fill_1 FILLER_78_342 ();
 sg13g2_fill_2 FILLER_78_370 ();
 sg13g2_fill_2 FILLER_78_377 ();
 sg13g2_fill_1 FILLER_78_379 ();
 sg13g2_fill_2 FILLER_78_407 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_168 ();
 sg13g2_decap_8 FILLER_79_175 ();
 sg13g2_decap_8 FILLER_79_182 ();
 sg13g2_decap_8 FILLER_79_189 ();
 sg13g2_fill_1 FILLER_79_239 ();
 sg13g2_fill_2 FILLER_79_268 ();
 sg13g2_fill_1 FILLER_79_270 ();
 sg13g2_fill_1 FILLER_79_276 ();
 sg13g2_decap_8 FILLER_79_280 ();
 sg13g2_fill_2 FILLER_79_287 ();
 sg13g2_fill_1 FILLER_79_292 ();
 sg13g2_decap_4 FILLER_79_298 ();
 sg13g2_fill_1 FILLER_79_302 ();
 sg13g2_fill_2 FILLER_79_309 ();
 sg13g2_fill_1 FILLER_79_311 ();
 sg13g2_fill_2 FILLER_79_340 ();
 sg13g2_fill_2 FILLER_79_378 ();
 sg13g2_fill_2 FILLER_79_407 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_8 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_139 ();
 sg13g2_fill_1 FILLER_80_143 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_201 ();
 sg13g2_decap_8 FILLER_80_208 ();
 sg13g2_decap_8 FILLER_80_215 ();
 sg13g2_fill_2 FILLER_80_222 ();
 sg13g2_fill_1 FILLER_80_224 ();
 sg13g2_decap_8 FILLER_80_234 ();
 sg13g2_fill_2 FILLER_80_241 ();
 sg13g2_decap_4 FILLER_80_255 ();
 sg13g2_decap_4 FILLER_80_268 ();
 sg13g2_decap_8 FILLER_80_277 ();
 sg13g2_decap_4 FILLER_80_284 ();
 sg13g2_fill_2 FILLER_80_293 ();
 sg13g2_fill_1 FILLER_80_295 ();
 sg13g2_fill_2 FILLER_80_300 ();
 sg13g2_fill_1 FILLER_80_302 ();
 sg13g2_fill_2 FILLER_80_349 ();
 sg13g2_fill_1 FILLER_80_351 ();
 sg13g2_fill_2 FILLER_80_365 ();
 sg13g2_fill_1 FILLER_80_367 ();
 sg13g2_decap_8 FILLER_80_372 ();
 sg13g2_decap_4 FILLER_80_379 ();
 sg13g2_fill_2 FILLER_80_383 ();
 sg13g2_decap_8 FILLER_80_397 ();
 sg13g2_decap_4 FILLER_80_404 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net14;
 assign uio_oe[1] = net15;
 assign uio_oe[2] = net16;
 assign uio_oe[3] = net17;
 assign uio_oe[4] = net18;
 assign uio_oe[5] = net138;
 assign uio_oe[6] = net19;
 assign uio_oe[7] = net20;
 assign uio_out[0] = net21;
 assign uio_out[1] = net22;
 assign uio_out[2] = net23;
 assign uio_out[3] = net24;
 assign uio_out[4] = net25;
 assign uio_out[6] = net26;
 assign uio_out[7] = net27;
endmodule
