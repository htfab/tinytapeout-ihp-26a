module tt_um_matth_fischer_vgaTT (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire clknet_0_clk;
 wire \abs_x[0] ;
 wire \abs_y[0] ;
 wire \anim_offset[1] ;
 wire \anim_offset[2] ;
 wire \anim_offset[3] ;
 wire \anim_offset[4] ;
 wire \anim_offset[5] ;
 wire \anim_offset[6] ;
 wire \anim_offset[7] ;
 wire \cx[1] ;
 wire \cx[2] ;
 wire \cx[3] ;
 wire \cx[4] ;
 wire \cx[5] ;
 wire \cy[1] ;
 wire \cy[2] ;
 wire \cy[3] ;
 wire \hpos[6] ;
 wire \hpos[7] ;
 wire \hpos[8] ;
 wire \hpos[9] ;
 wire hsync;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net1;
 wire net2;
 wire net3;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;

 sg13g2_inv_1 _296_ (.Y(_240_),
    .A(\cx[4] ));
 sg13g2_inv_2 _297_ (.Y(_241_),
    .A(net42));
 sg13g2_inv_2 _298_ (.Y(_242_),
    .A(net39));
 sg13g2_inv_1 _299_ (.Y(_243_),
    .A(net88));
 sg13g2_inv_1 _300_ (.Y(_244_),
    .A(net82));
 sg13g2_inv_1 _301_ (.Y(_245_),
    .A(\anim_offset[1] ));
 sg13g2_inv_1 _302_ (.Y(_246_),
    .A(net2));
 sg13g2_and2_1 _303_ (.A(net84),
    .B(net37),
    .X(_247_));
 sg13g2_nand3_1 _304_ (.B(net71),
    .C(_247_),
    .A(net38),
    .Y(_248_));
 sg13g2_nand2_1 _305_ (.Y(_249_),
    .A(net80),
    .B(net76));
 sg13g2_nor2_1 _306_ (.A(net39),
    .B(net68),
    .Y(_250_));
 sg13g2_nand4_1 _307_ (.B(net80),
    .C(_249_),
    .A(net40),
    .Y(_251_),
    .D(_250_));
 sg13g2_nor2_1 _308_ (.A(_248_),
    .B(net90),
    .Y(_001_));
 sg13g2_nor2_1 _309_ (.A(\cx[4] ),
    .B(\cx[5] ),
    .Y(_252_));
 sg13g2_nor3_1 _310_ (.A(\cx[4] ),
    .B(\cx[5] ),
    .C(net44),
    .Y(_253_));
 sg13g2_nand2_1 _311_ (.Y(_254_),
    .A(net73),
    .B(net42));
 sg13g2_and4_1 _312_ (.A(net92),
    .B(net86),
    .C(net73),
    .D(net44),
    .X(_255_));
 sg13g2_nor4_1 _313_ (.A(net43),
    .B(_253_),
    .C(net74),
    .D(_255_),
    .Y(_000_));
 sg13g2_and2_1 _314_ (.A(net39),
    .B(net38),
    .X(_256_));
 sg13g2_and4_1 _315_ (.A(net39),
    .B(net38),
    .C(\hvsync_gen.vpos[7] ),
    .D(net37),
    .X(_257_));
 sg13g2_nand4_1 _316_ (.B(net38),
    .C(\hvsync_gen.vpos[7] ),
    .A(net39),
    .Y(_258_),
    .D(net37));
 sg13g2_nor2_1 _317_ (.A(\hvsync_gen.vpos[8] ),
    .B(\hvsync_gen.vpos[9] ),
    .Y(_259_));
 sg13g2_or2_1 _318_ (.X(_260_),
    .B(\hvsync_gen.vpos[9] ),
    .A(\hvsync_gen.vpos[8] ));
 sg13g2_nor2_1 _319_ (.A(_257_),
    .B(net36),
    .Y(_261_));
 sg13g2_or2_1 _320_ (.X(_262_),
    .B(net40),
    .A(net41));
 sg13g2_nor3_1 _321_ (.A(net41),
    .B(net40),
    .C(\cy[2] ),
    .Y(_263_));
 sg13g2_nor4_2 _322_ (.A(net41),
    .B(net40),
    .C(\cy[3] ),
    .Y(_264_),
    .D(\cy[2] ));
 sg13g2_nor3_1 _323_ (.A(_257_),
    .B(net36),
    .C(_264_),
    .Y(_265_));
 sg13g2_nand2_1 _324_ (.Y(_266_),
    .A(_256_),
    .B(_264_));
 sg13g2_xor2_1 _325_ (.B(net38),
    .A(net39),
    .X(_267_));
 sg13g2_a221oi_1 _326_ (.B2(net39),
    .C1(net36),
    .B1(_264_),
    .A1(_247_),
    .Y(_268_),
    .A2(_256_));
 sg13g2_xnor2_1 _327_ (.Y(_269_),
    .A(_267_),
    .B(_268_));
 sg13g2_or2_1 _328_ (.X(_270_),
    .B(net44),
    .A(\hpos[7] ));
 sg13g2_o21ai_1 _329_ (.B1(net43),
    .Y(_271_),
    .A1(\hpos[7] ),
    .A2(net44));
 sg13g2_and2_1 _330_ (.A(_241_),
    .B(_271_),
    .X(_272_));
 sg13g2_or2_1 _331_ (.X(_273_),
    .B(\cx[1] ),
    .A(net45));
 sg13g2_or3_1 _332_ (.A(net45),
    .B(\cx[1] ),
    .C(\cx[2] ),
    .X(_029_));
 sg13g2_nor4_2 _333_ (.A(net45),
    .B(\cx[1] ),
    .C(\cx[3] ),
    .Y(_030_),
    .D(\cx[2] ));
 sg13g2_or4_1 _334_ (.A(net45),
    .B(\cx[1] ),
    .C(\cx[3] ),
    .D(\cx[2] ),
    .X(_031_));
 sg13g2_nand3_1 _335_ (.B(_271_),
    .C(_031_),
    .A(_241_),
    .Y(_032_));
 sg13g2_a221oi_1 _336_ (.B2(_240_),
    .C1(net42),
    .B1(_030_),
    .A1(net43),
    .Y(_033_),
    .A2(_270_));
 sg13g2_xor2_1 _337_ (.B(_033_),
    .A(\cx[5] ),
    .X(_034_));
 sg13g2_nor2_1 _338_ (.A(_269_),
    .B(_034_),
    .Y(_035_));
 sg13g2_nand3_1 _339_ (.B(_271_),
    .C(_273_),
    .A(_241_),
    .Y(_036_));
 sg13g2_xor2_1 _340_ (.B(_036_),
    .A(\cx[2] ),
    .X(_037_));
 sg13g2_nand3_1 _341_ (.B(_259_),
    .C(_262_),
    .A(_258_),
    .Y(_038_));
 sg13g2_xnor2_1 _342_ (.Y(_039_),
    .A(\cy[2] ),
    .B(_038_));
 sg13g2_nor2_1 _343_ (.A(_037_),
    .B(_039_),
    .Y(_040_));
 sg13g2_nand3_1 _344_ (.B(_271_),
    .C(_029_),
    .A(_241_),
    .Y(_041_));
 sg13g2_xor2_1 _345_ (.B(_041_),
    .A(\cx[3] ),
    .X(_042_));
 sg13g2_xnor2_1 _346_ (.Y(_043_),
    .A(\cx[3] ),
    .B(_041_));
 sg13g2_nor3_1 _347_ (.A(_257_),
    .B(net36),
    .C(_263_),
    .Y(_044_));
 sg13g2_xor2_1 _348_ (.B(_044_),
    .A(\cy[3] ),
    .X(_045_));
 sg13g2_xnor2_1 _349_ (.Y(_046_),
    .A(\cy[3] ),
    .B(_044_));
 sg13g2_or4_1 _350_ (.A(_037_),
    .B(_039_),
    .C(_043_),
    .D(_046_),
    .X(_047_));
 sg13g2_xnor2_1 _351_ (.Y(_048_),
    .A(\cx[4] ),
    .B(_032_));
 sg13g2_xnor2_1 _352_ (.Y(_049_),
    .A(_242_),
    .B(_265_));
 sg13g2_nor2_1 _353_ (.A(_048_),
    .B(_049_),
    .Y(_050_));
 sg13g2_nand3_1 _354_ (.B(net38),
    .C(net37),
    .A(\hvsync_gen.vpos[4] ),
    .Y(_051_));
 sg13g2_and2_1 _355_ (.A(net36),
    .B(_051_),
    .X(_052_));
 sg13g2_nor4_1 _356_ (.A(_257_),
    .B(_260_),
    .C(_264_),
    .D(_051_),
    .Y(_053_));
 sg13g2_o21ai_1 _357_ (.B1(\hvsync_gen.vpos[7] ),
    .Y(_054_),
    .A1(_052_),
    .A2(_053_));
 sg13g2_or3_1 _358_ (.A(\hvsync_gen.vpos[7] ),
    .B(_052_),
    .C(_053_),
    .X(_055_));
 sg13g2_xnor2_1 _359_ (.Y(_056_),
    .A(\hpos[7] ),
    .B(net44));
 sg13g2_nand3_1 _360_ (.B(_252_),
    .C(_030_),
    .A(net44),
    .Y(_057_));
 sg13g2_nand3_1 _361_ (.B(_056_),
    .C(_057_),
    .A(_272_),
    .Y(_058_));
 sg13g2_a21o_2 _362_ (.A2(_057_),
    .A1(_272_),
    .B1(_056_),
    .X(_059_));
 sg13g2_and2_1 _363_ (.A(_058_),
    .B(_059_),
    .X(_060_));
 sg13g2_a22oi_1 _364_ (.Y(_061_),
    .B1(_058_),
    .B2(_059_),
    .A2(_055_),
    .A1(_054_));
 sg13g2_a22oi_1 _365_ (.Y(_062_),
    .B1(_048_),
    .B2(_049_),
    .A2(_034_),
    .A1(_269_));
 sg13g2_nand2_1 _366_ (.Y(_063_),
    .A(net41),
    .B(\cy[1] ));
 sg13g2_xor2_1 _367_ (.B(net40),
    .A(net41),
    .X(_064_));
 sg13g2_nor3_1 _368_ (.A(_257_),
    .B(net36),
    .C(_064_),
    .Y(_065_));
 sg13g2_a21oi_1 _369_ (.A1(_258_),
    .A2(_259_),
    .Y(_066_),
    .B1(net40));
 sg13g2_xnor2_1 _370_ (.Y(_067_),
    .A(net45),
    .B(net103));
 sg13g2_nand3_1 _371_ (.B(_271_),
    .C(_067_),
    .A(_241_),
    .Y(_068_));
 sg13g2_o21ai_1 _372_ (.B1(_068_),
    .Y(_069_),
    .A1(\cx[1] ),
    .A2(_272_));
 sg13g2_nand2b_1 _373_ (.Y(_070_),
    .B(\abs_y[0] ),
    .A_N(\abs_x[0] ));
 sg13g2_a22oi_1 _374_ (.Y(_071_),
    .B1(_042_),
    .B2(_045_),
    .A2(_039_),
    .A1(_037_));
 sg13g2_nor3_1 _375_ (.A(_065_),
    .B(_066_),
    .C(_070_),
    .Y(_072_));
 sg13g2_o21ai_1 _376_ (.B1(_070_),
    .Y(_073_),
    .A1(_065_),
    .A2(_066_));
 sg13g2_o21ai_1 _377_ (.B1(_073_),
    .Y(_074_),
    .A1(_069_),
    .A2(_072_));
 sg13g2_a221oi_1 _378_ (.B2(_074_),
    .C1(_040_),
    .B1(_071_),
    .A1(_043_),
    .Y(_075_),
    .A2(_046_));
 sg13g2_and4_1 _379_ (.A(_054_),
    .B(_055_),
    .C(_058_),
    .D(_059_),
    .X(_076_));
 sg13g2_nand4_1 _380_ (.B(_055_),
    .C(_058_),
    .A(_054_),
    .Y(_077_),
    .D(_059_));
 sg13g2_a221oi_1 _381_ (.B2(_252_),
    .C1(net42),
    .B1(_030_),
    .A1(net43),
    .Y(_078_),
    .A2(_270_));
 sg13g2_xnor2_1 _382_ (.Y(_079_),
    .A(\hpos[6] ),
    .B(_078_));
 sg13g2_xnor2_1 _383_ (.Y(_080_),
    .A(net37),
    .B(_256_));
 sg13g2_nand3_1 _384_ (.B(_266_),
    .C(_080_),
    .A(_261_),
    .Y(_081_));
 sg13g2_a21o_2 _385_ (.A2(_266_),
    .A1(_261_),
    .B1(_080_),
    .X(_082_));
 sg13g2_nand2_1 _386_ (.Y(_083_),
    .A(_081_),
    .B(_082_));
 sg13g2_and3_1 _387_ (.X(_084_),
    .A(_079_),
    .B(_081_),
    .C(_082_));
 sg13g2_nand3_1 _388_ (.B(_081_),
    .C(_082_),
    .A(_079_),
    .Y(_085_));
 sg13g2_a21oi_1 _389_ (.A1(_081_),
    .A2(_082_),
    .Y(_086_),
    .B1(_079_));
 sg13g2_nor4_1 _390_ (.A(_061_),
    .B(_076_),
    .C(_084_),
    .D(_086_),
    .Y(_087_));
 sg13g2_or4_1 _391_ (.A(_061_),
    .B(_076_),
    .C(_084_),
    .D(_086_),
    .X(_088_));
 sg13g2_nand3b_1 _392_ (.B(_047_),
    .C(_062_),
    .Y(_089_),
    .A_N(_035_));
 sg13g2_or4_1 _393_ (.A(_050_),
    .B(_075_),
    .C(_088_),
    .D(_089_),
    .X(_090_));
 sg13g2_nor2_1 _394_ (.A(_035_),
    .B(_062_),
    .Y(_091_));
 sg13g2_a21oi_1 _395_ (.A1(_077_),
    .A2(_085_),
    .Y(_092_),
    .B1(_061_));
 sg13g2_a21oi_1 _396_ (.A1(_087_),
    .A2(_091_),
    .Y(_093_),
    .B1(_092_));
 sg13g2_nand2_1 _397_ (.Y(_094_),
    .A(net43),
    .B(\hpos[9] ));
 sg13g2_nor2_1 _398_ (.A(_241_),
    .B(_271_),
    .Y(_095_));
 sg13g2_or2_1 _399_ (.X(_096_),
    .B(_271_),
    .A(_241_));
 sg13g2_o21ai_1 _400_ (.B1(\hvsync_gen.vpos[9] ),
    .Y(_097_),
    .A1(\hvsync_gen.vpos[8] ),
    .A2(_257_));
 sg13g2_nor2_1 _401_ (.A(_095_),
    .B(_097_),
    .Y(_098_));
 sg13g2_inv_1 _402_ (.Y(_099_),
    .A(_098_));
 sg13g2_nor2_1 _403_ (.A(net43),
    .B(_270_),
    .Y(_100_));
 sg13g2_nor2_1 _404_ (.A(net42),
    .B(_100_),
    .Y(_101_));
 sg13g2_o21ai_1 _405_ (.B1(_101_),
    .Y(_102_),
    .A1(\hpos[7] ),
    .A2(_057_));
 sg13g2_nand2_1 _406_ (.Y(_103_),
    .A(\hpos[9] ),
    .B(_100_));
 sg13g2_and3_1 _407_ (.X(_104_),
    .A(_271_),
    .B(_102_),
    .C(_103_));
 sg13g2_xnor2_1 _408_ (.Y(_105_),
    .A(\hvsync_gen.vpos[8] ),
    .B(_257_));
 sg13g2_nand2_1 _409_ (.Y(_106_),
    .A(net36),
    .B(_105_));
 sg13g2_o21ai_1 _410_ (.B1(_099_),
    .Y(_107_),
    .A1(_104_),
    .A2(_106_));
 sg13g2_a21oi_2 _411_ (.B1(_107_),
    .Y(_108_),
    .A2(_093_),
    .A1(_090_));
 sg13g2_a21o_1 _412_ (.A2(_093_),
    .A1(_090_),
    .B1(_107_),
    .X(_109_));
 sg13g2_nand2_1 _413_ (.Y(_110_),
    .A(_095_),
    .B(_097_));
 sg13g2_nand2_1 _414_ (.Y(_111_),
    .A(_104_),
    .B(_106_));
 sg13g2_a21o_1 _415_ (.A2(_111_),
    .A1(_110_),
    .B1(_098_),
    .X(_112_));
 sg13g2_a21oi_2 _416_ (.B1(_098_),
    .Y(_113_),
    .A2(_111_),
    .A1(_110_));
 sg13g2_nor2_1 _417_ (.A(_108_),
    .B(_113_),
    .Y(_114_));
 sg13g2_a21oi_1 _418_ (.A1(_109_),
    .A2(_112_),
    .Y(_115_),
    .B1(\abs_x[0] ));
 sg13g2_nor3_1 _419_ (.A(\abs_y[0] ),
    .B(_108_),
    .C(_113_),
    .Y(_116_));
 sg13g2_nor4_2 _420_ (.A(_096_),
    .B(_097_),
    .C(_115_),
    .Y(_117_),
    .D(_116_));
 sg13g2_or4_1 _421_ (.A(_065_),
    .B(_066_),
    .C(_108_),
    .D(_113_),
    .X(_118_));
 sg13g2_o21ai_1 _422_ (.B1(_118_),
    .Y(_119_),
    .A1(_069_),
    .A2(net33));
 sg13g2_nand2_1 _423_ (.Y(_120_),
    .A(_117_),
    .B(_119_));
 sg13g2_nor3_1 _424_ (.A(_039_),
    .B(_108_),
    .C(_113_),
    .Y(_121_));
 sg13g2_o21ai_1 _425_ (.B1(_037_),
    .Y(_122_),
    .A1(_108_),
    .A2(_113_));
 sg13g2_nor2b_2 _426_ (.A(_121_),
    .B_N(_122_),
    .Y(_123_));
 sg13g2_nand3_1 _427_ (.B(_119_),
    .C(_123_),
    .A(_117_),
    .Y(_124_));
 sg13g2_mux2_1 _428_ (.A0(_043_),
    .A1(_045_),
    .S(net33),
    .X(_125_));
 sg13g2_nand4_1 _429_ (.B(_119_),
    .C(_123_),
    .A(_117_),
    .Y(_126_),
    .D(_125_));
 sg13g2_nand2_1 _430_ (.Y(_127_),
    .A(_049_),
    .B(net33));
 sg13g2_o21ai_1 _431_ (.B1(_127_),
    .Y(_128_),
    .A1(_048_),
    .A2(net33));
 sg13g2_nor2_1 _432_ (.A(_126_),
    .B(_128_),
    .Y(_129_));
 sg13g2_xor2_1 _433_ (.B(_128_),
    .A(_126_),
    .X(_130_));
 sg13g2_nor2_1 _434_ (.A(\anim_offset[2] ),
    .B(\anim_offset[1] ),
    .Y(_131_));
 sg13g2_nor2_1 _435_ (.A(_245_),
    .B(net2),
    .Y(_132_));
 sg13g2_nor2_1 _436_ (.A(net2),
    .B(_131_),
    .Y(_133_));
 sg13g2_a21oi_1 _437_ (.A1(_244_),
    .A2(_131_),
    .Y(_134_),
    .B1(net2));
 sg13g2_xnor2_1 _438_ (.Y(_135_),
    .A(\anim_offset[4] ),
    .B(_134_));
 sg13g2_nand2_1 _439_ (.Y(_136_),
    .A(_130_),
    .B(_135_));
 sg13g2_xor2_1 _440_ (.B(_135_),
    .A(_130_),
    .X(_137_));
 sg13g2_xor2_1 _441_ (.B(_125_),
    .A(_124_),
    .X(_138_));
 sg13g2_xnor2_1 _442_ (.Y(_139_),
    .A(\anim_offset[3] ),
    .B(_133_));
 sg13g2_inv_1 _443_ (.Y(_140_),
    .A(_139_));
 sg13g2_xnor2_1 _444_ (.Y(_141_),
    .A(\anim_offset[2] ),
    .B(_132_));
 sg13g2_xor2_1 _445_ (.B(_123_),
    .A(_120_),
    .X(_142_));
 sg13g2_xor2_1 _446_ (.B(_119_),
    .A(_117_),
    .X(_143_));
 sg13g2_nor2_1 _447_ (.A(_138_),
    .B(_140_),
    .Y(_144_));
 sg13g2_o21ai_1 _448_ (.B1(_141_),
    .Y(_145_),
    .A1(_245_),
    .A2(_143_));
 sg13g2_nor3_1 _449_ (.A(_245_),
    .B(_141_),
    .C(_143_),
    .Y(_146_));
 sg13g2_a221oi_1 _450_ (.B2(_145_),
    .C1(_146_),
    .B1(_142_),
    .A1(_138_),
    .Y(_147_),
    .A2(_140_));
 sg13g2_o21ai_1 _451_ (.B1(_137_),
    .Y(_148_),
    .A1(_144_),
    .A2(_147_));
 sg13g2_nor3_1 _452_ (.A(_137_),
    .B(_144_),
    .C(_147_),
    .Y(_149_));
 sg13g2_o21ai_1 _453_ (.B1(\hpos[9] ),
    .Y(_150_),
    .A1(\hpos[7] ),
    .A2(\hpos[8] ));
 sg13g2_nand3b_1 _454_ (.B(_248_),
    .C(_150_),
    .Y(_151_),
    .A_N(\hvsync_gen.vpos[9] ));
 sg13g2_nor2_1 _455_ (.A(_149_),
    .B(_151_),
    .Y(_152_));
 sg13g2_and2_1 _456_ (.A(_148_),
    .B(_152_),
    .X(uo_out[4]));
 sg13g2_nand2_1 _457_ (.Y(_153_),
    .A(_269_),
    .B(net33));
 sg13g2_o21ai_1 _458_ (.B1(_153_),
    .Y(_154_),
    .A1(_034_),
    .A2(net33));
 sg13g2_nor3_1 _459_ (.A(_126_),
    .B(_128_),
    .C(_154_),
    .Y(_155_));
 sg13g2_xnor2_1 _460_ (.Y(_156_),
    .A(_129_),
    .B(_154_));
 sg13g2_nor3_1 _461_ (.A(\anim_offset[4] ),
    .B(\anim_offset[3] ),
    .C(_133_),
    .Y(_157_));
 sg13g2_nor2_1 _462_ (.A(net2),
    .B(_157_),
    .Y(_158_));
 sg13g2_xnor2_1 _463_ (.Y(_159_),
    .A(\anim_offset[5] ),
    .B(_158_));
 sg13g2_and2_1 _464_ (.A(_156_),
    .B(_159_),
    .X(_160_));
 sg13g2_xnor2_1 _465_ (.Y(_161_),
    .A(_156_),
    .B(_159_));
 sg13g2_and3_1 _466_ (.X(_162_),
    .A(_136_),
    .B(_148_),
    .C(_161_));
 sg13g2_a21oi_1 _467_ (.A1(_136_),
    .A2(_148_),
    .Y(_163_),
    .B1(_161_));
 sg13g2_nor3_2 _468_ (.A(_151_),
    .B(_162_),
    .C(_163_),
    .Y(uo_out[5]));
 sg13g2_mux2_1 _469_ (.A0(_079_),
    .A1(_083_),
    .S(net33),
    .X(_164_));
 sg13g2_nand2_1 _470_ (.Y(_165_),
    .A(_155_),
    .B(_164_));
 sg13g2_xor2_1 _471_ (.B(_164_),
    .A(_155_),
    .X(_166_));
 sg13g2_a21oi_1 _472_ (.A1(_243_),
    .A2(_157_),
    .Y(_167_),
    .B1(net2));
 sg13g2_xor2_1 _473_ (.B(_167_),
    .A(\anim_offset[6] ),
    .X(_168_));
 sg13g2_nand2b_1 _474_ (.Y(_169_),
    .B(_166_),
    .A_N(_168_));
 sg13g2_xnor2_1 _475_ (.Y(_170_),
    .A(_166_),
    .B(_168_));
 sg13g2_nor3_1 _476_ (.A(_160_),
    .B(_163_),
    .C(_170_),
    .Y(_171_));
 sg13g2_o21ai_1 _477_ (.B1(_170_),
    .Y(_172_),
    .A1(_160_),
    .A2(_163_));
 sg13g2_nand2b_1 _478_ (.Y(_173_),
    .B(_172_),
    .A_N(_171_));
 sg13g2_nor2_2 _479_ (.A(_151_),
    .B(_173_),
    .Y(uo_out[6]));
 sg13g2_o21ai_1 _480_ (.B1(_246_),
    .Y(_174_),
    .A1(\anim_offset[6] ),
    .A2(_167_));
 sg13g2_xnor2_1 _481_ (.Y(_175_),
    .A(\anim_offset[7] ),
    .B(_174_));
 sg13g2_nand3_1 _482_ (.B(_055_),
    .C(net33),
    .A(_054_),
    .Y(_176_));
 sg13g2_o21ai_1 _483_ (.B1(_176_),
    .Y(_177_),
    .A1(_060_),
    .A2(_114_));
 sg13g2_xnor2_1 _484_ (.Y(_178_),
    .A(_175_),
    .B(_177_));
 sg13g2_xnor2_1 _485_ (.Y(_179_),
    .A(_165_),
    .B(_178_));
 sg13g2_and3_1 _486_ (.X(_180_),
    .A(_169_),
    .B(_172_),
    .C(_179_));
 sg13g2_a21oi_1 _487_ (.A1(_169_),
    .A2(_172_),
    .Y(_181_),
    .B1(_179_));
 sg13g2_nor3_1 _488_ (.A(_151_),
    .B(_180_),
    .C(_181_),
    .Y(uo_out[2]));
 sg13g2_and3_1 _489_ (.X(_182_),
    .A(net45),
    .B(\cx[1] ),
    .C(net65));
 sg13g2_and2_1 _490_ (.A(net95),
    .B(_182_),
    .X(_183_));
 sg13g2_and2_1 _491_ (.A(net92),
    .B(_183_),
    .X(_184_));
 sg13g2_nor3_1 _492_ (.A(\cx[5] ),
    .B(_270_),
    .C(_094_),
    .Y(_185_));
 sg13g2_and2_1 _493_ (.A(_184_),
    .B(_185_),
    .X(_186_));
 sg13g2_nor2b_2 _494_ (.A(_186_),
    .B_N(net46),
    .Y(_187_));
 sg13g2_nand2b_2 _495_ (.Y(_188_),
    .B(net46),
    .A_N(_186_));
 sg13g2_nor2_1 _496_ (.A(net45),
    .B(_188_),
    .Y(_002_));
 sg13g2_nor2_1 _497_ (.A(_067_),
    .B(_188_),
    .Y(_003_));
 sg13g2_a21oi_1 _498_ (.A1(net45),
    .A2(\cx[1] ),
    .Y(_189_),
    .B1(net65));
 sg13g2_nor3_1 _499_ (.A(_182_),
    .B(_188_),
    .C(net66),
    .Y(_004_));
 sg13g2_o21ai_1 _500_ (.B1(net46),
    .Y(_190_),
    .A1(net95),
    .A2(_182_));
 sg13g2_nor2_1 _501_ (.A(_183_),
    .B(net96),
    .Y(_005_));
 sg13g2_o21ai_1 _502_ (.B1(net46),
    .Y(_191_),
    .A1(net92),
    .A2(_183_));
 sg13g2_nor2_1 _503_ (.A(_184_),
    .B(net93),
    .Y(_006_));
 sg13g2_and2_1 _504_ (.A(net86),
    .B(_184_),
    .X(_192_));
 sg13g2_nor2_1 _505_ (.A(net86),
    .B(_184_),
    .Y(_193_));
 sg13g2_nor3_1 _506_ (.A(_188_),
    .B(_192_),
    .C(net87),
    .Y(_007_));
 sg13g2_xnor2_1 _507_ (.Y(_194_),
    .A(net44),
    .B(_192_));
 sg13g2_nor2_1 _508_ (.A(_188_),
    .B(_194_),
    .Y(_008_));
 sg13g2_a21oi_1 _509_ (.A1(net44),
    .A2(_192_),
    .Y(_195_),
    .B1(net73));
 sg13g2_and2_1 _510_ (.A(_255_),
    .B(_183_),
    .X(_196_));
 sg13g2_nor3_1 _511_ (.A(_188_),
    .B(net79),
    .C(_196_),
    .Y(_009_));
 sg13g2_nor2_1 _512_ (.A(net43),
    .B(_196_),
    .Y(_197_));
 sg13g2_and2_1 _513_ (.A(net43),
    .B(_196_),
    .X(_198_));
 sg13g2_nor3_1 _514_ (.A(_188_),
    .B(_197_),
    .C(_198_),
    .Y(_010_));
 sg13g2_o21ai_1 _515_ (.B1(net35),
    .Y(_199_),
    .A1(net42),
    .A2(_198_));
 sg13g2_a21oi_1 _516_ (.A1(net42),
    .A2(_198_),
    .Y(_011_),
    .B1(_199_));
 sg13g2_or4_1 _517_ (.A(\hvsync_gen.vpos[4] ),
    .B(\hvsync_gen.vpos[5] ),
    .C(\hvsync_gen.vpos[7] ),
    .D(net37),
    .X(_200_));
 sg13g2_nor4_1 _518_ (.A(\hpos[8] ),
    .B(net42),
    .C(net36),
    .D(_270_),
    .Y(_201_));
 sg13g2_nand4_1 _519_ (.B(_264_),
    .C(_030_),
    .A(_252_),
    .Y(_202_),
    .D(_201_));
 sg13g2_or3_1 _520_ (.A(net1),
    .B(_200_),
    .C(_202_),
    .X(_203_));
 sg13g2_xnor2_1 _521_ (.Y(_012_),
    .A(net56),
    .B(_203_));
 sg13g2_nor2_1 _522_ (.A(net1),
    .B(net56),
    .Y(_204_));
 sg13g2_nor3_1 _523_ (.A(_200_),
    .B(_202_),
    .C(_204_),
    .Y(_205_));
 sg13g2_and2_1 _524_ (.A(net58),
    .B(_205_),
    .X(_206_));
 sg13g2_xor2_1 _525_ (.B(_205_),
    .A(net58),
    .X(_013_));
 sg13g2_and2_1 _526_ (.A(net82),
    .B(_206_),
    .X(_207_));
 sg13g2_xnor2_1 _527_ (.Y(_014_),
    .A(_244_),
    .B(_206_));
 sg13g2_and2_1 _528_ (.A(net60),
    .B(_207_),
    .X(_208_));
 sg13g2_xor2_1 _529_ (.B(_207_),
    .A(net60),
    .X(_015_));
 sg13g2_xnor2_1 _530_ (.Y(_016_),
    .A(_243_),
    .B(_208_));
 sg13g2_nand3_1 _531_ (.B(net97),
    .C(_208_),
    .A(net88),
    .Y(_209_));
 sg13g2_a21o_1 _532_ (.A2(_208_),
    .A1(net88),
    .B1(net97),
    .X(_210_));
 sg13g2_and2_1 _533_ (.A(_209_),
    .B(_210_),
    .X(_017_));
 sg13g2_xnor2_1 _534_ (.Y(_018_),
    .A(net62),
    .B(_209_));
 sg13g2_nand2_1 _535_ (.Y(_211_),
    .A(net46),
    .B(_186_));
 sg13g2_inv_1 _536_ (.Y(_212_),
    .A(_211_));
 sg13g2_nor4_1 _537_ (.A(_249_),
    .B(_262_),
    .C(_106_),
    .D(_200_),
    .Y(_213_));
 sg13g2_or2_1 _538_ (.X(_214_),
    .B(_213_),
    .A(_211_));
 sg13g2_inv_1 _539_ (.Y(_215_),
    .A(net34));
 sg13g2_nand2_1 _540_ (.Y(_216_),
    .A(net41),
    .B(net35));
 sg13g2_o21ai_1 _541_ (.B1(_216_),
    .Y(_019_),
    .A1(net41),
    .A2(net34));
 sg13g2_a22oi_1 _542_ (.Y(_217_),
    .B1(_212_),
    .B2(_064_),
    .A2(net35),
    .A1(net40));
 sg13g2_inv_1 _543_ (.Y(_020_),
    .A(_217_));
 sg13g2_nand2_1 _544_ (.Y(_218_),
    .A(net76),
    .B(net35));
 sg13g2_nand3_1 _545_ (.B(net40),
    .C(net76),
    .A(net41),
    .Y(_219_));
 sg13g2_xor2_1 _546_ (.B(_063_),
    .A(net76),
    .X(_220_));
 sg13g2_o21ai_1 _547_ (.B1(_218_),
    .Y(_021_),
    .A1(net34),
    .A2(_220_));
 sg13g2_nand2_1 _548_ (.Y(_221_),
    .A(net80),
    .B(net35));
 sg13g2_or2_1 _549_ (.X(_222_),
    .B(_063_),
    .A(_249_));
 sg13g2_xor2_1 _550_ (.B(_219_),
    .A(net80),
    .X(_223_));
 sg13g2_o21ai_1 _551_ (.B1(_221_),
    .Y(_022_),
    .A1(net34),
    .A2(_223_));
 sg13g2_nand2_1 _552_ (.Y(_224_),
    .A(net39),
    .B(net35));
 sg13g2_nor2_1 _553_ (.A(_242_),
    .B(_222_),
    .Y(_225_));
 sg13g2_xnor2_1 _554_ (.Y(_226_),
    .A(_242_),
    .B(_222_));
 sg13g2_o21ai_1 _555_ (.B1(_224_),
    .Y(_023_),
    .A1(net34),
    .A2(_226_));
 sg13g2_nand2_1 _556_ (.Y(_227_),
    .A(net64),
    .B(net35));
 sg13g2_and2_1 _557_ (.A(net38),
    .B(_225_),
    .X(_228_));
 sg13g2_xnor2_1 _558_ (.Y(_229_),
    .A(net38),
    .B(_225_));
 sg13g2_o21ai_1 _559_ (.B1(_227_),
    .Y(_024_),
    .A1(net34),
    .A2(_229_));
 sg13g2_nand2_1 _560_ (.Y(_230_),
    .A(net37),
    .B(net35));
 sg13g2_xnor2_1 _561_ (.Y(_231_),
    .A(net37),
    .B(_228_));
 sg13g2_o21ai_1 _562_ (.B1(_230_),
    .Y(_025_),
    .A1(net34),
    .A2(_231_));
 sg13g2_a21oi_1 _563_ (.A1(\hvsync_gen.vpos[6] ),
    .A2(_228_),
    .Y(_232_),
    .B1(net84));
 sg13g2_nor2_2 _564_ (.A(_258_),
    .B(_222_),
    .Y(_233_));
 sg13g2_nor3_1 _565_ (.A(net34),
    .B(_232_),
    .C(_233_),
    .Y(_234_));
 sg13g2_a21o_1 _566_ (.A2(_187_),
    .A1(net84),
    .B1(_234_),
    .X(_026_));
 sg13g2_a21oi_1 _567_ (.A1(net71),
    .A2(_233_),
    .Y(_235_),
    .B1(_214_));
 sg13g2_nor2_1 _568_ (.A(_187_),
    .B(_235_),
    .Y(_236_));
 sg13g2_a21oi_1 _569_ (.A1(_215_),
    .A2(_233_),
    .Y(_237_),
    .B1(net71));
 sg13g2_nor2_1 _570_ (.A(_236_),
    .B(net72),
    .Y(_027_));
 sg13g2_o21ai_1 _571_ (.B1(net68),
    .Y(_238_),
    .A1(_187_),
    .A2(_235_));
 sg13g2_nand3b_1 _572_ (.B(_233_),
    .C(\hvsync_gen.vpos[8] ),
    .Y(_239_),
    .A_N(net68));
 sg13g2_o21ai_1 _573_ (.B1(net69),
    .Y(_028_),
    .A1(_214_),
    .A2(_239_));
 sg13g2_dfrbpq_2 _574_ (.RESET_B(net49),
    .D(_002_),
    .Q(\abs_x[0] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _575_ (.RESET_B(net21),
    .D(_003_),
    .Q(\cx[1] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _576_ (.RESET_B(net20),
    .D(net67),
    .Q(\cx[2] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _577_ (.RESET_B(net19),
    .D(_005_),
    .Q(\cx[3] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _578_ (.RESET_B(net55),
    .D(_006_),
    .Q(\cx[4] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_2 _579_ (.RESET_B(net54),
    .D(_007_),
    .Q(\cx[5] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _580_ (.RESET_B(net53),
    .D(_008_),
    .Q(\hpos[6] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_2 _581_ (.RESET_B(net52),
    .D(_009_),
    .Q(\hpos[7] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _582_ (.RESET_B(net51),
    .D(_010_),
    .Q(\hpos[8] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _583_ (.RESET_B(net50),
    .D(net99),
    .Q(\hpos[9] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _584_ (.RESET_B(net46),
    .D(net57),
    .Q(\anim_offset[1] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_2 _585_ (.RESET_B(net46),
    .D(net59),
    .Q(\anim_offset[2] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_2 _586_ (.RESET_B(net46),
    .D(_014_),
    .Q(\anim_offset[3] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_2 _587_ (.RESET_B(net47),
    .D(net61),
    .Q(\anim_offset[4] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_2 _588_ (.RESET_B(net47),
    .D(_016_),
    .Q(\anim_offset[5] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_2 _589_ (.RESET_B(net47),
    .D(_017_),
    .Q(\anim_offset[6] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _590_ (.RESET_B(net47),
    .D(net63),
    .Q(\anim_offset[7] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _591_ (.RESET_B(net48),
    .D(net75),
    .Q(hsync),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_2 _592_ (.RESET_B(net32),
    .D(_019_),
    .Q(\abs_y[0] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_1 _593_ (.RESET_B(net30),
    .D(_020_),
    .Q(\cy[1] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_2 _594_ (.RESET_B(net28),
    .D(net77),
    .Q(\cy[2] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_2 _595_ (.RESET_B(net26),
    .D(net81),
    .Q(\cy[3] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_2 _596_ (.RESET_B(net24),
    .D(net101),
    .Q(\hvsync_gen.vpos[4] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _597_ (.RESET_B(net22),
    .D(_024_),
    .Q(\hvsync_gen.vpos[5] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_1 _598_ (.RESET_B(net29),
    .D(_025_),
    .Q(\hvsync_gen.vpos[6] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_2 _599_ (.RESET_B(net25),
    .D(net85),
    .Q(\hvsync_gen.vpos[7] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _600_ (.RESET_B(net31),
    .D(_027_),
    .Q(\hvsync_gen.vpos[8] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _601_ (.RESET_B(net27),
    .D(net70),
    .Q(\hvsync_gen.vpos[9] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_1 _602_ (.RESET_B(net23),
    .D(net91),
    .Q(\hvsync_gen.vsync ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_tiehi _576__20 (.L_HI(net20));
 sg13g2_tiehi _575__21 (.L_HI(net21));
 sg13g2_tiehi _597__22 (.L_HI(net22));
 sg13g2_tiehi _602__23 (.L_HI(net23));
 sg13g2_tiehi _596__24 (.L_HI(net24));
 sg13g2_tiehi _599__25 (.L_HI(net25));
 sg13g2_tiehi _595__26 (.L_HI(net26));
 sg13g2_tiehi _601__27 (.L_HI(net27));
 sg13g2_tiehi _594__28 (.L_HI(net28));
 sg13g2_tiehi _598__29 (.L_HI(net29));
 sg13g2_tiehi _593__30 (.L_HI(net30));
 sg13g2_tiehi _600__31 (.L_HI(net31));
 sg13g2_tiehi _592__32 (.L_HI(net32));
 sg13g2_tiehi _591__33 (.L_HI(net48));
 sg13g2_tiehi _574__34 (.L_HI(net49));
 sg13g2_tiehi _583__35 (.L_HI(net50));
 sg13g2_tiehi _582__36 (.L_HI(net51));
 sg13g2_tiehi _581__37 (.L_HI(net52));
 sg13g2_tiehi _580__38 (.L_HI(net53));
 sg13g2_tiehi _579__39 (.L_HI(net54));
 sg13g2_tiehi _578__40 (.L_HI(net55));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_matth_fischer_vgaTT_4 (.L_LO(net4));
 sg13g2_tielo tt_um_matth_fischer_vgaTT_5 (.L_LO(net5));
 sg13g2_tielo tt_um_matth_fischer_vgaTT_6 (.L_LO(net6));
 sg13g2_tielo tt_um_matth_fischer_vgaTT_7 (.L_LO(net7));
 sg13g2_tielo tt_um_matth_fischer_vgaTT_8 (.L_LO(net8));
 sg13g2_tielo tt_um_matth_fischer_vgaTT_9 (.L_LO(net9));
 sg13g2_tielo tt_um_matth_fischer_vgaTT_10 (.L_LO(net10));
 sg13g2_tielo tt_um_matth_fischer_vgaTT_11 (.L_LO(net11));
 sg13g2_tielo tt_um_matth_fischer_vgaTT_12 (.L_LO(net12));
 sg13g2_tielo tt_um_matth_fischer_vgaTT_13 (.L_LO(net13));
 sg13g2_tielo tt_um_matth_fischer_vgaTT_14 (.L_LO(net14));
 sg13g2_tielo tt_um_matth_fischer_vgaTT_15 (.L_LO(net15));
 sg13g2_tielo tt_um_matth_fischer_vgaTT_16 (.L_LO(net16));
 sg13g2_tielo tt_um_matth_fischer_vgaTT_17 (.L_LO(net17));
 sg13g2_tielo tt_um_matth_fischer_vgaTT_18 (.L_LO(net18));
 sg13g2_tiehi _577__19 (.L_HI(net19));
 sg13g2_buf_1 _641_ (.A(uo_out[5]),
    .X(uo_out[0]));
 sg13g2_buf_1 _642_ (.A(uo_out[6]),
    .X(uo_out[1]));
 sg13g2_buf_1 _643_ (.A(\hvsync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _644_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout33 (.A(_114_),
    .X(net33));
 sg13g2_buf_8 fanout34 (.A(_214_),
    .X(net34));
 sg13g2_buf_8 fanout35 (.A(_187_),
    .X(net35));
 sg13g2_buf_8 fanout36 (.A(_260_),
    .X(net36));
 sg13g2_buf_8 fanout37 (.A(net102),
    .X(net37));
 sg13g2_buf_8 fanout38 (.A(net64),
    .X(net38));
 sg13g2_buf_8 fanout39 (.A(net100),
    .X(net39));
 sg13g2_buf_8 fanout40 (.A(net89),
    .X(net40));
 sg13g2_buf_8 fanout41 (.A(net94),
    .X(net41));
 sg13g2_buf_8 fanout42 (.A(net98),
    .X(net42));
 sg13g2_buf_8 fanout43 (.A(net104),
    .X(net43));
 sg13g2_buf_8 fanout44 (.A(net78),
    .X(net44));
 sg13g2_buf_8 fanout45 (.A(net83),
    .X(net45));
 sg13g2_buf_8 fanout46 (.A(rst_n),
    .X(net46));
 sg13g2_buf_1 fanout47 (.A(rst_n),
    .X(net47));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_tielo tt_um_matth_fischer_vgaTT_3 (.L_LO(net3));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_3__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_3_6__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\anim_offset[1] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold2 (.A(_012_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold3 (.A(\anim_offset[2] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold4 (.A(_013_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold5 (.A(\anim_offset[4] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold6 (.A(_015_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold7 (.A(\anim_offset[7] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold8 (.A(_018_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold9 (.A(\hvsync_gen.vpos[5] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold10 (.A(\cx[2] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold11 (.A(_189_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold12 (.A(_004_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold13 (.A(\hvsync_gen.vpos[9] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold14 (.A(_238_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold15 (.A(_028_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold16 (.A(\hvsync_gen.vpos[8] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold17 (.A(_237_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold18 (.A(\hpos[7] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold19 (.A(_254_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold20 (.A(_000_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold21 (.A(\cy[2] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold22 (.A(_021_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold23 (.A(\hpos[6] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold24 (.A(_195_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold25 (.A(\cy[3] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold26 (.A(_022_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold27 (.A(\anim_offset[3] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold28 (.A(\abs_x[0] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold29 (.A(\hvsync_gen.vpos[7] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold30 (.A(_026_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold31 (.A(\cx[5] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold32 (.A(_193_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold33 (.A(\anim_offset[5] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold34 (.A(\cy[1] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold35 (.A(_251_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold36 (.A(_001_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold37 (.A(\cx[4] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold38 (.A(_191_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold39 (.A(\abs_y[0] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold40 (.A(\cx[3] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold41 (.A(_190_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold42 (.A(\anim_offset[6] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold43 (.A(\hpos[9] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold44 (.A(_011_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold45 (.A(\hvsync_gen.vpos[4] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold46 (.A(_023_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold47 (.A(\hvsync_gen.vpos[6] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold48 (.A(\cx[1] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold49 (.A(\hpos[8] ),
    .X(net104));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_4 FILLER_22_140 ();
 sg13g2_fill_2 FILLER_22_144 ();
 sg13g2_decap_8 FILLER_22_150 ();
 sg13g2_decap_8 FILLER_22_157 ();
 sg13g2_decap_8 FILLER_22_164 ();
 sg13g2_decap_8 FILLER_22_171 ();
 sg13g2_decap_8 FILLER_22_178 ();
 sg13g2_fill_2 FILLER_22_185 ();
 sg13g2_decap_8 FILLER_22_191 ();
 sg13g2_decap_8 FILLER_22_198 ();
 sg13g2_decap_4 FILLER_22_205 ();
 sg13g2_fill_2 FILLER_22_209 ();
 sg13g2_decap_8 FILLER_22_246 ();
 sg13g2_decap_8 FILLER_22_253 ();
 sg13g2_decap_8 FILLER_22_260 ();
 sg13g2_decap_8 FILLER_22_267 ();
 sg13g2_decap_8 FILLER_22_274 ();
 sg13g2_decap_8 FILLER_22_281 ();
 sg13g2_decap_8 FILLER_22_288 ();
 sg13g2_decap_8 FILLER_22_295 ();
 sg13g2_decap_8 FILLER_22_302 ();
 sg13g2_decap_8 FILLER_22_309 ();
 sg13g2_decap_8 FILLER_22_316 ();
 sg13g2_decap_8 FILLER_22_323 ();
 sg13g2_decap_8 FILLER_22_330 ();
 sg13g2_decap_8 FILLER_22_337 ();
 sg13g2_decap_8 FILLER_22_344 ();
 sg13g2_decap_8 FILLER_22_351 ();
 sg13g2_decap_8 FILLER_22_358 ();
 sg13g2_decap_8 FILLER_22_365 ();
 sg13g2_decap_8 FILLER_22_372 ();
 sg13g2_decap_8 FILLER_22_379 ();
 sg13g2_decap_8 FILLER_22_386 ();
 sg13g2_decap_8 FILLER_22_393 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_fill_1 FILLER_23_140 ();
 sg13g2_fill_2 FILLER_23_169 ();
 sg13g2_fill_2 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_293 ();
 sg13g2_decap_8 FILLER_23_300 ();
 sg13g2_decap_8 FILLER_23_307 ();
 sg13g2_decap_8 FILLER_23_314 ();
 sg13g2_decap_8 FILLER_23_321 ();
 sg13g2_decap_8 FILLER_23_328 ();
 sg13g2_decap_8 FILLER_23_335 ();
 sg13g2_decap_8 FILLER_23_342 ();
 sg13g2_decap_8 FILLER_23_349 ();
 sg13g2_decap_8 FILLER_23_356 ();
 sg13g2_decap_8 FILLER_23_363 ();
 sg13g2_decap_8 FILLER_23_370 ();
 sg13g2_decap_8 FILLER_23_377 ();
 sg13g2_decap_8 FILLER_23_384 ();
 sg13g2_decap_8 FILLER_23_391 ();
 sg13g2_decap_8 FILLER_23_398 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_4 FILLER_24_133 ();
 sg13g2_fill_1 FILLER_24_137 ();
 sg13g2_decap_4 FILLER_24_141 ();
 sg13g2_fill_1 FILLER_24_145 ();
 sg13g2_fill_2 FILLER_24_160 ();
 sg13g2_fill_2 FILLER_24_179 ();
 sg13g2_fill_1 FILLER_24_181 ();
 sg13g2_fill_2 FILLER_24_195 ();
 sg13g2_decap_4 FILLER_24_219 ();
 sg13g2_fill_2 FILLER_24_276 ();
 sg13g2_fill_1 FILLER_24_300 ();
 sg13g2_decap_8 FILLER_24_314 ();
 sg13g2_decap_8 FILLER_24_321 ();
 sg13g2_decap_8 FILLER_24_328 ();
 sg13g2_decap_8 FILLER_24_335 ();
 sg13g2_decap_8 FILLER_24_342 ();
 sg13g2_decap_8 FILLER_24_349 ();
 sg13g2_decap_8 FILLER_24_356 ();
 sg13g2_decap_8 FILLER_24_363 ();
 sg13g2_decap_8 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_377 ();
 sg13g2_decap_8 FILLER_24_384 ();
 sg13g2_decap_8 FILLER_24_391 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_fill_2 FILLER_25_119 ();
 sg13g2_decap_4 FILLER_25_195 ();
 sg13g2_fill_1 FILLER_25_199 ();
 sg13g2_fill_1 FILLER_25_240 ();
 sg13g2_fill_2 FILLER_25_296 ();
 sg13g2_decap_8 FILLER_25_326 ();
 sg13g2_decap_8 FILLER_25_333 ();
 sg13g2_decap_8 FILLER_25_340 ();
 sg13g2_decap_8 FILLER_25_347 ();
 sg13g2_decap_8 FILLER_25_354 ();
 sg13g2_decap_8 FILLER_25_361 ();
 sg13g2_decap_8 FILLER_25_368 ();
 sg13g2_decap_8 FILLER_25_375 ();
 sg13g2_decap_8 FILLER_25_382 ();
 sg13g2_decap_8 FILLER_25_389 ();
 sg13g2_decap_8 FILLER_25_396 ();
 sg13g2_decap_4 FILLER_25_403 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_fill_2 FILLER_26_137 ();
 sg13g2_decap_8 FILLER_26_143 ();
 sg13g2_decap_4 FILLER_26_150 ();
 sg13g2_fill_1 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_181 ();
 sg13g2_decap_4 FILLER_26_188 ();
 sg13g2_decap_4 FILLER_26_223 ();
 sg13g2_fill_1 FILLER_26_227 ();
 sg13g2_fill_2 FILLER_26_238 ();
 sg13g2_fill_1 FILLER_26_246 ();
 sg13g2_fill_2 FILLER_26_252 ();
 sg13g2_fill_1 FILLER_26_254 ();
 sg13g2_fill_2 FILLER_26_259 ();
 sg13g2_decap_4 FILLER_26_266 ();
 sg13g2_fill_1 FILLER_26_270 ();
 sg13g2_decap_8 FILLER_26_296 ();
 sg13g2_fill_2 FILLER_26_303 ();
 sg13g2_fill_1 FILLER_26_305 ();
 sg13g2_decap_8 FILLER_26_310 ();
 sg13g2_decap_8 FILLER_26_317 ();
 sg13g2_decap_8 FILLER_26_324 ();
 sg13g2_decap_8 FILLER_26_331 ();
 sg13g2_decap_8 FILLER_26_338 ();
 sg13g2_decap_8 FILLER_26_345 ();
 sg13g2_decap_8 FILLER_26_352 ();
 sg13g2_decap_8 FILLER_26_359 ();
 sg13g2_decap_8 FILLER_26_366 ();
 sg13g2_decap_8 FILLER_26_373 ();
 sg13g2_decap_8 FILLER_26_380 ();
 sg13g2_decap_8 FILLER_26_387 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_fill_2 FILLER_27_98 ();
 sg13g2_fill_1 FILLER_27_100 ();
 sg13g2_decap_8 FILLER_27_106 ();
 sg13g2_decap_8 FILLER_27_113 ();
 sg13g2_fill_2 FILLER_27_120 ();
 sg13g2_fill_1 FILLER_27_122 ();
 sg13g2_decap_8 FILLER_27_131 ();
 sg13g2_decap_8 FILLER_27_138 ();
 sg13g2_decap_8 FILLER_27_145 ();
 sg13g2_fill_1 FILLER_27_152 ();
 sg13g2_decap_4 FILLER_27_175 ();
 sg13g2_fill_2 FILLER_27_179 ();
 sg13g2_fill_2 FILLER_27_198 ();
 sg13g2_fill_1 FILLER_27_200 ();
 sg13g2_decap_8 FILLER_27_209 ();
 sg13g2_decap_4 FILLER_27_238 ();
 sg13g2_fill_2 FILLER_27_274 ();
 sg13g2_fill_2 FILLER_27_285 ();
 sg13g2_decap_8 FILLER_27_327 ();
 sg13g2_decap_8 FILLER_27_334 ();
 sg13g2_decap_8 FILLER_27_341 ();
 sg13g2_decap_8 FILLER_27_348 ();
 sg13g2_decap_8 FILLER_27_355 ();
 sg13g2_decap_8 FILLER_27_362 ();
 sg13g2_decap_8 FILLER_27_369 ();
 sg13g2_decap_8 FILLER_27_376 ();
 sg13g2_decap_8 FILLER_27_383 ();
 sg13g2_decap_8 FILLER_27_390 ();
 sg13g2_decap_8 FILLER_27_397 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_fill_2 FILLER_28_112 ();
 sg13g2_fill_1 FILLER_28_114 ();
 sg13g2_decap_4 FILLER_28_147 ();
 sg13g2_fill_2 FILLER_28_205 ();
 sg13g2_decap_4 FILLER_28_224 ();
 sg13g2_decap_4 FILLER_28_239 ();
 sg13g2_fill_2 FILLER_28_243 ();
 sg13g2_fill_1 FILLER_28_250 ();
 sg13g2_decap_8 FILLER_28_256 ();
 sg13g2_decap_8 FILLER_28_300 ();
 sg13g2_fill_2 FILLER_28_307 ();
 sg13g2_fill_2 FILLER_28_321 ();
 sg13g2_decap_8 FILLER_28_341 ();
 sg13g2_decap_8 FILLER_28_348 ();
 sg13g2_decap_8 FILLER_28_355 ();
 sg13g2_decap_8 FILLER_28_362 ();
 sg13g2_decap_8 FILLER_28_369 ();
 sg13g2_decap_8 FILLER_28_376 ();
 sg13g2_decap_8 FILLER_28_383 ();
 sg13g2_decap_8 FILLER_28_390 ();
 sg13g2_decap_8 FILLER_28_397 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_4 FILLER_29_70 ();
 sg13g2_fill_1 FILLER_29_74 ();
 sg13g2_fill_2 FILLER_29_96 ();
 sg13g2_fill_1 FILLER_29_98 ();
 sg13g2_fill_2 FILLER_29_121 ();
 sg13g2_fill_1 FILLER_29_123 ();
 sg13g2_decap_8 FILLER_29_128 ();
 sg13g2_fill_2 FILLER_29_135 ();
 sg13g2_fill_1 FILLER_29_173 ();
 sg13g2_fill_2 FILLER_29_193 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_fill_2 FILLER_29_217 ();
 sg13g2_fill_1 FILLER_29_235 ();
 sg13g2_decap_4 FILLER_29_254 ();
 sg13g2_fill_2 FILLER_29_266 ();
 sg13g2_fill_2 FILLER_29_272 ();
 sg13g2_decap_8 FILLER_29_279 ();
 sg13g2_fill_2 FILLER_29_329 ();
 sg13g2_fill_1 FILLER_29_331 ();
 sg13g2_fill_1 FILLER_29_341 ();
 sg13g2_decap_8 FILLER_29_351 ();
 sg13g2_decap_8 FILLER_29_358 ();
 sg13g2_decap_8 FILLER_29_365 ();
 sg13g2_decap_8 FILLER_29_372 ();
 sg13g2_decap_8 FILLER_29_379 ();
 sg13g2_decap_8 FILLER_29_386 ();
 sg13g2_decap_8 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_400 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_fill_1 FILLER_30_70 ();
 sg13g2_fill_2 FILLER_30_99 ();
 sg13g2_fill_1 FILLER_30_101 ();
 sg13g2_fill_2 FILLER_30_111 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_fill_1 FILLER_30_133 ();
 sg13g2_fill_2 FILLER_30_142 ();
 sg13g2_decap_4 FILLER_30_173 ();
 sg13g2_fill_1 FILLER_30_187 ();
 sg13g2_fill_2 FILLER_30_196 ();
 sg13g2_fill_1 FILLER_30_198 ();
 sg13g2_fill_1 FILLER_30_209 ();
 sg13g2_fill_2 FILLER_30_220 ();
 sg13g2_decap_8 FILLER_30_235 ();
 sg13g2_decap_4 FILLER_30_242 ();
 sg13g2_fill_1 FILLER_30_246 ();
 sg13g2_fill_2 FILLER_30_255 ();
 sg13g2_decap_8 FILLER_30_265 ();
 sg13g2_fill_2 FILLER_30_272 ();
 sg13g2_decap_8 FILLER_30_282 ();
 sg13g2_fill_2 FILLER_30_289 ();
 sg13g2_fill_1 FILLER_30_291 ();
 sg13g2_fill_1 FILLER_30_297 ();
 sg13g2_fill_2 FILLER_30_310 ();
 sg13g2_fill_2 FILLER_30_321 ();
 sg13g2_fill_1 FILLER_30_323 ();
 sg13g2_decap_8 FILLER_30_360 ();
 sg13g2_decap_8 FILLER_30_367 ();
 sg13g2_decap_8 FILLER_30_374 ();
 sg13g2_decap_8 FILLER_30_381 ();
 sg13g2_decap_8 FILLER_30_388 ();
 sg13g2_decap_8 FILLER_30_395 ();
 sg13g2_decap_8 FILLER_30_402 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_fill_2 FILLER_31_77 ();
 sg13g2_fill_1 FILLER_31_79 ();
 sg13g2_decap_4 FILLER_31_108 ();
 sg13g2_decap_8 FILLER_31_159 ();
 sg13g2_decap_8 FILLER_31_166 ();
 sg13g2_decap_4 FILLER_31_173 ();
 sg13g2_fill_1 FILLER_31_177 ();
 sg13g2_fill_2 FILLER_31_183 ();
 sg13g2_decap_4 FILLER_31_190 ();
 sg13g2_fill_1 FILLER_31_194 ();
 sg13g2_fill_2 FILLER_31_240 ();
 sg13g2_fill_1 FILLER_31_242 ();
 sg13g2_decap_4 FILLER_31_260 ();
 sg13g2_fill_1 FILLER_31_264 ();
 sg13g2_decap_8 FILLER_31_282 ();
 sg13g2_decap_4 FILLER_31_289 ();
 sg13g2_fill_1 FILLER_31_293 ();
 sg13g2_fill_2 FILLER_31_304 ();
 sg13g2_fill_2 FILLER_31_318 ();
 sg13g2_decap_8 FILLER_31_324 ();
 sg13g2_decap_8 FILLER_31_367 ();
 sg13g2_decap_8 FILLER_31_374 ();
 sg13g2_decap_8 FILLER_31_381 ();
 sg13g2_decap_8 FILLER_31_388 ();
 sg13g2_decap_8 FILLER_31_395 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_4 FILLER_32_70 ();
 sg13g2_fill_1 FILLER_32_74 ();
 sg13g2_decap_4 FILLER_32_79 ();
 sg13g2_fill_2 FILLER_32_83 ();
 sg13g2_decap_4 FILLER_32_89 ();
 sg13g2_fill_2 FILLER_32_93 ();
 sg13g2_fill_2 FILLER_32_130 ();
 sg13g2_decap_8 FILLER_32_136 ();
 sg13g2_fill_2 FILLER_32_143 ();
 sg13g2_decap_8 FILLER_32_159 ();
 sg13g2_fill_1 FILLER_32_166 ();
 sg13g2_decap_4 FILLER_32_178 ();
 sg13g2_fill_2 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_fill_2 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_fill_2 FILLER_32_231 ();
 sg13g2_decap_4 FILLER_32_237 ();
 sg13g2_decap_4 FILLER_32_245 ();
 sg13g2_fill_2 FILLER_32_253 ();
 sg13g2_fill_1 FILLER_32_255 ();
 sg13g2_decap_4 FILLER_32_260 ();
 sg13g2_fill_2 FILLER_32_264 ();
 sg13g2_fill_1 FILLER_32_272 ();
 sg13g2_decap_8 FILLER_32_281 ();
 sg13g2_fill_1 FILLER_32_288 ();
 sg13g2_decap_8 FILLER_32_301 ();
 sg13g2_fill_2 FILLER_32_308 ();
 sg13g2_fill_1 FILLER_32_333 ();
 sg13g2_fill_1 FILLER_32_339 ();
 sg13g2_decap_8 FILLER_32_365 ();
 sg13g2_decap_8 FILLER_32_372 ();
 sg13g2_decap_8 FILLER_32_379 ();
 sg13g2_decap_8 FILLER_32_386 ();
 sg13g2_decap_8 FILLER_32_393 ();
 sg13g2_decap_8 FILLER_32_400 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_4 FILLER_33_98 ();
 sg13g2_fill_2 FILLER_33_134 ();
 sg13g2_fill_2 FILLER_33_143 ();
 sg13g2_fill_1 FILLER_33_145 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_fill_2 FILLER_33_161 ();
 sg13g2_fill_2 FILLER_33_178 ();
 sg13g2_fill_1 FILLER_33_180 ();
 sg13g2_fill_2 FILLER_33_204 ();
 sg13g2_decap_4 FILLER_33_221 ();
 sg13g2_fill_2 FILLER_33_240 ();
 sg13g2_fill_1 FILLER_33_242 ();
 sg13g2_fill_1 FILLER_33_253 ();
 sg13g2_fill_2 FILLER_33_263 ();
 sg13g2_decap_8 FILLER_33_270 ();
 sg13g2_decap_8 FILLER_33_277 ();
 sg13g2_fill_1 FILLER_33_284 ();
 sg13g2_decap_8 FILLER_33_307 ();
 sg13g2_fill_2 FILLER_33_314 ();
 sg13g2_decap_8 FILLER_33_329 ();
 sg13g2_fill_2 FILLER_33_336 ();
 sg13g2_fill_1 FILLER_33_346 ();
 sg13g2_decap_8 FILLER_33_375 ();
 sg13g2_decap_8 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_33_389 ();
 sg13g2_decap_8 FILLER_33_396 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_fill_1 FILLER_34_70 ();
 sg13g2_fill_2 FILLER_34_129 ();
 sg13g2_fill_2 FILLER_34_147 ();
 sg13g2_fill_1 FILLER_34_149 ();
 sg13g2_decap_8 FILLER_34_178 ();
 sg13g2_fill_1 FILLER_34_185 ();
 sg13g2_fill_2 FILLER_34_194 ();
 sg13g2_fill_1 FILLER_34_196 ();
 sg13g2_decap_4 FILLER_34_206 ();
 sg13g2_fill_2 FILLER_34_214 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_decap_8 FILLER_34_237 ();
 sg13g2_decap_8 FILLER_34_244 ();
 sg13g2_decap_4 FILLER_34_251 ();
 sg13g2_fill_1 FILLER_34_255 ();
 sg13g2_fill_1 FILLER_34_261 ();
 sg13g2_decap_8 FILLER_34_278 ();
 sg13g2_fill_2 FILLER_34_285 ();
 sg13g2_fill_1 FILLER_34_287 ();
 sg13g2_decap_8 FILLER_34_304 ();
 sg13g2_decap_8 FILLER_34_311 ();
 sg13g2_decap_8 FILLER_34_318 ();
 sg13g2_fill_1 FILLER_34_341 ();
 sg13g2_decap_8 FILLER_34_373 ();
 sg13g2_decap_8 FILLER_34_380 ();
 sg13g2_decap_8 FILLER_34_387 ();
 sg13g2_decap_8 FILLER_34_394 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_4 FILLER_35_70 ();
 sg13g2_fill_2 FILLER_35_74 ();
 sg13g2_decap_4 FILLER_35_80 ();
 sg13g2_fill_1 FILLER_35_84 ();
 sg13g2_fill_2 FILLER_35_135 ();
 sg13g2_fill_2 FILLER_35_145 ();
 sg13g2_fill_1 FILLER_35_147 ();
 sg13g2_fill_1 FILLER_35_167 ();
 sg13g2_fill_2 FILLER_35_181 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_4 FILLER_35_203 ();
 sg13g2_fill_1 FILLER_35_207 ();
 sg13g2_decap_4 FILLER_35_213 ();
 sg13g2_fill_1 FILLER_35_229 ();
 sg13g2_fill_2 FILLER_35_238 ();
 sg13g2_decap_8 FILLER_35_257 ();
 sg13g2_decap_4 FILLER_35_264 ();
 sg13g2_decap_8 FILLER_35_272 ();
 sg13g2_decap_4 FILLER_35_279 ();
 sg13g2_fill_2 FILLER_35_283 ();
 sg13g2_fill_2 FILLER_35_293 ();
 sg13g2_decap_4 FILLER_35_308 ();
 sg13g2_fill_1 FILLER_35_312 ();
 sg13g2_fill_1 FILLER_35_330 ();
 sg13g2_fill_2 FILLER_35_339 ();
 sg13g2_decap_8 FILLER_35_373 ();
 sg13g2_decap_8 FILLER_35_380 ();
 sg13g2_decap_8 FILLER_35_387 ();
 sg13g2_decap_8 FILLER_35_394 ();
 sg13g2_decap_8 FILLER_35_401 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_fill_1 FILLER_36_70 ();
 sg13g2_fill_1 FILLER_36_99 ();
 sg13g2_fill_2 FILLER_36_124 ();
 sg13g2_fill_2 FILLER_36_135 ();
 sg13g2_fill_1 FILLER_36_137 ();
 sg13g2_fill_2 FILLER_36_147 ();
 sg13g2_fill_2 FILLER_36_180 ();
 sg13g2_decap_8 FILLER_36_190 ();
 sg13g2_decap_8 FILLER_36_197 ();
 sg13g2_fill_1 FILLER_36_204 ();
 sg13g2_decap_4 FILLER_36_218 ();
 sg13g2_decap_8 FILLER_36_235 ();
 sg13g2_decap_4 FILLER_36_242 ();
 sg13g2_fill_1 FILLER_36_246 ();
 sg13g2_decap_4 FILLER_36_261 ();
 sg13g2_fill_1 FILLER_36_265 ();
 sg13g2_decap_4 FILLER_36_274 ();
 sg13g2_fill_2 FILLER_36_278 ();
 sg13g2_fill_2 FILLER_36_285 ();
 sg13g2_fill_1 FILLER_36_292 ();
 sg13g2_decap_8 FILLER_36_298 ();
 sg13g2_decap_8 FILLER_36_305 ();
 sg13g2_decap_4 FILLER_36_344 ();
 sg13g2_fill_1 FILLER_36_348 ();
 sg13g2_decap_8 FILLER_36_367 ();
 sg13g2_decap_8 FILLER_36_374 ();
 sg13g2_decap_8 FILLER_36_381 ();
 sg13g2_decap_8 FILLER_36_388 ();
 sg13g2_decap_8 FILLER_36_395 ();
 sg13g2_decap_8 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_fill_2 FILLER_37_63 ();
 sg13g2_fill_1 FILLER_37_65 ();
 sg13g2_fill_2 FILLER_37_124 ();
 sg13g2_fill_1 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_4 FILLER_37_210 ();
 sg13g2_decap_4 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_232 ();
 sg13g2_decap_8 FILLER_37_239 ();
 sg13g2_decap_8 FILLER_37_246 ();
 sg13g2_decap_4 FILLER_37_253 ();
 sg13g2_fill_2 FILLER_37_273 ();
 sg13g2_fill_1 FILLER_37_275 ();
 sg13g2_fill_2 FILLER_37_281 ();
 sg13g2_fill_1 FILLER_37_283 ();
 sg13g2_decap_4 FILLER_37_307 ();
 sg13g2_fill_1 FILLER_37_311 ();
 sg13g2_fill_1 FILLER_37_320 ();
 sg13g2_fill_2 FILLER_37_344 ();
 sg13g2_fill_1 FILLER_37_346 ();
 sg13g2_decap_8 FILLER_37_375 ();
 sg13g2_decap_8 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_37_396 ();
 sg13g2_decap_4 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_fill_2 FILLER_38_49 ();
 sg13g2_fill_2 FILLER_38_115 ();
 sg13g2_fill_2 FILLER_38_126 ();
 sg13g2_fill_2 FILLER_38_148 ();
 sg13g2_fill_2 FILLER_38_158 ();
 sg13g2_fill_2 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_218 ();
 sg13g2_fill_1 FILLER_38_222 ();
 sg13g2_decap_8 FILLER_38_254 ();
 sg13g2_fill_2 FILLER_38_261 ();
 sg13g2_fill_1 FILLER_38_263 ();
 sg13g2_fill_2 FILLER_38_268 ();
 sg13g2_decap_8 FILLER_38_282 ();
 sg13g2_decap_8 FILLER_38_289 ();
 sg13g2_fill_2 FILLER_38_296 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_315 ();
 sg13g2_decap_4 FILLER_38_322 ();
 sg13g2_decap_4 FILLER_38_330 ();
 sg13g2_decap_8 FILLER_38_378 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net3;
 assign uio_oe[1] = net4;
 assign uio_oe[2] = net5;
 assign uio_oe[3] = net6;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_oe[7] = net10;
 assign uio_out[0] = net11;
 assign uio_out[1] = net12;
 assign uio_out[2] = net13;
 assign uio_out[3] = net14;
 assign uio_out[4] = net15;
 assign uio_out[5] = net16;
 assign uio_out[6] = net17;
 assign uio_out[7] = net18;
endmodule
