module tt_um_not_a_dinosaur (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire clknet_0_clk;
 wire \dinosaur_y_pos[0] ;
 wire \dinosaur_y_pos[1] ;
 wire \dinosaur_y_pos[2] ;
 wire \dinosaur_y_pos[3] ;
 wire \dinosaur_y_pos[4] ;
 wire \dinosaur_y_pos[5] ;
 wire \dinosaur_y_pos[6] ;
 wire \dinosaur_y_pos[7] ;
 wire \dinosaur_y_pos[8] ;
 wire \dinosaur_y_pos[9] ;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire \jump_counter[0] ;
 wire \jump_counter[10] ;
 wire \jump_counter[11] ;
 wire \jump_counter[12] ;
 wire \jump_counter[13] ;
 wire \jump_counter[14] ;
 wire \jump_counter[15] ;
 wire \jump_counter[16] ;
 wire \jump_counter[17] ;
 wire \jump_counter[18] ;
 wire \jump_counter[19] ;
 wire \jump_counter[1] ;
 wire \jump_counter[20] ;
 wire \jump_counter[21] ;
 wire \jump_counter[22] ;
 wire \jump_counter[23] ;
 wire \jump_counter[2] ;
 wire \jump_counter[3] ;
 wire \jump_counter[4] ;
 wire \jump_counter[5] ;
 wire \jump_counter[6] ;
 wire \jump_counter[7] ;
 wire \jump_counter[8] ;
 wire \jump_counter[9] ;
 wire \jump_state[0] ;
 wire \jump_state[1] ;
 wire \jump_state[2] ;
 wire \jump_state[3] ;
 wire prev_button_state;
 wire \square_counter[0] ;
 wire \square_counter[10] ;
 wire \square_counter[11] ;
 wire \square_counter[12] ;
 wire \square_counter[13] ;
 wire \square_counter[14] ;
 wire \square_counter[15] ;
 wire \square_counter[16] ;
 wire \square_counter[17] ;
 wire \square_counter[18] ;
 wire \square_counter[19] ;
 wire \square_counter[1] ;
 wire \square_counter[20] ;
 wire \square_counter[21] ;
 wire \square_counter[22] ;
 wire \square_counter[23] ;
 wire \square_counter[2] ;
 wire \square_counter[3] ;
 wire \square_counter[4] ;
 wire \square_counter[5] ;
 wire \square_counter[6] ;
 wire \square_counter[7] ;
 wire \square_counter[8] ;
 wire \square_counter[9] ;
 wire \square_x_pos[0] ;
 wire \square_x_pos[1] ;
 wire \square_x_pos[2] ;
 wire \square_x_pos[3] ;
 wire \square_x_pos[4] ;
 wire \square_x_pos[5] ;
 wire \square_x_pos[6] ;
 wire \square_x_pos[7] ;
 wire \square_x_pos[8] ;
 wire \square_x_pos[9] ;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net1;
 wire net2;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;

 sg13g2_inv_1 _0615_ (.Y(_0094_),
    .A(net194));
 sg13g2_inv_1 _0616_ (.Y(_0095_),
    .A(net234));
 sg13g2_inv_2 _0617_ (.Y(_0096_),
    .A(\square_x_pos[6] ));
 sg13g2_inv_1 _0618_ (.Y(_0097_),
    .A(\square_x_pos[5] ));
 sg13g2_inv_2 _0619_ (.Y(_0098_),
    .A(net303));
 sg13g2_inv_1 _0620_ (.Y(_0099_),
    .A(\square_x_pos[3] ));
 sg13g2_inv_1 _0621_ (.Y(_0100_),
    .A(net297));
 sg13g2_inv_1 _0622_ (.Y(_0101_),
    .A(net187));
 sg13g2_inv_1 _0623_ (.Y(_0102_),
    .A(net200));
 sg13g2_inv_1 _0624_ (.Y(_0103_),
    .A(net214));
 sg13g2_inv_2 _0625_ (.Y(_0104_),
    .A(net298));
 sg13g2_inv_1 _0626_ (.Y(_0105_),
    .A(\jump_counter[9] ));
 sg13g2_inv_1 _0627_ (.Y(_0106_),
    .A(net261));
 sg13g2_inv_2 _0628_ (.Y(_0107_),
    .A(\dinosaur_y_pos[7] ));
 sg13g2_inv_2 _0629_ (.Y(_0108_),
    .A(\dinosaur_y_pos[6] ));
 sg13g2_inv_1 _0630_ (.Y(_0109_),
    .A(\dinosaur_y_pos[4] ));
 sg13g2_inv_1 _0631_ (.Y(_0110_),
    .A(\dinosaur_y_pos[3] ));
 sg13g2_inv_1 _0632_ (.Y(_0111_),
    .A(net275));
 sg13g2_inv_1 _0633_ (.Y(_0112_),
    .A(\square_counter[15] ));
 sg13g2_inv_1 _0634_ (.Y(_0113_),
    .A(\square_counter[11] ));
 sg13g2_inv_1 _0635_ (.Y(_0114_),
    .A(net300));
 sg13g2_inv_1 _0636_ (.Y(_0115_),
    .A(net204));
 sg13g2_inv_1 _0637_ (.Y(_0116_),
    .A(net156));
 sg13g2_inv_1 _0638_ (.Y(_0117_),
    .A(net62));
 sg13g2_inv_2 _0639_ (.Y(_0118_),
    .A(net279));
 sg13g2_inv_2 _0640_ (.Y(_0119_),
    .A(net263));
 sg13g2_inv_1 _0641_ (.Y(_0120_),
    .A(net211));
 sg13g2_inv_2 _0642_ (.Y(_0121_),
    .A(net232));
 sg13g2_inv_1 _0643_ (.Y(_0122_),
    .A(\hvsync_gen.hpos[1] ));
 sg13g2_inv_1 _0644_ (.Y(_0123_),
    .A(net56));
 sg13g2_inv_4 _0645_ (.A(\hvsync_gen.hpos[2] ),
    .Y(_0124_));
 sg13g2_inv_1 _0646_ (.Y(_0125_),
    .A(\hvsync_gen.hpos[7] ));
 sg13g2_inv_1 _0647_ (.Y(_0126_),
    .A(\hvsync_gen.hpos[6] ));
 sg13g2_inv_1 _0648_ (.Y(_0127_),
    .A(\hvsync_gen.hpos[4] ));
 sg13g2_nand3_1 _0649_ (.B(net52),
    .C(net211),
    .A(net263),
    .Y(_0128_));
 sg13g2_and2_1 _0650_ (.A(net267),
    .B(net245),
    .X(_0129_));
 sg13g2_o21ai_1 _0651_ (.B1(net267),
    .Y(_0130_),
    .A1(net245),
    .A2(net53));
 sg13g2_or4_1 _0652_ (.A(net232),
    .B(net209),
    .C(_0129_),
    .D(_0130_),
    .X(_0131_));
 sg13g2_nor3_1 _0653_ (.A(_0118_),
    .B(_0128_),
    .C(_0131_),
    .Y(_0001_));
 sg13g2_and3_1 _0654_ (.X(_0132_),
    .A(\hvsync_gen.hpos[6] ),
    .B(net55),
    .C(\hvsync_gen.hpos[4] ));
 sg13g2_nor3_1 _0655_ (.A(\hvsync_gen.hpos[6] ),
    .B(net55),
    .C(\hvsync_gen.hpos[4] ),
    .Y(_0133_));
 sg13g2_nand2_1 _0656_ (.Y(_0134_),
    .A(\hvsync_gen.hpos[9] ),
    .B(\hvsync_gen.hpos[7] ));
 sg13g2_nor4_1 _0657_ (.A(net198),
    .B(_0132_),
    .C(_0133_),
    .D(_0134_),
    .Y(_0000_));
 sg13g2_and2_1 _0658_ (.A(\dinosaur_y_pos[5] ),
    .B(\dinosaur_y_pos[4] ),
    .X(_0135_));
 sg13g2_nand3_1 _0659_ (.B(\dinosaur_y_pos[5] ),
    .C(\dinosaur_y_pos[4] ),
    .A(\dinosaur_y_pos[6] ),
    .Y(_0136_));
 sg13g2_xnor2_1 _0660_ (.Y(_0137_),
    .A(\dinosaur_y_pos[6] ),
    .B(_0135_));
 sg13g2_or2_1 _0661_ (.X(_0138_),
    .B(_0137_),
    .A(net52));
 sg13g2_nor2_1 _0662_ (.A(\dinosaur_y_pos[5] ),
    .B(\dinosaur_y_pos[4] ),
    .Y(_0139_));
 sg13g2_o21ai_1 _0663_ (.B1(\hvsync_gen.vpos[5] ),
    .Y(_0140_),
    .A1(_0135_),
    .A2(_0139_));
 sg13g2_xor2_1 _0664_ (.B(\hvsync_gen.vpos[4] ),
    .A(\dinosaur_y_pos[4] ),
    .X(_0141_));
 sg13g2_or3_1 _0665_ (.A(\hvsync_gen.vpos[5] ),
    .B(_0135_),
    .C(_0139_),
    .X(_0142_));
 sg13g2_nand3_1 _0666_ (.B(_0141_),
    .C(_0142_),
    .A(_0140_),
    .Y(_0143_));
 sg13g2_nor2_1 _0667_ (.A(_0110_),
    .B(\hvsync_gen.vpos[3] ),
    .Y(_0144_));
 sg13g2_nor2b_1 _0668_ (.A(\dinosaur_y_pos[2] ),
    .B_N(\hvsync_gen.vpos[2] ),
    .Y(_0145_));
 sg13g2_xnor2_1 _0669_ (.Y(_0146_),
    .A(\dinosaur_y_pos[2] ),
    .B(\hvsync_gen.vpos[2] ));
 sg13g2_nor2b_1 _0670_ (.A(\dinosaur_y_pos[1] ),
    .B_N(net53),
    .Y(_0147_));
 sg13g2_nand2b_2 _0671_ (.Y(_0148_),
    .B(\dinosaur_y_pos[0] ),
    .A_N(net54));
 sg13g2_xnor2_1 _0672_ (.Y(_0149_),
    .A(\dinosaur_y_pos[1] ),
    .B(net53));
 sg13g2_a21o_2 _0673_ (.A2(_0149_),
    .A1(_0148_),
    .B1(_0147_),
    .X(_0150_));
 sg13g2_a21o_1 _0674_ (.A2(_0150_),
    .A1(_0146_),
    .B1(_0145_),
    .X(_0151_));
 sg13g2_a221oi_1 _0675_ (.B2(_0150_),
    .C1(_0145_),
    .B1(_0146_),
    .A1(_0110_),
    .Y(_0152_),
    .A2(\hvsync_gen.vpos[3] ));
 sg13g2_nor3_1 _0676_ (.A(_0143_),
    .B(_0144_),
    .C(_0152_),
    .Y(_0153_));
 sg13g2_o21ai_1 _0677_ (.B1(_0140_),
    .Y(_0154_),
    .A1(_0109_),
    .A2(_0121_));
 sg13g2_and2_1 _0678_ (.A(_0142_),
    .B(_0154_),
    .X(_0155_));
 sg13g2_o21ai_1 _0679_ (.B1(_0138_),
    .Y(_0156_),
    .A1(_0153_),
    .A2(_0155_));
 sg13g2_nor2_2 _0680_ (.A(_0107_),
    .B(_0136_),
    .Y(_0157_));
 sg13g2_xnor2_1 _0681_ (.Y(_0158_),
    .A(_0107_),
    .B(_0136_));
 sg13g2_a22oi_1 _0682_ (.Y(_0159_),
    .B1(_0158_),
    .B2(\hvsync_gen.vpos[7] ),
    .A2(_0137_),
    .A1(net52));
 sg13g2_nand2_1 _0683_ (.Y(_0160_),
    .A(net57),
    .B(_0157_));
 sg13g2_xnor2_1 _0684_ (.Y(_0161_),
    .A(net57),
    .B(_0157_));
 sg13g2_nand2b_1 _0685_ (.Y(_0162_),
    .B(_0119_),
    .A_N(_0158_));
 sg13g2_o21ai_1 _0686_ (.B1(_0162_),
    .Y(_0163_),
    .A1(\hvsync_gen.vpos[8] ),
    .A2(_0161_));
 sg13g2_a21o_1 _0687_ (.A2(_0159_),
    .A1(_0156_),
    .B1(_0163_),
    .X(_0164_));
 sg13g2_xnor2_1 _0688_ (.Y(_0165_),
    .A(_0106_),
    .B(_0160_));
 sg13g2_a22oi_1 _0689_ (.Y(_0166_),
    .B1(_0165_),
    .B2(\hvsync_gen.vpos[9] ),
    .A2(_0161_),
    .A1(\hvsync_gen.vpos[8] ));
 sg13g2_nor2b_1 _0690_ (.A(\dinosaur_y_pos[9] ),
    .B_N(\hvsync_gen.vpos[9] ),
    .Y(_0167_));
 sg13g2_nor2_1 _0691_ (.A(_0160_),
    .B(_0167_),
    .Y(_0168_));
 sg13g2_nor2_1 _0692_ (.A(_0106_),
    .B(\hvsync_gen.vpos[9] ),
    .Y(_0169_));
 sg13g2_or2_1 _0693_ (.X(_0170_),
    .B(_0169_),
    .A(_0168_));
 sg13g2_a21o_1 _0694_ (.A2(_0166_),
    .A1(_0164_),
    .B1(_0170_),
    .X(_0171_));
 sg13g2_o21ai_1 _0695_ (.B1(\hvsync_gen.hpos[9] ),
    .Y(_0172_),
    .A1(\hvsync_gen.hpos[8] ),
    .A2(\hvsync_gen.hpos[7] ));
 sg13g2_nor2b_1 _0696_ (.A(\hvsync_gen.vpos[9] ),
    .B_N(_0172_),
    .Y(_0173_));
 sg13g2_o21ai_1 _0697_ (.B1(_0173_),
    .Y(_0174_),
    .A1(_0118_),
    .A2(_0128_));
 sg13g2_and2_1 _0698_ (.A(net177),
    .B(net285),
    .X(_0175_));
 sg13g2_and3_2 _0699_ (.X(_0176_),
    .A(net56),
    .B(net196),
    .C(_0175_));
 sg13g2_nor2_1 _0700_ (.A(net57),
    .B(_0118_),
    .Y(_0177_));
 sg13g2_a21oi_1 _0701_ (.A1(_0169_),
    .A2(_0177_),
    .Y(_0178_),
    .B1(\hvsync_gen.hpos[7] ));
 sg13g2_nand2_1 _0702_ (.Y(_0179_),
    .A(\hvsync_gen.hpos[8] ),
    .B(\hvsync_gen.hpos[6] ));
 sg13g2_nor4_1 _0703_ (.A(\hvsync_gen.hpos[9] ),
    .B(net55),
    .C(\hvsync_gen.hpos[4] ),
    .D(_0179_),
    .Y(_0180_));
 sg13g2_nand2_1 _0704_ (.Y(_0181_),
    .A(_0178_),
    .B(_0180_));
 sg13g2_or3_1 _0705_ (.A(_0174_),
    .B(_0176_),
    .C(_0181_),
    .X(_0182_));
 sg13g2_or3_1 _0706_ (.A(_0141_),
    .B(_0144_),
    .C(_0152_),
    .X(_0183_));
 sg13g2_nand2b_1 _0707_ (.Y(_0184_),
    .B(\hvsync_gen.vpos[5] ),
    .A_N(\dinosaur_y_pos[5] ));
 sg13g2_and2_1 _0708_ (.A(_0143_),
    .B(_0184_),
    .X(_0185_));
 sg13g2_nor2_1 _0709_ (.A(_0108_),
    .B(net52),
    .Y(_0186_));
 sg13g2_a221oi_1 _0710_ (.B2(_0185_),
    .C1(_0186_),
    .B1(_0183_),
    .A1(\dinosaur_y_pos[5] ),
    .Y(_0187_),
    .A2(_0120_));
 sg13g2_nand2_1 _0711_ (.Y(_0188_),
    .A(_0108_),
    .B(net52));
 sg13g2_o21ai_1 _0712_ (.B1(_0188_),
    .Y(_0189_),
    .A1(\dinosaur_y_pos[7] ),
    .A2(_0119_));
 sg13g2_a221oi_1 _0713_ (.B2(\dinosaur_y_pos[7] ),
    .C1(_0169_),
    .B1(_0119_),
    .A1(net57),
    .Y(_0190_),
    .A2(_0118_));
 sg13g2_o21ai_1 _0714_ (.B1(_0190_),
    .Y(_0191_),
    .A1(_0187_),
    .A2(_0189_));
 sg13g2_nor2_1 _0715_ (.A(_0167_),
    .B(_0177_),
    .Y(_0192_));
 sg13g2_a21oi_1 _0716_ (.A1(_0191_),
    .A2(_0192_),
    .Y(_0193_),
    .B1(_0182_));
 sg13g2_xor2_1 _0717_ (.B(_0150_),
    .A(_0146_),
    .X(_0194_));
 sg13g2_xnor2_1 _0718_ (.Y(_0195_),
    .A(_0146_),
    .B(_0150_));
 sg13g2_xor2_1 _0719_ (.B(_0149_),
    .A(_0148_),
    .X(_0196_));
 sg13g2_xnor2_1 _0720_ (.Y(_0197_),
    .A(_0148_),
    .B(_0149_));
 sg13g2_o21ai_1 _0721_ (.B1(\hvsync_gen.hpos[0] ),
    .Y(_0198_),
    .A1(_0194_),
    .A2(_0196_));
 sg13g2_xor2_1 _0722_ (.B(net54),
    .A(\dinosaur_y_pos[0] ),
    .X(_0199_));
 sg13g2_nand3_1 _0723_ (.B(_0196_),
    .C(_0199_),
    .A(_0194_),
    .Y(_0200_));
 sg13g2_nand2b_1 _0724_ (.Y(_0201_),
    .B(_0124_),
    .A_N(_0200_));
 sg13g2_xnor2_1 _0725_ (.Y(_0202_),
    .A(\dinosaur_y_pos[3] ),
    .B(\hvsync_gen.vpos[3] ));
 sg13g2_xnor2_1 _0726_ (.Y(_0203_),
    .A(_0151_),
    .B(_0202_));
 sg13g2_a21oi_1 _0727_ (.A1(_0198_),
    .A2(_0201_),
    .Y(_0204_),
    .B1(_0203_));
 sg13g2_and2_1 _0728_ (.A(_0196_),
    .B(_0199_),
    .X(_0205_));
 sg13g2_nand3b_1 _0729_ (.B(\hvsync_gen.hpos[0] ),
    .C(_0195_),
    .Y(_0206_),
    .A_N(_0205_));
 sg13g2_a21oi_1 _0730_ (.A1(_0124_),
    .A2(_0206_),
    .Y(_0207_),
    .B1(net56));
 sg13g2_nor3_1 _0731_ (.A(_0194_),
    .B(_0196_),
    .C(_0199_),
    .Y(_0208_));
 sg13g2_nor4_1 _0732_ (.A(_0122_),
    .B(_0194_),
    .C(_0196_),
    .D(_0199_),
    .Y(_0209_));
 sg13g2_o21ai_1 _0733_ (.B1(_0203_),
    .Y(_0210_),
    .A1(_0124_),
    .A2(_0209_));
 sg13g2_o21ai_1 _0734_ (.B1(_0210_),
    .Y(_0211_),
    .A1(\hvsync_gen.hpos[1] ),
    .A2(_0207_));
 sg13g2_o21ai_1 _0735_ (.B1(_0211_),
    .Y(_0212_),
    .A1(_0123_),
    .A2(_0204_));
 sg13g2_mux2_1 _0736_ (.A0(_0197_),
    .A1(_0205_),
    .S(_0195_),
    .X(_0213_));
 sg13g2_o21ai_1 _0737_ (.B1(_0203_),
    .Y(_0214_),
    .A1(\hvsync_gen.hpos[0] ),
    .A2(_0213_));
 sg13g2_nor2_2 _0738_ (.A(net177),
    .B(net285),
    .Y(_0215_));
 sg13g2_a21oi_1 _0739_ (.A1(_0195_),
    .A2(_0197_),
    .Y(_0216_),
    .B1(\hvsync_gen.hpos[1] ));
 sg13g2_a21oi_1 _0740_ (.A1(_0200_),
    .A2(_0216_),
    .Y(_0217_),
    .B1(_0215_));
 sg13g2_and2_1 _0741_ (.A(net56),
    .B(_0203_),
    .X(_0218_));
 sg13g2_a221oi_1 _0742_ (.B2(_0208_),
    .C1(_0217_),
    .B1(_0218_),
    .A1(_0123_),
    .Y(_0219_),
    .A2(_0214_));
 sg13g2_nand3b_1 _0743_ (.B(_0203_),
    .C(_0213_),
    .Y(_0220_),
    .A_N(\hvsync_gen.hpos[0] ));
 sg13g2_a21oi_1 _0744_ (.A1(\hvsync_gen.hpos[3] ),
    .A2(_0220_),
    .Y(_0221_),
    .B1(_0122_));
 sg13g2_or3_1 _0745_ (.A(_0124_),
    .B(_0219_),
    .C(_0221_),
    .X(_0222_));
 sg13g2_and4_1 _0746_ (.A(_0171_),
    .B(_0193_),
    .C(_0212_),
    .D(_0222_),
    .X(uo_out[6]));
 sg13g2_nor2b_1 _0747_ (.A(\square_x_pos[9] ),
    .B_N(\hvsync_gen.hpos[9] ),
    .Y(_0223_));
 sg13g2_a21oi_1 _0748_ (.A1(_0094_),
    .A2(\hvsync_gen.hpos[8] ),
    .Y(_0224_),
    .B1(_0223_));
 sg13g2_o21ai_1 _0749_ (.B1(_0224_),
    .Y(_0225_),
    .A1(\square_x_pos[7] ),
    .A2(_0125_));
 sg13g2_nand2b_1 _0750_ (.Y(_0226_),
    .B(\square_x_pos[0] ),
    .A_N(\hvsync_gen.hpos[0] ));
 sg13g2_nor2_1 _0751_ (.A(\square_x_pos[2] ),
    .B(_0124_),
    .Y(_0227_));
 sg13g2_nand2_1 _0752_ (.Y(_0228_),
    .A(\hvsync_gen.hpos[1] ),
    .B(_0226_));
 sg13g2_a22oi_1 _0753_ (.Y(_0229_),
    .B1(_0228_),
    .B2(\square_x_pos[1] ),
    .A2(_0215_),
    .A1(\square_x_pos[0] ));
 sg13g2_a22oi_1 _0754_ (.Y(_0230_),
    .B1(_0124_),
    .B2(\square_x_pos[2] ),
    .A2(_0123_),
    .A1(\square_x_pos[3] ));
 sg13g2_o21ai_1 _0755_ (.B1(_0230_),
    .Y(_0231_),
    .A1(_0227_),
    .A2(_0229_));
 sg13g2_a22oi_1 _0756_ (.Y(_0232_),
    .B1(\hvsync_gen.hpos[4] ),
    .B2(_0098_),
    .A2(net56),
    .A1(_0099_));
 sg13g2_a22oi_1 _0757_ (.Y(_0233_),
    .B1(_0231_),
    .B2(_0232_),
    .A2(_0127_),
    .A1(\square_x_pos[4] ));
 sg13g2_o21ai_1 _0758_ (.B1(_0233_),
    .Y(_0234_),
    .A1(_0097_),
    .A2(net55));
 sg13g2_a22oi_1 _0759_ (.Y(_0235_),
    .B1(net55),
    .B2(_0097_),
    .A2(\hvsync_gen.hpos[6] ),
    .A1(_0096_));
 sg13g2_nor2_1 _0760_ (.A(_0095_),
    .B(\hvsync_gen.hpos[7] ),
    .Y(_0236_));
 sg13g2_a221oi_1 _0761_ (.B2(_0235_),
    .C1(_0236_),
    .B1(_0234_),
    .A1(\square_x_pos[6] ),
    .Y(_0237_),
    .A2(_0126_));
 sg13g2_or2_1 _0762_ (.X(_0238_),
    .B(_0237_),
    .A(_0225_));
 sg13g2_a21o_2 _0763_ (.A2(\square_x_pos[1] ),
    .A1(\square_x_pos[2] ),
    .B1(\square_x_pos[3] ),
    .X(_0239_));
 sg13g2_nand3_1 _0764_ (.B(\square_x_pos[4] ),
    .C(_0239_),
    .A(\square_x_pos[5] ),
    .Y(_0240_));
 sg13g2_or2_1 _0765_ (.X(_0241_),
    .B(_0240_),
    .A(_0096_));
 sg13g2_a21oi_1 _0766_ (.A1(\hvsync_gen.hpos[1] ),
    .A2(_0226_),
    .Y(_0242_),
    .B1(\square_x_pos[1] ));
 sg13g2_xor2_1 _0767_ (.B(\square_x_pos[1] ),
    .A(\square_x_pos[2] ),
    .X(_0243_));
 sg13g2_a22oi_1 _0768_ (.Y(_0244_),
    .B1(_0243_),
    .B2(_0124_),
    .A2(_0215_),
    .A1(\square_x_pos[0] ));
 sg13g2_nand2b_1 _0769_ (.Y(_0245_),
    .B(_0244_),
    .A_N(_0242_));
 sg13g2_nand3_1 _0770_ (.B(\square_x_pos[2] ),
    .C(\square_x_pos[1] ),
    .A(\square_x_pos[3] ),
    .Y(_0246_));
 sg13g2_and2_1 _0771_ (.A(_0239_),
    .B(_0246_),
    .X(_0247_));
 sg13g2_nor2_1 _0772_ (.A(_0124_),
    .B(_0243_),
    .Y(_0248_));
 sg13g2_a21oi_1 _0773_ (.A1(net56),
    .A2(_0247_),
    .Y(_0249_),
    .B1(_0248_));
 sg13g2_xnor2_1 _0774_ (.Y(_0250_),
    .A(_0098_),
    .B(_0239_));
 sg13g2_nor2_1 _0775_ (.A(net56),
    .B(_0247_),
    .Y(_0251_));
 sg13g2_a221oi_1 _0776_ (.B2(_0127_),
    .C1(_0251_),
    .B1(_0250_),
    .A1(_0245_),
    .Y(_0252_),
    .A2(_0249_));
 sg13g2_nor2_1 _0777_ (.A(_0127_),
    .B(_0250_),
    .Y(_0253_));
 sg13g2_a21o_1 _0778_ (.A2(_0239_),
    .A1(\square_x_pos[4] ),
    .B1(\square_x_pos[5] ),
    .X(_0254_));
 sg13g2_nand2_1 _0779_ (.Y(_0255_),
    .A(_0240_),
    .B(_0254_));
 sg13g2_a21oi_1 _0780_ (.A1(net55),
    .A2(_0255_),
    .Y(_0256_),
    .B1(_0253_));
 sg13g2_nor2b_1 _0781_ (.A(_0252_),
    .B_N(_0256_),
    .Y(_0257_));
 sg13g2_xnor2_1 _0782_ (.Y(_0258_),
    .A(_0096_),
    .B(_0240_));
 sg13g2_nand2b_1 _0783_ (.Y(_0259_),
    .B(_0126_),
    .A_N(_0258_));
 sg13g2_o21ai_1 _0784_ (.B1(_0259_),
    .Y(_0260_),
    .A1(net55),
    .A2(_0255_));
 sg13g2_nand2b_1 _0785_ (.Y(_0261_),
    .B(\square_x_pos[8] ),
    .A_N(\hvsync_gen.hpos[8] ));
 sg13g2_o21ai_1 _0786_ (.B1(_0261_),
    .Y(_0262_),
    .A1(\square_x_pos[8] ),
    .A2(_0223_));
 sg13g2_a21oi_1 _0787_ (.A1(_0236_),
    .A2(_0262_),
    .Y(_0263_),
    .B1(_0224_));
 sg13g2_a21oi_1 _0788_ (.A1(\hvsync_gen.hpos[6] ),
    .A2(_0258_),
    .Y(_0264_),
    .B1(_0263_));
 sg13g2_o21ai_1 _0789_ (.B1(_0264_),
    .Y(_0265_),
    .A1(_0257_),
    .A2(_0260_));
 sg13g2_o21ai_1 _0790_ (.B1(_0265_),
    .Y(_0266_),
    .A1(_0225_),
    .A2(_0241_));
 sg13g2_and2_1 _0791_ (.A(_0225_),
    .B(_0241_),
    .X(_0267_));
 sg13g2_nor4_1 _0792_ (.A(\hvsync_gen.vpos[8] ),
    .B(_0121_),
    .C(_0128_),
    .D(_0130_),
    .Y(_0268_));
 sg13g2_nor4_1 _0793_ (.A(\hvsync_gen.vpos[7] ),
    .B(net52),
    .C(\hvsync_gen.vpos[5] ),
    .D(\hvsync_gen.vpos[4] ),
    .Y(_0269_));
 sg13g2_nor3_1 _0794_ (.A(_0118_),
    .B(\hvsync_gen.vpos[3] ),
    .C(\hvsync_gen.vpos[2] ),
    .Y(_0270_));
 sg13g2_a21oi_1 _0795_ (.A1(_0269_),
    .A2(_0270_),
    .Y(_0271_),
    .B1(_0268_));
 sg13g2_nand2b_1 _0796_ (.Y(_0272_),
    .B(\square_x_pos[9] ),
    .A_N(\hvsync_gen.hpos[9] ));
 sg13g2_o21ai_1 _0797_ (.B1(_0272_),
    .Y(_0273_),
    .A1(_0223_),
    .A2(_0261_));
 sg13g2_nor4_1 _0798_ (.A(_0174_),
    .B(_0267_),
    .C(_0271_),
    .D(_0273_),
    .Y(_0274_));
 sg13g2_and2_1 _0799_ (.A(_0266_),
    .B(_0274_),
    .X(_0275_));
 sg13g2_a21o_1 _0800_ (.A2(_0275_),
    .A1(_0238_),
    .B1(uo_out[6]),
    .X(uo_out[4]));
 sg13g2_nor4_1 _0801_ (.A(net135),
    .B(net141),
    .C(net139),
    .D(net137),
    .Y(_0276_));
 sg13g2_nor3_1 _0802_ (.A(\jump_counter[8] ),
    .B(\jump_counter[7] ),
    .C(\jump_counter[6] ),
    .Y(_0277_));
 sg13g2_nor4_1 _0803_ (.A(\jump_counter[13] ),
    .B(\jump_counter[12] ),
    .C(\jump_counter[11] ),
    .D(\jump_counter[10] ),
    .Y(_0278_));
 sg13g2_o21ai_1 _0804_ (.B1(_0278_),
    .Y(_0279_),
    .A1(_0105_),
    .A2(_0277_));
 sg13g2_a21oi_1 _0805_ (.A1(\jump_counter[14] ),
    .A2(_0279_),
    .Y(_0280_),
    .B1(\jump_counter[15] ));
 sg13g2_nand4_1 _0806_ (.B(\jump_counter[18] ),
    .C(\jump_counter[17] ),
    .A(\jump_counter[19] ),
    .Y(_0281_),
    .D(\jump_counter[16] ));
 sg13g2_o21ai_1 _0807_ (.B1(_0276_),
    .Y(_0282_),
    .A1(_0280_),
    .A2(_0281_));
 sg13g2_inv_1 _0808_ (.Y(_0283_),
    .A(_0282_));
 sg13g2_nor3_2 _0809_ (.A(net290),
    .B(net190),
    .C(net189),
    .Y(_0284_));
 sg13g2_nand2_1 _0810_ (.Y(_0285_),
    .A(net225),
    .B(_0284_));
 sg13g2_and2_1 _0811_ (.A(\dinosaur_y_pos[1] ),
    .B(\dinosaur_y_pos[0] ),
    .X(_0286_));
 sg13g2_nor4_1 _0812_ (.A(\dinosaur_y_pos[5] ),
    .B(\dinosaur_y_pos[3] ),
    .C(\dinosaur_y_pos[2] ),
    .D(_0286_),
    .Y(_0287_));
 sg13g2_nor4_1 _0813_ (.A(_0107_),
    .B(_0108_),
    .C(_0139_),
    .D(_0287_),
    .Y(_0288_));
 sg13g2_nor3_1 _0814_ (.A(net261),
    .B(net57),
    .C(_0288_),
    .Y(_0289_));
 sg13g2_nand2b_1 _0815_ (.Y(_0290_),
    .B(_0289_),
    .A_N(_0285_));
 sg13g2_nor3_2 _0816_ (.A(\jump_state[0] ),
    .B(\jump_state[3] ),
    .C(\jump_state[2] ),
    .Y(_0291_));
 sg13g2_nand2_1 _0817_ (.Y(_0292_),
    .A(\jump_state[1] ),
    .B(_0291_));
 sg13g2_nor4_1 _0818_ (.A(net261),
    .B(net57),
    .C(_0157_),
    .D(net50),
    .Y(_0293_));
 sg13g2_a21oi_1 _0819_ (.A1(\jump_state[0] ),
    .A2(_0284_),
    .Y(_0294_),
    .B1(_0293_));
 sg13g2_inv_1 _0820_ (.Y(_0295_),
    .A(_0294_));
 sg13g2_and3_2 _0821_ (.X(_0296_),
    .A(_0282_),
    .B(_0290_),
    .C(_0295_));
 sg13g2_nand3_1 _0822_ (.B(_0290_),
    .C(_0295_),
    .A(_0282_),
    .Y(_0297_));
 sg13g2_xnor2_1 _0823_ (.Y(_0298_),
    .A(net287),
    .B(_0296_));
 sg13g2_nor2_1 _0824_ (.A(net58),
    .B(_0298_),
    .Y(_0002_));
 sg13g2_a21oi_1 _0825_ (.A1(\jump_state[1] ),
    .A2(_0291_),
    .Y(_0299_),
    .B1(_0111_));
 sg13g2_nand3_1 _0826_ (.B(\jump_state[1] ),
    .C(_0291_),
    .A(_0111_),
    .Y(_0300_));
 sg13g2_nor2b_1 _0827_ (.A(_0299_),
    .B_N(_0300_),
    .Y(_0301_));
 sg13g2_xor2_1 _0828_ (.B(_0301_),
    .A(\dinosaur_y_pos[0] ),
    .X(_0302_));
 sg13g2_o21ai_1 _0829_ (.B1(net59),
    .Y(_0303_),
    .A1(net49),
    .A2(_0302_));
 sg13g2_a21oi_1 _0830_ (.A1(_0111_),
    .A2(net49),
    .Y(_0003_),
    .B1(_0303_));
 sg13g2_and2_1 _0831_ (.A(net288),
    .B(net50),
    .X(_0304_));
 sg13g2_xor2_1 _0832_ (.B(net50),
    .A(net288),
    .X(_0305_));
 sg13g2_a21o_1 _0833_ (.A2(_0300_),
    .A1(net287),
    .B1(_0299_),
    .X(_0306_));
 sg13g2_xnor2_1 _0834_ (.Y(_0307_),
    .A(_0305_),
    .B(_0306_));
 sg13g2_o21ai_1 _0835_ (.B1(net59),
    .Y(_0308_),
    .A1(net288),
    .A2(_0296_));
 sg13g2_a21oi_1 _0836_ (.A1(_0296_),
    .A2(_0307_),
    .Y(_0004_),
    .B1(_0308_));
 sg13g2_nor2_1 _0837_ (.A(\dinosaur_y_pos[3] ),
    .B(net51),
    .Y(_0309_));
 sg13g2_xnor2_1 _0838_ (.Y(_0310_),
    .A(net299),
    .B(net50));
 sg13g2_a21oi_1 _0839_ (.A1(_0305_),
    .A2(_0306_),
    .Y(_0311_),
    .B1(_0304_));
 sg13g2_xnor2_1 _0840_ (.Y(_0312_),
    .A(_0310_),
    .B(_0311_));
 sg13g2_o21ai_1 _0841_ (.B1(net59),
    .Y(_0313_),
    .A1(net299),
    .A2(_0296_));
 sg13g2_a21oi_1 _0842_ (.A1(_0296_),
    .A2(_0312_),
    .Y(_0005_),
    .B1(_0313_));
 sg13g2_xnor2_1 _0843_ (.Y(_0314_),
    .A(\dinosaur_y_pos[4] ),
    .B(net51));
 sg13g2_a221oi_1 _0844_ (.B2(_0306_),
    .C1(_0304_),
    .B1(_0305_),
    .A1(\dinosaur_y_pos[3] ),
    .Y(_0315_),
    .A2(net51));
 sg13g2_o21ai_1 _0845_ (.B1(_0314_),
    .Y(_0316_),
    .A1(_0309_),
    .A2(_0315_));
 sg13g2_nor3_1 _0846_ (.A(_0309_),
    .B(_0314_),
    .C(_0315_),
    .Y(_0317_));
 sg13g2_nor2_1 _0847_ (.A(net49),
    .B(_0317_),
    .Y(_0318_));
 sg13g2_a22oi_1 _0848_ (.Y(_0319_),
    .B1(_0316_),
    .B2(_0318_),
    .A2(net49),
    .A1(net304));
 sg13g2_nand2_1 _0849_ (.Y(_0006_),
    .A(net61),
    .B(_0319_));
 sg13g2_a21oi_1 _0850_ (.A1(\dinosaur_y_pos[4] ),
    .A2(net51),
    .Y(_0320_),
    .B1(_0317_));
 sg13g2_xnor2_1 _0851_ (.Y(_0321_),
    .A(net292),
    .B(net51));
 sg13g2_xnor2_1 _0852_ (.Y(_0322_),
    .A(_0320_),
    .B(_0321_));
 sg13g2_a21oi_1 _0853_ (.A1(net292),
    .A2(net49),
    .Y(_0323_),
    .B1(net58));
 sg13g2_o21ai_1 _0854_ (.B1(_0323_),
    .Y(_0007_),
    .A1(net49),
    .A2(_0322_));
 sg13g2_a21oi_1 _0855_ (.A1(\jump_state[1] ),
    .A2(_0291_),
    .Y(_0324_),
    .B1(_0108_));
 sg13g2_xnor2_1 _0856_ (.Y(_0325_),
    .A(_0108_),
    .B(net50));
 sg13g2_inv_1 _0857_ (.Y(_0326_),
    .A(_0325_));
 sg13g2_or4_1 _0858_ (.A(_0309_),
    .B(_0314_),
    .C(_0315_),
    .D(_0321_),
    .X(_0327_));
 sg13g2_nand2b_1 _0859_ (.Y(_0328_),
    .B(net50),
    .A_N(_0139_));
 sg13g2_nand3_1 _0860_ (.B(_0327_),
    .C(_0328_),
    .A(_0326_),
    .Y(_0329_));
 sg13g2_a21o_1 _0861_ (.A2(_0328_),
    .A1(_0327_),
    .B1(_0326_),
    .X(_0330_));
 sg13g2_nand3_1 _0862_ (.B(_0329_),
    .C(_0330_),
    .A(_0296_),
    .Y(_0331_));
 sg13g2_a21oi_1 _0863_ (.A1(net278),
    .A2(net49),
    .Y(_0332_),
    .B1(net58));
 sg13g2_nand2_1 _0864_ (.Y(_0008_),
    .A(_0331_),
    .B(_0332_));
 sg13g2_xnor2_1 _0865_ (.Y(_0333_),
    .A(_0107_),
    .B(net50));
 sg13g2_nand2b_1 _0866_ (.Y(_0334_),
    .B(_0330_),
    .A_N(_0324_));
 sg13g2_xnor2_1 _0867_ (.Y(_0335_),
    .A(_0333_),
    .B(_0334_));
 sg13g2_a21oi_1 _0868_ (.A1(net282),
    .A2(net49),
    .Y(_0336_),
    .B1(net58));
 sg13g2_o21ai_1 _0869_ (.B1(_0336_),
    .Y(_0009_),
    .A1(_0297_),
    .A2(_0335_));
 sg13g2_nand2_1 _0870_ (.Y(_0337_),
    .A(_0325_),
    .B(_0333_));
 sg13g2_nand2b_1 _0871_ (.Y(_0338_),
    .B(_0328_),
    .A_N(_0324_));
 sg13g2_a21oi_1 _0872_ (.A1(\dinosaur_y_pos[7] ),
    .A2(net51),
    .Y(_0339_),
    .B1(_0338_));
 sg13g2_o21ai_1 _0873_ (.B1(_0339_),
    .Y(_0340_),
    .A1(_0327_),
    .A2(_0337_));
 sg13g2_xor2_1 _0874_ (.B(_0340_),
    .A(net50),
    .X(_0341_));
 sg13g2_a21oi_1 _0875_ (.A1(_0296_),
    .A2(_0341_),
    .Y(_0342_),
    .B1(net57));
 sg13g2_and3_1 _0876_ (.X(_0343_),
    .A(net57),
    .B(_0296_),
    .C(_0341_));
 sg13g2_nor3_1 _0877_ (.A(net58),
    .B(_0342_),
    .C(_0343_),
    .Y(_0010_));
 sg13g2_nor3_1 _0878_ (.A(\dinosaur_y_pos[8] ),
    .B(_0297_),
    .C(_0340_),
    .Y(_0344_));
 sg13g2_nor3_1 _0879_ (.A(_0106_),
    .B(_0117_),
    .C(_0344_),
    .Y(_0011_));
 sg13g2_and2_1 _0880_ (.A(net280),
    .B(_0176_),
    .X(_0345_));
 sg13g2_nor3_1 _0881_ (.A(\hvsync_gen.hpos[7] ),
    .B(\hvsync_gen.hpos[6] ),
    .C(net55),
    .Y(_0346_));
 sg13g2_nand4_1 _0882_ (.B(\hvsync_gen.hpos[8] ),
    .C(_0345_),
    .A(\hvsync_gen.hpos[9] ),
    .Y(_0347_),
    .D(_0346_));
 sg13g2_inv_1 _0883_ (.Y(_0348_),
    .A(_0347_));
 sg13g2_nor2_2 _0884_ (.A(net58),
    .B(_0348_),
    .Y(_0349_));
 sg13g2_nand2_2 _0885_ (.Y(_0350_),
    .A(net62),
    .B(_0347_));
 sg13g2_nor2_1 _0886_ (.A(net177),
    .B(_0350_),
    .Y(_0012_));
 sg13g2_nor3_1 _0887_ (.A(_0175_),
    .B(_0215_),
    .C(_0350_),
    .Y(_0013_));
 sg13g2_o21ai_1 _0888_ (.B1(net62),
    .Y(_0351_),
    .A1(net196),
    .A2(_0175_));
 sg13g2_a21oi_1 _0889_ (.A1(net196),
    .A2(_0175_),
    .Y(_0014_),
    .B1(_0351_));
 sg13g2_a21oi_1 _0890_ (.A1(net196),
    .A2(_0175_),
    .Y(_0352_),
    .B1(net56));
 sg13g2_nor3_1 _0891_ (.A(net58),
    .B(_0176_),
    .C(net272),
    .Y(_0015_));
 sg13g2_o21ai_1 _0892_ (.B1(net62),
    .Y(_0353_),
    .A1(net280),
    .A2(_0176_));
 sg13g2_nor2_1 _0893_ (.A(_0345_),
    .B(_0353_),
    .Y(_0016_));
 sg13g2_and2_1 _0894_ (.A(net241),
    .B(_0345_),
    .X(_0354_));
 sg13g2_nor2_1 _0895_ (.A(net241),
    .B(_0345_),
    .Y(_0355_));
 sg13g2_nor3_1 _0896_ (.A(_0350_),
    .B(_0354_),
    .C(net242),
    .Y(_0017_));
 sg13g2_xnor2_1 _0897_ (.Y(_0356_),
    .A(net286),
    .B(_0354_));
 sg13g2_nor2_1 _0898_ (.A(_0350_),
    .B(_0356_),
    .Y(_0018_));
 sg13g2_and3_1 _0899_ (.X(_0357_),
    .A(net256),
    .B(_0132_),
    .C(_0176_));
 sg13g2_a21oi_1 _0900_ (.A1(_0132_),
    .A2(_0176_),
    .Y(_0358_),
    .B1(net256));
 sg13g2_nor3_1 _0901_ (.A(_0350_),
    .B(_0357_),
    .C(net257),
    .Y(_0019_));
 sg13g2_nor2_1 _0902_ (.A(net198),
    .B(_0357_),
    .Y(_0359_));
 sg13g2_and2_1 _0903_ (.A(net198),
    .B(_0357_),
    .X(_0360_));
 sg13g2_nor3_1 _0904_ (.A(_0350_),
    .B(_0359_),
    .C(_0360_),
    .Y(_0020_));
 sg13g2_a21oi_1 _0905_ (.A1(net289),
    .A2(_0360_),
    .Y(_0361_),
    .B1(_0350_));
 sg13g2_o21ai_1 _0906_ (.B1(_0361_),
    .Y(_0362_),
    .A1(net289),
    .A2(_0360_));
 sg13g2_inv_1 _0907_ (.Y(_0021_),
    .A(_0362_));
 sg13g2_nor2b_2 _0908_ (.A(\jump_state[0] ),
    .B_N(_0284_),
    .Y(_0363_));
 sg13g2_or4_1 _0909_ (.A(net225),
    .B(net305),
    .C(net190),
    .D(net189),
    .X(_0364_));
 sg13g2_o21ai_1 _0910_ (.B1(net60),
    .Y(_0365_),
    .A1(_0283_),
    .A2(_0363_));
 sg13g2_inv_4 _0911_ (.A(net48),
    .Y(_0366_));
 sg13g2_nor2_1 _0912_ (.A(net230),
    .B(_0364_),
    .Y(_0367_));
 sg13g2_and2_1 _0913_ (.A(net230),
    .B(_0364_),
    .X(_0368_));
 sg13g2_nor3_1 _0914_ (.A(net47),
    .B(net231),
    .C(_0368_),
    .Y(_0022_));
 sg13g2_o21ai_1 _0915_ (.B1(_0366_),
    .Y(_0369_),
    .A1(net158),
    .A2(_0368_));
 sg13g2_a21oi_1 _0916_ (.A1(net158),
    .A2(_0368_),
    .Y(_0023_),
    .B1(_0369_));
 sg13g2_and4_1 _0917_ (.A(net149),
    .B(net158),
    .C(\jump_counter[0] ),
    .D(_0364_),
    .X(_0370_));
 sg13g2_a21oi_1 _0918_ (.A1(\jump_counter[1] ),
    .A2(_0368_),
    .Y(_0371_),
    .B1(net149));
 sg13g2_nor3_1 _0919_ (.A(net48),
    .B(_0370_),
    .C(net150),
    .Y(_0024_));
 sg13g2_and2_1 _0920_ (.A(net202),
    .B(_0370_),
    .X(_0372_));
 sg13g2_nor2_1 _0921_ (.A(net202),
    .B(_0370_),
    .Y(_0373_));
 sg13g2_nor3_1 _0922_ (.A(net47),
    .B(_0372_),
    .C(net203),
    .Y(_0025_));
 sg13g2_o21ai_1 _0923_ (.B1(_0366_),
    .Y(_0374_),
    .A1(net160),
    .A2(_0372_));
 sg13g2_a21oi_1 _0924_ (.A1(net160),
    .A2(_0372_),
    .Y(_0026_),
    .B1(_0374_));
 sg13g2_and2_1 _0925_ (.A(net143),
    .B(net160),
    .X(_0375_));
 sg13g2_and2_1 _0926_ (.A(_0372_),
    .B(_0375_),
    .X(_0376_));
 sg13g2_a21oi_1 _0927_ (.A1(\jump_counter[4] ),
    .A2(_0372_),
    .Y(_0377_),
    .B1(net143));
 sg13g2_nor3_1 _0928_ (.A(net48),
    .B(_0376_),
    .C(net144),
    .Y(_0027_));
 sg13g2_nor2_1 _0929_ (.A(net213),
    .B(_0376_),
    .Y(_0378_));
 sg13g2_and4_1 _0930_ (.A(net213),
    .B(net202),
    .C(_0370_),
    .D(_0375_),
    .X(_0379_));
 sg13g2_nor3_1 _0931_ (.A(net48),
    .B(_0378_),
    .C(_0379_),
    .Y(_0028_));
 sg13g2_and2_1 _0932_ (.A(net236),
    .B(_0379_),
    .X(_0380_));
 sg13g2_nor2_1 _0933_ (.A(net236),
    .B(_0379_),
    .Y(_0381_));
 sg13g2_nor3_1 _0934_ (.A(net48),
    .B(_0380_),
    .C(_0381_),
    .Y(_0029_));
 sg13g2_o21ai_1 _0935_ (.B1(_0366_),
    .Y(_0382_),
    .A1(net152),
    .A2(_0380_));
 sg13g2_a21oi_1 _0936_ (.A1(net152),
    .A2(_0380_),
    .Y(_0030_),
    .B1(_0382_));
 sg13g2_a21oi_1 _0937_ (.A1(net152),
    .A2(_0380_),
    .Y(_0383_),
    .B1(net168));
 sg13g2_nand4_1 _0938_ (.B(net152),
    .C(net236),
    .A(net168),
    .Y(_0384_),
    .D(_0379_));
 sg13g2_nand2_1 _0939_ (.Y(_0385_),
    .A(_0366_),
    .B(_0384_));
 sg13g2_nor2_1 _0940_ (.A(net169),
    .B(_0385_),
    .Y(_0031_));
 sg13g2_and2_1 _0941_ (.A(_0104_),
    .B(_0384_),
    .X(_0386_));
 sg13g2_nor2_1 _0942_ (.A(_0104_),
    .B(_0384_),
    .Y(_0387_));
 sg13g2_nor3_1 _0943_ (.A(net47),
    .B(_0386_),
    .C(_0387_),
    .Y(_0032_));
 sg13g2_nor2_1 _0944_ (.A(net214),
    .B(_0387_),
    .Y(_0388_));
 sg13g2_nor3_2 _0945_ (.A(_0103_),
    .B(_0104_),
    .C(_0384_),
    .Y(_0389_));
 sg13g2_nor3_1 _0946_ (.A(net47),
    .B(net215),
    .C(_0389_),
    .Y(_0033_));
 sg13g2_o21ai_1 _0947_ (.B1(_0366_),
    .Y(_0390_),
    .A1(net154),
    .A2(_0389_));
 sg13g2_a21oi_1 _0948_ (.A1(net154),
    .A2(_0389_),
    .Y(_0034_),
    .B1(_0390_));
 sg13g2_a21oi_1 _0949_ (.A1(net154),
    .A2(_0389_),
    .Y(_0391_),
    .B1(net181));
 sg13g2_nand2_1 _0950_ (.Y(_0392_),
    .A(net181),
    .B(net154));
 sg13g2_nor4_1 _0951_ (.A(_0103_),
    .B(_0104_),
    .C(_0384_),
    .D(_0392_),
    .Y(_0393_));
 sg13g2_nor3_1 _0952_ (.A(net47),
    .B(net182),
    .C(_0393_),
    .Y(_0035_));
 sg13g2_nor2_1 _0953_ (.A(net239),
    .B(_0393_),
    .Y(_0394_));
 sg13g2_and2_1 _0954_ (.A(net239),
    .B(_0393_),
    .X(_0395_));
 sg13g2_nor3_1 _0955_ (.A(net47),
    .B(net240),
    .C(_0395_),
    .Y(_0036_));
 sg13g2_nor2_1 _0956_ (.A(net219),
    .B(_0395_),
    .Y(_0396_));
 sg13g2_and3_2 _0957_ (.X(_0397_),
    .A(net219),
    .B(net239),
    .C(_0393_));
 sg13g2_nor3_1 _0958_ (.A(net47),
    .B(net220),
    .C(_0397_),
    .Y(_0037_));
 sg13g2_nand2_1 _0959_ (.Y(_0398_),
    .A(\jump_counter[16] ),
    .B(_0397_));
 sg13g2_a21oi_1 _0960_ (.A1(net284),
    .A2(_0397_),
    .Y(_0399_),
    .B1(net47));
 sg13g2_o21ai_1 _0961_ (.B1(_0399_),
    .Y(_0400_),
    .A1(net284),
    .A2(_0397_));
 sg13g2_inv_1 _0962_ (.Y(_0038_),
    .A(_0400_));
 sg13g2_nand3_1 _0963_ (.B(\jump_counter[16] ),
    .C(_0397_),
    .A(net200),
    .Y(_0401_));
 sg13g2_nand2_1 _0964_ (.Y(_0402_),
    .A(_0366_),
    .B(_0401_));
 sg13g2_a21oi_1 _0965_ (.A1(_0102_),
    .A2(_0398_),
    .Y(_0039_),
    .B1(_0402_));
 sg13g2_or2_1 _0966_ (.X(_0403_),
    .B(_0401_),
    .A(_0282_));
 sg13g2_nand4_1 _0967_ (.B(\jump_counter[17] ),
    .C(\jump_counter[16] ),
    .A(net187),
    .Y(_0404_),
    .D(_0397_));
 sg13g2_nand2_1 _0968_ (.Y(_0405_),
    .A(_0366_),
    .B(_0404_));
 sg13g2_a21oi_1 _0969_ (.A1(_0101_),
    .A2(_0403_),
    .Y(_0040_),
    .B1(_0405_));
 sg13g2_nand3_1 _0970_ (.B(_0366_),
    .C(_0404_),
    .A(net191),
    .Y(_0406_));
 sg13g2_nand3b_1 _0971_ (.B(net59),
    .C(_0276_),
    .Y(_0407_),
    .A_N(net191));
 sg13g2_o21ai_1 _0972_ (.B1(net192),
    .Y(_0041_),
    .A1(_0404_),
    .A2(_0407_));
 sg13g2_and3_1 _0973_ (.X(_0042_),
    .A(net137),
    .B(net59),
    .C(_0363_));
 sg13g2_and3_1 _0974_ (.X(_0043_),
    .A(net139),
    .B(net59),
    .C(_0363_));
 sg13g2_and3_1 _0975_ (.X(_0044_),
    .A(net141),
    .B(net59),
    .C(_0363_));
 sg13g2_and3_1 _0976_ (.X(_0045_),
    .A(net135),
    .B(net59),
    .C(_0363_));
 sg13g2_nor2_1 _0977_ (.A(\square_counter[7] ),
    .B(\square_counter[8] ),
    .Y(_0408_));
 sg13g2_nand2_1 _0978_ (.Y(_0409_),
    .A(net146),
    .B(\square_counter[9] ));
 sg13g2_o21ai_1 _0979_ (.B1(_0113_),
    .Y(_0410_),
    .A1(_0408_),
    .A2(_0409_));
 sg13g2_or2_1 _0980_ (.X(_0411_),
    .B(\square_counter[13] ),
    .A(\square_counter[14] ));
 sg13g2_a21oi_1 _0981_ (.A1(\square_counter[12] ),
    .A2(_0410_),
    .Y(_0412_),
    .B1(_0411_));
 sg13g2_nor3_1 _0982_ (.A(\square_counter[18] ),
    .B(\square_counter[17] ),
    .C(\square_counter[16] ),
    .Y(_0413_));
 sg13g2_o21ai_1 _0983_ (.B1(_0413_),
    .Y(_0414_),
    .A1(_0112_),
    .A2(_0412_));
 sg13g2_and2_1 _0984_ (.A(\square_counter[20] ),
    .B(\square_counter[19] ),
    .X(_0415_));
 sg13g2_or2_1 _0985_ (.X(_0416_),
    .B(\square_counter[21] ),
    .A(\square_counter[22] ));
 sg13g2_a21oi_1 _0986_ (.A1(_0414_),
    .A2(_0415_),
    .Y(_0417_),
    .B1(_0416_));
 sg13g2_or2_1 _0987_ (.X(_0418_),
    .B(\square_x_pos[2] ),
    .A(\square_x_pos[3] ));
 sg13g2_nand2b_1 _0988_ (.Y(_0419_),
    .B(_0098_),
    .A_N(_0418_));
 sg13g2_or4_1 _0989_ (.A(net234),
    .B(\square_x_pos[6] ),
    .C(\square_x_pos[5] ),
    .D(_0419_),
    .X(_0420_));
 sg13g2_nand2b_1 _0990_ (.Y(_0421_),
    .B(_0094_),
    .A_N(_0420_));
 sg13g2_nor3_1 _0991_ (.A(net259),
    .B(\square_x_pos[1] ),
    .C(_0421_),
    .Y(_0422_));
 sg13g2_or4_1 _0992_ (.A(net297),
    .B(_0116_),
    .C(_0417_),
    .D(_0422_),
    .X(_0423_));
 sg13g2_o21ai_1 _0993_ (.B1(net62),
    .Y(_0424_),
    .A1(_0116_),
    .A2(_0417_));
 sg13g2_or2_1 _0994_ (.X(_0425_),
    .B(net46),
    .A(_0100_));
 sg13g2_o21ai_1 _0995_ (.B1(_0425_),
    .Y(_0046_),
    .A1(net58),
    .A2(_0423_));
 sg13g2_nor2_1 _0996_ (.A(net253),
    .B(\square_x_pos[0] ),
    .Y(_0426_));
 sg13g2_nand3b_1 _0997_ (.B(_0426_),
    .C(net156),
    .Y(_0427_),
    .A_N(_0417_));
 sg13g2_nand2b_1 _0998_ (.Y(_0428_),
    .B(net62),
    .A_N(_0422_));
 sg13g2_nand3_1 _0999_ (.B(net62),
    .C(_0423_),
    .A(net253),
    .Y(_0429_));
 sg13g2_o21ai_1 _1000_ (.B1(net254),
    .Y(_0047_),
    .A1(_0427_),
    .A2(_0428_));
 sg13g2_and2_1 _1001_ (.A(net46),
    .B(_0428_),
    .X(_0430_));
 sg13g2_nor2_1 _1002_ (.A(\square_x_pos[2] ),
    .B(_0427_),
    .Y(_0431_));
 sg13g2_xor2_1 _1003_ (.B(_0427_),
    .A(net295),
    .X(_0432_));
 sg13g2_nor2_1 _1004_ (.A(_0430_),
    .B(net296),
    .Y(_0048_));
 sg13g2_xnor2_1 _1005_ (.Y(_0433_),
    .A(net269),
    .B(_0431_));
 sg13g2_nor2_1 _1006_ (.A(_0430_),
    .B(net270),
    .Y(_0049_));
 sg13g2_nor2_1 _1007_ (.A(_0419_),
    .B(_0427_),
    .Y(_0434_));
 sg13g2_o21ai_1 _1008_ (.B1(net303),
    .Y(_0435_),
    .A1(_0418_),
    .A2(_0427_));
 sg13g2_nor2b_1 _1009_ (.A(_0434_),
    .B_N(_0435_),
    .Y(_0436_));
 sg13g2_nor2_1 _1010_ (.A(_0430_),
    .B(_0436_),
    .Y(_0050_));
 sg13g2_nor3_1 _1011_ (.A(\square_x_pos[5] ),
    .B(_0419_),
    .C(_0427_),
    .Y(_0437_));
 sg13g2_xnor2_1 _1012_ (.Y(_0438_),
    .A(net273),
    .B(_0434_));
 sg13g2_nor2_1 _1013_ (.A(_0430_),
    .B(net274),
    .Y(_0051_));
 sg13g2_and2_1 _1014_ (.A(_0096_),
    .B(_0437_),
    .X(_0439_));
 sg13g2_xnor2_1 _1015_ (.Y(_0440_),
    .A(net265),
    .B(_0437_));
 sg13g2_nor2_1 _1016_ (.A(_0430_),
    .B(net266),
    .Y(_0052_));
 sg13g2_nor2b_1 _1017_ (.A(_0420_),
    .B_N(_0426_),
    .Y(_0441_));
 sg13g2_o21ai_1 _1018_ (.B1(net46),
    .Y(_0442_),
    .A1(_0428_),
    .A2(_0441_));
 sg13g2_o21ai_1 _1019_ (.B1(_0442_),
    .Y(_0053_),
    .A1(_0095_),
    .A2(_0439_));
 sg13g2_nand2_1 _1020_ (.Y(_0443_),
    .A(net194),
    .B(_0442_));
 sg13g2_or2_1 _1021_ (.X(_0444_),
    .B(_0427_),
    .A(_0421_));
 sg13g2_nand2_1 _1022_ (.Y(_0445_),
    .A(\square_x_pos[9] ),
    .B(net62));
 sg13g2_o21ai_1 _1023_ (.B1(_0443_),
    .Y(_0054_),
    .A1(_0444_),
    .A2(_0445_));
 sg13g2_a21o_1 _1024_ (.A2(_0444_),
    .A1(net259),
    .B1(_0430_),
    .X(_0055_));
 sg13g2_nor2b_1 _1025_ (.A(prev_button_state),
    .B_N(net1),
    .Y(_0446_));
 sg13g2_a21oi_1 _1026_ (.A1(_0284_),
    .A2(_0446_),
    .Y(_0447_),
    .B1(net225));
 sg13g2_o21ai_1 _1027_ (.B1(net60),
    .Y(_0448_),
    .A1(_0283_),
    .A2(_0290_));
 sg13g2_nor2_1 _1028_ (.A(net226),
    .B(_0448_),
    .Y(_0056_));
 sg13g2_a21oi_1 _1029_ (.A1(_0285_),
    .A2(net51),
    .Y(_0449_),
    .B1(_0283_));
 sg13g2_nor2_1 _1030_ (.A(_0289_),
    .B(_0293_),
    .Y(_0450_));
 sg13g2_o21ai_1 _1031_ (.B1(net60),
    .Y(_0451_),
    .A1(net290),
    .A2(_0449_));
 sg13g2_a21oi_1 _1032_ (.A1(_0449_),
    .A2(_0450_),
    .Y(_0057_),
    .B1(_0451_));
 sg13g2_and2_1 _1033_ (.A(net60),
    .B(net189),
    .X(_0058_));
 sg13g2_and2_1 _1034_ (.A(net60),
    .B(net190),
    .X(_0059_));
 sg13g2_nand2_1 _1035_ (.Y(_0452_),
    .A(net54),
    .B(_0349_));
 sg13g2_nor3_1 _1036_ (.A(net54),
    .B(\hvsync_gen.vpos[8] ),
    .C(net53),
    .Y(_0453_));
 sg13g2_nand4_1 _1037_ (.B(_0129_),
    .C(_0269_),
    .A(\hvsync_gen.vpos[9] ),
    .Y(_0454_),
    .D(_0453_));
 sg13g2_nand3_1 _1038_ (.B(_0348_),
    .C(_0454_),
    .A(net61),
    .Y(_0455_));
 sg13g2_o21ai_1 _1039_ (.B1(_0452_),
    .Y(_0060_),
    .A1(net54),
    .A2(net42));
 sg13g2_nand2_1 _1040_ (.Y(_0456_),
    .A(net53),
    .B(_0349_));
 sg13g2_xnor2_1 _1041_ (.Y(_0457_),
    .A(net54),
    .B(net53));
 sg13g2_o21ai_1 _1042_ (.B1(_0456_),
    .Y(_0061_),
    .A1(net42),
    .A2(_0457_));
 sg13g2_nand2_1 _1043_ (.Y(_0458_),
    .A(net245),
    .B(_0349_));
 sg13g2_a21oi_1 _1044_ (.A1(net54),
    .A2(net53),
    .Y(_0459_),
    .B1(net245));
 sg13g2_nand3_1 _1045_ (.B(net245),
    .C(net53),
    .A(net54),
    .Y(_0460_));
 sg13g2_nand2b_1 _1046_ (.Y(_0461_),
    .B(_0460_),
    .A_N(_0459_));
 sg13g2_o21ai_1 _1047_ (.B1(_0458_),
    .Y(_0062_),
    .A1(net42),
    .A2(_0461_));
 sg13g2_nand2_1 _1048_ (.Y(_0462_),
    .A(net267),
    .B(_0349_));
 sg13g2_nand3_1 _1049_ (.B(\hvsync_gen.vpos[1] ),
    .C(_0129_),
    .A(\hvsync_gen.vpos[0] ),
    .Y(_0463_));
 sg13g2_xor2_1 _1050_ (.B(_0460_),
    .A(net267),
    .X(_0464_));
 sg13g2_o21ai_1 _1051_ (.B1(_0462_),
    .Y(_0063_),
    .A1(net42),
    .A2(_0464_));
 sg13g2_nand2_1 _1052_ (.Y(_0465_),
    .A(net232),
    .B(_0349_));
 sg13g2_or2_1 _1053_ (.X(_0466_),
    .B(_0463_),
    .A(_0121_));
 sg13g2_xnor2_1 _1054_ (.Y(_0467_),
    .A(_0121_),
    .B(_0463_));
 sg13g2_o21ai_1 _1055_ (.B1(_0465_),
    .Y(_0064_),
    .A1(net42),
    .A2(_0467_));
 sg13g2_nand2_1 _1056_ (.Y(_0468_),
    .A(net211),
    .B(_0349_));
 sg13g2_nor2_1 _1057_ (.A(_0120_),
    .B(_0466_),
    .Y(_0469_));
 sg13g2_xnor2_1 _1058_ (.Y(_0470_),
    .A(_0120_),
    .B(_0466_));
 sg13g2_o21ai_1 _1059_ (.B1(_0468_),
    .Y(_0065_),
    .A1(_0455_),
    .A2(_0470_));
 sg13g2_nand2_1 _1060_ (.Y(_0471_),
    .A(net52),
    .B(_0349_));
 sg13g2_xnor2_1 _1061_ (.Y(_0472_),
    .A(net52),
    .B(_0469_));
 sg13g2_o21ai_1 _1062_ (.B1(_0471_),
    .Y(_0066_),
    .A1(net42),
    .A2(_0472_));
 sg13g2_nor2_1 _1063_ (.A(_0128_),
    .B(_0466_),
    .Y(_0473_));
 sg13g2_a21oi_1 _1064_ (.A1(\hvsync_gen.vpos[6] ),
    .A2(_0469_),
    .Y(_0474_),
    .B1(net263));
 sg13g2_or3_1 _1065_ (.A(_0455_),
    .B(_0473_),
    .C(_0474_),
    .X(_0475_));
 sg13g2_o21ai_1 _1066_ (.B1(_0475_),
    .Y(_0067_),
    .A1(_0119_),
    .A2(_0350_));
 sg13g2_a21oi_1 _1067_ (.A1(net279),
    .A2(_0473_),
    .Y(_0476_),
    .B1(net42));
 sg13g2_nor2_1 _1068_ (.A(_0349_),
    .B(_0476_),
    .Y(_0477_));
 sg13g2_nor2b_1 _1069_ (.A(net42),
    .B_N(_0473_),
    .Y(_0478_));
 sg13g2_nor2_1 _1070_ (.A(net279),
    .B(_0478_),
    .Y(_0479_));
 sg13g2_nor2_1 _1071_ (.A(_0477_),
    .B(_0479_),
    .Y(_0068_));
 sg13g2_a21oi_1 _1072_ (.A1(\hvsync_gen.vpos[8] ),
    .A2(_0478_),
    .Y(_0480_),
    .B1(net209));
 sg13g2_a21oi_1 _1073_ (.A1(net209),
    .A2(_0477_),
    .Y(_0069_),
    .B1(_0480_));
 sg13g2_nor2_1 _1074_ (.A(net134),
    .B(net44),
    .Y(_0070_));
 sg13g2_xnor2_1 _1075_ (.Y(_0481_),
    .A(net134),
    .B(net258));
 sg13g2_nor2_1 _1076_ (.A(net44),
    .B(_0481_),
    .Y(_0071_));
 sg13g2_and3_1 _1077_ (.X(_0482_),
    .A(net134),
    .B(\square_counter[1] ),
    .C(net162));
 sg13g2_a21oi_1 _1078_ (.A1(net134),
    .A2(\square_counter[1] ),
    .Y(_0483_),
    .B1(net162));
 sg13g2_nor3_1 _1079_ (.A(net44),
    .B(_0482_),
    .C(net163),
    .Y(_0072_));
 sg13g2_and4_1 _1080_ (.A(net134),
    .B(\square_counter[1] ),
    .C(net162),
    .D(net184),
    .X(_0484_));
 sg13g2_nor2_1 _1081_ (.A(net184),
    .B(_0482_),
    .Y(_0485_));
 sg13g2_nor3_1 _1082_ (.A(net44),
    .B(_0484_),
    .C(net185),
    .Y(_0073_));
 sg13g2_and2_1 _1083_ (.A(net207),
    .B(_0484_),
    .X(_0486_));
 sg13g2_nor2_1 _1084_ (.A(net207),
    .B(_0484_),
    .Y(_0487_));
 sg13g2_nor3_1 _1085_ (.A(net45),
    .B(_0486_),
    .C(net208),
    .Y(_0074_));
 sg13g2_xnor2_1 _1086_ (.Y(_0488_),
    .A(net247),
    .B(_0486_));
 sg13g2_nor2_1 _1087_ (.A(_0424_),
    .B(_0488_),
    .Y(_0075_));
 sg13g2_nand4_1 _1088_ (.B(net247),
    .C(net277),
    .A(net207),
    .Y(_0489_),
    .D(_0484_));
 sg13g2_a21oi_1 _1089_ (.A1(net247),
    .A2(_0486_),
    .Y(_0490_),
    .B1(net277));
 sg13g2_nor2_1 _1090_ (.A(net45),
    .B(_0490_),
    .Y(_0491_));
 sg13g2_and2_1 _1091_ (.A(_0489_),
    .B(_0491_),
    .X(_0076_));
 sg13g2_nor2_1 _1092_ (.A(_0114_),
    .B(_0489_),
    .Y(_0492_));
 sg13g2_and2_1 _1093_ (.A(_0114_),
    .B(_0489_),
    .X(_0493_));
 sg13g2_nor3_1 _1094_ (.A(net44),
    .B(_0492_),
    .C(_0493_),
    .Y(_0077_));
 sg13g2_nor3_1 _1095_ (.A(_0114_),
    .B(_0115_),
    .C(_0489_),
    .Y(_0494_));
 sg13g2_nor2_1 _1096_ (.A(net204),
    .B(_0492_),
    .Y(_0495_));
 sg13g2_nor3_1 _1097_ (.A(net44),
    .B(_0494_),
    .C(net205),
    .Y(_0078_));
 sg13g2_xnor2_1 _1098_ (.Y(_0496_),
    .A(net237),
    .B(_0494_));
 sg13g2_nor2_1 _1099_ (.A(net44),
    .B(net238),
    .Y(_0079_));
 sg13g2_nor4_1 _1100_ (.A(_0114_),
    .B(_0115_),
    .C(_0409_),
    .D(_0489_),
    .Y(_0497_));
 sg13g2_a21oi_1 _1101_ (.A1(\square_counter[9] ),
    .A2(_0494_),
    .Y(_0498_),
    .B1(net146));
 sg13g2_nor3_1 _1102_ (.A(net44),
    .B(_0497_),
    .C(net147),
    .Y(_0080_));
 sg13g2_and2_1 _1103_ (.A(net217),
    .B(_0497_),
    .X(_0499_));
 sg13g2_nor2_1 _1104_ (.A(net217),
    .B(_0497_),
    .Y(_0500_));
 sg13g2_nor3_1 _1105_ (.A(net43),
    .B(_0499_),
    .C(net218),
    .Y(_0081_));
 sg13g2_xnor2_1 _1106_ (.Y(_0501_),
    .A(net251),
    .B(_0499_));
 sg13g2_nor2_1 _1107_ (.A(net43),
    .B(_0501_),
    .Y(_0082_));
 sg13g2_a21oi_1 _1108_ (.A1(\square_counter[12] ),
    .A2(_0499_),
    .Y(_0502_),
    .B1(net178));
 sg13g2_and4_1 _1109_ (.A(net178),
    .B(\square_counter[12] ),
    .C(net217),
    .D(_0497_),
    .X(_0503_));
 sg13g2_nor3_1 _1110_ (.A(net43),
    .B(net179),
    .C(_0503_),
    .Y(_0083_));
 sg13g2_nor2_1 _1111_ (.A(net228),
    .B(_0503_),
    .Y(_0504_));
 sg13g2_and2_1 _1112_ (.A(net228),
    .B(_0503_),
    .X(_0505_));
 sg13g2_nor3_1 _1113_ (.A(net43),
    .B(net229),
    .C(_0505_),
    .Y(_0084_));
 sg13g2_xnor2_1 _1114_ (.Y(_0506_),
    .A(net252),
    .B(_0505_));
 sg13g2_nor2_1 _1115_ (.A(net43),
    .B(_0506_),
    .Y(_0085_));
 sg13g2_a21oi_1 _1116_ (.A1(\square_counter[15] ),
    .A2(_0505_),
    .Y(_0507_),
    .B1(net165));
 sg13g2_and4_1 _1117_ (.A(net165),
    .B(\square_counter[15] ),
    .C(net228),
    .D(_0503_),
    .X(_0508_));
 sg13g2_nor3_1 _1118_ (.A(net43),
    .B(net166),
    .C(_0508_),
    .Y(_0086_));
 sg13g2_nor2_1 _1119_ (.A(net249),
    .B(_0508_),
    .Y(_0509_));
 sg13g2_and2_1 _1120_ (.A(net249),
    .B(_0508_),
    .X(_0510_));
 sg13g2_nor3_1 _1121_ (.A(net43),
    .B(net250),
    .C(_0510_),
    .Y(_0087_));
 sg13g2_xnor2_1 _1122_ (.Y(_0511_),
    .A(net260),
    .B(_0510_));
 sg13g2_nor2_1 _1123_ (.A(net45),
    .B(_0511_),
    .Y(_0088_));
 sg13g2_a21oi_1 _1124_ (.A1(\square_counter[18] ),
    .A2(_0510_),
    .Y(_0512_),
    .B1(net171));
 sg13g2_and4_1 _1125_ (.A(net171),
    .B(\square_counter[18] ),
    .C(\square_counter[17] ),
    .D(_0508_),
    .X(_0513_));
 sg13g2_nor3_1 _1126_ (.A(net43),
    .B(net172),
    .C(_0513_),
    .Y(_0089_));
 sg13g2_xnor2_1 _1127_ (.Y(_0514_),
    .A(net243),
    .B(_0513_));
 sg13g2_nor2_1 _1128_ (.A(net46),
    .B(net244),
    .Y(_0090_));
 sg13g2_a21oi_1 _1129_ (.A1(\square_counter[20] ),
    .A2(_0513_),
    .Y(_0515_),
    .B1(net174));
 sg13g2_and3_2 _1130_ (.X(_0516_),
    .A(net174),
    .B(\square_counter[20] ),
    .C(_0513_));
 sg13g2_nor3_1 _1131_ (.A(net46),
    .B(net175),
    .C(_0516_),
    .Y(_0091_));
 sg13g2_nor2_1 _1132_ (.A(net222),
    .B(_0516_),
    .Y(_0517_));
 sg13g2_a21oi_1 _1133_ (.A1(net222),
    .A2(_0516_),
    .Y(_0518_),
    .B1(net46));
 sg13g2_nor2b_1 _1134_ (.A(net223),
    .B_N(_0518_),
    .Y(_0092_));
 sg13g2_a21oi_1 _1135_ (.A1(\square_counter[22] ),
    .A2(_0516_),
    .Y(_0519_),
    .B1(net156));
 sg13g2_nor2_1 _1136_ (.A(net46),
    .B(net157),
    .Y(_0093_));
 sg13g2_dfrbpq_2 _1137_ (.RESET_B(net97),
    .D(_0002_),
    .Q(\dinosaur_y_pos[0] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _1138_ (.RESET_B(net78),
    .D(net276),
    .Q(\dinosaur_y_pos[1] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _1139_ (.RESET_B(net76),
    .D(_0004_),
    .Q(\dinosaur_y_pos[2] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _1140_ (.RESET_B(net74),
    .D(_0005_),
    .Q(\dinosaur_y_pos[3] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _1141_ (.RESET_B(net72),
    .D(_0006_),
    .Q(\dinosaur_y_pos[4] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _1142_ (.RESET_B(net70),
    .D(net293),
    .Q(\dinosaur_y_pos[5] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _1143_ (.RESET_B(net68),
    .D(_0008_),
    .Q(\dinosaur_y_pos[6] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _1144_ (.RESET_B(net66),
    .D(net283),
    .Q(\dinosaur_y_pos[7] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_1 _1145_ (.RESET_B(net64),
    .D(_0010_),
    .Q(\dinosaur_y_pos[8] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _1146_ (.RESET_B(net41),
    .D(net262),
    .Q(\dinosaur_y_pos[9] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _1147_ (.RESET_B(net39),
    .D(_0012_),
    .Q(\hvsync_gen.hpos[0] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _1148_ (.RESET_B(net38),
    .D(_0013_),
    .Q(\hvsync_gen.hpos[1] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _1149_ (.RESET_B(net37),
    .D(net197),
    .Q(\hvsync_gen.hpos[2] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_1 _1150_ (.RESET_B(net36),
    .D(_0015_),
    .Q(\hvsync_gen.hpos[3] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _1151_ (.RESET_B(net35),
    .D(_0016_),
    .Q(\hvsync_gen.hpos[4] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _1152_ (.RESET_B(net34),
    .D(_0017_),
    .Q(\hvsync_gen.hpos[5] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_2 _1153_ (.RESET_B(net33),
    .D(_0018_),
    .Q(\hvsync_gen.hpos[6] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_2 _1154_ (.RESET_B(net32),
    .D(_0019_),
    .Q(\hvsync_gen.hpos[7] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _1155_ (.RESET_B(net31),
    .D(_0020_),
    .Q(\hvsync_gen.hpos[8] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_2 _1156_ (.RESET_B(net30),
    .D(_0021_),
    .Q(\hvsync_gen.hpos[9] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_1 _1157_ (.RESET_B(net29),
    .D(_0022_),
    .Q(\jump_counter[0] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_1 _1158_ (.RESET_B(net27),
    .D(net159),
    .Q(\jump_counter[1] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _1159_ (.RESET_B(net25),
    .D(net151),
    .Q(\jump_counter[2] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_1 _1160_ (.RESET_B(net23),
    .D(_0025_),
    .Q(\jump_counter[3] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _1161_ (.RESET_B(net21),
    .D(net161),
    .Q(\jump_counter[4] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _1162_ (.RESET_B(net19),
    .D(net145),
    .Q(\jump_counter[5] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _1163_ (.RESET_B(net133),
    .D(_0028_),
    .Q(\jump_counter[6] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _1164_ (.RESET_B(net131),
    .D(_0029_),
    .Q(\jump_counter[7] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_2 _1165_ (.RESET_B(net129),
    .D(net153),
    .Q(\jump_counter[8] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _1166_ (.RESET_B(net127),
    .D(net170),
    .Q(\jump_counter[9] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _1167_ (.RESET_B(net125),
    .D(_0032_),
    .Q(\jump_counter[10] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _1168_ (.RESET_B(net123),
    .D(net216),
    .Q(\jump_counter[11] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _1169_ (.RESET_B(net121),
    .D(net155),
    .Q(\jump_counter[12] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _1170_ (.RESET_B(net119),
    .D(net183),
    .Q(\jump_counter[13] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _1171_ (.RESET_B(net117),
    .D(_0036_),
    .Q(\jump_counter[14] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _1172_ (.RESET_B(net115),
    .D(net221),
    .Q(\jump_counter[15] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _1173_ (.RESET_B(net113),
    .D(_0038_),
    .Q(\jump_counter[16] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_1 _1174_ (.RESET_B(net111),
    .D(net201),
    .Q(\jump_counter[17] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _1175_ (.RESET_B(net108),
    .D(net188),
    .Q(\jump_counter[18] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _1176_ (.RESET_B(net106),
    .D(net193),
    .Q(\jump_counter[19] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_1 _1177_ (.RESET_B(net104),
    .D(net138),
    .Q(\jump_counter[20] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_1 _1178_ (.RESET_B(net102),
    .D(net140),
    .Q(\jump_counter[21] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_1 _1179_ (.RESET_B(net100),
    .D(net142),
    .Q(\jump_counter[22] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_1 _1180_ (.RESET_B(net96),
    .D(net136),
    .Q(\jump_counter[23] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _1181_ (.RESET_B(net94),
    .D(_0046_),
    .Q(\square_x_pos[0] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _1182_ (.RESET_B(net92),
    .D(net255),
    .Q(\square_x_pos[1] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_2 _1183_ (.RESET_B(net90),
    .D(_0048_),
    .Q(\square_x_pos[2] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_2 _1184_ (.RESET_B(net88),
    .D(_0049_),
    .Q(\square_x_pos[3] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_2 _1185_ (.RESET_B(net86),
    .D(_0050_),
    .Q(\square_x_pos[4] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_2 _1186_ (.RESET_B(net84),
    .D(_0051_),
    .Q(\square_x_pos[5] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_2 _1187_ (.RESET_B(net82),
    .D(_0052_),
    .Q(\square_x_pos[6] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_1 _1188_ (.RESET_B(net80),
    .D(net235),
    .Q(\square_x_pos[7] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_1 _1189_ (.RESET_B(net77),
    .D(net195),
    .Q(\square_x_pos[8] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_2 _1190_ (.RESET_B(net73),
    .D(_0055_),
    .Q(\square_x_pos[9] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_2 _1191_ (.RESET_B(net69),
    .D(net227),
    .Q(\jump_state[0] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _1192_ (.RESET_B(net67),
    .D(net291),
    .Q(\jump_state[1] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _1193_ (.RESET_B(net65),
    .D(_0058_),
    .Q(\jump_state[2] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _1194_ (.RESET_B(net98),
    .D(_0059_),
    .Q(\jump_state[3] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_1 _1195_ (.RESET_B(net109),
    .D(net1),
    .Q(prev_button_state),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_1 _1196_ (.RESET_B(net63),
    .D(net199),
    .Q(hsync),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_1 _1197_ (.RESET_B(net40),
    .D(_0060_),
    .Q(\hvsync_gen.vpos[0] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_1 _1198_ (.RESET_B(net26),
    .D(_0061_),
    .Q(\hvsync_gen.vpos[1] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_2 _1199_ (.RESET_B(net22),
    .D(net246),
    .Q(\hvsync_gen.vpos[2] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _1200_ (.RESET_B(net18),
    .D(net268),
    .Q(\hvsync_gen.vpos[3] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _1201_ (.RESET_B(net130),
    .D(net233),
    .Q(\hvsync_gen.vpos[4] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _1202_ (.RESET_B(net126),
    .D(net212),
    .Q(\hvsync_gen.vpos[5] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_1 _1203_ (.RESET_B(net122),
    .D(_0066_),
    .Q(\hvsync_gen.vpos[6] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _1204_ (.RESET_B(net118),
    .D(net264),
    .Q(\hvsync_gen.vpos[7] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_2 _1205_ (.RESET_B(net114),
    .D(_0068_),
    .Q(\hvsync_gen.vpos[8] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_2 _1206_ (.RESET_B(net107),
    .D(net210),
    .Q(\hvsync_gen.vpos[9] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_1 _1207_ (.RESET_B(net110),
    .D(_0001_),
    .Q(\hvsync_gen.vsync ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_2 _1208_ (.RESET_B(net105),
    .D(_0070_),
    .Q(\square_counter[0] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _1209_ (.RESET_B(net103),
    .D(_0071_),
    .Q(\square_counter[1] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_1 _1210_ (.RESET_B(net101),
    .D(net164),
    .Q(\square_counter[2] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_1 _1211_ (.RESET_B(net99),
    .D(net186),
    .Q(\square_counter[3] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_1 _1212_ (.RESET_B(net95),
    .D(_0074_),
    .Q(\square_counter[4] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_1 _1213_ (.RESET_B(net93),
    .D(net248),
    .Q(\square_counter[5] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_1 _1214_ (.RESET_B(net91),
    .D(_0076_),
    .Q(\square_counter[6] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_1 _1215_ (.RESET_B(net89),
    .D(_0077_),
    .Q(\square_counter[7] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_1 _1216_ (.RESET_B(net87),
    .D(net206),
    .Q(\square_counter[8] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _1217_ (.RESET_B(net85),
    .D(_0079_),
    .Q(\square_counter[9] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _1218_ (.RESET_B(net83),
    .D(net148),
    .Q(\square_counter[10] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _1219_ (.RESET_B(net81),
    .D(_0081_),
    .Q(\square_counter[11] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_2 _1220_ (.RESET_B(net79),
    .D(_0082_),
    .Q(\square_counter[12] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _1221_ (.RESET_B(net75),
    .D(net180),
    .Q(\square_counter[13] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _1222_ (.RESET_B(net71),
    .D(_0084_),
    .Q(\square_counter[14] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_2 _1223_ (.RESET_B(net28),
    .D(_0085_),
    .Q(\square_counter[15] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _1224_ (.RESET_B(net24),
    .D(net167),
    .Q(\square_counter[16] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _1225_ (.RESET_B(net20),
    .D(_0087_),
    .Q(\square_counter[17] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_2 _1226_ (.RESET_B(net132),
    .D(_0088_),
    .Q(\square_counter[18] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_1 _1227_ (.RESET_B(net128),
    .D(net173),
    .Q(\square_counter[19] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_2 _1228_ (.RESET_B(net124),
    .D(_0090_),
    .Q(\square_counter[20] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_1 _1229_ (.RESET_B(net120),
    .D(net176),
    .Q(\square_counter[21] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_1 _1230_ (.RESET_B(net116),
    .D(net224),
    .Q(\square_counter[22] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_1 _1231_ (.RESET_B(net112),
    .D(_0093_),
    .Q(\square_counter[23] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_tiehi _1162__19 (.L_HI(net19));
 sg13g2_tiehi _1225__20 (.L_HI(net20));
 sg13g2_tiehi _1161__21 (.L_HI(net21));
 sg13g2_tiehi _1199__22 (.L_HI(net22));
 sg13g2_tiehi _1160__23 (.L_HI(net23));
 sg13g2_tiehi _1224__24 (.L_HI(net24));
 sg13g2_tiehi _1159__25 (.L_HI(net25));
 sg13g2_tiehi _1198__26 (.L_HI(net26));
 sg13g2_tiehi _1158__27 (.L_HI(net27));
 sg13g2_tiehi _1223__28 (.L_HI(net28));
 sg13g2_tiehi _1157__29 (.L_HI(net29));
 sg13g2_tiehi _1156__30 (.L_HI(net30));
 sg13g2_tiehi _1155__31 (.L_HI(net31));
 sg13g2_tiehi _1154__32 (.L_HI(net32));
 sg13g2_tiehi _1153__33 (.L_HI(net33));
 sg13g2_tiehi _1152__34 (.L_HI(net34));
 sg13g2_tiehi _1151__35 (.L_HI(net35));
 sg13g2_tiehi _1150__36 (.L_HI(net36));
 sg13g2_tiehi _1149__37 (.L_HI(net37));
 sg13g2_tiehi _1148__38 (.L_HI(net38));
 sg13g2_tiehi _1147__39 (.L_HI(net39));
 sg13g2_tiehi _1197__40 (.L_HI(net40));
 sg13g2_tiehi _1146__41 (.L_HI(net41));
 sg13g2_tiehi _1196__42 (.L_HI(net63));
 sg13g2_tiehi _1145__43 (.L_HI(net64));
 sg13g2_tiehi _1193__44 (.L_HI(net65));
 sg13g2_tiehi _1144__45 (.L_HI(net66));
 sg13g2_tiehi _1192__46 (.L_HI(net67));
 sg13g2_tiehi _1143__47 (.L_HI(net68));
 sg13g2_tiehi _1191__48 (.L_HI(net69));
 sg13g2_tiehi _1142__49 (.L_HI(net70));
 sg13g2_tiehi _1222__50 (.L_HI(net71));
 sg13g2_tiehi _1141__51 (.L_HI(net72));
 sg13g2_tiehi _1190__52 (.L_HI(net73));
 sg13g2_tiehi _1140__53 (.L_HI(net74));
 sg13g2_tiehi _1221__54 (.L_HI(net75));
 sg13g2_tiehi _1139__55 (.L_HI(net76));
 sg13g2_tiehi _1189__56 (.L_HI(net77));
 sg13g2_tiehi _1138__57 (.L_HI(net78));
 sg13g2_tiehi _1220__58 (.L_HI(net79));
 sg13g2_tiehi _1188__59 (.L_HI(net80));
 sg13g2_tiehi _1219__60 (.L_HI(net81));
 sg13g2_tiehi _1187__61 (.L_HI(net82));
 sg13g2_tiehi _1218__62 (.L_HI(net83));
 sg13g2_tiehi _1186__63 (.L_HI(net84));
 sg13g2_tiehi _1217__64 (.L_HI(net85));
 sg13g2_tiehi _1185__65 (.L_HI(net86));
 sg13g2_tiehi _1216__66 (.L_HI(net87));
 sg13g2_tiehi _1184__67 (.L_HI(net88));
 sg13g2_tiehi _1215__68 (.L_HI(net89));
 sg13g2_tiehi _1183__69 (.L_HI(net90));
 sg13g2_tiehi _1214__70 (.L_HI(net91));
 sg13g2_tiehi _1182__71 (.L_HI(net92));
 sg13g2_tiehi _1213__72 (.L_HI(net93));
 sg13g2_tiehi _1181__73 (.L_HI(net94));
 sg13g2_tiehi _1212__74 (.L_HI(net95));
 sg13g2_tiehi _1180__75 (.L_HI(net96));
 sg13g2_tiehi _1137__76 (.L_HI(net97));
 sg13g2_tiehi _1194__77 (.L_HI(net98));
 sg13g2_tiehi _1211__78 (.L_HI(net99));
 sg13g2_tiehi _1179__79 (.L_HI(net100));
 sg13g2_tiehi _1210__80 (.L_HI(net101));
 sg13g2_tiehi _1178__81 (.L_HI(net102));
 sg13g2_tiehi _1209__82 (.L_HI(net103));
 sg13g2_tiehi _1177__83 (.L_HI(net104));
 sg13g2_tiehi _1208__84 (.L_HI(net105));
 sg13g2_tiehi _1176__85 (.L_HI(net106));
 sg13g2_tiehi _1206__86 (.L_HI(net107));
 sg13g2_tiehi _1175__87 (.L_HI(net108));
 sg13g2_tiehi _1195__88 (.L_HI(net109));
 sg13g2_tiehi _1207__89 (.L_HI(net110));
 sg13g2_tiehi _1174__90 (.L_HI(net111));
 sg13g2_tiehi _1231__91 (.L_HI(net112));
 sg13g2_tiehi _1173__92 (.L_HI(net113));
 sg13g2_tiehi _1205__93 (.L_HI(net114));
 sg13g2_tiehi _1172__94 (.L_HI(net115));
 sg13g2_tiehi _1230__95 (.L_HI(net116));
 sg13g2_tiehi _1171__96 (.L_HI(net117));
 sg13g2_tiehi _1204__97 (.L_HI(net118));
 sg13g2_tiehi _1170__98 (.L_HI(net119));
 sg13g2_tiehi _1229__99 (.L_HI(net120));
 sg13g2_tiehi _1169__100 (.L_HI(net121));
 sg13g2_tiehi _1203__101 (.L_HI(net122));
 sg13g2_tiehi _1168__102 (.L_HI(net123));
 sg13g2_tiehi _1228__103 (.L_HI(net124));
 sg13g2_tiehi _1167__104 (.L_HI(net125));
 sg13g2_tiehi _1202__105 (.L_HI(net126));
 sg13g2_tiehi _1166__106 (.L_HI(net127));
 sg13g2_tiehi _1227__107 (.L_HI(net128));
 sg13g2_tiehi _1165__108 (.L_HI(net129));
 sg13g2_tiehi _1201__109 (.L_HI(net130));
 sg13g2_tiehi _1164__110 (.L_HI(net131));
 sg13g2_tiehi _1226__111 (.L_HI(net132));
 sg13g2_tiehi _1163__112 (.L_HI(net133));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_not_a_dinosaur_3 (.L_LO(net3));
 sg13g2_tielo tt_um_not_a_dinosaur_4 (.L_LO(net4));
 sg13g2_tielo tt_um_not_a_dinosaur_5 (.L_LO(net5));
 sg13g2_tielo tt_um_not_a_dinosaur_6 (.L_LO(net6));
 sg13g2_tielo tt_um_not_a_dinosaur_7 (.L_LO(net7));
 sg13g2_tielo tt_um_not_a_dinosaur_8 (.L_LO(net8));
 sg13g2_tielo tt_um_not_a_dinosaur_9 (.L_LO(net9));
 sg13g2_tielo tt_um_not_a_dinosaur_10 (.L_LO(net10));
 sg13g2_tielo tt_um_not_a_dinosaur_11 (.L_LO(net11));
 sg13g2_tielo tt_um_not_a_dinosaur_12 (.L_LO(net12));
 sg13g2_tielo tt_um_not_a_dinosaur_13 (.L_LO(net13));
 sg13g2_tielo tt_um_not_a_dinosaur_14 (.L_LO(net14));
 sg13g2_tielo tt_um_not_a_dinosaur_15 (.L_LO(net15));
 sg13g2_tielo tt_um_not_a_dinosaur_16 (.L_LO(net16));
 sg13g2_tielo tt_um_not_a_dinosaur_17 (.L_LO(net17));
 sg13g2_tiehi _1200__18 (.L_HI(net18));
 sg13g2_buf_1 _1343_ (.A(uo_out[4]),
    .X(uo_out[0]));
 sg13g2_buf_1 _1344_ (.A(uo_out[6]),
    .X(uo_out[1]));
 sg13g2_buf_1 _1345_ (.A(uo_out[6]),
    .X(uo_out[2]));
 sg13g2_buf_1 _1346_ (.A(\hvsync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _1347_ (.A(uo_out[6]),
    .X(uo_out[5]));
 sg13g2_buf_1 _1348_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout42 (.A(_0455_),
    .X(net42));
 sg13g2_buf_8 fanout43 (.A(net45),
    .X(net43));
 sg13g2_buf_8 fanout44 (.A(net45),
    .X(net44));
 sg13g2_buf_8 fanout45 (.A(net46),
    .X(net45));
 sg13g2_buf_8 fanout46 (.A(_0424_),
    .X(net46));
 sg13g2_buf_8 fanout47 (.A(_0365_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0365_),
    .X(net48));
 sg13g2_buf_8 fanout49 (.A(_0297_),
    .X(net49));
 sg13g2_buf_8 fanout50 (.A(net51),
    .X(net50));
 sg13g2_buf_8 fanout51 (.A(_0292_),
    .X(net51));
 sg13g2_buf_8 fanout52 (.A(net281),
    .X(net52));
 sg13g2_buf_8 fanout53 (.A(net302),
    .X(net53));
 sg13g2_buf_8 fanout54 (.A(net294),
    .X(net54));
 sg13g2_buf_8 fanout55 (.A(net241),
    .X(net55));
 sg13g2_buf_8 fanout56 (.A(net271),
    .X(net56));
 sg13g2_buf_8 fanout57 (.A(net301),
    .X(net57));
 sg13g2_buf_8 fanout58 (.A(_0117_),
    .X(net58));
 sg13g2_buf_8 fanout59 (.A(net61),
    .X(net59));
 sg13g2_buf_1 fanout60 (.A(net61),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(rst_n),
    .X(net61));
 sg13g2_buf_8 fanout62 (.A(rst_n),
    .X(net62));
 sg13g2_buf_1 input1 (.A(ui_in[1]),
    .X(net1));
 sg13g2_tielo tt_um_not_a_dinosaur_2 (.L_LO(net2));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_4_0_0_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_4_1_0_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_4_2_0_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_4_3_0_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_4_4_0_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_4_5_0_clk));
 sg13g2_buf_1 clkload6 (.A(clknet_4_7_0_clk));
 sg13g2_buf_1 clkload7 (.A(clknet_4_8_0_clk));
 sg13g2_buf_1 clkload8 (.A(clknet_4_9_0_clk));
 sg13g2_buf_1 clkload9 (.A(clknet_4_10_0_clk));
 sg13g2_buf_1 clkload10 (.A(clknet_4_11_0_clk));
 sg13g2_buf_1 clkload11 (.A(clknet_4_12_0_clk));
 sg13g2_buf_1 clkload12 (.A(clknet_4_13_0_clk));
 sg13g2_buf_1 clkload13 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\square_counter[0] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold2 (.A(\jump_counter[23] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0045_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold4 (.A(\jump_counter[20] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0042_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold6 (.A(\jump_counter[21] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0043_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold8 (.A(\jump_counter[22] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0044_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold10 (.A(\jump_counter[5] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0377_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0027_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold13 (.A(\square_counter[10] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0498_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0080_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold16 (.A(\jump_counter[2] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0371_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0024_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold19 (.A(\jump_counter[8] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0030_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold21 (.A(\jump_counter[12] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0034_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold23 (.A(\square_counter[23] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0519_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold25 (.A(\jump_counter[1] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0023_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold27 (.A(\jump_counter[4] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0026_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold29 (.A(\square_counter[2] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0483_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0072_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold32 (.A(\square_counter[16] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0507_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0086_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold35 (.A(\jump_counter[9] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0383_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0031_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold38 (.A(\square_counter[19] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0512_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0089_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold41 (.A(\square_counter[21] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0515_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0091_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold44 (.A(\hvsync_gen.hpos[0] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold45 (.A(\square_counter[13] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0502_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0083_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold48 (.A(\jump_counter[13] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0391_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0035_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold51 (.A(\square_counter[3] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0485_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0073_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold54 (.A(\jump_counter[18] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0040_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold56 (.A(\jump_state[2] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold57 (.A(\jump_state[3] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold58 (.A(\jump_counter[19] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0406_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0041_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold61 (.A(\square_x_pos[8] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0054_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold63 (.A(\hvsync_gen.hpos[2] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0014_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold65 (.A(\hvsync_gen.hpos[8] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0000_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold67 (.A(\jump_counter[17] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0039_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold69 (.A(\jump_counter[3] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0373_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold71 (.A(\square_counter[8] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0495_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0078_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold74 (.A(\square_counter[4] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0487_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold76 (.A(\hvsync_gen.vpos[9] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0069_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold78 (.A(\hvsync_gen.vpos[5] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0065_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold80 (.A(\jump_counter[6] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold81 (.A(\jump_counter[11] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0388_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0033_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold84 (.A(\square_counter[11] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0500_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold86 (.A(\jump_counter[15] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0396_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0037_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold89 (.A(\square_counter[22] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0517_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0092_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold92 (.A(\jump_state[0] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0447_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0056_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold95 (.A(\square_counter[14] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0504_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold97 (.A(\jump_counter[0] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0367_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold99 (.A(\hvsync_gen.vpos[4] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0064_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold101 (.A(\square_x_pos[7] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0053_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold103 (.A(\jump_counter[7] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold104 (.A(\square_counter[9] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0496_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold106 (.A(\jump_counter[14] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0394_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold108 (.A(\hvsync_gen.hpos[5] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0355_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold110 (.A(\square_counter[20] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0514_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold112 (.A(\hvsync_gen.vpos[2] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0062_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold114 (.A(\square_counter[5] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0075_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold116 (.A(\square_counter[17] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0509_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold118 (.A(\square_counter[12] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold119 (.A(\square_counter[15] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold120 (.A(\square_x_pos[1] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0429_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0047_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold123 (.A(\hvsync_gen.hpos[7] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0358_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold125 (.A(\square_counter[1] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold126 (.A(\square_x_pos[9] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold127 (.A(\square_counter[18] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold128 (.A(\dinosaur_y_pos[9] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0011_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold130 (.A(\hvsync_gen.vpos[7] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0067_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold132 (.A(\square_x_pos[6] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0440_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold134 (.A(\hvsync_gen.vpos[3] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0063_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold136 (.A(\square_x_pos[3] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0433_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold138 (.A(\hvsync_gen.hpos[3] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0352_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold140 (.A(\square_x_pos[5] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0438_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold142 (.A(\dinosaur_y_pos[1] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0003_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold144 (.A(\square_counter[6] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold145 (.A(\dinosaur_y_pos[6] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold146 (.A(\hvsync_gen.vpos[8] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold147 (.A(\hvsync_gen.hpos[4] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold148 (.A(\hvsync_gen.vpos[6] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold149 (.A(\dinosaur_y_pos[7] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0009_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold151 (.A(\jump_counter[16] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold152 (.A(\hvsync_gen.hpos[1] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold153 (.A(\hvsync_gen.hpos[6] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold154 (.A(\dinosaur_y_pos[0] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold155 (.A(\dinosaur_y_pos[2] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold156 (.A(\hvsync_gen.hpos[9] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold157 (.A(\jump_state[1] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0057_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold159 (.A(\dinosaur_y_pos[5] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0007_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold161 (.A(\hvsync_gen.vpos[0] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold162 (.A(\square_x_pos[2] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0432_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold164 (.A(\square_x_pos[0] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold165 (.A(\jump_counter[10] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold166 (.A(\dinosaur_y_pos[3] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold167 (.A(\square_counter[7] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold168 (.A(\dinosaur_y_pos[8] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold169 (.A(\hvsync_gen.vpos[1] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold170 (.A(\square_x_pos[4] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold171 (.A(\dinosaur_y_pos[4] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold172 (.A(\jump_state[1] ),
    .X(net305));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_fill_2 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_4 FILLER_6_308 ();
 sg13g2_fill_2 FILLER_6_312 ();
 sg13g2_decap_8 FILLER_6_319 ();
 sg13g2_decap_8 FILLER_6_326 ();
 sg13g2_decap_8 FILLER_6_333 ();
 sg13g2_decap_8 FILLER_6_340 ();
 sg13g2_decap_8 FILLER_6_347 ();
 sg13g2_decap_8 FILLER_6_354 ();
 sg13g2_decap_8 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_368 ();
 sg13g2_decap_8 FILLER_6_375 ();
 sg13g2_decap_8 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_6_389 ();
 sg13g2_decap_8 FILLER_6_396 ();
 sg13g2_decap_4 FILLER_6_403 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_4 FILLER_7_238 ();
 sg13g2_fill_2 FILLER_7_242 ();
 sg13g2_decap_4 FILLER_7_275 ();
 sg13g2_decap_8 FILLER_7_283 ();
 sg13g2_decap_8 FILLER_7_290 ();
 sg13g2_decap_4 FILLER_7_297 ();
 sg13g2_fill_2 FILLER_7_301 ();
 sg13g2_decap_4 FILLER_7_316 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_4 FILLER_7_350 ();
 sg13g2_fill_1 FILLER_7_354 ();
 sg13g2_decap_4 FILLER_7_359 ();
 sg13g2_fill_1 FILLER_7_363 ();
 sg13g2_decap_8 FILLER_7_379 ();
 sg13g2_decap_8 FILLER_7_386 ();
 sg13g2_decap_8 FILLER_7_393 ();
 sg13g2_decap_8 FILLER_7_400 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_fill_2 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_149 ();
 sg13g2_decap_8 FILLER_8_156 ();
 sg13g2_decap_8 FILLER_8_163 ();
 sg13g2_decap_8 FILLER_8_170 ();
 sg13g2_decap_8 FILLER_8_177 ();
 sg13g2_decap_8 FILLER_8_184 ();
 sg13g2_decap_8 FILLER_8_191 ();
 sg13g2_decap_8 FILLER_8_198 ();
 sg13g2_decap_8 FILLER_8_205 ();
 sg13g2_decap_8 FILLER_8_212 ();
 sg13g2_decap_8 FILLER_8_219 ();
 sg13g2_decap_8 FILLER_8_226 ();
 sg13g2_decap_8 FILLER_8_233 ();
 sg13g2_fill_2 FILLER_8_267 ();
 sg13g2_fill_1 FILLER_8_269 ();
 sg13g2_fill_1 FILLER_8_325 ();
 sg13g2_fill_2 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_395 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_4 FILLER_9_98 ();
 sg13g2_fill_1 FILLER_9_102 ();
 sg13g2_fill_2 FILLER_9_107 ();
 sg13g2_decap_8 FILLER_9_113 ();
 sg13g2_decap_4 FILLER_9_120 ();
 sg13g2_fill_1 FILLER_9_132 ();
 sg13g2_decap_8 FILLER_9_151 ();
 sg13g2_decap_8 FILLER_9_158 ();
 sg13g2_decap_8 FILLER_9_165 ();
 sg13g2_decap_4 FILLER_9_172 ();
 sg13g2_fill_2 FILLER_9_176 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_fill_1 FILLER_9_217 ();
 sg13g2_fill_2 FILLER_9_251 ();
 sg13g2_fill_1 FILLER_9_253 ();
 sg13g2_fill_1 FILLER_9_265 ();
 sg13g2_fill_2 FILLER_9_284 ();
 sg13g2_fill_1 FILLER_9_286 ();
 sg13g2_decap_4 FILLER_9_309 ();
 sg13g2_decap_4 FILLER_9_323 ();
 sg13g2_fill_1 FILLER_9_332 ();
 sg13g2_fill_2 FILLER_9_341 ();
 sg13g2_fill_1 FILLER_9_343 ();
 sg13g2_fill_2 FILLER_9_353 ();
 sg13g2_fill_2 FILLER_9_364 ();
 sg13g2_fill_1 FILLER_9_366 ();
 sg13g2_fill_1 FILLER_9_381 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_4 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_78 ();
 sg13g2_decap_4 FILLER_10_85 ();
 sg13g2_fill_1 FILLER_10_89 ();
 sg13g2_decap_4 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_4 FILLER_10_217 ();
 sg13g2_fill_2 FILLER_10_221 ();
 sg13g2_decap_4 FILLER_10_227 ();
 sg13g2_fill_2 FILLER_10_231 ();
 sg13g2_fill_2 FILLER_10_256 ();
 sg13g2_fill_1 FILLER_10_286 ();
 sg13g2_decap_4 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_4 FILLER_11_63 ();
 sg13g2_fill_1 FILLER_11_67 ();
 sg13g2_fill_2 FILLER_11_96 ();
 sg13g2_fill_2 FILLER_11_116 ();
 sg13g2_fill_2 FILLER_11_136 ();
 sg13g2_fill_1 FILLER_11_155 ();
 sg13g2_fill_1 FILLER_11_183 ();
 sg13g2_fill_1 FILLER_11_201 ();
 sg13g2_fill_1 FILLER_11_256 ();
 sg13g2_decap_4 FILLER_11_287 ();
 sg13g2_fill_1 FILLER_11_313 ();
 sg13g2_decap_8 FILLER_11_321 ();
 sg13g2_decap_8 FILLER_11_328 ();
 sg13g2_fill_2 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_4 FILLER_12_84 ();
 sg13g2_fill_2 FILLER_12_106 ();
 sg13g2_fill_1 FILLER_12_140 ();
 sg13g2_decap_4 FILLER_12_154 ();
 sg13g2_fill_1 FILLER_12_158 ();
 sg13g2_fill_2 FILLER_12_178 ();
 sg13g2_fill_1 FILLER_12_180 ();
 sg13g2_fill_2 FILLER_12_195 ();
 sg13g2_fill_1 FILLER_12_197 ();
 sg13g2_decap_8 FILLER_12_220 ();
 sg13g2_decap_4 FILLER_12_227 ();
 sg13g2_fill_2 FILLER_12_231 ();
 sg13g2_decap_4 FILLER_12_237 ();
 sg13g2_fill_2 FILLER_12_241 ();
 sg13g2_fill_1 FILLER_12_320 ();
 sg13g2_decap_4 FILLER_12_330 ();
 sg13g2_fill_1 FILLER_12_334 ();
 sg13g2_fill_2 FILLER_12_376 ();
 sg13g2_fill_1 FILLER_12_378 ();
 sg13g2_decap_4 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_fill_1 FILLER_13_70 ();
 sg13g2_fill_2 FILLER_13_153 ();
 sg13g2_fill_1 FILLER_13_155 ();
 sg13g2_fill_1 FILLER_13_168 ();
 sg13g2_decap_4 FILLER_13_173 ();
 sg13g2_fill_1 FILLER_13_177 ();
 sg13g2_fill_2 FILLER_13_222 ();
 sg13g2_fill_2 FILLER_13_233 ();
 sg13g2_fill_1 FILLER_13_275 ();
 sg13g2_fill_1 FILLER_13_308 ();
 sg13g2_fill_2 FILLER_13_336 ();
 sg13g2_fill_1 FILLER_13_338 ();
 sg13g2_fill_2 FILLER_13_345 ();
 sg13g2_fill_2 FILLER_13_379 ();
 sg13g2_fill_1 FILLER_13_381 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_fill_2 FILLER_14_70 ();
 sg13g2_fill_1 FILLER_14_72 ();
 sg13g2_decap_4 FILLER_14_147 ();
 sg13g2_decap_4 FILLER_14_164 ();
 sg13g2_decap_4 FILLER_14_173 ();
 sg13g2_fill_2 FILLER_14_195 ();
 sg13g2_fill_1 FILLER_14_206 ();
 sg13g2_fill_1 FILLER_14_239 ();
 sg13g2_decap_8 FILLER_14_244 ();
 sg13g2_decap_4 FILLER_14_251 ();
 sg13g2_fill_2 FILLER_14_255 ();
 sg13g2_decap_4 FILLER_14_271 ();
 sg13g2_fill_2 FILLER_14_294 ();
 sg13g2_fill_1 FILLER_14_296 ();
 sg13g2_fill_1 FILLER_14_308 ();
 sg13g2_fill_2 FILLER_14_322 ();
 sg13g2_fill_1 FILLER_14_324 ();
 sg13g2_fill_2 FILLER_14_344 ();
 sg13g2_fill_1 FILLER_14_358 ();
 sg13g2_fill_1 FILLER_14_363 ();
 sg13g2_fill_2 FILLER_14_382 ();
 sg13g2_fill_1 FILLER_14_384 ();
 sg13g2_decap_4 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_fill_2 FILLER_15_70 ();
 sg13g2_fill_1 FILLER_15_100 ();
 sg13g2_fill_2 FILLER_15_145 ();
 sg13g2_decap_4 FILLER_15_174 ();
 sg13g2_fill_2 FILLER_15_178 ();
 sg13g2_decap_4 FILLER_15_188 ();
 sg13g2_fill_2 FILLER_15_242 ();
 sg13g2_fill_2 FILLER_15_302 ();
 sg13g2_fill_1 FILLER_15_322 ();
 sg13g2_fill_2 FILLER_15_328 ();
 sg13g2_fill_1 FILLER_15_357 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_fill_2 FILLER_16_70 ();
 sg13g2_fill_1 FILLER_16_72 ();
 sg13g2_fill_2 FILLER_16_105 ();
 sg13g2_fill_1 FILLER_16_146 ();
 sg13g2_fill_1 FILLER_16_155 ();
 sg13g2_fill_1 FILLER_16_206 ();
 sg13g2_fill_2 FILLER_16_330 ();
 sg13g2_fill_1 FILLER_16_394 ();
 sg13g2_decap_4 FILLER_16_404 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_fill_1 FILLER_17_124 ();
 sg13g2_fill_1 FILLER_17_134 ();
 sg13g2_fill_1 FILLER_17_162 ();
 sg13g2_decap_8 FILLER_17_186 ();
 sg13g2_fill_2 FILLER_17_202 ();
 sg13g2_fill_1 FILLER_17_253 ();
 sg13g2_fill_2 FILLER_17_290 ();
 sg13g2_fill_1 FILLER_17_292 ();
 sg13g2_fill_2 FILLER_17_302 ();
 sg13g2_fill_1 FILLER_17_327 ();
 sg13g2_fill_2 FILLER_17_343 ();
 sg13g2_fill_1 FILLER_17_362 ();
 sg13g2_decap_8 FILLER_17_394 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_4 FILLER_18_70 ();
 sg13g2_fill_1 FILLER_18_74 ();
 sg13g2_decap_8 FILLER_18_79 ();
 sg13g2_fill_1 FILLER_18_129 ();
 sg13g2_fill_1 FILLER_18_147 ();
 sg13g2_fill_1 FILLER_18_157 ();
 sg13g2_fill_2 FILLER_18_234 ();
 sg13g2_fill_1 FILLER_18_236 ();
 sg13g2_fill_2 FILLER_18_291 ();
 sg13g2_decap_4 FILLER_18_320 ();
 sg13g2_fill_1 FILLER_18_333 ();
 sg13g2_fill_2 FILLER_18_349 ();
 sg13g2_fill_2 FILLER_18_360 ();
 sg13g2_fill_1 FILLER_18_362 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_fill_2 FILLER_19_107 ();
 sg13g2_decap_8 FILLER_19_190 ();
 sg13g2_decap_8 FILLER_19_197 ();
 sg13g2_fill_2 FILLER_19_204 ();
 sg13g2_fill_1 FILLER_19_206 ();
 sg13g2_fill_2 FILLER_19_228 ();
 sg13g2_decap_4 FILLER_19_239 ();
 sg13g2_decap_8 FILLER_19_247 ();
 sg13g2_decap_4 FILLER_19_254 ();
 sg13g2_fill_2 FILLER_19_258 ();
 sg13g2_fill_2 FILLER_19_300 ();
 sg13g2_fill_1 FILLER_19_302 ();
 sg13g2_decap_4 FILLER_19_312 ();
 sg13g2_fill_1 FILLER_19_348 ();
 sg13g2_fill_1 FILLER_19_363 ();
 sg13g2_fill_2 FILLER_19_382 ();
 sg13g2_fill_1 FILLER_19_393 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_fill_2 FILLER_20_77 ();
 sg13g2_fill_2 FILLER_20_97 ();
 sg13g2_fill_1 FILLER_20_99 ();
 sg13g2_fill_2 FILLER_20_114 ();
 sg13g2_fill_2 FILLER_20_125 ();
 sg13g2_fill_1 FILLER_20_136 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_4 FILLER_20_168 ();
 sg13g2_fill_1 FILLER_20_172 ();
 sg13g2_fill_1 FILLER_20_201 ();
 sg13g2_fill_2 FILLER_20_229 ();
 sg13g2_fill_1 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_4 FILLER_20_252 ();
 sg13g2_fill_1 FILLER_20_256 ();
 sg13g2_fill_1 FILLER_20_284 ();
 sg13g2_decap_8 FILLER_20_318 ();
 sg13g2_decap_4 FILLER_20_325 ();
 sg13g2_fill_1 FILLER_20_333 ();
 sg13g2_fill_1 FILLER_20_367 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_4 FILLER_21_70 ();
 sg13g2_fill_1 FILLER_21_74 ();
 sg13g2_fill_2 FILLER_21_120 ();
 sg13g2_fill_1 FILLER_21_131 ();
 sg13g2_fill_1 FILLER_21_135 ();
 sg13g2_fill_2 FILLER_21_141 ();
 sg13g2_fill_1 FILLER_21_143 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_4 FILLER_21_154 ();
 sg13g2_fill_1 FILLER_21_158 ();
 sg13g2_decap_4 FILLER_21_172 ();
 sg13g2_fill_1 FILLER_21_176 ();
 sg13g2_fill_2 FILLER_21_195 ();
 sg13g2_fill_1 FILLER_21_197 ();
 sg13g2_decap_8 FILLER_21_216 ();
 sg13g2_fill_2 FILLER_21_223 ();
 sg13g2_fill_1 FILLER_21_225 ();
 sg13g2_decap_8 FILLER_21_254 ();
 sg13g2_fill_1 FILLER_21_261 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_4 FILLER_21_280 ();
 sg13g2_fill_1 FILLER_21_284 ();
 sg13g2_decap_8 FILLER_21_304 ();
 sg13g2_decap_8 FILLER_21_311 ();
 sg13g2_fill_1 FILLER_21_318 ();
 sg13g2_decap_4 FILLER_21_335 ();
 sg13g2_fill_2 FILLER_21_339 ();
 sg13g2_fill_1 FILLER_21_354 ();
 sg13g2_fill_1 FILLER_21_363 ();
 sg13g2_decap_4 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_4 FILLER_22_84 ();
 sg13g2_fill_2 FILLER_22_132 ();
 sg13g2_fill_1 FILLER_22_134 ();
 sg13g2_fill_1 FILLER_22_153 ();
 sg13g2_decap_8 FILLER_22_213 ();
 sg13g2_fill_2 FILLER_22_220 ();
 sg13g2_fill_2 FILLER_22_238 ();
 sg13g2_decap_4 FILLER_22_247 ();
 sg13g2_fill_2 FILLER_22_251 ();
 sg13g2_fill_1 FILLER_22_285 ();
 sg13g2_decap_4 FILLER_22_295 ();
 sg13g2_fill_2 FILLER_22_299 ();
 sg13g2_decap_8 FILLER_22_320 ();
 sg13g2_decap_4 FILLER_22_327 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_fill_1 FILLER_22_350 ();
 sg13g2_fill_1 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_fill_2 FILLER_23_119 ();
 sg13g2_fill_2 FILLER_23_154 ();
 sg13g2_fill_1 FILLER_23_156 ();
 sg13g2_decap_8 FILLER_23_166 ();
 sg13g2_decap_4 FILLER_23_173 ();
 sg13g2_fill_2 FILLER_23_192 ();
 sg13g2_fill_2 FILLER_23_221 ();
 sg13g2_fill_1 FILLER_23_223 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_fill_2 FILLER_23_273 ();
 sg13g2_fill_1 FILLER_23_275 ();
 sg13g2_decap_4 FILLER_23_284 ();
 sg13g2_fill_2 FILLER_23_288 ();
 sg13g2_decap_4 FILLER_23_351 ();
 sg13g2_fill_2 FILLER_23_355 ();
 sg13g2_fill_2 FILLER_23_367 ();
 sg13g2_decap_8 FILLER_23_391 ();
 sg13g2_decap_8 FILLER_23_398 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_fill_2 FILLER_24_84 ();
 sg13g2_fill_1 FILLER_24_86 ();
 sg13g2_fill_2 FILLER_24_125 ();
 sg13g2_decap_4 FILLER_24_174 ();
 sg13g2_fill_1 FILLER_24_178 ();
 sg13g2_decap_4 FILLER_24_184 ();
 sg13g2_decap_8 FILLER_24_199 ();
 sg13g2_decap_8 FILLER_24_206 ();
 sg13g2_fill_2 FILLER_24_213 ();
 sg13g2_fill_1 FILLER_24_215 ();
 sg13g2_fill_1 FILLER_24_231 ();
 sg13g2_fill_2 FILLER_24_262 ();
 sg13g2_fill_1 FILLER_24_264 ();
 sg13g2_decap_8 FILLER_24_289 ();
 sg13g2_fill_2 FILLER_24_301 ();
 sg13g2_fill_1 FILLER_24_303 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_fill_2 FILLER_24_322 ();
 sg13g2_fill_2 FILLER_24_332 ();
 sg13g2_fill_2 FILLER_24_339 ();
 sg13g2_fill_1 FILLER_24_341 ();
 sg13g2_decap_4 FILLER_24_350 ();
 sg13g2_fill_1 FILLER_24_354 ();
 sg13g2_decap_8 FILLER_24_363 ();
 sg13g2_decap_8 FILLER_24_370 ();
 sg13g2_fill_2 FILLER_24_391 ();
 sg13g2_fill_1 FILLER_24_393 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_4 FILLER_25_70 ();
 sg13g2_fill_1 FILLER_25_74 ();
 sg13g2_fill_2 FILLER_25_103 ();
 sg13g2_fill_2 FILLER_25_122 ();
 sg13g2_fill_1 FILLER_25_129 ();
 sg13g2_fill_1 FILLER_25_140 ();
 sg13g2_decap_4 FILLER_25_150 ();
 sg13g2_fill_2 FILLER_25_154 ();
 sg13g2_decap_4 FILLER_25_169 ();
 sg13g2_decap_8 FILLER_25_187 ();
 sg13g2_fill_1 FILLER_25_194 ();
 sg13g2_decap_4 FILLER_25_199 ();
 sg13g2_fill_1 FILLER_25_203 ();
 sg13g2_decap_4 FILLER_25_207 ();
 sg13g2_fill_2 FILLER_25_211 ();
 sg13g2_fill_2 FILLER_25_248 ();
 sg13g2_fill_1 FILLER_25_250 ();
 sg13g2_decap_8 FILLER_25_267 ();
 sg13g2_fill_2 FILLER_25_290 ();
 sg13g2_decap_8 FILLER_25_339 ();
 sg13g2_fill_2 FILLER_25_346 ();
 sg13g2_decap_4 FILLER_25_374 ();
 sg13g2_fill_1 FILLER_25_396 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_fill_2 FILLER_26_77 ();
 sg13g2_fill_1 FILLER_26_79 ();
 sg13g2_fill_2 FILLER_26_84 ();
 sg13g2_fill_2 FILLER_26_124 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_166 ();
 sg13g2_decap_4 FILLER_26_173 ();
 sg13g2_decap_4 FILLER_26_184 ();
 sg13g2_fill_2 FILLER_26_188 ();
 sg13g2_decap_8 FILLER_26_207 ();
 sg13g2_decap_4 FILLER_26_214 ();
 sg13g2_fill_1 FILLER_26_218 ();
 sg13g2_decap_8 FILLER_26_234 ();
 sg13g2_decap_4 FILLER_26_241 ();
 sg13g2_fill_2 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_268 ();
 sg13g2_fill_2 FILLER_26_275 ();
 sg13g2_fill_1 FILLER_26_277 ();
 sg13g2_fill_1 FILLER_26_283 ();
 sg13g2_decap_4 FILLER_26_316 ();
 sg13g2_fill_2 FILLER_26_320 ();
 sg13g2_decap_8 FILLER_26_342 ();
 sg13g2_decap_4 FILLER_26_349 ();
 sg13g2_fill_2 FILLER_26_353 ();
 sg13g2_decap_8 FILLER_26_365 ();
 sg13g2_decap_8 FILLER_26_372 ();
 sg13g2_fill_2 FILLER_26_384 ();
 sg13g2_fill_1 FILLER_26_386 ();
 sg13g2_decap_4 FILLER_26_404 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_fill_1 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_82 ();
 sg13g2_fill_2 FILLER_27_89 ();
 sg13g2_fill_1 FILLER_27_91 ();
 sg13g2_fill_2 FILLER_27_137 ();
 sg13g2_fill_2 FILLER_27_144 ();
 sg13g2_decap_4 FILLER_27_150 ();
 sg13g2_decap_8 FILLER_27_169 ();
 sg13g2_fill_1 FILLER_27_188 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_4 FILLER_27_203 ();
 sg13g2_fill_2 FILLER_27_207 ();
 sg13g2_fill_2 FILLER_27_282 ();
 sg13g2_fill_2 FILLER_27_316 ();
 sg13g2_decap_4 FILLER_27_329 ();
 sg13g2_decap_8 FILLER_27_352 ();
 sg13g2_fill_2 FILLER_27_367 ();
 sg13g2_fill_1 FILLER_27_369 ();
 sg13g2_fill_1 FILLER_27_380 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_fill_2 FILLER_28_70 ();
 sg13g2_fill_1 FILLER_28_72 ();
 sg13g2_fill_1 FILLER_28_101 ();
 sg13g2_fill_1 FILLER_28_111 ();
 sg13g2_decap_4 FILLER_28_121 ();
 sg13g2_fill_1 FILLER_28_125 ();
 sg13g2_fill_2 FILLER_28_158 ();
 sg13g2_fill_1 FILLER_28_180 ();
 sg13g2_fill_2 FILLER_28_186 ();
 sg13g2_fill_1 FILLER_28_188 ();
 sg13g2_decap_8 FILLER_28_204 ();
 sg13g2_decap_8 FILLER_28_211 ();
 sg13g2_fill_2 FILLER_28_222 ();
 sg13g2_fill_1 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_234 ();
 sg13g2_decap_8 FILLER_28_241 ();
 sg13g2_decap_8 FILLER_28_248 ();
 sg13g2_decap_8 FILLER_28_282 ();
 sg13g2_decap_8 FILLER_28_289 ();
 sg13g2_fill_2 FILLER_28_296 ();
 sg13g2_fill_1 FILLER_28_298 ();
 sg13g2_decap_8 FILLER_28_304 ();
 sg13g2_decap_4 FILLER_28_311 ();
 sg13g2_decap_8 FILLER_28_319 ();
 sg13g2_fill_2 FILLER_28_344 ();
 sg13g2_fill_1 FILLER_28_346 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_fill_2 FILLER_29_95 ();
 sg13g2_fill_1 FILLER_29_118 ();
 sg13g2_decap_8 FILLER_29_142 ();
 sg13g2_fill_2 FILLER_29_152 ();
 sg13g2_fill_1 FILLER_29_160 ();
 sg13g2_fill_2 FILLER_29_182 ();
 sg13g2_fill_2 FILLER_29_212 ();
 sg13g2_fill_1 FILLER_29_214 ();
 sg13g2_decap_8 FILLER_29_235 ();
 sg13g2_fill_2 FILLER_29_242 ();
 sg13g2_fill_1 FILLER_29_244 ();
 sg13g2_fill_1 FILLER_29_249 ();
 sg13g2_fill_2 FILLER_29_274 ();
 sg13g2_fill_1 FILLER_29_276 ();
 sg13g2_decap_4 FILLER_29_290 ();
 sg13g2_fill_1 FILLER_29_312 ();
 sg13g2_fill_1 FILLER_29_317 ();
 sg13g2_decap_8 FILLER_29_332 ();
 sg13g2_decap_4 FILLER_29_339 ();
 sg13g2_fill_1 FILLER_29_343 ();
 sg13g2_fill_1 FILLER_29_392 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_fill_2 FILLER_30_84 ();
 sg13g2_decap_4 FILLER_30_123 ();
 sg13g2_fill_1 FILLER_30_127 ();
 sg13g2_fill_1 FILLER_30_155 ();
 sg13g2_fill_2 FILLER_30_165 ();
 sg13g2_fill_1 FILLER_30_180 ();
 sg13g2_fill_2 FILLER_30_188 ();
 sg13g2_fill_2 FILLER_30_200 ();
 sg13g2_decap_8 FILLER_30_218 ();
 sg13g2_fill_1 FILLER_30_225 ();
 sg13g2_fill_1 FILLER_30_237 ();
 sg13g2_fill_2 FILLER_30_248 ();
 sg13g2_decap_4 FILLER_30_254 ();
 sg13g2_fill_1 FILLER_30_258 ();
 sg13g2_decap_8 FILLER_30_263 ();
 sg13g2_decap_4 FILLER_30_270 ();
 sg13g2_fill_1 FILLER_30_274 ();
 sg13g2_decap_4 FILLER_30_304 ();
 sg13g2_fill_1 FILLER_30_308 ();
 sg13g2_fill_2 FILLER_30_315 ();
 sg13g2_fill_1 FILLER_30_317 ();
 sg13g2_decap_8 FILLER_30_333 ();
 sg13g2_fill_1 FILLER_30_340 ();
 sg13g2_fill_1 FILLER_30_361 ();
 sg13g2_fill_2 FILLER_30_371 ();
 sg13g2_fill_1 FILLER_30_373 ();
 sg13g2_fill_2 FILLER_30_378 ();
 sg13g2_fill_1 FILLER_30_380 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_fill_2 FILLER_31_118 ();
 sg13g2_fill_2 FILLER_31_133 ();
 sg13g2_fill_1 FILLER_31_149 ();
 sg13g2_fill_2 FILLER_31_159 ();
 sg13g2_fill_1 FILLER_31_180 ();
 sg13g2_decap_8 FILLER_31_194 ();
 sg13g2_fill_2 FILLER_31_201 ();
 sg13g2_decap_4 FILLER_31_209 ();
 sg13g2_decap_8 FILLER_31_223 ();
 sg13g2_decap_8 FILLER_31_230 ();
 sg13g2_decap_4 FILLER_31_237 ();
 sg13g2_fill_1 FILLER_31_241 ();
 sg13g2_fill_2 FILLER_31_252 ();
 sg13g2_decap_4 FILLER_31_276 ();
 sg13g2_fill_2 FILLER_31_285 ();
 sg13g2_fill_1 FILLER_31_287 ();
 sg13g2_decap_8 FILLER_31_304 ();
 sg13g2_decap_8 FILLER_31_311 ();
 sg13g2_fill_1 FILLER_31_323 ();
 sg13g2_decap_4 FILLER_31_337 ();
 sg13g2_fill_2 FILLER_31_359 ();
 sg13g2_decap_4 FILLER_31_365 ();
 sg13g2_fill_1 FILLER_31_369 ();
 sg13g2_decap_4 FILLER_31_374 ();
 sg13g2_fill_1 FILLER_31_378 ();
 sg13g2_decap_4 FILLER_31_383 ();
 sg13g2_decap_8 FILLER_31_391 ();
 sg13g2_decap_8 FILLER_31_398 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_160 ();
 sg13g2_fill_2 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_197 ();
 sg13g2_decap_8 FILLER_32_204 ();
 sg13g2_decap_4 FILLER_32_211 ();
 sg13g2_decap_4 FILLER_32_231 ();
 sg13g2_decap_8 FILLER_32_244 ();
 sg13g2_fill_2 FILLER_32_251 ();
 sg13g2_decap_4 FILLER_32_258 ();
 sg13g2_decap_4 FILLER_32_267 ();
 sg13g2_decap_8 FILLER_32_277 ();
 sg13g2_decap_8 FILLER_32_303 ();
 sg13g2_fill_1 FILLER_32_310 ();
 sg13g2_fill_1 FILLER_32_322 ();
 sg13g2_fill_2 FILLER_32_327 ();
 sg13g2_fill_1 FILLER_32_337 ();
 sg13g2_decap_4 FILLER_32_342 ();
 sg13g2_fill_2 FILLER_32_351 ();
 sg13g2_decap_8 FILLER_32_370 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_4 FILLER_33_98 ();
 sg13g2_fill_1 FILLER_33_102 ();
 sg13g2_decap_8 FILLER_33_107 ();
 sg13g2_decap_8 FILLER_33_114 ();
 sg13g2_decap_8 FILLER_33_121 ();
 sg13g2_decap_8 FILLER_33_128 ();
 sg13g2_fill_2 FILLER_33_135 ();
 sg13g2_fill_2 FILLER_33_145 ();
 sg13g2_decap_8 FILLER_33_151 ();
 sg13g2_decap_8 FILLER_33_158 ();
 sg13g2_fill_1 FILLER_33_165 ();
 sg13g2_fill_2 FILLER_33_185 ();
 sg13g2_fill_1 FILLER_33_187 ();
 sg13g2_decap_4 FILLER_33_225 ();
 sg13g2_fill_1 FILLER_33_229 ();
 sg13g2_fill_2 FILLER_33_258 ();
 sg13g2_fill_1 FILLER_33_260 ();
 sg13g2_fill_2 FILLER_33_288 ();
 sg13g2_fill_1 FILLER_33_295 ();
 sg13g2_fill_2 FILLER_33_345 ();
 sg13g2_fill_1 FILLER_33_347 ();
 sg13g2_fill_2 FILLER_33_353 ();
 sg13g2_fill_2 FILLER_33_383 ();
 sg13g2_fill_1 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_391 ();
 sg13g2_decap_8 FILLER_33_398 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_fill_1 FILLER_34_140 ();
 sg13g2_fill_1 FILLER_34_169 ();
 sg13g2_fill_2 FILLER_34_218 ();
 sg13g2_fill_1 FILLER_34_220 ();
 sg13g2_decap_4 FILLER_34_230 ();
 sg13g2_fill_2 FILLER_34_234 ();
 sg13g2_decap_4 FILLER_34_240 ();
 sg13g2_fill_2 FILLER_34_244 ();
 sg13g2_fill_1 FILLER_34_292 ();
 sg13g2_decap_8 FILLER_34_333 ();
 sg13g2_decap_4 FILLER_34_365 ();
 sg13g2_fill_2 FILLER_34_369 ();
 sg13g2_fill_2 FILLER_34_380 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_fill_2 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_153 ();
 sg13g2_decap_4 FILLER_35_160 ();
 sg13g2_fill_1 FILLER_35_164 ();
 sg13g2_decap_4 FILLER_35_177 ();
 sg13g2_fill_2 FILLER_35_181 ();
 sg13g2_decap_4 FILLER_35_187 ();
 sg13g2_fill_2 FILLER_35_191 ();
 sg13g2_fill_1 FILLER_35_200 ();
 sg13g2_fill_2 FILLER_35_210 ();
 sg13g2_fill_1 FILLER_35_212 ();
 sg13g2_decap_8 FILLER_35_241 ();
 sg13g2_decap_8 FILLER_35_248 ();
 sg13g2_decap_4 FILLER_35_255 ();
 sg13g2_fill_2 FILLER_35_259 ();
 sg13g2_decap_8 FILLER_35_269 ();
 sg13g2_decap_8 FILLER_35_276 ();
 sg13g2_fill_1 FILLER_35_283 ();
 sg13g2_decap_4 FILLER_35_293 ();
 sg13g2_decap_4 FILLER_35_301 ();
 sg13g2_decap_8 FILLER_35_309 ();
 sg13g2_decap_8 FILLER_35_316 ();
 sg13g2_decap_4 FILLER_35_323 ();
 sg13g2_decap_8 FILLER_35_332 ();
 sg13g2_fill_1 FILLER_35_339 ();
 sg13g2_fill_2 FILLER_35_384 ();
 sg13g2_fill_1 FILLER_35_386 ();
 sg13g2_decap_8 FILLER_35_391 ();
 sg13g2_decap_8 FILLER_35_398 ();
 sg13g2_decap_4 FILLER_35_405 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_4 FILLER_36_140 ();
 sg13g2_fill_2 FILLER_36_186 ();
 sg13g2_fill_1 FILLER_36_188 ();
 sg13g2_fill_1 FILLER_36_199 ();
 sg13g2_fill_2 FILLER_36_205 ();
 sg13g2_fill_2 FILLER_36_213 ();
 sg13g2_fill_1 FILLER_36_215 ();
 sg13g2_decap_8 FILLER_36_229 ();
 sg13g2_fill_2 FILLER_36_236 ();
 sg13g2_decap_4 FILLER_36_269 ();
 sg13g2_fill_1 FILLER_36_273 ();
 sg13g2_fill_2 FILLER_36_286 ();
 sg13g2_fill_2 FILLER_36_311 ();
 sg13g2_fill_1 FILLER_36_313 ();
 sg13g2_fill_2 FILLER_36_324 ();
 sg13g2_fill_1 FILLER_36_335 ();
 sg13g2_fill_2 FILLER_36_344 ();
 sg13g2_fill_1 FILLER_36_359 ();
 sg13g2_fill_2 FILLER_36_373 ();
 sg13g2_decap_4 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_4 FILLER_37_168 ();
 sg13g2_fill_1 FILLER_37_197 ();
 sg13g2_decap_8 FILLER_37_235 ();
 sg13g2_fill_1 FILLER_37_242 ();
 sg13g2_decap_8 FILLER_37_247 ();
 sg13g2_fill_2 FILLER_37_254 ();
 sg13g2_fill_1 FILLER_37_256 ();
 sg13g2_decap_8 FILLER_37_261 ();
 sg13g2_decap_8 FILLER_37_268 ();
 sg13g2_fill_2 FILLER_37_275 ();
 sg13g2_fill_1 FILLER_37_282 ();
 sg13g2_decap_8 FILLER_37_301 ();
 sg13g2_fill_2 FILLER_37_326 ();
 sg13g2_fill_1 FILLER_37_328 ();
 sg13g2_fill_1 FILLER_37_342 ();
 sg13g2_fill_2 FILLER_37_352 ();
 sg13g2_fill_2 FILLER_37_372 ();
 sg13g2_fill_1 FILLER_37_374 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_208 ();
 sg13g2_fill_2 FILLER_38_212 ();
 sg13g2_fill_2 FILLER_38_249 ();
 sg13g2_fill_1 FILLER_38_251 ();
 sg13g2_decap_8 FILLER_38_279 ();
 sg13g2_fill_2 FILLER_38_286 ();
 sg13g2_fill_2 FILLER_38_324 ();
 sg13g2_fill_1 FILLER_38_326 ();
 sg13g2_fill_1 FILLER_38_355 ();
 sg13g2_decap_8 FILLER_38_397 ();
 sg13g2_decap_4 FILLER_38_404 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
endmodule
