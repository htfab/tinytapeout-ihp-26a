module tt_um_dranoel06_SAP1 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire clknet_0_clk;
 wire \cpu0.a_reg[0] ;
 wire \cpu0.a_reg[1] ;
 wire \cpu0.a_reg[2] ;
 wire \cpu0.a_reg[3] ;
 wire \cpu0.a_reg[4] ;
 wire \cpu0.a_reg[5] ;
 wire \cpu0.a_reg[6] ;
 wire \cpu0.a_reg[7] ;
 wire \cpu0.b_reg[0] ;
 wire \cpu0.b_reg[1] ;
 wire \cpu0.b_reg[2] ;
 wire \cpu0.b_reg[3] ;
 wire \cpu0.b_reg[4] ;
 wire \cpu0.b_reg[5] ;
 wire \cpu0.b_reg[6] ;
 wire \cpu0.b_reg[7] ;
 wire \cpu0.carry_flag ;
 wire \cpu0.ir[0] ;
 wire \cpu0.ir[1] ;
 wire \cpu0.ir[2] ;
 wire \cpu0.ir[3] ;
 wire \cpu0.ir[4] ;
 wire \cpu0.ir[5] ;
 wire \cpu0.ir[6] ;
 wire \cpu0.ir[7] ;
 wire \cpu0.mar[0] ;
 wire \cpu0.mar[1] ;
 wire \cpu0.mar[2] ;
 wire \cpu0.mar[3] ;
 wire \cpu0.pc[0] ;
 wire \cpu0.pc[1] ;
 wire \cpu0.pc[2] ;
 wire \cpu0.pc[3] ;
 wire \cpu0.ram[0][0] ;
 wire \cpu0.ram[0][1] ;
 wire \cpu0.ram[0][2] ;
 wire \cpu0.ram[0][3] ;
 wire \cpu0.ram[0][4] ;
 wire \cpu0.ram[0][5] ;
 wire \cpu0.ram[0][6] ;
 wire \cpu0.ram[0][7] ;
 wire \cpu0.ram[10][0] ;
 wire \cpu0.ram[10][1] ;
 wire \cpu0.ram[10][2] ;
 wire \cpu0.ram[10][3] ;
 wire \cpu0.ram[10][4] ;
 wire \cpu0.ram[10][5] ;
 wire \cpu0.ram[10][6] ;
 wire \cpu0.ram[10][7] ;
 wire \cpu0.ram[11][0] ;
 wire \cpu0.ram[11][1] ;
 wire \cpu0.ram[11][2] ;
 wire \cpu0.ram[11][3] ;
 wire \cpu0.ram[11][4] ;
 wire \cpu0.ram[11][5] ;
 wire \cpu0.ram[11][6] ;
 wire \cpu0.ram[11][7] ;
 wire \cpu0.ram[12][0] ;
 wire \cpu0.ram[12][1] ;
 wire \cpu0.ram[12][2] ;
 wire \cpu0.ram[12][3] ;
 wire \cpu0.ram[12][4] ;
 wire \cpu0.ram[12][5] ;
 wire \cpu0.ram[12][6] ;
 wire \cpu0.ram[12][7] ;
 wire \cpu0.ram[13][0] ;
 wire \cpu0.ram[13][1] ;
 wire \cpu0.ram[13][2] ;
 wire \cpu0.ram[13][3] ;
 wire \cpu0.ram[13][4] ;
 wire \cpu0.ram[13][5] ;
 wire \cpu0.ram[13][6] ;
 wire \cpu0.ram[13][7] ;
 wire \cpu0.ram[14][0] ;
 wire \cpu0.ram[14][1] ;
 wire \cpu0.ram[14][2] ;
 wire \cpu0.ram[14][3] ;
 wire \cpu0.ram[14][4] ;
 wire \cpu0.ram[14][5] ;
 wire \cpu0.ram[14][6] ;
 wire \cpu0.ram[14][7] ;
 wire \cpu0.ram[15][0] ;
 wire \cpu0.ram[15][1] ;
 wire \cpu0.ram[15][2] ;
 wire \cpu0.ram[15][3] ;
 wire \cpu0.ram[15][4] ;
 wire \cpu0.ram[15][5] ;
 wire \cpu0.ram[15][6] ;
 wire \cpu0.ram[15][7] ;
 wire \cpu0.ram[1][0] ;
 wire \cpu0.ram[1][1] ;
 wire \cpu0.ram[1][2] ;
 wire \cpu0.ram[1][3] ;
 wire \cpu0.ram[1][4] ;
 wire \cpu0.ram[1][5] ;
 wire \cpu0.ram[1][6] ;
 wire \cpu0.ram[1][7] ;
 wire \cpu0.ram[2][0] ;
 wire \cpu0.ram[2][1] ;
 wire \cpu0.ram[2][2] ;
 wire \cpu0.ram[2][3] ;
 wire \cpu0.ram[2][4] ;
 wire \cpu0.ram[2][5] ;
 wire \cpu0.ram[2][6] ;
 wire \cpu0.ram[2][7] ;
 wire \cpu0.ram[3][0] ;
 wire \cpu0.ram[3][1] ;
 wire \cpu0.ram[3][2] ;
 wire \cpu0.ram[3][3] ;
 wire \cpu0.ram[3][4] ;
 wire \cpu0.ram[3][5] ;
 wire \cpu0.ram[3][6] ;
 wire \cpu0.ram[3][7] ;
 wire \cpu0.ram[4][0] ;
 wire \cpu0.ram[4][1] ;
 wire \cpu0.ram[4][2] ;
 wire \cpu0.ram[4][3] ;
 wire \cpu0.ram[4][4] ;
 wire \cpu0.ram[4][5] ;
 wire \cpu0.ram[4][6] ;
 wire \cpu0.ram[4][7] ;
 wire \cpu0.ram[5][0] ;
 wire \cpu0.ram[5][1] ;
 wire \cpu0.ram[5][2] ;
 wire \cpu0.ram[5][3] ;
 wire \cpu0.ram[5][4] ;
 wire \cpu0.ram[5][5] ;
 wire \cpu0.ram[5][6] ;
 wire \cpu0.ram[5][7] ;
 wire \cpu0.ram[6][0] ;
 wire \cpu0.ram[6][1] ;
 wire \cpu0.ram[6][2] ;
 wire \cpu0.ram[6][3] ;
 wire \cpu0.ram[6][4] ;
 wire \cpu0.ram[6][5] ;
 wire \cpu0.ram[6][6] ;
 wire \cpu0.ram[6][7] ;
 wire \cpu0.ram[7][0] ;
 wire \cpu0.ram[7][1] ;
 wire \cpu0.ram[7][2] ;
 wire \cpu0.ram[7][3] ;
 wire \cpu0.ram[7][4] ;
 wire \cpu0.ram[7][5] ;
 wire \cpu0.ram[7][6] ;
 wire \cpu0.ram[7][7] ;
 wire \cpu0.ram[8][0] ;
 wire \cpu0.ram[8][1] ;
 wire \cpu0.ram[8][2] ;
 wire \cpu0.ram[8][3] ;
 wire \cpu0.ram[8][4] ;
 wire \cpu0.ram[8][5] ;
 wire \cpu0.ram[8][6] ;
 wire \cpu0.ram[8][7] ;
 wire \cpu0.ram[9][0] ;
 wire \cpu0.ram[9][1] ;
 wire \cpu0.ram[9][2] ;
 wire \cpu0.ram[9][3] ;
 wire \cpu0.ram[9][4] ;
 wire \cpu0.ram[9][5] ;
 wire \cpu0.ram[9][6] ;
 wire \cpu0.ram[9][7] ;
 wire \cpu0.step[0] ;
 wire \cpu0.step[1] ;
 wire \cpu0.step[2] ;
 wire \cpu0.zero_flag ;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;

 sg13g2_inv_1 _0761_ (.Y(_0181_),
    .A(\cpu0.step[0] ));
 sg13g2_inv_2 _0762_ (.Y(_0182_),
    .A(net179));
 sg13g2_inv_1 _0763_ (.Y(_0183_),
    .A(net161));
 sg13g2_inv_4 _0764_ (.A(net159),
    .Y(_0184_));
 sg13g2_inv_1 _0765_ (.Y(_0185_),
    .A(net268));
 sg13g2_inv_1 _0766_ (.Y(_0186_),
    .A(net273));
 sg13g2_inv_1 _0767_ (.Y(_0187_),
    .A(\cpu0.ram[4][2] ));
 sg13g2_inv_1 _0768_ (.Y(_0188_),
    .A(net272));
 sg13g2_inv_1 _0769_ (.Y(_0189_),
    .A(\cpu0.ram[4][3] ));
 sg13g2_inv_1 _0770_ (.Y(_0190_),
    .A(net270));
 sg13g2_inv_1 _0771_ (.Y(_0191_),
    .A(\cpu0.ram[13][4] ));
 sg13g2_inv_1 _0772_ (.Y(_0192_),
    .A(\cpu0.ram[11][5] ));
 sg13g2_inv_1 _0773_ (.Y(_0193_),
    .A(\cpu0.ram[13][5] ));
 sg13g2_inv_1 _0774_ (.Y(_0194_),
    .A(\cpu0.ram[12][6] ));
 sg13g2_nor2b_1 _0775_ (.A(\cpu0.ir[7] ),
    .B_N(\cpu0.ir[6] ),
    .Y(_0195_));
 sg13g2_nand2b_1 _0776_ (.Y(_0196_),
    .B(\cpu0.ir[6] ),
    .A_N(\cpu0.ir[7] ));
 sg13g2_nand2_1 _0777_ (.Y(_0197_),
    .A(net154),
    .B(net179));
 sg13g2_nor3_1 _0778_ (.A(\cpu0.step[0] ),
    .B(\cpu0.step[1] ),
    .C(_0197_),
    .Y(_0198_));
 sg13g2_nor2b_1 _0779_ (.A(net153),
    .B_N(\cpu0.ir[4] ),
    .Y(_0199_));
 sg13g2_nand2b_2 _0780_ (.Y(_0200_),
    .B(\cpu0.ir[4] ),
    .A_N(net153));
 sg13g2_nand3_1 _0781_ (.B(_0198_),
    .C(_0199_),
    .A(_0195_),
    .Y(_0201_));
 sg13g2_nand2b_1 _0782_ (.Y(_0202_),
    .B(_0201_),
    .A_N(net13));
 sg13g2_nor2_1 _0783_ (.A(net13),
    .B(_0201_),
    .Y(_0203_));
 sg13g2_mux2_1 _0784_ (.A0(net11),
    .A1(\cpu0.mar[2] ),
    .S(net146),
    .X(_0204_));
 sg13g2_mux2_1 _0785_ (.A0(net12),
    .A1(\cpu0.mar[3] ),
    .S(net146),
    .X(_0205_));
 sg13g2_nand3b_1 _0786_ (.B(_0204_),
    .C(_0202_),
    .Y(_0206_),
    .A_N(_0205_));
 sg13g2_mux2_1 _0787_ (.A0(net9),
    .A1(\cpu0.mar[0] ),
    .S(net146),
    .X(_0207_));
 sg13g2_mux2_1 _0788_ (.A0(net10),
    .A1(\cpu0.mar[1] ),
    .S(net146),
    .X(_0208_));
 sg13g2_nand2b_2 _0789_ (.Y(_0209_),
    .B(_0207_),
    .A_N(_0208_));
 sg13g2_or2_1 _0790_ (.X(_0210_),
    .B(_0209_),
    .A(_0206_));
 sg13g2_nand3b_1 _0791_ (.B(net179),
    .C(net437),
    .Y(_0211_),
    .A_N(net432));
 sg13g2_nor2_2 _0792_ (.A(net154),
    .B(_0211_),
    .Y(_0212_));
 sg13g2_or2_1 _0793_ (.X(_0213_),
    .B(_0211_),
    .A(net154));
 sg13g2_and2_1 _0794_ (.A(net437),
    .B(net432),
    .X(_0214_));
 sg13g2_nor2b_2 _0795_ (.A(net154),
    .B_N(_0214_),
    .Y(_0215_));
 sg13g2_inv_1 _0796_ (.Y(_0216_),
    .A(_0215_));
 sg13g2_nand2b_1 _0797_ (.Y(_0217_),
    .B(\cpu0.ir[7] ),
    .A_N(\cpu0.ir[6] ));
 sg13g2_nor2_1 _0798_ (.A(_0200_),
    .B(_0217_),
    .Y(_0218_));
 sg13g2_nor3_1 _0799_ (.A(net153),
    .B(\cpu0.ir[4] ),
    .C(_0196_),
    .Y(_0219_));
 sg13g2_nor2b_1 _0800_ (.A(net153),
    .B_N(\cpu0.zero_flag ),
    .Y(_0220_));
 sg13g2_a21oi_1 _0801_ (.A1(\cpu0.carry_flag ),
    .A2(net153),
    .Y(_0221_),
    .B1(_0220_));
 sg13g2_nor4_1 _0802_ (.A(\cpu0.ir[4] ),
    .B(_0216_),
    .C(_0217_),
    .D(_0221_),
    .Y(_0222_));
 sg13g2_mux2_1 _0803_ (.A0(_0222_),
    .A1(_0215_),
    .S(_0219_),
    .X(_0223_));
 sg13g2_nand2_1 _0804_ (.Y(_0224_),
    .A(\cpu0.ir[6] ),
    .B(net153));
 sg13g2_a21oi_1 _0805_ (.A1(_0200_),
    .A2(_0224_),
    .Y(_0225_),
    .B1(\cpu0.ir[7] ));
 sg13g2_a21oi_1 _0806_ (.A1(_0215_),
    .A2(_0218_),
    .Y(_0226_),
    .B1(_0223_));
 sg13g2_nor2_1 _0807_ (.A(\cpu0.ir[7] ),
    .B(\cpu0.ir[6] ),
    .Y(_0227_));
 sg13g2_nand2b_1 _0808_ (.Y(_0228_),
    .B(net153),
    .A_N(\cpu0.ir[4] ));
 sg13g2_nor3_1 _0809_ (.A(\cpu0.ir[7] ),
    .B(\cpu0.ir[6] ),
    .C(_0228_),
    .Y(_0229_));
 sg13g2_a21oi_1 _0810_ (.A1(_0215_),
    .A2(_0225_),
    .Y(_0230_),
    .B1(_0229_));
 sg13g2_nand2_2 _0811_ (.Y(_0231_),
    .A(net179),
    .B(_0215_));
 sg13g2_a221oi_1 _0812_ (.B2(_0226_),
    .C1(_0182_),
    .B1(_0230_),
    .A1(_0216_),
    .Y(_0232_),
    .A2(_0229_));
 sg13g2_inv_1 _0813_ (.Y(_0233_),
    .A(_0232_));
 sg13g2_nand2_1 _0814_ (.Y(_0234_),
    .A(\cpu0.ir[0] ),
    .B(_0232_));
 sg13g2_mux4_1 _0815_ (.S0(net166),
    .A0(\cpu0.ram[4][0] ),
    .A1(\cpu0.ram[5][0] ),
    .A2(\cpu0.ram[6][0] ),
    .A3(\cpu0.ram[7][0] ),
    .S1(net160),
    .X(_0235_));
 sg13g2_mux4_1 _0816_ (.S0(net170),
    .A0(\cpu0.ram[0][0] ),
    .A1(\cpu0.ram[1][0] ),
    .A2(\cpu0.ram[2][0] ),
    .A3(\cpu0.ram[3][0] ),
    .S1(net161),
    .X(_0236_));
 sg13g2_and3_2 _0817_ (.X(_0237_),
    .A(net153),
    .B(\cpu0.ir[4] ),
    .C(_0195_));
 sg13g2_nor2_1 _0818_ (.A(_0229_),
    .B(_0237_),
    .Y(_0238_));
 sg13g2_inv_1 _0819_ (.Y(_0239_),
    .A(_0238_));
 sg13g2_o21ai_1 _0820_ (.B1(_0198_),
    .Y(_0240_),
    .A1(_0218_),
    .A2(_0239_));
 sg13g2_nor2b_1 _0821_ (.A(net437),
    .B_N(net432),
    .Y(_0241_));
 sg13g2_nand2_1 _0822_ (.Y(_0242_),
    .A(net179),
    .B(_0241_));
 sg13g2_nor2_2 _0823_ (.A(net154),
    .B(_0242_),
    .Y(_0243_));
 sg13g2_or2_1 _0824_ (.X(_0244_),
    .B(_0242_),
    .A(net154));
 sg13g2_nand3_1 _0825_ (.B(_0199_),
    .C(_0227_),
    .A(_0198_),
    .Y(_0245_));
 sg13g2_inv_2 _0826_ (.Y(_0246_),
    .A(_0245_));
 sg13g2_and3_2 _0827_ (.X(_0247_),
    .A(net143),
    .B(net149),
    .C(_0245_));
 sg13g2_nand3_1 _0828_ (.B(net149),
    .C(_0245_),
    .A(net143),
    .Y(_0248_));
 sg13g2_mux4_1 _0829_ (.S0(net168),
    .A0(\cpu0.ram[12][0] ),
    .A1(\cpu0.ram[13][0] ),
    .A2(\cpu0.ram[14][0] ),
    .A3(\cpu0.ram[15][0] ),
    .S1(net163),
    .X(_0249_));
 sg13g2_mux4_1 _0830_ (.S0(net176),
    .A0(\cpu0.ram[8][0] ),
    .A1(\cpu0.ram[9][0] ),
    .A2(\cpu0.ram[10][0] ),
    .A3(\cpu0.ram[11][0] ),
    .S1(net165),
    .X(_0250_));
 sg13g2_mux4_1 _0831_ (.S0(_0184_),
    .A0(_0235_),
    .A1(_0236_),
    .A2(_0249_),
    .A3(_0250_),
    .S1(net155),
    .X(_0251_));
 sg13g2_nand3_1 _0832_ (.B(\cpu0.ir[4] ),
    .C(_0227_),
    .A(net271),
    .Y(_0252_));
 sg13g2_or2_1 _0833_ (.X(_0253_),
    .B(_0252_),
    .A(_0231_));
 sg13g2_nand2_2 _0834_ (.Y(_0254_),
    .A(_0201_),
    .B(net145));
 sg13g2_nor2b_1 _0835_ (.A(\cpu0.a_reg[0] ),
    .B_N(\cpu0.b_reg[0] ),
    .Y(_0255_));
 sg13g2_xor2_1 _0836_ (.B(\cpu0.a_reg[0] ),
    .A(\cpu0.b_reg[0] ),
    .X(_0256_));
 sg13g2_nand2_2 _0837_ (.Y(_0257_),
    .A(net154),
    .B(_0241_));
 sg13g2_nor2_1 _0838_ (.A(_0238_),
    .B(_0257_),
    .Y(_0258_));
 sg13g2_nor3_2 _0839_ (.A(_0182_),
    .B(_0238_),
    .C(_0257_),
    .Y(_0259_));
 sg13g2_a22oi_1 _0840_ (.Y(_0260_),
    .B1(_0256_),
    .B2(net144),
    .A2(_0254_),
    .A1(\cpu0.a_reg[0] ));
 sg13g2_a21oi_1 _0841_ (.A1(_0248_),
    .A2(_0251_),
    .Y(_0261_),
    .B1(_0212_));
 sg13g2_nand3_1 _0842_ (.B(_0260_),
    .C(_0261_),
    .A(_0234_),
    .Y(_0262_));
 sg13g2_o21ai_1 _0843_ (.B1(_0262_),
    .Y(_0263_),
    .A1(\cpu0.pc[0] ),
    .A2(_0213_));
 sg13g2_nor2_1 _0844_ (.A(net1),
    .B(net147),
    .Y(_0264_));
 sg13g2_a21oi_2 _0845_ (.B1(_0264_),
    .Y(_0265_),
    .A2(_0263_),
    .A1(net148));
 sg13g2_mux2_1 _0846_ (.A0(net136),
    .A1(net428),
    .S(_0210_),
    .X(_0004_));
 sg13g2_nand3b_1 _0847_ (.B(net154),
    .C(\cpu0.step[0] ),
    .Y(_0266_),
    .A_N(\cpu0.step[1] ));
 sg13g2_nor3_1 _0848_ (.A(_0200_),
    .B(_0217_),
    .C(_0266_),
    .Y(_0267_));
 sg13g2_nor2_2 _0849_ (.A(_0237_),
    .B(_0267_),
    .Y(_0268_));
 sg13g2_a21o_2 _0850_ (.A2(_0257_),
    .A1(_0237_),
    .B1(_0182_),
    .X(_0269_));
 sg13g2_or2_1 _0851_ (.X(_0270_),
    .B(_0269_),
    .A(_0268_));
 sg13g2_o21ai_1 _0852_ (.B1(\cpu0.b_reg[0] ),
    .Y(_0271_),
    .A1(_0268_),
    .A2(_0269_));
 sg13g2_xor2_1 _0853_ (.B(_0271_),
    .A(\cpu0.b_reg[1] ),
    .X(_0272_));
 sg13g2_nand2_1 _0854_ (.Y(_0273_),
    .A(\cpu0.a_reg[1] ),
    .B(_0272_));
 sg13g2_xnor2_1 _0855_ (.Y(_0274_),
    .A(\cpu0.a_reg[1] ),
    .B(_0272_));
 sg13g2_xor2_1 _0856_ (.B(_0274_),
    .A(_0255_),
    .X(_0275_));
 sg13g2_a22oi_1 _0857_ (.Y(_0276_),
    .B1(net144),
    .B2(_0275_),
    .A2(_0254_),
    .A1(\cpu0.a_reg[1] ));
 sg13g2_a21oi_1 _0858_ (.A1(\cpu0.ir[1] ),
    .A2(_0232_),
    .Y(_0277_),
    .B1(_0248_));
 sg13g2_nand2_1 _0859_ (.Y(_0278_),
    .A(_0276_),
    .B(_0277_));
 sg13g2_mux4_1 _0860_ (.S0(net170),
    .A0(\cpu0.ram[0][1] ),
    .A1(\cpu0.ram[1][1] ),
    .A2(\cpu0.ram[2][1] ),
    .A3(\cpu0.ram[3][1] ),
    .S1(net161),
    .X(_0279_));
 sg13g2_mux2_1 _0861_ (.A0(\cpu0.ram[4][1] ),
    .A1(\cpu0.ram[5][1] ),
    .S(net168),
    .X(_0280_));
 sg13g2_mux2_1 _0862_ (.A0(\cpu0.ram[6][1] ),
    .A1(\cpu0.ram[7][1] ),
    .S(net168),
    .X(_0281_));
 sg13g2_nand2_1 _0863_ (.Y(_0282_),
    .A(net161),
    .B(_0281_));
 sg13g2_a21oi_1 _0864_ (.A1(net151),
    .A2(_0280_),
    .Y(_0283_),
    .B1(_0184_));
 sg13g2_a21oi_1 _0865_ (.A1(_0282_),
    .A2(_0283_),
    .Y(_0284_),
    .B1(net155));
 sg13g2_o21ai_1 _0866_ (.B1(_0284_),
    .Y(_0285_),
    .A1(net157),
    .A2(_0279_));
 sg13g2_nand2b_1 _0867_ (.Y(_0286_),
    .B(net172),
    .A_N(\cpu0.ram[13][1] ));
 sg13g2_o21ai_1 _0868_ (.B1(_0286_),
    .Y(_0287_),
    .A1(net172),
    .A2(\cpu0.ram[12][1] ));
 sg13g2_o21ai_1 _0869_ (.B1(net163),
    .Y(_0288_),
    .A1(net173),
    .A2(\cpu0.ram[14][1] ));
 sg13g2_a21oi_1 _0870_ (.A1(net172),
    .A2(_0186_),
    .Y(_0289_),
    .B1(_0288_));
 sg13g2_o21ai_1 _0871_ (.B1(net158),
    .Y(_0290_),
    .A1(net164),
    .A2(_0287_));
 sg13g2_a21oi_1 _0872_ (.A1(net176),
    .A2(_0185_),
    .Y(_0291_),
    .B1(net163));
 sg13g2_o21ai_1 _0873_ (.B1(_0291_),
    .Y(_0292_),
    .A1(net176),
    .A2(\cpu0.ram[8][1] ));
 sg13g2_mux2_1 _0874_ (.A0(\cpu0.ram[10][1] ),
    .A1(\cpu0.ram[11][1] ),
    .S(net176),
    .X(_0293_));
 sg13g2_a21oi_1 _0875_ (.A1(net165),
    .A2(_0293_),
    .Y(_0294_),
    .B1(net158));
 sg13g2_o21ai_1 _0876_ (.B1(net156),
    .Y(_0295_),
    .A1(_0289_),
    .A2(_0290_));
 sg13g2_a21oi_1 _0877_ (.A1(_0292_),
    .A2(_0294_),
    .Y(_0296_),
    .B1(_0295_));
 sg13g2_nor2_1 _0878_ (.A(_0247_),
    .B(_0296_),
    .Y(_0297_));
 sg13g2_a21oi_1 _0879_ (.A1(_0285_),
    .A2(_0297_),
    .Y(_0298_),
    .B1(_0212_));
 sg13g2_a22oi_1 _0880_ (.Y(_0299_),
    .B1(_0278_),
    .B2(_0298_),
    .A2(_0212_),
    .A1(\cpu0.pc[1] ));
 sg13g2_nor2_1 _0881_ (.A(net2),
    .B(net147),
    .Y(_0300_));
 sg13g2_a21oi_2 _0882_ (.B1(_0300_),
    .Y(_0301_),
    .A2(_0299_),
    .A1(net147));
 sg13g2_mux2_1 _0883_ (.A0(net134),
    .A1(net411),
    .S(_0210_),
    .X(_0005_));
 sg13g2_o21ai_1 _0884_ (.B1(_0273_),
    .Y(_0302_),
    .A1(_0255_),
    .A2(_0274_));
 sg13g2_or2_1 _0885_ (.X(_0303_),
    .B(\cpu0.b_reg[0] ),
    .A(\cpu0.b_reg[1] ));
 sg13g2_o21ai_1 _0886_ (.B1(_0303_),
    .Y(_0304_),
    .A1(_0268_),
    .A2(_0269_));
 sg13g2_xor2_1 _0887_ (.B(_0304_),
    .A(\cpu0.b_reg[2] ),
    .X(_0305_));
 sg13g2_or2_1 _0888_ (.X(_0306_),
    .B(_0305_),
    .A(\cpu0.a_reg[2] ));
 sg13g2_and2_1 _0889_ (.A(\cpu0.a_reg[2] ),
    .B(_0305_),
    .X(_0307_));
 sg13g2_xnor2_1 _0890_ (.Y(_0308_),
    .A(\cpu0.a_reg[2] ),
    .B(_0305_));
 sg13g2_xnor2_1 _0891_ (.Y(_0309_),
    .A(_0302_),
    .B(_0308_));
 sg13g2_a221oi_1 _0892_ (.B2(_0309_),
    .C1(_0232_),
    .B1(_0259_),
    .A1(\cpu0.a_reg[2] ),
    .Y(_0310_),
    .A2(_0254_));
 sg13g2_o21ai_1 _0893_ (.B1(_0247_),
    .Y(_0311_),
    .A1(\cpu0.ir[2] ),
    .A2(_0233_));
 sg13g2_nor2b_1 _0894_ (.A(net174),
    .B_N(\cpu0.ram[8][2] ),
    .Y(_0312_));
 sg13g2_a21oi_1 _0895_ (.A1(net174),
    .A2(\cpu0.ram[9][2] ),
    .Y(_0313_),
    .B1(_0312_));
 sg13g2_nand2b_1 _0896_ (.Y(_0314_),
    .B(\cpu0.ram[10][2] ),
    .A_N(net175));
 sg13g2_a21oi_1 _0897_ (.A1(net175),
    .A2(\cpu0.ram[11][2] ),
    .Y(_0315_),
    .B1(net151));
 sg13g2_a221oi_1 _0898_ (.B2(_0315_),
    .C1(net158),
    .B1(_0314_),
    .A1(net152),
    .Y(_0316_),
    .A2(_0313_));
 sg13g2_mux2_1 _0899_ (.A0(\cpu0.ram[12][2] ),
    .A1(\cpu0.ram[13][2] ),
    .S(net172),
    .X(_0317_));
 sg13g2_o21ai_1 _0900_ (.B1(net164),
    .Y(_0318_),
    .A1(net173),
    .A2(_0188_));
 sg13g2_a21oi_1 _0901_ (.A1(net173),
    .A2(\cpu0.ram[15][2] ),
    .Y(_0319_),
    .B1(_0318_));
 sg13g2_o21ai_1 _0902_ (.B1(net158),
    .Y(_0320_),
    .A1(net164),
    .A2(_0317_));
 sg13g2_o21ai_1 _0903_ (.B1(net156),
    .Y(_0321_),
    .A1(_0319_),
    .A2(_0320_));
 sg13g2_nor2_1 _0904_ (.A(_0316_),
    .B(_0321_),
    .Y(_0322_));
 sg13g2_mux4_1 _0905_ (.S0(net170),
    .A0(\cpu0.ram[0][2] ),
    .A1(\cpu0.ram[1][2] ),
    .A2(\cpu0.ram[2][2] ),
    .A3(\cpu0.ram[3][2] ),
    .S1(net162),
    .X(_0323_));
 sg13g2_a21oi_1 _0906_ (.A1(net167),
    .A2(\cpu0.ram[5][2] ),
    .Y(_0324_),
    .B1(net160));
 sg13g2_o21ai_1 _0907_ (.B1(_0324_),
    .Y(_0325_),
    .A1(net166),
    .A2(_0187_));
 sg13g2_nor2b_1 _0908_ (.A(net166),
    .B_N(\cpu0.ram[6][2] ),
    .Y(_0326_));
 sg13g2_a21oi_1 _0909_ (.A1(net166),
    .A2(\cpu0.ram[7][2] ),
    .Y(_0327_),
    .B1(_0326_));
 sg13g2_a21oi_1 _0910_ (.A1(net160),
    .A2(_0327_),
    .Y(_0328_),
    .B1(_0184_));
 sg13g2_a221oi_1 _0911_ (.B2(_0328_),
    .C1(net155),
    .B1(_0325_),
    .A1(_0184_),
    .Y(_0329_),
    .A2(_0323_));
 sg13g2_nor2_1 _0912_ (.A(_0322_),
    .B(_0329_),
    .Y(_0330_));
 sg13g2_a21oi_1 _0913_ (.A1(_0248_),
    .A2(_0330_),
    .Y(_0331_),
    .B1(_0212_));
 sg13g2_o21ai_1 _0914_ (.B1(_0331_),
    .Y(_0332_),
    .A1(_0310_),
    .A2(_0311_));
 sg13g2_o21ai_1 _0915_ (.B1(_0332_),
    .Y(_0333_),
    .A1(\cpu0.pc[2] ),
    .A2(_0213_));
 sg13g2_nor2_1 _0916_ (.A(net3),
    .B(net147),
    .Y(_0334_));
 sg13g2_a21oi_2 _0917_ (.B1(_0334_),
    .Y(_0335_),
    .A2(_0333_),
    .A1(net147));
 sg13g2_mux2_1 _0918_ (.A0(net132),
    .A1(net343),
    .S(_0210_),
    .X(_0006_));
 sg13g2_or2_1 _0919_ (.X(_0336_),
    .B(_0303_),
    .A(\cpu0.b_reg[2] ));
 sg13g2_o21ai_1 _0920_ (.B1(_0336_),
    .Y(_0337_),
    .A1(_0268_),
    .A2(_0269_));
 sg13g2_xor2_1 _0921_ (.B(_0337_),
    .A(\cpu0.b_reg[3] ),
    .X(_0338_));
 sg13g2_or2_1 _0922_ (.X(_0339_),
    .B(_0338_),
    .A(\cpu0.a_reg[3] ));
 sg13g2_and2_1 _0923_ (.A(\cpu0.a_reg[3] ),
    .B(_0338_),
    .X(_0340_));
 sg13g2_xor2_1 _0924_ (.B(_0338_),
    .A(\cpu0.a_reg[3] ),
    .X(_0341_));
 sg13g2_a21oi_1 _0925_ (.A1(_0302_),
    .A2(_0306_),
    .Y(_0342_),
    .B1(_0307_));
 sg13g2_xnor2_1 _0926_ (.Y(_0343_),
    .A(_0341_),
    .B(_0342_));
 sg13g2_a221oi_1 _0927_ (.B2(_0343_),
    .C1(_0232_),
    .B1(_0259_),
    .A1(\cpu0.a_reg[3] ),
    .Y(_0344_),
    .A2(_0254_));
 sg13g2_o21ai_1 _0928_ (.B1(_0247_),
    .Y(_0345_),
    .A1(\cpu0.ir[3] ),
    .A2(_0233_));
 sg13g2_mux2_1 _0929_ (.A0(\cpu0.ram[12][3] ),
    .A1(\cpu0.ram[13][3] ),
    .S(net171),
    .X(_0346_));
 sg13g2_o21ai_1 _0930_ (.B1(net164),
    .Y(_0347_),
    .A1(net172),
    .A2(_0190_));
 sg13g2_a21oi_1 _0931_ (.A1(net172),
    .A2(\cpu0.ram[15][3] ),
    .Y(_0348_),
    .B1(_0347_));
 sg13g2_o21ai_1 _0932_ (.B1(net158),
    .Y(_0349_),
    .A1(net163),
    .A2(_0346_));
 sg13g2_nor2b_1 _0933_ (.A(net177),
    .B_N(\cpu0.ram[8][3] ),
    .Y(_0350_));
 sg13g2_a21oi_1 _0934_ (.A1(net174),
    .A2(\cpu0.ram[9][3] ),
    .Y(_0351_),
    .B1(_0350_));
 sg13g2_nand2b_1 _0935_ (.Y(_0352_),
    .B(\cpu0.ram[10][3] ),
    .A_N(net174));
 sg13g2_a21oi_1 _0936_ (.A1(net174),
    .A2(\cpu0.ram[11][3] ),
    .Y(_0353_),
    .B1(net152));
 sg13g2_a221oi_1 _0937_ (.B2(_0353_),
    .C1(net158),
    .B1(_0352_),
    .A1(net152),
    .Y(_0354_),
    .A2(_0351_));
 sg13g2_o21ai_1 _0938_ (.B1(net156),
    .Y(_0355_),
    .A1(_0348_),
    .A2(_0349_));
 sg13g2_nor2_1 _0939_ (.A(_0354_),
    .B(_0355_),
    .Y(_0356_));
 sg13g2_mux4_1 _0940_ (.S0(net170),
    .A0(\cpu0.ram[0][3] ),
    .A1(\cpu0.ram[1][3] ),
    .A2(\cpu0.ram[2][3] ),
    .A3(\cpu0.ram[3][3] ),
    .S1(net162),
    .X(_0357_));
 sg13g2_a21oi_1 _0941_ (.A1(net167),
    .A2(\cpu0.ram[5][3] ),
    .Y(_0358_),
    .B1(net160));
 sg13g2_o21ai_1 _0942_ (.B1(_0358_),
    .Y(_0359_),
    .A1(net166),
    .A2(_0189_));
 sg13g2_nor2b_1 _0943_ (.A(net166),
    .B_N(\cpu0.ram[6][3] ),
    .Y(_0360_));
 sg13g2_a21oi_1 _0944_ (.A1(net166),
    .A2(\cpu0.ram[7][3] ),
    .Y(_0361_),
    .B1(_0360_));
 sg13g2_a21oi_1 _0945_ (.A1(net160),
    .A2(_0361_),
    .Y(_0362_),
    .B1(_0184_));
 sg13g2_a221oi_1 _0946_ (.B2(_0362_),
    .C1(net155),
    .B1(_0359_),
    .A1(_0184_),
    .Y(_0363_),
    .A2(_0357_));
 sg13g2_nor2_1 _0947_ (.A(_0356_),
    .B(_0363_),
    .Y(_0364_));
 sg13g2_a21oi_1 _0948_ (.A1(_0248_),
    .A2(_0364_),
    .Y(_0365_),
    .B1(_0212_));
 sg13g2_o21ai_1 _0949_ (.B1(_0365_),
    .Y(_0366_),
    .A1(_0344_),
    .A2(_0345_));
 sg13g2_o21ai_1 _0950_ (.B1(_0366_),
    .Y(_0367_),
    .A1(\cpu0.pc[3] ),
    .A2(_0213_));
 sg13g2_nor2_1 _0951_ (.A(net4),
    .B(net147),
    .Y(_0368_));
 sg13g2_a21oi_2 _0952_ (.B1(_0368_),
    .Y(_0369_),
    .A2(_0367_),
    .A1(net147));
 sg13g2_mux2_1 _0953_ (.A0(net128),
    .A1(net329),
    .S(_0210_),
    .X(_0007_));
 sg13g2_nor2_1 _0954_ (.A(net5),
    .B(net147),
    .Y(_0370_));
 sg13g2_nor2b_1 _0955_ (.A(_0308_),
    .B_N(_0341_),
    .Y(_0371_));
 sg13g2_a221oi_1 _0956_ (.B2(_0302_),
    .C1(_0340_),
    .B1(_0371_),
    .A1(_0307_),
    .Y(_0372_),
    .A2(_0339_));
 sg13g2_o21ai_1 _0957_ (.B1(_0270_),
    .Y(_0373_),
    .A1(\cpu0.b_reg[3] ),
    .A2(_0336_));
 sg13g2_xor2_1 _0958_ (.B(_0373_),
    .A(\cpu0.b_reg[4] ),
    .X(_0374_));
 sg13g2_nand2_1 _0959_ (.Y(_0375_),
    .A(\cpu0.a_reg[4] ),
    .B(_0374_));
 sg13g2_xor2_1 _0960_ (.B(_0374_),
    .A(\cpu0.a_reg[4] ),
    .X(_0376_));
 sg13g2_nand2b_1 _0961_ (.Y(_0377_),
    .B(_0376_),
    .A_N(_0372_));
 sg13g2_xnor2_1 _0962_ (.Y(_0378_),
    .A(_0372_),
    .B(_0376_));
 sg13g2_a221oi_1 _0963_ (.B2(_0378_),
    .C1(_0248_),
    .B1(net144),
    .A1(\cpu0.a_reg[4] ),
    .Y(_0379_),
    .A2(_0254_));
 sg13g2_o21ai_1 _0964_ (.B1(net152),
    .Y(_0380_),
    .A1(net172),
    .A2(\cpu0.ram[12][4] ));
 sg13g2_a21oi_1 _0965_ (.A1(net172),
    .A2(_0191_),
    .Y(_0381_),
    .B1(_0380_));
 sg13g2_nor2b_1 _0966_ (.A(\cpu0.ram[15][4] ),
    .B_N(net173),
    .Y(_0382_));
 sg13g2_o21ai_1 _0967_ (.B1(net164),
    .Y(_0383_),
    .A1(net173),
    .A2(\cpu0.ram[14][4] ));
 sg13g2_o21ai_1 _0968_ (.B1(net158),
    .Y(_0384_),
    .A1(_0382_),
    .A2(_0383_));
 sg13g2_mux4_1 _0969_ (.S0(net176),
    .A0(\cpu0.ram[8][4] ),
    .A1(\cpu0.ram[9][4] ),
    .A2(\cpu0.ram[10][4] ),
    .A3(\cpu0.ram[11][4] ),
    .S1(net165),
    .X(_0385_));
 sg13g2_nor2_1 _0970_ (.A(net159),
    .B(_0385_),
    .Y(_0386_));
 sg13g2_o21ai_1 _0971_ (.B1(net156),
    .Y(_0387_),
    .A1(_0381_),
    .A2(_0384_));
 sg13g2_mux4_1 _0972_ (.S0(net170),
    .A0(\cpu0.ram[0][4] ),
    .A1(\cpu0.ram[1][4] ),
    .A2(\cpu0.ram[2][4] ),
    .A3(\cpu0.ram[3][4] ),
    .S1(net161),
    .X(_0388_));
 sg13g2_nor2_1 _0973_ (.A(net157),
    .B(_0388_),
    .Y(_0389_));
 sg13g2_mux2_1 _0974_ (.A0(\cpu0.ram[4][4] ),
    .A1(\cpu0.ram[5][4] ),
    .S(net168),
    .X(_0390_));
 sg13g2_nor2b_1 _0975_ (.A(\cpu0.ram[7][4] ),
    .B_N(net168),
    .Y(_0391_));
 sg13g2_o21ai_1 _0976_ (.B1(net160),
    .Y(_0392_),
    .A1(net168),
    .A2(\cpu0.ram[6][4] ));
 sg13g2_o21ai_1 _0977_ (.B1(net157),
    .Y(_0393_),
    .A1(_0391_),
    .A2(_0392_));
 sg13g2_a21oi_1 _0978_ (.A1(net151),
    .A2(_0390_),
    .Y(_0394_),
    .B1(_0393_));
 sg13g2_nor3_1 _0979_ (.A(net156),
    .B(_0389_),
    .C(_0394_),
    .Y(_0395_));
 sg13g2_nor2_1 _0980_ (.A(_0247_),
    .B(_0395_),
    .Y(_0396_));
 sg13g2_o21ai_1 _0981_ (.B1(_0396_),
    .Y(_0397_),
    .A1(_0386_),
    .A2(_0387_));
 sg13g2_nand2b_2 _0982_ (.Y(_0398_),
    .B(_0397_),
    .A_N(_0379_));
 sg13g2_a21oi_2 _0983_ (.B1(_0370_),
    .Y(_0399_),
    .A2(_0398_),
    .A1(net146));
 sg13g2_mux2_1 _0984_ (.A0(net130),
    .A1(net422),
    .S(_0210_),
    .X(_0008_));
 sg13g2_or3_1 _0985_ (.A(\cpu0.b_reg[4] ),
    .B(\cpu0.b_reg[3] ),
    .C(_0336_),
    .X(_0400_));
 sg13g2_nand2_1 _0986_ (.Y(_0401_),
    .A(_0270_),
    .B(_0400_));
 sg13g2_xor2_1 _0987_ (.B(_0401_),
    .A(\cpu0.b_reg[5] ),
    .X(_0402_));
 sg13g2_nand2_1 _0988_ (.Y(_0403_),
    .A(\cpu0.a_reg[5] ),
    .B(_0402_));
 sg13g2_xor2_1 _0989_ (.B(_0402_),
    .A(\cpu0.a_reg[5] ),
    .X(_0404_));
 sg13g2_inv_1 _0990_ (.Y(_0405_),
    .A(_0404_));
 sg13g2_nand3_1 _0991_ (.B(_0377_),
    .C(_0405_),
    .A(_0375_),
    .Y(_0406_));
 sg13g2_and2_1 _0992_ (.A(_0376_),
    .B(_0404_),
    .X(_0407_));
 sg13g2_nor2b_1 _0993_ (.A(_0372_),
    .B_N(_0407_),
    .Y(_0408_));
 sg13g2_o21ai_1 _0994_ (.B1(net144),
    .Y(_0409_),
    .A1(_0375_),
    .A2(_0405_));
 sg13g2_nor2_1 _0995_ (.A(_0408_),
    .B(_0409_),
    .Y(_0410_));
 sg13g2_a221oi_1 _0996_ (.B2(_0410_),
    .C1(_0248_),
    .B1(_0406_),
    .A1(\cpu0.a_reg[5] ),
    .Y(_0411_),
    .A2(_0254_));
 sg13g2_mux4_1 _0997_ (.S0(net170),
    .A0(\cpu0.ram[0][5] ),
    .A1(\cpu0.ram[1][5] ),
    .A2(\cpu0.ram[2][5] ),
    .A3(\cpu0.ram[3][5] ),
    .S1(net162),
    .X(_0412_));
 sg13g2_and2_1 _0998_ (.A(_0184_),
    .B(_0412_),
    .X(_0413_));
 sg13g2_mux4_1 _0999_ (.S0(net166),
    .A0(\cpu0.ram[4][5] ),
    .A1(\cpu0.ram[5][5] ),
    .A2(\cpu0.ram[6][5] ),
    .A3(\cpu0.ram[7][5] ),
    .S1(net160),
    .X(_0414_));
 sg13g2_a21oi_1 _1000_ (.A1(net159),
    .A2(_0414_),
    .Y(_0415_),
    .B1(_0413_));
 sg13g2_mux2_1 _1001_ (.A0(\cpu0.ram[8][5] ),
    .A1(\cpu0.ram[9][5] ),
    .S(net168),
    .X(_0416_));
 sg13g2_nand2_1 _1002_ (.Y(_0417_),
    .A(net151),
    .B(_0416_));
 sg13g2_o21ai_1 _1003_ (.B1(net163),
    .Y(_0418_),
    .A1(net171),
    .A2(\cpu0.ram[10][5] ));
 sg13g2_a21oi_1 _1004_ (.A1(net171),
    .A2(_0192_),
    .Y(_0419_),
    .B1(_0418_));
 sg13g2_nor2_1 _1005_ (.A(net157),
    .B(_0419_),
    .Y(_0420_));
 sg13g2_o21ai_1 _1006_ (.B1(net151),
    .Y(_0421_),
    .A1(net171),
    .A2(\cpu0.ram[12][5] ));
 sg13g2_a21oi_1 _1007_ (.A1(net171),
    .A2(_0193_),
    .Y(_0422_),
    .B1(_0421_));
 sg13g2_nor2b_1 _1008_ (.A(\cpu0.ram[15][5] ),
    .B_N(net171),
    .Y(_0423_));
 sg13g2_o21ai_1 _1009_ (.B1(net163),
    .Y(_0424_),
    .A1(net171),
    .A2(\cpu0.ram[14][5] ));
 sg13g2_o21ai_1 _1010_ (.B1(net157),
    .Y(_0425_),
    .A1(_0423_),
    .A2(_0424_));
 sg13g2_o21ai_1 _1011_ (.B1(net155),
    .Y(_0426_),
    .A1(_0422_),
    .A2(_0425_));
 sg13g2_a21oi_1 _1012_ (.A1(_0417_),
    .A2(_0420_),
    .Y(_0427_),
    .B1(_0426_));
 sg13g2_nor2_1 _1013_ (.A(_0247_),
    .B(_0427_),
    .Y(_0428_));
 sg13g2_o21ai_1 _1014_ (.B1(_0428_),
    .Y(_0429_),
    .A1(net155),
    .A2(_0415_));
 sg13g2_nand2b_2 _1015_ (.Y(_0430_),
    .B(_0429_),
    .A_N(_0411_));
 sg13g2_nor2_1 _1016_ (.A(net6),
    .B(net146),
    .Y(_0431_));
 sg13g2_a21oi_2 _1017_ (.B1(_0431_),
    .Y(_0432_),
    .A2(_0430_),
    .A1(net146));
 sg13g2_mux2_1 _1018_ (.A0(net126),
    .A1(net398),
    .S(_0210_),
    .X(_0009_));
 sg13g2_o21ai_1 _1019_ (.B1(_0270_),
    .Y(_0433_),
    .A1(\cpu0.b_reg[5] ),
    .A2(_0400_));
 sg13g2_xor2_1 _1020_ (.B(_0433_),
    .A(\cpu0.b_reg[6] ),
    .X(_0434_));
 sg13g2_nand2_1 _1021_ (.Y(_0435_),
    .A(\cpu0.a_reg[6] ),
    .B(_0434_));
 sg13g2_xor2_1 _1022_ (.B(_0434_),
    .A(net294),
    .X(_0436_));
 sg13g2_o21ai_1 _1023_ (.B1(_0403_),
    .Y(_0437_),
    .A1(_0375_),
    .A2(_0405_));
 sg13g2_o21ai_1 _1024_ (.B1(_0436_),
    .Y(_0438_),
    .A1(_0408_),
    .A2(_0437_));
 sg13g2_nor3_1 _1025_ (.A(_0408_),
    .B(_0436_),
    .C(_0437_),
    .Y(_0439_));
 sg13g2_nor2b_1 _1026_ (.A(_0439_),
    .B_N(net144),
    .Y(_0440_));
 sg13g2_a221oi_1 _1027_ (.B2(_0440_),
    .C1(_0248_),
    .B1(_0438_),
    .A1(\cpu0.a_reg[6] ),
    .Y(_0441_),
    .A2(_0254_));
 sg13g2_nand2b_1 _1028_ (.Y(_0442_),
    .B(net176),
    .A_N(\cpu0.ram[11][6] ));
 sg13g2_mux2_1 _1029_ (.A0(\cpu0.ram[8][6] ),
    .A1(\cpu0.ram[9][6] ),
    .S(net176),
    .X(_0443_));
 sg13g2_o21ai_1 _1030_ (.B1(_0442_),
    .Y(_0444_),
    .A1(net177),
    .A2(\cpu0.ram[10][6] ));
 sg13g2_a21oi_1 _1031_ (.A1(net165),
    .A2(_0444_),
    .Y(_0445_),
    .B1(net159));
 sg13g2_o21ai_1 _1032_ (.B1(_0445_),
    .Y(_0446_),
    .A1(net163),
    .A2(_0443_));
 sg13g2_o21ai_1 _1033_ (.B1(net151),
    .Y(_0447_),
    .A1(net174),
    .A2(_0194_));
 sg13g2_a21oi_1 _1034_ (.A1(net174),
    .A2(\cpu0.ram[13][6] ),
    .Y(_0448_),
    .B1(_0447_));
 sg13g2_mux2_1 _1035_ (.A0(\cpu0.ram[14][6] ),
    .A1(\cpu0.ram[15][6] ),
    .S(net174),
    .X(_0449_));
 sg13g2_o21ai_1 _1036_ (.B1(net158),
    .Y(_0450_),
    .A1(net152),
    .A2(_0449_));
 sg13g2_o21ai_1 _1037_ (.B1(_0446_),
    .Y(_0451_),
    .A1(_0448_),
    .A2(_0450_));
 sg13g2_mux4_1 _1038_ (.S0(_0000_),
    .A0(\cpu0.ram[0][6] ),
    .A1(\cpu0.ram[1][6] ),
    .A2(\cpu0.ram[2][6] ),
    .A3(\cpu0.ram[3][6] ),
    .S1(net161),
    .X(_0452_));
 sg13g2_mux2_1 _1039_ (.A0(\cpu0.ram[4][6] ),
    .A1(\cpu0.ram[5][6] ),
    .S(net168),
    .X(_0453_));
 sg13g2_nor2b_1 _1040_ (.A(\cpu0.ram[7][6] ),
    .B_N(net169),
    .Y(_0454_));
 sg13g2_o21ai_1 _1041_ (.B1(net161),
    .Y(_0455_),
    .A1(net169),
    .A2(\cpu0.ram[6][6] ));
 sg13g2_o21ai_1 _1042_ (.B1(net157),
    .Y(_0456_),
    .A1(_0454_),
    .A2(_0455_));
 sg13g2_a21oi_1 _1043_ (.A1(net151),
    .A2(_0453_),
    .Y(_0457_),
    .B1(_0456_));
 sg13g2_nor2_1 _1044_ (.A(net156),
    .B(_0457_),
    .Y(_0458_));
 sg13g2_o21ai_1 _1045_ (.B1(_0458_),
    .Y(_0459_),
    .A1(net157),
    .A2(_0452_));
 sg13g2_a21oi_1 _1046_ (.A1(net156),
    .A2(_0451_),
    .Y(_0460_),
    .B1(_0247_));
 sg13g2_a21o_2 _1047_ (.A2(_0460_),
    .A1(_0459_),
    .B1(_0441_),
    .X(_0461_));
 sg13g2_nor2_1 _1048_ (.A(net7),
    .B(net148),
    .Y(_0462_));
 sg13g2_a21oi_2 _1049_ (.B1(_0462_),
    .Y(_0463_),
    .A2(_0461_),
    .A1(net146));
 sg13g2_mux2_1 _1050_ (.A0(net124),
    .A1(net342),
    .S(_0210_),
    .X(_0010_));
 sg13g2_nor2_1 _1051_ (.A(net8),
    .B(net148),
    .Y(_0464_));
 sg13g2_nand2_1 _1052_ (.Y(_0465_),
    .A(\cpu0.b_reg[6] ),
    .B(_0270_));
 sg13g2_nand2_1 _1053_ (.Y(_0466_),
    .A(_0433_),
    .B(_0465_));
 sg13g2_xnor2_1 _1054_ (.Y(_0467_),
    .A(\cpu0.b_reg[7] ),
    .B(_0466_));
 sg13g2_nor2_1 _1055_ (.A(\cpu0.a_reg[7] ),
    .B(_0467_),
    .Y(_0468_));
 sg13g2_xnor2_1 _1056_ (.Y(_0469_),
    .A(net424),
    .B(_0467_));
 sg13g2_nand3_1 _1057_ (.B(_0438_),
    .C(_0469_),
    .A(_0435_),
    .Y(_0470_));
 sg13g2_a21o_1 _1058_ (.A2(_0438_),
    .A1(_0435_),
    .B1(_0469_),
    .X(_0471_));
 sg13g2_nand3_1 _1059_ (.B(_0470_),
    .C(_0471_),
    .A(net144),
    .Y(_0472_));
 sg13g2_a21oi_1 _1060_ (.A1(net424),
    .A2(_0254_),
    .Y(_0473_),
    .B1(_0248_));
 sg13g2_mux4_1 _1061_ (.S0(net170),
    .A0(\cpu0.ram[0][7] ),
    .A1(\cpu0.ram[1][7] ),
    .A2(\cpu0.ram[2][7] ),
    .A3(\cpu0.ram[3][7] ),
    .S1(net162),
    .X(_0474_));
 sg13g2_nand2b_1 _1062_ (.Y(_0475_),
    .B(_0184_),
    .A_N(_0474_));
 sg13g2_mux2_1 _1063_ (.A0(\cpu0.ram[4][7] ),
    .A1(\cpu0.ram[5][7] ),
    .S(net167),
    .X(_0476_));
 sg13g2_nor2b_1 _1064_ (.A(\cpu0.ram[7][7] ),
    .B_N(net167),
    .Y(_0477_));
 sg13g2_o21ai_1 _1065_ (.B1(net160),
    .Y(_0478_),
    .A1(net167),
    .A2(\cpu0.ram[6][7] ));
 sg13g2_o21ai_1 _1066_ (.B1(net157),
    .Y(_0479_),
    .A1(_0477_),
    .A2(_0478_));
 sg13g2_a21oi_1 _1067_ (.A1(net151),
    .A2(_0476_),
    .Y(_0480_),
    .B1(_0479_));
 sg13g2_nor2_1 _1068_ (.A(net155),
    .B(_0480_),
    .Y(_0481_));
 sg13g2_mux4_1 _1069_ (.S0(net176),
    .A0(\cpu0.ram[8][7] ),
    .A1(\cpu0.ram[9][7] ),
    .A2(\cpu0.ram[10][7] ),
    .A3(\cpu0.ram[11][7] ),
    .S1(net165),
    .X(_0482_));
 sg13g2_mux4_1 _1070_ (.S0(net171),
    .A0(\cpu0.ram[12][7] ),
    .A1(\cpu0.ram[13][7] ),
    .A2(\cpu0.ram[14][7] ),
    .A3(\cpu0.ram[15][7] ),
    .S1(net163),
    .X(_0483_));
 sg13g2_mux2_1 _1071_ (.A0(_0482_),
    .A1(_0483_),
    .S(net159),
    .X(_0484_));
 sg13g2_a221oi_1 _1072_ (.B2(net155),
    .C1(_0247_),
    .B1(_0484_),
    .A1(_0475_),
    .Y(_0485_),
    .A2(_0481_));
 sg13g2_a21o_2 _1073_ (.A2(_0473_),
    .A1(_0472_),
    .B1(_0485_),
    .X(_0486_));
 sg13g2_a21oi_2 _1074_ (.B1(_0464_),
    .Y(_0487_),
    .A2(_0486_),
    .A1(net148));
 sg13g2_mux2_1 _1075_ (.A0(net122),
    .A1(net390),
    .S(_0210_),
    .X(_0011_));
 sg13g2_a21oi_1 _1076_ (.A1(\cpu0.ir[7] ),
    .A2(\cpu0.ir[6] ),
    .Y(_0488_),
    .B1(_0200_));
 sg13g2_nor2_1 _1077_ (.A(_0239_),
    .B(_0488_),
    .Y(_0489_));
 sg13g2_o21ai_1 _1078_ (.B1(_0213_),
    .Y(_0490_),
    .A1(_0231_),
    .A2(_0489_));
 sg13g2_o21ai_1 _1079_ (.B1(net178),
    .Y(_0491_),
    .A1(net443),
    .A2(net141));
 sg13g2_a21oi_1 _1080_ (.A1(_0263_),
    .A2(net141),
    .Y(_0012_),
    .B1(_0491_));
 sg13g2_o21ai_1 _1081_ (.B1(net178),
    .Y(_0492_),
    .A1(net440),
    .A2(net141));
 sg13g2_a21oi_1 _1082_ (.A1(_0299_),
    .A2(net141),
    .Y(_0013_),
    .B1(_0492_));
 sg13g2_o21ai_1 _1083_ (.B1(net178),
    .Y(_0493_),
    .A1(net438),
    .A2(net141));
 sg13g2_a21oi_1 _1084_ (.A1(_0333_),
    .A2(net141),
    .Y(_0014_),
    .B1(_0493_));
 sg13g2_o21ai_1 _1085_ (.B1(net178),
    .Y(_0494_),
    .A1(net439),
    .A2(net142));
 sg13g2_a21oi_1 _1086_ (.A1(_0367_),
    .A2(net142),
    .Y(_0015_),
    .B1(_0494_));
 sg13g2_nand2b_2 _1087_ (.Y(_0495_),
    .B(_0208_),
    .A_N(_0207_));
 sg13g2_nor2b_1 _1088_ (.A(_0204_),
    .B_N(_0202_),
    .Y(_0496_));
 sg13g2_nand2b_1 _1089_ (.Y(_0497_),
    .B(_0496_),
    .A_N(_0205_));
 sg13g2_or2_1 _1090_ (.X(_0498_),
    .B(_0497_),
    .A(_0495_));
 sg13g2_mux2_1 _1091_ (.A0(net136),
    .A1(net363),
    .S(_0498_),
    .X(_0016_));
 sg13g2_mux2_1 _1092_ (.A0(net134),
    .A1(net386),
    .S(_0498_),
    .X(_0017_));
 sg13g2_mux2_1 _1093_ (.A0(net132),
    .A1(net349),
    .S(_0498_),
    .X(_0018_));
 sg13g2_mux2_1 _1094_ (.A0(net128),
    .A1(net346),
    .S(_0498_),
    .X(_0019_));
 sg13g2_mux2_1 _1095_ (.A0(net130),
    .A1(net415),
    .S(_0498_),
    .X(_0020_));
 sg13g2_mux2_1 _1096_ (.A0(net126),
    .A1(net356),
    .S(_0498_),
    .X(_0021_));
 sg13g2_mux2_1 _1097_ (.A0(net124),
    .A1(net409),
    .S(_0498_),
    .X(_0022_));
 sg13g2_mux2_1 _1098_ (.A0(net122),
    .A1(net378),
    .S(_0498_),
    .X(_0023_));
 sg13g2_nand2_1 _1099_ (.Y(_0024_),
    .A(_0211_),
    .B(_0242_));
 sg13g2_o21ai_1 _1100_ (.B1(_0231_),
    .Y(_0025_),
    .A1(_0197_),
    .A2(_0214_));
 sg13g2_nand3_1 _1101_ (.B(_0204_),
    .C(_0205_),
    .A(_0202_),
    .Y(_0499_));
 sg13g2_or2_1 _1102_ (.X(_0500_),
    .B(_0499_),
    .A(_0495_));
 sg13g2_mux2_1 _1103_ (.A0(net137),
    .A1(net338),
    .S(net140),
    .X(_0026_));
 sg13g2_mux2_1 _1104_ (.A0(net135),
    .A1(net403),
    .S(net140),
    .X(_0027_));
 sg13g2_nor2_1 _1105_ (.A(net133),
    .B(net140),
    .Y(_0501_));
 sg13g2_a21oi_1 _1106_ (.A1(_0188_),
    .A2(net140),
    .Y(_0028_),
    .B1(_0501_));
 sg13g2_nor2_1 _1107_ (.A(net129),
    .B(net140),
    .Y(_0502_));
 sg13g2_a21oi_1 _1108_ (.A1(_0190_),
    .A2(net140),
    .Y(_0029_),
    .B1(_0502_));
 sg13g2_mux2_1 _1109_ (.A0(net131),
    .A1(net365),
    .S(_0500_),
    .X(_0030_));
 sg13g2_mux2_1 _1110_ (.A0(net127),
    .A1(net379),
    .S(net140),
    .X(_0031_));
 sg13g2_mux2_1 _1111_ (.A0(net125),
    .A1(net324),
    .S(_0500_),
    .X(_0032_));
 sg13g2_mux2_1 _1112_ (.A0(net123),
    .A1(net350),
    .S(net140),
    .X(_0033_));
 sg13g2_a21oi_1 _1113_ (.A1(net432),
    .A2(\cpu0.step[2] ),
    .Y(_0503_),
    .B1(_0181_));
 sg13g2_nor2_1 _1114_ (.A(_0182_),
    .B(net433),
    .Y(_0034_));
 sg13g2_nor2_2 _1115_ (.A(_0207_),
    .B(_0208_),
    .Y(_0504_));
 sg13g2_nand2b_2 _1116_ (.Y(_0505_),
    .B(_0504_),
    .A_N(_0206_));
 sg13g2_mux2_1 _1117_ (.A0(net136),
    .A1(net407),
    .S(_0505_),
    .X(_0035_));
 sg13g2_mux2_1 _1118_ (.A0(net134),
    .A1(net298),
    .S(_0505_),
    .X(_0036_));
 sg13g2_mux2_1 _1119_ (.A0(net132),
    .A1(net326),
    .S(_0505_),
    .X(_0037_));
 sg13g2_mux2_1 _1120_ (.A0(net128),
    .A1(net371),
    .S(_0505_),
    .X(_0038_));
 sg13g2_mux2_1 _1121_ (.A0(net130),
    .A1(net408),
    .S(_0505_),
    .X(_0039_));
 sg13g2_mux2_1 _1122_ (.A0(net126),
    .A1(net362),
    .S(_0505_),
    .X(_0040_));
 sg13g2_mux2_1 _1123_ (.A0(net124),
    .A1(net396),
    .S(_0505_),
    .X(_0041_));
 sg13g2_mux2_1 _1124_ (.A0(net122),
    .A1(net323),
    .S(_0505_),
    .X(_0042_));
 sg13g2_nand2_2 _1125_ (.Y(_0506_),
    .A(_0207_),
    .B(_0208_));
 sg13g2_or2_1 _1126_ (.X(_0507_),
    .B(_0506_),
    .A(_0497_));
 sg13g2_mux2_1 _1127_ (.A0(net136),
    .A1(net339),
    .S(_0507_),
    .X(_0043_));
 sg13g2_mux2_1 _1128_ (.A0(net134),
    .A1(net315),
    .S(_0507_),
    .X(_0044_));
 sg13g2_mux2_1 _1129_ (.A0(net132),
    .A1(net367),
    .S(_0507_),
    .X(_0045_));
 sg13g2_mux2_1 _1130_ (.A0(net128),
    .A1(net316),
    .S(_0507_),
    .X(_0046_));
 sg13g2_mux2_1 _1131_ (.A0(net130),
    .A1(net401),
    .S(_0507_),
    .X(_0047_));
 sg13g2_mux2_1 _1132_ (.A0(net126),
    .A1(net388),
    .S(_0507_),
    .X(_0048_));
 sg13g2_mux2_1 _1133_ (.A0(net124),
    .A1(net314),
    .S(_0507_),
    .X(_0049_));
 sg13g2_mux2_1 _1134_ (.A0(net122),
    .A1(net325),
    .S(_0507_),
    .X(_0050_));
 sg13g2_or2_1 _1135_ (.X(_0508_),
    .B(_0497_),
    .A(_0209_));
 sg13g2_mux2_1 _1136_ (.A0(net136),
    .A1(net344),
    .S(_0508_),
    .X(_0051_));
 sg13g2_mux2_1 _1137_ (.A0(net134),
    .A1(net383),
    .S(_0508_),
    .X(_0052_));
 sg13g2_mux2_1 _1138_ (.A0(net132),
    .A1(net427),
    .S(_0508_),
    .X(_0053_));
 sg13g2_mux2_1 _1139_ (.A0(net128),
    .A1(net394),
    .S(_0508_),
    .X(_0054_));
 sg13g2_mux2_1 _1140_ (.A0(net130),
    .A1(net413),
    .S(_0508_),
    .X(_0055_));
 sg13g2_mux2_1 _1141_ (.A0(net126),
    .A1(net307),
    .S(_0508_),
    .X(_0056_));
 sg13g2_mux2_1 _1142_ (.A0(net124),
    .A1(net423),
    .S(_0508_),
    .X(_0057_));
 sg13g2_mux2_1 _1143_ (.A0(net122),
    .A1(net360),
    .S(_0508_),
    .X(_0058_));
 sg13g2_or2_1 _1144_ (.X(_0509_),
    .B(_0506_),
    .A(_0499_));
 sg13g2_mux2_1 _1145_ (.A0(net137),
    .A1(net406),
    .S(net139),
    .X(_0059_));
 sg13g2_nor2_1 _1146_ (.A(net135),
    .B(net139),
    .Y(_0510_));
 sg13g2_a21oi_1 _1147_ (.A1(_0186_),
    .A2(net139),
    .Y(_0060_),
    .B1(_0510_));
 sg13g2_mux2_1 _1148_ (.A0(net133),
    .A1(net321),
    .S(net139),
    .X(_0061_));
 sg13g2_mux2_1 _1149_ (.A0(net129),
    .A1(net376),
    .S(net139),
    .X(_0062_));
 sg13g2_mux2_1 _1150_ (.A0(net131),
    .A1(net353),
    .S(net139),
    .X(_0063_));
 sg13g2_mux2_1 _1151_ (.A0(net127),
    .A1(net359),
    .S(net139),
    .X(_0064_));
 sg13g2_mux2_1 _1152_ (.A0(net125),
    .A1(net412),
    .S(_0509_),
    .X(_0065_));
 sg13g2_mux2_1 _1153_ (.A0(net123),
    .A1(net421),
    .S(net139),
    .X(_0066_));
 sg13g2_nor2_2 _1154_ (.A(_0246_),
    .B(net144),
    .Y(_0511_));
 sg13g2_nor3_1 _1155_ (.A(_0196_),
    .B(_0228_),
    .C(_0231_),
    .Y(_0512_));
 sg13g2_nor3_2 _1156_ (.A(_0246_),
    .B(net144),
    .C(_0512_),
    .Y(_0513_));
 sg13g2_and2_1 _1157_ (.A(net180),
    .B(_0513_),
    .X(_0514_));
 sg13g2_nand2_1 _1158_ (.Y(_0515_),
    .A(net285),
    .B(_0514_));
 sg13g2_o21ai_1 _1159_ (.B1(_0515_),
    .Y(_0067_),
    .A1(_0263_),
    .A2(_0513_));
 sg13g2_nand2_1 _1160_ (.Y(_0516_),
    .A(net300),
    .B(_0514_));
 sg13g2_o21ai_1 _1161_ (.B1(_0516_),
    .Y(_0068_),
    .A1(_0299_),
    .A2(_0513_));
 sg13g2_nand2_1 _1162_ (.Y(_0517_),
    .A(net351),
    .B(_0514_));
 sg13g2_o21ai_1 _1163_ (.B1(_0517_),
    .Y(_0069_),
    .A1(_0333_),
    .A2(_0513_));
 sg13g2_nand2_1 _1164_ (.Y(_0518_),
    .A(net425),
    .B(_0514_));
 sg13g2_o21ai_1 _1165_ (.B1(_0518_),
    .Y(_0070_),
    .A1(_0367_),
    .A2(_0513_));
 sg13g2_nand2_1 _1166_ (.Y(_0519_),
    .A(net295),
    .B(_0514_));
 sg13g2_o21ai_1 _1167_ (.B1(_0519_),
    .Y(_0071_),
    .A1(_0398_),
    .A2(_0511_));
 sg13g2_nand2_1 _1168_ (.Y(_0520_),
    .A(net286),
    .B(_0514_));
 sg13g2_o21ai_1 _1169_ (.B1(_0520_),
    .Y(_0072_),
    .A1(_0430_),
    .A2(_0511_));
 sg13g2_nand2_1 _1170_ (.Y(_0521_),
    .A(net294),
    .B(_0514_));
 sg13g2_o21ai_1 _1171_ (.B1(_0521_),
    .Y(_0073_),
    .A1(_0461_),
    .A2(_0511_));
 sg13g2_nand2_1 _1172_ (.Y(_0522_),
    .A(net424),
    .B(_0514_));
 sg13g2_o21ai_1 _1173_ (.B1(_0522_),
    .Y(_0074_),
    .A1(_0486_),
    .A2(_0511_));
 sg13g2_nor2_2 _1174_ (.A(_0182_),
    .B(_0243_),
    .Y(_0523_));
 sg13g2_nand2_1 _1175_ (.Y(_0524_),
    .A(net267),
    .B(_0523_));
 sg13g2_o21ai_1 _1176_ (.B1(_0524_),
    .Y(_0075_),
    .A1(net149),
    .A2(_0263_));
 sg13g2_nand2_1 _1177_ (.Y(_0525_),
    .A(net266),
    .B(_0523_));
 sg13g2_o21ai_1 _1178_ (.B1(_0525_),
    .Y(_0076_),
    .A1(net149),
    .A2(_0299_));
 sg13g2_nand2_1 _1179_ (.Y(_0526_),
    .A(net274),
    .B(_0523_));
 sg13g2_o21ai_1 _1180_ (.B1(_0526_),
    .Y(_0077_),
    .A1(net149),
    .A2(_0333_));
 sg13g2_nand2_1 _1181_ (.Y(_0527_),
    .A(net269),
    .B(_0523_));
 sg13g2_o21ai_1 _1182_ (.B1(_0527_),
    .Y(_0078_),
    .A1(net149),
    .A2(_0367_));
 sg13g2_nand2_1 _1183_ (.Y(_0528_),
    .A(net434),
    .B(_0523_));
 sg13g2_o21ai_1 _1184_ (.B1(_0528_),
    .Y(_0079_),
    .A1(net149),
    .A2(_0398_));
 sg13g2_nand2_1 _1185_ (.Y(_0529_),
    .A(net271),
    .B(_0523_));
 sg13g2_o21ai_1 _1186_ (.B1(_0529_),
    .Y(_0080_),
    .A1(net149),
    .A2(_0430_));
 sg13g2_nand2_1 _1187_ (.Y(_0530_),
    .A(net429),
    .B(_0523_));
 sg13g2_o21ai_1 _1188_ (.B1(_0530_),
    .Y(_0081_),
    .A1(net150),
    .A2(_0461_));
 sg13g2_nand2_1 _1189_ (.Y(_0531_),
    .A(net435),
    .B(_0523_));
 sg13g2_o21ai_1 _1190_ (.B1(_0531_),
    .Y(_0082_),
    .A1(net150),
    .A2(_0486_));
 sg13g2_nand2_2 _1191_ (.Y(_0532_),
    .A(net179),
    .B(_0223_));
 sg13g2_xnor2_1 _1192_ (.Y(_0533_),
    .A(net444),
    .B(net150));
 sg13g2_nand3_1 _1193_ (.B(_0532_),
    .C(_0533_),
    .A(net178),
    .Y(_0534_));
 sg13g2_o21ai_1 _1194_ (.B1(_0534_),
    .Y(_0087_),
    .A1(_0263_),
    .A2(_0532_));
 sg13g2_nand3_1 _1195_ (.B(net444),
    .C(_0243_),
    .A(net442),
    .Y(_0535_));
 sg13g2_a21o_1 _1196_ (.A2(_0243_),
    .A1(net444),
    .B1(net442),
    .X(_0536_));
 sg13g2_nand4_1 _1197_ (.B(_0532_),
    .C(_0535_),
    .A(net178),
    .Y(_0537_),
    .D(_0536_));
 sg13g2_o21ai_1 _1198_ (.B1(_0537_),
    .Y(_0088_),
    .A1(_0299_),
    .A2(_0532_));
 sg13g2_nand3_1 _1199_ (.B(_0532_),
    .C(_0535_),
    .A(net441),
    .Y(_0538_));
 sg13g2_o21ai_1 _1200_ (.B1(_0538_),
    .Y(_0539_),
    .A1(net441),
    .A2(_0535_));
 sg13g2_nand2_1 _1201_ (.Y(_0540_),
    .A(net178),
    .B(_0539_));
 sg13g2_o21ai_1 _1202_ (.B1(_0540_),
    .Y(_0089_),
    .A1(_0333_),
    .A2(_0532_));
 sg13g2_nand4_1 _1203_ (.B(net442),
    .C(net444),
    .A(net441),
    .Y(_0541_),
    .D(_0243_));
 sg13g2_xnor2_1 _1204_ (.Y(_0542_),
    .A(net445),
    .B(_0541_));
 sg13g2_nand3_1 _1205_ (.B(_0532_),
    .C(_0542_),
    .A(net178),
    .Y(_0543_));
 sg13g2_o21ai_1 _1206_ (.B1(_0543_),
    .Y(_0090_),
    .A1(_0367_),
    .A2(_0532_));
 sg13g2_or2_1 _1207_ (.X(_0544_),
    .B(_0499_),
    .A(_0209_));
 sg13g2_mux2_1 _1208_ (.A0(net137),
    .A1(net340),
    .S(_0544_),
    .X(_0091_));
 sg13g2_mux2_1 _1209_ (.A0(net135),
    .A1(net303),
    .S(_0544_),
    .X(_0092_));
 sg13g2_mux2_1 _1210_ (.A0(net133),
    .A1(net334),
    .S(_0544_),
    .X(_0093_));
 sg13g2_mux2_1 _1211_ (.A0(net129),
    .A1(net364),
    .S(_0544_),
    .X(_0094_));
 sg13g2_mux2_1 _1212_ (.A0(net131),
    .A1(net302),
    .S(_0544_),
    .X(_0095_));
 sg13g2_mux2_1 _1213_ (.A0(net127),
    .A1(net366),
    .S(_0544_),
    .X(_0096_));
 sg13g2_mux2_1 _1214_ (.A0(net125),
    .A1(net385),
    .S(_0544_),
    .X(_0097_));
 sg13g2_mux2_1 _1215_ (.A0(net123),
    .A1(net404),
    .S(_0544_),
    .X(_0098_));
 sg13g2_and2_1 _1216_ (.A(net180),
    .B(net145),
    .X(_0545_));
 sg13g2_nand2_1 _1217_ (.Y(_0546_),
    .A(net275),
    .B(_0545_));
 sg13g2_o21ai_1 _1218_ (.B1(_0546_),
    .Y(_0099_),
    .A1(net145),
    .A2(_0263_));
 sg13g2_nand2_1 _1219_ (.Y(_0547_),
    .A(net277),
    .B(_0545_));
 sg13g2_o21ai_1 _1220_ (.B1(_0547_),
    .Y(_0100_),
    .A1(_0253_),
    .A2(_0299_));
 sg13g2_nand2_1 _1221_ (.Y(_0548_),
    .A(net283),
    .B(_0545_));
 sg13g2_o21ai_1 _1222_ (.B1(_0548_),
    .Y(_0101_),
    .A1(_0253_),
    .A2(_0333_));
 sg13g2_nand2_1 _1223_ (.Y(_0549_),
    .A(net291),
    .B(_0545_));
 sg13g2_o21ai_1 _1224_ (.B1(_0549_),
    .Y(_0102_),
    .A1(net145),
    .A2(_0367_));
 sg13g2_nand2_1 _1225_ (.Y(_0550_),
    .A(net281),
    .B(_0545_));
 sg13g2_o21ai_1 _1226_ (.B1(_0550_),
    .Y(_0103_),
    .A1(net145),
    .A2(_0398_));
 sg13g2_nand2_1 _1227_ (.Y(_0551_),
    .A(net282),
    .B(_0545_));
 sg13g2_o21ai_1 _1228_ (.B1(_0551_),
    .Y(_0104_),
    .A1(net145),
    .A2(_0430_));
 sg13g2_nand2_1 _1229_ (.Y(_0552_),
    .A(net293),
    .B(_0545_));
 sg13g2_o21ai_1 _1230_ (.B1(_0552_),
    .Y(_0105_),
    .A1(net145),
    .A2(_0461_));
 sg13g2_nand2_1 _1231_ (.Y(_0553_),
    .A(net279),
    .B(_0545_));
 sg13g2_o21ai_1 _1232_ (.B1(_0553_),
    .Y(_0106_),
    .A1(net145),
    .A2(_0486_));
 sg13g2_nand2_1 _1233_ (.Y(_0554_),
    .A(_0205_),
    .B(_0496_));
 sg13g2_nand3_1 _1234_ (.B(_0496_),
    .C(_0504_),
    .A(_0205_),
    .Y(_0555_));
 sg13g2_mux2_1 _1235_ (.A0(net137),
    .A1(net348),
    .S(_0555_),
    .X(_0107_));
 sg13g2_mux2_1 _1236_ (.A0(net135),
    .A1(net320),
    .S(_0555_),
    .X(_0108_));
 sg13g2_mux2_1 _1237_ (.A0(net133),
    .A1(net297),
    .S(_0555_),
    .X(_0109_));
 sg13g2_mux2_1 _1238_ (.A0(net129),
    .A1(net296),
    .S(_0555_),
    .X(_0110_));
 sg13g2_mux2_1 _1239_ (.A0(net131),
    .A1(net330),
    .S(_0555_),
    .X(_0111_));
 sg13g2_mux2_1 _1240_ (.A0(net127),
    .A1(net419),
    .S(_0555_),
    .X(_0112_));
 sg13g2_mux2_1 _1241_ (.A0(net125),
    .A1(net313),
    .S(_0555_),
    .X(_0113_));
 sg13g2_mux2_1 _1242_ (.A0(net123),
    .A1(net328),
    .S(_0555_),
    .X(_0114_));
 sg13g2_or2_1 _1243_ (.X(_0556_),
    .B(_0495_),
    .A(_0206_));
 sg13g2_mux2_1 _1244_ (.A0(net136),
    .A1(net418),
    .S(_0556_),
    .X(_0115_));
 sg13g2_mux2_1 _1245_ (.A0(net134),
    .A1(net361),
    .S(_0556_),
    .X(_0116_));
 sg13g2_mux2_1 _1246_ (.A0(net132),
    .A1(net304),
    .S(_0556_),
    .X(_0117_));
 sg13g2_mux2_1 _1247_ (.A0(net128),
    .A1(net341),
    .S(_0556_),
    .X(_0118_));
 sg13g2_mux2_1 _1248_ (.A0(net130),
    .A1(net357),
    .S(_0556_),
    .X(_0119_));
 sg13g2_mux2_1 _1249_ (.A0(net126),
    .A1(net337),
    .S(_0556_),
    .X(_0120_));
 sg13g2_mux2_1 _1250_ (.A0(net124),
    .A1(net384),
    .S(_0556_),
    .X(_0121_));
 sg13g2_mux2_1 _1251_ (.A0(net122),
    .A1(net414),
    .S(_0556_),
    .X(_0122_));
 sg13g2_or2_1 _1252_ (.X(_0557_),
    .B(_0506_),
    .A(_0206_));
 sg13g2_mux2_1 _1253_ (.A0(net136),
    .A1(net392),
    .S(_0557_),
    .X(_0123_));
 sg13g2_mux2_1 _1254_ (.A0(net134),
    .A1(net368),
    .S(_0557_),
    .X(_0124_));
 sg13g2_mux2_1 _1255_ (.A0(net132),
    .A1(net397),
    .S(_0557_),
    .X(_0125_));
 sg13g2_mux2_1 _1256_ (.A0(net128),
    .A1(net374),
    .S(_0557_),
    .X(_0126_));
 sg13g2_mux2_1 _1257_ (.A0(net130),
    .A1(net331),
    .S(_0557_),
    .X(_0127_));
 sg13g2_mux2_1 _1258_ (.A0(net126),
    .A1(net395),
    .S(_0557_),
    .X(_0128_));
 sg13g2_mux2_1 _1259_ (.A0(net124),
    .A1(net336),
    .S(_0557_),
    .X(_0129_));
 sg13g2_mux2_1 _1260_ (.A0(net122),
    .A1(net332),
    .S(_0557_),
    .X(_0130_));
 sg13g2_nand2b_2 _1261_ (.Y(_0558_),
    .B(_0504_),
    .A_N(_0497_));
 sg13g2_mux2_1 _1262_ (.A0(net136),
    .A1(net405),
    .S(_0558_),
    .X(_0131_));
 sg13g2_mux2_1 _1263_ (.A0(net134),
    .A1(net317),
    .S(_0558_),
    .X(_0132_));
 sg13g2_mux2_1 _1264_ (.A0(net132),
    .A1(net372),
    .S(_0558_),
    .X(_0133_));
 sg13g2_mux2_1 _1265_ (.A0(net128),
    .A1(net420),
    .S(_0558_),
    .X(_0134_));
 sg13g2_mux2_1 _1266_ (.A0(net130),
    .A1(net327),
    .S(_0558_),
    .X(_0135_));
 sg13g2_mux2_1 _1267_ (.A0(net126),
    .A1(net375),
    .S(_0558_),
    .X(_0136_));
 sg13g2_mux2_1 _1268_ (.A0(net124),
    .A1(net333),
    .S(_0558_),
    .X(_0137_));
 sg13g2_mux2_1 _1269_ (.A0(net122),
    .A1(net309),
    .S(_0558_),
    .X(_0138_));
 sg13g2_or2_1 _1270_ (.X(_0559_),
    .B(_0554_),
    .A(_0495_));
 sg13g2_mux2_1 _1271_ (.A0(net137),
    .A1(net347),
    .S(_0559_),
    .X(_0139_));
 sg13g2_mux2_1 _1272_ (.A0(net135),
    .A1(net308),
    .S(_0559_),
    .X(_0140_));
 sg13g2_mux2_1 _1273_ (.A0(net133),
    .A1(net319),
    .S(_0559_),
    .X(_0141_));
 sg13g2_mux2_1 _1274_ (.A0(net129),
    .A1(net377),
    .S(_0559_),
    .X(_0142_));
 sg13g2_mux2_1 _1275_ (.A0(net131),
    .A1(net426),
    .S(_0559_),
    .X(_0143_));
 sg13g2_mux2_1 _1276_ (.A0(net127),
    .A1(net373),
    .S(_0559_),
    .X(_0144_));
 sg13g2_mux2_1 _1277_ (.A0(net125),
    .A1(net370),
    .S(_0559_),
    .X(_0145_));
 sg13g2_mux2_1 _1278_ (.A0(net123),
    .A1(net311),
    .S(_0559_),
    .X(_0146_));
 sg13g2_or2_1 _1279_ (.X(_0560_),
    .B(_0554_),
    .A(_0506_));
 sg13g2_mux2_1 _1280_ (.A0(net137),
    .A1(net312),
    .S(_0560_),
    .X(_0147_));
 sg13g2_mux2_1 _1281_ (.A0(net135),
    .A1(net380),
    .S(_0560_),
    .X(_0148_));
 sg13g2_mux2_1 _1282_ (.A0(net133),
    .A1(net382),
    .S(_0560_),
    .X(_0149_));
 sg13g2_mux2_1 _1283_ (.A0(net129),
    .A1(net354),
    .S(_0560_),
    .X(_0150_));
 sg13g2_mux2_1 _1284_ (.A0(net131),
    .A1(net402),
    .S(_0560_),
    .X(_0151_));
 sg13g2_mux2_1 _1285_ (.A0(net127),
    .A1(net335),
    .S(_0560_),
    .X(_0152_));
 sg13g2_mux2_1 _1286_ (.A0(net125),
    .A1(net381),
    .S(_0560_),
    .X(_0153_));
 sg13g2_mux2_1 _1287_ (.A0(net123),
    .A1(net369),
    .S(_0560_),
    .X(_0154_));
 sg13g2_or2_1 _1288_ (.X(_0561_),
    .B(_0554_),
    .A(_0209_));
 sg13g2_mux2_1 _1289_ (.A0(net137),
    .A1(net322),
    .S(net138),
    .X(_0155_));
 sg13g2_nor2_1 _1290_ (.A(net135),
    .B(net138),
    .Y(_0562_));
 sg13g2_a21oi_1 _1291_ (.A1(_0185_),
    .A2(net138),
    .Y(_0156_),
    .B1(_0562_));
 sg13g2_mux2_1 _1292_ (.A0(net133),
    .A1(net416),
    .S(net138),
    .X(_0157_));
 sg13g2_mux2_1 _1293_ (.A0(net129),
    .A1(net358),
    .S(net138),
    .X(_0158_));
 sg13g2_mux2_1 _1294_ (.A0(net131),
    .A1(net389),
    .S(net138),
    .X(_0159_));
 sg13g2_mux2_1 _1295_ (.A0(net127),
    .A1(net391),
    .S(net138),
    .X(_0160_));
 sg13g2_mux2_1 _1296_ (.A0(net125),
    .A1(net352),
    .S(_0561_),
    .X(_0161_));
 sg13g2_mux2_1 _1297_ (.A0(net123),
    .A1(net410),
    .S(net138),
    .X(_0162_));
 sg13g2_and2_1 _1298_ (.A(net180),
    .B(_0240_),
    .X(_0563_));
 sg13g2_nand2_1 _1299_ (.Y(_0564_),
    .A(net399),
    .B(_0563_));
 sg13g2_o21ai_1 _1300_ (.B1(_0564_),
    .Y(_0163_),
    .A1(_0240_),
    .A2(_0263_));
 sg13g2_nand2_1 _1301_ (.Y(_0565_),
    .A(net289),
    .B(_0563_));
 sg13g2_o21ai_1 _1302_ (.B1(_0565_),
    .Y(_0164_),
    .A1(_0240_),
    .A2(_0299_));
 sg13g2_nand2_1 _1303_ (.Y(_0566_),
    .A(net276),
    .B(_0563_));
 sg13g2_o21ai_1 _1304_ (.B1(_0566_),
    .Y(_0165_),
    .A1(net143),
    .A2(_0333_));
 sg13g2_nand2_1 _1305_ (.Y(_0567_),
    .A(net292),
    .B(_0563_));
 sg13g2_o21ai_1 _1306_ (.B1(_0567_),
    .Y(_0166_),
    .A1(net143),
    .A2(_0367_));
 sg13g2_nand2_1 _1307_ (.Y(_0568_),
    .A(net299),
    .B(_0563_));
 sg13g2_o21ai_1 _1308_ (.B1(_0568_),
    .Y(_0167_),
    .A1(net143),
    .A2(_0398_));
 sg13g2_nand2_1 _1309_ (.Y(_0569_),
    .A(net310),
    .B(_0563_));
 sg13g2_o21ai_1 _1310_ (.B1(_0569_),
    .Y(_0168_),
    .A1(net143),
    .A2(_0430_));
 sg13g2_nand2_1 _1311_ (.Y(_0570_),
    .A(net305),
    .B(_0563_));
 sg13g2_o21ai_1 _1312_ (.B1(_0570_),
    .Y(_0169_),
    .A1(net143),
    .A2(_0461_));
 sg13g2_nand2_1 _1313_ (.Y(_0571_),
    .A(net287),
    .B(_0563_));
 sg13g2_o21ai_1 _1314_ (.B1(_0571_),
    .Y(_0170_),
    .A1(net143),
    .A2(_0486_));
 sg13g2_nor2_1 _1315_ (.A(_0258_),
    .B(_0267_),
    .Y(_0572_));
 sg13g2_or2_1 _1316_ (.X(_0573_),
    .B(_0267_),
    .A(_0258_));
 sg13g2_nand2_1 _1317_ (.Y(_0574_),
    .A(net436),
    .B(_0572_));
 sg13g2_nor3_1 _1318_ (.A(_0256_),
    .B(_0274_),
    .C(_0572_),
    .Y(_0575_));
 sg13g2_nand4_1 _1319_ (.B(_0407_),
    .C(_0436_),
    .A(_0371_),
    .Y(_0576_),
    .D(_0575_));
 sg13g2_o21ai_1 _1320_ (.B1(_0574_),
    .Y(_0577_),
    .A1(_0469_),
    .A2(_0576_));
 sg13g2_and2_1 _1321_ (.A(net180),
    .B(_0577_),
    .X(_0171_));
 sg13g2_o21ai_1 _1322_ (.B1(_0270_),
    .Y(_0578_),
    .A1(net287),
    .A2(_0466_));
 sg13g2_a21oi_1 _1323_ (.A1(_0435_),
    .A2(_0438_),
    .Y(_0579_),
    .B1(_0468_));
 sg13g2_a21o_1 _1324_ (.A2(_0467_),
    .A1(net424),
    .B1(_0579_),
    .X(_0580_));
 sg13g2_xnor2_1 _1325_ (.Y(_0581_),
    .A(_0578_),
    .B(_0580_));
 sg13g2_o21ai_1 _1326_ (.B1(net180),
    .Y(_0582_),
    .A1(net430),
    .A2(_0573_));
 sg13g2_a21oi_1 _1327_ (.A1(_0573_),
    .A2(_0581_),
    .Y(_0172_),
    .B1(_0582_));
 sg13g2_nand2b_2 _1328_ (.Y(_0583_),
    .B(_0504_),
    .A_N(_0499_));
 sg13g2_mux2_1 _1329_ (.A0(net137),
    .A1(net306),
    .S(_0583_),
    .X(_0173_));
 sg13g2_mux2_1 _1330_ (.A0(net135),
    .A1(net318),
    .S(_0583_),
    .X(_0174_));
 sg13g2_mux2_1 _1331_ (.A0(net133),
    .A1(net387),
    .S(_0583_),
    .X(_0175_));
 sg13g2_mux2_1 _1332_ (.A0(net129),
    .A1(net301),
    .S(_0583_),
    .X(_0176_));
 sg13g2_mux2_1 _1333_ (.A0(net131),
    .A1(net417),
    .S(_0583_),
    .X(_0177_));
 sg13g2_mux2_1 _1334_ (.A0(net127),
    .A1(net345),
    .S(_0583_),
    .X(_0178_));
 sg13g2_mux2_1 _1335_ (.A0(net125),
    .A1(net393),
    .S(_0583_),
    .X(_0179_));
 sg13g2_mux2_1 _1336_ (.A0(net123),
    .A1(net355),
    .S(_0583_),
    .X(_0180_));
 sg13g2_a21oi_1 _1337_ (.A1(_0263_),
    .A2(net141),
    .Y(_0083_),
    .B1(_0491_));
 sg13g2_a21oi_1 _1338_ (.A1(_0299_),
    .A2(net141),
    .Y(_0084_),
    .B1(_0492_));
 sg13g2_a21oi_1 _1339_ (.A1(_0333_),
    .A2(net142),
    .Y(_0085_),
    .B1(_0493_));
 sg13g2_a21oi_1 _1340_ (.A1(_0367_),
    .A2(net142),
    .Y(_0086_),
    .B1(_0494_));
 sg13g2_dfrbpq_1 _1341_ (.RESET_B(net92),
    .D(_0004_),
    .Q(\cpu0.ram[5][0] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1342_ (.RESET_B(net242),
    .D(_0005_),
    .Q(\cpu0.ram[5][1] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1343_ (.RESET_B(net241),
    .D(_0006_),
    .Q(\cpu0.ram[5][2] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1344_ (.RESET_B(net240),
    .D(_0007_),
    .Q(\cpu0.ram[5][3] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1345_ (.RESET_B(net239),
    .D(_0008_),
    .Q(\cpu0.ram[5][4] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1346_ (.RESET_B(net238),
    .D(_0009_),
    .Q(\cpu0.ram[5][5] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1347_ (.RESET_B(net237),
    .D(_0010_),
    .Q(\cpu0.ram[5][6] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1348_ (.RESET_B(net236),
    .D(_0011_),
    .Q(\cpu0.ram[5][7] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_2 _1349_ (.RESET_B(net235),
    .D(_0012_),
    .Q(_0000_),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_2 _1350_ (.RESET_B(net234),
    .D(_0013_),
    .Q(_0001_),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1351_ (.RESET_B(net233),
    .D(_0014_),
    .Q(_0002_),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1352_ (.RESET_B(net232),
    .D(_0015_),
    .Q(_0003_),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1353_ (.RESET_B(net231),
    .D(_0016_),
    .Q(\cpu0.ram[2][0] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1354_ (.RESET_B(net230),
    .D(_0017_),
    .Q(\cpu0.ram[2][1] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1355_ (.RESET_B(net229),
    .D(_0018_),
    .Q(\cpu0.ram[2][2] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1356_ (.RESET_B(net228),
    .D(_0019_),
    .Q(\cpu0.ram[2][3] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1357_ (.RESET_B(net227),
    .D(_0020_),
    .Q(\cpu0.ram[2][4] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1358_ (.RESET_B(net226),
    .D(_0021_),
    .Q(\cpu0.ram[2][5] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1359_ (.RESET_B(net225),
    .D(_0022_),
    .Q(\cpu0.ram[2][6] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1360_ (.RESET_B(net224),
    .D(_0023_),
    .Q(\cpu0.ram[2][7] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_2 _1361_ (.RESET_B(net223),
    .D(_0024_),
    .Q(\cpu0.step[1] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1362_ (.RESET_B(net222),
    .D(_0025_),
    .Q(\cpu0.step[2] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1363_ (.RESET_B(net221),
    .D(_0026_),
    .Q(\cpu0.ram[14][0] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1364_ (.RESET_B(net220),
    .D(_0027_),
    .Q(\cpu0.ram[14][1] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1365_ (.RESET_B(net219),
    .D(_0028_),
    .Q(\cpu0.ram[14][2] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1366_ (.RESET_B(net218),
    .D(_0029_),
    .Q(\cpu0.ram[14][3] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1367_ (.RESET_B(net217),
    .D(_0030_),
    .Q(\cpu0.ram[14][4] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1368_ (.RESET_B(net216),
    .D(_0031_),
    .Q(\cpu0.ram[14][5] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1369_ (.RESET_B(net215),
    .D(_0032_),
    .Q(\cpu0.ram[14][6] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1370_ (.RESET_B(net214),
    .D(_0033_),
    .Q(\cpu0.ram[14][7] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _1371_ (.RESET_B(net213),
    .D(_0034_),
    .Q(\cpu0.step[0] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1372_ (.RESET_B(net212),
    .D(_0035_),
    .Q(\cpu0.ram[4][0] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1373_ (.RESET_B(net211),
    .D(_0036_),
    .Q(\cpu0.ram[4][1] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1374_ (.RESET_B(net210),
    .D(_0037_),
    .Q(\cpu0.ram[4][2] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1375_ (.RESET_B(net209),
    .D(_0038_),
    .Q(\cpu0.ram[4][3] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1376_ (.RESET_B(net208),
    .D(_0039_),
    .Q(\cpu0.ram[4][4] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1377_ (.RESET_B(net207),
    .D(_0040_),
    .Q(\cpu0.ram[4][5] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1378_ (.RESET_B(net206),
    .D(_0041_),
    .Q(\cpu0.ram[4][6] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1379_ (.RESET_B(net205),
    .D(_0042_),
    .Q(\cpu0.ram[4][7] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1380_ (.RESET_B(net204),
    .D(_0043_),
    .Q(\cpu0.ram[3][0] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1381_ (.RESET_B(net203),
    .D(_0044_),
    .Q(\cpu0.ram[3][1] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1382_ (.RESET_B(net202),
    .D(_0045_),
    .Q(\cpu0.ram[3][2] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1383_ (.RESET_B(net201),
    .D(_0046_),
    .Q(\cpu0.ram[3][3] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1384_ (.RESET_B(net200),
    .D(_0047_),
    .Q(\cpu0.ram[3][4] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1385_ (.RESET_B(net199),
    .D(_0048_),
    .Q(\cpu0.ram[3][5] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1386_ (.RESET_B(net198),
    .D(_0049_),
    .Q(\cpu0.ram[3][6] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1387_ (.RESET_B(net197),
    .D(_0050_),
    .Q(\cpu0.ram[3][7] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1388_ (.RESET_B(net196),
    .D(_0051_),
    .Q(\cpu0.ram[1][0] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1389_ (.RESET_B(net195),
    .D(_0052_),
    .Q(\cpu0.ram[1][1] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1390_ (.RESET_B(net194),
    .D(_0053_),
    .Q(\cpu0.ram[1][2] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1391_ (.RESET_B(net193),
    .D(_0054_),
    .Q(\cpu0.ram[1][3] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1392_ (.RESET_B(net192),
    .D(_0055_),
    .Q(\cpu0.ram[1][4] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1393_ (.RESET_B(net191),
    .D(_0056_),
    .Q(\cpu0.ram[1][5] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1394_ (.RESET_B(net190),
    .D(_0057_),
    .Q(\cpu0.ram[1][6] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1395_ (.RESET_B(net189),
    .D(_0058_),
    .Q(\cpu0.ram[1][7] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1396_ (.RESET_B(net188),
    .D(_0059_),
    .Q(\cpu0.ram[15][0] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1397_ (.RESET_B(net187),
    .D(_0060_),
    .Q(\cpu0.ram[15][1] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1398_ (.RESET_B(net186),
    .D(_0061_),
    .Q(\cpu0.ram[15][2] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1399_ (.RESET_B(net185),
    .D(_0062_),
    .Q(\cpu0.ram[15][3] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1400_ (.RESET_B(net184),
    .D(_0063_),
    .Q(\cpu0.ram[15][4] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1401_ (.RESET_B(net183),
    .D(_0064_),
    .Q(\cpu0.ram[15][5] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1402_ (.RESET_B(net182),
    .D(_0065_),
    .Q(\cpu0.ram[15][6] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1403_ (.RESET_B(net181),
    .D(_0066_),
    .Q(\cpu0.ram[15][7] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _1404_ (.RESET_B(net121),
    .D(_0067_),
    .Q(\cpu0.a_reg[0] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 _1405_ (.RESET_B(net119),
    .D(_0068_),
    .Q(\cpu0.a_reg[1] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _1406_ (.RESET_B(net117),
    .D(_0069_),
    .Q(\cpu0.a_reg[2] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _1407_ (.RESET_B(net115),
    .D(_0070_),
    .Q(\cpu0.a_reg[3] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _1408_ (.RESET_B(net113),
    .D(_0071_),
    .Q(\cpu0.a_reg[4] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 _1409_ (.RESET_B(net111),
    .D(_0072_),
    .Q(\cpu0.a_reg[5] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 _1410_ (.RESET_B(net109),
    .D(_0073_),
    .Q(\cpu0.a_reg[6] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 _1411_ (.RESET_B(net107),
    .D(_0074_),
    .Q(\cpu0.a_reg[7] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1412_ (.RESET_B(net105),
    .D(_0075_),
    .Q(\cpu0.ir[0] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1413_ (.RESET_B(net103),
    .D(_0076_),
    .Q(\cpu0.ir[1] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1414_ (.RESET_B(net101),
    .D(_0077_),
    .Q(\cpu0.ir[2] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1415_ (.RESET_B(net99),
    .D(_0078_),
    .Q(\cpu0.ir[3] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 _1416_ (.RESET_B(net97),
    .D(_0079_),
    .Q(\cpu0.ir[4] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1417_ (.RESET_B(net95),
    .D(_0080_),
    .Q(\cpu0.ir[5] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _1418_ (.RESET_B(net93),
    .D(_0081_),
    .Q(\cpu0.ir[6] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _1419_ (.RESET_B(net91),
    .D(_0082_),
    .Q(\cpu0.ir[7] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1420_ (.RESET_B(net89),
    .D(_0083_),
    .Q(\cpu0.mar[0] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1421_ (.RESET_B(net87),
    .D(_0084_),
    .Q(\cpu0.mar[1] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1422_ (.RESET_B(net85),
    .D(_0085_),
    .Q(\cpu0.mar[2] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1423_ (.RESET_B(net83),
    .D(_0086_),
    .Q(\cpu0.mar[3] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 _1424_ (.RESET_B(net81),
    .D(_0087_),
    .Q(\cpu0.pc[0] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _1425_ (.RESET_B(net79),
    .D(_0088_),
    .Q(\cpu0.pc[1] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _1426_ (.RESET_B(net77),
    .D(_0089_),
    .Q(\cpu0.pc[2] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1427_ (.RESET_B(net75),
    .D(_0090_),
    .Q(\cpu0.pc[3] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1428_ (.RESET_B(net73),
    .D(_0091_),
    .Q(\cpu0.ram[13][0] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1429_ (.RESET_B(net72),
    .D(_0092_),
    .Q(\cpu0.ram[13][1] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1430_ (.RESET_B(net71),
    .D(_0093_),
    .Q(\cpu0.ram[13][2] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1431_ (.RESET_B(net70),
    .D(_0094_),
    .Q(\cpu0.ram[13][3] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1432_ (.RESET_B(net69),
    .D(_0095_),
    .Q(\cpu0.ram[13][4] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1433_ (.RESET_B(net68),
    .D(_0096_),
    .Q(\cpu0.ram[13][5] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1434_ (.RESET_B(net67),
    .D(_0097_),
    .Q(\cpu0.ram[13][6] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1435_ (.RESET_B(net66),
    .D(_0098_),
    .Q(\cpu0.ram[13][7] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1436_ (.RESET_B(net65),
    .D(_0099_),
    .Q(uo_out[0]),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1437_ (.RESET_B(net63),
    .D(net278),
    .Q(uo_out[1]),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1438_ (.RESET_B(net61),
    .D(net284),
    .Q(uo_out[2]),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1439_ (.RESET_B(net59),
    .D(_0102_),
    .Q(uo_out[3]),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1440_ (.RESET_B(net57),
    .D(_0103_),
    .Q(uo_out[4]),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1441_ (.RESET_B(net55),
    .D(_0104_),
    .Q(uo_out[5]),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1442_ (.RESET_B(net53),
    .D(_0105_),
    .Q(uo_out[6]),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1443_ (.RESET_B(net51),
    .D(net280),
    .Q(uo_out[7]),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1444_ (.RESET_B(net49),
    .D(_0107_),
    .Q(\cpu0.ram[8][0] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1445_ (.RESET_B(net48),
    .D(_0108_),
    .Q(\cpu0.ram[8][1] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1446_ (.RESET_B(net47),
    .D(_0109_),
    .Q(\cpu0.ram[8][2] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1447_ (.RESET_B(net46),
    .D(_0110_),
    .Q(\cpu0.ram[8][3] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1448_ (.RESET_B(net45),
    .D(_0111_),
    .Q(\cpu0.ram[8][4] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1449_ (.RESET_B(net44),
    .D(_0112_),
    .Q(\cpu0.ram[8][5] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1450_ (.RESET_B(net43),
    .D(_0113_),
    .Q(\cpu0.ram[8][6] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1451_ (.RESET_B(net42),
    .D(_0114_),
    .Q(\cpu0.ram[8][7] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1452_ (.RESET_B(net41),
    .D(_0115_),
    .Q(\cpu0.ram[6][0] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1453_ (.RESET_B(net40),
    .D(_0116_),
    .Q(\cpu0.ram[6][1] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1454_ (.RESET_B(net39),
    .D(_0117_),
    .Q(\cpu0.ram[6][2] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1455_ (.RESET_B(net38),
    .D(_0118_),
    .Q(\cpu0.ram[6][3] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1456_ (.RESET_B(net37),
    .D(_0119_),
    .Q(\cpu0.ram[6][4] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1457_ (.RESET_B(net36),
    .D(_0120_),
    .Q(\cpu0.ram[6][5] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1458_ (.RESET_B(net35),
    .D(_0121_),
    .Q(\cpu0.ram[6][6] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1459_ (.RESET_B(net34),
    .D(_0122_),
    .Q(\cpu0.ram[6][7] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1460_ (.RESET_B(net33),
    .D(_0123_),
    .Q(\cpu0.ram[7][0] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1461_ (.RESET_B(net32),
    .D(_0124_),
    .Q(\cpu0.ram[7][1] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1462_ (.RESET_B(net31),
    .D(_0125_),
    .Q(\cpu0.ram[7][2] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1463_ (.RESET_B(net30),
    .D(_0126_),
    .Q(\cpu0.ram[7][3] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1464_ (.RESET_B(net265),
    .D(_0127_),
    .Q(\cpu0.ram[7][4] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1465_ (.RESET_B(net264),
    .D(_0128_),
    .Q(\cpu0.ram[7][5] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1466_ (.RESET_B(net263),
    .D(_0129_),
    .Q(\cpu0.ram[7][6] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1467_ (.RESET_B(net262),
    .D(_0130_),
    .Q(\cpu0.ram[7][7] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1468_ (.RESET_B(net261),
    .D(_0131_),
    .Q(\cpu0.ram[0][0] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1469_ (.RESET_B(net260),
    .D(_0132_),
    .Q(\cpu0.ram[0][1] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1470_ (.RESET_B(net259),
    .D(_0133_),
    .Q(\cpu0.ram[0][2] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1471_ (.RESET_B(net258),
    .D(_0134_),
    .Q(\cpu0.ram[0][3] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1472_ (.RESET_B(net257),
    .D(_0135_),
    .Q(\cpu0.ram[0][4] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1473_ (.RESET_B(net256),
    .D(_0136_),
    .Q(\cpu0.ram[0][5] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1474_ (.RESET_B(net255),
    .D(_0137_),
    .Q(\cpu0.ram[0][6] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1475_ (.RESET_B(net254),
    .D(_0138_),
    .Q(\cpu0.ram[0][7] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1476_ (.RESET_B(net253),
    .D(_0139_),
    .Q(\cpu0.ram[10][0] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1477_ (.RESET_B(net252),
    .D(_0140_),
    .Q(\cpu0.ram[10][1] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1478_ (.RESET_B(net251),
    .D(_0141_),
    .Q(\cpu0.ram[10][2] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1479_ (.RESET_B(net250),
    .D(_0142_),
    .Q(\cpu0.ram[10][3] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1480_ (.RESET_B(net249),
    .D(_0143_),
    .Q(\cpu0.ram[10][4] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1481_ (.RESET_B(net248),
    .D(_0144_),
    .Q(\cpu0.ram[10][5] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1482_ (.RESET_B(net247),
    .D(_0145_),
    .Q(\cpu0.ram[10][6] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1483_ (.RESET_B(net246),
    .D(_0146_),
    .Q(\cpu0.ram[10][7] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1484_ (.RESET_B(net245),
    .D(_0147_),
    .Q(\cpu0.ram[11][0] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1485_ (.RESET_B(net244),
    .D(_0148_),
    .Q(\cpu0.ram[11][1] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1486_ (.RESET_B(net243),
    .D(_0149_),
    .Q(\cpu0.ram[11][2] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1487_ (.RESET_B(net120),
    .D(_0150_),
    .Q(\cpu0.ram[11][3] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1488_ (.RESET_B(net118),
    .D(_0151_),
    .Q(\cpu0.ram[11][4] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1489_ (.RESET_B(net116),
    .D(_0152_),
    .Q(\cpu0.ram[11][5] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1490_ (.RESET_B(net114),
    .D(_0153_),
    .Q(\cpu0.ram[11][6] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1491_ (.RESET_B(net112),
    .D(_0154_),
    .Q(\cpu0.ram[11][7] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1492_ (.RESET_B(net110),
    .D(_0155_),
    .Q(\cpu0.ram[9][0] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1493_ (.RESET_B(net108),
    .D(_0156_),
    .Q(\cpu0.ram[9][1] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1494_ (.RESET_B(net106),
    .D(_0157_),
    .Q(\cpu0.ram[9][2] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1495_ (.RESET_B(net104),
    .D(_0158_),
    .Q(\cpu0.ram[9][3] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1496_ (.RESET_B(net102),
    .D(_0159_),
    .Q(\cpu0.ram[9][4] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1497_ (.RESET_B(net100),
    .D(_0160_),
    .Q(\cpu0.ram[9][5] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1498_ (.RESET_B(net98),
    .D(_0161_),
    .Q(\cpu0.ram[9][6] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1499_ (.RESET_B(net96),
    .D(_0162_),
    .Q(\cpu0.ram[9][7] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _1500_ (.RESET_B(net94),
    .D(net400),
    .Q(\cpu0.b_reg[0] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1501_ (.RESET_B(net90),
    .D(net290),
    .Q(\cpu0.b_reg[1] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1502_ (.RESET_B(net86),
    .D(_0165_),
    .Q(\cpu0.b_reg[2] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _1503_ (.RESET_B(net82),
    .D(_0166_),
    .Q(\cpu0.b_reg[3] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1504_ (.RESET_B(net78),
    .D(_0167_),
    .Q(\cpu0.b_reg[4] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1505_ (.RESET_B(net74),
    .D(_0168_),
    .Q(\cpu0.b_reg[5] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1506_ (.RESET_B(net62),
    .D(_0169_),
    .Q(\cpu0.b_reg[6] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1507_ (.RESET_B(net58),
    .D(net288),
    .Q(\cpu0.b_reg[7] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1508_ (.RESET_B(net54),
    .D(_0171_),
    .Q(\cpu0.zero_flag ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1509_ (.RESET_B(net50),
    .D(net431),
    .Q(\cpu0.carry_flag ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1510_ (.RESET_B(net88),
    .D(_0173_),
    .Q(\cpu0.ram[12][0] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1511_ (.RESET_B(net84),
    .D(_0174_),
    .Q(\cpu0.ram[12][1] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1512_ (.RESET_B(net80),
    .D(_0175_),
    .Q(\cpu0.ram[12][2] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1513_ (.RESET_B(net76),
    .D(_0176_),
    .Q(\cpu0.ram[12][3] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1514_ (.RESET_B(net64),
    .D(_0177_),
    .Q(\cpu0.ram[12][4] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1515_ (.RESET_B(net60),
    .D(_0178_),
    .Q(\cpu0.ram[12][5] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1516_ (.RESET_B(net56),
    .D(_0179_),
    .Q(\cpu0.ram[12][6] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1517_ (.RESET_B(net52),
    .D(_0180_),
    .Q(\cpu0.ram[12][7] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_tiehi _1462__31 (.L_HI(net31));
 sg13g2_tiehi _1461__32 (.L_HI(net32));
 sg13g2_tiehi _1460__33 (.L_HI(net33));
 sg13g2_tiehi _1459__34 (.L_HI(net34));
 sg13g2_tiehi _1458__35 (.L_HI(net35));
 sg13g2_tiehi _1457__36 (.L_HI(net36));
 sg13g2_tiehi _1456__37 (.L_HI(net37));
 sg13g2_tiehi _1455__38 (.L_HI(net38));
 sg13g2_tiehi _1454__39 (.L_HI(net39));
 sg13g2_tiehi _1453__40 (.L_HI(net40));
 sg13g2_tiehi _1452__41 (.L_HI(net41));
 sg13g2_tiehi _1451__42 (.L_HI(net42));
 sg13g2_tiehi _1450__43 (.L_HI(net43));
 sg13g2_tiehi _1449__44 (.L_HI(net44));
 sg13g2_tiehi _1448__45 (.L_HI(net45));
 sg13g2_tiehi _1447__46 (.L_HI(net46));
 sg13g2_tiehi _1446__47 (.L_HI(net47));
 sg13g2_tiehi _1445__48 (.L_HI(net48));
 sg13g2_tiehi _1444__49 (.L_HI(net49));
 sg13g2_tiehi _1509__50 (.L_HI(net50));
 sg13g2_tiehi _1443__51 (.L_HI(net51));
 sg13g2_tiehi _1517__52 (.L_HI(net52));
 sg13g2_tiehi _1442__53 (.L_HI(net53));
 sg13g2_tiehi _1508__54 (.L_HI(net54));
 sg13g2_tiehi _1441__55 (.L_HI(net55));
 sg13g2_tiehi _1516__56 (.L_HI(net56));
 sg13g2_tiehi _1440__57 (.L_HI(net57));
 sg13g2_tiehi _1507__58 (.L_HI(net58));
 sg13g2_tiehi _1439__59 (.L_HI(net59));
 sg13g2_tiehi _1515__60 (.L_HI(net60));
 sg13g2_tiehi _1438__61 (.L_HI(net61));
 sg13g2_tiehi _1506__62 (.L_HI(net62));
 sg13g2_tiehi _1437__63 (.L_HI(net63));
 sg13g2_tiehi _1514__64 (.L_HI(net64));
 sg13g2_tiehi _1436__65 (.L_HI(net65));
 sg13g2_tiehi _1435__66 (.L_HI(net66));
 sg13g2_tiehi _1434__67 (.L_HI(net67));
 sg13g2_tiehi _1433__68 (.L_HI(net68));
 sg13g2_tiehi _1432__69 (.L_HI(net69));
 sg13g2_tiehi _1431__70 (.L_HI(net70));
 sg13g2_tiehi _1430__71 (.L_HI(net71));
 sg13g2_tiehi _1429__72 (.L_HI(net72));
 sg13g2_tiehi _1428__73 (.L_HI(net73));
 sg13g2_tiehi _1505__74 (.L_HI(net74));
 sg13g2_tiehi _1427__75 (.L_HI(net75));
 sg13g2_tiehi _1513__76 (.L_HI(net76));
 sg13g2_tiehi _1426__77 (.L_HI(net77));
 sg13g2_tiehi _1504__78 (.L_HI(net78));
 sg13g2_tiehi _1425__79 (.L_HI(net79));
 sg13g2_tiehi _1512__80 (.L_HI(net80));
 sg13g2_tiehi _1424__81 (.L_HI(net81));
 sg13g2_tiehi _1503__82 (.L_HI(net82));
 sg13g2_tiehi _1423__83 (.L_HI(net83));
 sg13g2_tiehi _1511__84 (.L_HI(net84));
 sg13g2_tiehi _1422__85 (.L_HI(net85));
 sg13g2_tiehi _1502__86 (.L_HI(net86));
 sg13g2_tiehi _1421__87 (.L_HI(net87));
 sg13g2_tiehi _1510__88 (.L_HI(net88));
 sg13g2_tiehi _1420__89 (.L_HI(net89));
 sg13g2_tiehi _1501__90 (.L_HI(net90));
 sg13g2_tiehi _1419__91 (.L_HI(net91));
 sg13g2_tiehi _1341__92 (.L_HI(net92));
 sg13g2_tiehi _1418__93 (.L_HI(net93));
 sg13g2_tiehi _1500__94 (.L_HI(net94));
 sg13g2_tiehi _1417__95 (.L_HI(net95));
 sg13g2_tiehi _1499__96 (.L_HI(net96));
 sg13g2_tiehi _1416__97 (.L_HI(net97));
 sg13g2_tiehi _1498__98 (.L_HI(net98));
 sg13g2_tiehi _1415__99 (.L_HI(net99));
 sg13g2_tiehi _1497__100 (.L_HI(net100));
 sg13g2_tiehi _1414__101 (.L_HI(net101));
 sg13g2_tiehi _1496__102 (.L_HI(net102));
 sg13g2_tiehi _1413__103 (.L_HI(net103));
 sg13g2_tiehi _1495__104 (.L_HI(net104));
 sg13g2_tiehi _1412__105 (.L_HI(net105));
 sg13g2_tiehi _1494__106 (.L_HI(net106));
 sg13g2_tiehi _1411__107 (.L_HI(net107));
 sg13g2_tiehi _1493__108 (.L_HI(net108));
 sg13g2_tiehi _1410__109 (.L_HI(net109));
 sg13g2_tiehi _1492__110 (.L_HI(net110));
 sg13g2_tiehi _1409__111 (.L_HI(net111));
 sg13g2_tiehi _1491__112 (.L_HI(net112));
 sg13g2_tiehi _1408__113 (.L_HI(net113));
 sg13g2_tiehi _1490__114 (.L_HI(net114));
 sg13g2_tiehi _1407__115 (.L_HI(net115));
 sg13g2_tiehi _1489__116 (.L_HI(net116));
 sg13g2_tiehi _1406__117 (.L_HI(net117));
 sg13g2_tiehi _1488__118 (.L_HI(net118));
 sg13g2_tiehi _1405__119 (.L_HI(net119));
 sg13g2_tiehi _1487__120 (.L_HI(net120));
 sg13g2_tiehi _1404__121 (.L_HI(net121));
 sg13g2_tiehi _1403__122 (.L_HI(net181));
 sg13g2_tiehi _1402__123 (.L_HI(net182));
 sg13g2_tiehi _1401__124 (.L_HI(net183));
 sg13g2_tiehi _1400__125 (.L_HI(net184));
 sg13g2_tiehi _1399__126 (.L_HI(net185));
 sg13g2_tiehi _1398__127 (.L_HI(net186));
 sg13g2_tiehi _1397__128 (.L_HI(net187));
 sg13g2_tiehi _1396__129 (.L_HI(net188));
 sg13g2_tiehi _1395__130 (.L_HI(net189));
 sg13g2_tiehi _1394__131 (.L_HI(net190));
 sg13g2_tiehi _1393__132 (.L_HI(net191));
 sg13g2_tiehi _1392__133 (.L_HI(net192));
 sg13g2_tiehi _1391__134 (.L_HI(net193));
 sg13g2_tiehi _1390__135 (.L_HI(net194));
 sg13g2_tiehi _1389__136 (.L_HI(net195));
 sg13g2_tiehi _1388__137 (.L_HI(net196));
 sg13g2_tiehi _1387__138 (.L_HI(net197));
 sg13g2_tiehi _1386__139 (.L_HI(net198));
 sg13g2_tiehi _1385__140 (.L_HI(net199));
 sg13g2_tiehi _1384__141 (.L_HI(net200));
 sg13g2_tiehi _1383__142 (.L_HI(net201));
 sg13g2_tiehi _1382__143 (.L_HI(net202));
 sg13g2_tiehi _1381__144 (.L_HI(net203));
 sg13g2_tiehi _1380__145 (.L_HI(net204));
 sg13g2_tiehi _1379__146 (.L_HI(net205));
 sg13g2_tiehi _1378__147 (.L_HI(net206));
 sg13g2_tiehi _1377__148 (.L_HI(net207));
 sg13g2_tiehi _1376__149 (.L_HI(net208));
 sg13g2_tiehi _1375__150 (.L_HI(net209));
 sg13g2_tiehi _1374__151 (.L_HI(net210));
 sg13g2_tiehi _1373__152 (.L_HI(net211));
 sg13g2_tiehi _1372__153 (.L_HI(net212));
 sg13g2_tiehi _1371__154 (.L_HI(net213));
 sg13g2_tiehi _1370__155 (.L_HI(net214));
 sg13g2_tiehi _1369__156 (.L_HI(net215));
 sg13g2_tiehi _1368__157 (.L_HI(net216));
 sg13g2_tiehi _1367__158 (.L_HI(net217));
 sg13g2_tiehi _1366__159 (.L_HI(net218));
 sg13g2_tiehi _1365__160 (.L_HI(net219));
 sg13g2_tiehi _1364__161 (.L_HI(net220));
 sg13g2_tiehi _1363__162 (.L_HI(net221));
 sg13g2_tiehi _1362__163 (.L_HI(net222));
 sg13g2_tiehi _1361__164 (.L_HI(net223));
 sg13g2_tiehi _1360__165 (.L_HI(net224));
 sg13g2_tiehi _1359__166 (.L_HI(net225));
 sg13g2_tiehi _1358__167 (.L_HI(net226));
 sg13g2_tiehi _1357__168 (.L_HI(net227));
 sg13g2_tiehi _1356__169 (.L_HI(net228));
 sg13g2_tiehi _1355__170 (.L_HI(net229));
 sg13g2_tiehi _1354__171 (.L_HI(net230));
 sg13g2_tiehi _1353__172 (.L_HI(net231));
 sg13g2_tiehi _1352__173 (.L_HI(net232));
 sg13g2_tiehi _1351__174 (.L_HI(net233));
 sg13g2_tiehi _1350__175 (.L_HI(net234));
 sg13g2_tiehi _1349__176 (.L_HI(net235));
 sg13g2_tiehi _1348__177 (.L_HI(net236));
 sg13g2_tiehi _1347__178 (.L_HI(net237));
 sg13g2_tiehi _1346__179 (.L_HI(net238));
 sg13g2_tiehi _1345__180 (.L_HI(net239));
 sg13g2_tiehi _1344__181 (.L_HI(net240));
 sg13g2_tiehi _1343__182 (.L_HI(net241));
 sg13g2_tiehi _1342__183 (.L_HI(net242));
 sg13g2_tiehi _1486__184 (.L_HI(net243));
 sg13g2_tiehi _1485__185 (.L_HI(net244));
 sg13g2_tiehi _1484__186 (.L_HI(net245));
 sg13g2_tiehi _1483__187 (.L_HI(net246));
 sg13g2_tiehi _1482__188 (.L_HI(net247));
 sg13g2_tiehi _1481__189 (.L_HI(net248));
 sg13g2_tiehi _1480__190 (.L_HI(net249));
 sg13g2_tiehi _1479__191 (.L_HI(net250));
 sg13g2_tiehi _1478__192 (.L_HI(net251));
 sg13g2_tiehi _1477__193 (.L_HI(net252));
 sg13g2_tiehi _1476__194 (.L_HI(net253));
 sg13g2_tiehi _1475__195 (.L_HI(net254));
 sg13g2_tiehi _1474__196 (.L_HI(net255));
 sg13g2_tiehi _1473__197 (.L_HI(net256));
 sg13g2_tiehi _1472__198 (.L_HI(net257));
 sg13g2_tiehi _1471__199 (.L_HI(net258));
 sg13g2_tiehi _1470__200 (.L_HI(net259));
 sg13g2_tiehi _1469__201 (.L_HI(net260));
 sg13g2_tiehi _1468__202 (.L_HI(net261));
 sg13g2_tiehi _1467__203 (.L_HI(net262));
 sg13g2_tiehi _1466__204 (.L_HI(net263));
 sg13g2_tiehi _1465__205 (.L_HI(net264));
 sg13g2_tiehi _1464__206 (.L_HI(net265));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_dranoel06_SAP1_15 (.L_LO(net15));
 sg13g2_tielo tt_um_dranoel06_SAP1_16 (.L_LO(net16));
 sg13g2_tielo tt_um_dranoel06_SAP1_17 (.L_LO(net17));
 sg13g2_tielo tt_um_dranoel06_SAP1_18 (.L_LO(net18));
 sg13g2_tielo tt_um_dranoel06_SAP1_19 (.L_LO(net19));
 sg13g2_tielo tt_um_dranoel06_SAP1_20 (.L_LO(net20));
 sg13g2_tielo tt_um_dranoel06_SAP1_21 (.L_LO(net21));
 sg13g2_tielo tt_um_dranoel06_SAP1_22 (.L_LO(net22));
 sg13g2_tielo tt_um_dranoel06_SAP1_23 (.L_LO(net23));
 sg13g2_tielo tt_um_dranoel06_SAP1_24 (.L_LO(net24));
 sg13g2_tielo tt_um_dranoel06_SAP1_25 (.L_LO(net25));
 sg13g2_tielo tt_um_dranoel06_SAP1_26 (.L_LO(net26));
 sg13g2_tielo tt_um_dranoel06_SAP1_27 (.L_LO(net27));
 sg13g2_tielo tt_um_dranoel06_SAP1_28 (.L_LO(net28));
 sg13g2_tielo tt_um_dranoel06_SAP1_29 (.L_LO(net29));
 sg13g2_tiehi _1463__30 (.L_HI(net30));
 sg13g2_buf_8 fanout122 (.A(_0487_),
    .X(net122));
 sg13g2_buf_8 fanout123 (.A(_0487_),
    .X(net123));
 sg13g2_buf_8 fanout124 (.A(_0463_),
    .X(net124));
 sg13g2_buf_8 fanout125 (.A(_0463_),
    .X(net125));
 sg13g2_buf_8 fanout126 (.A(_0432_),
    .X(net126));
 sg13g2_buf_8 fanout127 (.A(_0432_),
    .X(net127));
 sg13g2_buf_8 fanout128 (.A(_0369_),
    .X(net128));
 sg13g2_buf_8 fanout129 (.A(_0369_),
    .X(net129));
 sg13g2_buf_8 fanout130 (.A(_0399_),
    .X(net130));
 sg13g2_buf_8 fanout131 (.A(_0399_),
    .X(net131));
 sg13g2_buf_8 fanout132 (.A(_0335_),
    .X(net132));
 sg13g2_buf_8 fanout133 (.A(_0335_),
    .X(net133));
 sg13g2_buf_8 fanout134 (.A(_0301_),
    .X(net134));
 sg13g2_buf_8 fanout135 (.A(_0301_),
    .X(net135));
 sg13g2_buf_8 fanout136 (.A(_0265_),
    .X(net136));
 sg13g2_buf_8 fanout137 (.A(_0265_),
    .X(net137));
 sg13g2_buf_8 fanout138 (.A(_0561_),
    .X(net138));
 sg13g2_buf_8 fanout139 (.A(_0509_),
    .X(net139));
 sg13g2_buf_8 fanout140 (.A(_0500_),
    .X(net140));
 sg13g2_buf_8 fanout141 (.A(net142),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_0490_),
    .X(net142));
 sg13g2_buf_8 fanout143 (.A(_0240_),
    .X(net143));
 sg13g2_buf_8 fanout144 (.A(_0259_),
    .X(net144));
 sg13g2_buf_8 fanout145 (.A(_0253_),
    .X(net145));
 sg13g2_buf_8 fanout146 (.A(net148),
    .X(net146));
 sg13g2_buf_8 fanout147 (.A(net148),
    .X(net147));
 sg13g2_buf_8 fanout148 (.A(_0203_),
    .X(net148));
 sg13g2_buf_8 fanout149 (.A(net150),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_0244_),
    .X(net150));
 sg13g2_buf_8 fanout151 (.A(_0183_),
    .X(net151));
 sg13g2_buf_1 fanout152 (.A(_0183_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(\cpu0.ir[5] ),
    .X(net153));
 sg13g2_buf_8 fanout154 (.A(net446),
    .X(net154));
 sg13g2_buf_8 fanout155 (.A(net156),
    .X(net155));
 sg13g2_buf_8 fanout156 (.A(_0003_),
    .X(net156));
 sg13g2_buf_8 fanout157 (.A(net159),
    .X(net157));
 sg13g2_buf_8 fanout158 (.A(net159),
    .X(net158));
 sg13g2_buf_8 fanout159 (.A(_0002_),
    .X(net159));
 sg13g2_buf_8 fanout160 (.A(net161),
    .X(net160));
 sg13g2_buf_8 fanout161 (.A(_0001_),
    .X(net161));
 sg13g2_buf_8 fanout162 (.A(_0001_),
    .X(net162));
 sg13g2_buf_8 fanout163 (.A(net165),
    .X(net163));
 sg13g2_buf_1 fanout164 (.A(net165),
    .X(net164));
 sg13g2_buf_8 fanout165 (.A(_0001_),
    .X(net165));
 sg13g2_buf_8 fanout166 (.A(net169),
    .X(net166));
 sg13g2_buf_1 fanout167 (.A(net169),
    .X(net167));
 sg13g2_buf_8 fanout168 (.A(net169),
    .X(net168));
 sg13g2_buf_8 fanout169 (.A(net170),
    .X(net169));
 sg13g2_buf_8 fanout170 (.A(_0000_),
    .X(net170));
 sg13g2_buf_8 fanout171 (.A(net177),
    .X(net171));
 sg13g2_buf_8 fanout172 (.A(net175),
    .X(net172));
 sg13g2_buf_1 fanout173 (.A(net175),
    .X(net173));
 sg13g2_buf_8 fanout174 (.A(net175),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(net177),
    .X(net175));
 sg13g2_buf_8 fanout176 (.A(net177),
    .X(net176));
 sg13g2_buf_8 fanout177 (.A(_0000_),
    .X(net177));
 sg13g2_buf_8 fanout178 (.A(net179),
    .X(net178));
 sg13g2_buf_8 fanout179 (.A(net180),
    .X(net179));
 sg13g2_buf_8 fanout180 (.A(rst_n),
    .X(net180));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[7]),
    .X(net13));
 sg13g2_tielo tt_um_dranoel06_SAP1_14 (.L_LO(net14));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_8 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_8 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_8 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_8 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_8 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_8 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_8 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_8 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_8 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_8 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_8 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_8 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_8 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_8 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_8 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_8 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_8 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_8 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_8 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_8 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_8 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_8 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_8 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_8 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_8 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_8 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_8 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_8 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_8 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_8 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_8 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\cpu0.ir[1] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold2 (.A(\cpu0.ir[0] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold3 (.A(\cpu0.ram[9][1] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold4 (.A(\cpu0.ir[3] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold5 (.A(\cpu0.ram[14][3] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold6 (.A(\cpu0.ir[5] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold7 (.A(\cpu0.ram[14][2] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold8 (.A(\cpu0.ram[15][1] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold9 (.A(\cpu0.ir[2] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold10 (.A(uo_out[0]),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold11 (.A(\cpu0.b_reg[2] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold12 (.A(uo_out[1]),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0100_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold14 (.A(uo_out[7]),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0106_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold16 (.A(uo_out[4]),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold17 (.A(uo_out[5]),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold18 (.A(uo_out[2]),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0101_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold20 (.A(\cpu0.a_reg[0] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold21 (.A(\cpu0.a_reg[5] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold22 (.A(\cpu0.b_reg[7] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0170_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold24 (.A(\cpu0.b_reg[1] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0164_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold26 (.A(uo_out[3]),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold27 (.A(\cpu0.b_reg[3] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold28 (.A(uo_out[6]),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold29 (.A(\cpu0.a_reg[6] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold30 (.A(\cpu0.a_reg[4] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold31 (.A(\cpu0.ram[8][3] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold32 (.A(\cpu0.ram[8][2] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold33 (.A(\cpu0.ram[4][1] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold34 (.A(\cpu0.b_reg[4] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold35 (.A(\cpu0.a_reg[1] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold36 (.A(\cpu0.ram[12][3] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold37 (.A(\cpu0.ram[13][4] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold38 (.A(\cpu0.ram[13][1] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold39 (.A(\cpu0.ram[6][2] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold40 (.A(\cpu0.b_reg[6] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold41 (.A(\cpu0.ram[12][0] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold42 (.A(\cpu0.ram[1][5] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold43 (.A(\cpu0.ram[10][1] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold44 (.A(\cpu0.ram[0][7] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold45 (.A(\cpu0.b_reg[5] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold46 (.A(\cpu0.ram[10][7] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold47 (.A(\cpu0.ram[11][0] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold48 (.A(\cpu0.ram[8][6] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold49 (.A(\cpu0.ram[3][6] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold50 (.A(\cpu0.ram[3][1] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold51 (.A(\cpu0.ram[3][3] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold52 (.A(\cpu0.ram[0][1] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold53 (.A(\cpu0.ram[12][1] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold54 (.A(\cpu0.ram[10][2] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold55 (.A(\cpu0.ram[8][1] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold56 (.A(\cpu0.ram[15][2] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold57 (.A(\cpu0.ram[9][0] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold58 (.A(\cpu0.ram[4][7] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold59 (.A(\cpu0.ram[14][6] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold60 (.A(\cpu0.ram[3][7] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold61 (.A(\cpu0.ram[4][2] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold62 (.A(\cpu0.ram[0][4] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold63 (.A(\cpu0.ram[8][7] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold64 (.A(\cpu0.ram[5][3] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold65 (.A(\cpu0.ram[8][4] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold66 (.A(\cpu0.ram[7][4] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold67 (.A(\cpu0.ram[7][7] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold68 (.A(\cpu0.ram[0][6] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold69 (.A(\cpu0.ram[13][2] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold70 (.A(\cpu0.ram[11][5] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold71 (.A(\cpu0.ram[7][6] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold72 (.A(\cpu0.ram[6][5] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold73 (.A(\cpu0.ram[14][0] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold74 (.A(\cpu0.ram[3][0] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold75 (.A(\cpu0.ram[13][0] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold76 (.A(\cpu0.ram[6][3] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold77 (.A(\cpu0.ram[5][6] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold78 (.A(\cpu0.ram[5][2] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold79 (.A(\cpu0.ram[1][0] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold80 (.A(\cpu0.ram[12][5] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold81 (.A(\cpu0.ram[2][3] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold82 (.A(\cpu0.ram[10][0] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold83 (.A(\cpu0.ram[8][0] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold84 (.A(\cpu0.ram[2][2] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold85 (.A(\cpu0.ram[14][7] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold86 (.A(\cpu0.a_reg[2] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold87 (.A(\cpu0.ram[9][6] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold88 (.A(\cpu0.ram[15][4] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold89 (.A(\cpu0.ram[11][3] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold90 (.A(\cpu0.ram[12][7] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold91 (.A(\cpu0.ram[2][5] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold92 (.A(\cpu0.ram[6][4] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold93 (.A(\cpu0.ram[9][3] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold94 (.A(\cpu0.ram[15][5] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold95 (.A(\cpu0.ram[1][7] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold96 (.A(\cpu0.ram[6][1] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold97 (.A(\cpu0.ram[4][5] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold98 (.A(\cpu0.ram[2][0] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold99 (.A(\cpu0.ram[13][3] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold100 (.A(\cpu0.ram[14][4] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold101 (.A(\cpu0.ram[13][5] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold102 (.A(\cpu0.ram[3][2] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold103 (.A(\cpu0.ram[7][1] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold104 (.A(\cpu0.ram[11][7] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold105 (.A(\cpu0.ram[10][6] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold106 (.A(\cpu0.ram[4][3] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold107 (.A(\cpu0.ram[0][2] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold108 (.A(\cpu0.ram[10][5] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold109 (.A(\cpu0.ram[7][3] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold110 (.A(\cpu0.ram[0][5] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold111 (.A(\cpu0.ram[15][3] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold112 (.A(\cpu0.ram[10][3] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold113 (.A(\cpu0.ram[2][7] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold114 (.A(\cpu0.ram[14][5] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold115 (.A(\cpu0.ram[11][1] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold116 (.A(\cpu0.ram[11][6] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold117 (.A(\cpu0.ram[11][2] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold118 (.A(\cpu0.ram[1][1] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold119 (.A(\cpu0.ram[6][6] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold120 (.A(\cpu0.ram[13][6] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold121 (.A(\cpu0.ram[2][1] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold122 (.A(\cpu0.ram[12][2] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold123 (.A(\cpu0.ram[3][5] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold124 (.A(\cpu0.ram[9][4] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold125 (.A(\cpu0.ram[5][7] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold126 (.A(\cpu0.ram[9][5] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold127 (.A(\cpu0.ram[7][0] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold128 (.A(\cpu0.ram[12][6] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold129 (.A(\cpu0.ram[1][3] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold130 (.A(\cpu0.ram[7][5] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold131 (.A(\cpu0.ram[4][6] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold132 (.A(\cpu0.ram[7][2] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold133 (.A(\cpu0.ram[5][5] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold134 (.A(\cpu0.b_reg[0] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0163_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold136 (.A(\cpu0.ram[3][4] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold137 (.A(\cpu0.ram[11][4] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold138 (.A(\cpu0.ram[14][1] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold139 (.A(\cpu0.ram[13][7] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold140 (.A(\cpu0.ram[0][0] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold141 (.A(\cpu0.ram[15][0] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold142 (.A(\cpu0.ram[4][0] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold143 (.A(\cpu0.ram[4][4] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold144 (.A(\cpu0.ram[2][6] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold145 (.A(\cpu0.ram[9][7] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold146 (.A(\cpu0.ram[5][1] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold147 (.A(\cpu0.ram[15][6] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold148 (.A(\cpu0.ram[1][4] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold149 (.A(\cpu0.ram[6][7] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold150 (.A(\cpu0.ram[2][4] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold151 (.A(\cpu0.ram[9][2] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold152 (.A(\cpu0.ram[12][4] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold153 (.A(\cpu0.ram[6][0] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold154 (.A(\cpu0.ram[8][5] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold155 (.A(\cpu0.ram[0][3] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold156 (.A(\cpu0.ram[15][7] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold157 (.A(\cpu0.ram[5][4] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold158 (.A(\cpu0.ram[1][6] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold159 (.A(\cpu0.a_reg[7] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold160 (.A(\cpu0.a_reg[3] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold161 (.A(\cpu0.ram[10][4] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold162 (.A(\cpu0.ram[1][2] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold163 (.A(\cpu0.ram[5][0] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold164 (.A(\cpu0.ir[6] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold165 (.A(\cpu0.carry_flag ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0172_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold167 (.A(\cpu0.step[1] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0503_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold169 (.A(\cpu0.ir[4] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold170 (.A(\cpu0.ir[7] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold171 (.A(\cpu0.zero_flag ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold172 (.A(\cpu0.step[0] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold173 (.A(\cpu0.mar[2] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold174 (.A(\cpu0.mar[3] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold175 (.A(\cpu0.mar[1] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold176 (.A(\cpu0.pc[2] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold177 (.A(\cpu0.pc[1] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold178 (.A(\cpu0.mar[0] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold179 (.A(\cpu0.pc[0] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold180 (.A(\cpu0.pc[3] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold181 (.A(\cpu0.step[2] ),
    .X(net446));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_4 FILLER_0_84 ();
 sg13g2_fill_1 FILLER_0_88 ();
 sg13g2_decap_8 FILLER_0_102 ();
 sg13g2_decap_8 FILLER_0_109 ();
 sg13g2_decap_8 FILLER_0_116 ();
 sg13g2_decap_8 FILLER_0_123 ();
 sg13g2_decap_8 FILLER_0_130 ();
 sg13g2_decap_8 FILLER_0_137 ();
 sg13g2_fill_2 FILLER_0_144 ();
 sg13g2_fill_1 FILLER_0_146 ();
 sg13g2_decap_8 FILLER_0_156 ();
 sg13g2_decap_8 FILLER_0_172 ();
 sg13g2_decap_8 FILLER_0_179 ();
 sg13g2_decap_8 FILLER_0_186 ();
 sg13g2_decap_8 FILLER_0_193 ();
 sg13g2_fill_2 FILLER_0_200 ();
 sg13g2_fill_2 FILLER_0_215 ();
 sg13g2_fill_1 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_228 ();
 sg13g2_decap_8 FILLER_0_235 ();
 sg13g2_decap_8 FILLER_0_242 ();
 sg13g2_decap_8 FILLER_0_249 ();
 sg13g2_decap_8 FILLER_0_256 ();
 sg13g2_fill_2 FILLER_0_263 ();
 sg13g2_decap_8 FILLER_0_274 ();
 sg13g2_decap_8 FILLER_0_281 ();
 sg13g2_decap_4 FILLER_0_288 ();
 sg13g2_fill_2 FILLER_0_292 ();
 sg13g2_decap_8 FILLER_0_298 ();
 sg13g2_decap_8 FILLER_0_305 ();
 sg13g2_decap_8 FILLER_0_312 ();
 sg13g2_decap_8 FILLER_0_319 ();
 sg13g2_decap_8 FILLER_0_326 ();
 sg13g2_decap_8 FILLER_0_360 ();
 sg13g2_decap_8 FILLER_0_367 ();
 sg13g2_decap_4 FILLER_0_374 ();
 sg13g2_fill_2 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_383 ();
 sg13g2_decap_8 FILLER_0_390 ();
 sg13g2_decap_8 FILLER_0_397 ();
 sg13g2_decap_4 FILLER_0_404 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_4 FILLER_1_77 ();
 sg13g2_fill_2 FILLER_1_81 ();
 sg13g2_decap_8 FILLER_1_114 ();
 sg13g2_decap_8 FILLER_1_121 ();
 sg13g2_fill_2 FILLER_1_128 ();
 sg13g2_fill_1 FILLER_1_130 ();
 sg13g2_fill_2 FILLER_1_135 ();
 sg13g2_decap_8 FILLER_1_178 ();
 sg13g2_decap_4 FILLER_1_185 ();
 sg13g2_decap_8 FILLER_1_199 ();
 sg13g2_decap_8 FILLER_1_242 ();
 sg13g2_decap_4 FILLER_1_249 ();
 sg13g2_fill_2 FILLER_1_253 ();
 sg13g2_decap_4 FILLER_1_282 ();
 sg13g2_fill_1 FILLER_1_286 ();
 sg13g2_fill_2 FILLER_1_314 ();
 sg13g2_decap_8 FILLER_1_319 ();
 sg13g2_fill_2 FILLER_1_326 ();
 sg13g2_fill_2 FILLER_1_364 ();
 sg13g2_fill_1 FILLER_1_366 ();
 sg13g2_decap_4 FILLER_1_403 ();
 sg13g2_fill_2 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_62 ();
 sg13g2_decap_4 FILLER_2_69 ();
 sg13g2_fill_1 FILLER_2_73 ();
 sg13g2_decap_8 FILLER_2_115 ();
 sg13g2_fill_2 FILLER_2_242 ();
 sg13g2_fill_1 FILLER_2_244 ();
 sg13g2_fill_2 FILLER_2_282 ();
 sg13g2_fill_2 FILLER_2_325 ();
 sg13g2_decap_4 FILLER_2_356 ();
 sg13g2_decap_8 FILLER_2_400 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_fill_2 FILLER_3_28 ();
 sg13g2_fill_2 FILLER_3_50 ();
 sg13g2_fill_1 FILLER_3_52 ();
 sg13g2_decap_8 FILLER_3_62 ();
 sg13g2_decap_8 FILLER_3_69 ();
 sg13g2_fill_1 FILLER_3_76 ();
 sg13g2_fill_1 FILLER_3_104 ();
 sg13g2_decap_4 FILLER_3_195 ();
 sg13g2_fill_1 FILLER_3_199 ();
 sg13g2_decap_4 FILLER_3_251 ();
 sg13g2_fill_1 FILLER_3_288 ();
 sg13g2_fill_1 FILLER_3_313 ();
 sg13g2_fill_1 FILLER_3_337 ();
 sg13g2_fill_2 FILLER_3_356 ();
 sg13g2_fill_1 FILLER_3_366 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_4 FILLER_4_7 ();
 sg13g2_fill_2 FILLER_4_11 ();
 sg13g2_decap_8 FILLER_4_53 ();
 sg13g2_decap_8 FILLER_4_60 ();
 sg13g2_decap_4 FILLER_4_67 ();
 sg13g2_fill_2 FILLER_4_71 ();
 sg13g2_fill_2 FILLER_4_100 ();
 sg13g2_fill_1 FILLER_4_102 ();
 sg13g2_decap_8 FILLER_4_121 ();
 sg13g2_decap_4 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_241 ();
 sg13g2_decap_8 FILLER_4_248 ();
 sg13g2_decap_4 FILLER_4_255 ();
 sg13g2_fill_1 FILLER_4_259 ();
 sg13g2_fill_2 FILLER_4_271 ();
 sg13g2_fill_2 FILLER_4_286 ();
 sg13g2_fill_2 FILLER_4_301 ();
 sg13g2_fill_1 FILLER_4_303 ();
 sg13g2_decap_4 FILLER_4_309 ();
 sg13g2_fill_2 FILLER_4_358 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_57 ();
 sg13g2_decap_8 FILLER_5_64 ();
 sg13g2_fill_2 FILLER_5_71 ();
 sg13g2_fill_1 FILLER_5_73 ();
 sg13g2_fill_2 FILLER_5_88 ();
 sg13g2_decap_4 FILLER_5_124 ();
 sg13g2_fill_2 FILLER_5_128 ();
 sg13g2_fill_2 FILLER_5_205 ();
 sg13g2_fill_2 FILLER_5_243 ();
 sg13g2_fill_2 FILLER_5_257 ();
 sg13g2_fill_1 FILLER_5_259 ();
 sg13g2_fill_1 FILLER_5_265 ();
 sg13g2_fill_1 FILLER_5_293 ();
 sg13g2_fill_1 FILLER_5_299 ();
 sg13g2_decap_8 FILLER_5_305 ();
 sg13g2_fill_2 FILLER_5_312 ();
 sg13g2_fill_1 FILLER_5_314 ();
 sg13g2_fill_1 FILLER_5_347 ();
 sg13g2_fill_2 FILLER_5_353 ();
 sg13g2_fill_2 FILLER_5_365 ();
 sg13g2_decap_4 FILLER_5_404 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_7 ();
 sg13g2_decap_4 FILLER_6_64 ();
 sg13g2_fill_2 FILLER_6_68 ();
 sg13g2_fill_2 FILLER_6_83 ();
 sg13g2_fill_1 FILLER_6_85 ();
 sg13g2_decap_8 FILLER_6_127 ();
 sg13g2_decap_4 FILLER_6_134 ();
 sg13g2_fill_2 FILLER_6_175 ();
 sg13g2_decap_4 FILLER_6_218 ();
 sg13g2_fill_2 FILLER_6_253 ();
 sg13g2_fill_2 FILLER_6_260 ();
 sg13g2_fill_2 FILLER_6_330 ();
 sg13g2_fill_1 FILLER_6_332 ();
 sg13g2_decap_8 FILLER_6_362 ();
 sg13g2_decap_8 FILLER_6_369 ();
 sg13g2_decap_4 FILLER_6_376 ();
 sg13g2_fill_2 FILLER_6_380 ();
 sg13g2_decap_4 FILLER_6_404 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_fill_2 FILLER_7_14 ();
 sg13g2_decap_4 FILLER_7_58 ();
 sg13g2_fill_1 FILLER_7_62 ();
 sg13g2_decap_4 FILLER_7_122 ();
 sg13g2_fill_1 FILLER_7_126 ();
 sg13g2_fill_1 FILLER_7_181 ();
 sg13g2_decap_8 FILLER_7_219 ();
 sg13g2_fill_2 FILLER_7_226 ();
 sg13g2_fill_1 FILLER_7_228 ();
 sg13g2_fill_2 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_323 ();
 sg13g2_decap_4 FILLER_7_330 ();
 sg13g2_fill_2 FILLER_7_347 ();
 sg13g2_fill_1 FILLER_7_349 ();
 sg13g2_fill_2 FILLER_7_363 ();
 sg13g2_fill_1 FILLER_7_365 ();
 sg13g2_decap_4 FILLER_7_403 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_4 FILLER_8_7 ();
 sg13g2_fill_1 FILLER_8_11 ();
 sg13g2_fill_1 FILLER_8_39 ();
 sg13g2_decap_4 FILLER_8_55 ();
 sg13g2_decap_8 FILLER_8_128 ();
 sg13g2_fill_2 FILLER_8_139 ();
 sg13g2_fill_2 FILLER_8_183 ();
 sg13g2_fill_2 FILLER_8_200 ();
 sg13g2_fill_1 FILLER_8_202 ();
 sg13g2_decap_8 FILLER_8_220 ();
 sg13g2_fill_2 FILLER_8_227 ();
 sg13g2_fill_1 FILLER_8_229 ();
 sg13g2_fill_2 FILLER_8_243 ();
 sg13g2_decap_8 FILLER_8_275 ();
 sg13g2_fill_1 FILLER_8_282 ();
 sg13g2_decap_4 FILLER_8_329 ();
 sg13g2_fill_1 FILLER_8_333 ();
 sg13g2_decap_4 FILLER_8_360 ();
 sg13g2_decap_8 FILLER_8_401 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_7 ();
 sg13g2_decap_4 FILLER_9_62 ();
 sg13g2_fill_1 FILLER_9_66 ();
 sg13g2_fill_1 FILLER_9_81 ();
 sg13g2_fill_2 FILLER_9_110 ();
 sg13g2_fill_1 FILLER_9_112 ();
 sg13g2_decap_4 FILLER_9_122 ();
 sg13g2_fill_2 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_141 ();
 sg13g2_fill_1 FILLER_9_148 ();
 sg13g2_decap_8 FILLER_9_177 ();
 sg13g2_decap_8 FILLER_9_184 ();
 sg13g2_fill_2 FILLER_9_207 ();
 sg13g2_fill_1 FILLER_9_209 ();
 sg13g2_decap_8 FILLER_9_219 ();
 sg13g2_decap_8 FILLER_9_226 ();
 sg13g2_decap_4 FILLER_9_233 ();
 sg13g2_fill_2 FILLER_9_237 ();
 sg13g2_decap_8 FILLER_9_271 ();
 sg13g2_decap_8 FILLER_9_278 ();
 sg13g2_fill_1 FILLER_9_285 ();
 sg13g2_fill_1 FILLER_9_332 ();
 sg13g2_fill_2 FILLER_9_369 ();
 sg13g2_fill_1 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_7 ();
 sg13g2_fill_2 FILLER_10_47 ();
 sg13g2_fill_1 FILLER_10_57 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_fill_1 FILLER_10_70 ();
 sg13g2_fill_2 FILLER_10_81 ();
 sg13g2_fill_1 FILLER_10_92 ();
 sg13g2_fill_2 FILLER_10_102 ();
 sg13g2_fill_1 FILLER_10_104 ();
 sg13g2_decap_4 FILLER_10_124 ();
 sg13g2_fill_2 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_187 ();
 sg13g2_fill_1 FILLER_10_194 ();
 sg13g2_fill_1 FILLER_10_236 ();
 sg13g2_fill_1 FILLER_10_249 ();
 sg13g2_decap_8 FILLER_10_272 ();
 sg13g2_fill_2 FILLER_10_279 ();
 sg13g2_fill_2 FILLER_10_295 ();
 sg13g2_fill_1 FILLER_10_297 ();
 sg13g2_decap_4 FILLER_10_339 ();
 sg13g2_fill_2 FILLER_10_355 ();
 sg13g2_fill_1 FILLER_10_357 ();
 sg13g2_decap_4 FILLER_10_368 ();
 sg13g2_fill_2 FILLER_10_372 ();
 sg13g2_decap_4 FILLER_10_404 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_fill_2 FILLER_11_14 ();
 sg13g2_fill_1 FILLER_11_20 ();
 sg13g2_fill_1 FILLER_11_58 ();
 sg13g2_fill_1 FILLER_11_72 ();
 sg13g2_fill_2 FILLER_11_100 ();
 sg13g2_fill_1 FILLER_11_102 ();
 sg13g2_decap_8 FILLER_11_130 ();
 sg13g2_fill_2 FILLER_11_137 ();
 sg13g2_fill_1 FILLER_11_139 ();
 sg13g2_fill_1 FILLER_11_281 ();
 sg13g2_fill_2 FILLER_11_314 ();
 sg13g2_fill_1 FILLER_11_316 ();
 sg13g2_fill_2 FILLER_11_331 ();
 sg13g2_fill_1 FILLER_11_333 ();
 sg13g2_fill_2 FILLER_11_361 ();
 sg13g2_decap_4 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_fill_1 FILLER_12_21 ();
 sg13g2_fill_1 FILLER_12_31 ();
 sg13g2_fill_2 FILLER_12_68 ();
 sg13g2_fill_2 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_234 ();
 sg13g2_decap_4 FILLER_12_241 ();
 sg13g2_fill_2 FILLER_12_245 ();
 sg13g2_fill_2 FILLER_12_297 ();
 sg13g2_fill_1 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_353 ();
 sg13g2_decap_4 FILLER_12_360 ();
 sg13g2_fill_1 FILLER_12_364 ();
 sg13g2_fill_2 FILLER_12_379 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_7 ();
 sg13g2_fill_1 FILLER_13_36 ();
 sg13g2_fill_1 FILLER_13_55 ();
 sg13g2_fill_1 FILLER_13_73 ();
 sg13g2_fill_2 FILLER_13_88 ();
 sg13g2_decap_8 FILLER_13_137 ();
 sg13g2_decap_4 FILLER_13_144 ();
 sg13g2_fill_2 FILLER_13_152 ();
 sg13g2_fill_1 FILLER_13_154 ();
 sg13g2_decap_4 FILLER_13_165 ();
 sg13g2_fill_2 FILLER_13_195 ();
 sg13g2_decap_8 FILLER_13_234 ();
 sg13g2_decap_4 FILLER_13_241 ();
 sg13g2_fill_2 FILLER_13_269 ();
 sg13g2_decap_8 FILLER_13_284 ();
 sg13g2_decap_8 FILLER_13_291 ();
 sg13g2_fill_2 FILLER_13_303 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_fill_1 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_decap_4 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_66 ();
 sg13g2_fill_2 FILLER_14_90 ();
 sg13g2_decap_8 FILLER_14_137 ();
 sg13g2_fill_1 FILLER_14_144 ();
 sg13g2_decap_8 FILLER_14_149 ();
 sg13g2_decap_4 FILLER_14_156 ();
 sg13g2_fill_2 FILLER_14_160 ();
 sg13g2_fill_1 FILLER_14_172 ();
 sg13g2_fill_2 FILLER_14_200 ();
 sg13g2_fill_1 FILLER_14_202 ();
 sg13g2_decap_8 FILLER_14_221 ();
 sg13g2_decap_8 FILLER_14_228 ();
 sg13g2_decap_4 FILLER_14_235 ();
 sg13g2_fill_2 FILLER_14_239 ();
 sg13g2_decap_4 FILLER_14_251 ();
 sg13g2_fill_1 FILLER_14_264 ();
 sg13g2_fill_1 FILLER_14_274 ();
 sg13g2_decap_8 FILLER_14_284 ();
 sg13g2_decap_8 FILLER_14_291 ();
 sg13g2_fill_1 FILLER_14_298 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_fill_2 FILLER_14_329 ();
 sg13g2_decap_4 FILLER_14_338 ();
 sg13g2_decap_8 FILLER_14_351 ();
 sg13g2_fill_1 FILLER_14_358 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_4 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_51 ();
 sg13g2_fill_1 FILLER_15_79 ();
 sg13g2_fill_2 FILLER_15_84 ();
 sg13g2_fill_2 FILLER_15_92 ();
 sg13g2_decap_8 FILLER_15_138 ();
 sg13g2_decap_4 FILLER_15_145 ();
 sg13g2_fill_1 FILLER_15_149 ();
 sg13g2_decap_4 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_214 ();
 sg13g2_decap_8 FILLER_15_221 ();
 sg13g2_decap_4 FILLER_15_228 ();
 sg13g2_fill_2 FILLER_15_232 ();
 sg13g2_decap_4 FILLER_15_265 ();
 sg13g2_fill_2 FILLER_15_289 ();
 sg13g2_fill_1 FILLER_15_291 ();
 sg13g2_decap_4 FILLER_15_361 ();
 sg13g2_fill_2 FILLER_15_397 ();
 sg13g2_fill_1 FILLER_15_399 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_4 ();
 sg13g2_fill_1 FILLER_16_63 ();
 sg13g2_decap_4 FILLER_16_69 ();
 sg13g2_fill_2 FILLER_16_73 ();
 sg13g2_decap_4 FILLER_16_80 ();
 sg13g2_fill_1 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_145 ();
 sg13g2_decap_4 FILLER_16_152 ();
 sg13g2_fill_1 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_220 ();
 sg13g2_decap_4 FILLER_16_227 ();
 sg13g2_decap_4 FILLER_16_272 ();
 sg13g2_fill_2 FILLER_16_276 ();
 sg13g2_fill_2 FILLER_16_339 ();
 sg13g2_fill_1 FILLER_16_341 ();
 sg13g2_decap_4 FILLER_16_369 ();
 sg13g2_decap_4 FILLER_16_404 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_47 ();
 sg13g2_decap_4 FILLER_17_54 ();
 sg13g2_fill_1 FILLER_17_58 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_4 FILLER_17_168 ();
 sg13g2_fill_2 FILLER_17_172 ();
 sg13g2_decap_8 FILLER_17_216 ();
 sg13g2_decap_4 FILLER_17_223 ();
 sg13g2_fill_1 FILLER_17_227 ();
 sg13g2_fill_2 FILLER_17_291 ();
 sg13g2_decap_8 FILLER_17_320 ();
 sg13g2_decap_8 FILLER_17_358 ();
 sg13g2_fill_1 FILLER_17_365 ();
 sg13g2_decap_4 FILLER_17_403 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_decap_4 FILLER_18_59 ();
 sg13g2_fill_1 FILLER_18_63 ();
 sg13g2_fill_2 FILLER_18_114 ();
 sg13g2_fill_1 FILLER_18_116 ();
 sg13g2_fill_1 FILLER_18_122 ();
 sg13g2_decap_8 FILLER_18_142 ();
 sg13g2_decap_8 FILLER_18_149 ();
 sg13g2_decap_8 FILLER_18_156 ();
 sg13g2_decap_8 FILLER_18_163 ();
 sg13g2_fill_1 FILLER_18_175 ();
 sg13g2_fill_1 FILLER_18_204 ();
 sg13g2_decap_8 FILLER_18_214 ();
 sg13g2_decap_8 FILLER_18_221 ();
 sg13g2_fill_2 FILLER_18_245 ();
 sg13g2_fill_1 FILLER_18_276 ();
 sg13g2_decap_4 FILLER_18_286 ();
 sg13g2_fill_1 FILLER_18_290 ();
 sg13g2_fill_2 FILLER_18_295 ();
 sg13g2_fill_1 FILLER_18_297 ();
 sg13g2_decap_4 FILLER_18_311 ();
 sg13g2_fill_1 FILLER_18_315 ();
 sg13g2_decap_4 FILLER_18_329 ();
 sg13g2_fill_1 FILLER_18_333 ();
 sg13g2_fill_1 FILLER_18_366 ();
 sg13g2_decap_4 FILLER_18_377 ();
 sg13g2_fill_1 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_4 FILLER_19_54 ();
 sg13g2_fill_2 FILLER_19_58 ();
 sg13g2_fill_2 FILLER_19_86 ();
 sg13g2_fill_1 FILLER_19_88 ();
 sg13g2_fill_2 FILLER_19_108 ();
 sg13g2_fill_1 FILLER_19_110 ();
 sg13g2_decap_8 FILLER_19_129 ();
 sg13g2_decap_8 FILLER_19_136 ();
 sg13g2_decap_8 FILLER_19_143 ();
 sg13g2_fill_2 FILLER_19_176 ();
 sg13g2_decap_4 FILLER_19_199 ();
 sg13g2_fill_1 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_208 ();
 sg13g2_fill_2 FILLER_19_215 ();
 sg13g2_decap_4 FILLER_19_221 ();
 sg13g2_fill_1 FILLER_19_225 ();
 sg13g2_decap_4 FILLER_19_239 ();
 sg13g2_fill_1 FILLER_19_253 ();
 sg13g2_decap_4 FILLER_19_269 ();
 sg13g2_fill_2 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_302 ();
 sg13g2_decap_8 FILLER_19_309 ();
 sg13g2_fill_1 FILLER_19_356 ();
 sg13g2_decap_8 FILLER_19_361 ();
 sg13g2_decap_4 FILLER_19_380 ();
 sg13g2_fill_1 FILLER_19_384 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_4 FILLER_19_403 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_47 ();
 sg13g2_decap_8 FILLER_20_62 ();
 sg13g2_fill_2 FILLER_20_69 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_fill_1 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_104 ();
 sg13g2_fill_2 FILLER_20_120 ();
 sg13g2_fill_1 FILLER_20_122 ();
 sg13g2_decap_4 FILLER_20_136 ();
 sg13g2_fill_2 FILLER_20_158 ();
 sg13g2_fill_1 FILLER_20_160 ();
 sg13g2_decap_8 FILLER_20_193 ();
 sg13g2_decap_8 FILLER_20_200 ();
 sg13g2_fill_1 FILLER_20_220 ();
 sg13g2_fill_2 FILLER_20_263 ();
 sg13g2_fill_1 FILLER_20_265 ();
 sg13g2_decap_8 FILLER_20_305 ();
 sg13g2_decap_4 FILLER_20_312 ();
 sg13g2_fill_2 FILLER_20_316 ();
 sg13g2_decap_4 FILLER_20_335 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_4 FILLER_20_357 ();
 sg13g2_fill_1 FILLER_20_361 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_4 FILLER_21_7 ();
 sg13g2_fill_1 FILLER_21_11 ();
 sg13g2_decap_8 FILLER_21_53 ();
 sg13g2_fill_2 FILLER_21_60 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_fill_2 FILLER_21_135 ();
 sg13g2_decap_8 FILLER_21_150 ();
 sg13g2_fill_2 FILLER_21_157 ();
 sg13g2_decap_8 FILLER_21_195 ();
 sg13g2_decap_8 FILLER_21_202 ();
 sg13g2_decap_4 FILLER_21_209 ();
 sg13g2_fill_2 FILLER_21_249 ();
 sg13g2_fill_1 FILLER_21_251 ();
 sg13g2_fill_1 FILLER_21_265 ();
 sg13g2_decap_8 FILLER_21_311 ();
 sg13g2_decap_8 FILLER_21_318 ();
 sg13g2_decap_8 FILLER_21_325 ();
 sg13g2_fill_2 FILLER_21_332 ();
 sg13g2_fill_1 FILLER_21_334 ();
 sg13g2_decap_8 FILLER_21_340 ();
 sg13g2_decap_4 FILLER_21_347 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_fill_1 FILLER_22_31 ();
 sg13g2_decap_8 FILLER_22_41 ();
 sg13g2_decap_8 FILLER_22_48 ();
 sg13g2_decap_8 FILLER_22_55 ();
 sg13g2_fill_2 FILLER_22_62 ();
 sg13g2_decap_8 FILLER_22_101 ();
 sg13g2_fill_1 FILLER_22_108 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_fill_2 FILLER_22_147 ();
 sg13g2_fill_1 FILLER_22_149 ();
 sg13g2_decap_4 FILLER_22_203 ();
 sg13g2_fill_2 FILLER_22_207 ();
 sg13g2_fill_2 FILLER_22_246 ();
 sg13g2_decap_4 FILLER_22_308 ();
 sg13g2_fill_2 FILLER_22_312 ();
 sg13g2_fill_2 FILLER_22_357 ();
 sg13g2_fill_1 FILLER_22_359 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_4 FILLER_23_14 ();
 sg13g2_fill_2 FILLER_23_18 ();
 sg13g2_decap_8 FILLER_23_40 ();
 sg13g2_decap_8 FILLER_23_47 ();
 sg13g2_decap_4 FILLER_23_54 ();
 sg13g2_fill_1 FILLER_23_58 ();
 sg13g2_decap_8 FILLER_23_104 ();
 sg13g2_decap_4 FILLER_23_111 ();
 sg13g2_decap_8 FILLER_23_136 ();
 sg13g2_decap_8 FILLER_23_143 ();
 sg13g2_decap_4 FILLER_23_150 ();
 sg13g2_fill_1 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_198 ();
 sg13g2_fill_1 FILLER_23_236 ();
 sg13g2_decap_4 FILLER_23_259 ();
 sg13g2_fill_1 FILLER_23_263 ();
 sg13g2_fill_2 FILLER_23_268 ();
 sg13g2_fill_1 FILLER_23_270 ();
 sg13g2_decap_4 FILLER_23_275 ();
 sg13g2_fill_2 FILLER_23_279 ();
 sg13g2_fill_2 FILLER_23_285 ();
 sg13g2_decap_8 FILLER_23_296 ();
 sg13g2_decap_4 FILLER_23_303 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_4 FILLER_24_7 ();
 sg13g2_fill_1 FILLER_24_59 ();
 sg13g2_decap_8 FILLER_24_104 ();
 sg13g2_decap_4 FILLER_24_111 ();
 sg13g2_fill_2 FILLER_24_115 ();
 sg13g2_fill_1 FILLER_24_127 ();
 sg13g2_decap_8 FILLER_24_149 ();
 sg13g2_decap_8 FILLER_24_156 ();
 sg13g2_fill_1 FILLER_24_163 ();
 sg13g2_decap_8 FILLER_24_193 ();
 sg13g2_decap_8 FILLER_24_200 ();
 sg13g2_decap_4 FILLER_24_207 ();
 sg13g2_fill_1 FILLER_24_211 ();
 sg13g2_fill_1 FILLER_24_249 ();
 sg13g2_decap_4 FILLER_24_255 ();
 sg13g2_fill_1 FILLER_24_259 ();
 sg13g2_fill_2 FILLER_24_265 ();
 sg13g2_fill_1 FILLER_24_267 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_fill_2 FILLER_24_349 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_fill_1 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_59 ();
 sg13g2_decap_4 FILLER_25_102 ();
 sg13g2_fill_2 FILLER_25_106 ();
 sg13g2_decap_8 FILLER_25_149 ();
 sg13g2_decap_8 FILLER_25_156 ();
 sg13g2_decap_8 FILLER_25_163 ();
 sg13g2_fill_1 FILLER_25_170 ();
 sg13g2_fill_1 FILLER_25_183 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_4 FILLER_25_217 ();
 sg13g2_fill_2 FILLER_25_221 ();
 sg13g2_decap_8 FILLER_25_232 ();
 sg13g2_fill_2 FILLER_25_239 ();
 sg13g2_decap_4 FILLER_25_249 ();
 sg13g2_fill_2 FILLER_25_253 ();
 sg13g2_decap_8 FILLER_25_305 ();
 sg13g2_fill_2 FILLER_25_312 ();
 sg13g2_fill_1 FILLER_25_314 ();
 sg13g2_fill_2 FILLER_25_329 ();
 sg13g2_fill_1 FILLER_25_331 ();
 sg13g2_fill_1 FILLER_25_337 ();
 sg13g2_fill_1 FILLER_25_352 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_4 ();
 sg13g2_decap_8 FILLER_26_54 ();
 sg13g2_decap_8 FILLER_26_61 ();
 sg13g2_fill_2 FILLER_26_68 ();
 sg13g2_decap_8 FILLER_26_93 ();
 sg13g2_decap_4 FILLER_26_165 ();
 sg13g2_fill_1 FILLER_26_169 ();
 sg13g2_fill_2 FILLER_26_198 ();
 sg13g2_decap_8 FILLER_26_204 ();
 sg13g2_decap_8 FILLER_26_211 ();
 sg13g2_fill_1 FILLER_26_218 ();
 sg13g2_decap_8 FILLER_26_236 ();
 sg13g2_decap_8 FILLER_26_243 ();
 sg13g2_decap_4 FILLER_26_250 ();
 sg13g2_fill_1 FILLER_26_282 ();
 sg13g2_fill_2 FILLER_26_305 ();
 sg13g2_decap_8 FILLER_26_313 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_4 FILLER_27_56 ();
 sg13g2_fill_1 FILLER_27_60 ();
 sg13g2_fill_2 FILLER_27_65 ();
 sg13g2_fill_2 FILLER_27_90 ();
 sg13g2_fill_1 FILLER_27_92 ();
 sg13g2_fill_2 FILLER_27_113 ();
 sg13g2_fill_1 FILLER_27_115 ();
 sg13g2_decap_8 FILLER_27_152 ();
 sg13g2_decap_8 FILLER_27_159 ();
 sg13g2_fill_1 FILLER_27_166 ();
 sg13g2_fill_1 FILLER_27_209 ();
 sg13g2_decap_8 FILLER_27_243 ();
 sg13g2_decap_8 FILLER_27_250 ();
 sg13g2_fill_2 FILLER_27_257 ();
 sg13g2_fill_2 FILLER_27_263 ();
 sg13g2_decap_4 FILLER_27_324 ();
 sg13g2_fill_2 FILLER_27_338 ();
 sg13g2_fill_1 FILLER_27_373 ();
 sg13g2_decap_8 FILLER_27_396 ();
 sg13g2_decap_4 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_14 ();
 sg13g2_fill_1 FILLER_28_64 ();
 sg13g2_decap_8 FILLER_28_92 ();
 sg13g2_decap_4 FILLER_28_99 ();
 sg13g2_fill_1 FILLER_28_103 ();
 sg13g2_fill_1 FILLER_28_114 ();
 sg13g2_decap_8 FILLER_28_142 ();
 sg13g2_decap_8 FILLER_28_149 ();
 sg13g2_fill_2 FILLER_28_156 ();
 sg13g2_fill_1 FILLER_28_189 ();
 sg13g2_fill_2 FILLER_28_203 ();
 sg13g2_fill_1 FILLER_28_205 ();
 sg13g2_fill_2 FILLER_28_214 ();
 sg13g2_fill_1 FILLER_28_216 ();
 sg13g2_decap_8 FILLER_28_248 ();
 sg13g2_decap_8 FILLER_28_255 ();
 sg13g2_fill_1 FILLER_28_262 ();
 sg13g2_fill_2 FILLER_28_272 ();
 sg13g2_fill_1 FILLER_28_274 ();
 sg13g2_decap_8 FILLER_28_328 ();
 sg13g2_fill_2 FILLER_28_335 ();
 sg13g2_fill_1 FILLER_28_337 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_7 ();
 sg13g2_decap_4 FILLER_29_45 ();
 sg13g2_fill_2 FILLER_29_49 ();
 sg13g2_fill_2 FILLER_29_112 ();
 sg13g2_fill_1 FILLER_29_114 ();
 sg13g2_decap_8 FILLER_29_150 ();
 sg13g2_decap_8 FILLER_29_157 ();
 sg13g2_fill_1 FILLER_29_164 ();
 sg13g2_fill_1 FILLER_29_220 ();
 sg13g2_decap_8 FILLER_29_245 ();
 sg13g2_decap_4 FILLER_29_252 ();
 sg13g2_fill_1 FILLER_29_310 ();
 sg13g2_decap_8 FILLER_29_319 ();
 sg13g2_decap_8 FILLER_29_326 ();
 sg13g2_decap_8 FILLER_29_333 ();
 sg13g2_decap_4 FILLER_29_340 ();
 sg13g2_fill_2 FILLER_29_344 ();
 sg13g2_fill_2 FILLER_29_360 ();
 sg13g2_fill_1 FILLER_29_362 ();
 sg13g2_fill_2 FILLER_29_369 ();
 sg13g2_fill_1 FILLER_29_371 ();
 sg13g2_fill_1 FILLER_29_379 ();
 sg13g2_decap_4 FILLER_29_393 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_fill_2 FILLER_30_60 ();
 sg13g2_decap_4 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_137 ();
 sg13g2_decap_4 FILLER_30_144 ();
 sg13g2_fill_2 FILLER_30_148 ();
 sg13g2_fill_2 FILLER_30_191 ();
 sg13g2_decap_8 FILLER_30_236 ();
 sg13g2_decap_8 FILLER_30_243 ();
 sg13g2_fill_2 FILLER_30_250 ();
 sg13g2_fill_1 FILLER_30_252 ();
 sg13g2_fill_2 FILLER_30_312 ();
 sg13g2_fill_1 FILLER_30_326 ();
 sg13g2_fill_2 FILLER_30_361 ();
 sg13g2_fill_1 FILLER_30_363 ();
 sg13g2_fill_2 FILLER_30_387 ();
 sg13g2_decap_8 FILLER_30_402 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_50 ();
 sg13g2_decap_8 FILLER_31_57 ();
 sg13g2_fill_1 FILLER_31_81 ();
 sg13g2_decap_8 FILLER_31_101 ();
 sg13g2_decap_4 FILLER_31_145 ();
 sg13g2_fill_1 FILLER_31_149 ();
 sg13g2_fill_2 FILLER_31_163 ();
 sg13g2_fill_1 FILLER_31_165 ();
 sg13g2_decap_8 FILLER_31_174 ();
 sg13g2_decap_8 FILLER_31_181 ();
 sg13g2_fill_2 FILLER_31_188 ();
 sg13g2_fill_1 FILLER_31_190 ();
 sg13g2_fill_2 FILLER_31_211 ();
 sg13g2_decap_8 FILLER_31_239 ();
 sg13g2_decap_8 FILLER_31_246 ();
 sg13g2_decap_8 FILLER_31_253 ();
 sg13g2_fill_1 FILLER_31_260 ();
 sg13g2_decap_4 FILLER_31_266 ();
 sg13g2_fill_1 FILLER_31_285 ();
 sg13g2_decap_8 FILLER_31_291 ();
 sg13g2_decap_8 FILLER_31_310 ();
 sg13g2_fill_1 FILLER_31_321 ();
 sg13g2_fill_2 FILLER_31_334 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_4 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_11 ();
 sg13g2_decap_8 FILLER_32_52 ();
 sg13g2_fill_2 FILLER_32_59 ();
 sg13g2_fill_2 FILLER_32_71 ();
 sg13g2_decap_4 FILLER_32_83 ();
 sg13g2_fill_2 FILLER_32_87 ();
 sg13g2_fill_2 FILLER_32_116 ();
 sg13g2_decap_8 FILLER_32_149 ();
 sg13g2_decap_8 FILLER_32_156 ();
 sg13g2_fill_2 FILLER_32_163 ();
 sg13g2_fill_1 FILLER_32_165 ();
 sg13g2_fill_1 FILLER_32_202 ();
 sg13g2_decap_8 FILLER_32_236 ();
 sg13g2_decap_8 FILLER_32_243 ();
 sg13g2_decap_4 FILLER_32_250 ();
 sg13g2_fill_2 FILLER_32_254 ();
 sg13g2_fill_2 FILLER_32_269 ();
 sg13g2_fill_1 FILLER_32_271 ();
 sg13g2_fill_2 FILLER_32_280 ();
 sg13g2_fill_2 FILLER_32_329 ();
 sg13g2_fill_1 FILLER_32_331 ();
 sg13g2_decap_4 FILLER_32_344 ();
 sg13g2_fill_1 FILLER_32_399 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_7 ();
 sg13g2_fill_2 FILLER_33_11 ();
 sg13g2_fill_2 FILLER_33_53 ();
 sg13g2_fill_1 FILLER_33_55 ();
 sg13g2_fill_1 FILLER_33_105 ();
 sg13g2_fill_1 FILLER_33_115 ();
 sg13g2_decap_8 FILLER_33_150 ();
 sg13g2_decap_4 FILLER_33_157 ();
 sg13g2_fill_1 FILLER_33_165 ();
 sg13g2_fill_2 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_236 ();
 sg13g2_decap_4 FILLER_33_247 ();
 sg13g2_fill_1 FILLER_33_251 ();
 sg13g2_fill_1 FILLER_33_284 ();
 sg13g2_decap_8 FILLER_33_312 ();
 sg13g2_decap_8 FILLER_33_319 ();
 sg13g2_fill_2 FILLER_33_331 ();
 sg13g2_fill_2 FILLER_33_343 ();
 sg13g2_fill_2 FILLER_33_351 ();
 sg13g2_fill_1 FILLER_33_376 ();
 sg13g2_fill_2 FILLER_33_385 ();
 sg13g2_fill_1 FILLER_33_387 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_4 FILLER_34_75 ();
 sg13g2_fill_1 FILLER_34_118 ();
 sg13g2_fill_1 FILLER_34_138 ();
 sg13g2_fill_1 FILLER_34_192 ();
 sg13g2_fill_2 FILLER_34_198 ();
 sg13g2_fill_1 FILLER_34_200 ();
 sg13g2_fill_1 FILLER_34_205 ();
 sg13g2_fill_1 FILLER_34_210 ();
 sg13g2_decap_4 FILLER_34_229 ();
 sg13g2_fill_2 FILLER_34_233 ();
 sg13g2_fill_2 FILLER_34_244 ();
 sg13g2_fill_1 FILLER_34_246 ();
 sg13g2_fill_1 FILLER_34_283 ();
 sg13g2_fill_2 FILLER_34_306 ();
 sg13g2_fill_1 FILLER_34_308 ();
 sg13g2_decap_4 FILLER_34_333 ();
 sg13g2_fill_1 FILLER_34_337 ();
 sg13g2_decap_4 FILLER_34_372 ();
 sg13g2_fill_1 FILLER_34_376 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_14 ();
 sg13g2_fill_1 FILLER_35_16 ();
 sg13g2_decap_4 FILLER_35_57 ();
 sg13g2_decap_8 FILLER_35_115 ();
 sg13g2_decap_4 FILLER_35_122 ();
 sg13g2_fill_2 FILLER_35_126 ();
 sg13g2_fill_2 FILLER_35_145 ();
 sg13g2_fill_1 FILLER_35_191 ();
 sg13g2_fill_2 FILLER_35_243 ();
 sg13g2_fill_2 FILLER_35_276 ();
 sg13g2_fill_2 FILLER_35_296 ();
 sg13g2_fill_1 FILLER_35_298 ();
 sg13g2_fill_2 FILLER_35_312 ();
 sg13g2_fill_2 FILLER_35_340 ();
 sg13g2_decap_4 FILLER_35_357 ();
 sg13g2_fill_1 FILLER_35_361 ();
 sg13g2_fill_2 FILLER_35_376 ();
 sg13g2_fill_1 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_401 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_fill_1 FILLER_36_50 ();
 sg13g2_fill_1 FILLER_36_64 ();
 sg13g2_decap_8 FILLER_36_123 ();
 sg13g2_fill_2 FILLER_36_130 ();
 sg13g2_fill_1 FILLER_36_132 ();
 sg13g2_fill_2 FILLER_36_160 ();
 sg13g2_fill_2 FILLER_36_171 ();
 sg13g2_fill_2 FILLER_36_178 ();
 sg13g2_decap_4 FILLER_36_184 ();
 sg13g2_fill_1 FILLER_36_188 ();
 sg13g2_fill_1 FILLER_36_216 ();
 sg13g2_fill_2 FILLER_36_226 ();
 sg13g2_fill_2 FILLER_36_282 ();
 sg13g2_fill_2 FILLER_36_338 ();
 sg13g2_fill_1 FILLER_36_340 ();
 sg13g2_decap_4 FILLER_36_404 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_4 FILLER_37_21 ();
 sg13g2_fill_1 FILLER_37_25 ();
 sg13g2_decap_8 FILLER_37_30 ();
 sg13g2_fill_2 FILLER_37_37 ();
 sg13g2_fill_1 FILLER_37_66 ();
 sg13g2_fill_1 FILLER_37_116 ();
 sg13g2_fill_1 FILLER_37_164 ();
 sg13g2_fill_1 FILLER_37_192 ();
 sg13g2_fill_2 FILLER_37_322 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_4 FILLER_38_28 ();
 sg13g2_fill_1 FILLER_38_32 ();
 sg13g2_fill_2 FILLER_38_50 ();
 sg13g2_fill_1 FILLER_38_52 ();
 sg13g2_fill_1 FILLER_38_100 ();
 sg13g2_fill_1 FILLER_38_110 ();
 sg13g2_fill_2 FILLER_38_184 ();
 sg13g2_fill_1 FILLER_38_186 ();
 sg13g2_decap_4 FILLER_38_196 ();
 sg13g2_fill_2 FILLER_38_200 ();
 sg13g2_fill_1 FILLER_38_206 ();
 sg13g2_decap_8 FILLER_38_211 ();
 sg13g2_decap_8 FILLER_38_218 ();
 sg13g2_decap_8 FILLER_38_225 ();
 sg13g2_fill_1 FILLER_38_232 ();
 sg13g2_fill_2 FILLER_38_237 ();
 sg13g2_fill_1 FILLER_38_274 ();
 sg13g2_fill_1 FILLER_38_292 ();
 sg13g2_fill_2 FILLER_38_306 ();
 sg13g2_fill_1 FILLER_38_308 ();
 sg13g2_fill_2 FILLER_38_350 ();
 sg13g2_decap_4 FILLER_38_356 ();
 sg13g2_decap_4 FILLER_38_364 ();
 sg13g2_decap_4 FILLER_38_372 ();
 sg13g2_fill_1 FILLER_38_384 ();
 sg13g2_decap_8 FILLER_38_394 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net14;
 assign uio_oe[1] = net15;
 assign uio_oe[2] = net16;
 assign uio_oe[3] = net17;
 assign uio_oe[4] = net18;
 assign uio_oe[5] = net19;
 assign uio_oe[6] = net20;
 assign uio_oe[7] = net21;
 assign uio_out[0] = net22;
 assign uio_out[1] = net23;
 assign uio_out[2] = net24;
 assign uio_out[3] = net25;
 assign uio_out[4] = net26;
 assign uio_out[5] = net27;
 assign uio_out[6] = net28;
 assign uio_out[7] = net29;
endmodule
